module basic_750_5000_1000_10_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_409,In_730);
and U1 (N_1,In_370,In_378);
xnor U2 (N_2,In_293,In_694);
or U3 (N_3,In_718,In_736);
xor U4 (N_4,In_534,In_123);
or U5 (N_5,In_400,In_383);
xor U6 (N_6,In_650,In_433);
nand U7 (N_7,In_360,In_125);
nor U8 (N_8,In_604,In_605);
and U9 (N_9,In_476,In_46);
and U10 (N_10,In_707,In_492);
and U11 (N_11,In_682,In_175);
xnor U12 (N_12,In_167,In_714);
nand U13 (N_13,In_516,In_171);
or U14 (N_14,In_111,In_273);
or U15 (N_15,In_284,In_2);
nand U16 (N_16,In_681,In_633);
or U17 (N_17,In_398,In_311);
nor U18 (N_18,In_7,In_572);
or U19 (N_19,In_238,In_532);
and U20 (N_20,In_13,In_388);
xor U21 (N_21,In_723,In_50);
or U22 (N_22,In_313,In_287);
or U23 (N_23,In_137,In_524);
xnor U24 (N_24,In_598,In_72);
or U25 (N_25,In_402,In_57);
and U26 (N_26,In_157,In_468);
xnor U27 (N_27,In_322,In_429);
and U28 (N_28,In_419,In_478);
xor U29 (N_29,In_336,In_744);
nand U30 (N_30,In_65,In_526);
and U31 (N_31,In_37,In_455);
and U32 (N_32,In_298,In_415);
nand U33 (N_33,In_477,In_69);
nand U34 (N_34,In_216,In_579);
xnor U35 (N_35,In_466,In_458);
xor U36 (N_36,In_99,In_249);
or U37 (N_37,In_363,In_326);
xnor U38 (N_38,In_106,In_571);
or U39 (N_39,In_735,In_602);
nand U40 (N_40,In_306,In_183);
and U41 (N_41,In_303,In_49);
xnor U42 (N_42,In_554,In_747);
or U43 (N_43,In_725,In_422);
and U44 (N_44,In_709,In_275);
xnor U45 (N_45,In_342,In_295);
or U46 (N_46,In_577,In_635);
or U47 (N_47,In_401,In_717);
and U48 (N_48,In_653,In_426);
xor U49 (N_49,In_348,In_404);
and U50 (N_50,In_496,In_277);
nand U51 (N_51,In_460,In_300);
xnor U52 (N_52,In_209,In_701);
nand U53 (N_53,In_439,In_634);
nor U54 (N_54,In_552,In_228);
nor U55 (N_55,In_290,In_715);
nor U56 (N_56,In_237,In_555);
and U57 (N_57,In_217,In_90);
nor U58 (N_58,In_620,In_66);
or U59 (N_59,In_39,In_28);
nor U60 (N_60,In_365,In_456);
xnor U61 (N_61,In_230,In_465);
nor U62 (N_62,In_140,In_549);
xor U63 (N_63,In_188,In_358);
nor U64 (N_64,In_589,In_133);
and U65 (N_65,In_254,In_142);
and U66 (N_66,In_655,In_722);
nand U67 (N_67,In_193,In_145);
xor U68 (N_68,In_22,In_472);
xor U69 (N_69,In_127,In_522);
xnor U70 (N_70,In_27,In_412);
and U71 (N_71,In_76,In_489);
nor U72 (N_72,In_606,In_220);
and U73 (N_73,In_566,In_474);
nand U74 (N_74,In_252,In_109);
xnor U75 (N_75,In_518,In_340);
nor U76 (N_76,In_712,In_420);
nand U77 (N_77,In_73,In_379);
nor U78 (N_78,In_449,In_459);
xnor U79 (N_79,In_246,In_481);
and U80 (N_80,In_189,In_208);
or U81 (N_81,In_366,In_55);
nor U82 (N_82,In_721,In_450);
nand U83 (N_83,In_148,In_622);
nor U84 (N_84,In_685,In_235);
or U85 (N_85,In_704,In_291);
nor U86 (N_86,In_45,In_67);
xnor U87 (N_87,In_505,In_130);
and U88 (N_88,In_194,In_461);
nor U89 (N_89,In_386,In_615);
nor U90 (N_90,In_32,In_62);
and U91 (N_91,In_218,In_475);
nand U92 (N_92,In_574,In_202);
nand U93 (N_93,In_488,In_191);
xnor U94 (N_94,In_393,In_104);
nand U95 (N_95,In_616,In_211);
and U96 (N_96,In_312,In_21);
nor U97 (N_97,In_196,In_173);
xor U98 (N_98,In_150,In_138);
and U99 (N_99,In_699,In_100);
and U100 (N_100,In_234,In_700);
nor U101 (N_101,In_91,In_541);
nand U102 (N_102,In_101,In_158);
and U103 (N_103,In_647,In_502);
or U104 (N_104,In_517,In_660);
xor U105 (N_105,In_705,In_212);
nor U106 (N_106,In_159,In_227);
nand U107 (N_107,In_656,In_676);
or U108 (N_108,In_359,In_551);
nand U109 (N_109,In_165,In_247);
nor U110 (N_110,In_546,In_223);
nor U111 (N_111,In_24,In_19);
nor U112 (N_112,In_177,In_338);
or U113 (N_113,In_529,In_179);
xor U114 (N_114,In_29,In_713);
xor U115 (N_115,In_600,In_396);
nor U116 (N_116,In_25,In_328);
xor U117 (N_117,In_564,In_144);
nor U118 (N_118,In_20,In_527);
nand U119 (N_119,In_71,In_623);
and U120 (N_120,In_282,In_486);
nor U121 (N_121,In_151,In_64);
and U122 (N_122,In_498,In_637);
xnor U123 (N_123,In_156,In_431);
nor U124 (N_124,In_662,In_116);
nand U125 (N_125,In_178,In_397);
nand U126 (N_126,In_658,In_557);
or U127 (N_127,In_181,In_703);
and U128 (N_128,In_163,In_274);
or U129 (N_129,In_501,In_248);
nand U130 (N_130,In_110,In_60);
nand U131 (N_131,In_40,In_535);
and U132 (N_132,In_688,In_573);
or U133 (N_133,In_103,In_129);
nand U134 (N_134,In_14,In_443);
xor U135 (N_135,In_683,In_446);
xnor U136 (N_136,In_418,In_464);
nand U137 (N_137,In_687,In_95);
xor U138 (N_138,In_444,In_543);
or U139 (N_139,In_737,In_176);
xnor U140 (N_140,In_327,In_644);
xnor U141 (N_141,In_480,In_425);
nor U142 (N_142,In_441,In_599);
and U143 (N_143,In_430,In_152);
xnor U144 (N_144,In_266,In_558);
nor U145 (N_145,In_684,In_270);
or U146 (N_146,In_587,In_169);
or U147 (N_147,In_671,In_48);
or U148 (N_148,In_595,In_649);
xor U149 (N_149,In_533,In_413);
xnor U150 (N_150,In_190,In_53);
and U151 (N_151,In_584,In_262);
or U152 (N_152,In_79,In_531);
or U153 (N_153,In_520,In_41);
or U154 (N_154,In_4,In_463);
or U155 (N_155,In_626,In_315);
and U156 (N_156,In_343,In_453);
xor U157 (N_157,In_411,In_436);
and U158 (N_158,In_93,In_618);
xnor U159 (N_159,In_582,In_642);
nor U160 (N_160,In_207,In_745);
xnor U161 (N_161,In_500,In_585);
or U162 (N_162,In_628,In_83);
nor U163 (N_163,In_344,In_136);
nand U164 (N_164,In_357,In_204);
nand U165 (N_165,In_74,In_353);
or U166 (N_166,In_428,In_332);
and U167 (N_167,In_612,In_345);
and U168 (N_168,In_296,In_42);
nand U169 (N_169,In_105,In_294);
or U170 (N_170,In_259,In_567);
xnor U171 (N_171,In_485,In_180);
and U172 (N_172,In_427,In_673);
xnor U173 (N_173,In_155,In_18);
and U174 (N_174,In_253,In_371);
and U175 (N_175,In_319,In_504);
nand U176 (N_176,In_115,In_738);
and U177 (N_177,In_467,In_352);
nand U178 (N_178,In_447,In_497);
or U179 (N_179,In_668,In_696);
nor U180 (N_180,In_562,In_361);
xnor U181 (N_181,In_490,In_525);
or U182 (N_182,In_643,In_16);
and U183 (N_183,In_569,In_263);
and U184 (N_184,In_229,In_280);
nor U185 (N_185,In_384,In_128);
xnor U186 (N_186,In_203,In_354);
nand U187 (N_187,In_61,In_3);
nand U188 (N_188,In_575,In_337);
xnor U189 (N_189,In_614,In_385);
nor U190 (N_190,In_310,In_82);
xnor U191 (N_191,In_545,In_166);
xnor U192 (N_192,In_454,In_30);
nand U193 (N_193,In_667,In_629);
and U194 (N_194,In_749,In_596);
or U195 (N_195,In_31,In_33);
xor U196 (N_196,In_367,In_731);
nand U197 (N_197,In_182,In_267);
or U198 (N_198,In_278,In_56);
or U199 (N_199,In_670,In_364);
nor U200 (N_200,In_511,In_561);
and U201 (N_201,In_382,In_513);
and U202 (N_202,In_675,In_448);
nor U203 (N_203,In_139,In_36);
nand U204 (N_204,In_728,In_611);
and U205 (N_205,In_631,In_603);
nor U206 (N_206,In_452,In_222);
xnor U207 (N_207,In_576,In_677);
nor U208 (N_208,In_669,In_484);
xor U209 (N_209,In_686,In_88);
xor U210 (N_210,In_679,In_568);
nand U211 (N_211,In_399,In_205);
or U212 (N_212,In_350,In_421);
nor U213 (N_213,In_122,In_372);
or U214 (N_214,In_617,In_297);
xor U215 (N_215,In_395,In_434);
nand U216 (N_216,In_424,In_339);
xor U217 (N_217,In_563,In_355);
nand U218 (N_218,In_135,In_210);
nor U219 (N_219,In_632,In_307);
nor U220 (N_220,In_506,In_323);
nor U221 (N_221,In_609,In_610);
nand U222 (N_222,In_578,In_652);
nor U223 (N_223,In_646,In_11);
or U224 (N_224,In_732,In_215);
and U225 (N_225,In_519,In_523);
or U226 (N_226,In_59,In_70);
xnor U227 (N_227,In_321,In_377);
or U228 (N_228,In_316,In_119);
or U229 (N_229,In_271,In_292);
nor U230 (N_230,In_34,In_301);
and U231 (N_231,In_680,In_530);
and U232 (N_232,In_86,In_624);
and U233 (N_233,In_499,In_143);
nor U234 (N_234,In_43,In_268);
xor U235 (N_235,In_445,In_538);
xnor U236 (N_236,In_325,In_107);
xnor U237 (N_237,In_341,In_236);
nand U238 (N_238,In_547,In_743);
xnor U239 (N_239,In_12,In_423);
or U240 (N_240,In_470,In_394);
xor U241 (N_241,In_416,In_233);
nand U242 (N_242,In_318,In_724);
and U243 (N_243,In_317,In_432);
or U244 (N_244,In_225,In_588);
and U245 (N_245,In_410,In_601);
xor U246 (N_246,In_241,In_279);
nand U247 (N_247,In_373,In_548);
nor U248 (N_248,In_693,In_716);
xnor U249 (N_249,In_26,In_35);
xor U250 (N_250,In_58,In_94);
nor U251 (N_251,In_392,In_556);
or U252 (N_252,In_539,In_471);
and U253 (N_253,In_47,In_374);
nand U254 (N_254,In_147,In_17);
xnor U255 (N_255,In_195,In_164);
or U256 (N_256,In_442,In_134);
nor U257 (N_257,In_92,In_6);
nand U258 (N_258,In_232,In_243);
xnor U259 (N_259,In_691,In_437);
xor U260 (N_260,In_621,In_469);
nor U261 (N_261,In_78,In_308);
or U262 (N_262,In_114,In_174);
nand U263 (N_263,In_487,In_741);
xnor U264 (N_264,In_702,In_324);
nor U265 (N_265,In_224,In_665);
or U266 (N_266,In_406,In_329);
or U267 (N_267,In_560,In_514);
or U268 (N_268,In_356,In_347);
nor U269 (N_269,In_113,In_414);
nor U270 (N_270,In_651,In_544);
or U271 (N_271,In_89,In_407);
xnor U272 (N_272,In_638,In_168);
xor U273 (N_273,In_659,In_44);
nor U274 (N_274,In_240,In_245);
xor U275 (N_275,In_8,In_132);
or U276 (N_276,In_746,In_75);
xnor U277 (N_277,In_462,In_51);
nor U278 (N_278,In_0,In_457);
or U279 (N_279,In_528,In_663);
xnor U280 (N_280,In_23,In_593);
nand U281 (N_281,In_542,In_664);
or U282 (N_282,In_479,In_199);
and U283 (N_283,In_625,In_742);
xor U284 (N_284,In_666,In_242);
xnor U285 (N_285,In_473,In_405);
nand U286 (N_286,In_162,In_440);
nor U287 (N_287,In_200,In_314);
or U288 (N_288,In_692,In_510);
or U289 (N_289,In_221,In_260);
nand U290 (N_290,In_697,In_264);
xnor U291 (N_291,In_661,In_483);
xor U292 (N_292,In_187,In_640);
nor U293 (N_293,In_184,In_257);
and U294 (N_294,In_244,In_630);
and U295 (N_295,In_503,In_739);
nor U296 (N_296,In_198,In_251);
or U297 (N_297,In_52,In_206);
xor U298 (N_298,In_581,In_491);
xnor U299 (N_299,In_346,In_559);
and U300 (N_300,In_607,In_594);
nor U301 (N_301,In_154,In_387);
and U302 (N_302,In_495,In_10);
and U303 (N_303,In_320,In_403);
nand U304 (N_304,In_38,In_261);
or U305 (N_305,In_597,In_408);
nor U306 (N_306,In_126,In_170);
xor U307 (N_307,In_108,In_289);
nor U308 (N_308,In_592,In_87);
xor U309 (N_309,In_550,In_708);
nor U310 (N_310,In_63,In_239);
nand U311 (N_311,In_331,In_368);
xnor U312 (N_312,In_390,In_719);
nand U313 (N_313,In_580,In_54);
and U314 (N_314,In_77,In_231);
xor U315 (N_315,In_515,In_706);
xor U316 (N_316,In_186,In_98);
or U317 (N_317,In_281,In_309);
or U318 (N_318,In_219,In_639);
xnor U319 (N_319,In_507,In_96);
and U320 (N_320,In_214,In_258);
nand U321 (N_321,In_654,In_508);
and U322 (N_322,In_351,In_613);
or U323 (N_323,In_438,In_540);
and U324 (N_324,In_657,In_451);
xor U325 (N_325,In_226,In_674);
xor U326 (N_326,In_185,In_381);
and U327 (N_327,In_120,In_727);
nor U328 (N_328,In_286,In_678);
and U329 (N_329,In_591,In_192);
nand U330 (N_330,In_636,In_689);
or U331 (N_331,In_376,In_335);
xor U332 (N_332,In_362,In_161);
or U333 (N_333,In_349,In_80);
and U334 (N_334,In_118,In_153);
xor U335 (N_335,In_710,In_590);
nand U336 (N_336,In_698,In_330);
nand U337 (N_337,In_720,In_672);
nor U338 (N_338,In_389,In_81);
or U339 (N_339,In_250,In_9);
or U340 (N_340,In_112,In_146);
nor U341 (N_341,In_131,In_256);
xnor U342 (N_342,In_334,In_124);
nand U343 (N_343,In_302,In_197);
nand U344 (N_344,In_521,In_305);
and U345 (N_345,In_570,In_102);
nor U346 (N_346,In_512,In_97);
and U347 (N_347,In_333,In_272);
xnor U348 (N_348,In_748,In_375);
nand U349 (N_349,In_288,In_172);
nand U350 (N_350,In_304,In_494);
xor U351 (N_351,In_608,In_265);
xnor U352 (N_352,In_740,In_160);
nand U353 (N_353,In_68,In_417);
nor U354 (N_354,In_15,In_695);
or U355 (N_355,In_553,In_1);
nand U356 (N_356,In_269,In_141);
and U357 (N_357,In_729,In_149);
nor U358 (N_358,In_537,In_583);
nand U359 (N_359,In_117,In_627);
xor U360 (N_360,In_711,In_536);
nand U361 (N_361,In_213,In_299);
nor U362 (N_362,In_565,In_734);
xor U363 (N_363,In_726,In_5);
or U364 (N_364,In_586,In_121);
and U365 (N_365,In_201,In_255);
and U366 (N_366,In_482,In_733);
nand U367 (N_367,In_285,In_645);
nand U368 (N_368,In_84,In_648);
or U369 (N_369,In_380,In_641);
nand U370 (N_370,In_85,In_509);
or U371 (N_371,In_276,In_619);
nand U372 (N_372,In_690,In_391);
xnor U373 (N_373,In_283,In_369);
xnor U374 (N_374,In_493,In_435);
xnor U375 (N_375,In_527,In_687);
xor U376 (N_376,In_289,In_246);
or U377 (N_377,In_303,In_265);
or U378 (N_378,In_621,In_550);
and U379 (N_379,In_41,In_130);
xor U380 (N_380,In_128,In_553);
and U381 (N_381,In_221,In_52);
or U382 (N_382,In_374,In_473);
xor U383 (N_383,In_688,In_421);
and U384 (N_384,In_84,In_265);
or U385 (N_385,In_724,In_430);
xnor U386 (N_386,In_707,In_498);
nand U387 (N_387,In_613,In_244);
nor U388 (N_388,In_596,In_638);
nor U389 (N_389,In_644,In_126);
or U390 (N_390,In_138,In_620);
nor U391 (N_391,In_564,In_323);
xor U392 (N_392,In_434,In_34);
nor U393 (N_393,In_737,In_524);
and U394 (N_394,In_461,In_230);
and U395 (N_395,In_424,In_243);
and U396 (N_396,In_85,In_21);
nor U397 (N_397,In_546,In_398);
nor U398 (N_398,In_423,In_19);
or U399 (N_399,In_504,In_218);
nand U400 (N_400,In_464,In_710);
and U401 (N_401,In_575,In_396);
nor U402 (N_402,In_168,In_103);
nand U403 (N_403,In_373,In_621);
nand U404 (N_404,In_552,In_199);
nand U405 (N_405,In_162,In_234);
nand U406 (N_406,In_167,In_563);
and U407 (N_407,In_32,In_309);
or U408 (N_408,In_227,In_629);
xor U409 (N_409,In_289,In_476);
or U410 (N_410,In_339,In_703);
xor U411 (N_411,In_237,In_411);
or U412 (N_412,In_420,In_552);
nand U413 (N_413,In_428,In_164);
nand U414 (N_414,In_22,In_264);
nand U415 (N_415,In_211,In_437);
or U416 (N_416,In_159,In_333);
nor U417 (N_417,In_275,In_241);
xor U418 (N_418,In_416,In_346);
xnor U419 (N_419,In_29,In_393);
nor U420 (N_420,In_747,In_189);
or U421 (N_421,In_418,In_390);
or U422 (N_422,In_65,In_164);
nor U423 (N_423,In_585,In_52);
or U424 (N_424,In_251,In_39);
or U425 (N_425,In_202,In_302);
xnor U426 (N_426,In_134,In_504);
and U427 (N_427,In_253,In_714);
nand U428 (N_428,In_280,In_411);
xnor U429 (N_429,In_387,In_632);
nor U430 (N_430,In_475,In_344);
xnor U431 (N_431,In_709,In_579);
and U432 (N_432,In_577,In_701);
xnor U433 (N_433,In_105,In_107);
and U434 (N_434,In_401,In_535);
nand U435 (N_435,In_253,In_409);
nand U436 (N_436,In_525,In_609);
xnor U437 (N_437,In_236,In_369);
and U438 (N_438,In_56,In_474);
nor U439 (N_439,In_354,In_174);
nor U440 (N_440,In_78,In_18);
nor U441 (N_441,In_215,In_496);
or U442 (N_442,In_378,In_589);
nand U443 (N_443,In_178,In_555);
xor U444 (N_444,In_735,In_71);
nand U445 (N_445,In_57,In_410);
nor U446 (N_446,In_189,In_692);
nor U447 (N_447,In_631,In_418);
nand U448 (N_448,In_743,In_433);
nor U449 (N_449,In_651,In_373);
xor U450 (N_450,In_426,In_227);
nor U451 (N_451,In_644,In_232);
xnor U452 (N_452,In_385,In_144);
and U453 (N_453,In_95,In_629);
nand U454 (N_454,In_99,In_143);
and U455 (N_455,In_29,In_259);
nor U456 (N_456,In_575,In_193);
and U457 (N_457,In_340,In_180);
or U458 (N_458,In_418,In_495);
nand U459 (N_459,In_517,In_314);
and U460 (N_460,In_116,In_176);
nand U461 (N_461,In_674,In_622);
or U462 (N_462,In_364,In_214);
or U463 (N_463,In_402,In_613);
xor U464 (N_464,In_625,In_477);
xor U465 (N_465,In_715,In_257);
and U466 (N_466,In_35,In_132);
and U467 (N_467,In_292,In_158);
nor U468 (N_468,In_248,In_485);
xor U469 (N_469,In_473,In_650);
and U470 (N_470,In_80,In_680);
or U471 (N_471,In_232,In_695);
and U472 (N_472,In_412,In_668);
nor U473 (N_473,In_695,In_346);
or U474 (N_474,In_158,In_177);
and U475 (N_475,In_686,In_271);
xnor U476 (N_476,In_538,In_267);
and U477 (N_477,In_531,In_136);
xor U478 (N_478,In_437,In_387);
nor U479 (N_479,In_536,In_369);
xnor U480 (N_480,In_712,In_180);
xor U481 (N_481,In_501,In_418);
xnor U482 (N_482,In_441,In_14);
xor U483 (N_483,In_53,In_358);
xnor U484 (N_484,In_748,In_596);
nand U485 (N_485,In_397,In_707);
nor U486 (N_486,In_367,In_711);
nand U487 (N_487,In_88,In_520);
and U488 (N_488,In_506,In_528);
xor U489 (N_489,In_454,In_620);
nand U490 (N_490,In_591,In_339);
and U491 (N_491,In_507,In_625);
xor U492 (N_492,In_314,In_469);
nand U493 (N_493,In_405,In_337);
xor U494 (N_494,In_25,In_307);
xnor U495 (N_495,In_2,In_728);
or U496 (N_496,In_566,In_404);
nor U497 (N_497,In_306,In_676);
nand U498 (N_498,In_619,In_93);
nor U499 (N_499,In_678,In_504);
nor U500 (N_500,N_206,N_239);
or U501 (N_501,N_115,N_60);
xor U502 (N_502,N_54,N_492);
and U503 (N_503,N_138,N_495);
nor U504 (N_504,N_373,N_333);
nor U505 (N_505,N_277,N_378);
nor U506 (N_506,N_123,N_202);
nand U507 (N_507,N_6,N_235);
or U508 (N_508,N_321,N_433);
and U509 (N_509,N_361,N_29);
nor U510 (N_510,N_344,N_400);
and U511 (N_511,N_141,N_210);
and U512 (N_512,N_69,N_9);
or U513 (N_513,N_301,N_350);
and U514 (N_514,N_352,N_150);
nand U515 (N_515,N_47,N_313);
nor U516 (N_516,N_20,N_471);
and U517 (N_517,N_309,N_121);
xnor U518 (N_518,N_16,N_459);
nand U519 (N_519,N_230,N_367);
nand U520 (N_520,N_311,N_62);
and U521 (N_521,N_261,N_215);
xor U522 (N_522,N_448,N_70);
nand U523 (N_523,N_369,N_442);
nor U524 (N_524,N_385,N_273);
or U525 (N_525,N_95,N_186);
or U526 (N_526,N_165,N_351);
and U527 (N_527,N_94,N_209);
nor U528 (N_528,N_372,N_86);
nand U529 (N_529,N_270,N_197);
and U530 (N_530,N_79,N_424);
and U531 (N_531,N_478,N_458);
nor U532 (N_532,N_90,N_208);
or U533 (N_533,N_377,N_469);
nor U534 (N_534,N_101,N_49);
xnor U535 (N_535,N_304,N_320);
nand U536 (N_536,N_430,N_97);
nor U537 (N_537,N_59,N_189);
nand U538 (N_538,N_251,N_269);
xor U539 (N_539,N_272,N_256);
nand U540 (N_540,N_19,N_98);
and U541 (N_541,N_218,N_331);
nand U542 (N_542,N_399,N_162);
and U543 (N_543,N_125,N_499);
xnor U544 (N_544,N_45,N_63);
and U545 (N_545,N_220,N_418);
nor U546 (N_546,N_308,N_249);
nor U547 (N_547,N_420,N_444);
xnor U548 (N_548,N_314,N_435);
or U549 (N_549,N_130,N_196);
nand U550 (N_550,N_395,N_116);
or U551 (N_551,N_490,N_384);
and U552 (N_552,N_383,N_267);
or U553 (N_553,N_477,N_419);
or U554 (N_554,N_61,N_149);
xnor U555 (N_555,N_494,N_167);
and U556 (N_556,N_353,N_366);
nand U557 (N_557,N_410,N_257);
nand U558 (N_558,N_135,N_255);
nor U559 (N_559,N_204,N_286);
nor U560 (N_560,N_24,N_36);
nor U561 (N_561,N_40,N_71);
nor U562 (N_562,N_145,N_75);
xnor U563 (N_563,N_429,N_114);
or U564 (N_564,N_339,N_466);
nand U565 (N_565,N_200,N_474);
and U566 (N_566,N_169,N_451);
nand U567 (N_567,N_342,N_405);
or U568 (N_568,N_391,N_96);
xor U569 (N_569,N_401,N_393);
or U570 (N_570,N_51,N_462);
xor U571 (N_571,N_346,N_276);
xor U572 (N_572,N_334,N_179);
and U573 (N_573,N_232,N_248);
and U574 (N_574,N_148,N_456);
or U575 (N_575,N_496,N_28);
nand U576 (N_576,N_485,N_11);
xnor U577 (N_577,N_214,N_13);
xor U578 (N_578,N_404,N_275);
xnor U579 (N_579,N_132,N_285);
or U580 (N_580,N_422,N_25);
nor U581 (N_581,N_359,N_180);
or U582 (N_582,N_32,N_128);
and U583 (N_583,N_475,N_39);
or U584 (N_584,N_472,N_241);
nand U585 (N_585,N_408,N_406);
nor U586 (N_586,N_183,N_152);
xnor U587 (N_587,N_362,N_139);
and U588 (N_588,N_182,N_274);
and U589 (N_589,N_368,N_154);
or U590 (N_590,N_280,N_319);
or U591 (N_591,N_349,N_355);
and U592 (N_592,N_85,N_497);
and U593 (N_593,N_74,N_425);
nor U594 (N_594,N_7,N_175);
or U595 (N_595,N_279,N_194);
xor U596 (N_596,N_438,N_450);
xnor U597 (N_597,N_21,N_443);
or U598 (N_598,N_498,N_452);
xor U599 (N_599,N_306,N_168);
nor U600 (N_600,N_35,N_467);
and U601 (N_601,N_161,N_268);
nor U602 (N_602,N_108,N_463);
xor U603 (N_603,N_282,N_465);
and U604 (N_604,N_348,N_188);
and U605 (N_605,N_445,N_44);
or U606 (N_606,N_106,N_177);
nand U607 (N_607,N_482,N_436);
or U608 (N_608,N_126,N_300);
nand U609 (N_609,N_104,N_253);
and U610 (N_610,N_338,N_297);
nand U611 (N_611,N_50,N_439);
and U612 (N_612,N_153,N_335);
xor U613 (N_613,N_192,N_224);
xnor U614 (N_614,N_302,N_244);
nor U615 (N_615,N_129,N_22);
xor U616 (N_616,N_64,N_226);
xor U617 (N_617,N_441,N_66);
nor U618 (N_618,N_387,N_17);
nand U619 (N_619,N_187,N_65);
and U620 (N_620,N_146,N_262);
nor U621 (N_621,N_227,N_172);
xor U622 (N_622,N_489,N_379);
xnor U623 (N_623,N_155,N_281);
and U624 (N_624,N_403,N_158);
nand U625 (N_625,N_18,N_437);
and U626 (N_626,N_263,N_205);
or U627 (N_627,N_303,N_449);
and U628 (N_628,N_53,N_317);
and U629 (N_629,N_229,N_231);
and U630 (N_630,N_105,N_330);
and U631 (N_631,N_112,N_102);
nand U632 (N_632,N_414,N_91);
or U633 (N_633,N_398,N_250);
xor U634 (N_634,N_191,N_341);
and U635 (N_635,N_143,N_72);
xnor U636 (N_636,N_142,N_212);
nand U637 (N_637,N_487,N_382);
and U638 (N_638,N_325,N_416);
nand U639 (N_639,N_431,N_233);
xor U640 (N_640,N_120,N_78);
and U641 (N_641,N_423,N_15);
xnor U642 (N_642,N_271,N_396);
xor U643 (N_643,N_31,N_415);
and U644 (N_644,N_181,N_493);
nor U645 (N_645,N_390,N_26);
nor U646 (N_646,N_80,N_296);
or U647 (N_647,N_329,N_266);
or U648 (N_648,N_340,N_119);
xor U649 (N_649,N_41,N_455);
nand U650 (N_650,N_163,N_225);
xor U651 (N_651,N_38,N_473);
nand U652 (N_652,N_176,N_293);
nand U653 (N_653,N_190,N_460);
nand U654 (N_654,N_221,N_323);
nor U655 (N_655,N_245,N_413);
and U656 (N_656,N_371,N_43);
and U657 (N_657,N_488,N_417);
or U658 (N_658,N_357,N_312);
nand U659 (N_659,N_37,N_476);
nand U660 (N_660,N_3,N_411);
xnor U661 (N_661,N_203,N_328);
and U662 (N_662,N_107,N_77);
nor U663 (N_663,N_73,N_111);
or U664 (N_664,N_428,N_228);
nor U665 (N_665,N_461,N_122);
xor U666 (N_666,N_364,N_4);
xnor U667 (N_667,N_134,N_82);
or U668 (N_668,N_185,N_491);
nor U669 (N_669,N_117,N_289);
nor U670 (N_670,N_389,N_58);
nand U671 (N_671,N_219,N_386);
and U672 (N_672,N_365,N_110);
and U673 (N_673,N_480,N_81);
xor U674 (N_674,N_57,N_93);
nor U675 (N_675,N_322,N_332);
nand U676 (N_676,N_464,N_345);
xor U677 (N_677,N_216,N_88);
and U678 (N_678,N_374,N_343);
nand U679 (N_679,N_380,N_124);
nand U680 (N_680,N_113,N_222);
and U681 (N_681,N_326,N_242);
and U682 (N_682,N_201,N_42);
nor U683 (N_683,N_375,N_174);
nand U684 (N_684,N_193,N_136);
xnor U685 (N_685,N_170,N_427);
xor U686 (N_686,N_184,N_237);
xor U687 (N_687,N_432,N_207);
nand U688 (N_688,N_178,N_337);
xnor U689 (N_689,N_376,N_87);
nand U690 (N_690,N_409,N_223);
and U691 (N_691,N_265,N_100);
or U692 (N_692,N_315,N_48);
nor U693 (N_693,N_260,N_434);
or U694 (N_694,N_246,N_2);
or U695 (N_695,N_5,N_447);
or U696 (N_696,N_12,N_283);
xor U697 (N_697,N_195,N_23);
nor U698 (N_698,N_254,N_173);
and U699 (N_699,N_10,N_347);
or U700 (N_700,N_316,N_55);
and U701 (N_701,N_33,N_358);
nor U702 (N_702,N_133,N_481);
nor U703 (N_703,N_213,N_440);
nand U704 (N_704,N_147,N_336);
nor U705 (N_705,N_307,N_166);
or U706 (N_706,N_144,N_137);
and U707 (N_707,N_360,N_295);
xor U708 (N_708,N_247,N_402);
and U709 (N_709,N_483,N_164);
nand U710 (N_710,N_67,N_127);
and U711 (N_711,N_83,N_397);
xnor U712 (N_712,N_156,N_486);
nand U713 (N_713,N_240,N_363);
or U714 (N_714,N_292,N_171);
xor U715 (N_715,N_34,N_92);
nand U716 (N_716,N_421,N_252);
and U717 (N_717,N_457,N_27);
nand U718 (N_718,N_198,N_259);
nand U719 (N_719,N_278,N_211);
xor U720 (N_720,N_118,N_287);
and U721 (N_721,N_103,N_264);
xnor U722 (N_722,N_89,N_1);
nor U723 (N_723,N_236,N_46);
nor U724 (N_724,N_238,N_84);
nand U725 (N_725,N_56,N_318);
nand U726 (N_726,N_327,N_356);
or U727 (N_727,N_76,N_140);
nand U728 (N_728,N_68,N_426);
or U729 (N_729,N_131,N_381);
nand U730 (N_730,N_199,N_52);
nand U731 (N_731,N_324,N_109);
xnor U732 (N_732,N_234,N_392);
and U733 (N_733,N_217,N_354);
xor U734 (N_734,N_151,N_0);
or U735 (N_735,N_299,N_291);
and U736 (N_736,N_446,N_468);
and U737 (N_737,N_454,N_258);
xor U738 (N_738,N_30,N_8);
and U739 (N_739,N_484,N_290);
and U740 (N_740,N_388,N_453);
and U741 (N_741,N_288,N_284);
xor U742 (N_742,N_394,N_310);
or U743 (N_743,N_99,N_305);
nand U744 (N_744,N_243,N_157);
nand U745 (N_745,N_407,N_160);
and U746 (N_746,N_298,N_370);
nor U747 (N_747,N_294,N_159);
nand U748 (N_748,N_470,N_479);
and U749 (N_749,N_412,N_14);
and U750 (N_750,N_340,N_352);
and U751 (N_751,N_132,N_145);
nand U752 (N_752,N_171,N_289);
xor U753 (N_753,N_106,N_480);
xor U754 (N_754,N_448,N_64);
nor U755 (N_755,N_201,N_254);
or U756 (N_756,N_196,N_169);
or U757 (N_757,N_106,N_284);
and U758 (N_758,N_134,N_387);
or U759 (N_759,N_445,N_219);
nor U760 (N_760,N_291,N_429);
or U761 (N_761,N_251,N_205);
nand U762 (N_762,N_183,N_250);
nor U763 (N_763,N_271,N_352);
xnor U764 (N_764,N_123,N_326);
and U765 (N_765,N_498,N_404);
nor U766 (N_766,N_250,N_408);
or U767 (N_767,N_119,N_124);
and U768 (N_768,N_80,N_465);
xor U769 (N_769,N_12,N_132);
xnor U770 (N_770,N_329,N_291);
nand U771 (N_771,N_386,N_81);
nand U772 (N_772,N_270,N_431);
or U773 (N_773,N_239,N_385);
or U774 (N_774,N_181,N_48);
nand U775 (N_775,N_290,N_337);
or U776 (N_776,N_271,N_380);
xor U777 (N_777,N_308,N_208);
or U778 (N_778,N_100,N_378);
or U779 (N_779,N_233,N_123);
nand U780 (N_780,N_337,N_210);
xor U781 (N_781,N_363,N_278);
xor U782 (N_782,N_260,N_121);
xnor U783 (N_783,N_69,N_176);
xor U784 (N_784,N_487,N_27);
and U785 (N_785,N_80,N_320);
xor U786 (N_786,N_56,N_496);
or U787 (N_787,N_167,N_203);
or U788 (N_788,N_246,N_385);
or U789 (N_789,N_462,N_168);
nand U790 (N_790,N_327,N_55);
xor U791 (N_791,N_231,N_147);
or U792 (N_792,N_29,N_339);
nand U793 (N_793,N_88,N_191);
nand U794 (N_794,N_495,N_3);
and U795 (N_795,N_100,N_386);
or U796 (N_796,N_121,N_314);
and U797 (N_797,N_228,N_456);
and U798 (N_798,N_132,N_288);
and U799 (N_799,N_359,N_107);
nand U800 (N_800,N_432,N_339);
and U801 (N_801,N_471,N_211);
nor U802 (N_802,N_164,N_170);
xnor U803 (N_803,N_158,N_55);
and U804 (N_804,N_196,N_427);
nor U805 (N_805,N_273,N_51);
xnor U806 (N_806,N_337,N_56);
and U807 (N_807,N_409,N_49);
nor U808 (N_808,N_94,N_21);
or U809 (N_809,N_117,N_132);
nand U810 (N_810,N_183,N_445);
nand U811 (N_811,N_295,N_142);
nand U812 (N_812,N_264,N_365);
or U813 (N_813,N_265,N_331);
nor U814 (N_814,N_407,N_184);
xnor U815 (N_815,N_105,N_181);
nor U816 (N_816,N_261,N_486);
or U817 (N_817,N_134,N_206);
nor U818 (N_818,N_441,N_65);
or U819 (N_819,N_286,N_81);
or U820 (N_820,N_101,N_351);
and U821 (N_821,N_478,N_237);
nand U822 (N_822,N_362,N_425);
or U823 (N_823,N_494,N_96);
nor U824 (N_824,N_25,N_115);
nand U825 (N_825,N_229,N_298);
nor U826 (N_826,N_255,N_305);
and U827 (N_827,N_42,N_178);
or U828 (N_828,N_193,N_6);
xnor U829 (N_829,N_163,N_444);
and U830 (N_830,N_64,N_263);
xor U831 (N_831,N_472,N_66);
nor U832 (N_832,N_291,N_460);
nor U833 (N_833,N_160,N_482);
nand U834 (N_834,N_72,N_278);
nand U835 (N_835,N_242,N_345);
xnor U836 (N_836,N_480,N_173);
or U837 (N_837,N_454,N_131);
or U838 (N_838,N_147,N_109);
and U839 (N_839,N_465,N_238);
nand U840 (N_840,N_322,N_209);
or U841 (N_841,N_9,N_21);
nor U842 (N_842,N_14,N_46);
xnor U843 (N_843,N_283,N_188);
nor U844 (N_844,N_472,N_190);
nor U845 (N_845,N_20,N_407);
or U846 (N_846,N_366,N_347);
or U847 (N_847,N_195,N_290);
and U848 (N_848,N_382,N_163);
xnor U849 (N_849,N_141,N_153);
xor U850 (N_850,N_54,N_432);
nand U851 (N_851,N_17,N_6);
nor U852 (N_852,N_356,N_102);
and U853 (N_853,N_397,N_98);
and U854 (N_854,N_157,N_22);
nor U855 (N_855,N_328,N_121);
or U856 (N_856,N_310,N_267);
xnor U857 (N_857,N_263,N_327);
and U858 (N_858,N_392,N_325);
and U859 (N_859,N_151,N_75);
nor U860 (N_860,N_8,N_493);
and U861 (N_861,N_280,N_12);
xnor U862 (N_862,N_442,N_103);
nand U863 (N_863,N_154,N_149);
or U864 (N_864,N_412,N_473);
and U865 (N_865,N_134,N_337);
nor U866 (N_866,N_129,N_120);
or U867 (N_867,N_154,N_478);
xnor U868 (N_868,N_498,N_238);
and U869 (N_869,N_289,N_424);
nor U870 (N_870,N_74,N_492);
nand U871 (N_871,N_379,N_301);
nand U872 (N_872,N_175,N_313);
and U873 (N_873,N_430,N_361);
and U874 (N_874,N_170,N_460);
and U875 (N_875,N_349,N_312);
nor U876 (N_876,N_226,N_284);
xnor U877 (N_877,N_346,N_375);
xor U878 (N_878,N_80,N_443);
nor U879 (N_879,N_260,N_136);
nor U880 (N_880,N_300,N_23);
and U881 (N_881,N_495,N_196);
xnor U882 (N_882,N_52,N_68);
and U883 (N_883,N_379,N_12);
and U884 (N_884,N_435,N_144);
or U885 (N_885,N_402,N_455);
nor U886 (N_886,N_69,N_369);
xnor U887 (N_887,N_228,N_414);
nand U888 (N_888,N_290,N_155);
and U889 (N_889,N_68,N_184);
nor U890 (N_890,N_65,N_98);
and U891 (N_891,N_135,N_271);
nor U892 (N_892,N_392,N_483);
nand U893 (N_893,N_442,N_90);
nor U894 (N_894,N_235,N_478);
xnor U895 (N_895,N_263,N_285);
and U896 (N_896,N_214,N_326);
nor U897 (N_897,N_350,N_318);
nor U898 (N_898,N_245,N_289);
and U899 (N_899,N_245,N_241);
nand U900 (N_900,N_110,N_281);
and U901 (N_901,N_11,N_211);
nor U902 (N_902,N_482,N_370);
or U903 (N_903,N_381,N_427);
and U904 (N_904,N_25,N_103);
nor U905 (N_905,N_209,N_279);
xor U906 (N_906,N_98,N_43);
xor U907 (N_907,N_412,N_393);
and U908 (N_908,N_443,N_171);
nor U909 (N_909,N_396,N_97);
and U910 (N_910,N_47,N_436);
and U911 (N_911,N_247,N_144);
or U912 (N_912,N_347,N_162);
nand U913 (N_913,N_119,N_376);
or U914 (N_914,N_359,N_315);
xor U915 (N_915,N_402,N_111);
or U916 (N_916,N_12,N_486);
xor U917 (N_917,N_363,N_356);
or U918 (N_918,N_349,N_304);
nor U919 (N_919,N_492,N_50);
nor U920 (N_920,N_176,N_482);
nand U921 (N_921,N_293,N_206);
nand U922 (N_922,N_444,N_66);
xor U923 (N_923,N_112,N_275);
and U924 (N_924,N_374,N_78);
and U925 (N_925,N_314,N_396);
nor U926 (N_926,N_197,N_126);
or U927 (N_927,N_365,N_71);
or U928 (N_928,N_24,N_221);
nand U929 (N_929,N_86,N_334);
nor U930 (N_930,N_122,N_466);
nand U931 (N_931,N_107,N_453);
xor U932 (N_932,N_316,N_426);
xor U933 (N_933,N_73,N_291);
xnor U934 (N_934,N_64,N_412);
nand U935 (N_935,N_55,N_288);
and U936 (N_936,N_373,N_151);
and U937 (N_937,N_50,N_235);
or U938 (N_938,N_453,N_297);
or U939 (N_939,N_390,N_412);
and U940 (N_940,N_487,N_233);
nor U941 (N_941,N_99,N_383);
and U942 (N_942,N_483,N_180);
nand U943 (N_943,N_335,N_389);
nor U944 (N_944,N_384,N_432);
or U945 (N_945,N_144,N_340);
nor U946 (N_946,N_495,N_198);
xnor U947 (N_947,N_99,N_344);
nand U948 (N_948,N_24,N_422);
and U949 (N_949,N_127,N_156);
nand U950 (N_950,N_4,N_327);
nor U951 (N_951,N_184,N_497);
nor U952 (N_952,N_198,N_54);
xnor U953 (N_953,N_405,N_167);
xor U954 (N_954,N_429,N_73);
or U955 (N_955,N_183,N_276);
and U956 (N_956,N_189,N_45);
nor U957 (N_957,N_386,N_354);
nor U958 (N_958,N_34,N_357);
xnor U959 (N_959,N_468,N_397);
xnor U960 (N_960,N_390,N_274);
and U961 (N_961,N_313,N_379);
and U962 (N_962,N_266,N_21);
and U963 (N_963,N_167,N_439);
or U964 (N_964,N_1,N_311);
nand U965 (N_965,N_434,N_54);
nand U966 (N_966,N_142,N_487);
or U967 (N_967,N_173,N_287);
or U968 (N_968,N_263,N_336);
xor U969 (N_969,N_341,N_195);
xnor U970 (N_970,N_373,N_452);
xor U971 (N_971,N_356,N_16);
or U972 (N_972,N_221,N_324);
or U973 (N_973,N_194,N_20);
xnor U974 (N_974,N_163,N_344);
nor U975 (N_975,N_201,N_264);
or U976 (N_976,N_156,N_70);
and U977 (N_977,N_381,N_207);
nand U978 (N_978,N_307,N_303);
or U979 (N_979,N_290,N_81);
nor U980 (N_980,N_343,N_223);
nand U981 (N_981,N_330,N_404);
xnor U982 (N_982,N_448,N_229);
and U983 (N_983,N_43,N_54);
nor U984 (N_984,N_397,N_378);
nand U985 (N_985,N_78,N_289);
nor U986 (N_986,N_308,N_87);
xor U987 (N_987,N_236,N_244);
or U988 (N_988,N_380,N_379);
and U989 (N_989,N_417,N_262);
or U990 (N_990,N_361,N_341);
or U991 (N_991,N_263,N_101);
xnor U992 (N_992,N_219,N_321);
nor U993 (N_993,N_201,N_413);
or U994 (N_994,N_409,N_2);
nand U995 (N_995,N_35,N_137);
nor U996 (N_996,N_429,N_332);
xnor U997 (N_997,N_88,N_195);
and U998 (N_998,N_204,N_479);
xnor U999 (N_999,N_105,N_129);
nor U1000 (N_1000,N_812,N_943);
nor U1001 (N_1001,N_517,N_821);
or U1002 (N_1002,N_506,N_775);
and U1003 (N_1003,N_614,N_705);
xnor U1004 (N_1004,N_771,N_648);
nand U1005 (N_1005,N_865,N_670);
nor U1006 (N_1006,N_518,N_950);
and U1007 (N_1007,N_562,N_537);
xnor U1008 (N_1008,N_658,N_822);
and U1009 (N_1009,N_684,N_825);
xnor U1010 (N_1010,N_785,N_897);
nand U1011 (N_1011,N_667,N_853);
or U1012 (N_1012,N_982,N_665);
nor U1013 (N_1013,N_528,N_948);
xnor U1014 (N_1014,N_998,N_792);
or U1015 (N_1015,N_552,N_883);
or U1016 (N_1016,N_762,N_920);
or U1017 (N_1017,N_615,N_979);
xnor U1018 (N_1018,N_902,N_734);
xor U1019 (N_1019,N_931,N_851);
and U1020 (N_1020,N_643,N_758);
nand U1021 (N_1021,N_940,N_676);
nand U1022 (N_1022,N_561,N_895);
or U1023 (N_1023,N_704,N_923);
and U1024 (N_1024,N_873,N_970);
xnor U1025 (N_1025,N_657,N_740);
nand U1026 (N_1026,N_933,N_859);
xnor U1027 (N_1027,N_509,N_751);
xnor U1028 (N_1028,N_627,N_513);
or U1029 (N_1029,N_701,N_815);
nand U1030 (N_1030,N_857,N_663);
nor U1031 (N_1031,N_869,N_942);
nor U1032 (N_1032,N_829,N_955);
nand U1033 (N_1033,N_557,N_721);
xnor U1034 (N_1034,N_660,N_972);
and U1035 (N_1035,N_907,N_661);
xnor U1036 (N_1036,N_674,N_796);
or U1037 (N_1037,N_656,N_534);
and U1038 (N_1038,N_682,N_951);
and U1039 (N_1039,N_543,N_739);
and U1040 (N_1040,N_754,N_995);
nand U1041 (N_1041,N_727,N_742);
and U1042 (N_1042,N_504,N_863);
nand U1043 (N_1043,N_713,N_579);
and U1044 (N_1044,N_949,N_626);
nand U1045 (N_1045,N_725,N_699);
and U1046 (N_1046,N_596,N_935);
nand U1047 (N_1047,N_524,N_582);
nor U1048 (N_1048,N_761,N_500);
or U1049 (N_1049,N_813,N_989);
or U1050 (N_1050,N_885,N_635);
nand U1051 (N_1051,N_847,N_550);
and U1052 (N_1052,N_718,N_954);
or U1053 (N_1053,N_508,N_924);
xor U1054 (N_1054,N_957,N_575);
and U1055 (N_1055,N_953,N_590);
xor U1056 (N_1056,N_547,N_545);
nand U1057 (N_1057,N_605,N_880);
or U1058 (N_1058,N_720,N_722);
nor U1059 (N_1059,N_782,N_572);
and U1060 (N_1060,N_914,N_686);
or U1061 (N_1061,N_881,N_738);
xnor U1062 (N_1062,N_669,N_968);
nand U1063 (N_1063,N_843,N_542);
or U1064 (N_1064,N_811,N_799);
or U1065 (N_1065,N_841,N_803);
nor U1066 (N_1066,N_903,N_532);
or U1067 (N_1067,N_818,N_861);
or U1068 (N_1068,N_872,N_918);
nand U1069 (N_1069,N_555,N_678);
or U1070 (N_1070,N_809,N_616);
xnor U1071 (N_1071,N_639,N_706);
nor U1072 (N_1072,N_697,N_976);
or U1073 (N_1073,N_618,N_574);
xnor U1074 (N_1074,N_934,N_512);
xor U1075 (N_1075,N_988,N_541);
nor U1076 (N_1076,N_798,N_898);
nand U1077 (N_1077,N_717,N_606);
or U1078 (N_1078,N_971,N_571);
or U1079 (N_1079,N_609,N_858);
xor U1080 (N_1080,N_556,N_832);
and U1081 (N_1081,N_905,N_564);
nand U1082 (N_1082,N_689,N_939);
and U1083 (N_1083,N_800,N_620);
nor U1084 (N_1084,N_969,N_780);
xor U1085 (N_1085,N_947,N_553);
nand U1086 (N_1086,N_700,N_752);
nor U1087 (N_1087,N_593,N_788);
xnor U1088 (N_1088,N_756,N_680);
nor U1089 (N_1089,N_549,N_877);
xnor U1090 (N_1090,N_566,N_691);
xor U1091 (N_1091,N_875,N_929);
nand U1092 (N_1092,N_878,N_588);
nor U1093 (N_1093,N_879,N_502);
xnor U1094 (N_1094,N_837,N_540);
xor U1095 (N_1095,N_838,N_709);
and U1096 (N_1096,N_797,N_589);
nand U1097 (N_1097,N_624,N_884);
nand U1098 (N_1098,N_522,N_889);
or U1099 (N_1099,N_833,N_586);
xnor U1100 (N_1100,N_655,N_828);
nor U1101 (N_1101,N_967,N_927);
xor U1102 (N_1102,N_960,N_628);
xnor U1103 (N_1103,N_783,N_594);
xor U1104 (N_1104,N_791,N_505);
and U1105 (N_1105,N_819,N_621);
xnor U1106 (N_1106,N_631,N_787);
or U1107 (N_1107,N_874,N_563);
and U1108 (N_1108,N_985,N_687);
and U1109 (N_1109,N_625,N_611);
nand U1110 (N_1110,N_514,N_850);
or U1111 (N_1111,N_677,N_926);
nand U1112 (N_1112,N_679,N_915);
and U1113 (N_1113,N_731,N_804);
nor U1114 (N_1114,N_852,N_896);
and U1115 (N_1115,N_584,N_745);
nand U1116 (N_1116,N_604,N_735);
xnor U1117 (N_1117,N_781,N_937);
nand U1118 (N_1118,N_793,N_922);
xor U1119 (N_1119,N_784,N_671);
nor U1120 (N_1120,N_645,N_688);
or U1121 (N_1121,N_601,N_710);
or U1122 (N_1122,N_743,N_824);
nor U1123 (N_1123,N_981,N_530);
xnor U1124 (N_1124,N_794,N_632);
nor U1125 (N_1125,N_610,N_629);
nor U1126 (N_1126,N_597,N_892);
nand U1127 (N_1127,N_652,N_741);
nor U1128 (N_1128,N_765,N_980);
nand U1129 (N_1129,N_666,N_723);
nor U1130 (N_1130,N_577,N_757);
and U1131 (N_1131,N_816,N_826);
nor U1132 (N_1132,N_997,N_978);
or U1133 (N_1133,N_580,N_567);
xnor U1134 (N_1134,N_763,N_692);
and U1135 (N_1135,N_591,N_855);
or U1136 (N_1136,N_592,N_759);
xnor U1137 (N_1137,N_768,N_503);
xor U1138 (N_1138,N_559,N_888);
nor U1139 (N_1139,N_844,N_527);
or U1140 (N_1140,N_977,N_846);
nand U1141 (N_1141,N_962,N_983);
nor U1142 (N_1142,N_917,N_755);
nor U1143 (N_1143,N_640,N_866);
nand U1144 (N_1144,N_945,N_776);
nor U1145 (N_1145,N_702,N_786);
nor U1146 (N_1146,N_778,N_636);
nor U1147 (N_1147,N_807,N_908);
or U1148 (N_1148,N_840,N_901);
nor U1149 (N_1149,N_521,N_644);
nand U1150 (N_1150,N_906,N_696);
and U1151 (N_1151,N_569,N_619);
and U1152 (N_1152,N_820,N_726);
or U1153 (N_1153,N_769,N_890);
nand U1154 (N_1154,N_693,N_544);
nor U1155 (N_1155,N_810,N_675);
nand U1156 (N_1156,N_694,N_959);
nand U1157 (N_1157,N_737,N_539);
nand U1158 (N_1158,N_952,N_790);
nor U1159 (N_1159,N_876,N_827);
or U1160 (N_1160,N_930,N_641);
and U1161 (N_1161,N_899,N_685);
and U1162 (N_1162,N_817,N_690);
nand U1163 (N_1163,N_871,N_913);
nand U1164 (N_1164,N_975,N_712);
nor U1165 (N_1165,N_538,N_845);
and U1166 (N_1166,N_507,N_729);
and U1167 (N_1167,N_617,N_573);
and U1168 (N_1168,N_623,N_515);
nor U1169 (N_1169,N_576,N_650);
nand U1170 (N_1170,N_554,N_996);
nor U1171 (N_1171,N_747,N_613);
and U1172 (N_1172,N_568,N_802);
or U1173 (N_1173,N_622,N_766);
or U1174 (N_1174,N_707,N_649);
and U1175 (N_1175,N_744,N_990);
and U1176 (N_1176,N_711,N_984);
or U1177 (N_1177,N_634,N_728);
or U1178 (N_1178,N_773,N_638);
xor U1179 (N_1179,N_991,N_664);
and U1180 (N_1180,N_719,N_642);
xor U1181 (N_1181,N_647,N_633);
nor U1182 (N_1182,N_900,N_830);
nor U1183 (N_1183,N_578,N_839);
xor U1184 (N_1184,N_795,N_925);
and U1185 (N_1185,N_546,N_854);
xor U1186 (N_1186,N_748,N_753);
nand U1187 (N_1187,N_912,N_864);
xor U1188 (N_1188,N_867,N_662);
and U1189 (N_1189,N_558,N_834);
or U1190 (N_1190,N_520,N_630);
or U1191 (N_1191,N_986,N_548);
nand U1192 (N_1192,N_767,N_886);
xor U1193 (N_1193,N_535,N_603);
or U1194 (N_1194,N_746,N_993);
nand U1195 (N_1195,N_992,N_668);
xnor U1196 (N_1196,N_695,N_585);
nor U1197 (N_1197,N_510,N_772);
nor U1198 (N_1198,N_893,N_501);
or U1199 (N_1199,N_806,N_570);
and U1200 (N_1200,N_525,N_760);
nand U1201 (N_1201,N_919,N_715);
or U1202 (N_1202,N_789,N_973);
nor U1203 (N_1203,N_921,N_598);
and U1204 (N_1204,N_904,N_511);
nor U1205 (N_1205,N_836,N_966);
and U1206 (N_1206,N_681,N_910);
or U1207 (N_1207,N_560,N_956);
nor U1208 (N_1208,N_963,N_909);
nor U1209 (N_1209,N_831,N_523);
and U1210 (N_1210,N_730,N_736);
and U1211 (N_1211,N_974,N_607);
nand U1212 (N_1212,N_938,N_958);
and U1213 (N_1213,N_911,N_946);
or U1214 (N_1214,N_551,N_862);
or U1215 (N_1215,N_529,N_999);
nand U1216 (N_1216,N_531,N_987);
nor U1217 (N_1217,N_749,N_961);
and U1218 (N_1218,N_887,N_637);
and U1219 (N_1219,N_870,N_882);
xnor U1220 (N_1220,N_849,N_519);
or U1221 (N_1221,N_608,N_703);
nor U1222 (N_1222,N_894,N_595);
xnor U1223 (N_1223,N_774,N_856);
or U1224 (N_1224,N_891,N_994);
nor U1225 (N_1225,N_928,N_808);
xor U1226 (N_1226,N_733,N_651);
nand U1227 (N_1227,N_750,N_714);
nand U1228 (N_1228,N_565,N_823);
or U1229 (N_1229,N_932,N_835);
or U1230 (N_1230,N_777,N_965);
nor U1231 (N_1231,N_716,N_805);
or U1232 (N_1232,N_916,N_599);
nor U1233 (N_1233,N_654,N_941);
and U1234 (N_1234,N_944,N_653);
or U1235 (N_1235,N_672,N_516);
nor U1236 (N_1236,N_536,N_587);
and U1237 (N_1237,N_698,N_814);
nand U1238 (N_1238,N_732,N_801);
nand U1239 (N_1239,N_581,N_724);
nand U1240 (N_1240,N_868,N_673);
xnor U1241 (N_1241,N_708,N_860);
and U1242 (N_1242,N_659,N_583);
nand U1243 (N_1243,N_842,N_848);
nor U1244 (N_1244,N_683,N_612);
and U1245 (N_1245,N_764,N_770);
nand U1246 (N_1246,N_602,N_936);
nor U1247 (N_1247,N_600,N_964);
and U1248 (N_1248,N_779,N_533);
nand U1249 (N_1249,N_646,N_526);
nor U1250 (N_1250,N_665,N_709);
nand U1251 (N_1251,N_842,N_834);
nand U1252 (N_1252,N_819,N_862);
or U1253 (N_1253,N_734,N_798);
or U1254 (N_1254,N_869,N_835);
nor U1255 (N_1255,N_532,N_665);
nor U1256 (N_1256,N_831,N_881);
nor U1257 (N_1257,N_560,N_665);
xnor U1258 (N_1258,N_974,N_878);
and U1259 (N_1259,N_576,N_547);
or U1260 (N_1260,N_825,N_996);
and U1261 (N_1261,N_587,N_661);
xnor U1262 (N_1262,N_983,N_699);
and U1263 (N_1263,N_564,N_890);
or U1264 (N_1264,N_508,N_860);
and U1265 (N_1265,N_922,N_740);
xnor U1266 (N_1266,N_524,N_889);
nor U1267 (N_1267,N_514,N_511);
nand U1268 (N_1268,N_637,N_735);
and U1269 (N_1269,N_935,N_706);
xor U1270 (N_1270,N_733,N_783);
xnor U1271 (N_1271,N_575,N_518);
and U1272 (N_1272,N_993,N_621);
or U1273 (N_1273,N_630,N_553);
nand U1274 (N_1274,N_966,N_529);
nor U1275 (N_1275,N_729,N_761);
nand U1276 (N_1276,N_926,N_757);
or U1277 (N_1277,N_984,N_878);
xnor U1278 (N_1278,N_586,N_564);
or U1279 (N_1279,N_614,N_735);
or U1280 (N_1280,N_574,N_694);
nor U1281 (N_1281,N_656,N_541);
or U1282 (N_1282,N_916,N_895);
or U1283 (N_1283,N_572,N_828);
and U1284 (N_1284,N_829,N_923);
and U1285 (N_1285,N_996,N_880);
nor U1286 (N_1286,N_619,N_526);
or U1287 (N_1287,N_763,N_968);
and U1288 (N_1288,N_683,N_547);
xnor U1289 (N_1289,N_713,N_596);
nand U1290 (N_1290,N_544,N_977);
nor U1291 (N_1291,N_713,N_765);
or U1292 (N_1292,N_547,N_531);
or U1293 (N_1293,N_634,N_802);
or U1294 (N_1294,N_603,N_932);
nor U1295 (N_1295,N_775,N_865);
nor U1296 (N_1296,N_841,N_738);
or U1297 (N_1297,N_513,N_660);
or U1298 (N_1298,N_692,N_634);
nor U1299 (N_1299,N_913,N_532);
nor U1300 (N_1300,N_950,N_960);
and U1301 (N_1301,N_561,N_754);
xnor U1302 (N_1302,N_667,N_918);
nor U1303 (N_1303,N_745,N_987);
xnor U1304 (N_1304,N_664,N_794);
or U1305 (N_1305,N_712,N_917);
nand U1306 (N_1306,N_749,N_660);
or U1307 (N_1307,N_645,N_869);
or U1308 (N_1308,N_678,N_558);
nand U1309 (N_1309,N_817,N_604);
nor U1310 (N_1310,N_858,N_780);
nand U1311 (N_1311,N_858,N_723);
nand U1312 (N_1312,N_740,N_926);
nor U1313 (N_1313,N_797,N_967);
and U1314 (N_1314,N_551,N_899);
and U1315 (N_1315,N_754,N_715);
and U1316 (N_1316,N_683,N_789);
nor U1317 (N_1317,N_535,N_820);
or U1318 (N_1318,N_701,N_743);
xnor U1319 (N_1319,N_905,N_648);
nor U1320 (N_1320,N_624,N_763);
or U1321 (N_1321,N_812,N_774);
nor U1322 (N_1322,N_680,N_769);
or U1323 (N_1323,N_848,N_672);
or U1324 (N_1324,N_895,N_781);
nand U1325 (N_1325,N_959,N_749);
or U1326 (N_1326,N_823,N_770);
and U1327 (N_1327,N_548,N_518);
nand U1328 (N_1328,N_600,N_806);
or U1329 (N_1329,N_954,N_577);
xor U1330 (N_1330,N_788,N_842);
or U1331 (N_1331,N_799,N_977);
or U1332 (N_1332,N_980,N_922);
or U1333 (N_1333,N_759,N_577);
nand U1334 (N_1334,N_882,N_583);
nand U1335 (N_1335,N_639,N_774);
xnor U1336 (N_1336,N_787,N_648);
nor U1337 (N_1337,N_850,N_805);
and U1338 (N_1338,N_588,N_989);
or U1339 (N_1339,N_549,N_989);
and U1340 (N_1340,N_836,N_795);
nand U1341 (N_1341,N_763,N_735);
nand U1342 (N_1342,N_540,N_553);
and U1343 (N_1343,N_696,N_996);
nand U1344 (N_1344,N_735,N_503);
or U1345 (N_1345,N_864,N_887);
nand U1346 (N_1346,N_716,N_919);
nand U1347 (N_1347,N_799,N_859);
xnor U1348 (N_1348,N_522,N_833);
or U1349 (N_1349,N_913,N_557);
xnor U1350 (N_1350,N_762,N_713);
nand U1351 (N_1351,N_959,N_521);
and U1352 (N_1352,N_541,N_652);
xnor U1353 (N_1353,N_826,N_920);
and U1354 (N_1354,N_530,N_829);
and U1355 (N_1355,N_803,N_617);
xor U1356 (N_1356,N_703,N_725);
nor U1357 (N_1357,N_666,N_713);
and U1358 (N_1358,N_785,N_635);
xnor U1359 (N_1359,N_952,N_924);
nand U1360 (N_1360,N_857,N_574);
nor U1361 (N_1361,N_709,N_969);
xor U1362 (N_1362,N_630,N_533);
or U1363 (N_1363,N_905,N_757);
nand U1364 (N_1364,N_659,N_951);
nand U1365 (N_1365,N_775,N_786);
nand U1366 (N_1366,N_738,N_769);
xor U1367 (N_1367,N_577,N_675);
xor U1368 (N_1368,N_706,N_694);
xnor U1369 (N_1369,N_922,N_635);
or U1370 (N_1370,N_752,N_851);
xnor U1371 (N_1371,N_878,N_544);
xnor U1372 (N_1372,N_527,N_510);
xnor U1373 (N_1373,N_514,N_551);
nor U1374 (N_1374,N_961,N_899);
and U1375 (N_1375,N_790,N_882);
or U1376 (N_1376,N_684,N_956);
xor U1377 (N_1377,N_607,N_677);
or U1378 (N_1378,N_654,N_963);
nand U1379 (N_1379,N_895,N_850);
and U1380 (N_1380,N_513,N_833);
nand U1381 (N_1381,N_913,N_820);
and U1382 (N_1382,N_606,N_602);
and U1383 (N_1383,N_794,N_898);
or U1384 (N_1384,N_630,N_626);
or U1385 (N_1385,N_713,N_864);
nand U1386 (N_1386,N_949,N_812);
nor U1387 (N_1387,N_617,N_838);
or U1388 (N_1388,N_938,N_968);
xnor U1389 (N_1389,N_837,N_694);
or U1390 (N_1390,N_544,N_545);
nand U1391 (N_1391,N_514,N_746);
xor U1392 (N_1392,N_897,N_577);
xor U1393 (N_1393,N_960,N_585);
nand U1394 (N_1394,N_925,N_735);
nor U1395 (N_1395,N_656,N_642);
nand U1396 (N_1396,N_563,N_521);
or U1397 (N_1397,N_862,N_593);
xor U1398 (N_1398,N_729,N_905);
and U1399 (N_1399,N_680,N_746);
nand U1400 (N_1400,N_668,N_888);
and U1401 (N_1401,N_596,N_816);
nand U1402 (N_1402,N_888,N_774);
xnor U1403 (N_1403,N_878,N_903);
or U1404 (N_1404,N_774,N_509);
xor U1405 (N_1405,N_886,N_578);
nand U1406 (N_1406,N_628,N_657);
nor U1407 (N_1407,N_903,N_868);
xnor U1408 (N_1408,N_631,N_981);
xnor U1409 (N_1409,N_522,N_870);
nand U1410 (N_1410,N_919,N_587);
and U1411 (N_1411,N_609,N_714);
nor U1412 (N_1412,N_641,N_942);
or U1413 (N_1413,N_652,N_938);
nor U1414 (N_1414,N_602,N_539);
nor U1415 (N_1415,N_669,N_972);
xnor U1416 (N_1416,N_759,N_897);
or U1417 (N_1417,N_528,N_726);
nor U1418 (N_1418,N_540,N_838);
nor U1419 (N_1419,N_844,N_953);
xor U1420 (N_1420,N_778,N_723);
nor U1421 (N_1421,N_540,N_598);
nand U1422 (N_1422,N_796,N_926);
nor U1423 (N_1423,N_709,N_981);
nor U1424 (N_1424,N_877,N_824);
nand U1425 (N_1425,N_567,N_627);
nand U1426 (N_1426,N_614,N_834);
nor U1427 (N_1427,N_693,N_961);
nor U1428 (N_1428,N_510,N_640);
nand U1429 (N_1429,N_997,N_707);
nor U1430 (N_1430,N_968,N_640);
or U1431 (N_1431,N_608,N_754);
nor U1432 (N_1432,N_563,N_549);
nand U1433 (N_1433,N_859,N_778);
or U1434 (N_1434,N_697,N_858);
and U1435 (N_1435,N_868,N_590);
nand U1436 (N_1436,N_716,N_559);
nor U1437 (N_1437,N_900,N_790);
xor U1438 (N_1438,N_747,N_579);
nor U1439 (N_1439,N_949,N_980);
and U1440 (N_1440,N_877,N_509);
nand U1441 (N_1441,N_831,N_651);
nor U1442 (N_1442,N_775,N_873);
nand U1443 (N_1443,N_741,N_862);
xor U1444 (N_1444,N_674,N_706);
nor U1445 (N_1445,N_554,N_648);
and U1446 (N_1446,N_604,N_780);
nor U1447 (N_1447,N_829,N_746);
nand U1448 (N_1448,N_563,N_815);
or U1449 (N_1449,N_998,N_631);
and U1450 (N_1450,N_677,N_509);
nand U1451 (N_1451,N_994,N_585);
xnor U1452 (N_1452,N_572,N_838);
or U1453 (N_1453,N_835,N_506);
or U1454 (N_1454,N_597,N_879);
nand U1455 (N_1455,N_780,N_795);
xnor U1456 (N_1456,N_516,N_898);
or U1457 (N_1457,N_851,N_551);
nor U1458 (N_1458,N_510,N_949);
nor U1459 (N_1459,N_736,N_501);
or U1460 (N_1460,N_922,N_890);
xor U1461 (N_1461,N_689,N_903);
nor U1462 (N_1462,N_996,N_888);
or U1463 (N_1463,N_511,N_952);
and U1464 (N_1464,N_804,N_961);
xnor U1465 (N_1465,N_984,N_628);
or U1466 (N_1466,N_685,N_572);
and U1467 (N_1467,N_555,N_657);
or U1468 (N_1468,N_845,N_743);
xor U1469 (N_1469,N_815,N_618);
or U1470 (N_1470,N_727,N_923);
or U1471 (N_1471,N_511,N_731);
and U1472 (N_1472,N_532,N_694);
nor U1473 (N_1473,N_647,N_631);
and U1474 (N_1474,N_716,N_894);
or U1475 (N_1475,N_961,N_567);
nor U1476 (N_1476,N_893,N_866);
and U1477 (N_1477,N_680,N_695);
and U1478 (N_1478,N_770,N_992);
and U1479 (N_1479,N_580,N_594);
nor U1480 (N_1480,N_887,N_918);
or U1481 (N_1481,N_881,N_788);
xor U1482 (N_1482,N_984,N_835);
xor U1483 (N_1483,N_840,N_777);
and U1484 (N_1484,N_670,N_577);
or U1485 (N_1485,N_915,N_504);
nor U1486 (N_1486,N_773,N_878);
nand U1487 (N_1487,N_847,N_793);
nand U1488 (N_1488,N_699,N_702);
nand U1489 (N_1489,N_994,N_653);
nand U1490 (N_1490,N_703,N_592);
nand U1491 (N_1491,N_697,N_884);
or U1492 (N_1492,N_830,N_524);
nand U1493 (N_1493,N_678,N_663);
nor U1494 (N_1494,N_595,N_856);
and U1495 (N_1495,N_716,N_690);
nor U1496 (N_1496,N_834,N_900);
and U1497 (N_1497,N_644,N_688);
xnor U1498 (N_1498,N_990,N_780);
nand U1499 (N_1499,N_721,N_700);
xnor U1500 (N_1500,N_1201,N_1479);
xor U1501 (N_1501,N_1040,N_1128);
nor U1502 (N_1502,N_1134,N_1209);
xor U1503 (N_1503,N_1308,N_1327);
and U1504 (N_1504,N_1016,N_1068);
nand U1505 (N_1505,N_1026,N_1458);
nor U1506 (N_1506,N_1385,N_1136);
and U1507 (N_1507,N_1153,N_1064);
nor U1508 (N_1508,N_1324,N_1426);
xor U1509 (N_1509,N_1462,N_1244);
or U1510 (N_1510,N_1216,N_1012);
xnor U1511 (N_1511,N_1157,N_1151);
or U1512 (N_1512,N_1264,N_1230);
nor U1513 (N_1513,N_1352,N_1088);
nor U1514 (N_1514,N_1343,N_1160);
nand U1515 (N_1515,N_1059,N_1311);
and U1516 (N_1516,N_1172,N_1204);
or U1517 (N_1517,N_1250,N_1115);
nor U1518 (N_1518,N_1390,N_1326);
xnor U1519 (N_1519,N_1333,N_1362);
nand U1520 (N_1520,N_1213,N_1152);
or U1521 (N_1521,N_1120,N_1183);
or U1522 (N_1522,N_1382,N_1232);
or U1523 (N_1523,N_1018,N_1001);
or U1524 (N_1524,N_1484,N_1102);
and U1525 (N_1525,N_1010,N_1089);
or U1526 (N_1526,N_1450,N_1144);
and U1527 (N_1527,N_1127,N_1052);
or U1528 (N_1528,N_1117,N_1242);
and U1529 (N_1529,N_1286,N_1495);
xor U1530 (N_1530,N_1021,N_1061);
and U1531 (N_1531,N_1175,N_1181);
nor U1532 (N_1532,N_1218,N_1268);
or U1533 (N_1533,N_1245,N_1258);
and U1534 (N_1534,N_1474,N_1078);
or U1535 (N_1535,N_1377,N_1491);
xor U1536 (N_1536,N_1079,N_1101);
nand U1537 (N_1537,N_1416,N_1289);
and U1538 (N_1538,N_1497,N_1256);
nor U1539 (N_1539,N_1345,N_1374);
or U1540 (N_1540,N_1186,N_1187);
nor U1541 (N_1541,N_1370,N_1276);
xor U1542 (N_1542,N_1036,N_1116);
xor U1543 (N_1543,N_1174,N_1348);
and U1544 (N_1544,N_1193,N_1130);
nand U1545 (N_1545,N_1364,N_1022);
xor U1546 (N_1546,N_1277,N_1257);
nor U1547 (N_1547,N_1274,N_1284);
or U1548 (N_1548,N_1261,N_1035);
or U1549 (N_1549,N_1192,N_1231);
nand U1550 (N_1550,N_1372,N_1243);
nand U1551 (N_1551,N_1240,N_1017);
or U1552 (N_1552,N_1471,N_1486);
or U1553 (N_1553,N_1060,N_1341);
or U1554 (N_1554,N_1007,N_1143);
xnor U1555 (N_1555,N_1464,N_1415);
xor U1556 (N_1556,N_1019,N_1205);
nand U1557 (N_1557,N_1373,N_1161);
nand U1558 (N_1558,N_1121,N_1470);
nor U1559 (N_1559,N_1493,N_1321);
nor U1560 (N_1560,N_1452,N_1169);
nand U1561 (N_1561,N_1400,N_1113);
xor U1562 (N_1562,N_1328,N_1401);
nor U1563 (N_1563,N_1198,N_1297);
nor U1564 (N_1564,N_1330,N_1062);
nand U1565 (N_1565,N_1338,N_1190);
and U1566 (N_1566,N_1032,N_1002);
xor U1567 (N_1567,N_1265,N_1421);
or U1568 (N_1568,N_1315,N_1476);
and U1569 (N_1569,N_1309,N_1389);
nand U1570 (N_1570,N_1070,N_1069);
xnor U1571 (N_1571,N_1428,N_1106);
xor U1572 (N_1572,N_1039,N_1044);
and U1573 (N_1573,N_1425,N_1149);
or U1574 (N_1574,N_1446,N_1472);
nand U1575 (N_1575,N_1383,N_1422);
nor U1576 (N_1576,N_1434,N_1033);
or U1577 (N_1577,N_1260,N_1394);
nor U1578 (N_1578,N_1312,N_1133);
xnor U1579 (N_1579,N_1015,N_1063);
and U1580 (N_1580,N_1357,N_1456);
xor U1581 (N_1581,N_1168,N_1483);
and U1582 (N_1582,N_1359,N_1272);
and U1583 (N_1583,N_1030,N_1222);
nand U1584 (N_1584,N_1498,N_1057);
or U1585 (N_1585,N_1131,N_1455);
nand U1586 (N_1586,N_1004,N_1013);
xor U1587 (N_1587,N_1259,N_1378);
or U1588 (N_1588,N_1356,N_1165);
and U1589 (N_1589,N_1454,N_1171);
nand U1590 (N_1590,N_1103,N_1110);
nand U1591 (N_1591,N_1191,N_1184);
nand U1592 (N_1592,N_1212,N_1478);
and U1593 (N_1593,N_1066,N_1282);
nor U1594 (N_1594,N_1252,N_1273);
nor U1595 (N_1595,N_1140,N_1298);
nand U1596 (N_1596,N_1367,N_1405);
and U1597 (N_1597,N_1448,N_1224);
xnor U1598 (N_1598,N_1053,N_1482);
nor U1599 (N_1599,N_1047,N_1473);
nand U1600 (N_1600,N_1429,N_1229);
xor U1601 (N_1601,N_1323,N_1339);
xor U1602 (N_1602,N_1335,N_1351);
nand U1603 (N_1603,N_1366,N_1095);
xnor U1604 (N_1604,N_1177,N_1319);
xnor U1605 (N_1605,N_1379,N_1443);
or U1606 (N_1606,N_1275,N_1210);
xnor U1607 (N_1607,N_1307,N_1305);
xnor U1608 (N_1608,N_1148,N_1225);
or U1609 (N_1609,N_1246,N_1402);
nor U1610 (N_1610,N_1361,N_1028);
nor U1611 (N_1611,N_1023,N_1034);
xor U1612 (N_1612,N_1189,N_1251);
or U1613 (N_1613,N_1353,N_1176);
and U1614 (N_1614,N_1269,N_1159);
and U1615 (N_1615,N_1111,N_1219);
nand U1616 (N_1616,N_1197,N_1093);
xnor U1617 (N_1617,N_1238,N_1475);
nand U1618 (N_1618,N_1188,N_1295);
nand U1619 (N_1619,N_1100,N_1334);
and U1620 (N_1620,N_1112,N_1406);
nor U1621 (N_1621,N_1280,N_1027);
nor U1622 (N_1622,N_1099,N_1008);
nor U1623 (N_1623,N_1081,N_1397);
or U1624 (N_1624,N_1077,N_1435);
nor U1625 (N_1625,N_1020,N_1300);
nand U1626 (N_1626,N_1090,N_1006);
and U1627 (N_1627,N_1108,N_1453);
nor U1628 (N_1628,N_1132,N_1185);
or U1629 (N_1629,N_1031,N_1322);
and U1630 (N_1630,N_1166,N_1067);
xnor U1631 (N_1631,N_1221,N_1051);
nor U1632 (N_1632,N_1125,N_1396);
nor U1633 (N_1633,N_1431,N_1045);
xor U1634 (N_1634,N_1096,N_1388);
nor U1635 (N_1635,N_1439,N_1214);
nor U1636 (N_1636,N_1239,N_1387);
nor U1637 (N_1637,N_1075,N_1331);
nand U1638 (N_1638,N_1233,N_1271);
nor U1639 (N_1639,N_1316,N_1228);
nor U1640 (N_1640,N_1043,N_1104);
or U1641 (N_1641,N_1146,N_1349);
xnor U1642 (N_1642,N_1097,N_1417);
and U1643 (N_1643,N_1082,N_1118);
and U1644 (N_1644,N_1485,N_1003);
xnor U1645 (N_1645,N_1206,N_1457);
nand U1646 (N_1646,N_1419,N_1369);
nand U1647 (N_1647,N_1279,N_1332);
and U1648 (N_1648,N_1145,N_1442);
and U1649 (N_1649,N_1365,N_1142);
nand U1650 (N_1650,N_1170,N_1432);
nand U1651 (N_1651,N_1105,N_1314);
xor U1652 (N_1652,N_1156,N_1488);
nor U1653 (N_1653,N_1433,N_1241);
or U1654 (N_1654,N_1194,N_1438);
or U1655 (N_1655,N_1445,N_1226);
and U1656 (N_1656,N_1091,N_1296);
nand U1657 (N_1657,N_1011,N_1107);
and U1658 (N_1658,N_1000,N_1463);
and U1659 (N_1659,N_1492,N_1092);
nand U1660 (N_1660,N_1403,N_1342);
nor U1661 (N_1661,N_1071,N_1267);
and U1662 (N_1662,N_1360,N_1009);
nand U1663 (N_1663,N_1292,N_1025);
nor U1664 (N_1664,N_1293,N_1302);
nand U1665 (N_1665,N_1147,N_1380);
or U1666 (N_1666,N_1014,N_1024);
or U1667 (N_1667,N_1109,N_1072);
xor U1668 (N_1668,N_1208,N_1247);
nand U1669 (N_1669,N_1306,N_1195);
nand U1670 (N_1670,N_1480,N_1150);
xnor U1671 (N_1671,N_1179,N_1469);
nand U1672 (N_1672,N_1126,N_1123);
nor U1673 (N_1673,N_1467,N_1376);
and U1674 (N_1674,N_1227,N_1283);
nor U1675 (N_1675,N_1073,N_1202);
or U1676 (N_1676,N_1310,N_1167);
nor U1677 (N_1677,N_1211,N_1304);
nor U1678 (N_1678,N_1466,N_1220);
xor U1679 (N_1679,N_1249,N_1291);
nor U1680 (N_1680,N_1138,N_1384);
nand U1681 (N_1681,N_1460,N_1158);
nand U1682 (N_1682,N_1329,N_1200);
or U1683 (N_1683,N_1398,N_1420);
xnor U1684 (N_1684,N_1058,N_1355);
nor U1685 (N_1685,N_1489,N_1083);
xnor U1686 (N_1686,N_1203,N_1122);
or U1687 (N_1687,N_1255,N_1087);
or U1688 (N_1688,N_1164,N_1318);
nor U1689 (N_1689,N_1301,N_1325);
xor U1690 (N_1690,N_1029,N_1162);
xor U1691 (N_1691,N_1094,N_1235);
nor U1692 (N_1692,N_1049,N_1487);
nor U1693 (N_1693,N_1371,N_1412);
nand U1694 (N_1694,N_1444,N_1135);
or U1695 (N_1695,N_1119,N_1076);
and U1696 (N_1696,N_1074,N_1410);
nand U1697 (N_1697,N_1358,N_1290);
or U1698 (N_1698,N_1129,N_1395);
and U1699 (N_1699,N_1375,N_1137);
nand U1700 (N_1700,N_1451,N_1281);
nor U1701 (N_1701,N_1368,N_1391);
nor U1702 (N_1702,N_1499,N_1336);
xor U1703 (N_1703,N_1248,N_1465);
xnor U1704 (N_1704,N_1299,N_1354);
and U1705 (N_1705,N_1303,N_1468);
and U1706 (N_1706,N_1163,N_1350);
xor U1707 (N_1707,N_1278,N_1139);
xor U1708 (N_1708,N_1178,N_1447);
nand U1709 (N_1709,N_1337,N_1196);
xor U1710 (N_1710,N_1437,N_1086);
or U1711 (N_1711,N_1477,N_1363);
or U1712 (N_1712,N_1234,N_1423);
xor U1713 (N_1713,N_1223,N_1408);
or U1714 (N_1714,N_1392,N_1217);
nor U1715 (N_1715,N_1461,N_1294);
nor U1716 (N_1716,N_1490,N_1005);
and U1717 (N_1717,N_1114,N_1346);
xor U1718 (N_1718,N_1182,N_1386);
xnor U1719 (N_1719,N_1084,N_1407);
nand U1720 (N_1720,N_1496,N_1347);
or U1721 (N_1721,N_1494,N_1124);
xnor U1722 (N_1722,N_1413,N_1048);
or U1723 (N_1723,N_1055,N_1427);
nor U1724 (N_1724,N_1037,N_1253);
nor U1725 (N_1725,N_1154,N_1270);
or U1726 (N_1726,N_1287,N_1141);
xor U1727 (N_1727,N_1065,N_1424);
or U1728 (N_1728,N_1215,N_1393);
xor U1729 (N_1729,N_1041,N_1038);
and U1730 (N_1730,N_1436,N_1199);
nand U1731 (N_1731,N_1046,N_1263);
xor U1732 (N_1732,N_1414,N_1098);
nor U1733 (N_1733,N_1180,N_1340);
xnor U1734 (N_1734,N_1430,N_1320);
or U1735 (N_1735,N_1155,N_1317);
nand U1736 (N_1736,N_1481,N_1262);
xor U1737 (N_1737,N_1441,N_1050);
xor U1738 (N_1738,N_1404,N_1440);
nor U1739 (N_1739,N_1056,N_1459);
and U1740 (N_1740,N_1054,N_1042);
xor U1741 (N_1741,N_1449,N_1173);
or U1742 (N_1742,N_1085,N_1418);
or U1743 (N_1743,N_1285,N_1381);
nand U1744 (N_1744,N_1313,N_1409);
xnor U1745 (N_1745,N_1236,N_1266);
or U1746 (N_1746,N_1254,N_1344);
nor U1747 (N_1747,N_1080,N_1288);
or U1748 (N_1748,N_1411,N_1399);
and U1749 (N_1749,N_1237,N_1207);
xnor U1750 (N_1750,N_1437,N_1198);
nand U1751 (N_1751,N_1489,N_1136);
nor U1752 (N_1752,N_1030,N_1491);
xor U1753 (N_1753,N_1248,N_1403);
xnor U1754 (N_1754,N_1334,N_1061);
and U1755 (N_1755,N_1065,N_1480);
and U1756 (N_1756,N_1060,N_1313);
and U1757 (N_1757,N_1224,N_1430);
or U1758 (N_1758,N_1294,N_1099);
and U1759 (N_1759,N_1267,N_1293);
nor U1760 (N_1760,N_1143,N_1350);
nand U1761 (N_1761,N_1115,N_1105);
and U1762 (N_1762,N_1323,N_1458);
nor U1763 (N_1763,N_1203,N_1421);
nand U1764 (N_1764,N_1399,N_1267);
and U1765 (N_1765,N_1303,N_1416);
xnor U1766 (N_1766,N_1448,N_1143);
xnor U1767 (N_1767,N_1429,N_1407);
nor U1768 (N_1768,N_1206,N_1448);
xnor U1769 (N_1769,N_1153,N_1444);
and U1770 (N_1770,N_1397,N_1276);
xor U1771 (N_1771,N_1368,N_1079);
nor U1772 (N_1772,N_1169,N_1256);
xnor U1773 (N_1773,N_1048,N_1363);
and U1774 (N_1774,N_1177,N_1050);
or U1775 (N_1775,N_1390,N_1017);
xnor U1776 (N_1776,N_1485,N_1470);
nor U1777 (N_1777,N_1225,N_1416);
nand U1778 (N_1778,N_1172,N_1082);
and U1779 (N_1779,N_1049,N_1306);
xnor U1780 (N_1780,N_1037,N_1428);
nand U1781 (N_1781,N_1018,N_1238);
nand U1782 (N_1782,N_1209,N_1318);
nor U1783 (N_1783,N_1085,N_1017);
xor U1784 (N_1784,N_1276,N_1471);
nor U1785 (N_1785,N_1215,N_1375);
or U1786 (N_1786,N_1195,N_1259);
nor U1787 (N_1787,N_1367,N_1110);
or U1788 (N_1788,N_1177,N_1458);
or U1789 (N_1789,N_1194,N_1464);
nor U1790 (N_1790,N_1312,N_1059);
nand U1791 (N_1791,N_1471,N_1286);
or U1792 (N_1792,N_1004,N_1005);
xor U1793 (N_1793,N_1431,N_1255);
nor U1794 (N_1794,N_1355,N_1487);
or U1795 (N_1795,N_1352,N_1130);
and U1796 (N_1796,N_1233,N_1163);
xor U1797 (N_1797,N_1359,N_1388);
nor U1798 (N_1798,N_1017,N_1252);
nor U1799 (N_1799,N_1133,N_1453);
nand U1800 (N_1800,N_1214,N_1147);
nand U1801 (N_1801,N_1330,N_1192);
or U1802 (N_1802,N_1038,N_1279);
nor U1803 (N_1803,N_1466,N_1166);
nand U1804 (N_1804,N_1404,N_1445);
and U1805 (N_1805,N_1424,N_1415);
xnor U1806 (N_1806,N_1346,N_1393);
or U1807 (N_1807,N_1189,N_1047);
and U1808 (N_1808,N_1231,N_1435);
and U1809 (N_1809,N_1144,N_1329);
nand U1810 (N_1810,N_1099,N_1036);
and U1811 (N_1811,N_1289,N_1425);
nor U1812 (N_1812,N_1153,N_1349);
and U1813 (N_1813,N_1392,N_1179);
or U1814 (N_1814,N_1498,N_1245);
or U1815 (N_1815,N_1388,N_1347);
nand U1816 (N_1816,N_1202,N_1147);
nand U1817 (N_1817,N_1256,N_1065);
nor U1818 (N_1818,N_1238,N_1035);
and U1819 (N_1819,N_1059,N_1083);
nor U1820 (N_1820,N_1122,N_1431);
xor U1821 (N_1821,N_1191,N_1024);
or U1822 (N_1822,N_1391,N_1163);
and U1823 (N_1823,N_1024,N_1362);
nor U1824 (N_1824,N_1473,N_1160);
or U1825 (N_1825,N_1377,N_1463);
and U1826 (N_1826,N_1404,N_1089);
or U1827 (N_1827,N_1350,N_1011);
or U1828 (N_1828,N_1013,N_1441);
or U1829 (N_1829,N_1427,N_1109);
xor U1830 (N_1830,N_1174,N_1113);
or U1831 (N_1831,N_1198,N_1260);
nor U1832 (N_1832,N_1252,N_1259);
xnor U1833 (N_1833,N_1059,N_1328);
and U1834 (N_1834,N_1245,N_1444);
xor U1835 (N_1835,N_1348,N_1164);
and U1836 (N_1836,N_1247,N_1352);
xor U1837 (N_1837,N_1372,N_1279);
nor U1838 (N_1838,N_1440,N_1030);
or U1839 (N_1839,N_1489,N_1333);
or U1840 (N_1840,N_1385,N_1286);
or U1841 (N_1841,N_1044,N_1276);
nand U1842 (N_1842,N_1044,N_1311);
or U1843 (N_1843,N_1358,N_1287);
nor U1844 (N_1844,N_1368,N_1076);
or U1845 (N_1845,N_1337,N_1351);
nor U1846 (N_1846,N_1193,N_1492);
nor U1847 (N_1847,N_1275,N_1375);
or U1848 (N_1848,N_1073,N_1078);
nor U1849 (N_1849,N_1361,N_1212);
or U1850 (N_1850,N_1146,N_1262);
xnor U1851 (N_1851,N_1098,N_1454);
nand U1852 (N_1852,N_1257,N_1382);
or U1853 (N_1853,N_1281,N_1484);
nand U1854 (N_1854,N_1211,N_1437);
nand U1855 (N_1855,N_1021,N_1318);
nor U1856 (N_1856,N_1247,N_1293);
nor U1857 (N_1857,N_1485,N_1125);
xnor U1858 (N_1858,N_1445,N_1021);
or U1859 (N_1859,N_1429,N_1056);
xnor U1860 (N_1860,N_1185,N_1273);
and U1861 (N_1861,N_1435,N_1147);
and U1862 (N_1862,N_1172,N_1203);
and U1863 (N_1863,N_1086,N_1095);
xnor U1864 (N_1864,N_1271,N_1354);
nor U1865 (N_1865,N_1299,N_1292);
nor U1866 (N_1866,N_1103,N_1346);
xnor U1867 (N_1867,N_1323,N_1011);
and U1868 (N_1868,N_1334,N_1030);
and U1869 (N_1869,N_1008,N_1172);
nor U1870 (N_1870,N_1418,N_1205);
nand U1871 (N_1871,N_1400,N_1158);
and U1872 (N_1872,N_1307,N_1243);
nand U1873 (N_1873,N_1317,N_1111);
and U1874 (N_1874,N_1448,N_1423);
nand U1875 (N_1875,N_1367,N_1134);
nand U1876 (N_1876,N_1284,N_1146);
nor U1877 (N_1877,N_1003,N_1122);
xnor U1878 (N_1878,N_1262,N_1157);
or U1879 (N_1879,N_1076,N_1341);
xnor U1880 (N_1880,N_1427,N_1331);
nand U1881 (N_1881,N_1019,N_1107);
nor U1882 (N_1882,N_1297,N_1325);
xor U1883 (N_1883,N_1262,N_1143);
nand U1884 (N_1884,N_1108,N_1477);
or U1885 (N_1885,N_1375,N_1212);
xnor U1886 (N_1886,N_1263,N_1111);
and U1887 (N_1887,N_1380,N_1101);
or U1888 (N_1888,N_1116,N_1350);
xnor U1889 (N_1889,N_1203,N_1488);
xor U1890 (N_1890,N_1372,N_1143);
nor U1891 (N_1891,N_1161,N_1408);
xnor U1892 (N_1892,N_1366,N_1440);
nand U1893 (N_1893,N_1239,N_1270);
nor U1894 (N_1894,N_1371,N_1451);
nand U1895 (N_1895,N_1027,N_1392);
or U1896 (N_1896,N_1202,N_1171);
or U1897 (N_1897,N_1235,N_1157);
nand U1898 (N_1898,N_1093,N_1264);
or U1899 (N_1899,N_1487,N_1154);
nor U1900 (N_1900,N_1414,N_1221);
nor U1901 (N_1901,N_1251,N_1269);
and U1902 (N_1902,N_1024,N_1094);
nand U1903 (N_1903,N_1362,N_1398);
xnor U1904 (N_1904,N_1218,N_1161);
nor U1905 (N_1905,N_1257,N_1124);
and U1906 (N_1906,N_1245,N_1421);
xnor U1907 (N_1907,N_1177,N_1333);
and U1908 (N_1908,N_1229,N_1280);
xor U1909 (N_1909,N_1309,N_1477);
and U1910 (N_1910,N_1107,N_1238);
nand U1911 (N_1911,N_1436,N_1308);
nor U1912 (N_1912,N_1247,N_1360);
nand U1913 (N_1913,N_1208,N_1328);
nand U1914 (N_1914,N_1271,N_1052);
and U1915 (N_1915,N_1198,N_1209);
nor U1916 (N_1916,N_1215,N_1181);
or U1917 (N_1917,N_1136,N_1429);
nand U1918 (N_1918,N_1319,N_1030);
and U1919 (N_1919,N_1222,N_1483);
xor U1920 (N_1920,N_1081,N_1176);
and U1921 (N_1921,N_1310,N_1235);
or U1922 (N_1922,N_1028,N_1125);
or U1923 (N_1923,N_1418,N_1268);
and U1924 (N_1924,N_1019,N_1186);
xor U1925 (N_1925,N_1042,N_1351);
nor U1926 (N_1926,N_1044,N_1063);
or U1927 (N_1927,N_1008,N_1144);
xor U1928 (N_1928,N_1247,N_1120);
nor U1929 (N_1929,N_1222,N_1092);
nor U1930 (N_1930,N_1215,N_1402);
or U1931 (N_1931,N_1390,N_1325);
or U1932 (N_1932,N_1046,N_1232);
xor U1933 (N_1933,N_1420,N_1215);
or U1934 (N_1934,N_1089,N_1240);
and U1935 (N_1935,N_1291,N_1421);
and U1936 (N_1936,N_1046,N_1422);
and U1937 (N_1937,N_1443,N_1294);
or U1938 (N_1938,N_1435,N_1438);
nand U1939 (N_1939,N_1341,N_1358);
xnor U1940 (N_1940,N_1461,N_1348);
nor U1941 (N_1941,N_1240,N_1111);
xor U1942 (N_1942,N_1266,N_1111);
and U1943 (N_1943,N_1287,N_1290);
xnor U1944 (N_1944,N_1278,N_1350);
or U1945 (N_1945,N_1109,N_1309);
xor U1946 (N_1946,N_1483,N_1357);
and U1947 (N_1947,N_1058,N_1020);
or U1948 (N_1948,N_1227,N_1020);
xor U1949 (N_1949,N_1194,N_1130);
and U1950 (N_1950,N_1395,N_1270);
or U1951 (N_1951,N_1348,N_1008);
xnor U1952 (N_1952,N_1490,N_1338);
and U1953 (N_1953,N_1330,N_1390);
nand U1954 (N_1954,N_1086,N_1130);
nor U1955 (N_1955,N_1457,N_1253);
nor U1956 (N_1956,N_1171,N_1195);
xor U1957 (N_1957,N_1480,N_1379);
xor U1958 (N_1958,N_1342,N_1212);
and U1959 (N_1959,N_1006,N_1198);
xnor U1960 (N_1960,N_1238,N_1177);
nand U1961 (N_1961,N_1263,N_1170);
or U1962 (N_1962,N_1177,N_1002);
and U1963 (N_1963,N_1122,N_1486);
or U1964 (N_1964,N_1424,N_1281);
xnor U1965 (N_1965,N_1443,N_1284);
and U1966 (N_1966,N_1368,N_1331);
and U1967 (N_1967,N_1012,N_1327);
and U1968 (N_1968,N_1449,N_1051);
nand U1969 (N_1969,N_1335,N_1027);
and U1970 (N_1970,N_1396,N_1048);
xor U1971 (N_1971,N_1020,N_1395);
nor U1972 (N_1972,N_1277,N_1022);
nand U1973 (N_1973,N_1219,N_1080);
nor U1974 (N_1974,N_1244,N_1292);
or U1975 (N_1975,N_1483,N_1079);
and U1976 (N_1976,N_1347,N_1472);
nand U1977 (N_1977,N_1325,N_1478);
and U1978 (N_1978,N_1392,N_1237);
or U1979 (N_1979,N_1377,N_1172);
xor U1980 (N_1980,N_1149,N_1400);
xor U1981 (N_1981,N_1483,N_1086);
nor U1982 (N_1982,N_1309,N_1179);
and U1983 (N_1983,N_1429,N_1042);
xor U1984 (N_1984,N_1246,N_1480);
nand U1985 (N_1985,N_1421,N_1310);
xor U1986 (N_1986,N_1321,N_1154);
xor U1987 (N_1987,N_1347,N_1314);
nor U1988 (N_1988,N_1489,N_1250);
xor U1989 (N_1989,N_1473,N_1404);
and U1990 (N_1990,N_1316,N_1412);
nand U1991 (N_1991,N_1049,N_1443);
nand U1992 (N_1992,N_1455,N_1383);
or U1993 (N_1993,N_1139,N_1250);
xnor U1994 (N_1994,N_1369,N_1062);
nand U1995 (N_1995,N_1307,N_1124);
and U1996 (N_1996,N_1041,N_1448);
nor U1997 (N_1997,N_1417,N_1441);
nor U1998 (N_1998,N_1438,N_1400);
nor U1999 (N_1999,N_1167,N_1430);
nor U2000 (N_2000,N_1802,N_1901);
or U2001 (N_2001,N_1669,N_1970);
or U2002 (N_2002,N_1830,N_1768);
xor U2003 (N_2003,N_1755,N_1639);
xor U2004 (N_2004,N_1825,N_1561);
nor U2005 (N_2005,N_1957,N_1573);
nand U2006 (N_2006,N_1935,N_1955);
xnor U2007 (N_2007,N_1542,N_1622);
xnor U2008 (N_2008,N_1878,N_1933);
xnor U2009 (N_2009,N_1869,N_1505);
nand U2010 (N_2010,N_1585,N_1983);
or U2011 (N_2011,N_1562,N_1555);
nor U2012 (N_2012,N_1579,N_1833);
and U2013 (N_2013,N_1919,N_1884);
and U2014 (N_2014,N_1532,N_1899);
or U2015 (N_2015,N_1740,N_1932);
xnor U2016 (N_2016,N_1984,N_1625);
nor U2017 (N_2017,N_1784,N_1868);
and U2018 (N_2018,N_1888,N_1920);
xnor U2019 (N_2019,N_1818,N_1671);
nand U2020 (N_2020,N_1862,N_1841);
or U2021 (N_2021,N_1670,N_1914);
nor U2022 (N_2022,N_1592,N_1891);
nor U2023 (N_2023,N_1599,N_1791);
and U2024 (N_2024,N_1857,N_1781);
and U2025 (N_2025,N_1769,N_1712);
xnor U2026 (N_2026,N_1780,N_1750);
nand U2027 (N_2027,N_1779,N_1703);
or U2028 (N_2028,N_1626,N_1500);
or U2029 (N_2029,N_1510,N_1597);
xnor U2030 (N_2030,N_1689,N_1913);
xnor U2031 (N_2031,N_1978,N_1649);
xor U2032 (N_2032,N_1591,N_1916);
nor U2033 (N_2033,N_1588,N_1745);
xnor U2034 (N_2034,N_1560,N_1654);
and U2035 (N_2035,N_1771,N_1726);
nor U2036 (N_2036,N_1600,N_1937);
and U2037 (N_2037,N_1509,N_1861);
and U2038 (N_2038,N_1507,N_1644);
or U2039 (N_2039,N_1679,N_1613);
nor U2040 (N_2040,N_1590,N_1722);
nand U2041 (N_2041,N_1981,N_1998);
and U2042 (N_2042,N_1986,N_1720);
nand U2043 (N_2043,N_1617,N_1821);
nor U2044 (N_2044,N_1690,N_1959);
and U2045 (N_2045,N_1807,N_1666);
or U2046 (N_2046,N_1525,N_1805);
nor U2047 (N_2047,N_1570,N_1814);
or U2048 (N_2048,N_1929,N_1820);
nand U2049 (N_2049,N_1554,N_1587);
xnor U2050 (N_2050,N_1876,N_1700);
nor U2051 (N_2051,N_1894,N_1730);
xnor U2052 (N_2052,N_1893,N_1607);
xor U2053 (N_2053,N_1871,N_1604);
and U2054 (N_2054,N_1902,N_1598);
nor U2055 (N_2055,N_1563,N_1971);
or U2056 (N_2056,N_1724,N_1685);
or U2057 (N_2057,N_1514,N_1708);
nand U2058 (N_2058,N_1503,N_1909);
xnor U2059 (N_2059,N_1832,N_1538);
xnor U2060 (N_2060,N_1774,N_1628);
xnor U2061 (N_2061,N_1886,N_1976);
nor U2062 (N_2062,N_1803,N_1875);
nor U2063 (N_2063,N_1918,N_1758);
or U2064 (N_2064,N_1898,N_1954);
nand U2065 (N_2065,N_1731,N_1760);
xor U2066 (N_2066,N_1537,N_1564);
nor U2067 (N_2067,N_1974,N_1668);
and U2068 (N_2068,N_1962,N_1522);
and U2069 (N_2069,N_1782,N_1698);
or U2070 (N_2070,N_1717,N_1808);
nor U2071 (N_2071,N_1797,N_1969);
xor U2072 (N_2072,N_1866,N_1867);
and U2073 (N_2073,N_1930,N_1855);
nand U2074 (N_2074,N_1879,N_1991);
xor U2075 (N_2075,N_1941,N_1860);
nor U2076 (N_2076,N_1578,N_1870);
and U2077 (N_2077,N_1544,N_1534);
nor U2078 (N_2078,N_1729,N_1580);
nand U2079 (N_2079,N_1925,N_1934);
nor U2080 (N_2080,N_1582,N_1952);
and U2081 (N_2081,N_1776,N_1743);
or U2082 (N_2082,N_1853,N_1519);
and U2083 (N_2083,N_1787,N_1765);
or U2084 (N_2084,N_1880,N_1695);
xnor U2085 (N_2085,N_1967,N_1754);
nand U2086 (N_2086,N_1852,N_1882);
xor U2087 (N_2087,N_1569,N_1912);
xor U2088 (N_2088,N_1546,N_1715);
xor U2089 (N_2089,N_1831,N_1517);
nand U2090 (N_2090,N_1718,N_1692);
or U2091 (N_2091,N_1602,N_1660);
or U2092 (N_2092,N_1535,N_1665);
xor U2093 (N_2093,N_1951,N_1516);
or U2094 (N_2094,N_1801,N_1611);
nor U2095 (N_2095,N_1848,N_1636);
xor U2096 (N_2096,N_1798,N_1647);
and U2097 (N_2097,N_1696,N_1761);
and U2098 (N_2098,N_1577,N_1748);
and U2099 (N_2099,N_1817,N_1789);
and U2100 (N_2100,N_1631,N_1683);
nand U2101 (N_2101,N_1742,N_1924);
nand U2102 (N_2102,N_1629,N_1550);
or U2103 (N_2103,N_1652,N_1872);
xor U2104 (N_2104,N_1594,N_1677);
nor U2105 (N_2105,N_1826,N_1975);
or U2106 (N_2106,N_1972,N_1586);
nand U2107 (N_2107,N_1711,N_1980);
and U2108 (N_2108,N_1908,N_1843);
nor U2109 (N_2109,N_1574,N_1645);
nand U2110 (N_2110,N_1827,N_1530);
xnor U2111 (N_2111,N_1713,N_1950);
nand U2112 (N_2112,N_1583,N_1557);
and U2113 (N_2113,N_1940,N_1896);
xnor U2114 (N_2114,N_1844,N_1783);
nor U2115 (N_2115,N_1630,N_1738);
or U2116 (N_2116,N_1620,N_1839);
or U2117 (N_2117,N_1744,N_1531);
nand U2118 (N_2118,N_1709,N_1721);
xor U2119 (N_2119,N_1863,N_1627);
nor U2120 (N_2120,N_1956,N_1526);
or U2121 (N_2121,N_1667,N_1949);
or U2122 (N_2122,N_1682,N_1567);
or U2123 (N_2123,N_1650,N_1850);
xnor U2124 (N_2124,N_1741,N_1606);
nor U2125 (N_2125,N_1751,N_1816);
nand U2126 (N_2126,N_1632,N_1800);
xor U2127 (N_2127,N_1999,N_1795);
nand U2128 (N_2128,N_1979,N_1566);
or U2129 (N_2129,N_1553,N_1746);
xnor U2130 (N_2130,N_1699,N_1887);
and U2131 (N_2131,N_1702,N_1985);
nor U2132 (N_2132,N_1788,N_1739);
nand U2133 (N_2133,N_1733,N_1958);
xor U2134 (N_2134,N_1838,N_1938);
nor U2135 (N_2135,N_1944,N_1549);
or U2136 (N_2136,N_1504,N_1885);
and U2137 (N_2137,N_1993,N_1813);
nor U2138 (N_2138,N_1736,N_1643);
or U2139 (N_2139,N_1523,N_1856);
or U2140 (N_2140,N_1551,N_1995);
xor U2141 (N_2141,N_1508,N_1704);
nand U2142 (N_2142,N_1656,N_1638);
nor U2143 (N_2143,N_1936,N_1524);
and U2144 (N_2144,N_1520,N_1637);
or U2145 (N_2145,N_1728,N_1928);
nand U2146 (N_2146,N_1996,N_1829);
or U2147 (N_2147,N_1911,N_1759);
nand U2148 (N_2148,N_1897,N_1994);
nand U2149 (N_2149,N_1877,N_1687);
and U2150 (N_2150,N_1697,N_1548);
or U2151 (N_2151,N_1904,N_1921);
xor U2152 (N_2152,N_1605,N_1595);
xor U2153 (N_2153,N_1786,N_1641);
nand U2154 (N_2154,N_1915,N_1710);
and U2155 (N_2155,N_1987,N_1533);
or U2156 (N_2156,N_1655,N_1714);
and U2157 (N_2157,N_1501,N_1942);
or U2158 (N_2158,N_1927,N_1757);
nand U2159 (N_2159,N_1865,N_1812);
or U2160 (N_2160,N_1939,N_1608);
or U2161 (N_2161,N_1662,N_1763);
nand U2162 (N_2162,N_1540,N_1640);
nand U2163 (N_2163,N_1559,N_1684);
nor U2164 (N_2164,N_1547,N_1545);
or U2165 (N_2165,N_1823,N_1905);
nand U2166 (N_2166,N_1778,N_1663);
nand U2167 (N_2167,N_1945,N_1633);
nor U2168 (N_2168,N_1571,N_1749);
xor U2169 (N_2169,N_1874,N_1576);
xor U2170 (N_2170,N_1646,N_1527);
or U2171 (N_2171,N_1601,N_1965);
and U2172 (N_2172,N_1809,N_1515);
and U2173 (N_2173,N_1661,N_1948);
and U2174 (N_2174,N_1926,N_1735);
nor U2175 (N_2175,N_1753,N_1794);
and U2176 (N_2176,N_1834,N_1734);
or U2177 (N_2177,N_1799,N_1552);
nor U2178 (N_2178,N_1943,N_1623);
or U2179 (N_2179,N_1614,N_1982);
xor U2180 (N_2180,N_1988,N_1737);
and U2181 (N_2181,N_1764,N_1790);
nand U2182 (N_2182,N_1845,N_1792);
or U2183 (N_2183,N_1997,N_1906);
nand U2184 (N_2184,N_1725,N_1811);
and U2185 (N_2185,N_1675,N_1858);
and U2186 (N_2186,N_1947,N_1881);
nand U2187 (N_2187,N_1681,N_1900);
nor U2188 (N_2188,N_1558,N_1989);
xnor U2189 (N_2189,N_1785,N_1873);
or U2190 (N_2190,N_1556,N_1946);
or U2191 (N_2191,N_1575,N_1851);
nor U2192 (N_2192,N_1716,N_1521);
xnor U2193 (N_2193,N_1973,N_1609);
xor U2194 (N_2194,N_1589,N_1634);
xor U2195 (N_2195,N_1766,N_1772);
nand U2196 (N_2196,N_1770,N_1543);
or U2197 (N_2197,N_1835,N_1892);
or U2198 (N_2198,N_1678,N_1664);
or U2199 (N_2199,N_1864,N_1992);
nand U2200 (N_2200,N_1842,N_1840);
or U2201 (N_2201,N_1635,N_1529);
nand U2202 (N_2202,N_1624,N_1732);
xnor U2203 (N_2203,N_1568,N_1694);
nor U2204 (N_2204,N_1931,N_1890);
nand U2205 (N_2205,N_1747,N_1806);
and U2206 (N_2206,N_1688,N_1658);
or U2207 (N_2207,N_1691,N_1966);
nor U2208 (N_2208,N_1565,N_1836);
xor U2209 (N_2209,N_1968,N_1651);
and U2210 (N_2210,N_1672,N_1593);
and U2211 (N_2211,N_1854,N_1777);
and U2212 (N_2212,N_1707,N_1964);
or U2213 (N_2213,N_1511,N_1701);
or U2214 (N_2214,N_1528,N_1512);
or U2215 (N_2215,N_1536,N_1773);
nand U2216 (N_2216,N_1706,N_1686);
nand U2217 (N_2217,N_1963,N_1917);
nand U2218 (N_2218,N_1796,N_1619);
nor U2219 (N_2219,N_1752,N_1847);
xnor U2220 (N_2220,N_1584,N_1596);
nand U2221 (N_2221,N_1775,N_1990);
and U2222 (N_2222,N_1615,N_1793);
nand U2223 (N_2223,N_1756,N_1603);
or U2224 (N_2224,N_1923,N_1616);
nor U2225 (N_2225,N_1903,N_1648);
or U2226 (N_2226,N_1506,N_1815);
and U2227 (N_2227,N_1889,N_1659);
and U2228 (N_2228,N_1621,N_1518);
xor U2229 (N_2229,N_1653,N_1705);
xor U2230 (N_2230,N_1977,N_1819);
and U2231 (N_2231,N_1910,N_1723);
xor U2232 (N_2232,N_1859,N_1539);
and U2233 (N_2233,N_1657,N_1719);
xor U2234 (N_2234,N_1676,N_1727);
nor U2235 (N_2235,N_1961,N_1572);
or U2236 (N_2236,N_1618,N_1849);
and U2237 (N_2237,N_1953,N_1846);
xor U2238 (N_2238,N_1502,N_1673);
and U2239 (N_2239,N_1822,N_1581);
and U2240 (N_2240,N_1883,N_1907);
nor U2241 (N_2241,N_1922,N_1837);
or U2242 (N_2242,N_1895,N_1810);
nand U2243 (N_2243,N_1642,N_1541);
and U2244 (N_2244,N_1674,N_1828);
nor U2245 (N_2245,N_1767,N_1960);
nor U2246 (N_2246,N_1804,N_1693);
and U2247 (N_2247,N_1824,N_1762);
and U2248 (N_2248,N_1610,N_1612);
xor U2249 (N_2249,N_1513,N_1680);
xnor U2250 (N_2250,N_1507,N_1907);
nor U2251 (N_2251,N_1705,N_1846);
xnor U2252 (N_2252,N_1703,N_1836);
xnor U2253 (N_2253,N_1678,N_1975);
xor U2254 (N_2254,N_1502,N_1525);
nor U2255 (N_2255,N_1543,N_1532);
nand U2256 (N_2256,N_1695,N_1928);
and U2257 (N_2257,N_1709,N_1808);
nor U2258 (N_2258,N_1604,N_1647);
or U2259 (N_2259,N_1810,N_1961);
or U2260 (N_2260,N_1512,N_1691);
and U2261 (N_2261,N_1597,N_1935);
or U2262 (N_2262,N_1823,N_1620);
nor U2263 (N_2263,N_1524,N_1680);
xor U2264 (N_2264,N_1756,N_1922);
xnor U2265 (N_2265,N_1856,N_1837);
or U2266 (N_2266,N_1831,N_1953);
nand U2267 (N_2267,N_1711,N_1844);
nor U2268 (N_2268,N_1733,N_1748);
or U2269 (N_2269,N_1950,N_1669);
or U2270 (N_2270,N_1840,N_1656);
xnor U2271 (N_2271,N_1941,N_1771);
nand U2272 (N_2272,N_1992,N_1530);
nand U2273 (N_2273,N_1648,N_1553);
nand U2274 (N_2274,N_1742,N_1986);
or U2275 (N_2275,N_1993,N_1829);
nand U2276 (N_2276,N_1528,N_1953);
nand U2277 (N_2277,N_1678,N_1803);
nand U2278 (N_2278,N_1793,N_1962);
xor U2279 (N_2279,N_1631,N_1519);
nor U2280 (N_2280,N_1987,N_1877);
and U2281 (N_2281,N_1989,N_1563);
nand U2282 (N_2282,N_1975,N_1547);
and U2283 (N_2283,N_1638,N_1886);
xor U2284 (N_2284,N_1833,N_1619);
nor U2285 (N_2285,N_1569,N_1822);
and U2286 (N_2286,N_1888,N_1881);
nand U2287 (N_2287,N_1757,N_1610);
or U2288 (N_2288,N_1864,N_1705);
xnor U2289 (N_2289,N_1924,N_1649);
and U2290 (N_2290,N_1804,N_1905);
nand U2291 (N_2291,N_1845,N_1678);
or U2292 (N_2292,N_1534,N_1838);
or U2293 (N_2293,N_1773,N_1552);
nor U2294 (N_2294,N_1518,N_1862);
nor U2295 (N_2295,N_1893,N_1634);
nor U2296 (N_2296,N_1891,N_1705);
nor U2297 (N_2297,N_1680,N_1663);
and U2298 (N_2298,N_1891,N_1816);
nand U2299 (N_2299,N_1856,N_1788);
and U2300 (N_2300,N_1986,N_1911);
nand U2301 (N_2301,N_1638,N_1648);
and U2302 (N_2302,N_1558,N_1784);
and U2303 (N_2303,N_1801,N_1797);
nor U2304 (N_2304,N_1624,N_1801);
and U2305 (N_2305,N_1547,N_1974);
and U2306 (N_2306,N_1734,N_1900);
nor U2307 (N_2307,N_1637,N_1631);
nor U2308 (N_2308,N_1921,N_1790);
xor U2309 (N_2309,N_1851,N_1742);
and U2310 (N_2310,N_1849,N_1948);
nand U2311 (N_2311,N_1718,N_1689);
or U2312 (N_2312,N_1669,N_1609);
xor U2313 (N_2313,N_1920,N_1638);
nand U2314 (N_2314,N_1650,N_1744);
nand U2315 (N_2315,N_1618,N_1944);
xor U2316 (N_2316,N_1503,N_1661);
xor U2317 (N_2317,N_1581,N_1599);
and U2318 (N_2318,N_1675,N_1708);
nand U2319 (N_2319,N_1833,N_1561);
nor U2320 (N_2320,N_1977,N_1947);
and U2321 (N_2321,N_1968,N_1625);
nand U2322 (N_2322,N_1690,N_1766);
xor U2323 (N_2323,N_1895,N_1510);
xor U2324 (N_2324,N_1544,N_1668);
or U2325 (N_2325,N_1581,N_1935);
xnor U2326 (N_2326,N_1864,N_1847);
nand U2327 (N_2327,N_1539,N_1695);
nor U2328 (N_2328,N_1983,N_1567);
and U2329 (N_2329,N_1699,N_1549);
and U2330 (N_2330,N_1650,N_1675);
and U2331 (N_2331,N_1714,N_1580);
nand U2332 (N_2332,N_1615,N_1655);
and U2333 (N_2333,N_1602,N_1794);
nor U2334 (N_2334,N_1597,N_1723);
or U2335 (N_2335,N_1511,N_1509);
nand U2336 (N_2336,N_1936,N_1593);
and U2337 (N_2337,N_1544,N_1609);
nand U2338 (N_2338,N_1889,N_1846);
nand U2339 (N_2339,N_1780,N_1638);
nor U2340 (N_2340,N_1970,N_1817);
nand U2341 (N_2341,N_1711,N_1900);
nor U2342 (N_2342,N_1587,N_1758);
xnor U2343 (N_2343,N_1840,N_1967);
nand U2344 (N_2344,N_1588,N_1778);
and U2345 (N_2345,N_1694,N_1717);
xnor U2346 (N_2346,N_1577,N_1977);
or U2347 (N_2347,N_1728,N_1749);
nor U2348 (N_2348,N_1959,N_1938);
and U2349 (N_2349,N_1587,N_1966);
xnor U2350 (N_2350,N_1603,N_1670);
nor U2351 (N_2351,N_1953,N_1703);
xnor U2352 (N_2352,N_1527,N_1520);
nor U2353 (N_2353,N_1742,N_1665);
or U2354 (N_2354,N_1730,N_1873);
nor U2355 (N_2355,N_1935,N_1921);
xnor U2356 (N_2356,N_1662,N_1669);
nor U2357 (N_2357,N_1932,N_1638);
and U2358 (N_2358,N_1510,N_1874);
and U2359 (N_2359,N_1807,N_1945);
xor U2360 (N_2360,N_1792,N_1559);
or U2361 (N_2361,N_1755,N_1972);
and U2362 (N_2362,N_1543,N_1853);
xor U2363 (N_2363,N_1736,N_1614);
and U2364 (N_2364,N_1977,N_1779);
or U2365 (N_2365,N_1938,N_1916);
and U2366 (N_2366,N_1608,N_1714);
nor U2367 (N_2367,N_1780,N_1711);
nor U2368 (N_2368,N_1900,N_1764);
and U2369 (N_2369,N_1712,N_1502);
and U2370 (N_2370,N_1763,N_1881);
nand U2371 (N_2371,N_1546,N_1587);
xor U2372 (N_2372,N_1522,N_1566);
nor U2373 (N_2373,N_1889,N_1626);
or U2374 (N_2374,N_1948,N_1622);
nand U2375 (N_2375,N_1504,N_1945);
and U2376 (N_2376,N_1703,N_1847);
nand U2377 (N_2377,N_1888,N_1908);
nor U2378 (N_2378,N_1949,N_1626);
or U2379 (N_2379,N_1579,N_1674);
or U2380 (N_2380,N_1614,N_1878);
nor U2381 (N_2381,N_1628,N_1671);
xor U2382 (N_2382,N_1777,N_1675);
xnor U2383 (N_2383,N_1578,N_1888);
and U2384 (N_2384,N_1507,N_1686);
nand U2385 (N_2385,N_1683,N_1607);
xor U2386 (N_2386,N_1745,N_1873);
or U2387 (N_2387,N_1820,N_1826);
nor U2388 (N_2388,N_1867,N_1885);
nor U2389 (N_2389,N_1662,N_1831);
and U2390 (N_2390,N_1871,N_1969);
nor U2391 (N_2391,N_1985,N_1790);
or U2392 (N_2392,N_1664,N_1622);
xor U2393 (N_2393,N_1516,N_1874);
xor U2394 (N_2394,N_1577,N_1883);
nand U2395 (N_2395,N_1945,N_1694);
and U2396 (N_2396,N_1855,N_1653);
and U2397 (N_2397,N_1553,N_1533);
and U2398 (N_2398,N_1535,N_1960);
nand U2399 (N_2399,N_1671,N_1807);
xnor U2400 (N_2400,N_1570,N_1532);
or U2401 (N_2401,N_1581,N_1943);
nor U2402 (N_2402,N_1554,N_1714);
or U2403 (N_2403,N_1722,N_1916);
nand U2404 (N_2404,N_1944,N_1787);
xnor U2405 (N_2405,N_1698,N_1789);
and U2406 (N_2406,N_1854,N_1864);
nand U2407 (N_2407,N_1729,N_1715);
nor U2408 (N_2408,N_1809,N_1545);
or U2409 (N_2409,N_1545,N_1720);
or U2410 (N_2410,N_1565,N_1532);
and U2411 (N_2411,N_1648,N_1603);
nor U2412 (N_2412,N_1750,N_1517);
nor U2413 (N_2413,N_1868,N_1598);
and U2414 (N_2414,N_1597,N_1904);
xor U2415 (N_2415,N_1681,N_1623);
and U2416 (N_2416,N_1897,N_1796);
or U2417 (N_2417,N_1584,N_1626);
and U2418 (N_2418,N_1512,N_1647);
nand U2419 (N_2419,N_1562,N_1783);
and U2420 (N_2420,N_1911,N_1520);
or U2421 (N_2421,N_1514,N_1618);
xor U2422 (N_2422,N_1796,N_1714);
xnor U2423 (N_2423,N_1667,N_1833);
or U2424 (N_2424,N_1895,N_1940);
and U2425 (N_2425,N_1781,N_1899);
nand U2426 (N_2426,N_1984,N_1594);
or U2427 (N_2427,N_1985,N_1521);
or U2428 (N_2428,N_1527,N_1725);
nor U2429 (N_2429,N_1923,N_1645);
and U2430 (N_2430,N_1822,N_1651);
and U2431 (N_2431,N_1599,N_1700);
nor U2432 (N_2432,N_1516,N_1721);
or U2433 (N_2433,N_1620,N_1829);
and U2434 (N_2434,N_1792,N_1843);
nor U2435 (N_2435,N_1755,N_1687);
and U2436 (N_2436,N_1764,N_1923);
or U2437 (N_2437,N_1971,N_1581);
xnor U2438 (N_2438,N_1854,N_1694);
and U2439 (N_2439,N_1949,N_1836);
nor U2440 (N_2440,N_1585,N_1504);
nor U2441 (N_2441,N_1969,N_1668);
nor U2442 (N_2442,N_1515,N_1847);
and U2443 (N_2443,N_1848,N_1918);
xor U2444 (N_2444,N_1807,N_1659);
nand U2445 (N_2445,N_1665,N_1834);
nand U2446 (N_2446,N_1900,N_1980);
xor U2447 (N_2447,N_1675,N_1985);
nor U2448 (N_2448,N_1599,N_1947);
nor U2449 (N_2449,N_1783,N_1606);
nor U2450 (N_2450,N_1736,N_1846);
xnor U2451 (N_2451,N_1684,N_1585);
nor U2452 (N_2452,N_1602,N_1775);
nand U2453 (N_2453,N_1991,N_1872);
xnor U2454 (N_2454,N_1801,N_1883);
nand U2455 (N_2455,N_1542,N_1793);
nand U2456 (N_2456,N_1882,N_1544);
and U2457 (N_2457,N_1808,N_1609);
xor U2458 (N_2458,N_1609,N_1934);
and U2459 (N_2459,N_1987,N_1658);
or U2460 (N_2460,N_1823,N_1533);
xnor U2461 (N_2461,N_1577,N_1575);
xor U2462 (N_2462,N_1688,N_1930);
xnor U2463 (N_2463,N_1807,N_1687);
and U2464 (N_2464,N_1735,N_1736);
xnor U2465 (N_2465,N_1894,N_1858);
nand U2466 (N_2466,N_1604,N_1948);
and U2467 (N_2467,N_1702,N_1619);
nand U2468 (N_2468,N_1683,N_1991);
nand U2469 (N_2469,N_1649,N_1712);
nor U2470 (N_2470,N_1653,N_1621);
and U2471 (N_2471,N_1668,N_1980);
xnor U2472 (N_2472,N_1704,N_1590);
or U2473 (N_2473,N_1626,N_1677);
xnor U2474 (N_2474,N_1659,N_1827);
or U2475 (N_2475,N_1579,N_1566);
or U2476 (N_2476,N_1553,N_1679);
xnor U2477 (N_2477,N_1551,N_1790);
and U2478 (N_2478,N_1751,N_1888);
xnor U2479 (N_2479,N_1874,N_1730);
and U2480 (N_2480,N_1874,N_1562);
nand U2481 (N_2481,N_1808,N_1525);
nor U2482 (N_2482,N_1615,N_1870);
nand U2483 (N_2483,N_1713,N_1721);
nand U2484 (N_2484,N_1643,N_1997);
or U2485 (N_2485,N_1880,N_1812);
xor U2486 (N_2486,N_1713,N_1760);
or U2487 (N_2487,N_1707,N_1518);
or U2488 (N_2488,N_1663,N_1888);
and U2489 (N_2489,N_1848,N_1712);
nand U2490 (N_2490,N_1856,N_1781);
nand U2491 (N_2491,N_1609,N_1616);
or U2492 (N_2492,N_1857,N_1827);
and U2493 (N_2493,N_1871,N_1869);
and U2494 (N_2494,N_1830,N_1725);
nand U2495 (N_2495,N_1611,N_1667);
nand U2496 (N_2496,N_1986,N_1719);
or U2497 (N_2497,N_1658,N_1941);
or U2498 (N_2498,N_1555,N_1932);
nand U2499 (N_2499,N_1885,N_1517);
and U2500 (N_2500,N_2145,N_2286);
or U2501 (N_2501,N_2116,N_2210);
xor U2502 (N_2502,N_2473,N_2250);
nor U2503 (N_2503,N_2403,N_2494);
and U2504 (N_2504,N_2127,N_2486);
xnor U2505 (N_2505,N_2090,N_2164);
or U2506 (N_2506,N_2226,N_2076);
xnor U2507 (N_2507,N_2008,N_2024);
and U2508 (N_2508,N_2374,N_2029);
nand U2509 (N_2509,N_2098,N_2153);
nor U2510 (N_2510,N_2327,N_2215);
and U2511 (N_2511,N_2357,N_2208);
xor U2512 (N_2512,N_2453,N_2430);
or U2513 (N_2513,N_2012,N_2368);
or U2514 (N_2514,N_2052,N_2310);
or U2515 (N_2515,N_2379,N_2092);
and U2516 (N_2516,N_2059,N_2365);
nand U2517 (N_2517,N_2172,N_2466);
nand U2518 (N_2518,N_2382,N_2235);
xnor U2519 (N_2519,N_2030,N_2221);
nand U2520 (N_2520,N_2497,N_2232);
and U2521 (N_2521,N_2114,N_2380);
and U2522 (N_2522,N_2271,N_2387);
xnor U2523 (N_2523,N_2077,N_2170);
or U2524 (N_2524,N_2465,N_2464);
xor U2525 (N_2525,N_2353,N_2418);
or U2526 (N_2526,N_2134,N_2176);
xnor U2527 (N_2527,N_2106,N_2407);
xor U2528 (N_2528,N_2456,N_2390);
or U2529 (N_2529,N_2443,N_2496);
or U2530 (N_2530,N_2230,N_2067);
and U2531 (N_2531,N_2213,N_2259);
xor U2532 (N_2532,N_2050,N_2202);
nor U2533 (N_2533,N_2332,N_2203);
nor U2534 (N_2534,N_2169,N_2243);
xor U2535 (N_2535,N_2180,N_2007);
nand U2536 (N_2536,N_2107,N_2450);
xnor U2537 (N_2537,N_2063,N_2436);
xor U2538 (N_2538,N_2483,N_2423);
nand U2539 (N_2539,N_2157,N_2140);
or U2540 (N_2540,N_2411,N_2001);
xor U2541 (N_2541,N_2046,N_2248);
xor U2542 (N_2542,N_2021,N_2476);
nor U2543 (N_2543,N_2425,N_2412);
nor U2544 (N_2544,N_2246,N_2254);
nand U2545 (N_2545,N_2378,N_2069);
or U2546 (N_2546,N_2424,N_2333);
and U2547 (N_2547,N_2178,N_2207);
and U2548 (N_2548,N_2071,N_2151);
nand U2549 (N_2549,N_2188,N_2343);
nor U2550 (N_2550,N_2081,N_2439);
nor U2551 (N_2551,N_2391,N_2272);
nand U2552 (N_2552,N_2319,N_2091);
nor U2553 (N_2553,N_2303,N_2110);
nand U2554 (N_2554,N_2014,N_2227);
nand U2555 (N_2555,N_2467,N_2020);
or U2556 (N_2556,N_2186,N_2233);
and U2557 (N_2557,N_2410,N_2335);
or U2558 (N_2558,N_2009,N_2371);
xor U2559 (N_2559,N_2237,N_2028);
or U2560 (N_2560,N_2426,N_2301);
nor U2561 (N_2561,N_2499,N_2452);
and U2562 (N_2562,N_2458,N_2193);
nor U2563 (N_2563,N_2179,N_2449);
nor U2564 (N_2564,N_2320,N_2209);
nor U2565 (N_2565,N_2428,N_2274);
nor U2566 (N_2566,N_2267,N_2204);
nand U2567 (N_2567,N_2468,N_2305);
nand U2568 (N_2568,N_2264,N_2370);
nand U2569 (N_2569,N_2137,N_2064);
nor U2570 (N_2570,N_2018,N_2057);
nand U2571 (N_2571,N_2032,N_2103);
xnor U2572 (N_2572,N_2401,N_2121);
and U2573 (N_2573,N_2461,N_2026);
nand U2574 (N_2574,N_2045,N_2108);
nand U2575 (N_2575,N_2437,N_2058);
or U2576 (N_2576,N_2404,N_2173);
nand U2577 (N_2577,N_2120,N_2493);
nand U2578 (N_2578,N_2212,N_2201);
xnor U2579 (N_2579,N_2383,N_2280);
or U2580 (N_2580,N_2276,N_2240);
and U2581 (N_2581,N_2396,N_2068);
or U2582 (N_2582,N_2073,N_2054);
and U2583 (N_2583,N_2150,N_2220);
and U2584 (N_2584,N_2298,N_2119);
nand U2585 (N_2585,N_2460,N_2448);
or U2586 (N_2586,N_2457,N_2435);
and U2587 (N_2587,N_2102,N_2263);
or U2588 (N_2588,N_2080,N_2388);
xor U2589 (N_2589,N_2031,N_2469);
or U2590 (N_2590,N_2147,N_2287);
or U2591 (N_2591,N_2075,N_2495);
or U2592 (N_2592,N_2013,N_2115);
or U2593 (N_2593,N_2345,N_2347);
nand U2594 (N_2594,N_2002,N_2109);
nand U2595 (N_2595,N_2143,N_2060);
and U2596 (N_2596,N_2366,N_2348);
and U2597 (N_2597,N_2163,N_2277);
or U2598 (N_2598,N_2440,N_2189);
or U2599 (N_2599,N_2405,N_2249);
or U2600 (N_2600,N_2022,N_2268);
and U2601 (N_2601,N_2384,N_2329);
or U2602 (N_2602,N_2346,N_2089);
or U2603 (N_2603,N_2304,N_2218);
nor U2604 (N_2604,N_2341,N_2487);
xor U2605 (N_2605,N_2400,N_2300);
nand U2606 (N_2606,N_2048,N_2442);
xnor U2607 (N_2607,N_2043,N_2123);
and U2608 (N_2608,N_2491,N_2217);
or U2609 (N_2609,N_2314,N_2372);
or U2610 (N_2610,N_2344,N_2244);
nor U2611 (N_2611,N_2385,N_2182);
or U2612 (N_2612,N_2299,N_2142);
nor U2613 (N_2613,N_2196,N_2222);
xor U2614 (N_2614,N_2125,N_2402);
nor U2615 (N_2615,N_2006,N_2283);
and U2616 (N_2616,N_2431,N_2165);
nand U2617 (N_2617,N_2459,N_2255);
or U2618 (N_2618,N_2337,N_2160);
nor U2619 (N_2619,N_2105,N_2079);
and U2620 (N_2620,N_2262,N_2141);
nand U2621 (N_2621,N_2036,N_2311);
or U2622 (N_2622,N_2242,N_2434);
and U2623 (N_2623,N_2392,N_2354);
nand U2624 (N_2624,N_2490,N_2306);
nor U2625 (N_2625,N_2148,N_2085);
and U2626 (N_2626,N_2338,N_2138);
or U2627 (N_2627,N_2482,N_2433);
nor U2628 (N_2628,N_2316,N_2214);
nor U2629 (N_2629,N_2313,N_2185);
xnor U2630 (N_2630,N_2463,N_2399);
xor U2631 (N_2631,N_2289,N_2190);
nor U2632 (N_2632,N_2016,N_2111);
xnor U2633 (N_2633,N_2023,N_2297);
or U2634 (N_2634,N_2187,N_2270);
and U2635 (N_2635,N_2238,N_2133);
or U2636 (N_2636,N_2168,N_2011);
and U2637 (N_2637,N_2038,N_2062);
nand U2638 (N_2638,N_2219,N_2295);
and U2639 (N_2639,N_2285,N_2171);
xor U2640 (N_2640,N_2393,N_2361);
nor U2641 (N_2641,N_2154,N_2290);
or U2642 (N_2642,N_2447,N_2231);
or U2643 (N_2643,N_2136,N_2397);
nand U2644 (N_2644,N_2416,N_2088);
nand U2645 (N_2645,N_2258,N_2377);
and U2646 (N_2646,N_2471,N_2409);
nor U2647 (N_2647,N_2129,N_2158);
xnor U2648 (N_2648,N_2236,N_2275);
nor U2649 (N_2649,N_2177,N_2003);
nand U2650 (N_2650,N_2083,N_2192);
or U2651 (N_2651,N_2175,N_2294);
xor U2652 (N_2652,N_2200,N_2478);
or U2653 (N_2653,N_2017,N_2099);
or U2654 (N_2654,N_2122,N_2094);
xnor U2655 (N_2655,N_2161,N_2315);
and U2656 (N_2656,N_2144,N_2135);
xor U2657 (N_2657,N_2369,N_2454);
and U2658 (N_2658,N_2049,N_2095);
nand U2659 (N_2659,N_2113,N_2253);
xnor U2660 (N_2660,N_2441,N_2056);
nor U2661 (N_2661,N_2066,N_2162);
xnor U2662 (N_2662,N_2166,N_2395);
xnor U2663 (N_2663,N_2257,N_2093);
and U2664 (N_2664,N_2055,N_2130);
and U2665 (N_2665,N_2475,N_2037);
nand U2666 (N_2666,N_2398,N_2061);
nand U2667 (N_2667,N_2477,N_2472);
or U2668 (N_2668,N_2317,N_2184);
nand U2669 (N_2669,N_2307,N_2100);
nor U2670 (N_2670,N_2474,N_2406);
nand U2671 (N_2671,N_2413,N_2118);
nor U2672 (N_2672,N_2096,N_2330);
nor U2673 (N_2673,N_2375,N_2389);
or U2674 (N_2674,N_2070,N_2010);
xnor U2675 (N_2675,N_2223,N_2386);
xnor U2676 (N_2676,N_2376,N_2101);
nor U2677 (N_2677,N_2041,N_2211);
or U2678 (N_2678,N_2360,N_2446);
nor U2679 (N_2679,N_2322,N_2266);
nor U2680 (N_2680,N_2252,N_2342);
or U2681 (N_2681,N_2117,N_2381);
or U2682 (N_2682,N_2191,N_2362);
nand U2683 (N_2683,N_2027,N_2097);
nand U2684 (N_2684,N_2181,N_2084);
nand U2685 (N_2685,N_2336,N_2429);
nor U2686 (N_2686,N_2086,N_2451);
nand U2687 (N_2687,N_2216,N_2183);
xnor U2688 (N_2688,N_2005,N_2364);
xnor U2689 (N_2689,N_2205,N_2308);
nand U2690 (N_2690,N_2131,N_2149);
nand U2691 (N_2691,N_2174,N_2312);
or U2692 (N_2692,N_2078,N_2195);
and U2693 (N_2693,N_2245,N_2112);
xor U2694 (N_2694,N_2194,N_2321);
or U2695 (N_2695,N_2485,N_2481);
nor U2696 (N_2696,N_2355,N_2044);
or U2697 (N_2697,N_2489,N_2082);
or U2698 (N_2698,N_2484,N_2488);
and U2699 (N_2699,N_2065,N_2087);
nand U2700 (N_2700,N_2128,N_2273);
nand U2701 (N_2701,N_2318,N_2265);
nor U2702 (N_2702,N_2394,N_2039);
nand U2703 (N_2703,N_2225,N_2198);
nand U2704 (N_2704,N_2349,N_2234);
and U2705 (N_2705,N_2291,N_2139);
xor U2706 (N_2706,N_2260,N_2278);
nor U2707 (N_2707,N_2373,N_2480);
or U2708 (N_2708,N_2419,N_2241);
nand U2709 (N_2709,N_2339,N_2279);
xnor U2710 (N_2710,N_2156,N_2296);
or U2711 (N_2711,N_2053,N_2000);
xnor U2712 (N_2712,N_2051,N_2229);
or U2713 (N_2713,N_2159,N_2199);
and U2714 (N_2714,N_2197,N_2422);
nand U2715 (N_2715,N_2025,N_2438);
or U2716 (N_2716,N_2356,N_2146);
and U2717 (N_2717,N_2309,N_2358);
xnor U2718 (N_2718,N_2256,N_2417);
nor U2719 (N_2719,N_2019,N_2293);
nand U2720 (N_2720,N_2126,N_2334);
nand U2721 (N_2721,N_2152,N_2479);
nand U2722 (N_2722,N_2074,N_2206);
or U2723 (N_2723,N_2340,N_2420);
and U2724 (N_2724,N_2352,N_2363);
xnor U2725 (N_2725,N_2167,N_2492);
or U2726 (N_2726,N_2033,N_2445);
xor U2727 (N_2727,N_2034,N_2324);
nor U2728 (N_2728,N_2155,N_2247);
or U2729 (N_2729,N_2421,N_2015);
nor U2730 (N_2730,N_2004,N_2132);
nand U2731 (N_2731,N_2408,N_2331);
xor U2732 (N_2732,N_2284,N_2415);
or U2733 (N_2733,N_2282,N_2498);
and U2734 (N_2734,N_2228,N_2326);
nor U2735 (N_2735,N_2325,N_2288);
and U2736 (N_2736,N_2261,N_2328);
and U2737 (N_2737,N_2444,N_2224);
or U2738 (N_2738,N_2367,N_2104);
nand U2739 (N_2739,N_2455,N_2462);
or U2740 (N_2740,N_2414,N_2269);
nand U2741 (N_2741,N_2351,N_2040);
nand U2742 (N_2742,N_2350,N_2359);
and U2743 (N_2743,N_2239,N_2323);
nand U2744 (N_2744,N_2042,N_2281);
nand U2745 (N_2745,N_2432,N_2427);
or U2746 (N_2746,N_2072,N_2302);
and U2747 (N_2747,N_2251,N_2047);
or U2748 (N_2748,N_2124,N_2292);
nor U2749 (N_2749,N_2470,N_2035);
nor U2750 (N_2750,N_2045,N_2313);
xnor U2751 (N_2751,N_2110,N_2483);
xor U2752 (N_2752,N_2141,N_2286);
nor U2753 (N_2753,N_2109,N_2352);
or U2754 (N_2754,N_2306,N_2489);
xnor U2755 (N_2755,N_2244,N_2023);
nor U2756 (N_2756,N_2315,N_2178);
nor U2757 (N_2757,N_2099,N_2493);
nor U2758 (N_2758,N_2190,N_2435);
and U2759 (N_2759,N_2297,N_2106);
nor U2760 (N_2760,N_2385,N_2132);
xnor U2761 (N_2761,N_2466,N_2139);
xnor U2762 (N_2762,N_2335,N_2318);
and U2763 (N_2763,N_2132,N_2361);
nand U2764 (N_2764,N_2111,N_2265);
xor U2765 (N_2765,N_2117,N_2092);
xor U2766 (N_2766,N_2327,N_2117);
and U2767 (N_2767,N_2298,N_2054);
nor U2768 (N_2768,N_2483,N_2033);
or U2769 (N_2769,N_2267,N_2348);
xnor U2770 (N_2770,N_2275,N_2332);
or U2771 (N_2771,N_2220,N_2061);
or U2772 (N_2772,N_2408,N_2207);
xor U2773 (N_2773,N_2029,N_2289);
nand U2774 (N_2774,N_2462,N_2250);
or U2775 (N_2775,N_2118,N_2293);
and U2776 (N_2776,N_2007,N_2328);
or U2777 (N_2777,N_2240,N_2119);
xnor U2778 (N_2778,N_2149,N_2181);
nor U2779 (N_2779,N_2241,N_2160);
or U2780 (N_2780,N_2193,N_2482);
and U2781 (N_2781,N_2471,N_2477);
or U2782 (N_2782,N_2272,N_2430);
and U2783 (N_2783,N_2459,N_2332);
nor U2784 (N_2784,N_2010,N_2034);
xor U2785 (N_2785,N_2348,N_2227);
nand U2786 (N_2786,N_2247,N_2328);
or U2787 (N_2787,N_2493,N_2405);
xnor U2788 (N_2788,N_2257,N_2361);
nand U2789 (N_2789,N_2064,N_2213);
nor U2790 (N_2790,N_2158,N_2009);
xnor U2791 (N_2791,N_2473,N_2134);
xnor U2792 (N_2792,N_2032,N_2064);
nand U2793 (N_2793,N_2317,N_2186);
nand U2794 (N_2794,N_2352,N_2019);
xor U2795 (N_2795,N_2456,N_2082);
and U2796 (N_2796,N_2039,N_2041);
or U2797 (N_2797,N_2403,N_2242);
xnor U2798 (N_2798,N_2435,N_2347);
nand U2799 (N_2799,N_2346,N_2132);
or U2800 (N_2800,N_2146,N_2157);
and U2801 (N_2801,N_2047,N_2120);
and U2802 (N_2802,N_2323,N_2302);
and U2803 (N_2803,N_2372,N_2435);
or U2804 (N_2804,N_2379,N_2447);
or U2805 (N_2805,N_2177,N_2295);
nor U2806 (N_2806,N_2342,N_2109);
xor U2807 (N_2807,N_2009,N_2377);
and U2808 (N_2808,N_2377,N_2059);
and U2809 (N_2809,N_2328,N_2211);
xor U2810 (N_2810,N_2266,N_2031);
xnor U2811 (N_2811,N_2029,N_2121);
nor U2812 (N_2812,N_2110,N_2306);
nand U2813 (N_2813,N_2028,N_2276);
nor U2814 (N_2814,N_2407,N_2297);
nand U2815 (N_2815,N_2381,N_2230);
and U2816 (N_2816,N_2202,N_2485);
nand U2817 (N_2817,N_2028,N_2293);
and U2818 (N_2818,N_2480,N_2000);
nand U2819 (N_2819,N_2039,N_2422);
nand U2820 (N_2820,N_2392,N_2341);
nand U2821 (N_2821,N_2472,N_2045);
nor U2822 (N_2822,N_2231,N_2052);
and U2823 (N_2823,N_2477,N_2425);
xor U2824 (N_2824,N_2398,N_2287);
xnor U2825 (N_2825,N_2076,N_2252);
xor U2826 (N_2826,N_2096,N_2288);
nor U2827 (N_2827,N_2195,N_2247);
and U2828 (N_2828,N_2153,N_2372);
or U2829 (N_2829,N_2408,N_2462);
xnor U2830 (N_2830,N_2476,N_2497);
or U2831 (N_2831,N_2167,N_2439);
and U2832 (N_2832,N_2465,N_2440);
nor U2833 (N_2833,N_2055,N_2358);
nand U2834 (N_2834,N_2262,N_2154);
or U2835 (N_2835,N_2426,N_2181);
and U2836 (N_2836,N_2394,N_2376);
and U2837 (N_2837,N_2405,N_2228);
nor U2838 (N_2838,N_2063,N_2458);
and U2839 (N_2839,N_2077,N_2221);
nor U2840 (N_2840,N_2030,N_2427);
xor U2841 (N_2841,N_2324,N_2379);
xnor U2842 (N_2842,N_2465,N_2458);
or U2843 (N_2843,N_2403,N_2456);
or U2844 (N_2844,N_2379,N_2180);
nand U2845 (N_2845,N_2112,N_2162);
nor U2846 (N_2846,N_2345,N_2161);
nand U2847 (N_2847,N_2347,N_2354);
or U2848 (N_2848,N_2419,N_2200);
and U2849 (N_2849,N_2326,N_2394);
xnor U2850 (N_2850,N_2356,N_2262);
and U2851 (N_2851,N_2295,N_2149);
xor U2852 (N_2852,N_2186,N_2465);
nor U2853 (N_2853,N_2311,N_2077);
and U2854 (N_2854,N_2443,N_2420);
nand U2855 (N_2855,N_2343,N_2217);
nand U2856 (N_2856,N_2264,N_2081);
nand U2857 (N_2857,N_2082,N_2441);
nor U2858 (N_2858,N_2019,N_2111);
nor U2859 (N_2859,N_2261,N_2372);
or U2860 (N_2860,N_2271,N_2033);
xor U2861 (N_2861,N_2458,N_2417);
or U2862 (N_2862,N_2444,N_2155);
nand U2863 (N_2863,N_2424,N_2431);
xnor U2864 (N_2864,N_2262,N_2145);
or U2865 (N_2865,N_2320,N_2051);
xor U2866 (N_2866,N_2224,N_2435);
and U2867 (N_2867,N_2376,N_2065);
or U2868 (N_2868,N_2419,N_2267);
nor U2869 (N_2869,N_2338,N_2478);
nor U2870 (N_2870,N_2035,N_2234);
and U2871 (N_2871,N_2060,N_2353);
or U2872 (N_2872,N_2277,N_2028);
and U2873 (N_2873,N_2073,N_2011);
and U2874 (N_2874,N_2433,N_2173);
and U2875 (N_2875,N_2272,N_2264);
or U2876 (N_2876,N_2120,N_2293);
nor U2877 (N_2877,N_2253,N_2345);
nand U2878 (N_2878,N_2079,N_2340);
or U2879 (N_2879,N_2059,N_2391);
and U2880 (N_2880,N_2345,N_2223);
or U2881 (N_2881,N_2060,N_2492);
and U2882 (N_2882,N_2043,N_2448);
xnor U2883 (N_2883,N_2099,N_2083);
nor U2884 (N_2884,N_2195,N_2414);
nand U2885 (N_2885,N_2273,N_2091);
xnor U2886 (N_2886,N_2440,N_2172);
nand U2887 (N_2887,N_2401,N_2266);
nand U2888 (N_2888,N_2428,N_2334);
nand U2889 (N_2889,N_2073,N_2124);
xor U2890 (N_2890,N_2438,N_2434);
nand U2891 (N_2891,N_2379,N_2046);
nor U2892 (N_2892,N_2392,N_2251);
and U2893 (N_2893,N_2465,N_2269);
nand U2894 (N_2894,N_2110,N_2258);
or U2895 (N_2895,N_2322,N_2499);
and U2896 (N_2896,N_2207,N_2001);
nor U2897 (N_2897,N_2273,N_2349);
and U2898 (N_2898,N_2332,N_2330);
nor U2899 (N_2899,N_2141,N_2006);
xor U2900 (N_2900,N_2034,N_2486);
or U2901 (N_2901,N_2088,N_2379);
nor U2902 (N_2902,N_2242,N_2377);
or U2903 (N_2903,N_2288,N_2350);
or U2904 (N_2904,N_2152,N_2278);
or U2905 (N_2905,N_2362,N_2101);
xor U2906 (N_2906,N_2041,N_2348);
nor U2907 (N_2907,N_2409,N_2185);
xor U2908 (N_2908,N_2356,N_2275);
nand U2909 (N_2909,N_2170,N_2432);
or U2910 (N_2910,N_2269,N_2439);
xor U2911 (N_2911,N_2260,N_2231);
nor U2912 (N_2912,N_2236,N_2062);
or U2913 (N_2913,N_2472,N_2385);
nand U2914 (N_2914,N_2009,N_2036);
or U2915 (N_2915,N_2063,N_2260);
or U2916 (N_2916,N_2212,N_2221);
and U2917 (N_2917,N_2138,N_2179);
xor U2918 (N_2918,N_2367,N_2106);
nor U2919 (N_2919,N_2264,N_2166);
nor U2920 (N_2920,N_2035,N_2265);
xnor U2921 (N_2921,N_2332,N_2326);
nor U2922 (N_2922,N_2206,N_2128);
nor U2923 (N_2923,N_2398,N_2351);
and U2924 (N_2924,N_2279,N_2427);
nor U2925 (N_2925,N_2176,N_2497);
xnor U2926 (N_2926,N_2266,N_2335);
and U2927 (N_2927,N_2301,N_2195);
xnor U2928 (N_2928,N_2047,N_2289);
nor U2929 (N_2929,N_2120,N_2177);
and U2930 (N_2930,N_2091,N_2139);
and U2931 (N_2931,N_2167,N_2320);
xnor U2932 (N_2932,N_2357,N_2156);
nor U2933 (N_2933,N_2231,N_2163);
nor U2934 (N_2934,N_2497,N_2048);
xnor U2935 (N_2935,N_2347,N_2488);
and U2936 (N_2936,N_2021,N_2213);
and U2937 (N_2937,N_2244,N_2289);
nor U2938 (N_2938,N_2256,N_2423);
nor U2939 (N_2939,N_2001,N_2028);
nor U2940 (N_2940,N_2210,N_2045);
and U2941 (N_2941,N_2333,N_2384);
nand U2942 (N_2942,N_2449,N_2413);
or U2943 (N_2943,N_2016,N_2446);
and U2944 (N_2944,N_2066,N_2086);
nor U2945 (N_2945,N_2259,N_2372);
and U2946 (N_2946,N_2366,N_2363);
nand U2947 (N_2947,N_2128,N_2160);
or U2948 (N_2948,N_2394,N_2340);
xor U2949 (N_2949,N_2375,N_2326);
or U2950 (N_2950,N_2259,N_2201);
xnor U2951 (N_2951,N_2261,N_2475);
xnor U2952 (N_2952,N_2342,N_2485);
xor U2953 (N_2953,N_2238,N_2318);
xor U2954 (N_2954,N_2475,N_2296);
nor U2955 (N_2955,N_2486,N_2196);
and U2956 (N_2956,N_2214,N_2157);
nand U2957 (N_2957,N_2065,N_2107);
nand U2958 (N_2958,N_2191,N_2399);
and U2959 (N_2959,N_2005,N_2362);
nand U2960 (N_2960,N_2296,N_2083);
and U2961 (N_2961,N_2139,N_2342);
nand U2962 (N_2962,N_2334,N_2201);
nor U2963 (N_2963,N_2097,N_2205);
xor U2964 (N_2964,N_2079,N_2158);
nor U2965 (N_2965,N_2230,N_2294);
nand U2966 (N_2966,N_2276,N_2262);
xnor U2967 (N_2967,N_2215,N_2232);
nor U2968 (N_2968,N_2360,N_2295);
or U2969 (N_2969,N_2326,N_2468);
and U2970 (N_2970,N_2190,N_2141);
and U2971 (N_2971,N_2107,N_2056);
nor U2972 (N_2972,N_2406,N_2479);
or U2973 (N_2973,N_2353,N_2141);
xnor U2974 (N_2974,N_2304,N_2431);
nor U2975 (N_2975,N_2383,N_2282);
and U2976 (N_2976,N_2180,N_2001);
nor U2977 (N_2977,N_2147,N_2326);
or U2978 (N_2978,N_2400,N_2287);
xor U2979 (N_2979,N_2121,N_2164);
xnor U2980 (N_2980,N_2140,N_2223);
or U2981 (N_2981,N_2065,N_2289);
xor U2982 (N_2982,N_2465,N_2313);
nand U2983 (N_2983,N_2172,N_2344);
or U2984 (N_2984,N_2279,N_2036);
or U2985 (N_2985,N_2172,N_2176);
or U2986 (N_2986,N_2021,N_2100);
nor U2987 (N_2987,N_2466,N_2234);
nand U2988 (N_2988,N_2488,N_2144);
or U2989 (N_2989,N_2227,N_2060);
nor U2990 (N_2990,N_2330,N_2457);
or U2991 (N_2991,N_2326,N_2417);
and U2992 (N_2992,N_2122,N_2079);
nor U2993 (N_2993,N_2046,N_2324);
and U2994 (N_2994,N_2320,N_2436);
nand U2995 (N_2995,N_2088,N_2256);
nand U2996 (N_2996,N_2269,N_2015);
nand U2997 (N_2997,N_2352,N_2406);
and U2998 (N_2998,N_2323,N_2240);
nand U2999 (N_2999,N_2207,N_2069);
or U3000 (N_3000,N_2540,N_2920);
nor U3001 (N_3001,N_2564,N_2940);
and U3002 (N_3002,N_2896,N_2771);
nand U3003 (N_3003,N_2763,N_2908);
and U3004 (N_3004,N_2938,N_2834);
and U3005 (N_3005,N_2934,N_2755);
nand U3006 (N_3006,N_2904,N_2567);
and U3007 (N_3007,N_2827,N_2963);
nand U3008 (N_3008,N_2628,N_2669);
or U3009 (N_3009,N_2914,N_2508);
xnor U3010 (N_3010,N_2910,N_2792);
nor U3011 (N_3011,N_2525,N_2702);
xnor U3012 (N_3012,N_2560,N_2593);
nand U3013 (N_3013,N_2521,N_2821);
and U3014 (N_3014,N_2987,N_2616);
nand U3015 (N_3015,N_2740,N_2909);
xnor U3016 (N_3016,N_2955,N_2655);
or U3017 (N_3017,N_2637,N_2966);
or U3018 (N_3018,N_2681,N_2583);
nand U3019 (N_3019,N_2667,N_2603);
nand U3020 (N_3020,N_2953,N_2861);
or U3021 (N_3021,N_2836,N_2777);
or U3022 (N_3022,N_2986,N_2787);
nand U3023 (N_3023,N_2510,N_2585);
or U3024 (N_3024,N_2766,N_2578);
and U3025 (N_3025,N_2846,N_2634);
and U3026 (N_3026,N_2710,N_2964);
and U3027 (N_3027,N_2544,N_2689);
xor U3028 (N_3028,N_2644,N_2847);
and U3029 (N_3029,N_2725,N_2588);
nand U3030 (N_3030,N_2767,N_2942);
xor U3031 (N_3031,N_2842,N_2611);
nand U3032 (N_3032,N_2607,N_2675);
and U3033 (N_3033,N_2780,N_2784);
nand U3034 (N_3034,N_2595,N_2992);
and U3035 (N_3035,N_2706,N_2608);
xnor U3036 (N_3036,N_2764,N_2793);
xor U3037 (N_3037,N_2639,N_2811);
xnor U3038 (N_3038,N_2994,N_2860);
nor U3039 (N_3039,N_2885,N_2712);
and U3040 (N_3040,N_2800,N_2517);
nand U3041 (N_3041,N_2529,N_2858);
nor U3042 (N_3042,N_2527,N_2519);
nor U3043 (N_3043,N_2602,N_2956);
and U3044 (N_3044,N_2946,N_2817);
xnor U3045 (N_3045,N_2818,N_2636);
or U3046 (N_3046,N_2932,N_2654);
nand U3047 (N_3047,N_2633,N_2918);
nor U3048 (N_3048,N_2900,N_2622);
and U3049 (N_3049,N_2822,N_2664);
and U3050 (N_3050,N_2586,N_2795);
xnor U3051 (N_3051,N_2699,N_2548);
and U3052 (N_3052,N_2625,N_2516);
nand U3053 (N_3053,N_2748,N_2754);
nor U3054 (N_3054,N_2627,N_2899);
nor U3055 (N_3055,N_2666,N_2980);
nor U3056 (N_3056,N_2883,N_2974);
or U3057 (N_3057,N_2645,N_2785);
xnor U3058 (N_3058,N_2662,N_2761);
nand U3059 (N_3059,N_2514,N_2684);
xor U3060 (N_3060,N_2572,N_2647);
nor U3061 (N_3061,N_2686,N_2976);
and U3062 (N_3062,N_2897,N_2906);
or U3063 (N_3063,N_2709,N_2642);
xor U3064 (N_3064,N_2977,N_2503);
xor U3065 (N_3065,N_2965,N_2750);
xnor U3066 (N_3066,N_2786,N_2804);
xnor U3067 (N_3067,N_2659,N_2923);
nor U3068 (N_3068,N_2889,N_2555);
nor U3069 (N_3069,N_2687,N_2872);
xor U3070 (N_3070,N_2613,N_2879);
nand U3071 (N_3071,N_2797,N_2794);
and U3072 (N_3072,N_2682,N_2554);
nor U3073 (N_3073,N_2531,N_2762);
nor U3074 (N_3074,N_2704,N_2758);
or U3075 (N_3075,N_2500,N_2988);
nor U3076 (N_3076,N_2577,N_2542);
nand U3077 (N_3077,N_2550,N_2851);
or U3078 (N_3078,N_2590,N_2913);
xor U3079 (N_3079,N_2968,N_2925);
and U3080 (N_3080,N_2535,N_2806);
or U3081 (N_3081,N_2975,N_2971);
nor U3082 (N_3082,N_2703,N_2892);
nand U3083 (N_3083,N_2638,N_2957);
nand U3084 (N_3084,N_2632,N_2753);
and U3085 (N_3085,N_2856,N_2717);
nand U3086 (N_3086,N_2715,N_2587);
or U3087 (N_3087,N_2926,N_2594);
nand U3088 (N_3088,N_2640,N_2835);
or U3089 (N_3089,N_2618,N_2573);
xnor U3090 (N_3090,N_2841,N_2930);
or U3091 (N_3091,N_2837,N_2924);
and U3092 (N_3092,N_2781,N_2803);
or U3093 (N_3093,N_2562,N_2936);
xor U3094 (N_3094,N_2949,N_2522);
or U3095 (N_3095,N_2808,N_2597);
nand U3096 (N_3096,N_2958,N_2770);
xor U3097 (N_3097,N_2657,N_2724);
and U3098 (N_3098,N_2919,N_2893);
or U3099 (N_3099,N_2504,N_2671);
or U3100 (N_3100,N_2996,N_2759);
and U3101 (N_3101,N_2502,N_2673);
or U3102 (N_3102,N_2849,N_2839);
or U3103 (N_3103,N_2898,N_2871);
or U3104 (N_3104,N_2576,N_2511);
or U3105 (N_3105,N_2912,N_2962);
xnor U3106 (N_3106,N_2937,N_2944);
and U3107 (N_3107,N_2928,N_2723);
nand U3108 (N_3108,N_2850,N_2814);
and U3109 (N_3109,N_2870,N_2840);
nand U3110 (N_3110,N_2538,N_2716);
nand U3111 (N_3111,N_2782,N_2737);
and U3112 (N_3112,N_2545,N_2624);
or U3113 (N_3113,N_2886,N_2742);
nor U3114 (N_3114,N_2981,N_2729);
nor U3115 (N_3115,N_2697,N_2884);
nand U3116 (N_3116,N_2894,N_2609);
nand U3117 (N_3117,N_2549,N_2990);
nand U3118 (N_3118,N_2660,N_2863);
xnor U3119 (N_3119,N_2679,N_2751);
nand U3120 (N_3120,N_2880,N_2907);
or U3121 (N_3121,N_2619,N_2816);
or U3122 (N_3122,N_2776,N_2713);
and U3123 (N_3123,N_2700,N_2739);
and U3124 (N_3124,N_2789,N_2552);
and U3125 (N_3125,N_2999,N_2783);
nor U3126 (N_3126,N_2569,N_2695);
and U3127 (N_3127,N_2959,N_2825);
and U3128 (N_3128,N_2623,N_2929);
nor U3129 (N_3129,N_2635,N_2888);
and U3130 (N_3130,N_2604,N_2612);
nand U3131 (N_3131,N_2556,N_2916);
nand U3132 (N_3132,N_2891,N_2580);
nand U3133 (N_3133,N_2939,N_2969);
xor U3134 (N_3134,N_2997,N_2546);
and U3135 (N_3135,N_2651,N_2558);
and U3136 (N_3136,N_2512,N_2813);
nor U3137 (N_3137,N_2905,N_2857);
nor U3138 (N_3138,N_2769,N_2553);
and U3139 (N_3139,N_2539,N_2757);
nand U3140 (N_3140,N_2855,N_2665);
nand U3141 (N_3141,N_2656,N_2967);
xnor U3142 (N_3142,N_2668,N_2887);
xor U3143 (N_3143,N_2532,N_2534);
nor U3144 (N_3144,N_2756,N_2678);
nor U3145 (N_3145,N_2674,N_2917);
xnor U3146 (N_3146,N_2582,N_2993);
xor U3147 (N_3147,N_2945,N_2864);
and U3148 (N_3148,N_2952,N_2865);
nand U3149 (N_3149,N_2829,N_2985);
or U3150 (N_3150,N_2747,N_2693);
nand U3151 (N_3151,N_2903,N_2960);
xor U3152 (N_3152,N_2833,N_2895);
and U3153 (N_3153,N_2868,N_2875);
nor U3154 (N_3154,N_2877,N_2584);
or U3155 (N_3155,N_2705,N_2866);
or U3156 (N_3156,N_2819,N_2973);
and U3157 (N_3157,N_2820,N_2557);
or U3158 (N_3158,N_2809,N_2852);
nor U3159 (N_3159,N_2882,N_2600);
nand U3160 (N_3160,N_2848,N_2581);
and U3161 (N_3161,N_2648,N_2722);
nor U3162 (N_3162,N_2915,N_2601);
nand U3163 (N_3163,N_2726,N_2736);
xor U3164 (N_3164,N_2773,N_2641);
nor U3165 (N_3165,N_2620,N_2935);
or U3166 (N_3166,N_2670,N_2614);
nand U3167 (N_3167,N_2843,N_2592);
and U3168 (N_3168,N_2530,N_2526);
or U3169 (N_3169,N_2881,N_2561);
nor U3170 (N_3170,N_2862,N_2890);
nor U3171 (N_3171,N_2505,N_2649);
nand U3172 (N_3172,N_2509,N_2501);
and U3173 (N_3173,N_2646,N_2805);
and U3174 (N_3174,N_2772,N_2859);
nand U3175 (N_3175,N_2815,N_2831);
and U3176 (N_3176,N_2830,N_2680);
nand U3177 (N_3177,N_2570,N_2650);
xor U3178 (N_3178,N_2661,N_2563);
nor U3179 (N_3179,N_2676,N_2610);
xor U3180 (N_3180,N_2774,N_2995);
xor U3181 (N_3181,N_2571,N_2801);
nor U3182 (N_3182,N_2707,N_2902);
nor U3183 (N_3183,N_2523,N_2790);
xor U3184 (N_3184,N_2765,N_2989);
nand U3185 (N_3185,N_2869,N_2826);
nand U3186 (N_3186,N_2943,N_2998);
nor U3187 (N_3187,N_2802,N_2853);
or U3188 (N_3188,N_2921,N_2845);
nor U3189 (N_3189,N_2690,N_2796);
xnor U3190 (N_3190,N_2559,N_2984);
nand U3191 (N_3191,N_2807,N_2515);
nand U3192 (N_3192,N_2685,N_2524);
xor U3193 (N_3193,N_2970,N_2513);
xor U3194 (N_3194,N_2749,N_2599);
nand U3195 (N_3195,N_2692,N_2824);
nand U3196 (N_3196,N_2536,N_2652);
xnor U3197 (N_3197,N_2728,N_2854);
or U3198 (N_3198,N_2566,N_2779);
and U3199 (N_3199,N_2874,N_2617);
nor U3200 (N_3200,N_2683,N_2543);
nor U3201 (N_3201,N_2746,N_2694);
nand U3202 (N_3202,N_2978,N_2507);
xor U3203 (N_3203,N_2951,N_2954);
and U3204 (N_3204,N_2691,N_2768);
or U3205 (N_3205,N_2541,N_2760);
and U3206 (N_3206,N_2752,N_2911);
nand U3207 (N_3207,N_2828,N_2631);
nand U3208 (N_3208,N_2972,N_2711);
nor U3209 (N_3209,N_2727,N_2547);
nand U3210 (N_3210,N_2696,N_2941);
and U3211 (N_3211,N_2931,N_2721);
nor U3212 (N_3212,N_2688,N_2672);
and U3213 (N_3213,N_2579,N_2775);
or U3214 (N_3214,N_2948,N_2606);
xnor U3215 (N_3215,N_2698,N_2810);
nand U3216 (N_3216,N_2982,N_2798);
xor U3217 (N_3217,N_2743,N_2537);
or U3218 (N_3218,N_2718,N_2629);
nor U3219 (N_3219,N_2663,N_2701);
or U3220 (N_3220,N_2844,N_2734);
nor U3221 (N_3221,N_2598,N_2878);
nand U3222 (N_3222,N_2605,N_2731);
nand U3223 (N_3223,N_2677,N_2643);
or U3224 (N_3224,N_2873,N_2799);
and U3225 (N_3225,N_2979,N_2735);
nor U3226 (N_3226,N_2927,N_2867);
nand U3227 (N_3227,N_2574,N_2947);
and U3228 (N_3228,N_2876,N_2732);
nand U3229 (N_3229,N_2745,N_2575);
or U3230 (N_3230,N_2615,N_2714);
nor U3231 (N_3231,N_2933,N_2788);
or U3232 (N_3232,N_2528,N_2591);
or U3233 (N_3233,N_2626,N_2922);
and U3234 (N_3234,N_2838,N_2658);
and U3235 (N_3235,N_2506,N_2589);
or U3236 (N_3236,N_2720,N_2812);
nor U3237 (N_3237,N_2596,N_2744);
and U3238 (N_3238,N_2708,N_2961);
nor U3239 (N_3239,N_2621,N_2568);
nand U3240 (N_3240,N_2741,N_2738);
nor U3241 (N_3241,N_2719,N_2832);
xnor U3242 (N_3242,N_2551,N_2533);
nor U3243 (N_3243,N_2950,N_2983);
or U3244 (N_3244,N_2733,N_2901);
nor U3245 (N_3245,N_2791,N_2565);
or U3246 (N_3246,N_2730,N_2991);
xnor U3247 (N_3247,N_2823,N_2778);
nand U3248 (N_3248,N_2520,N_2630);
or U3249 (N_3249,N_2518,N_2653);
xnor U3250 (N_3250,N_2583,N_2888);
nor U3251 (N_3251,N_2539,N_2709);
and U3252 (N_3252,N_2988,N_2521);
nor U3253 (N_3253,N_2861,N_2581);
nor U3254 (N_3254,N_2817,N_2944);
xnor U3255 (N_3255,N_2612,N_2512);
nand U3256 (N_3256,N_2725,N_2555);
or U3257 (N_3257,N_2684,N_2703);
or U3258 (N_3258,N_2820,N_2954);
or U3259 (N_3259,N_2999,N_2722);
and U3260 (N_3260,N_2695,N_2841);
nor U3261 (N_3261,N_2508,N_2534);
xor U3262 (N_3262,N_2659,N_2677);
xor U3263 (N_3263,N_2800,N_2631);
and U3264 (N_3264,N_2711,N_2719);
nand U3265 (N_3265,N_2578,N_2620);
nand U3266 (N_3266,N_2978,N_2500);
or U3267 (N_3267,N_2612,N_2949);
nand U3268 (N_3268,N_2720,N_2607);
and U3269 (N_3269,N_2601,N_2949);
xor U3270 (N_3270,N_2821,N_2685);
and U3271 (N_3271,N_2709,N_2871);
nor U3272 (N_3272,N_2693,N_2916);
xnor U3273 (N_3273,N_2787,N_2879);
or U3274 (N_3274,N_2738,N_2586);
or U3275 (N_3275,N_2562,N_2582);
or U3276 (N_3276,N_2755,N_2822);
and U3277 (N_3277,N_2695,N_2976);
and U3278 (N_3278,N_2910,N_2947);
nor U3279 (N_3279,N_2664,N_2570);
nor U3280 (N_3280,N_2713,N_2631);
xor U3281 (N_3281,N_2598,N_2638);
and U3282 (N_3282,N_2816,N_2564);
and U3283 (N_3283,N_2644,N_2749);
nor U3284 (N_3284,N_2932,N_2881);
or U3285 (N_3285,N_2836,N_2637);
nor U3286 (N_3286,N_2770,N_2744);
nand U3287 (N_3287,N_2726,N_2607);
and U3288 (N_3288,N_2918,N_2944);
or U3289 (N_3289,N_2927,N_2676);
xor U3290 (N_3290,N_2819,N_2665);
or U3291 (N_3291,N_2738,N_2756);
and U3292 (N_3292,N_2883,N_2678);
or U3293 (N_3293,N_2865,N_2687);
and U3294 (N_3294,N_2526,N_2747);
and U3295 (N_3295,N_2823,N_2572);
xnor U3296 (N_3296,N_2674,N_2998);
and U3297 (N_3297,N_2821,N_2707);
nand U3298 (N_3298,N_2669,N_2595);
and U3299 (N_3299,N_2879,N_2636);
and U3300 (N_3300,N_2870,N_2850);
nor U3301 (N_3301,N_2951,N_2606);
and U3302 (N_3302,N_2730,N_2728);
xnor U3303 (N_3303,N_2926,N_2774);
nand U3304 (N_3304,N_2514,N_2714);
nor U3305 (N_3305,N_2781,N_2750);
or U3306 (N_3306,N_2871,N_2720);
and U3307 (N_3307,N_2645,N_2551);
and U3308 (N_3308,N_2753,N_2624);
and U3309 (N_3309,N_2535,N_2699);
nor U3310 (N_3310,N_2577,N_2696);
or U3311 (N_3311,N_2757,N_2681);
nand U3312 (N_3312,N_2959,N_2535);
nand U3313 (N_3313,N_2739,N_2954);
nor U3314 (N_3314,N_2868,N_2557);
xor U3315 (N_3315,N_2651,N_2536);
xor U3316 (N_3316,N_2819,N_2810);
and U3317 (N_3317,N_2944,N_2674);
xnor U3318 (N_3318,N_2567,N_2919);
xnor U3319 (N_3319,N_2785,N_2741);
nor U3320 (N_3320,N_2828,N_2809);
xnor U3321 (N_3321,N_2866,N_2535);
xor U3322 (N_3322,N_2634,N_2665);
or U3323 (N_3323,N_2503,N_2887);
and U3324 (N_3324,N_2746,N_2625);
xor U3325 (N_3325,N_2795,N_2651);
nand U3326 (N_3326,N_2514,N_2749);
or U3327 (N_3327,N_2684,N_2687);
nand U3328 (N_3328,N_2557,N_2994);
xnor U3329 (N_3329,N_2770,N_2800);
nor U3330 (N_3330,N_2676,N_2893);
nand U3331 (N_3331,N_2924,N_2861);
or U3332 (N_3332,N_2525,N_2520);
or U3333 (N_3333,N_2961,N_2711);
xor U3334 (N_3334,N_2714,N_2931);
or U3335 (N_3335,N_2585,N_2720);
nand U3336 (N_3336,N_2703,N_2521);
and U3337 (N_3337,N_2662,N_2658);
xnor U3338 (N_3338,N_2937,N_2703);
or U3339 (N_3339,N_2807,N_2604);
nand U3340 (N_3340,N_2761,N_2906);
nand U3341 (N_3341,N_2967,N_2538);
and U3342 (N_3342,N_2673,N_2503);
xor U3343 (N_3343,N_2964,N_2762);
nand U3344 (N_3344,N_2506,N_2937);
or U3345 (N_3345,N_2741,N_2524);
or U3346 (N_3346,N_2534,N_2793);
nand U3347 (N_3347,N_2653,N_2744);
and U3348 (N_3348,N_2500,N_2659);
nor U3349 (N_3349,N_2991,N_2579);
nand U3350 (N_3350,N_2951,N_2699);
or U3351 (N_3351,N_2548,N_2738);
nor U3352 (N_3352,N_2820,N_2950);
nor U3353 (N_3353,N_2797,N_2936);
nor U3354 (N_3354,N_2806,N_2573);
xnor U3355 (N_3355,N_2815,N_2806);
nand U3356 (N_3356,N_2824,N_2503);
nor U3357 (N_3357,N_2831,N_2507);
or U3358 (N_3358,N_2803,N_2962);
nor U3359 (N_3359,N_2561,N_2694);
xnor U3360 (N_3360,N_2621,N_2982);
and U3361 (N_3361,N_2559,N_2796);
xnor U3362 (N_3362,N_2829,N_2930);
nor U3363 (N_3363,N_2691,N_2510);
or U3364 (N_3364,N_2928,N_2826);
nand U3365 (N_3365,N_2877,N_2526);
xnor U3366 (N_3366,N_2979,N_2698);
or U3367 (N_3367,N_2530,N_2561);
xnor U3368 (N_3368,N_2525,N_2504);
xor U3369 (N_3369,N_2838,N_2626);
nor U3370 (N_3370,N_2512,N_2934);
and U3371 (N_3371,N_2821,N_2706);
or U3372 (N_3372,N_2994,N_2955);
and U3373 (N_3373,N_2766,N_2575);
and U3374 (N_3374,N_2501,N_2584);
and U3375 (N_3375,N_2577,N_2558);
nand U3376 (N_3376,N_2515,N_2808);
nand U3377 (N_3377,N_2689,N_2615);
nor U3378 (N_3378,N_2827,N_2713);
or U3379 (N_3379,N_2510,N_2864);
nand U3380 (N_3380,N_2524,N_2816);
nor U3381 (N_3381,N_2562,N_2944);
nor U3382 (N_3382,N_2884,N_2981);
nand U3383 (N_3383,N_2527,N_2904);
nor U3384 (N_3384,N_2633,N_2648);
nand U3385 (N_3385,N_2793,N_2795);
nor U3386 (N_3386,N_2574,N_2835);
xnor U3387 (N_3387,N_2971,N_2601);
or U3388 (N_3388,N_2914,N_2919);
and U3389 (N_3389,N_2579,N_2724);
or U3390 (N_3390,N_2951,N_2547);
or U3391 (N_3391,N_2826,N_2787);
and U3392 (N_3392,N_2548,N_2868);
xnor U3393 (N_3393,N_2525,N_2532);
and U3394 (N_3394,N_2906,N_2733);
nor U3395 (N_3395,N_2892,N_2798);
xor U3396 (N_3396,N_2841,N_2898);
nand U3397 (N_3397,N_2747,N_2724);
nand U3398 (N_3398,N_2870,N_2916);
and U3399 (N_3399,N_2939,N_2545);
and U3400 (N_3400,N_2873,N_2824);
nor U3401 (N_3401,N_2750,N_2572);
nand U3402 (N_3402,N_2565,N_2789);
or U3403 (N_3403,N_2860,N_2625);
xor U3404 (N_3404,N_2815,N_2931);
or U3405 (N_3405,N_2683,N_2610);
nand U3406 (N_3406,N_2595,N_2981);
nor U3407 (N_3407,N_2697,N_2872);
nand U3408 (N_3408,N_2804,N_2549);
and U3409 (N_3409,N_2816,N_2972);
xor U3410 (N_3410,N_2709,N_2695);
and U3411 (N_3411,N_2924,N_2866);
nor U3412 (N_3412,N_2754,N_2948);
nand U3413 (N_3413,N_2990,N_2551);
and U3414 (N_3414,N_2916,N_2738);
or U3415 (N_3415,N_2723,N_2590);
and U3416 (N_3416,N_2898,N_2633);
or U3417 (N_3417,N_2573,N_2722);
nor U3418 (N_3418,N_2790,N_2852);
nor U3419 (N_3419,N_2701,N_2653);
xnor U3420 (N_3420,N_2531,N_2861);
nand U3421 (N_3421,N_2575,N_2836);
nand U3422 (N_3422,N_2902,N_2555);
nand U3423 (N_3423,N_2986,N_2946);
nor U3424 (N_3424,N_2718,N_2860);
nor U3425 (N_3425,N_2925,N_2972);
xor U3426 (N_3426,N_2949,N_2873);
xnor U3427 (N_3427,N_2552,N_2946);
and U3428 (N_3428,N_2832,N_2521);
nor U3429 (N_3429,N_2770,N_2887);
nor U3430 (N_3430,N_2872,N_2986);
and U3431 (N_3431,N_2983,N_2563);
nor U3432 (N_3432,N_2633,N_2767);
nand U3433 (N_3433,N_2931,N_2578);
xnor U3434 (N_3434,N_2523,N_2691);
xor U3435 (N_3435,N_2982,N_2931);
and U3436 (N_3436,N_2956,N_2823);
nor U3437 (N_3437,N_2869,N_2562);
nand U3438 (N_3438,N_2733,N_2623);
nand U3439 (N_3439,N_2944,N_2753);
and U3440 (N_3440,N_2982,N_2624);
xnor U3441 (N_3441,N_2730,N_2664);
or U3442 (N_3442,N_2690,N_2829);
or U3443 (N_3443,N_2693,N_2841);
and U3444 (N_3444,N_2602,N_2751);
nor U3445 (N_3445,N_2742,N_2904);
or U3446 (N_3446,N_2895,N_2653);
and U3447 (N_3447,N_2708,N_2613);
or U3448 (N_3448,N_2935,N_2734);
nand U3449 (N_3449,N_2702,N_2898);
or U3450 (N_3450,N_2660,N_2810);
nand U3451 (N_3451,N_2569,N_2573);
nand U3452 (N_3452,N_2935,N_2618);
and U3453 (N_3453,N_2692,N_2999);
and U3454 (N_3454,N_2977,N_2758);
and U3455 (N_3455,N_2941,N_2911);
nor U3456 (N_3456,N_2586,N_2632);
and U3457 (N_3457,N_2548,N_2817);
nor U3458 (N_3458,N_2860,N_2786);
nand U3459 (N_3459,N_2977,N_2541);
nand U3460 (N_3460,N_2809,N_2925);
or U3461 (N_3461,N_2755,N_2859);
xnor U3462 (N_3462,N_2781,N_2809);
xor U3463 (N_3463,N_2666,N_2671);
nand U3464 (N_3464,N_2852,N_2853);
nor U3465 (N_3465,N_2684,N_2756);
nand U3466 (N_3466,N_2958,N_2665);
and U3467 (N_3467,N_2900,N_2966);
or U3468 (N_3468,N_2554,N_2750);
xor U3469 (N_3469,N_2924,N_2881);
or U3470 (N_3470,N_2778,N_2639);
nor U3471 (N_3471,N_2880,N_2850);
xnor U3472 (N_3472,N_2757,N_2622);
xnor U3473 (N_3473,N_2553,N_2906);
xnor U3474 (N_3474,N_2687,N_2759);
nor U3475 (N_3475,N_2810,N_2602);
nand U3476 (N_3476,N_2653,N_2769);
and U3477 (N_3477,N_2517,N_2600);
xor U3478 (N_3478,N_2731,N_2927);
and U3479 (N_3479,N_2649,N_2624);
nand U3480 (N_3480,N_2952,N_2832);
nor U3481 (N_3481,N_2552,N_2508);
nand U3482 (N_3482,N_2953,N_2769);
nor U3483 (N_3483,N_2656,N_2570);
or U3484 (N_3484,N_2591,N_2618);
nor U3485 (N_3485,N_2608,N_2510);
nor U3486 (N_3486,N_2740,N_2884);
nand U3487 (N_3487,N_2697,N_2658);
and U3488 (N_3488,N_2852,N_2635);
nor U3489 (N_3489,N_2617,N_2928);
or U3490 (N_3490,N_2537,N_2876);
nand U3491 (N_3491,N_2939,N_2522);
or U3492 (N_3492,N_2802,N_2708);
or U3493 (N_3493,N_2655,N_2990);
or U3494 (N_3494,N_2752,N_2904);
or U3495 (N_3495,N_2806,N_2653);
nand U3496 (N_3496,N_2521,N_2894);
and U3497 (N_3497,N_2642,N_2673);
nand U3498 (N_3498,N_2714,N_2564);
nand U3499 (N_3499,N_2637,N_2931);
or U3500 (N_3500,N_3413,N_3316);
and U3501 (N_3501,N_3027,N_3350);
nand U3502 (N_3502,N_3432,N_3305);
and U3503 (N_3503,N_3425,N_3035);
or U3504 (N_3504,N_3000,N_3160);
nor U3505 (N_3505,N_3203,N_3284);
nand U3506 (N_3506,N_3463,N_3459);
xnor U3507 (N_3507,N_3393,N_3013);
nand U3508 (N_3508,N_3171,N_3270);
nor U3509 (N_3509,N_3483,N_3254);
xnor U3510 (N_3510,N_3398,N_3217);
nand U3511 (N_3511,N_3045,N_3351);
nand U3512 (N_3512,N_3208,N_3046);
nand U3513 (N_3513,N_3093,N_3477);
and U3514 (N_3514,N_3016,N_3190);
nor U3515 (N_3515,N_3226,N_3201);
nor U3516 (N_3516,N_3253,N_3052);
nand U3517 (N_3517,N_3380,N_3352);
or U3518 (N_3518,N_3448,N_3139);
and U3519 (N_3519,N_3499,N_3136);
or U3520 (N_3520,N_3358,N_3024);
or U3521 (N_3521,N_3230,N_3296);
nor U3522 (N_3522,N_3435,N_3472);
xnor U3523 (N_3523,N_3144,N_3141);
and U3524 (N_3524,N_3229,N_3241);
nor U3525 (N_3525,N_3222,N_3408);
nor U3526 (N_3526,N_3334,N_3388);
nor U3527 (N_3527,N_3247,N_3063);
xor U3528 (N_3528,N_3064,N_3044);
and U3529 (N_3529,N_3366,N_3414);
or U3530 (N_3530,N_3025,N_3486);
nand U3531 (N_3531,N_3126,N_3062);
xor U3532 (N_3532,N_3231,N_3436);
and U3533 (N_3533,N_3119,N_3251);
nand U3534 (N_3534,N_3315,N_3466);
and U3535 (N_3535,N_3225,N_3422);
or U3536 (N_3536,N_3240,N_3209);
and U3537 (N_3537,N_3485,N_3043);
and U3538 (N_3538,N_3452,N_3238);
nand U3539 (N_3539,N_3451,N_3146);
nor U3540 (N_3540,N_3474,N_3470);
xor U3541 (N_3541,N_3127,N_3212);
nand U3542 (N_3542,N_3234,N_3220);
nand U3543 (N_3543,N_3419,N_3172);
nor U3544 (N_3544,N_3376,N_3018);
xor U3545 (N_3545,N_3424,N_3345);
and U3546 (N_3546,N_3496,N_3204);
xor U3547 (N_3547,N_3105,N_3367);
xnor U3548 (N_3548,N_3069,N_3362);
xnor U3549 (N_3549,N_3030,N_3487);
or U3550 (N_3550,N_3088,N_3070);
and U3551 (N_3551,N_3218,N_3087);
or U3552 (N_3552,N_3465,N_3423);
or U3553 (N_3553,N_3417,N_3154);
xnor U3554 (N_3554,N_3492,N_3498);
nor U3555 (N_3555,N_3009,N_3323);
xor U3556 (N_3556,N_3041,N_3262);
nor U3557 (N_3557,N_3246,N_3040);
and U3558 (N_3558,N_3078,N_3294);
and U3559 (N_3559,N_3329,N_3196);
or U3560 (N_3560,N_3082,N_3180);
or U3561 (N_3561,N_3076,N_3148);
xor U3562 (N_3562,N_3047,N_3245);
nand U3563 (N_3563,N_3428,N_3276);
nand U3564 (N_3564,N_3134,N_3031);
xor U3565 (N_3565,N_3214,N_3322);
and U3566 (N_3566,N_3489,N_3162);
or U3567 (N_3567,N_3060,N_3383);
xor U3568 (N_3568,N_3301,N_3454);
or U3569 (N_3569,N_3447,N_3017);
nand U3570 (N_3570,N_3051,N_3281);
or U3571 (N_3571,N_3143,N_3104);
nand U3572 (N_3572,N_3020,N_3364);
nor U3573 (N_3573,N_3418,N_3372);
and U3574 (N_3574,N_3166,N_3079);
nor U3575 (N_3575,N_3153,N_3444);
and U3576 (N_3576,N_3327,N_3330);
nand U3577 (N_3577,N_3400,N_3083);
nand U3578 (N_3578,N_3033,N_3395);
xor U3579 (N_3579,N_3023,N_3191);
xnor U3580 (N_3580,N_3197,N_3168);
xor U3581 (N_3581,N_3150,N_3390);
or U3582 (N_3582,N_3115,N_3289);
nand U3583 (N_3583,N_3147,N_3198);
and U3584 (N_3584,N_3488,N_3125);
nand U3585 (N_3585,N_3462,N_3122);
xor U3586 (N_3586,N_3346,N_3494);
and U3587 (N_3587,N_3210,N_3271);
or U3588 (N_3588,N_3178,N_3058);
nor U3589 (N_3589,N_3363,N_3103);
and U3590 (N_3590,N_3159,N_3244);
nand U3591 (N_3591,N_3194,N_3003);
and U3592 (N_3592,N_3137,N_3348);
and U3593 (N_3593,N_3286,N_3067);
xnor U3594 (N_3594,N_3096,N_3261);
or U3595 (N_3595,N_3090,N_3443);
nor U3596 (N_3596,N_3193,N_3406);
or U3597 (N_3597,N_3291,N_3184);
nor U3598 (N_3598,N_3108,N_3442);
or U3599 (N_3599,N_3396,N_3453);
and U3600 (N_3600,N_3333,N_3319);
xor U3601 (N_3601,N_3439,N_3002);
nor U3602 (N_3602,N_3310,N_3264);
or U3603 (N_3603,N_3389,N_3258);
nor U3604 (N_3604,N_3365,N_3293);
nand U3605 (N_3605,N_3106,N_3213);
nand U3606 (N_3606,N_3098,N_3384);
nor U3607 (N_3607,N_3121,N_3309);
and U3608 (N_3608,N_3278,N_3192);
and U3609 (N_3609,N_3133,N_3421);
xor U3610 (N_3610,N_3048,N_3361);
or U3611 (N_3611,N_3438,N_3054);
or U3612 (N_3612,N_3131,N_3124);
xor U3613 (N_3613,N_3155,N_3303);
nor U3614 (N_3614,N_3404,N_3337);
and U3615 (N_3615,N_3359,N_3100);
nand U3616 (N_3616,N_3449,N_3074);
xnor U3617 (N_3617,N_3324,N_3109);
nand U3618 (N_3618,N_3138,N_3407);
and U3619 (N_3619,N_3170,N_3469);
xnor U3620 (N_3620,N_3183,N_3297);
or U3621 (N_3621,N_3415,N_3326);
nand U3622 (N_3622,N_3460,N_3292);
and U3623 (N_3623,N_3317,N_3445);
and U3624 (N_3624,N_3274,N_3290);
nand U3625 (N_3625,N_3263,N_3450);
xnor U3626 (N_3626,N_3032,N_3497);
nor U3627 (N_3627,N_3267,N_3354);
and U3628 (N_3628,N_3411,N_3369);
nor U3629 (N_3629,N_3416,N_3308);
nor U3630 (N_3630,N_3275,N_3304);
xor U3631 (N_3631,N_3332,N_3399);
and U3632 (N_3632,N_3368,N_3248);
xor U3633 (N_3633,N_3458,N_3099);
or U3634 (N_3634,N_3216,N_3280);
and U3635 (N_3635,N_3145,N_3176);
xor U3636 (N_3636,N_3233,N_3430);
nand U3637 (N_3637,N_3175,N_3114);
xor U3638 (N_3638,N_3205,N_3412);
nand U3639 (N_3639,N_3356,N_3331);
nor U3640 (N_3640,N_3207,N_3349);
xor U3641 (N_3641,N_3313,N_3397);
or U3642 (N_3642,N_3392,N_3373);
nor U3643 (N_3643,N_3173,N_3116);
nand U3644 (N_3644,N_3199,N_3446);
nand U3645 (N_3645,N_3341,N_3437);
or U3646 (N_3646,N_3336,N_3185);
or U3647 (N_3647,N_3287,N_3039);
xnor U3648 (N_3648,N_3468,N_3312);
or U3649 (N_3649,N_3174,N_3163);
xor U3650 (N_3650,N_3433,N_3236);
and U3651 (N_3651,N_3029,N_3471);
and U3652 (N_3652,N_3042,N_3482);
and U3653 (N_3653,N_3256,N_3490);
or U3654 (N_3654,N_3084,N_3110);
xor U3655 (N_3655,N_3132,N_3420);
or U3656 (N_3656,N_3227,N_3429);
or U3657 (N_3657,N_3091,N_3378);
nor U3658 (N_3658,N_3252,N_3034);
or U3659 (N_3659,N_3038,N_3097);
nor U3660 (N_3660,N_3129,N_3385);
or U3661 (N_3661,N_3357,N_3475);
nand U3662 (N_3662,N_3158,N_3255);
or U3663 (N_3663,N_3243,N_3285);
or U3664 (N_3664,N_3461,N_3375);
nor U3665 (N_3665,N_3335,N_3094);
nand U3666 (N_3666,N_3370,N_3391);
nand U3667 (N_3667,N_3320,N_3057);
nand U3668 (N_3668,N_3182,N_3484);
and U3669 (N_3669,N_3353,N_3379);
xor U3670 (N_3670,N_3250,N_3298);
and U3671 (N_3671,N_3339,N_3161);
nor U3672 (N_3672,N_3149,N_3004);
and U3673 (N_3673,N_3401,N_3065);
and U3674 (N_3674,N_3135,N_3342);
and U3675 (N_3675,N_3072,N_3242);
nand U3676 (N_3676,N_3478,N_3374);
nand U3677 (N_3677,N_3140,N_3405);
or U3678 (N_3678,N_3077,N_3071);
and U3679 (N_3679,N_3221,N_3202);
nor U3680 (N_3680,N_3328,N_3382);
xnor U3681 (N_3681,N_3050,N_3387);
or U3682 (N_3682,N_3228,N_3095);
nor U3683 (N_3683,N_3295,N_3306);
or U3684 (N_3684,N_3343,N_3409);
or U3685 (N_3685,N_3355,N_3179);
and U3686 (N_3686,N_3402,N_3006);
nor U3687 (N_3687,N_3495,N_3061);
or U3688 (N_3688,N_3089,N_3165);
nor U3689 (N_3689,N_3288,N_3169);
nor U3690 (N_3690,N_3427,N_3117);
nor U3691 (N_3691,N_3344,N_3235);
nand U3692 (N_3692,N_3037,N_3012);
xnor U3693 (N_3693,N_3219,N_3457);
nand U3694 (N_3694,N_3200,N_3403);
nor U3695 (N_3695,N_3476,N_3347);
and U3696 (N_3696,N_3410,N_3215);
and U3697 (N_3697,N_3273,N_3307);
and U3698 (N_3698,N_3377,N_3481);
nand U3699 (N_3699,N_3049,N_3426);
or U3700 (N_3700,N_3249,N_3102);
nor U3701 (N_3701,N_3279,N_3187);
nor U3702 (N_3702,N_3318,N_3480);
nand U3703 (N_3703,N_3130,N_3008);
nand U3704 (N_3704,N_3268,N_3272);
nor U3705 (N_3705,N_3101,N_3157);
or U3706 (N_3706,N_3302,N_3223);
xnor U3707 (N_3707,N_3015,N_3237);
and U3708 (N_3708,N_3022,N_3112);
xor U3709 (N_3709,N_3257,N_3282);
xnor U3710 (N_3710,N_3026,N_3239);
and U3711 (N_3711,N_3086,N_3007);
nand U3712 (N_3712,N_3011,N_3118);
nand U3713 (N_3713,N_3338,N_3195);
nand U3714 (N_3714,N_3181,N_3085);
or U3715 (N_3715,N_3265,N_3260);
nand U3716 (N_3716,N_3381,N_3269);
nand U3717 (N_3717,N_3434,N_3081);
nand U3718 (N_3718,N_3340,N_3001);
nand U3719 (N_3719,N_3467,N_3151);
nand U3720 (N_3720,N_3107,N_3299);
nor U3721 (N_3721,N_3113,N_3059);
and U3722 (N_3722,N_3111,N_3142);
or U3723 (N_3723,N_3189,N_3053);
or U3724 (N_3724,N_3073,N_3455);
or U3725 (N_3725,N_3056,N_3167);
or U3726 (N_3726,N_3186,N_3019);
xor U3727 (N_3727,N_3431,N_3479);
xor U3728 (N_3728,N_3164,N_3066);
xnor U3729 (N_3729,N_3055,N_3206);
and U3730 (N_3730,N_3441,N_3394);
or U3731 (N_3731,N_3360,N_3300);
or U3732 (N_3732,N_3120,N_3211);
nand U3733 (N_3733,N_3036,N_3277);
or U3734 (N_3734,N_3325,N_3440);
or U3735 (N_3735,N_3491,N_3232);
or U3736 (N_3736,N_3092,N_3068);
and U3737 (N_3737,N_3177,N_3075);
and U3738 (N_3738,N_3224,N_3128);
and U3739 (N_3739,N_3156,N_3314);
and U3740 (N_3740,N_3311,N_3493);
and U3741 (N_3741,N_3473,N_3283);
nand U3742 (N_3742,N_3005,N_3021);
or U3743 (N_3743,N_3028,N_3080);
nand U3744 (N_3744,N_3266,N_3188);
and U3745 (N_3745,N_3010,N_3464);
nand U3746 (N_3746,N_3456,N_3321);
or U3747 (N_3747,N_3123,N_3371);
and U3748 (N_3748,N_3386,N_3259);
nor U3749 (N_3749,N_3152,N_3014);
and U3750 (N_3750,N_3414,N_3064);
and U3751 (N_3751,N_3013,N_3006);
and U3752 (N_3752,N_3034,N_3156);
nor U3753 (N_3753,N_3407,N_3091);
or U3754 (N_3754,N_3024,N_3125);
or U3755 (N_3755,N_3081,N_3067);
xnor U3756 (N_3756,N_3410,N_3337);
nor U3757 (N_3757,N_3210,N_3316);
nand U3758 (N_3758,N_3420,N_3242);
xor U3759 (N_3759,N_3339,N_3395);
and U3760 (N_3760,N_3329,N_3147);
or U3761 (N_3761,N_3003,N_3303);
nand U3762 (N_3762,N_3093,N_3383);
nor U3763 (N_3763,N_3436,N_3443);
nand U3764 (N_3764,N_3317,N_3454);
nor U3765 (N_3765,N_3114,N_3299);
and U3766 (N_3766,N_3292,N_3305);
or U3767 (N_3767,N_3181,N_3167);
and U3768 (N_3768,N_3449,N_3364);
nand U3769 (N_3769,N_3111,N_3396);
nand U3770 (N_3770,N_3376,N_3213);
xnor U3771 (N_3771,N_3174,N_3146);
nand U3772 (N_3772,N_3078,N_3073);
nand U3773 (N_3773,N_3390,N_3187);
or U3774 (N_3774,N_3168,N_3259);
xor U3775 (N_3775,N_3187,N_3266);
xor U3776 (N_3776,N_3404,N_3306);
and U3777 (N_3777,N_3346,N_3303);
or U3778 (N_3778,N_3071,N_3059);
nand U3779 (N_3779,N_3402,N_3403);
nand U3780 (N_3780,N_3206,N_3016);
and U3781 (N_3781,N_3118,N_3064);
nor U3782 (N_3782,N_3479,N_3354);
xnor U3783 (N_3783,N_3354,N_3058);
nor U3784 (N_3784,N_3113,N_3004);
nor U3785 (N_3785,N_3363,N_3335);
nor U3786 (N_3786,N_3199,N_3376);
and U3787 (N_3787,N_3154,N_3036);
xor U3788 (N_3788,N_3426,N_3231);
and U3789 (N_3789,N_3118,N_3179);
nor U3790 (N_3790,N_3016,N_3247);
xor U3791 (N_3791,N_3450,N_3388);
xor U3792 (N_3792,N_3032,N_3081);
nand U3793 (N_3793,N_3070,N_3447);
and U3794 (N_3794,N_3440,N_3286);
nor U3795 (N_3795,N_3225,N_3099);
nor U3796 (N_3796,N_3437,N_3408);
nor U3797 (N_3797,N_3438,N_3378);
and U3798 (N_3798,N_3221,N_3096);
and U3799 (N_3799,N_3000,N_3478);
nor U3800 (N_3800,N_3288,N_3244);
or U3801 (N_3801,N_3211,N_3404);
nor U3802 (N_3802,N_3165,N_3325);
nand U3803 (N_3803,N_3242,N_3047);
xnor U3804 (N_3804,N_3057,N_3016);
or U3805 (N_3805,N_3274,N_3252);
or U3806 (N_3806,N_3102,N_3490);
xor U3807 (N_3807,N_3251,N_3380);
nand U3808 (N_3808,N_3032,N_3456);
or U3809 (N_3809,N_3154,N_3279);
nand U3810 (N_3810,N_3439,N_3029);
or U3811 (N_3811,N_3476,N_3410);
and U3812 (N_3812,N_3083,N_3015);
or U3813 (N_3813,N_3228,N_3454);
or U3814 (N_3814,N_3019,N_3398);
and U3815 (N_3815,N_3298,N_3166);
xor U3816 (N_3816,N_3009,N_3335);
nand U3817 (N_3817,N_3032,N_3060);
and U3818 (N_3818,N_3393,N_3274);
or U3819 (N_3819,N_3124,N_3098);
and U3820 (N_3820,N_3455,N_3017);
nor U3821 (N_3821,N_3196,N_3343);
xnor U3822 (N_3822,N_3227,N_3286);
or U3823 (N_3823,N_3276,N_3497);
nand U3824 (N_3824,N_3376,N_3217);
nand U3825 (N_3825,N_3355,N_3224);
nand U3826 (N_3826,N_3024,N_3494);
nor U3827 (N_3827,N_3061,N_3276);
and U3828 (N_3828,N_3047,N_3071);
nor U3829 (N_3829,N_3446,N_3088);
nand U3830 (N_3830,N_3473,N_3472);
or U3831 (N_3831,N_3374,N_3168);
nor U3832 (N_3832,N_3371,N_3282);
xor U3833 (N_3833,N_3261,N_3054);
nor U3834 (N_3834,N_3340,N_3072);
or U3835 (N_3835,N_3067,N_3319);
and U3836 (N_3836,N_3464,N_3161);
or U3837 (N_3837,N_3217,N_3105);
nand U3838 (N_3838,N_3102,N_3076);
or U3839 (N_3839,N_3240,N_3024);
nor U3840 (N_3840,N_3191,N_3056);
and U3841 (N_3841,N_3225,N_3285);
or U3842 (N_3842,N_3132,N_3320);
or U3843 (N_3843,N_3228,N_3227);
and U3844 (N_3844,N_3384,N_3133);
and U3845 (N_3845,N_3390,N_3027);
nor U3846 (N_3846,N_3310,N_3205);
or U3847 (N_3847,N_3227,N_3181);
nand U3848 (N_3848,N_3483,N_3226);
and U3849 (N_3849,N_3065,N_3454);
or U3850 (N_3850,N_3323,N_3344);
xor U3851 (N_3851,N_3016,N_3484);
nor U3852 (N_3852,N_3227,N_3230);
nand U3853 (N_3853,N_3188,N_3059);
and U3854 (N_3854,N_3464,N_3234);
and U3855 (N_3855,N_3294,N_3232);
nand U3856 (N_3856,N_3448,N_3033);
nand U3857 (N_3857,N_3241,N_3415);
nor U3858 (N_3858,N_3141,N_3100);
or U3859 (N_3859,N_3254,N_3445);
xnor U3860 (N_3860,N_3296,N_3022);
nor U3861 (N_3861,N_3348,N_3390);
xor U3862 (N_3862,N_3398,N_3372);
or U3863 (N_3863,N_3317,N_3248);
and U3864 (N_3864,N_3234,N_3192);
xnor U3865 (N_3865,N_3027,N_3392);
or U3866 (N_3866,N_3138,N_3041);
nor U3867 (N_3867,N_3011,N_3143);
nand U3868 (N_3868,N_3466,N_3242);
and U3869 (N_3869,N_3081,N_3485);
or U3870 (N_3870,N_3170,N_3259);
xnor U3871 (N_3871,N_3201,N_3446);
and U3872 (N_3872,N_3490,N_3116);
nor U3873 (N_3873,N_3366,N_3457);
nor U3874 (N_3874,N_3030,N_3375);
xnor U3875 (N_3875,N_3177,N_3213);
xnor U3876 (N_3876,N_3221,N_3277);
nand U3877 (N_3877,N_3069,N_3010);
nor U3878 (N_3878,N_3185,N_3172);
or U3879 (N_3879,N_3372,N_3083);
nand U3880 (N_3880,N_3355,N_3406);
nor U3881 (N_3881,N_3362,N_3489);
nand U3882 (N_3882,N_3150,N_3175);
and U3883 (N_3883,N_3134,N_3139);
and U3884 (N_3884,N_3358,N_3255);
nor U3885 (N_3885,N_3124,N_3239);
nand U3886 (N_3886,N_3254,N_3233);
and U3887 (N_3887,N_3469,N_3119);
nor U3888 (N_3888,N_3395,N_3418);
or U3889 (N_3889,N_3183,N_3119);
nor U3890 (N_3890,N_3057,N_3135);
nor U3891 (N_3891,N_3387,N_3409);
nand U3892 (N_3892,N_3102,N_3442);
and U3893 (N_3893,N_3117,N_3035);
nand U3894 (N_3894,N_3406,N_3224);
or U3895 (N_3895,N_3467,N_3195);
xnor U3896 (N_3896,N_3406,N_3240);
nor U3897 (N_3897,N_3162,N_3014);
xor U3898 (N_3898,N_3372,N_3392);
and U3899 (N_3899,N_3248,N_3250);
or U3900 (N_3900,N_3033,N_3009);
and U3901 (N_3901,N_3113,N_3389);
nor U3902 (N_3902,N_3352,N_3336);
and U3903 (N_3903,N_3075,N_3200);
nand U3904 (N_3904,N_3277,N_3332);
or U3905 (N_3905,N_3300,N_3171);
or U3906 (N_3906,N_3385,N_3408);
xor U3907 (N_3907,N_3134,N_3376);
and U3908 (N_3908,N_3354,N_3080);
nand U3909 (N_3909,N_3276,N_3256);
and U3910 (N_3910,N_3461,N_3116);
nor U3911 (N_3911,N_3047,N_3371);
nor U3912 (N_3912,N_3080,N_3339);
or U3913 (N_3913,N_3372,N_3299);
nor U3914 (N_3914,N_3085,N_3390);
nand U3915 (N_3915,N_3073,N_3464);
or U3916 (N_3916,N_3284,N_3457);
or U3917 (N_3917,N_3024,N_3117);
nand U3918 (N_3918,N_3160,N_3117);
nor U3919 (N_3919,N_3039,N_3235);
nor U3920 (N_3920,N_3205,N_3460);
and U3921 (N_3921,N_3068,N_3119);
or U3922 (N_3922,N_3109,N_3112);
xnor U3923 (N_3923,N_3296,N_3352);
and U3924 (N_3924,N_3422,N_3341);
and U3925 (N_3925,N_3123,N_3039);
nand U3926 (N_3926,N_3216,N_3374);
xnor U3927 (N_3927,N_3260,N_3099);
or U3928 (N_3928,N_3219,N_3163);
or U3929 (N_3929,N_3341,N_3210);
or U3930 (N_3930,N_3489,N_3337);
or U3931 (N_3931,N_3303,N_3074);
xor U3932 (N_3932,N_3044,N_3004);
nor U3933 (N_3933,N_3411,N_3431);
xnor U3934 (N_3934,N_3004,N_3350);
xnor U3935 (N_3935,N_3313,N_3074);
nor U3936 (N_3936,N_3406,N_3068);
xor U3937 (N_3937,N_3309,N_3431);
and U3938 (N_3938,N_3091,N_3102);
nor U3939 (N_3939,N_3088,N_3041);
xnor U3940 (N_3940,N_3304,N_3470);
nand U3941 (N_3941,N_3443,N_3054);
xnor U3942 (N_3942,N_3091,N_3075);
nand U3943 (N_3943,N_3316,N_3120);
and U3944 (N_3944,N_3441,N_3014);
nor U3945 (N_3945,N_3309,N_3358);
or U3946 (N_3946,N_3429,N_3461);
nand U3947 (N_3947,N_3354,N_3029);
or U3948 (N_3948,N_3029,N_3452);
nor U3949 (N_3949,N_3475,N_3147);
xnor U3950 (N_3950,N_3491,N_3430);
nor U3951 (N_3951,N_3023,N_3294);
nand U3952 (N_3952,N_3215,N_3402);
nor U3953 (N_3953,N_3169,N_3204);
xor U3954 (N_3954,N_3202,N_3475);
nand U3955 (N_3955,N_3255,N_3437);
nor U3956 (N_3956,N_3028,N_3035);
xor U3957 (N_3957,N_3149,N_3238);
nor U3958 (N_3958,N_3196,N_3471);
or U3959 (N_3959,N_3364,N_3013);
and U3960 (N_3960,N_3372,N_3252);
and U3961 (N_3961,N_3068,N_3172);
xor U3962 (N_3962,N_3478,N_3417);
xor U3963 (N_3963,N_3350,N_3419);
xor U3964 (N_3964,N_3214,N_3231);
or U3965 (N_3965,N_3283,N_3466);
nor U3966 (N_3966,N_3096,N_3165);
and U3967 (N_3967,N_3016,N_3049);
nand U3968 (N_3968,N_3203,N_3352);
xnor U3969 (N_3969,N_3013,N_3445);
xnor U3970 (N_3970,N_3358,N_3091);
or U3971 (N_3971,N_3269,N_3146);
nand U3972 (N_3972,N_3006,N_3127);
or U3973 (N_3973,N_3047,N_3459);
nor U3974 (N_3974,N_3303,N_3326);
xor U3975 (N_3975,N_3043,N_3072);
and U3976 (N_3976,N_3442,N_3192);
nor U3977 (N_3977,N_3237,N_3252);
nand U3978 (N_3978,N_3440,N_3174);
nand U3979 (N_3979,N_3186,N_3369);
and U3980 (N_3980,N_3391,N_3145);
nor U3981 (N_3981,N_3281,N_3452);
or U3982 (N_3982,N_3227,N_3193);
nor U3983 (N_3983,N_3008,N_3210);
nand U3984 (N_3984,N_3424,N_3417);
xnor U3985 (N_3985,N_3165,N_3382);
or U3986 (N_3986,N_3334,N_3464);
nand U3987 (N_3987,N_3219,N_3421);
xnor U3988 (N_3988,N_3422,N_3102);
nor U3989 (N_3989,N_3272,N_3153);
and U3990 (N_3990,N_3106,N_3372);
or U3991 (N_3991,N_3333,N_3099);
nor U3992 (N_3992,N_3388,N_3390);
nand U3993 (N_3993,N_3392,N_3164);
nor U3994 (N_3994,N_3364,N_3004);
nand U3995 (N_3995,N_3056,N_3196);
nand U3996 (N_3996,N_3357,N_3032);
or U3997 (N_3997,N_3481,N_3088);
nor U3998 (N_3998,N_3451,N_3271);
nor U3999 (N_3999,N_3492,N_3183);
nor U4000 (N_4000,N_3551,N_3730);
nor U4001 (N_4001,N_3563,N_3629);
and U4002 (N_4002,N_3699,N_3988);
xnor U4003 (N_4003,N_3689,N_3815);
nand U4004 (N_4004,N_3942,N_3915);
nand U4005 (N_4005,N_3644,N_3521);
or U4006 (N_4006,N_3986,N_3561);
xor U4007 (N_4007,N_3627,N_3976);
nor U4008 (N_4008,N_3820,N_3873);
or U4009 (N_4009,N_3672,N_3927);
or U4010 (N_4010,N_3603,N_3530);
nand U4011 (N_4011,N_3640,N_3651);
nor U4012 (N_4012,N_3859,N_3802);
nor U4013 (N_4013,N_3887,N_3958);
xor U4014 (N_4014,N_3749,N_3877);
and U4015 (N_4015,N_3991,N_3723);
nor U4016 (N_4016,N_3720,N_3557);
nand U4017 (N_4017,N_3940,N_3900);
or U4018 (N_4018,N_3786,N_3658);
nor U4019 (N_4019,N_3593,N_3770);
nand U4020 (N_4020,N_3606,N_3588);
or U4021 (N_4021,N_3715,N_3962);
xor U4022 (N_4022,N_3894,N_3743);
or U4023 (N_4023,N_3590,N_3684);
and U4024 (N_4024,N_3504,N_3577);
nand U4025 (N_4025,N_3949,N_3872);
nor U4026 (N_4026,N_3961,N_3729);
nor U4027 (N_4027,N_3703,N_3951);
or U4028 (N_4028,N_3954,N_3898);
nand U4029 (N_4029,N_3713,N_3569);
xor U4030 (N_4030,N_3666,N_3993);
xnor U4031 (N_4031,N_3550,N_3541);
xor U4032 (N_4032,N_3663,N_3555);
xor U4033 (N_4033,N_3646,N_3519);
or U4034 (N_4034,N_3548,N_3922);
nor U4035 (N_4035,N_3870,N_3762);
xnor U4036 (N_4036,N_3706,N_3570);
nand U4037 (N_4037,N_3682,N_3752);
nand U4038 (N_4038,N_3787,N_3805);
xnor U4039 (N_4039,N_3694,N_3889);
nand U4040 (N_4040,N_3585,N_3661);
or U4041 (N_4041,N_3858,N_3688);
or U4042 (N_4042,N_3533,N_3728);
and U4043 (N_4043,N_3866,N_3635);
or U4044 (N_4044,N_3824,N_3766);
xor U4045 (N_4045,N_3827,N_3578);
xnor U4046 (N_4046,N_3905,N_3617);
and U4047 (N_4047,N_3996,N_3586);
xnor U4048 (N_4048,N_3643,N_3734);
nor U4049 (N_4049,N_3972,N_3732);
and U4050 (N_4050,N_3819,N_3514);
nor U4051 (N_4051,N_3574,N_3837);
and U4052 (N_4052,N_3825,N_3607);
or U4053 (N_4053,N_3618,N_3552);
nor U4054 (N_4054,N_3980,N_3516);
xnor U4055 (N_4055,N_3681,N_3700);
nand U4056 (N_4056,N_3725,N_3526);
or U4057 (N_4057,N_3876,N_3613);
or U4058 (N_4058,N_3901,N_3920);
nand U4059 (N_4059,N_3930,N_3671);
or U4060 (N_4060,N_3724,N_3849);
xor U4061 (N_4061,N_3806,N_3636);
nand U4062 (N_4062,N_3763,N_3871);
xor U4063 (N_4063,N_3801,N_3685);
and U4064 (N_4064,N_3648,N_3829);
nand U4065 (N_4065,N_3518,N_3990);
and U4066 (N_4066,N_3669,N_3977);
xor U4067 (N_4067,N_3884,N_3941);
nand U4068 (N_4068,N_3793,N_3832);
or U4069 (N_4069,N_3931,N_3598);
xor U4070 (N_4070,N_3816,N_3864);
nand U4071 (N_4071,N_3874,N_3739);
or U4072 (N_4072,N_3722,N_3529);
or U4073 (N_4073,N_3934,N_3767);
xor U4074 (N_4074,N_3911,N_3788);
and U4075 (N_4075,N_3619,N_3926);
nand U4076 (N_4076,N_3836,N_3748);
or U4077 (N_4077,N_3830,N_3960);
and U4078 (N_4078,N_3620,N_3566);
nor U4079 (N_4079,N_3535,N_3674);
and U4080 (N_4080,N_3850,N_3537);
xor U4081 (N_4081,N_3584,N_3579);
and U4082 (N_4082,N_3846,N_3544);
xor U4083 (N_4083,N_3831,N_3969);
xor U4084 (N_4084,N_3853,N_3792);
nor U4085 (N_4085,N_3811,N_3841);
nand U4086 (N_4086,N_3891,N_3860);
nor U4087 (N_4087,N_3880,N_3800);
or U4088 (N_4088,N_3592,N_3842);
nand U4089 (N_4089,N_3676,N_3956);
nor U4090 (N_4090,N_3984,N_3594);
nor U4091 (N_4091,N_3978,N_3966);
xnor U4092 (N_4092,N_3721,N_3929);
nand U4093 (N_4093,N_3707,N_3974);
nand U4094 (N_4094,N_3946,N_3711);
or U4095 (N_4095,N_3667,N_3597);
xnor U4096 (N_4096,N_3791,N_3527);
nand U4097 (N_4097,N_3848,N_3686);
nand U4098 (N_4098,N_3695,N_3865);
xnor U4099 (N_4099,N_3675,N_3835);
and U4100 (N_4100,N_3639,N_3718);
xnor U4101 (N_4101,N_3596,N_3771);
nor U4102 (N_4102,N_3948,N_3742);
nand U4103 (N_4103,N_3807,N_3716);
and U4104 (N_4104,N_3632,N_3655);
xor U4105 (N_4105,N_3882,N_3572);
xor U4106 (N_4106,N_3808,N_3952);
xnor U4107 (N_4107,N_3895,N_3710);
or U4108 (N_4108,N_3520,N_3580);
nand U4109 (N_4109,N_3785,N_3509);
and U4110 (N_4110,N_3997,N_3945);
nand U4111 (N_4111,N_3925,N_3823);
xor U4112 (N_4112,N_3878,N_3531);
or U4113 (N_4113,N_3968,N_3928);
nor U4114 (N_4114,N_3589,N_3532);
nor U4115 (N_4115,N_3540,N_3575);
nor U4116 (N_4116,N_3818,N_3654);
nor U4117 (N_4117,N_3653,N_3546);
and U4118 (N_4118,N_3628,N_3776);
and U4119 (N_4119,N_3691,N_3868);
nand U4120 (N_4120,N_3558,N_3567);
xnor U4121 (N_4121,N_3896,N_3517);
and U4122 (N_4122,N_3804,N_3936);
nor U4123 (N_4123,N_3600,N_3565);
nor U4124 (N_4124,N_3981,N_3845);
xor U4125 (N_4125,N_3660,N_3549);
and U4126 (N_4126,N_3759,N_3528);
and U4127 (N_4127,N_3964,N_3697);
and U4128 (N_4128,N_3611,N_3963);
nand U4129 (N_4129,N_3781,N_3862);
and U4130 (N_4130,N_3615,N_3994);
and U4131 (N_4131,N_3547,N_3708);
or U4132 (N_4132,N_3851,N_3733);
or U4133 (N_4133,N_3799,N_3602);
xor U4134 (N_4134,N_3524,N_3614);
and U4135 (N_4135,N_3735,N_3794);
or U4136 (N_4136,N_3916,N_3812);
or U4137 (N_4137,N_3919,N_3538);
xnor U4138 (N_4138,N_3869,N_3634);
nor U4139 (N_4139,N_3624,N_3888);
nand U4140 (N_4140,N_3758,N_3918);
nor U4141 (N_4141,N_3505,N_3534);
xor U4142 (N_4142,N_3693,N_3638);
nor U4143 (N_4143,N_3965,N_3652);
xnor U4144 (N_4144,N_3731,N_3630);
nor U4145 (N_4145,N_3784,N_3844);
xor U4146 (N_4146,N_3959,N_3647);
and U4147 (N_4147,N_3992,N_3756);
and U4148 (N_4148,N_3626,N_3826);
and U4149 (N_4149,N_3625,N_3522);
xnor U4150 (N_4150,N_3863,N_3883);
and U4151 (N_4151,N_3668,N_3828);
xnor U4152 (N_4152,N_3503,N_3795);
and U4153 (N_4153,N_3744,N_3560);
or U4154 (N_4154,N_3501,N_3539);
xor U4155 (N_4155,N_3641,N_3857);
nor U4156 (N_4156,N_3803,N_3657);
nor U4157 (N_4157,N_3840,N_3559);
xnor U4158 (N_4158,N_3821,N_3678);
and U4159 (N_4159,N_3886,N_3995);
xor U4160 (N_4160,N_3543,N_3814);
xor U4161 (N_4161,N_3746,N_3692);
or U4162 (N_4162,N_3677,N_3750);
nand U4163 (N_4163,N_3698,N_3670);
xnor U4164 (N_4164,N_3616,N_3985);
and U4165 (N_4165,N_3664,N_3753);
or U4166 (N_4166,N_3642,N_3937);
nand U4167 (N_4167,N_3932,N_3604);
and U4168 (N_4168,N_3576,N_3975);
xnor U4169 (N_4169,N_3885,N_3912);
or U4170 (N_4170,N_3536,N_3847);
and U4171 (N_4171,N_3727,N_3983);
and U4172 (N_4172,N_3623,N_3854);
or U4173 (N_4173,N_3761,N_3513);
xnor U4174 (N_4174,N_3839,N_3704);
and U4175 (N_4175,N_3754,N_3921);
nor U4176 (N_4176,N_3745,N_3747);
or U4177 (N_4177,N_3998,N_3510);
xor U4178 (N_4178,N_3944,N_3525);
nand U4179 (N_4179,N_3571,N_3553);
xor U4180 (N_4180,N_3507,N_3789);
or U4181 (N_4181,N_3867,N_3659);
and U4182 (N_4182,N_3774,N_3765);
and U4183 (N_4183,N_3892,N_3971);
and U4184 (N_4184,N_3714,N_3938);
and U4185 (N_4185,N_3687,N_3612);
or U4186 (N_4186,N_3631,N_3610);
and U4187 (N_4187,N_3979,N_3738);
nor U4188 (N_4188,N_3508,N_3755);
and U4189 (N_4189,N_3554,N_3907);
and U4190 (N_4190,N_3798,N_3856);
and U4191 (N_4191,N_3621,N_3879);
or U4192 (N_4192,N_3982,N_3810);
and U4193 (N_4193,N_3909,N_3947);
nand U4194 (N_4194,N_3817,N_3701);
xor U4195 (N_4195,N_3855,N_3957);
or U4196 (N_4196,N_3768,N_3709);
and U4197 (N_4197,N_3897,N_3924);
and U4198 (N_4198,N_3568,N_3608);
nand U4199 (N_4199,N_3902,N_3783);
nand U4200 (N_4200,N_3906,N_3939);
and U4201 (N_4201,N_3782,N_3899);
and U4202 (N_4202,N_3757,N_3587);
xor U4203 (N_4203,N_3705,N_3773);
and U4204 (N_4204,N_3777,N_3970);
nor U4205 (N_4205,N_3601,N_3989);
nor U4206 (N_4206,N_3760,N_3893);
nand U4207 (N_4207,N_3999,N_3933);
and U4208 (N_4208,N_3573,N_3903);
nand U4209 (N_4209,N_3890,N_3910);
or U4210 (N_4210,N_3599,N_3583);
and U4211 (N_4211,N_3665,N_3737);
and U4212 (N_4212,N_3650,N_3605);
nor U4213 (N_4213,N_3502,N_3622);
nand U4214 (N_4214,N_3790,N_3736);
xor U4215 (N_4215,N_3778,N_3861);
nor U4216 (N_4216,N_3591,N_3796);
and U4217 (N_4217,N_3904,N_3769);
and U4218 (N_4218,N_3633,N_3834);
xnor U4219 (N_4219,N_3673,N_3581);
nor U4220 (N_4220,N_3843,N_3967);
or U4221 (N_4221,N_3953,N_3582);
nand U4222 (N_4222,N_3690,N_3719);
nor U4223 (N_4223,N_3833,N_3680);
or U4224 (N_4224,N_3511,N_3935);
or U4225 (N_4225,N_3809,N_3500);
nor U4226 (N_4226,N_3913,N_3515);
or U4227 (N_4227,N_3908,N_3564);
or U4228 (N_4228,N_3764,N_3813);
xor U4229 (N_4229,N_3943,N_3649);
or U4230 (N_4230,N_3726,N_3775);
and U4231 (N_4231,N_3545,N_3797);
xor U4232 (N_4232,N_3779,N_3751);
xnor U4233 (N_4233,N_3645,N_3955);
or U4234 (N_4234,N_3740,N_3875);
or U4235 (N_4235,N_3656,N_3512);
nand U4236 (N_4236,N_3881,N_3662);
xor U4237 (N_4237,N_3712,N_3987);
or U4238 (N_4238,N_3683,N_3923);
and U4239 (N_4239,N_3822,N_3702);
xor U4240 (N_4240,N_3852,N_3523);
xor U4241 (N_4241,N_3917,N_3562);
nand U4242 (N_4242,N_3609,N_3717);
xnor U4243 (N_4243,N_3696,N_3838);
xnor U4244 (N_4244,N_3973,N_3679);
nand U4245 (N_4245,N_3780,N_3506);
or U4246 (N_4246,N_3595,N_3950);
xnor U4247 (N_4247,N_3542,N_3772);
or U4248 (N_4248,N_3741,N_3637);
xor U4249 (N_4249,N_3914,N_3556);
nor U4250 (N_4250,N_3767,N_3971);
xnor U4251 (N_4251,N_3534,N_3779);
xnor U4252 (N_4252,N_3516,N_3773);
nor U4253 (N_4253,N_3866,N_3782);
nand U4254 (N_4254,N_3672,N_3554);
xor U4255 (N_4255,N_3979,N_3631);
nor U4256 (N_4256,N_3853,N_3689);
nor U4257 (N_4257,N_3721,N_3531);
nor U4258 (N_4258,N_3957,N_3963);
nor U4259 (N_4259,N_3621,N_3583);
and U4260 (N_4260,N_3506,N_3770);
and U4261 (N_4261,N_3726,N_3637);
nand U4262 (N_4262,N_3643,N_3776);
or U4263 (N_4263,N_3813,N_3561);
and U4264 (N_4264,N_3565,N_3860);
nand U4265 (N_4265,N_3982,N_3653);
nor U4266 (N_4266,N_3982,N_3710);
or U4267 (N_4267,N_3940,N_3590);
nor U4268 (N_4268,N_3951,N_3911);
nand U4269 (N_4269,N_3932,N_3721);
nand U4270 (N_4270,N_3599,N_3727);
nor U4271 (N_4271,N_3544,N_3751);
xor U4272 (N_4272,N_3899,N_3773);
nor U4273 (N_4273,N_3726,N_3977);
and U4274 (N_4274,N_3885,N_3593);
nor U4275 (N_4275,N_3968,N_3809);
nand U4276 (N_4276,N_3779,N_3604);
xor U4277 (N_4277,N_3613,N_3846);
or U4278 (N_4278,N_3975,N_3970);
nand U4279 (N_4279,N_3917,N_3753);
nand U4280 (N_4280,N_3867,N_3587);
or U4281 (N_4281,N_3883,N_3580);
nand U4282 (N_4282,N_3505,N_3922);
nor U4283 (N_4283,N_3865,N_3668);
and U4284 (N_4284,N_3507,N_3536);
xnor U4285 (N_4285,N_3795,N_3918);
and U4286 (N_4286,N_3640,N_3719);
nand U4287 (N_4287,N_3537,N_3945);
nand U4288 (N_4288,N_3678,N_3568);
nand U4289 (N_4289,N_3801,N_3548);
or U4290 (N_4290,N_3773,N_3790);
or U4291 (N_4291,N_3587,N_3803);
nor U4292 (N_4292,N_3683,N_3900);
nand U4293 (N_4293,N_3739,N_3695);
nor U4294 (N_4294,N_3645,N_3515);
nand U4295 (N_4295,N_3628,N_3644);
and U4296 (N_4296,N_3650,N_3510);
xor U4297 (N_4297,N_3987,N_3748);
and U4298 (N_4298,N_3820,N_3516);
xnor U4299 (N_4299,N_3897,N_3798);
nor U4300 (N_4300,N_3544,N_3584);
and U4301 (N_4301,N_3507,N_3538);
nor U4302 (N_4302,N_3530,N_3802);
and U4303 (N_4303,N_3545,N_3842);
or U4304 (N_4304,N_3945,N_3588);
or U4305 (N_4305,N_3770,N_3777);
nand U4306 (N_4306,N_3959,N_3825);
and U4307 (N_4307,N_3687,N_3645);
nor U4308 (N_4308,N_3625,N_3996);
xnor U4309 (N_4309,N_3754,N_3722);
or U4310 (N_4310,N_3836,N_3679);
or U4311 (N_4311,N_3598,N_3551);
or U4312 (N_4312,N_3759,N_3757);
nor U4313 (N_4313,N_3943,N_3645);
and U4314 (N_4314,N_3693,N_3554);
or U4315 (N_4315,N_3596,N_3697);
or U4316 (N_4316,N_3770,N_3756);
nor U4317 (N_4317,N_3994,N_3608);
and U4318 (N_4318,N_3532,N_3712);
and U4319 (N_4319,N_3788,N_3698);
or U4320 (N_4320,N_3628,N_3641);
and U4321 (N_4321,N_3666,N_3956);
and U4322 (N_4322,N_3576,N_3655);
nor U4323 (N_4323,N_3701,N_3769);
nand U4324 (N_4324,N_3585,N_3591);
nor U4325 (N_4325,N_3945,N_3969);
or U4326 (N_4326,N_3986,N_3506);
nand U4327 (N_4327,N_3818,N_3669);
and U4328 (N_4328,N_3982,N_3923);
nor U4329 (N_4329,N_3719,N_3621);
xor U4330 (N_4330,N_3954,N_3705);
xor U4331 (N_4331,N_3628,N_3651);
nor U4332 (N_4332,N_3816,N_3893);
and U4333 (N_4333,N_3803,N_3736);
nand U4334 (N_4334,N_3526,N_3875);
xnor U4335 (N_4335,N_3578,N_3834);
xnor U4336 (N_4336,N_3846,N_3695);
xnor U4337 (N_4337,N_3703,N_3590);
nor U4338 (N_4338,N_3796,N_3540);
or U4339 (N_4339,N_3977,N_3543);
or U4340 (N_4340,N_3598,N_3796);
xnor U4341 (N_4341,N_3555,N_3612);
nor U4342 (N_4342,N_3826,N_3846);
nor U4343 (N_4343,N_3971,N_3560);
nand U4344 (N_4344,N_3886,N_3854);
xor U4345 (N_4345,N_3598,N_3722);
or U4346 (N_4346,N_3778,N_3831);
or U4347 (N_4347,N_3735,N_3503);
or U4348 (N_4348,N_3857,N_3811);
and U4349 (N_4349,N_3772,N_3506);
nand U4350 (N_4350,N_3524,N_3694);
or U4351 (N_4351,N_3684,N_3501);
xor U4352 (N_4352,N_3827,N_3940);
xnor U4353 (N_4353,N_3843,N_3625);
nand U4354 (N_4354,N_3585,N_3682);
or U4355 (N_4355,N_3715,N_3932);
xor U4356 (N_4356,N_3992,N_3660);
xor U4357 (N_4357,N_3925,N_3768);
xnor U4358 (N_4358,N_3549,N_3902);
and U4359 (N_4359,N_3666,N_3892);
nand U4360 (N_4360,N_3541,N_3896);
and U4361 (N_4361,N_3653,N_3551);
or U4362 (N_4362,N_3884,N_3609);
xnor U4363 (N_4363,N_3519,N_3883);
nor U4364 (N_4364,N_3591,N_3761);
nor U4365 (N_4365,N_3881,N_3945);
or U4366 (N_4366,N_3747,N_3573);
and U4367 (N_4367,N_3622,N_3939);
or U4368 (N_4368,N_3659,N_3922);
or U4369 (N_4369,N_3714,N_3633);
nand U4370 (N_4370,N_3854,N_3602);
and U4371 (N_4371,N_3764,N_3529);
xnor U4372 (N_4372,N_3725,N_3860);
or U4373 (N_4373,N_3968,N_3953);
nand U4374 (N_4374,N_3913,N_3823);
and U4375 (N_4375,N_3682,N_3612);
nand U4376 (N_4376,N_3598,N_3750);
xor U4377 (N_4377,N_3867,N_3850);
and U4378 (N_4378,N_3636,N_3988);
xnor U4379 (N_4379,N_3923,N_3740);
or U4380 (N_4380,N_3959,N_3727);
and U4381 (N_4381,N_3904,N_3739);
nor U4382 (N_4382,N_3612,N_3702);
and U4383 (N_4383,N_3772,N_3794);
and U4384 (N_4384,N_3564,N_3806);
nand U4385 (N_4385,N_3688,N_3614);
nand U4386 (N_4386,N_3818,N_3620);
and U4387 (N_4387,N_3956,N_3565);
xor U4388 (N_4388,N_3912,N_3750);
xor U4389 (N_4389,N_3988,N_3808);
nand U4390 (N_4390,N_3941,N_3977);
and U4391 (N_4391,N_3904,N_3704);
and U4392 (N_4392,N_3692,N_3567);
nor U4393 (N_4393,N_3693,N_3883);
and U4394 (N_4394,N_3860,N_3747);
xor U4395 (N_4395,N_3829,N_3927);
nor U4396 (N_4396,N_3776,N_3957);
xnor U4397 (N_4397,N_3715,N_3845);
nor U4398 (N_4398,N_3610,N_3689);
and U4399 (N_4399,N_3581,N_3812);
nand U4400 (N_4400,N_3526,N_3661);
or U4401 (N_4401,N_3862,N_3597);
nand U4402 (N_4402,N_3968,N_3723);
nand U4403 (N_4403,N_3847,N_3540);
nor U4404 (N_4404,N_3622,N_3860);
and U4405 (N_4405,N_3688,N_3570);
xnor U4406 (N_4406,N_3682,N_3846);
nor U4407 (N_4407,N_3665,N_3514);
and U4408 (N_4408,N_3896,N_3727);
xor U4409 (N_4409,N_3903,N_3513);
and U4410 (N_4410,N_3599,N_3948);
nor U4411 (N_4411,N_3659,N_3765);
nor U4412 (N_4412,N_3556,N_3814);
nor U4413 (N_4413,N_3729,N_3978);
and U4414 (N_4414,N_3547,N_3629);
or U4415 (N_4415,N_3564,N_3655);
nor U4416 (N_4416,N_3735,N_3851);
xnor U4417 (N_4417,N_3854,N_3595);
or U4418 (N_4418,N_3853,N_3745);
nand U4419 (N_4419,N_3836,N_3742);
xor U4420 (N_4420,N_3752,N_3881);
xnor U4421 (N_4421,N_3952,N_3527);
nand U4422 (N_4422,N_3783,N_3991);
or U4423 (N_4423,N_3660,N_3633);
nor U4424 (N_4424,N_3656,N_3573);
or U4425 (N_4425,N_3972,N_3595);
or U4426 (N_4426,N_3937,N_3675);
xor U4427 (N_4427,N_3600,N_3914);
nand U4428 (N_4428,N_3905,N_3740);
or U4429 (N_4429,N_3512,N_3513);
nor U4430 (N_4430,N_3710,N_3868);
and U4431 (N_4431,N_3536,N_3758);
xor U4432 (N_4432,N_3686,N_3737);
xor U4433 (N_4433,N_3527,N_3899);
nor U4434 (N_4434,N_3540,N_3709);
or U4435 (N_4435,N_3816,N_3587);
and U4436 (N_4436,N_3583,N_3728);
or U4437 (N_4437,N_3505,N_3509);
or U4438 (N_4438,N_3518,N_3914);
nor U4439 (N_4439,N_3679,N_3943);
or U4440 (N_4440,N_3506,N_3511);
nand U4441 (N_4441,N_3705,N_3562);
nand U4442 (N_4442,N_3655,N_3850);
and U4443 (N_4443,N_3526,N_3701);
or U4444 (N_4444,N_3710,N_3906);
nor U4445 (N_4445,N_3952,N_3942);
nor U4446 (N_4446,N_3763,N_3906);
or U4447 (N_4447,N_3679,N_3739);
xnor U4448 (N_4448,N_3763,N_3829);
nor U4449 (N_4449,N_3925,N_3744);
and U4450 (N_4450,N_3905,N_3717);
nor U4451 (N_4451,N_3708,N_3926);
xnor U4452 (N_4452,N_3822,N_3806);
xnor U4453 (N_4453,N_3769,N_3922);
and U4454 (N_4454,N_3695,N_3572);
and U4455 (N_4455,N_3592,N_3838);
xnor U4456 (N_4456,N_3605,N_3804);
nand U4457 (N_4457,N_3528,N_3516);
xor U4458 (N_4458,N_3756,N_3928);
xnor U4459 (N_4459,N_3809,N_3789);
xor U4460 (N_4460,N_3869,N_3543);
nor U4461 (N_4461,N_3615,N_3875);
xor U4462 (N_4462,N_3979,N_3691);
or U4463 (N_4463,N_3652,N_3991);
nand U4464 (N_4464,N_3949,N_3871);
and U4465 (N_4465,N_3731,N_3513);
and U4466 (N_4466,N_3857,N_3822);
and U4467 (N_4467,N_3958,N_3729);
nor U4468 (N_4468,N_3813,N_3817);
xor U4469 (N_4469,N_3575,N_3970);
or U4470 (N_4470,N_3789,N_3934);
nor U4471 (N_4471,N_3862,N_3826);
and U4472 (N_4472,N_3698,N_3651);
or U4473 (N_4473,N_3974,N_3717);
nand U4474 (N_4474,N_3995,N_3850);
and U4475 (N_4475,N_3575,N_3974);
xor U4476 (N_4476,N_3992,N_3953);
and U4477 (N_4477,N_3880,N_3504);
and U4478 (N_4478,N_3865,N_3686);
nor U4479 (N_4479,N_3843,N_3591);
and U4480 (N_4480,N_3924,N_3832);
nor U4481 (N_4481,N_3659,N_3822);
or U4482 (N_4482,N_3750,N_3699);
or U4483 (N_4483,N_3744,N_3511);
or U4484 (N_4484,N_3819,N_3779);
nor U4485 (N_4485,N_3666,N_3577);
or U4486 (N_4486,N_3637,N_3820);
nand U4487 (N_4487,N_3605,N_3521);
or U4488 (N_4488,N_3724,N_3865);
nand U4489 (N_4489,N_3614,N_3800);
xor U4490 (N_4490,N_3536,N_3949);
and U4491 (N_4491,N_3629,N_3999);
or U4492 (N_4492,N_3922,N_3501);
or U4493 (N_4493,N_3786,N_3991);
nand U4494 (N_4494,N_3780,N_3532);
and U4495 (N_4495,N_3837,N_3950);
or U4496 (N_4496,N_3878,N_3615);
or U4497 (N_4497,N_3774,N_3932);
nand U4498 (N_4498,N_3561,N_3882);
nor U4499 (N_4499,N_3948,N_3882);
xor U4500 (N_4500,N_4204,N_4272);
nand U4501 (N_4501,N_4211,N_4045);
nor U4502 (N_4502,N_4406,N_4118);
nand U4503 (N_4503,N_4248,N_4217);
and U4504 (N_4504,N_4087,N_4444);
nand U4505 (N_4505,N_4119,N_4451);
nor U4506 (N_4506,N_4104,N_4323);
nor U4507 (N_4507,N_4455,N_4254);
or U4508 (N_4508,N_4458,N_4282);
nand U4509 (N_4509,N_4111,N_4441);
nand U4510 (N_4510,N_4416,N_4076);
and U4511 (N_4511,N_4348,N_4328);
nor U4512 (N_4512,N_4342,N_4338);
nand U4513 (N_4513,N_4401,N_4274);
nand U4514 (N_4514,N_4301,N_4378);
xnor U4515 (N_4515,N_4088,N_4051);
or U4516 (N_4516,N_4055,N_4412);
nor U4517 (N_4517,N_4271,N_4198);
nor U4518 (N_4518,N_4464,N_4242);
xor U4519 (N_4519,N_4083,N_4016);
nor U4520 (N_4520,N_4139,N_4168);
and U4521 (N_4521,N_4273,N_4465);
xor U4522 (N_4522,N_4292,N_4394);
nor U4523 (N_4523,N_4000,N_4108);
nand U4524 (N_4524,N_4288,N_4307);
xor U4525 (N_4525,N_4266,N_4240);
and U4526 (N_4526,N_4384,N_4259);
or U4527 (N_4527,N_4123,N_4079);
and U4528 (N_4528,N_4377,N_4106);
and U4529 (N_4529,N_4418,N_4120);
and U4530 (N_4530,N_4233,N_4194);
nor U4531 (N_4531,N_4166,N_4319);
xnor U4532 (N_4532,N_4435,N_4132);
and U4533 (N_4533,N_4480,N_4427);
or U4534 (N_4534,N_4226,N_4404);
and U4535 (N_4535,N_4115,N_4026);
xor U4536 (N_4536,N_4186,N_4320);
and U4537 (N_4537,N_4167,N_4158);
or U4538 (N_4538,N_4053,N_4413);
nand U4539 (N_4539,N_4131,N_4022);
nor U4540 (N_4540,N_4110,N_4380);
and U4541 (N_4541,N_4400,N_4381);
nand U4542 (N_4542,N_4239,N_4260);
nand U4543 (N_4543,N_4363,N_4298);
and U4544 (N_4544,N_4192,N_4302);
nand U4545 (N_4545,N_4483,N_4352);
or U4546 (N_4546,N_4177,N_4486);
xor U4547 (N_4547,N_4407,N_4372);
nand U4548 (N_4548,N_4414,N_4297);
or U4549 (N_4549,N_4442,N_4287);
or U4550 (N_4550,N_4366,N_4084);
nand U4551 (N_4551,N_4475,N_4382);
nand U4552 (N_4552,N_4452,N_4431);
nor U4553 (N_4553,N_4389,N_4246);
and U4554 (N_4554,N_4429,N_4430);
or U4555 (N_4555,N_4202,N_4457);
xnor U4556 (N_4556,N_4270,N_4150);
or U4557 (N_4557,N_4327,N_4059);
xnor U4558 (N_4558,N_4264,N_4344);
xor U4559 (N_4559,N_4080,N_4122);
xor U4560 (N_4560,N_4263,N_4471);
nor U4561 (N_4561,N_4296,N_4293);
or U4562 (N_4562,N_4175,N_4154);
nand U4563 (N_4563,N_4073,N_4280);
xnor U4564 (N_4564,N_4262,N_4481);
xor U4565 (N_4565,N_4215,N_4354);
nand U4566 (N_4566,N_4062,N_4017);
or U4567 (N_4567,N_4112,N_4438);
or U4568 (N_4568,N_4443,N_4456);
or U4569 (N_4569,N_4252,N_4420);
and U4570 (N_4570,N_4020,N_4070);
or U4571 (N_4571,N_4278,N_4487);
or U4572 (N_4572,N_4340,N_4074);
and U4573 (N_4573,N_4057,N_4317);
nand U4574 (N_4574,N_4245,N_4434);
or U4575 (N_4575,N_4379,N_4037);
and U4576 (N_4576,N_4305,N_4250);
nor U4577 (N_4577,N_4002,N_4089);
and U4578 (N_4578,N_4061,N_4490);
nor U4579 (N_4579,N_4228,N_4497);
nor U4580 (N_4580,N_4005,N_4311);
and U4581 (N_4581,N_4304,N_4161);
and U4582 (N_4582,N_4109,N_4035);
nand U4583 (N_4583,N_4256,N_4044);
xnor U4584 (N_4584,N_4001,N_4025);
nor U4585 (N_4585,N_4156,N_4056);
xor U4586 (N_4586,N_4386,N_4375);
xnor U4587 (N_4587,N_4063,N_4437);
or U4588 (N_4588,N_4399,N_4221);
xnor U4589 (N_4589,N_4135,N_4387);
or U4590 (N_4590,N_4402,N_4019);
or U4591 (N_4591,N_4180,N_4043);
nand U4592 (N_4592,N_4213,N_4459);
nand U4593 (N_4593,N_4197,N_4008);
or U4594 (N_4594,N_4157,N_4066);
and U4595 (N_4595,N_4355,N_4172);
nand U4596 (N_4596,N_4113,N_4183);
and U4597 (N_4597,N_4238,N_4454);
and U4598 (N_4598,N_4164,N_4388);
xor U4599 (N_4599,N_4127,N_4229);
and U4600 (N_4600,N_4102,N_4251);
nor U4601 (N_4601,N_4309,N_4212);
nor U4602 (N_4602,N_4145,N_4453);
nor U4603 (N_4603,N_4210,N_4257);
nor U4604 (N_4604,N_4163,N_4100);
or U4605 (N_4605,N_4470,N_4206);
and U4606 (N_4606,N_4247,N_4313);
and U4607 (N_4607,N_4173,N_4463);
nor U4608 (N_4608,N_4314,N_4281);
xor U4609 (N_4609,N_4195,N_4428);
or U4610 (N_4610,N_4013,N_4071);
nor U4611 (N_4611,N_4493,N_4138);
and U4612 (N_4612,N_4050,N_4149);
nor U4613 (N_4613,N_4306,N_4374);
or U4614 (N_4614,N_4201,N_4426);
nor U4615 (N_4615,N_4356,N_4114);
nand U4616 (N_4616,N_4393,N_4294);
and U4617 (N_4617,N_4343,N_4105);
or U4618 (N_4618,N_4143,N_4284);
and U4619 (N_4619,N_4027,N_4461);
and U4620 (N_4620,N_4411,N_4036);
xor U4621 (N_4621,N_4249,N_4015);
and U4622 (N_4622,N_4085,N_4449);
or U4623 (N_4623,N_4324,N_4003);
and U4624 (N_4624,N_4472,N_4170);
or U4625 (N_4625,N_4347,N_4205);
xor U4626 (N_4626,N_4290,N_4337);
or U4627 (N_4627,N_4326,N_4300);
and U4628 (N_4628,N_4383,N_4469);
nand U4629 (N_4629,N_4279,N_4286);
nor U4630 (N_4630,N_4422,N_4203);
or U4631 (N_4631,N_4092,N_4179);
nand U4632 (N_4632,N_4225,N_4448);
and U4633 (N_4633,N_4474,N_4390);
xor U4634 (N_4634,N_4339,N_4227);
and U4635 (N_4635,N_4049,N_4446);
xor U4636 (N_4636,N_4494,N_4146);
or U4637 (N_4637,N_4086,N_4152);
nand U4638 (N_4638,N_4098,N_4403);
or U4639 (N_4639,N_4128,N_4153);
and U4640 (N_4640,N_4365,N_4047);
nand U4641 (N_4641,N_4367,N_4243);
or U4642 (N_4642,N_4155,N_4346);
xor U4643 (N_4643,N_4216,N_4391);
and U4644 (N_4644,N_4207,N_4395);
and U4645 (N_4645,N_4144,N_4498);
nor U4646 (N_4646,N_4358,N_4174);
nand U4647 (N_4647,N_4253,N_4169);
nor U4648 (N_4648,N_4370,N_4136);
and U4649 (N_4649,N_4350,N_4090);
nand U4650 (N_4650,N_4335,N_4151);
nor U4651 (N_4651,N_4268,N_4265);
xor U4652 (N_4652,N_4477,N_4318);
nand U4653 (N_4653,N_4466,N_4409);
xor U4654 (N_4654,N_4368,N_4269);
and U4655 (N_4655,N_4478,N_4064);
nor U4656 (N_4656,N_4042,N_4489);
nor U4657 (N_4657,N_4039,N_4353);
xor U4658 (N_4658,N_4011,N_4329);
and U4659 (N_4659,N_4052,N_4078);
nor U4660 (N_4660,N_4436,N_4095);
xor U4661 (N_4661,N_4376,N_4024);
xor U4662 (N_4662,N_4236,N_4093);
xor U4663 (N_4663,N_4099,N_4275);
xnor U4664 (N_4664,N_4415,N_4065);
xnor U4665 (N_4665,N_4445,N_4142);
and U4666 (N_4666,N_4336,N_4012);
nor U4667 (N_4667,N_4291,N_4182);
xnor U4668 (N_4668,N_4495,N_4094);
nor U4669 (N_4669,N_4185,N_4315);
xnor U4670 (N_4670,N_4126,N_4218);
or U4671 (N_4671,N_4129,N_4014);
and U4672 (N_4672,N_4241,N_4398);
and U4673 (N_4673,N_4060,N_4034);
and U4674 (N_4674,N_4258,N_4492);
and U4675 (N_4675,N_4267,N_4231);
nor U4676 (N_4676,N_4234,N_4124);
nand U4677 (N_4677,N_4289,N_4408);
nand U4678 (N_4678,N_4488,N_4421);
or U4679 (N_4679,N_4176,N_4482);
xnor U4680 (N_4680,N_4331,N_4116);
xor U4681 (N_4681,N_4029,N_4360);
or U4682 (N_4682,N_4159,N_4148);
and U4683 (N_4683,N_4419,N_4160);
xor U4684 (N_4684,N_4069,N_4357);
xnor U4685 (N_4685,N_4308,N_4261);
and U4686 (N_4686,N_4189,N_4423);
nand U4687 (N_4687,N_4373,N_4165);
nor U4688 (N_4688,N_4187,N_4190);
xnor U4689 (N_4689,N_4209,N_4137);
nor U4690 (N_4690,N_4193,N_4230);
xnor U4691 (N_4691,N_4364,N_4303);
or U4692 (N_4692,N_4460,N_4316);
and U4693 (N_4693,N_4220,N_4075);
nor U4694 (N_4694,N_4397,N_4214);
xnor U4695 (N_4695,N_4021,N_4462);
nor U4696 (N_4696,N_4041,N_4067);
xor U4697 (N_4697,N_4058,N_4276);
and U4698 (N_4698,N_4223,N_4410);
or U4699 (N_4699,N_4018,N_4432);
xnor U4700 (N_4700,N_4341,N_4496);
nor U4701 (N_4701,N_4054,N_4068);
xor U4702 (N_4702,N_4499,N_4199);
nor U4703 (N_4703,N_4040,N_4244);
or U4704 (N_4704,N_4447,N_4082);
or U4705 (N_4705,N_4038,N_4191);
and U4706 (N_4706,N_4283,N_4219);
or U4707 (N_4707,N_4425,N_4184);
nand U4708 (N_4708,N_4107,N_4141);
nor U4709 (N_4709,N_4361,N_4222);
nor U4710 (N_4710,N_4031,N_4133);
or U4711 (N_4711,N_4332,N_4277);
nand U4712 (N_4712,N_4396,N_4371);
or U4713 (N_4713,N_4310,N_4030);
xor U4714 (N_4714,N_4023,N_4450);
and U4715 (N_4715,N_4134,N_4007);
and U4716 (N_4716,N_4046,N_4491);
nand U4717 (N_4717,N_4048,N_4010);
nor U4718 (N_4718,N_4424,N_4147);
or U4719 (N_4719,N_4476,N_4299);
or U4720 (N_4720,N_4072,N_4171);
nor U4721 (N_4721,N_4405,N_4121);
nor U4722 (N_4722,N_4091,N_4285);
xnor U4723 (N_4723,N_4334,N_4330);
nand U4724 (N_4724,N_4096,N_4130);
and U4725 (N_4725,N_4417,N_4385);
nand U4726 (N_4726,N_4117,N_4162);
and U4727 (N_4727,N_4140,N_4333);
xnor U4728 (N_4728,N_4103,N_4224);
xor U4729 (N_4729,N_4004,N_4077);
nor U4730 (N_4730,N_4188,N_4369);
nor U4731 (N_4731,N_4433,N_4295);
or U4732 (N_4732,N_4467,N_4312);
nor U4733 (N_4733,N_4232,N_4349);
nor U4734 (N_4734,N_4484,N_4009);
and U4735 (N_4735,N_4101,N_4028);
nand U4736 (N_4736,N_4439,N_4485);
nor U4737 (N_4737,N_4081,N_4440);
nand U4738 (N_4738,N_4125,N_4181);
xnor U4739 (N_4739,N_4359,N_4351);
and U4740 (N_4740,N_4392,N_4033);
nand U4741 (N_4741,N_4006,N_4196);
nor U4742 (N_4742,N_4362,N_4468);
nand U4743 (N_4743,N_4255,N_4322);
nor U4744 (N_4744,N_4200,N_4479);
nand U4745 (N_4745,N_4325,N_4032);
nand U4746 (N_4746,N_4473,N_4097);
xnor U4747 (N_4747,N_4178,N_4345);
nor U4748 (N_4748,N_4321,N_4208);
xnor U4749 (N_4749,N_4237,N_4235);
or U4750 (N_4750,N_4174,N_4476);
and U4751 (N_4751,N_4288,N_4160);
and U4752 (N_4752,N_4364,N_4144);
nand U4753 (N_4753,N_4087,N_4006);
and U4754 (N_4754,N_4004,N_4309);
nor U4755 (N_4755,N_4334,N_4243);
nor U4756 (N_4756,N_4205,N_4086);
xor U4757 (N_4757,N_4093,N_4133);
xnor U4758 (N_4758,N_4013,N_4480);
xor U4759 (N_4759,N_4248,N_4206);
xor U4760 (N_4760,N_4331,N_4303);
nand U4761 (N_4761,N_4253,N_4336);
or U4762 (N_4762,N_4173,N_4181);
and U4763 (N_4763,N_4127,N_4252);
nor U4764 (N_4764,N_4278,N_4070);
nor U4765 (N_4765,N_4119,N_4112);
nor U4766 (N_4766,N_4392,N_4354);
nand U4767 (N_4767,N_4038,N_4224);
xor U4768 (N_4768,N_4421,N_4270);
or U4769 (N_4769,N_4352,N_4294);
xor U4770 (N_4770,N_4262,N_4134);
xnor U4771 (N_4771,N_4173,N_4390);
and U4772 (N_4772,N_4402,N_4060);
nand U4773 (N_4773,N_4241,N_4084);
and U4774 (N_4774,N_4012,N_4083);
nand U4775 (N_4775,N_4442,N_4139);
xor U4776 (N_4776,N_4154,N_4024);
and U4777 (N_4777,N_4276,N_4483);
and U4778 (N_4778,N_4394,N_4210);
nand U4779 (N_4779,N_4084,N_4365);
or U4780 (N_4780,N_4083,N_4069);
or U4781 (N_4781,N_4216,N_4119);
xor U4782 (N_4782,N_4343,N_4406);
nor U4783 (N_4783,N_4454,N_4099);
nor U4784 (N_4784,N_4331,N_4432);
xor U4785 (N_4785,N_4253,N_4110);
or U4786 (N_4786,N_4085,N_4028);
xnor U4787 (N_4787,N_4206,N_4225);
nor U4788 (N_4788,N_4484,N_4239);
xor U4789 (N_4789,N_4237,N_4189);
xor U4790 (N_4790,N_4365,N_4432);
nor U4791 (N_4791,N_4051,N_4236);
nand U4792 (N_4792,N_4306,N_4230);
nor U4793 (N_4793,N_4483,N_4094);
xor U4794 (N_4794,N_4450,N_4347);
nand U4795 (N_4795,N_4351,N_4062);
and U4796 (N_4796,N_4356,N_4453);
or U4797 (N_4797,N_4413,N_4498);
and U4798 (N_4798,N_4095,N_4046);
nor U4799 (N_4799,N_4292,N_4059);
nand U4800 (N_4800,N_4074,N_4137);
and U4801 (N_4801,N_4089,N_4122);
or U4802 (N_4802,N_4265,N_4401);
or U4803 (N_4803,N_4249,N_4153);
or U4804 (N_4804,N_4133,N_4355);
nand U4805 (N_4805,N_4420,N_4025);
and U4806 (N_4806,N_4398,N_4000);
or U4807 (N_4807,N_4001,N_4297);
or U4808 (N_4808,N_4413,N_4041);
nor U4809 (N_4809,N_4112,N_4050);
and U4810 (N_4810,N_4430,N_4217);
nor U4811 (N_4811,N_4298,N_4331);
nor U4812 (N_4812,N_4168,N_4417);
nor U4813 (N_4813,N_4081,N_4068);
xor U4814 (N_4814,N_4323,N_4042);
and U4815 (N_4815,N_4142,N_4454);
nand U4816 (N_4816,N_4373,N_4408);
xnor U4817 (N_4817,N_4166,N_4088);
and U4818 (N_4818,N_4271,N_4470);
nor U4819 (N_4819,N_4385,N_4006);
xor U4820 (N_4820,N_4040,N_4154);
or U4821 (N_4821,N_4453,N_4033);
nand U4822 (N_4822,N_4437,N_4313);
xnor U4823 (N_4823,N_4470,N_4248);
xnor U4824 (N_4824,N_4297,N_4481);
and U4825 (N_4825,N_4037,N_4193);
and U4826 (N_4826,N_4126,N_4348);
xor U4827 (N_4827,N_4063,N_4259);
nand U4828 (N_4828,N_4382,N_4023);
and U4829 (N_4829,N_4038,N_4085);
nand U4830 (N_4830,N_4347,N_4315);
or U4831 (N_4831,N_4457,N_4150);
xnor U4832 (N_4832,N_4309,N_4110);
nand U4833 (N_4833,N_4046,N_4313);
and U4834 (N_4834,N_4373,N_4316);
nor U4835 (N_4835,N_4217,N_4147);
nand U4836 (N_4836,N_4421,N_4321);
nand U4837 (N_4837,N_4204,N_4439);
xnor U4838 (N_4838,N_4188,N_4384);
and U4839 (N_4839,N_4391,N_4316);
nand U4840 (N_4840,N_4383,N_4104);
nand U4841 (N_4841,N_4172,N_4314);
nor U4842 (N_4842,N_4224,N_4203);
nor U4843 (N_4843,N_4414,N_4006);
or U4844 (N_4844,N_4057,N_4410);
xnor U4845 (N_4845,N_4342,N_4439);
nand U4846 (N_4846,N_4349,N_4237);
and U4847 (N_4847,N_4081,N_4284);
or U4848 (N_4848,N_4440,N_4441);
or U4849 (N_4849,N_4244,N_4150);
nand U4850 (N_4850,N_4374,N_4283);
nor U4851 (N_4851,N_4274,N_4086);
or U4852 (N_4852,N_4227,N_4105);
nor U4853 (N_4853,N_4307,N_4119);
and U4854 (N_4854,N_4300,N_4427);
and U4855 (N_4855,N_4084,N_4116);
nor U4856 (N_4856,N_4395,N_4249);
or U4857 (N_4857,N_4449,N_4329);
or U4858 (N_4858,N_4484,N_4316);
and U4859 (N_4859,N_4256,N_4247);
nand U4860 (N_4860,N_4397,N_4254);
nor U4861 (N_4861,N_4138,N_4070);
or U4862 (N_4862,N_4226,N_4476);
nand U4863 (N_4863,N_4075,N_4413);
nand U4864 (N_4864,N_4436,N_4280);
xor U4865 (N_4865,N_4226,N_4365);
xor U4866 (N_4866,N_4358,N_4328);
or U4867 (N_4867,N_4031,N_4191);
and U4868 (N_4868,N_4479,N_4017);
xnor U4869 (N_4869,N_4063,N_4171);
nor U4870 (N_4870,N_4464,N_4195);
and U4871 (N_4871,N_4381,N_4064);
nand U4872 (N_4872,N_4292,N_4466);
nand U4873 (N_4873,N_4323,N_4354);
or U4874 (N_4874,N_4174,N_4149);
or U4875 (N_4875,N_4264,N_4023);
or U4876 (N_4876,N_4304,N_4155);
or U4877 (N_4877,N_4332,N_4446);
or U4878 (N_4878,N_4242,N_4170);
and U4879 (N_4879,N_4295,N_4001);
and U4880 (N_4880,N_4199,N_4254);
nor U4881 (N_4881,N_4012,N_4109);
nand U4882 (N_4882,N_4119,N_4219);
nor U4883 (N_4883,N_4094,N_4166);
xor U4884 (N_4884,N_4290,N_4251);
and U4885 (N_4885,N_4399,N_4119);
or U4886 (N_4886,N_4465,N_4269);
and U4887 (N_4887,N_4080,N_4199);
xnor U4888 (N_4888,N_4301,N_4104);
nand U4889 (N_4889,N_4142,N_4328);
or U4890 (N_4890,N_4171,N_4284);
nor U4891 (N_4891,N_4055,N_4070);
nand U4892 (N_4892,N_4262,N_4304);
nor U4893 (N_4893,N_4206,N_4474);
or U4894 (N_4894,N_4364,N_4390);
nand U4895 (N_4895,N_4227,N_4315);
nand U4896 (N_4896,N_4485,N_4014);
xnor U4897 (N_4897,N_4246,N_4282);
nor U4898 (N_4898,N_4445,N_4206);
and U4899 (N_4899,N_4492,N_4323);
nor U4900 (N_4900,N_4063,N_4147);
and U4901 (N_4901,N_4461,N_4378);
nand U4902 (N_4902,N_4312,N_4050);
or U4903 (N_4903,N_4022,N_4375);
or U4904 (N_4904,N_4374,N_4115);
xor U4905 (N_4905,N_4344,N_4146);
or U4906 (N_4906,N_4417,N_4158);
or U4907 (N_4907,N_4375,N_4352);
or U4908 (N_4908,N_4204,N_4209);
nor U4909 (N_4909,N_4431,N_4295);
nand U4910 (N_4910,N_4293,N_4227);
xnor U4911 (N_4911,N_4285,N_4040);
xor U4912 (N_4912,N_4388,N_4235);
or U4913 (N_4913,N_4347,N_4442);
nand U4914 (N_4914,N_4406,N_4247);
or U4915 (N_4915,N_4485,N_4220);
nor U4916 (N_4916,N_4358,N_4341);
nor U4917 (N_4917,N_4247,N_4455);
nand U4918 (N_4918,N_4375,N_4370);
nand U4919 (N_4919,N_4099,N_4381);
xor U4920 (N_4920,N_4261,N_4177);
nor U4921 (N_4921,N_4419,N_4491);
nor U4922 (N_4922,N_4068,N_4404);
nand U4923 (N_4923,N_4474,N_4158);
and U4924 (N_4924,N_4234,N_4056);
xnor U4925 (N_4925,N_4095,N_4426);
xnor U4926 (N_4926,N_4138,N_4281);
and U4927 (N_4927,N_4345,N_4187);
nor U4928 (N_4928,N_4456,N_4449);
and U4929 (N_4929,N_4071,N_4036);
and U4930 (N_4930,N_4215,N_4109);
or U4931 (N_4931,N_4409,N_4114);
or U4932 (N_4932,N_4081,N_4044);
or U4933 (N_4933,N_4399,N_4323);
and U4934 (N_4934,N_4471,N_4110);
nand U4935 (N_4935,N_4271,N_4444);
and U4936 (N_4936,N_4040,N_4134);
or U4937 (N_4937,N_4458,N_4256);
and U4938 (N_4938,N_4237,N_4152);
and U4939 (N_4939,N_4350,N_4212);
nor U4940 (N_4940,N_4032,N_4185);
or U4941 (N_4941,N_4491,N_4308);
and U4942 (N_4942,N_4185,N_4342);
nor U4943 (N_4943,N_4172,N_4108);
and U4944 (N_4944,N_4012,N_4088);
nor U4945 (N_4945,N_4252,N_4038);
nor U4946 (N_4946,N_4373,N_4471);
xor U4947 (N_4947,N_4226,N_4182);
xor U4948 (N_4948,N_4351,N_4051);
xor U4949 (N_4949,N_4312,N_4140);
and U4950 (N_4950,N_4329,N_4139);
xor U4951 (N_4951,N_4166,N_4307);
or U4952 (N_4952,N_4412,N_4226);
nor U4953 (N_4953,N_4288,N_4083);
and U4954 (N_4954,N_4196,N_4107);
nor U4955 (N_4955,N_4477,N_4145);
nand U4956 (N_4956,N_4316,N_4395);
nand U4957 (N_4957,N_4284,N_4046);
nor U4958 (N_4958,N_4141,N_4205);
nor U4959 (N_4959,N_4230,N_4196);
or U4960 (N_4960,N_4306,N_4075);
nor U4961 (N_4961,N_4471,N_4257);
or U4962 (N_4962,N_4052,N_4379);
xor U4963 (N_4963,N_4210,N_4073);
nand U4964 (N_4964,N_4453,N_4150);
nor U4965 (N_4965,N_4453,N_4380);
xor U4966 (N_4966,N_4018,N_4259);
xor U4967 (N_4967,N_4387,N_4066);
xnor U4968 (N_4968,N_4108,N_4308);
and U4969 (N_4969,N_4446,N_4021);
xor U4970 (N_4970,N_4053,N_4060);
nand U4971 (N_4971,N_4490,N_4131);
nand U4972 (N_4972,N_4139,N_4124);
and U4973 (N_4973,N_4304,N_4288);
nor U4974 (N_4974,N_4381,N_4132);
xor U4975 (N_4975,N_4367,N_4027);
nor U4976 (N_4976,N_4429,N_4233);
or U4977 (N_4977,N_4334,N_4409);
nor U4978 (N_4978,N_4185,N_4175);
or U4979 (N_4979,N_4188,N_4264);
xor U4980 (N_4980,N_4427,N_4414);
or U4981 (N_4981,N_4172,N_4234);
nand U4982 (N_4982,N_4210,N_4191);
nand U4983 (N_4983,N_4329,N_4138);
xor U4984 (N_4984,N_4132,N_4177);
and U4985 (N_4985,N_4173,N_4178);
and U4986 (N_4986,N_4178,N_4024);
xnor U4987 (N_4987,N_4458,N_4432);
nand U4988 (N_4988,N_4299,N_4099);
nor U4989 (N_4989,N_4154,N_4479);
nor U4990 (N_4990,N_4470,N_4143);
or U4991 (N_4991,N_4058,N_4450);
or U4992 (N_4992,N_4255,N_4221);
nor U4993 (N_4993,N_4280,N_4076);
or U4994 (N_4994,N_4349,N_4151);
and U4995 (N_4995,N_4250,N_4075);
and U4996 (N_4996,N_4339,N_4360);
xor U4997 (N_4997,N_4167,N_4213);
or U4998 (N_4998,N_4352,N_4259);
or U4999 (N_4999,N_4031,N_4041);
nand UO_0 (O_0,N_4547,N_4723);
xor UO_1 (O_1,N_4875,N_4678);
and UO_2 (O_2,N_4638,N_4615);
nor UO_3 (O_3,N_4741,N_4581);
nand UO_4 (O_4,N_4718,N_4505);
nor UO_5 (O_5,N_4567,N_4591);
and UO_6 (O_6,N_4577,N_4710);
nand UO_7 (O_7,N_4663,N_4646);
and UO_8 (O_8,N_4773,N_4534);
nand UO_9 (O_9,N_4884,N_4622);
or UO_10 (O_10,N_4636,N_4780);
and UO_11 (O_11,N_4905,N_4533);
or UO_12 (O_12,N_4782,N_4664);
nand UO_13 (O_13,N_4565,N_4894);
nand UO_14 (O_14,N_4624,N_4883);
and UO_15 (O_15,N_4521,N_4778);
and UO_16 (O_16,N_4698,N_4815);
or UO_17 (O_17,N_4775,N_4506);
and UO_18 (O_18,N_4938,N_4789);
or UO_19 (O_19,N_4986,N_4604);
nor UO_20 (O_20,N_4525,N_4669);
nand UO_21 (O_21,N_4770,N_4966);
or UO_22 (O_22,N_4602,N_4803);
nand UO_23 (O_23,N_4657,N_4955);
or UO_24 (O_24,N_4626,N_4942);
or UO_25 (O_25,N_4554,N_4779);
or UO_26 (O_26,N_4720,N_4732);
or UO_27 (O_27,N_4627,N_4594);
and UO_28 (O_28,N_4765,N_4761);
xnor UO_29 (O_29,N_4630,N_4569);
nand UO_30 (O_30,N_4724,N_4980);
or UO_31 (O_31,N_4994,N_4589);
xnor UO_32 (O_32,N_4650,N_4520);
nand UO_33 (O_33,N_4617,N_4914);
xor UO_34 (O_34,N_4674,N_4628);
nor UO_35 (O_35,N_4508,N_4652);
nand UO_36 (O_36,N_4595,N_4576);
nand UO_37 (O_37,N_4848,N_4606);
xor UO_38 (O_38,N_4828,N_4635);
and UO_39 (O_39,N_4748,N_4822);
xor UO_40 (O_40,N_4964,N_4693);
nand UO_41 (O_41,N_4965,N_4609);
xnor UO_42 (O_42,N_4621,N_4768);
xnor UO_43 (O_43,N_4578,N_4574);
and UO_44 (O_44,N_4679,N_4662);
or UO_45 (O_45,N_4752,N_4756);
xnor UO_46 (O_46,N_4751,N_4542);
nand UO_47 (O_47,N_4960,N_4537);
xnor UO_48 (O_48,N_4692,N_4642);
xor UO_49 (O_49,N_4711,N_4629);
nand UO_50 (O_50,N_4504,N_4551);
xor UO_51 (O_51,N_4561,N_4827);
nor UO_52 (O_52,N_4631,N_4854);
xnor UO_53 (O_53,N_4699,N_4946);
and UO_54 (O_54,N_4880,N_4634);
and UO_55 (O_55,N_4833,N_4536);
and UO_56 (O_56,N_4730,N_4516);
or UO_57 (O_57,N_4917,N_4588);
or UO_58 (O_58,N_4683,N_4998);
nand UO_59 (O_59,N_4802,N_4898);
nor UO_60 (O_60,N_4763,N_4715);
xor UO_61 (O_61,N_4788,N_4546);
nor UO_62 (O_62,N_4614,N_4685);
nor UO_63 (O_63,N_4835,N_4941);
and UO_64 (O_64,N_4840,N_4997);
or UO_65 (O_65,N_4821,N_4807);
or UO_66 (O_66,N_4540,N_4952);
nor UO_67 (O_67,N_4605,N_4743);
nand UO_68 (O_68,N_4819,N_4781);
nor UO_69 (O_69,N_4543,N_4675);
nor UO_70 (O_70,N_4535,N_4936);
nand UO_71 (O_71,N_4906,N_4859);
nor UO_72 (O_72,N_4796,N_4769);
and UO_73 (O_73,N_4616,N_4793);
nor UO_74 (O_74,N_4611,N_4868);
xnor UO_75 (O_75,N_4957,N_4697);
nand UO_76 (O_76,N_4947,N_4882);
nand UO_77 (O_77,N_4579,N_4747);
nor UO_78 (O_78,N_4829,N_4907);
nand UO_79 (O_79,N_4680,N_4864);
nor UO_80 (O_80,N_4716,N_4794);
and UO_81 (O_81,N_4590,N_4910);
nor UO_82 (O_82,N_4772,N_4943);
or UO_83 (O_83,N_4737,N_4786);
and UO_84 (O_84,N_4745,N_4904);
xor UO_85 (O_85,N_4700,N_4517);
nand UO_86 (O_86,N_4707,N_4774);
nor UO_87 (O_87,N_4948,N_4839);
or UO_88 (O_88,N_4637,N_4860);
nand UO_89 (O_89,N_4701,N_4872);
nand UO_90 (O_90,N_4584,N_4870);
nand UO_91 (O_91,N_4552,N_4528);
nand UO_92 (O_92,N_4593,N_4983);
nor UO_93 (O_93,N_4689,N_4961);
nand UO_94 (O_94,N_4726,N_4867);
nor UO_95 (O_95,N_4978,N_4973);
or UO_96 (O_96,N_4931,N_4513);
or UO_97 (O_97,N_4953,N_4792);
nor UO_98 (O_98,N_4580,N_4668);
and UO_99 (O_99,N_4811,N_4672);
nand UO_100 (O_100,N_4735,N_4874);
xor UO_101 (O_101,N_4509,N_4923);
nand UO_102 (O_102,N_4596,N_4977);
and UO_103 (O_103,N_4995,N_4556);
nand UO_104 (O_104,N_4808,N_4721);
nand UO_105 (O_105,N_4785,N_4688);
nand UO_106 (O_106,N_4645,N_4939);
nand UO_107 (O_107,N_4991,N_4684);
or UO_108 (O_108,N_4641,N_4510);
nand UO_109 (O_109,N_4557,N_4687);
or UO_110 (O_110,N_4930,N_4703);
and UO_111 (O_111,N_4826,N_4597);
and UO_112 (O_112,N_4690,N_4963);
or UO_113 (O_113,N_4704,N_4676);
xnor UO_114 (O_114,N_4824,N_4503);
or UO_115 (O_115,N_4992,N_4836);
nand UO_116 (O_116,N_4522,N_4893);
and UO_117 (O_117,N_4967,N_4575);
nor UO_118 (O_118,N_4853,N_4601);
and UO_119 (O_119,N_4981,N_4816);
and UO_120 (O_120,N_4862,N_4787);
nor UO_121 (O_121,N_4670,N_4759);
xor UO_122 (O_122,N_4795,N_4764);
and UO_123 (O_123,N_4585,N_4661);
xor UO_124 (O_124,N_4921,N_4784);
nand UO_125 (O_125,N_4909,N_4832);
or UO_126 (O_126,N_4996,N_4640);
and UO_127 (O_127,N_4878,N_4744);
or UO_128 (O_128,N_4753,N_4544);
xnor UO_129 (O_129,N_4813,N_4924);
and UO_130 (O_130,N_4705,N_4845);
nand UO_131 (O_131,N_4681,N_4582);
nand UO_132 (O_132,N_4993,N_4886);
and UO_133 (O_133,N_4916,N_4812);
nand UO_134 (O_134,N_4654,N_4709);
nand UO_135 (O_135,N_4559,N_4933);
xor UO_136 (O_136,N_4929,N_4990);
nor UO_137 (O_137,N_4856,N_4771);
nor UO_138 (O_138,N_4830,N_4975);
nand UO_139 (O_139,N_4648,N_4666);
nand UO_140 (O_140,N_4527,N_4889);
nand UO_141 (O_141,N_4740,N_4857);
nor UO_142 (O_142,N_4541,N_4702);
nand UO_143 (O_143,N_4600,N_4651);
nor UO_144 (O_144,N_4838,N_4956);
and UO_145 (O_145,N_4568,N_4712);
nand UO_146 (O_146,N_4608,N_4750);
xor UO_147 (O_147,N_4665,N_4810);
and UO_148 (O_148,N_4958,N_4817);
xor UO_149 (O_149,N_4677,N_4927);
nor UO_150 (O_150,N_4694,N_4691);
nor UO_151 (O_151,N_4866,N_4831);
and UO_152 (O_152,N_4937,N_4644);
and UO_153 (O_153,N_4500,N_4599);
nand UO_154 (O_154,N_4970,N_4954);
or UO_155 (O_155,N_4850,N_4982);
xor UO_156 (O_156,N_4800,N_4842);
and UO_157 (O_157,N_4887,N_4797);
nand UO_158 (O_158,N_4852,N_4524);
nand UO_159 (O_159,N_4671,N_4555);
xnor UO_160 (O_160,N_4545,N_4949);
or UO_161 (O_161,N_4731,N_4865);
nand UO_162 (O_162,N_4639,N_4777);
and UO_163 (O_163,N_4610,N_4655);
nand UO_164 (O_164,N_4658,N_4548);
nor UO_165 (O_165,N_4951,N_4550);
xnor UO_166 (O_166,N_4834,N_4592);
or UO_167 (O_167,N_4915,N_4901);
or UO_168 (O_168,N_4754,N_4526);
nand UO_169 (O_169,N_4729,N_4790);
nor UO_170 (O_170,N_4733,N_4673);
or UO_171 (O_171,N_4888,N_4935);
nand UO_172 (O_172,N_4656,N_4598);
and UO_173 (O_173,N_4871,N_4686);
nand UO_174 (O_174,N_4519,N_4767);
and UO_175 (O_175,N_4728,N_4749);
nor UO_176 (O_176,N_4653,N_4890);
nor UO_177 (O_177,N_4620,N_4783);
or UO_178 (O_178,N_4739,N_4719);
or UO_179 (O_179,N_4612,N_4563);
xor UO_180 (O_180,N_4558,N_4846);
nor UO_181 (O_181,N_4518,N_4932);
or UO_182 (O_182,N_4523,N_4757);
nand UO_183 (O_183,N_4607,N_4667);
nor UO_184 (O_184,N_4897,N_4549);
or UO_185 (O_185,N_4571,N_4979);
nand UO_186 (O_186,N_4633,N_4891);
nand UO_187 (O_187,N_4649,N_4892);
xnor UO_188 (O_188,N_4804,N_4573);
xnor UO_189 (O_189,N_4515,N_4799);
or UO_190 (O_190,N_4881,N_4643);
nor UO_191 (O_191,N_4805,N_4911);
xor UO_192 (O_192,N_4908,N_4972);
xnor UO_193 (O_193,N_4861,N_4706);
or UO_194 (O_194,N_4776,N_4974);
nand UO_195 (O_195,N_4849,N_4959);
nand UO_196 (O_196,N_4851,N_4841);
nor UO_197 (O_197,N_4798,N_4843);
and UO_198 (O_198,N_4945,N_4950);
nand UO_199 (O_199,N_4876,N_4603);
nand UO_200 (O_200,N_4879,N_4847);
nand UO_201 (O_201,N_4806,N_4746);
or UO_202 (O_202,N_4507,N_4758);
xnor UO_203 (O_203,N_4885,N_4660);
or UO_204 (O_204,N_4877,N_4722);
nor UO_205 (O_205,N_4825,N_4714);
nand UO_206 (O_206,N_4988,N_4944);
and UO_207 (O_207,N_4562,N_4999);
or UO_208 (O_208,N_4619,N_4919);
xnor UO_209 (O_209,N_4863,N_4586);
nor UO_210 (O_210,N_4736,N_4682);
and UO_211 (O_211,N_4734,N_4985);
or UO_212 (O_212,N_4962,N_4858);
xnor UO_213 (O_213,N_4902,N_4708);
or UO_214 (O_214,N_4583,N_4738);
nor UO_215 (O_215,N_4530,N_4514);
and UO_216 (O_216,N_4502,N_4566);
xnor UO_217 (O_217,N_4989,N_4532);
or UO_218 (O_218,N_4895,N_4968);
or UO_219 (O_219,N_4940,N_4766);
nor UO_220 (O_220,N_4837,N_4755);
nor UO_221 (O_221,N_4553,N_4934);
and UO_222 (O_222,N_4912,N_4529);
nor UO_223 (O_223,N_4613,N_4928);
or UO_224 (O_224,N_4713,N_4922);
nand UO_225 (O_225,N_4969,N_4791);
or UO_226 (O_226,N_4618,N_4623);
or UO_227 (O_227,N_4560,N_4873);
nand UO_228 (O_228,N_4727,N_4900);
and UO_229 (O_229,N_4903,N_4564);
nor UO_230 (O_230,N_4984,N_4570);
nand UO_231 (O_231,N_4760,N_4844);
xnor UO_232 (O_232,N_4539,N_4538);
xor UO_233 (O_233,N_4725,N_4918);
and UO_234 (O_234,N_4814,N_4572);
nor UO_235 (O_235,N_4925,N_4647);
or UO_236 (O_236,N_4625,N_4695);
or UO_237 (O_237,N_4587,N_4899);
xnor UO_238 (O_238,N_4762,N_4632);
xnor UO_239 (O_239,N_4913,N_4971);
nand UO_240 (O_240,N_4717,N_4926);
xor UO_241 (O_241,N_4920,N_4869);
xor UO_242 (O_242,N_4818,N_4809);
or UO_243 (O_243,N_4987,N_4659);
and UO_244 (O_244,N_4823,N_4696);
nor UO_245 (O_245,N_4820,N_4976);
nor UO_246 (O_246,N_4896,N_4511);
or UO_247 (O_247,N_4801,N_4531);
xor UO_248 (O_248,N_4855,N_4512);
xnor UO_249 (O_249,N_4501,N_4742);
nand UO_250 (O_250,N_4696,N_4882);
and UO_251 (O_251,N_4972,N_4598);
nand UO_252 (O_252,N_4795,N_4647);
xor UO_253 (O_253,N_4843,N_4661);
nand UO_254 (O_254,N_4710,N_4835);
nand UO_255 (O_255,N_4714,N_4785);
nor UO_256 (O_256,N_4924,N_4606);
nor UO_257 (O_257,N_4742,N_4847);
nand UO_258 (O_258,N_4902,N_4901);
xnor UO_259 (O_259,N_4909,N_4539);
and UO_260 (O_260,N_4725,N_4658);
and UO_261 (O_261,N_4871,N_4518);
nand UO_262 (O_262,N_4581,N_4818);
nand UO_263 (O_263,N_4540,N_4602);
or UO_264 (O_264,N_4562,N_4959);
or UO_265 (O_265,N_4730,N_4934);
xor UO_266 (O_266,N_4986,N_4922);
or UO_267 (O_267,N_4937,N_4979);
xnor UO_268 (O_268,N_4900,N_4568);
nand UO_269 (O_269,N_4916,N_4672);
or UO_270 (O_270,N_4994,N_4854);
and UO_271 (O_271,N_4801,N_4558);
and UO_272 (O_272,N_4623,N_4814);
or UO_273 (O_273,N_4673,N_4519);
nand UO_274 (O_274,N_4664,N_4737);
or UO_275 (O_275,N_4969,N_4736);
nor UO_276 (O_276,N_4958,N_4512);
or UO_277 (O_277,N_4522,N_4513);
or UO_278 (O_278,N_4862,N_4846);
xnor UO_279 (O_279,N_4969,N_4751);
xor UO_280 (O_280,N_4964,N_4873);
nand UO_281 (O_281,N_4816,N_4891);
nand UO_282 (O_282,N_4747,N_4778);
and UO_283 (O_283,N_4879,N_4553);
xnor UO_284 (O_284,N_4796,N_4666);
nor UO_285 (O_285,N_4864,N_4653);
xnor UO_286 (O_286,N_4977,N_4537);
nand UO_287 (O_287,N_4521,N_4691);
xor UO_288 (O_288,N_4721,N_4853);
nor UO_289 (O_289,N_4950,N_4998);
and UO_290 (O_290,N_4970,N_4989);
and UO_291 (O_291,N_4590,N_4811);
or UO_292 (O_292,N_4518,N_4767);
nand UO_293 (O_293,N_4698,N_4677);
xnor UO_294 (O_294,N_4520,N_4588);
nor UO_295 (O_295,N_4692,N_4693);
nand UO_296 (O_296,N_4752,N_4727);
nor UO_297 (O_297,N_4679,N_4768);
and UO_298 (O_298,N_4639,N_4633);
or UO_299 (O_299,N_4618,N_4806);
nand UO_300 (O_300,N_4714,N_4592);
or UO_301 (O_301,N_4965,N_4859);
nand UO_302 (O_302,N_4766,N_4530);
xor UO_303 (O_303,N_4967,N_4892);
or UO_304 (O_304,N_4774,N_4772);
nand UO_305 (O_305,N_4584,N_4660);
or UO_306 (O_306,N_4531,N_4939);
nor UO_307 (O_307,N_4633,N_4595);
or UO_308 (O_308,N_4798,N_4581);
xnor UO_309 (O_309,N_4723,N_4981);
and UO_310 (O_310,N_4864,N_4925);
nand UO_311 (O_311,N_4954,N_4597);
nor UO_312 (O_312,N_4939,N_4693);
nand UO_313 (O_313,N_4513,N_4523);
nor UO_314 (O_314,N_4602,N_4627);
xor UO_315 (O_315,N_4966,N_4942);
and UO_316 (O_316,N_4920,N_4886);
or UO_317 (O_317,N_4792,N_4635);
xor UO_318 (O_318,N_4950,N_4749);
nor UO_319 (O_319,N_4863,N_4550);
nor UO_320 (O_320,N_4664,N_4647);
and UO_321 (O_321,N_4549,N_4648);
nor UO_322 (O_322,N_4545,N_4834);
xor UO_323 (O_323,N_4795,N_4846);
or UO_324 (O_324,N_4881,N_4910);
nor UO_325 (O_325,N_4696,N_4526);
or UO_326 (O_326,N_4646,N_4741);
xor UO_327 (O_327,N_4882,N_4568);
and UO_328 (O_328,N_4597,N_4907);
or UO_329 (O_329,N_4645,N_4938);
nand UO_330 (O_330,N_4916,N_4674);
or UO_331 (O_331,N_4667,N_4961);
nand UO_332 (O_332,N_4610,N_4885);
nand UO_333 (O_333,N_4754,N_4877);
and UO_334 (O_334,N_4894,N_4878);
xnor UO_335 (O_335,N_4840,N_4939);
nor UO_336 (O_336,N_4575,N_4738);
xnor UO_337 (O_337,N_4715,N_4902);
nand UO_338 (O_338,N_4871,N_4592);
or UO_339 (O_339,N_4514,N_4834);
or UO_340 (O_340,N_4716,N_4669);
nand UO_341 (O_341,N_4828,N_4683);
nand UO_342 (O_342,N_4707,N_4795);
xnor UO_343 (O_343,N_4957,N_4892);
nand UO_344 (O_344,N_4588,N_4717);
and UO_345 (O_345,N_4997,N_4550);
or UO_346 (O_346,N_4628,N_4583);
nand UO_347 (O_347,N_4936,N_4958);
xnor UO_348 (O_348,N_4919,N_4565);
nor UO_349 (O_349,N_4944,N_4507);
nand UO_350 (O_350,N_4554,N_4689);
nand UO_351 (O_351,N_4536,N_4602);
or UO_352 (O_352,N_4981,N_4806);
nand UO_353 (O_353,N_4668,N_4809);
or UO_354 (O_354,N_4870,N_4859);
or UO_355 (O_355,N_4538,N_4784);
nand UO_356 (O_356,N_4951,N_4987);
and UO_357 (O_357,N_4500,N_4582);
and UO_358 (O_358,N_4657,N_4729);
xor UO_359 (O_359,N_4747,N_4532);
nand UO_360 (O_360,N_4732,N_4882);
nor UO_361 (O_361,N_4845,N_4668);
nor UO_362 (O_362,N_4972,N_4791);
or UO_363 (O_363,N_4558,N_4730);
xnor UO_364 (O_364,N_4802,N_4961);
nor UO_365 (O_365,N_4672,N_4994);
and UO_366 (O_366,N_4583,N_4652);
xnor UO_367 (O_367,N_4582,N_4827);
nand UO_368 (O_368,N_4828,N_4558);
or UO_369 (O_369,N_4589,N_4778);
nor UO_370 (O_370,N_4931,N_4716);
and UO_371 (O_371,N_4661,N_4981);
nor UO_372 (O_372,N_4779,N_4831);
and UO_373 (O_373,N_4520,N_4573);
nor UO_374 (O_374,N_4983,N_4767);
nor UO_375 (O_375,N_4765,N_4925);
and UO_376 (O_376,N_4793,N_4637);
nor UO_377 (O_377,N_4981,N_4789);
nor UO_378 (O_378,N_4673,N_4702);
or UO_379 (O_379,N_4570,N_4794);
nor UO_380 (O_380,N_4808,N_4529);
xnor UO_381 (O_381,N_4552,N_4827);
or UO_382 (O_382,N_4881,N_4571);
xor UO_383 (O_383,N_4993,N_4931);
and UO_384 (O_384,N_4619,N_4830);
nand UO_385 (O_385,N_4518,N_4774);
nand UO_386 (O_386,N_4819,N_4666);
nor UO_387 (O_387,N_4644,N_4529);
and UO_388 (O_388,N_4572,N_4866);
nor UO_389 (O_389,N_4902,N_4785);
nor UO_390 (O_390,N_4957,N_4674);
xor UO_391 (O_391,N_4564,N_4575);
or UO_392 (O_392,N_4824,N_4927);
nand UO_393 (O_393,N_4537,N_4733);
nand UO_394 (O_394,N_4700,N_4627);
xor UO_395 (O_395,N_4905,N_4714);
and UO_396 (O_396,N_4815,N_4699);
xor UO_397 (O_397,N_4605,N_4897);
nand UO_398 (O_398,N_4788,N_4825);
and UO_399 (O_399,N_4717,N_4531);
xor UO_400 (O_400,N_4517,N_4645);
nor UO_401 (O_401,N_4795,N_4837);
nand UO_402 (O_402,N_4801,N_4590);
or UO_403 (O_403,N_4979,N_4691);
or UO_404 (O_404,N_4762,N_4703);
nor UO_405 (O_405,N_4600,N_4620);
nor UO_406 (O_406,N_4593,N_4764);
or UO_407 (O_407,N_4946,N_4947);
nand UO_408 (O_408,N_4514,N_4835);
xnor UO_409 (O_409,N_4828,N_4572);
or UO_410 (O_410,N_4526,N_4996);
or UO_411 (O_411,N_4729,N_4867);
xor UO_412 (O_412,N_4800,N_4715);
nor UO_413 (O_413,N_4754,N_4896);
xor UO_414 (O_414,N_4937,N_4505);
and UO_415 (O_415,N_4960,N_4932);
xor UO_416 (O_416,N_4628,N_4595);
xor UO_417 (O_417,N_4818,N_4795);
xnor UO_418 (O_418,N_4590,N_4737);
and UO_419 (O_419,N_4907,N_4913);
nor UO_420 (O_420,N_4751,N_4664);
and UO_421 (O_421,N_4559,N_4687);
or UO_422 (O_422,N_4968,N_4991);
and UO_423 (O_423,N_4591,N_4619);
nand UO_424 (O_424,N_4995,N_4877);
nor UO_425 (O_425,N_4704,N_4517);
and UO_426 (O_426,N_4978,N_4954);
and UO_427 (O_427,N_4961,N_4754);
and UO_428 (O_428,N_4799,N_4732);
or UO_429 (O_429,N_4994,N_4586);
xor UO_430 (O_430,N_4954,N_4886);
nand UO_431 (O_431,N_4914,N_4990);
nand UO_432 (O_432,N_4715,N_4801);
and UO_433 (O_433,N_4876,N_4534);
or UO_434 (O_434,N_4794,N_4561);
and UO_435 (O_435,N_4580,N_4563);
nand UO_436 (O_436,N_4683,N_4617);
nor UO_437 (O_437,N_4869,N_4544);
nor UO_438 (O_438,N_4928,N_4971);
and UO_439 (O_439,N_4951,N_4958);
xor UO_440 (O_440,N_4899,N_4914);
and UO_441 (O_441,N_4954,N_4751);
nand UO_442 (O_442,N_4794,N_4582);
nand UO_443 (O_443,N_4737,N_4595);
nand UO_444 (O_444,N_4572,N_4816);
nand UO_445 (O_445,N_4843,N_4653);
nor UO_446 (O_446,N_4611,N_4517);
or UO_447 (O_447,N_4517,N_4534);
nand UO_448 (O_448,N_4782,N_4586);
xor UO_449 (O_449,N_4680,N_4971);
and UO_450 (O_450,N_4525,N_4633);
nor UO_451 (O_451,N_4759,N_4907);
or UO_452 (O_452,N_4650,N_4924);
and UO_453 (O_453,N_4628,N_4989);
xor UO_454 (O_454,N_4644,N_4810);
and UO_455 (O_455,N_4806,N_4677);
xor UO_456 (O_456,N_4986,N_4976);
xnor UO_457 (O_457,N_4681,N_4621);
and UO_458 (O_458,N_4976,N_4954);
or UO_459 (O_459,N_4594,N_4914);
nor UO_460 (O_460,N_4651,N_4661);
xor UO_461 (O_461,N_4826,N_4896);
nand UO_462 (O_462,N_4875,N_4563);
or UO_463 (O_463,N_4983,N_4966);
or UO_464 (O_464,N_4783,N_4716);
or UO_465 (O_465,N_4583,N_4716);
xnor UO_466 (O_466,N_4644,N_4849);
and UO_467 (O_467,N_4736,N_4946);
or UO_468 (O_468,N_4653,N_4791);
or UO_469 (O_469,N_4665,N_4770);
nor UO_470 (O_470,N_4503,N_4604);
and UO_471 (O_471,N_4772,N_4767);
and UO_472 (O_472,N_4668,N_4783);
nor UO_473 (O_473,N_4557,N_4935);
and UO_474 (O_474,N_4996,N_4675);
nand UO_475 (O_475,N_4760,N_4987);
or UO_476 (O_476,N_4650,N_4996);
xnor UO_477 (O_477,N_4775,N_4962);
nand UO_478 (O_478,N_4885,N_4856);
or UO_479 (O_479,N_4961,N_4731);
nand UO_480 (O_480,N_4938,N_4742);
and UO_481 (O_481,N_4998,N_4592);
nand UO_482 (O_482,N_4918,N_4645);
or UO_483 (O_483,N_4953,N_4659);
nor UO_484 (O_484,N_4541,N_4822);
nor UO_485 (O_485,N_4662,N_4572);
nand UO_486 (O_486,N_4556,N_4943);
nor UO_487 (O_487,N_4904,N_4937);
and UO_488 (O_488,N_4573,N_4541);
nor UO_489 (O_489,N_4523,N_4894);
or UO_490 (O_490,N_4795,N_4799);
nor UO_491 (O_491,N_4753,N_4816);
nor UO_492 (O_492,N_4500,N_4978);
nor UO_493 (O_493,N_4841,N_4964);
nand UO_494 (O_494,N_4887,N_4524);
and UO_495 (O_495,N_4782,N_4941);
nand UO_496 (O_496,N_4728,N_4600);
and UO_497 (O_497,N_4905,N_4599);
and UO_498 (O_498,N_4852,N_4542);
xor UO_499 (O_499,N_4886,N_4588);
xnor UO_500 (O_500,N_4732,N_4905);
and UO_501 (O_501,N_4588,N_4586);
nor UO_502 (O_502,N_4756,N_4810);
nor UO_503 (O_503,N_4985,N_4699);
or UO_504 (O_504,N_4502,N_4503);
nor UO_505 (O_505,N_4929,N_4546);
nand UO_506 (O_506,N_4621,N_4938);
nand UO_507 (O_507,N_4817,N_4781);
or UO_508 (O_508,N_4821,N_4668);
nand UO_509 (O_509,N_4582,N_4625);
or UO_510 (O_510,N_4702,N_4660);
xnor UO_511 (O_511,N_4642,N_4775);
xnor UO_512 (O_512,N_4687,N_4977);
or UO_513 (O_513,N_4844,N_4948);
or UO_514 (O_514,N_4820,N_4548);
and UO_515 (O_515,N_4744,N_4623);
nor UO_516 (O_516,N_4585,N_4987);
nor UO_517 (O_517,N_4581,N_4506);
or UO_518 (O_518,N_4884,N_4603);
nand UO_519 (O_519,N_4620,N_4719);
or UO_520 (O_520,N_4999,N_4559);
and UO_521 (O_521,N_4526,N_4746);
xnor UO_522 (O_522,N_4793,N_4758);
and UO_523 (O_523,N_4664,N_4671);
nor UO_524 (O_524,N_4863,N_4796);
and UO_525 (O_525,N_4814,N_4977);
xor UO_526 (O_526,N_4590,N_4822);
nor UO_527 (O_527,N_4693,N_4940);
nand UO_528 (O_528,N_4794,N_4924);
nor UO_529 (O_529,N_4781,N_4609);
nor UO_530 (O_530,N_4898,N_4920);
nand UO_531 (O_531,N_4506,N_4983);
nor UO_532 (O_532,N_4989,N_4788);
or UO_533 (O_533,N_4807,N_4747);
or UO_534 (O_534,N_4618,N_4877);
and UO_535 (O_535,N_4689,N_4806);
or UO_536 (O_536,N_4779,N_4901);
nor UO_537 (O_537,N_4714,N_4860);
xnor UO_538 (O_538,N_4882,N_4766);
nor UO_539 (O_539,N_4559,N_4738);
nor UO_540 (O_540,N_4737,N_4886);
nor UO_541 (O_541,N_4996,N_4610);
xnor UO_542 (O_542,N_4975,N_4963);
xor UO_543 (O_543,N_4936,N_4558);
xnor UO_544 (O_544,N_4656,N_4850);
xnor UO_545 (O_545,N_4885,N_4643);
and UO_546 (O_546,N_4618,N_4866);
and UO_547 (O_547,N_4614,N_4715);
nand UO_548 (O_548,N_4747,N_4635);
and UO_549 (O_549,N_4771,N_4528);
nand UO_550 (O_550,N_4953,N_4763);
nor UO_551 (O_551,N_4747,N_4799);
and UO_552 (O_552,N_4962,N_4854);
and UO_553 (O_553,N_4586,N_4680);
nand UO_554 (O_554,N_4821,N_4678);
nor UO_555 (O_555,N_4717,N_4748);
nand UO_556 (O_556,N_4954,N_4527);
and UO_557 (O_557,N_4503,N_4715);
and UO_558 (O_558,N_4608,N_4567);
xor UO_559 (O_559,N_4573,N_4883);
xor UO_560 (O_560,N_4764,N_4654);
nand UO_561 (O_561,N_4662,N_4776);
nand UO_562 (O_562,N_4714,N_4850);
xor UO_563 (O_563,N_4970,N_4861);
and UO_564 (O_564,N_4806,N_4736);
nand UO_565 (O_565,N_4625,N_4970);
xnor UO_566 (O_566,N_4529,N_4986);
nand UO_567 (O_567,N_4976,N_4773);
nand UO_568 (O_568,N_4787,N_4508);
nand UO_569 (O_569,N_4587,N_4862);
and UO_570 (O_570,N_4627,N_4813);
or UO_571 (O_571,N_4594,N_4929);
nor UO_572 (O_572,N_4560,N_4927);
nor UO_573 (O_573,N_4777,N_4920);
or UO_574 (O_574,N_4891,N_4726);
nand UO_575 (O_575,N_4888,N_4821);
nor UO_576 (O_576,N_4769,N_4523);
nand UO_577 (O_577,N_4671,N_4587);
xnor UO_578 (O_578,N_4546,N_4829);
and UO_579 (O_579,N_4694,N_4814);
nand UO_580 (O_580,N_4792,N_4634);
nor UO_581 (O_581,N_4754,N_4957);
xnor UO_582 (O_582,N_4747,N_4973);
nand UO_583 (O_583,N_4526,N_4902);
nor UO_584 (O_584,N_4961,N_4810);
or UO_585 (O_585,N_4941,N_4634);
nand UO_586 (O_586,N_4799,N_4939);
and UO_587 (O_587,N_4981,N_4655);
nand UO_588 (O_588,N_4772,N_4986);
or UO_589 (O_589,N_4842,N_4823);
nand UO_590 (O_590,N_4804,N_4953);
xnor UO_591 (O_591,N_4994,N_4735);
or UO_592 (O_592,N_4791,N_4959);
nand UO_593 (O_593,N_4502,N_4579);
nor UO_594 (O_594,N_4783,N_4573);
nand UO_595 (O_595,N_4652,N_4854);
xor UO_596 (O_596,N_4980,N_4599);
nand UO_597 (O_597,N_4991,N_4606);
xnor UO_598 (O_598,N_4612,N_4718);
nor UO_599 (O_599,N_4778,N_4803);
and UO_600 (O_600,N_4904,N_4658);
nor UO_601 (O_601,N_4657,N_4718);
xor UO_602 (O_602,N_4524,N_4760);
xor UO_603 (O_603,N_4876,N_4522);
or UO_604 (O_604,N_4980,N_4674);
or UO_605 (O_605,N_4543,N_4537);
xnor UO_606 (O_606,N_4701,N_4939);
or UO_607 (O_607,N_4512,N_4999);
or UO_608 (O_608,N_4814,N_4979);
nor UO_609 (O_609,N_4698,N_4914);
nand UO_610 (O_610,N_4768,N_4956);
or UO_611 (O_611,N_4747,N_4731);
nor UO_612 (O_612,N_4888,N_4840);
and UO_613 (O_613,N_4774,N_4829);
nand UO_614 (O_614,N_4601,N_4808);
nand UO_615 (O_615,N_4773,N_4752);
or UO_616 (O_616,N_4963,N_4839);
xnor UO_617 (O_617,N_4569,N_4682);
xnor UO_618 (O_618,N_4983,N_4772);
nor UO_619 (O_619,N_4847,N_4880);
and UO_620 (O_620,N_4594,N_4908);
xnor UO_621 (O_621,N_4586,N_4739);
or UO_622 (O_622,N_4598,N_4576);
nor UO_623 (O_623,N_4698,N_4817);
or UO_624 (O_624,N_4676,N_4813);
xnor UO_625 (O_625,N_4745,N_4750);
nand UO_626 (O_626,N_4862,N_4683);
xnor UO_627 (O_627,N_4630,N_4758);
and UO_628 (O_628,N_4751,N_4666);
xnor UO_629 (O_629,N_4596,N_4798);
nor UO_630 (O_630,N_4889,N_4724);
or UO_631 (O_631,N_4640,N_4690);
and UO_632 (O_632,N_4563,N_4551);
nand UO_633 (O_633,N_4868,N_4582);
nor UO_634 (O_634,N_4960,N_4564);
and UO_635 (O_635,N_4511,N_4735);
nand UO_636 (O_636,N_4522,N_4666);
nor UO_637 (O_637,N_4708,N_4543);
nor UO_638 (O_638,N_4525,N_4539);
xnor UO_639 (O_639,N_4627,N_4684);
or UO_640 (O_640,N_4768,N_4523);
and UO_641 (O_641,N_4570,N_4561);
nand UO_642 (O_642,N_4813,N_4552);
nand UO_643 (O_643,N_4632,N_4739);
nor UO_644 (O_644,N_4732,N_4933);
and UO_645 (O_645,N_4706,N_4988);
nand UO_646 (O_646,N_4515,N_4987);
nor UO_647 (O_647,N_4986,N_4507);
and UO_648 (O_648,N_4693,N_4874);
and UO_649 (O_649,N_4750,N_4592);
xor UO_650 (O_650,N_4525,N_4794);
nor UO_651 (O_651,N_4659,N_4973);
or UO_652 (O_652,N_4760,N_4632);
xor UO_653 (O_653,N_4729,N_4616);
xor UO_654 (O_654,N_4724,N_4627);
and UO_655 (O_655,N_4992,N_4663);
nor UO_656 (O_656,N_4849,N_4744);
or UO_657 (O_657,N_4678,N_4976);
xor UO_658 (O_658,N_4508,N_4999);
nand UO_659 (O_659,N_4707,N_4694);
nor UO_660 (O_660,N_4551,N_4743);
or UO_661 (O_661,N_4839,N_4565);
or UO_662 (O_662,N_4568,N_4949);
and UO_663 (O_663,N_4791,N_4618);
nor UO_664 (O_664,N_4963,N_4746);
and UO_665 (O_665,N_4998,N_4911);
or UO_666 (O_666,N_4733,N_4868);
nor UO_667 (O_667,N_4870,N_4996);
and UO_668 (O_668,N_4674,N_4723);
xnor UO_669 (O_669,N_4783,N_4714);
and UO_670 (O_670,N_4978,N_4651);
nor UO_671 (O_671,N_4559,N_4577);
or UO_672 (O_672,N_4994,N_4865);
nor UO_673 (O_673,N_4720,N_4824);
and UO_674 (O_674,N_4722,N_4580);
and UO_675 (O_675,N_4900,N_4890);
or UO_676 (O_676,N_4812,N_4503);
nor UO_677 (O_677,N_4611,N_4971);
nand UO_678 (O_678,N_4809,N_4930);
or UO_679 (O_679,N_4613,N_4635);
nor UO_680 (O_680,N_4983,N_4981);
and UO_681 (O_681,N_4841,N_4864);
xnor UO_682 (O_682,N_4889,N_4657);
and UO_683 (O_683,N_4639,N_4625);
nand UO_684 (O_684,N_4539,N_4681);
and UO_685 (O_685,N_4714,N_4538);
xnor UO_686 (O_686,N_4904,N_4614);
xor UO_687 (O_687,N_4804,N_4771);
nand UO_688 (O_688,N_4777,N_4997);
nor UO_689 (O_689,N_4738,N_4534);
nand UO_690 (O_690,N_4743,N_4570);
xor UO_691 (O_691,N_4972,N_4752);
and UO_692 (O_692,N_4695,N_4897);
or UO_693 (O_693,N_4862,N_4956);
and UO_694 (O_694,N_4582,N_4801);
or UO_695 (O_695,N_4871,N_4558);
nand UO_696 (O_696,N_4531,N_4786);
nor UO_697 (O_697,N_4663,N_4625);
or UO_698 (O_698,N_4957,N_4765);
and UO_699 (O_699,N_4892,N_4864);
and UO_700 (O_700,N_4583,N_4846);
and UO_701 (O_701,N_4937,N_4953);
or UO_702 (O_702,N_4957,N_4877);
xor UO_703 (O_703,N_4546,N_4696);
xor UO_704 (O_704,N_4666,N_4873);
nor UO_705 (O_705,N_4906,N_4893);
or UO_706 (O_706,N_4911,N_4526);
or UO_707 (O_707,N_4554,N_4712);
nand UO_708 (O_708,N_4882,N_4512);
or UO_709 (O_709,N_4779,N_4713);
xor UO_710 (O_710,N_4863,N_4785);
or UO_711 (O_711,N_4644,N_4676);
xor UO_712 (O_712,N_4642,N_4943);
nor UO_713 (O_713,N_4970,N_4770);
nor UO_714 (O_714,N_4692,N_4771);
nand UO_715 (O_715,N_4970,N_4571);
or UO_716 (O_716,N_4785,N_4970);
nor UO_717 (O_717,N_4590,N_4921);
xnor UO_718 (O_718,N_4930,N_4926);
or UO_719 (O_719,N_4511,N_4571);
nand UO_720 (O_720,N_4810,N_4668);
nor UO_721 (O_721,N_4891,N_4687);
nor UO_722 (O_722,N_4727,N_4921);
nand UO_723 (O_723,N_4528,N_4673);
or UO_724 (O_724,N_4841,N_4776);
or UO_725 (O_725,N_4877,N_4633);
or UO_726 (O_726,N_4758,N_4591);
nand UO_727 (O_727,N_4855,N_4572);
and UO_728 (O_728,N_4611,N_4788);
nor UO_729 (O_729,N_4789,N_4838);
and UO_730 (O_730,N_4842,N_4958);
or UO_731 (O_731,N_4814,N_4704);
or UO_732 (O_732,N_4958,N_4557);
or UO_733 (O_733,N_4853,N_4546);
or UO_734 (O_734,N_4837,N_4940);
xor UO_735 (O_735,N_4809,N_4716);
and UO_736 (O_736,N_4510,N_4638);
nor UO_737 (O_737,N_4853,N_4767);
or UO_738 (O_738,N_4888,N_4733);
nand UO_739 (O_739,N_4814,N_4992);
and UO_740 (O_740,N_4786,N_4955);
or UO_741 (O_741,N_4990,N_4715);
nor UO_742 (O_742,N_4996,N_4888);
nor UO_743 (O_743,N_4666,N_4504);
nand UO_744 (O_744,N_4690,N_4943);
nor UO_745 (O_745,N_4784,N_4898);
nand UO_746 (O_746,N_4804,N_4542);
nand UO_747 (O_747,N_4511,N_4787);
or UO_748 (O_748,N_4750,N_4718);
nand UO_749 (O_749,N_4655,N_4896);
or UO_750 (O_750,N_4669,N_4921);
nand UO_751 (O_751,N_4875,N_4778);
nand UO_752 (O_752,N_4823,N_4923);
nand UO_753 (O_753,N_4890,N_4954);
nand UO_754 (O_754,N_4809,N_4568);
and UO_755 (O_755,N_4574,N_4700);
nand UO_756 (O_756,N_4546,N_4855);
or UO_757 (O_757,N_4513,N_4567);
and UO_758 (O_758,N_4850,N_4544);
nand UO_759 (O_759,N_4645,N_4816);
nor UO_760 (O_760,N_4707,N_4747);
or UO_761 (O_761,N_4928,N_4867);
nor UO_762 (O_762,N_4779,N_4975);
or UO_763 (O_763,N_4734,N_4572);
nor UO_764 (O_764,N_4509,N_4514);
nand UO_765 (O_765,N_4798,N_4508);
and UO_766 (O_766,N_4840,N_4624);
nor UO_767 (O_767,N_4972,N_4697);
xnor UO_768 (O_768,N_4624,N_4929);
nand UO_769 (O_769,N_4560,N_4886);
nand UO_770 (O_770,N_4618,N_4541);
xor UO_771 (O_771,N_4503,N_4644);
or UO_772 (O_772,N_4537,N_4898);
xor UO_773 (O_773,N_4939,N_4556);
nand UO_774 (O_774,N_4571,N_4675);
nor UO_775 (O_775,N_4574,N_4535);
xor UO_776 (O_776,N_4786,N_4518);
nand UO_777 (O_777,N_4674,N_4773);
nor UO_778 (O_778,N_4603,N_4866);
and UO_779 (O_779,N_4930,N_4553);
nor UO_780 (O_780,N_4882,N_4671);
or UO_781 (O_781,N_4895,N_4693);
and UO_782 (O_782,N_4735,N_4529);
or UO_783 (O_783,N_4920,N_4954);
nand UO_784 (O_784,N_4563,N_4510);
nor UO_785 (O_785,N_4553,N_4618);
xor UO_786 (O_786,N_4771,N_4743);
and UO_787 (O_787,N_4902,N_4709);
nor UO_788 (O_788,N_4924,N_4910);
xor UO_789 (O_789,N_4623,N_4662);
and UO_790 (O_790,N_4702,N_4609);
nand UO_791 (O_791,N_4575,N_4775);
nand UO_792 (O_792,N_4617,N_4525);
or UO_793 (O_793,N_4907,N_4556);
nor UO_794 (O_794,N_4689,N_4528);
xnor UO_795 (O_795,N_4724,N_4939);
nor UO_796 (O_796,N_4601,N_4568);
xor UO_797 (O_797,N_4892,N_4990);
nor UO_798 (O_798,N_4691,N_4628);
xnor UO_799 (O_799,N_4762,N_4992);
or UO_800 (O_800,N_4745,N_4667);
nor UO_801 (O_801,N_4931,N_4868);
nand UO_802 (O_802,N_4976,N_4689);
nand UO_803 (O_803,N_4741,N_4588);
xor UO_804 (O_804,N_4897,N_4953);
xnor UO_805 (O_805,N_4547,N_4743);
xor UO_806 (O_806,N_4891,N_4932);
nand UO_807 (O_807,N_4528,N_4732);
and UO_808 (O_808,N_4755,N_4649);
nor UO_809 (O_809,N_4854,N_4948);
nor UO_810 (O_810,N_4588,N_4637);
nand UO_811 (O_811,N_4728,N_4790);
and UO_812 (O_812,N_4593,N_4953);
or UO_813 (O_813,N_4651,N_4672);
or UO_814 (O_814,N_4731,N_4708);
nand UO_815 (O_815,N_4935,N_4780);
and UO_816 (O_816,N_4521,N_4747);
nand UO_817 (O_817,N_4572,N_4993);
nor UO_818 (O_818,N_4773,N_4991);
or UO_819 (O_819,N_4604,N_4764);
xor UO_820 (O_820,N_4613,N_4874);
nor UO_821 (O_821,N_4640,N_4595);
or UO_822 (O_822,N_4621,N_4850);
and UO_823 (O_823,N_4755,N_4614);
nand UO_824 (O_824,N_4815,N_4642);
or UO_825 (O_825,N_4780,N_4585);
xnor UO_826 (O_826,N_4862,N_4742);
and UO_827 (O_827,N_4774,N_4587);
nor UO_828 (O_828,N_4995,N_4822);
or UO_829 (O_829,N_4737,N_4830);
nand UO_830 (O_830,N_4681,N_4983);
or UO_831 (O_831,N_4649,N_4608);
and UO_832 (O_832,N_4853,N_4541);
nand UO_833 (O_833,N_4926,N_4861);
nand UO_834 (O_834,N_4955,N_4943);
xor UO_835 (O_835,N_4859,N_4958);
nand UO_836 (O_836,N_4821,N_4559);
xnor UO_837 (O_837,N_4520,N_4827);
nor UO_838 (O_838,N_4648,N_4788);
nand UO_839 (O_839,N_4514,N_4941);
xor UO_840 (O_840,N_4623,N_4924);
nor UO_841 (O_841,N_4793,N_4940);
or UO_842 (O_842,N_4923,N_4972);
and UO_843 (O_843,N_4882,N_4851);
xor UO_844 (O_844,N_4640,N_4986);
nand UO_845 (O_845,N_4521,N_4820);
nor UO_846 (O_846,N_4780,N_4515);
xnor UO_847 (O_847,N_4896,N_4908);
nand UO_848 (O_848,N_4638,N_4723);
nor UO_849 (O_849,N_4605,N_4554);
xor UO_850 (O_850,N_4726,N_4756);
and UO_851 (O_851,N_4998,N_4808);
xnor UO_852 (O_852,N_4825,N_4541);
and UO_853 (O_853,N_4855,N_4727);
or UO_854 (O_854,N_4799,N_4517);
xor UO_855 (O_855,N_4715,N_4630);
nand UO_856 (O_856,N_4532,N_4520);
nor UO_857 (O_857,N_4880,N_4580);
nand UO_858 (O_858,N_4938,N_4648);
xnor UO_859 (O_859,N_4605,N_4760);
nor UO_860 (O_860,N_4628,N_4835);
or UO_861 (O_861,N_4838,N_4563);
nor UO_862 (O_862,N_4527,N_4944);
and UO_863 (O_863,N_4665,N_4958);
and UO_864 (O_864,N_4561,N_4595);
and UO_865 (O_865,N_4887,N_4956);
nor UO_866 (O_866,N_4971,N_4852);
nor UO_867 (O_867,N_4573,N_4542);
nand UO_868 (O_868,N_4879,N_4724);
nand UO_869 (O_869,N_4763,N_4672);
nand UO_870 (O_870,N_4566,N_4609);
and UO_871 (O_871,N_4814,N_4555);
nor UO_872 (O_872,N_4818,N_4814);
xnor UO_873 (O_873,N_4525,N_4703);
xnor UO_874 (O_874,N_4791,N_4569);
nand UO_875 (O_875,N_4682,N_4549);
and UO_876 (O_876,N_4504,N_4921);
xnor UO_877 (O_877,N_4795,N_4861);
or UO_878 (O_878,N_4511,N_4778);
nor UO_879 (O_879,N_4915,N_4840);
nor UO_880 (O_880,N_4549,N_4971);
nor UO_881 (O_881,N_4770,N_4742);
and UO_882 (O_882,N_4636,N_4690);
nor UO_883 (O_883,N_4899,N_4550);
nand UO_884 (O_884,N_4532,N_4945);
or UO_885 (O_885,N_4523,N_4718);
nor UO_886 (O_886,N_4674,N_4576);
or UO_887 (O_887,N_4664,N_4505);
nand UO_888 (O_888,N_4957,N_4511);
and UO_889 (O_889,N_4697,N_4580);
nor UO_890 (O_890,N_4866,N_4557);
xor UO_891 (O_891,N_4882,N_4931);
xor UO_892 (O_892,N_4754,N_4718);
xor UO_893 (O_893,N_4756,N_4949);
xor UO_894 (O_894,N_4615,N_4963);
and UO_895 (O_895,N_4819,N_4629);
xor UO_896 (O_896,N_4649,N_4500);
and UO_897 (O_897,N_4800,N_4808);
nor UO_898 (O_898,N_4837,N_4856);
nand UO_899 (O_899,N_4989,N_4553);
or UO_900 (O_900,N_4637,N_4832);
xnor UO_901 (O_901,N_4966,N_4837);
xor UO_902 (O_902,N_4833,N_4653);
nor UO_903 (O_903,N_4557,N_4782);
nand UO_904 (O_904,N_4839,N_4693);
xnor UO_905 (O_905,N_4762,N_4896);
xor UO_906 (O_906,N_4528,N_4860);
and UO_907 (O_907,N_4564,N_4532);
or UO_908 (O_908,N_4694,N_4944);
or UO_909 (O_909,N_4768,N_4504);
nor UO_910 (O_910,N_4674,N_4710);
xor UO_911 (O_911,N_4807,N_4721);
or UO_912 (O_912,N_4613,N_4912);
nor UO_913 (O_913,N_4979,N_4921);
nor UO_914 (O_914,N_4697,N_4671);
xor UO_915 (O_915,N_4709,N_4665);
and UO_916 (O_916,N_4519,N_4561);
nand UO_917 (O_917,N_4921,N_4745);
nor UO_918 (O_918,N_4648,N_4850);
or UO_919 (O_919,N_4796,N_4963);
xnor UO_920 (O_920,N_4745,N_4779);
nand UO_921 (O_921,N_4781,N_4929);
and UO_922 (O_922,N_4722,N_4595);
nand UO_923 (O_923,N_4809,N_4555);
nor UO_924 (O_924,N_4589,N_4817);
and UO_925 (O_925,N_4674,N_4884);
xor UO_926 (O_926,N_4825,N_4971);
and UO_927 (O_927,N_4833,N_4590);
xnor UO_928 (O_928,N_4906,N_4820);
nor UO_929 (O_929,N_4505,N_4823);
nand UO_930 (O_930,N_4700,N_4724);
nor UO_931 (O_931,N_4751,N_4599);
nand UO_932 (O_932,N_4736,N_4708);
and UO_933 (O_933,N_4928,N_4541);
and UO_934 (O_934,N_4513,N_4693);
and UO_935 (O_935,N_4873,N_4798);
or UO_936 (O_936,N_4652,N_4725);
nor UO_937 (O_937,N_4715,N_4862);
nor UO_938 (O_938,N_4555,N_4739);
xor UO_939 (O_939,N_4801,N_4568);
and UO_940 (O_940,N_4564,N_4649);
nand UO_941 (O_941,N_4987,N_4561);
xor UO_942 (O_942,N_4895,N_4852);
xnor UO_943 (O_943,N_4977,N_4933);
or UO_944 (O_944,N_4574,N_4530);
xor UO_945 (O_945,N_4936,N_4668);
nor UO_946 (O_946,N_4803,N_4830);
xnor UO_947 (O_947,N_4732,N_4619);
or UO_948 (O_948,N_4958,N_4715);
nand UO_949 (O_949,N_4505,N_4708);
xor UO_950 (O_950,N_4616,N_4809);
and UO_951 (O_951,N_4518,N_4975);
and UO_952 (O_952,N_4546,N_4972);
xor UO_953 (O_953,N_4802,N_4711);
and UO_954 (O_954,N_4992,N_4810);
or UO_955 (O_955,N_4929,N_4556);
nor UO_956 (O_956,N_4899,N_4511);
and UO_957 (O_957,N_4820,N_4860);
and UO_958 (O_958,N_4584,N_4526);
nor UO_959 (O_959,N_4654,N_4630);
xor UO_960 (O_960,N_4650,N_4529);
nand UO_961 (O_961,N_4748,N_4508);
xor UO_962 (O_962,N_4536,N_4822);
and UO_963 (O_963,N_4902,N_4814);
nor UO_964 (O_964,N_4963,N_4679);
nand UO_965 (O_965,N_4971,N_4731);
nand UO_966 (O_966,N_4644,N_4558);
nand UO_967 (O_967,N_4530,N_4587);
and UO_968 (O_968,N_4732,N_4909);
xnor UO_969 (O_969,N_4950,N_4875);
nand UO_970 (O_970,N_4915,N_4830);
xor UO_971 (O_971,N_4898,N_4731);
or UO_972 (O_972,N_4546,N_4577);
nor UO_973 (O_973,N_4550,N_4521);
and UO_974 (O_974,N_4859,N_4526);
nand UO_975 (O_975,N_4845,N_4560);
or UO_976 (O_976,N_4564,N_4652);
and UO_977 (O_977,N_4605,N_4730);
xor UO_978 (O_978,N_4805,N_4822);
or UO_979 (O_979,N_4564,N_4579);
nand UO_980 (O_980,N_4692,N_4793);
or UO_981 (O_981,N_4731,N_4900);
nor UO_982 (O_982,N_4985,N_4532);
nand UO_983 (O_983,N_4860,N_4564);
nand UO_984 (O_984,N_4837,N_4568);
nand UO_985 (O_985,N_4761,N_4737);
nand UO_986 (O_986,N_4901,N_4896);
nand UO_987 (O_987,N_4730,N_4735);
nand UO_988 (O_988,N_4688,N_4587);
and UO_989 (O_989,N_4553,N_4672);
or UO_990 (O_990,N_4897,N_4517);
nand UO_991 (O_991,N_4837,N_4948);
and UO_992 (O_992,N_4988,N_4747);
nand UO_993 (O_993,N_4990,N_4595);
and UO_994 (O_994,N_4941,N_4790);
and UO_995 (O_995,N_4813,N_4690);
xor UO_996 (O_996,N_4919,N_4693);
and UO_997 (O_997,N_4525,N_4989);
xnor UO_998 (O_998,N_4997,N_4917);
xor UO_999 (O_999,N_4811,N_4667);
endmodule