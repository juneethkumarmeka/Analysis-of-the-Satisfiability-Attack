module basic_1500_15000_2000_75_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_963,In_214);
and U1 (N_1,In_411,In_841);
nor U2 (N_2,In_84,In_1474);
xnor U3 (N_3,In_594,In_1355);
or U4 (N_4,In_800,In_29);
nand U5 (N_5,In_508,In_123);
nor U6 (N_6,In_336,In_636);
xnor U7 (N_7,In_1231,In_957);
xnor U8 (N_8,In_568,In_949);
nand U9 (N_9,In_779,In_937);
xor U10 (N_10,In_490,In_794);
nand U11 (N_11,In_1398,In_433);
and U12 (N_12,In_566,In_142);
or U13 (N_13,In_1167,In_589);
or U14 (N_14,In_1186,In_1115);
nor U15 (N_15,In_1470,In_138);
nor U16 (N_16,In_671,In_980);
or U17 (N_17,In_833,In_204);
and U18 (N_18,In_1255,In_1314);
nand U19 (N_19,In_1184,In_638);
nor U20 (N_20,In_557,In_639);
and U21 (N_21,In_1235,In_1183);
nand U22 (N_22,In_510,In_58);
or U23 (N_23,In_896,In_1360);
nor U24 (N_24,In_1440,In_1327);
and U25 (N_25,In_1047,In_1017);
nand U26 (N_26,In_1143,In_1204);
nand U27 (N_27,In_19,In_978);
xnor U28 (N_28,In_341,In_273);
or U29 (N_29,In_179,In_778);
xnor U30 (N_30,In_30,In_1237);
nand U31 (N_31,In_926,In_590);
nor U32 (N_32,In_1495,In_954);
or U33 (N_33,In_288,In_934);
or U34 (N_34,In_1034,In_651);
or U35 (N_35,In_665,In_378);
and U36 (N_36,In_400,In_1029);
xnor U37 (N_37,In_1304,In_921);
nand U38 (N_38,In_1272,In_1373);
nor U39 (N_39,In_164,In_753);
xnor U40 (N_40,In_1059,In_1309);
and U41 (N_41,In_34,In_967);
nor U42 (N_42,In_907,In_468);
xnor U43 (N_43,In_867,In_674);
xor U44 (N_44,In_1410,In_1072);
xor U45 (N_45,In_988,In_587);
xor U46 (N_46,In_1019,In_816);
or U47 (N_47,In_818,In_687);
xnor U48 (N_48,In_600,In_185);
and U49 (N_49,In_1101,In_976);
xnor U50 (N_50,In_1040,In_947);
nand U51 (N_51,In_1145,In_26);
nand U52 (N_52,In_1273,In_231);
or U53 (N_53,In_211,In_145);
xor U54 (N_54,In_1426,In_666);
and U55 (N_55,In_1238,In_785);
nor U56 (N_56,In_902,In_1176);
or U57 (N_57,In_243,In_802);
nand U58 (N_58,In_31,In_1246);
nand U59 (N_59,In_1009,In_565);
nand U60 (N_60,In_1413,In_783);
or U61 (N_61,In_956,In_768);
nand U62 (N_62,In_1378,In_745);
nand U63 (N_63,In_1486,In_1050);
or U64 (N_64,In_1032,In_321);
nand U65 (N_65,In_1036,In_1357);
nor U66 (N_66,In_175,In_1061);
nand U67 (N_67,In_1066,In_884);
xnor U68 (N_68,In_523,In_1347);
nor U69 (N_69,In_39,In_1431);
xor U70 (N_70,In_215,In_462);
nor U71 (N_71,In_40,In_407);
and U72 (N_72,In_168,In_1464);
or U73 (N_73,In_326,In_972);
or U74 (N_74,In_631,In_943);
or U75 (N_75,In_1039,In_1139);
xnor U76 (N_76,In_1142,In_1001);
or U77 (N_77,In_1316,In_358);
nor U78 (N_78,In_1102,In_419);
nor U79 (N_79,In_292,In_13);
xnor U80 (N_80,In_1094,In_556);
nand U81 (N_81,In_707,In_573);
or U82 (N_82,In_1498,In_235);
nand U83 (N_83,In_1092,In_78);
xnor U84 (N_84,In_901,In_71);
nor U85 (N_85,In_24,In_338);
nand U86 (N_86,In_852,In_1057);
and U87 (N_87,In_424,In_904);
xor U88 (N_88,In_1415,In_37);
nand U89 (N_89,In_45,In_881);
and U90 (N_90,In_552,In_363);
or U91 (N_91,In_1239,In_222);
nor U92 (N_92,In_483,In_1322);
or U93 (N_93,In_877,In_251);
and U94 (N_94,In_649,In_1229);
xor U95 (N_95,In_888,In_1450);
xnor U96 (N_96,In_1342,In_413);
nor U97 (N_97,In_193,In_1086);
or U98 (N_98,In_323,In_160);
xor U99 (N_99,In_828,In_208);
and U100 (N_100,In_613,In_1010);
nand U101 (N_101,In_197,In_1163);
and U102 (N_102,In_938,In_1307);
nor U103 (N_103,In_788,In_428);
nand U104 (N_104,In_445,In_1149);
nand U105 (N_105,In_1445,In_452);
nor U106 (N_106,In_6,In_619);
and U107 (N_107,In_1269,In_796);
or U108 (N_108,In_767,In_1211);
xnor U109 (N_109,In_908,In_758);
nand U110 (N_110,In_153,In_1244);
or U111 (N_111,In_1058,In_520);
and U112 (N_112,In_584,In_539);
xnor U113 (N_113,In_822,In_1110);
nor U114 (N_114,In_264,In_353);
and U115 (N_115,In_699,In_1003);
or U116 (N_116,In_1132,In_128);
or U117 (N_117,In_798,In_1114);
nand U118 (N_118,In_977,In_431);
and U119 (N_119,In_1449,In_731);
and U120 (N_120,In_1350,In_472);
or U121 (N_121,In_1321,In_1306);
and U122 (N_122,In_668,In_340);
xnor U123 (N_123,In_1218,In_79);
nor U124 (N_124,In_1120,In_293);
and U125 (N_125,In_1388,In_184);
and U126 (N_126,In_1397,In_70);
nor U127 (N_127,In_366,In_985);
or U128 (N_128,In_564,In_839);
or U129 (N_129,In_232,In_1024);
xnor U130 (N_130,In_1479,In_190);
or U131 (N_131,In_696,In_726);
or U132 (N_132,In_124,In_1080);
and U133 (N_133,In_152,In_405);
and U134 (N_134,In_494,In_5);
nand U135 (N_135,In_1077,In_922);
xnor U136 (N_136,In_530,In_1095);
xnor U137 (N_137,In_749,In_515);
or U138 (N_138,In_1436,In_862);
nor U139 (N_139,In_359,In_1326);
or U140 (N_140,In_398,In_391);
and U141 (N_141,In_1333,In_1344);
nor U142 (N_142,In_1267,In_1315);
nor U143 (N_143,In_1345,In_484);
xor U144 (N_144,In_681,In_174);
xor U145 (N_145,In_233,In_657);
and U146 (N_146,In_65,In_834);
xor U147 (N_147,In_1369,In_648);
xnor U148 (N_148,In_771,In_1295);
xor U149 (N_149,In_893,In_1113);
nand U150 (N_150,In_488,In_1282);
or U151 (N_151,In_534,In_1311);
nand U152 (N_152,In_698,In_919);
xnor U153 (N_153,In_1462,In_952);
nand U154 (N_154,In_74,In_1499);
or U155 (N_155,In_471,In_558);
nor U156 (N_156,In_955,In_1035);
nand U157 (N_157,In_249,In_1310);
nor U158 (N_158,In_969,In_968);
or U159 (N_159,In_772,In_429);
nand U160 (N_160,In_192,In_981);
xnor U161 (N_161,In_50,In_927);
and U162 (N_162,In_924,In_560);
xor U163 (N_163,In_1420,In_1290);
nor U164 (N_164,In_1334,In_202);
and U165 (N_165,In_171,In_1041);
nor U166 (N_166,In_1067,In_569);
nand U167 (N_167,In_1053,In_1361);
or U168 (N_168,In_1411,In_150);
and U169 (N_169,In_332,In_650);
and U170 (N_170,In_1002,In_143);
nor U171 (N_171,In_57,In_299);
nand U172 (N_172,In_607,In_252);
and U173 (N_173,In_1241,In_1414);
xnor U174 (N_174,In_456,In_825);
nand U175 (N_175,In_858,In_505);
and U176 (N_176,In_608,In_982);
nand U177 (N_177,In_38,In_1289);
xor U178 (N_178,In_1140,In_69);
and U179 (N_179,In_1324,In_1243);
nor U180 (N_180,In_664,In_795);
or U181 (N_181,In_319,In_513);
or U182 (N_182,In_1129,In_860);
xnor U183 (N_183,In_882,In_477);
nor U184 (N_184,In_387,In_1480);
nand U185 (N_185,In_1359,In_330);
and U186 (N_186,In_1060,In_502);
nand U187 (N_187,In_418,In_527);
nor U188 (N_188,In_770,In_482);
nor U189 (N_189,In_1141,In_9);
and U190 (N_190,In_894,In_261);
nor U191 (N_191,In_1427,In_1338);
nand U192 (N_192,In_129,In_914);
and U193 (N_193,In_618,In_1070);
or U194 (N_194,In_722,In_998);
nor U195 (N_195,In_507,In_1368);
and U196 (N_196,In_371,In_541);
nor U197 (N_197,In_642,In_318);
nor U198 (N_198,In_1494,In_1225);
nor U199 (N_199,In_1298,In_1021);
and U200 (N_200,In_63,N_153);
nand U201 (N_201,In_1429,In_492);
nor U202 (N_202,In_42,In_61);
and U203 (N_203,In_144,In_876);
nor U204 (N_204,In_1007,In_617);
nor U205 (N_205,In_658,In_1351);
nor U206 (N_206,In_803,In_535);
nand U207 (N_207,In_1276,N_159);
or U208 (N_208,In_633,In_1286);
or U209 (N_209,In_975,N_84);
nand U210 (N_210,In_172,N_147);
xnor U211 (N_211,In_368,In_889);
and U212 (N_212,N_34,In_1406);
nand U213 (N_213,In_903,In_1160);
and U214 (N_214,In_609,In_1089);
nand U215 (N_215,In_11,N_133);
or U216 (N_216,N_50,N_154);
nor U217 (N_217,In_109,In_322);
nand U218 (N_218,In_241,In_349);
xnor U219 (N_219,In_1493,In_1127);
xnor U220 (N_220,In_156,In_550);
or U221 (N_221,N_195,In_1245);
and U222 (N_222,In_700,In_1016);
nor U223 (N_223,In_266,In_146);
nand U224 (N_224,In_414,In_1485);
nand U225 (N_225,In_620,In_161);
nand U226 (N_226,In_103,In_1384);
or U227 (N_227,In_995,In_685);
nand U228 (N_228,In_166,In_364);
or U229 (N_229,In_1015,In_1006);
or U230 (N_230,In_849,N_8);
and U231 (N_231,In_1191,In_426);
or U232 (N_232,In_1097,In_842);
or U233 (N_233,In_1028,In_1228);
or U234 (N_234,N_48,In_522);
and U235 (N_235,In_821,In_1412);
xor U236 (N_236,In_1472,N_179);
and U237 (N_237,In_1386,In_1352);
or U238 (N_238,N_26,In_640);
nand U239 (N_239,In_1469,N_190);
or U240 (N_240,In_1135,In_46);
nand U241 (N_241,In_928,In_85);
xor U242 (N_242,In_1296,In_1328);
nand U243 (N_243,In_177,N_127);
and U244 (N_244,In_1161,In_278);
or U245 (N_245,In_401,In_1134);
xnor U246 (N_246,In_335,In_1288);
and U247 (N_247,In_693,In_1155);
nand U248 (N_248,In_131,N_102);
nand U249 (N_249,In_396,In_540);
or U250 (N_250,In_317,In_899);
nand U251 (N_251,In_17,In_1096);
and U252 (N_252,In_496,In_1483);
or U253 (N_253,In_602,In_945);
or U254 (N_254,In_994,In_809);
and U255 (N_255,N_30,In_760);
xnor U256 (N_256,In_100,In_582);
xnor U257 (N_257,In_290,N_72);
xnor U258 (N_258,In_845,In_104);
and U259 (N_259,In_1153,N_15);
and U260 (N_260,In_1170,In_1085);
nand U261 (N_261,In_936,In_258);
xnor U262 (N_262,In_271,N_188);
xnor U263 (N_263,N_31,In_571);
and U264 (N_264,In_1062,In_280);
and U265 (N_265,In_101,In_559);
xor U266 (N_266,In_1337,N_9);
or U267 (N_267,In_1091,In_1078);
nor U268 (N_268,In_561,In_422);
nand U269 (N_269,In_814,In_485);
and U270 (N_270,In_580,In_12);
nor U271 (N_271,N_199,In_352);
nand U272 (N_272,In_596,In_425);
nor U273 (N_273,N_14,N_107);
or U274 (N_274,In_734,In_495);
and U275 (N_275,N_135,In_1093);
xnor U276 (N_276,In_244,In_865);
or U277 (N_277,In_708,In_676);
or U278 (N_278,In_281,In_73);
xor U279 (N_279,In_738,In_1329);
and U280 (N_280,In_538,In_159);
nor U281 (N_281,In_227,In_764);
nor U282 (N_282,In_355,N_89);
nand U283 (N_283,In_312,In_686);
xor U284 (N_284,In_1022,In_1442);
xor U285 (N_285,In_1068,In_1150);
nor U286 (N_286,In_1433,In_1240);
nand U287 (N_287,N_18,In_1362);
nor U288 (N_288,In_1000,In_1477);
and U289 (N_289,In_993,In_545);
and U290 (N_290,In_824,In_1206);
nor U291 (N_291,In_1409,In_1222);
nand U292 (N_292,In_250,In_1216);
nor U293 (N_293,N_7,N_83);
and U294 (N_294,N_22,In_248);
nand U295 (N_295,In_1421,In_1205);
and U296 (N_296,In_132,In_7);
nand U297 (N_297,In_1199,In_122);
or U298 (N_298,In_586,N_21);
nor U299 (N_299,N_38,In_1490);
xor U300 (N_300,In_44,In_134);
nor U301 (N_301,In_757,In_1223);
or U302 (N_302,In_660,In_811);
xnor U303 (N_303,In_886,In_830);
xnor U304 (N_304,In_1179,In_1444);
or U305 (N_305,In_663,In_504);
xor U306 (N_306,N_35,N_181);
xor U307 (N_307,In_1382,In_498);
xnor U308 (N_308,N_139,In_1465);
and U309 (N_309,N_162,In_684);
or U310 (N_310,In_107,In_479);
xor U311 (N_311,In_1076,In_1247);
and U312 (N_312,In_544,In_991);
nand U313 (N_313,In_89,In_909);
or U314 (N_314,In_518,In_188);
or U315 (N_315,In_268,N_97);
and U316 (N_316,In_791,N_177);
or U317 (N_317,In_1291,In_467);
nor U318 (N_318,In_774,In_399);
or U319 (N_319,N_47,In_56);
and U320 (N_320,In_1012,In_380);
nand U321 (N_321,In_88,In_1377);
nand U322 (N_322,In_1020,In_1340);
or U323 (N_323,In_1082,In_1370);
nand U324 (N_324,N_100,In_20);
and U325 (N_325,In_18,In_334);
and U326 (N_326,In_461,In_115);
or U327 (N_327,In_1399,In_509);
nand U328 (N_328,In_1128,In_690);
or U329 (N_329,In_1187,N_191);
nand U330 (N_330,In_1111,In_86);
nor U331 (N_331,N_178,N_96);
nor U332 (N_332,In_324,In_158);
or U333 (N_333,In_555,In_548);
xor U334 (N_334,In_388,In_1270);
nand U335 (N_335,In_1083,In_735);
nor U336 (N_336,In_1122,In_1004);
or U337 (N_337,In_715,N_82);
nor U338 (N_338,In_76,In_66);
nor U339 (N_339,In_984,In_1230);
nand U340 (N_340,N_11,N_28);
or U341 (N_341,In_1044,In_781);
nand U342 (N_342,In_592,In_27);
nand U343 (N_343,In_603,In_1422);
or U344 (N_344,In_1073,In_283);
nor U345 (N_345,In_3,In_1242);
nor U346 (N_346,In_593,N_131);
nor U347 (N_347,In_256,In_1379);
nor U348 (N_348,In_294,In_1496);
nor U349 (N_349,In_379,N_71);
and U350 (N_350,In_793,In_1025);
nor U351 (N_351,In_1468,In_627);
nor U352 (N_352,In_848,In_1166);
nand U353 (N_353,In_105,In_375);
and U354 (N_354,In_1088,N_86);
nand U355 (N_355,In_688,In_176);
xor U356 (N_356,In_744,In_1013);
or U357 (N_357,In_1437,In_652);
xor U358 (N_358,In_597,In_1424);
or U359 (N_359,N_92,In_1210);
and U360 (N_360,In_282,In_986);
xor U361 (N_361,In_528,In_119);
xor U362 (N_362,N_91,In_1461);
nor U363 (N_363,In_577,In_567);
xnor U364 (N_364,In_1318,In_1374);
xor U365 (N_365,In_189,In_667);
xnor U366 (N_366,In_784,N_165);
nand U367 (N_367,N_41,In_412);
nand U368 (N_368,N_143,In_727);
nor U369 (N_369,In_910,In_1348);
nor U370 (N_370,In_221,In_112);
xor U371 (N_371,In_55,In_32);
nand U372 (N_372,In_1123,N_62);
or U373 (N_373,In_1201,In_90);
and U374 (N_374,In_581,In_1185);
nand U375 (N_375,In_216,In_598);
xor U376 (N_376,In_328,In_1391);
xor U377 (N_377,In_1109,N_180);
nand U378 (N_378,N_16,In_389);
nor U379 (N_379,In_1265,In_905);
nand U380 (N_380,In_140,In_213);
nand U381 (N_381,In_98,In_1215);
nor U382 (N_382,In_553,In_1174);
nor U383 (N_383,In_1214,In_762);
or U384 (N_384,In_1489,In_951);
nor U385 (N_385,In_1038,In_813);
or U386 (N_386,In_1079,In_831);
and U387 (N_387,In_935,N_136);
and U388 (N_388,In_840,In_827);
or U389 (N_389,In_916,In_1071);
xor U390 (N_390,In_992,In_661);
xor U391 (N_391,N_76,In_1484);
xor U392 (N_392,In_572,In_1193);
and U393 (N_393,In_615,In_611);
nor U394 (N_394,N_29,In_1301);
or U395 (N_395,In_716,In_342);
and U396 (N_396,In_236,N_148);
or U397 (N_397,N_80,In_230);
xnor U398 (N_398,In_372,In_224);
xnor U399 (N_399,In_501,N_160);
nor U400 (N_400,N_258,In_1432);
or U401 (N_401,In_878,In_365);
and U402 (N_402,In_469,N_207);
or U403 (N_403,In_1278,In_33);
and U404 (N_404,In_247,In_220);
nor U405 (N_405,N_224,N_370);
nor U406 (N_406,In_1281,N_205);
nand U407 (N_407,In_999,N_156);
xor U408 (N_408,In_157,In_1297);
or U409 (N_409,N_229,In_1250);
and U410 (N_410,In_741,N_237);
nand U411 (N_411,In_370,N_349);
xnor U412 (N_412,In_614,In_1353);
and U413 (N_413,In_1308,In_180);
and U414 (N_414,In_1380,In_421);
nand U415 (N_415,In_303,N_276);
nor U416 (N_416,In_162,N_351);
and U417 (N_417,In_1446,N_275);
and U418 (N_418,In_1147,In_705);
or U419 (N_419,In_973,In_1098);
nor U420 (N_420,N_232,In_191);
or U421 (N_421,In_72,In_67);
xnor U422 (N_422,N_64,In_1260);
nand U423 (N_423,In_912,N_388);
or U424 (N_424,In_1320,In_377);
xnor U425 (N_425,In_234,In_737);
or U426 (N_426,N_74,In_476);
or U427 (N_427,In_276,In_864);
and U428 (N_428,In_679,N_397);
nor U429 (N_429,In_782,In_773);
xor U430 (N_430,N_140,In_92);
nor U431 (N_431,In_201,In_838);
nor U432 (N_432,In_1118,N_120);
and U433 (N_433,In_531,In_310);
xnor U434 (N_434,N_290,In_628);
xnor U435 (N_435,In_742,N_253);
or U436 (N_436,In_210,In_16);
xor U437 (N_437,In_465,In_1148);
nand U438 (N_438,In_151,In_307);
nor U439 (N_439,In_1136,In_381);
nand U440 (N_440,N_341,In_1457);
nor U441 (N_441,In_1419,N_304);
xnor U442 (N_442,N_347,In_1045);
or U443 (N_443,In_308,N_386);
xor U444 (N_444,In_920,In_850);
nor U445 (N_445,In_446,N_98);
nor U446 (N_446,N_296,In_163);
nor U447 (N_447,N_196,In_929);
or U448 (N_448,In_362,In_1117);
or U449 (N_449,N_282,N_151);
nor U450 (N_450,In_843,N_245);
nand U451 (N_451,In_897,In_797);
nor U452 (N_452,N_361,In_547);
nor U453 (N_453,In_662,In_237);
nand U454 (N_454,In_302,N_350);
nand U455 (N_455,N_13,In_83);
nand U456 (N_456,N_381,In_1116);
xnor U457 (N_457,In_526,In_1317);
nor U458 (N_458,In_678,In_1387);
and U459 (N_459,In_1219,In_1323);
nand U460 (N_460,In_1452,In_198);
or U461 (N_461,In_1430,In_759);
or U462 (N_462,In_750,In_304);
or U463 (N_463,In_1325,In_887);
nor U464 (N_464,N_330,In_720);
and U465 (N_465,In_635,N_222);
and U466 (N_466,In_944,In_855);
and U467 (N_467,In_106,In_60);
and U468 (N_468,N_19,In_223);
or U469 (N_469,In_1356,N_17);
nor U470 (N_470,In_270,In_1178);
and U471 (N_471,In_1104,In_1405);
or U472 (N_472,In_354,In_459);
nor U473 (N_473,N_369,In_141);
and U474 (N_474,In_709,N_88);
xnor U475 (N_475,In_801,In_697);
and U476 (N_476,In_287,In_1343);
nand U477 (N_477,In_444,In_601);
nand U478 (N_478,In_478,In_82);
and U479 (N_479,In_1042,In_41);
nor U480 (N_480,In_1453,In_416);
or U481 (N_481,In_403,In_656);
xor U482 (N_482,In_390,In_563);
nand U483 (N_483,In_634,In_130);
nor U484 (N_484,In_1133,N_288);
or U485 (N_485,In_205,N_344);
nor U486 (N_486,In_574,In_1182);
nand U487 (N_487,In_917,N_273);
and U488 (N_488,In_1151,N_79);
and U489 (N_489,In_780,In_930);
or U490 (N_490,In_729,In_1418);
or U491 (N_491,In_807,In_448);
xnor U492 (N_492,N_90,In_890);
and U493 (N_493,In_173,N_103);
xor U494 (N_494,In_81,In_554);
nor U495 (N_495,In_212,In_1366);
xor U496 (N_496,In_805,In_1279);
nand U497 (N_497,In_595,N_161);
and U498 (N_498,In_1138,In_606);
and U499 (N_499,In_1376,N_109);
xor U500 (N_500,In_203,In_80);
nand U501 (N_501,In_361,N_37);
xor U502 (N_502,In_272,N_278);
nor U503 (N_503,In_313,In_1175);
and U504 (N_504,In_420,In_895);
or U505 (N_505,N_392,In_942);
nor U506 (N_506,In_1169,N_371);
xnor U507 (N_507,In_931,In_1030);
nand U508 (N_508,In_125,N_54);
xor U509 (N_509,In_1299,In_22);
xor U510 (N_510,In_1385,N_145);
xnor U511 (N_511,In_136,In_1300);
xnor U512 (N_512,In_1434,N_146);
nor U513 (N_513,In_493,N_68);
nand U514 (N_514,N_117,In_423);
xor U515 (N_515,In_1305,N_24);
xor U516 (N_516,In_1152,N_215);
nand U517 (N_517,In_1354,N_149);
xor U518 (N_518,In_1371,In_542);
nor U519 (N_519,In_116,In_675);
nor U520 (N_520,In_121,In_837);
nor U521 (N_521,N_189,N_315);
and U522 (N_522,In_408,In_939);
xnor U523 (N_523,In_546,In_497);
or U524 (N_524,N_32,N_326);
xor U525 (N_525,N_39,N_94);
nand U526 (N_526,In_746,In_219);
and U527 (N_527,N_69,In_376);
or U528 (N_528,N_216,In_305);
nand U529 (N_529,In_733,In_75);
or U530 (N_530,N_214,N_353);
xor U531 (N_531,In_883,In_300);
and U532 (N_532,In_395,N_391);
xor U533 (N_533,In_1221,In_351);
nand U534 (N_534,In_551,N_265);
or U535 (N_535,In_94,In_616);
xor U536 (N_536,In_1403,In_99);
nor U537 (N_537,In_591,In_622);
xnor U538 (N_538,In_820,In_932);
or U539 (N_539,In_306,In_1158);
nor U540 (N_540,In_970,In_286);
xnor U541 (N_541,N_281,In_427);
nand U542 (N_542,N_5,In_692);
or U543 (N_543,In_1257,In_77);
and U544 (N_544,N_269,N_362);
nor U545 (N_545,In_836,In_432);
or U546 (N_546,In_1125,In_1266);
nand U547 (N_547,In_357,In_409);
and U548 (N_548,In_1196,N_223);
nand U549 (N_549,In_347,N_220);
or U550 (N_550,In_1456,In_792);
and U551 (N_551,N_342,In_1106);
nand U552 (N_552,In_776,In_1026);
and U553 (N_553,In_1330,In_799);
nor U554 (N_554,N_208,In_933);
nor U555 (N_555,In_1084,In_1226);
xor U556 (N_556,In_102,In_1112);
or U557 (N_557,N_56,N_385);
nor U558 (N_558,In_1294,In_866);
xnor U559 (N_559,N_40,N_95);
nand U560 (N_560,N_157,N_142);
or U561 (N_561,N_312,In_512);
nand U562 (N_562,N_198,In_437);
nand U563 (N_563,N_263,In_1497);
nor U564 (N_564,N_65,In_491);
and U565 (N_565,N_67,N_320);
nor U566 (N_566,In_327,In_262);
and U567 (N_567,In_217,In_940);
xor U568 (N_568,In_1224,In_384);
nor U569 (N_569,In_714,In_1404);
nand U570 (N_570,In_1396,N_58);
and U571 (N_571,N_193,In_440);
or U572 (N_572,In_575,In_417);
or U573 (N_573,N_176,In_1087);
or U574 (N_574,In_49,N_211);
nor U575 (N_575,N_168,N_396);
nor U576 (N_576,In_182,In_148);
and U577 (N_577,In_804,N_164);
nand U578 (N_578,In_669,N_70);
and U579 (N_579,In_576,N_118);
and U580 (N_580,In_458,In_165);
and U581 (N_581,In_277,In_1458);
nor U582 (N_582,N_365,In_702);
and U583 (N_583,In_386,In_962);
and U584 (N_584,In_732,N_319);
nand U585 (N_585,N_10,In_360);
nand U586 (N_586,N_247,N_318);
nand U587 (N_587,In_506,N_375);
nor U588 (N_588,In_769,In_51);
xor U589 (N_589,In_285,In_404);
nand U590 (N_590,In_1400,In_521);
xnor U591 (N_591,In_1189,In_1287);
nand U592 (N_592,In_625,N_20);
xor U593 (N_593,N_125,In_1293);
nand U594 (N_594,N_212,In_1236);
nand U595 (N_595,In_314,N_87);
xnor U596 (N_596,N_358,N_206);
and U597 (N_597,In_1389,N_383);
or U598 (N_598,In_1335,In_186);
xor U599 (N_599,N_284,In_1435);
xnor U600 (N_600,N_345,N_512);
and U601 (N_601,N_217,N_169);
xor U602 (N_602,In_691,N_407);
nor U603 (N_603,N_563,In_487);
xor U604 (N_604,In_1075,N_412);
nor U605 (N_605,In_654,N_372);
nor U606 (N_606,N_504,N_438);
or U607 (N_607,N_510,N_402);
xor U608 (N_608,In_885,In_87);
and U609 (N_609,N_430,N_550);
or U610 (N_610,In_1402,N_368);
nand U611 (N_611,In_178,N_52);
nand U612 (N_612,N_441,N_481);
nand U613 (N_613,In_1146,In_630);
nand U614 (N_614,In_135,In_689);
nor U615 (N_615,In_736,N_2);
xnor U616 (N_616,In_1209,N_526);
or U617 (N_617,In_95,In_238);
nand U618 (N_618,N_558,In_632);
nor U619 (N_619,N_1,N_431);
and U620 (N_620,In_1263,N_339);
nor U621 (N_621,N_150,In_925);
or U622 (N_622,N_443,N_213);
nor U623 (N_623,In_170,In_394);
nor U624 (N_624,N_366,N_202);
or U625 (N_625,In_62,N_252);
or U626 (N_626,In_875,In_1475);
and U627 (N_627,In_1171,In_1);
or U628 (N_628,In_1208,N_389);
nor U629 (N_629,N_45,N_201);
nor U630 (N_630,N_433,In_525);
and U631 (N_631,In_643,N_590);
or U632 (N_632,In_644,In_356);
and U633 (N_633,N_230,In_345);
nand U634 (N_634,In_1381,N_582);
and U635 (N_635,N_194,In_410);
xor U636 (N_636,In_284,N_360);
or U637 (N_637,In_460,In_1048);
xor U638 (N_638,In_54,N_226);
and U639 (N_639,In_48,In_1212);
xnor U640 (N_640,N_587,In_672);
nor U641 (N_641,In_68,In_680);
or U642 (N_642,In_25,N_447);
nor U643 (N_643,N_417,N_44);
or U644 (N_644,In_1248,N_473);
and U645 (N_645,N_409,N_537);
nor U646 (N_646,In_997,In_1473);
xor U647 (N_647,N_513,In_406);
or U648 (N_648,N_432,In_1005);
nand U649 (N_649,N_171,N_144);
nand U650 (N_650,In_155,In_295);
and U651 (N_651,In_1023,In_466);
xnor U652 (N_652,In_1491,In_1011);
or U653 (N_653,In_1439,In_870);
or U654 (N_654,In_879,In_1177);
nand U655 (N_655,In_447,N_124);
nand U656 (N_656,N_551,In_486);
nand U657 (N_657,N_297,N_301);
and U658 (N_658,In_473,In_1285);
xnor U659 (N_659,N_170,In_1275);
or U660 (N_660,N_557,N_123);
or U661 (N_661,In_187,N_401);
xnor U662 (N_662,N_503,In_1194);
or U663 (N_663,N_277,N_423);
and U664 (N_664,In_35,In_655);
xnor U665 (N_665,N_321,In_263);
or U666 (N_666,N_3,N_367);
nand U667 (N_667,N_477,N_444);
nand U668 (N_668,In_154,In_1234);
xor U669 (N_669,N_323,N_501);
or U670 (N_670,N_121,N_434);
and U671 (N_671,N_254,N_152);
and U672 (N_672,N_519,In_1331);
and U673 (N_673,N_336,In_971);
xnor U674 (N_674,N_373,In_1162);
xor U675 (N_675,In_200,N_554);
or U676 (N_676,N_453,N_584);
and U677 (N_677,N_502,N_586);
or U678 (N_678,In_817,N_289);
nand U679 (N_679,In_1292,N_489);
or U680 (N_680,In_516,In_960);
and U681 (N_681,N_246,N_219);
nand U682 (N_682,In_1251,N_442);
nand U683 (N_683,In_950,In_740);
nand U684 (N_684,In_296,N_418);
or U685 (N_685,In_1126,In_108);
and U686 (N_686,N_174,In_367);
nor U687 (N_687,In_829,In_1081);
xor U688 (N_688,N_540,N_115);
nand U689 (N_689,In_291,In_748);
nand U690 (N_690,In_537,N_119);
nand U691 (N_691,N_307,N_185);
and U692 (N_692,In_500,In_397);
and U693 (N_693,In_118,N_414);
and U694 (N_694,N_267,N_60);
xnor U695 (N_695,In_52,N_454);
nor U696 (N_696,N_244,In_1033);
nand U697 (N_697,N_73,In_585);
nor U698 (N_698,N_186,N_594);
nor U699 (N_699,N_475,In_646);
or U700 (N_700,N_259,In_1392);
nand U701 (N_701,In_1232,N_343);
xor U702 (N_702,N_49,In_1264);
or U703 (N_703,In_269,N_183);
nand U704 (N_704,N_428,In_254);
or U705 (N_705,In_815,In_712);
nor U706 (N_706,In_532,In_1466);
and U707 (N_707,In_570,In_91);
nand U708 (N_708,In_441,N_187);
or U709 (N_709,In_311,In_605);
nand U710 (N_710,In_350,N_416);
or U711 (N_711,N_484,In_987);
xnor U712 (N_712,In_941,N_308);
and U713 (N_713,N_225,In_1460);
and U714 (N_714,N_547,In_673);
or U715 (N_715,In_2,N_487);
xnor U716 (N_716,In_1202,N_163);
xor U717 (N_717,In_259,N_427);
nor U718 (N_718,In_455,In_946);
nor U719 (N_719,In_133,N_6);
nand U720 (N_720,In_1258,N_236);
xnor U721 (N_721,N_104,In_1220);
xnor U722 (N_722,In_743,In_1198);
nor U723 (N_723,N_411,N_262);
nor U724 (N_724,In_806,N_77);
xor U725 (N_725,In_1173,N_184);
nand U726 (N_726,N_53,In_724);
and U727 (N_727,N_458,In_514);
nor U728 (N_728,In_1008,In_181);
and U729 (N_729,In_1451,N_497);
xor U730 (N_730,In_1303,N_55);
or U731 (N_731,N_243,In_517);
nand U732 (N_732,In_511,In_149);
and U733 (N_733,N_479,In_892);
or U734 (N_734,N_210,In_647);
and U735 (N_735,In_297,In_990);
nand U736 (N_736,In_763,In_209);
and U737 (N_737,N_376,In_369);
nor U738 (N_738,In_789,N_508);
xor U739 (N_739,N_337,In_621);
nand U740 (N_740,In_337,N_257);
nand U741 (N_741,In_1100,N_280);
xor U742 (N_742,N_589,In_183);
nand U743 (N_743,N_166,In_682);
nor U744 (N_744,In_1423,N_405);
nand U745 (N_745,In_1154,In_900);
nor U746 (N_746,In_374,In_64);
nand U747 (N_747,In_1014,In_579);
nor U748 (N_748,In_1375,In_1164);
and U749 (N_749,N_382,In_489);
or U750 (N_750,In_953,N_231);
or U751 (N_751,In_610,In_1031);
nand U752 (N_752,N_597,In_728);
nor U753 (N_753,In_844,In_1407);
xor U754 (N_754,In_333,In_1197);
or U755 (N_755,In_346,N_379);
xnor U756 (N_756,In_1284,In_343);
nand U757 (N_757,N_556,N_555);
and U758 (N_758,N_514,N_455);
nand U759 (N_759,In_1274,In_1302);
xnor U760 (N_760,In_1336,In_823);
nor U761 (N_761,N_380,N_81);
and U762 (N_762,N_486,N_209);
or U763 (N_763,N_425,In_339);
and U764 (N_764,N_299,In_1358);
nor U765 (N_765,N_528,N_105);
or U766 (N_766,In_857,N_421);
xor U767 (N_767,N_534,In_257);
xnor U768 (N_768,N_240,N_363);
xor U769 (N_769,In_1408,N_25);
or U770 (N_770,In_859,N_398);
xnor U771 (N_771,In_624,N_460);
xnor U772 (N_772,N_271,N_578);
xor U773 (N_773,In_1447,In_1108);
nand U774 (N_774,In_137,In_948);
nor U775 (N_775,In_645,N_527);
xor U776 (N_776,In_240,In_301);
and U777 (N_777,In_385,In_659);
nand U778 (N_778,N_130,N_328);
nor U779 (N_779,N_137,In_1107);
and U780 (N_780,In_1121,N_285);
nand U781 (N_781,N_437,N_302);
nor U782 (N_782,N_567,N_250);
or U783 (N_783,In_721,In_199);
xnor U784 (N_784,In_1131,In_218);
nand U785 (N_785,In_701,N_509);
nor U786 (N_786,N_0,N_451);
and U787 (N_787,In_812,In_1049);
nand U788 (N_788,N_112,In_958);
nand U789 (N_789,In_1065,In_761);
nand U790 (N_790,In_847,N_354);
nand U791 (N_791,N_274,N_394);
nor U792 (N_792,In_206,N_413);
xor U793 (N_793,N_482,In_435);
and U794 (N_794,N_251,N_445);
or U795 (N_795,In_1393,In_1192);
xor U796 (N_796,In_147,In_1052);
xnor U797 (N_797,In_454,N_134);
nor U798 (N_798,In_113,N_234);
nand U799 (N_799,In_1063,N_291);
xnor U800 (N_800,N_436,In_373);
nand U801 (N_801,In_863,In_1195);
xnor U802 (N_802,In_790,N_735);
and U803 (N_803,In_499,N_356);
nor U804 (N_804,N_694,N_678);
nor U805 (N_805,In_756,N_690);
nand U806 (N_806,In_965,N_724);
nand U807 (N_807,N_785,N_525);
and U808 (N_808,In_1254,In_434);
xor U809 (N_809,In_23,In_1492);
or U810 (N_810,N_769,N_741);
and U811 (N_811,In_239,In_583);
nor U812 (N_812,In_1056,N_172);
nand U813 (N_813,In_331,In_207);
xor U814 (N_814,N_762,In_964);
nor U815 (N_815,In_436,N_562);
and U816 (N_816,In_543,N_794);
nand U817 (N_817,N_703,N_238);
or U818 (N_818,In_725,In_1103);
nand U819 (N_819,N_322,N_292);
or U820 (N_820,In_775,N_598);
xor U821 (N_821,N_496,N_42);
nand U822 (N_822,N_305,N_553);
nand U823 (N_823,In_1172,N_571);
nand U824 (N_824,N_197,N_75);
nor U825 (N_825,N_766,N_764);
and U826 (N_826,In_393,N_780);
nand U827 (N_827,In_225,N_729);
nand U828 (N_828,In_117,In_979);
or U829 (N_829,N_331,N_577);
and U830 (N_830,N_492,In_15);
or U831 (N_831,In_653,N_659);
nand U832 (N_832,N_352,In_1233);
nand U833 (N_833,N_774,In_536);
nor U834 (N_834,N_731,In_966);
nand U835 (N_835,In_1482,N_751);
nor U836 (N_836,N_335,N_485);
or U837 (N_837,N_701,In_1130);
xnor U838 (N_838,N_338,N_552);
and U839 (N_839,N_627,In_996);
and U840 (N_840,N_723,N_293);
nor U841 (N_841,N_623,N_357);
or U842 (N_842,N_204,N_521);
xor U843 (N_843,In_706,In_229);
and U844 (N_844,N_378,N_755);
and U845 (N_845,In_1200,In_253);
or U846 (N_846,In_1018,N_736);
nand U847 (N_847,N_666,In_59);
nand U848 (N_848,N_543,N_758);
nand U849 (N_849,N_122,N_93);
and U850 (N_850,N_662,In_1339);
and U851 (N_851,N_691,N_753);
xnor U852 (N_852,N_778,N_515);
nor U853 (N_853,N_472,N_283);
and U854 (N_854,In_915,In_1417);
or U855 (N_855,In_167,N_720);
or U856 (N_856,N_505,In_819);
xnor U857 (N_857,N_781,N_531);
or U858 (N_858,In_765,N_768);
or U859 (N_859,N_286,In_755);
nand U860 (N_860,In_430,In_1099);
and U861 (N_861,In_694,N_618);
nor U862 (N_862,In_961,N_333);
xnor U863 (N_863,N_446,In_1487);
or U864 (N_864,N_182,In_1159);
or U865 (N_865,N_192,In_641);
nand U866 (N_866,In_8,N_671);
nand U867 (N_867,In_747,In_97);
or U868 (N_868,In_880,In_529);
nor U869 (N_869,N_689,In_751);
or U870 (N_870,In_1256,N_51);
or U871 (N_871,In_1349,In_787);
nand U872 (N_872,N_287,N_680);
xor U873 (N_873,N_529,N_708);
xor U874 (N_874,N_777,In_1365);
or U875 (N_875,In_869,In_0);
nor U876 (N_876,N_393,In_1459);
xnor U877 (N_877,In_1372,N_128);
and U878 (N_878,In_918,N_249);
xnor U879 (N_879,N_466,N_233);
xnor U880 (N_880,In_1367,In_898);
or U881 (N_881,N_334,In_325);
nor U882 (N_882,In_383,In_1467);
xor U883 (N_883,In_713,N_786);
and U884 (N_884,In_871,N_488);
nor U885 (N_885,N_653,In_96);
or U886 (N_886,N_429,N_340);
nor U887 (N_887,In_1395,N_324);
nand U888 (N_888,In_1252,N_595);
and U889 (N_889,N_476,N_573);
nand U890 (N_890,N_517,In_1313);
and U891 (N_891,N_709,N_663);
and U892 (N_892,In_1064,N_541);
and U893 (N_893,In_1144,N_116);
xor U894 (N_894,N_520,In_683);
and U895 (N_895,In_1262,N_260);
or U896 (N_896,N_621,In_766);
nor U897 (N_897,N_400,In_279);
and U898 (N_898,In_194,N_648);
nand U899 (N_899,N_110,N_524);
nand U900 (N_900,In_1037,In_835);
xor U901 (N_901,N_631,In_1165);
nand U902 (N_902,N_298,N_173);
or U903 (N_903,N_687,N_507);
nor U904 (N_904,In_1213,In_1090);
nor U905 (N_905,N_467,N_727);
xnor U906 (N_906,In_195,In_47);
xnor U907 (N_907,N_439,In_730);
nand U908 (N_908,N_743,In_872);
or U909 (N_909,N_765,N_698);
nor U910 (N_910,N_620,In_1463);
nor U911 (N_911,N_12,In_53);
xor U912 (N_912,N_59,In_853);
xnor U913 (N_913,In_1259,N_732);
xnor U914 (N_914,N_111,N_108);
or U915 (N_915,N_532,In_309);
and U916 (N_916,N_797,In_873);
and U917 (N_917,In_854,N_384);
or U918 (N_918,N_27,In_1074);
nand U919 (N_919,N_264,N_779);
and U920 (N_920,N_471,N_348);
or U921 (N_921,N_685,N_715);
xnor U922 (N_922,N_643,N_646);
and U923 (N_923,N_574,In_260);
or U924 (N_924,In_246,N_759);
or U925 (N_925,In_275,N_622);
nor U926 (N_926,N_422,N_462);
xnor U927 (N_927,N_493,N_592);
or U928 (N_928,N_635,N_763);
and U929 (N_929,N_456,N_523);
and U930 (N_930,N_511,N_682);
or U931 (N_931,N_616,N_410);
nor U932 (N_932,N_660,In_245);
nand U933 (N_933,In_599,N_716);
xor U934 (N_934,N_266,N_329);
nand U935 (N_935,In_906,N_677);
nor U936 (N_936,N_775,N_658);
nor U937 (N_937,N_637,N_463);
nor U938 (N_938,In_392,In_1390);
nand U939 (N_939,In_1119,In_1055);
nor U940 (N_940,N_539,N_702);
xor U941 (N_941,N_311,In_1332);
nand U942 (N_942,N_608,In_1277);
nand U943 (N_943,In_450,N_218);
or U944 (N_944,N_248,In_832);
or U945 (N_945,In_1181,In_1346);
or U946 (N_946,N_576,In_923);
nand U947 (N_947,In_519,N_772);
nand U948 (N_948,In_1455,N_560);
xnor U949 (N_949,In_1253,N_310);
xnor U950 (N_950,N_656,In_289);
and U951 (N_951,N_387,N_795);
xnor U952 (N_952,N_722,In_453);
nand U953 (N_953,In_524,In_255);
nand U954 (N_954,In_316,N_718);
nand U955 (N_955,In_226,N_377);
nor U956 (N_956,N_506,In_114);
nand U957 (N_957,In_911,N_664);
xor U958 (N_958,N_609,N_516);
nor U959 (N_959,In_612,N_650);
or U960 (N_960,In_464,N_565);
and U961 (N_961,In_1137,N_469);
nand U962 (N_962,In_1188,N_667);
xor U963 (N_963,In_475,In_442);
xnor U964 (N_964,N_681,N_657);
nand U965 (N_965,N_737,In_1051);
and U966 (N_966,In_382,N_672);
and U967 (N_967,N_522,In_562);
nand U968 (N_968,N_33,N_239);
or U969 (N_969,In_1157,N_66);
nand U970 (N_970,N_221,In_242);
and U971 (N_971,N_776,In_629);
nor U972 (N_972,N_495,N_754);
nand U973 (N_973,In_457,N_533);
xnor U974 (N_974,In_1448,N_538);
or U975 (N_975,N_426,N_669);
nand U976 (N_976,N_713,In_1054);
nor U977 (N_977,In_1271,In_111);
xor U978 (N_978,N_752,In_1441);
or U979 (N_979,N_734,N_63);
or U980 (N_980,N_601,N_491);
or U981 (N_981,N_798,In_1341);
nand U982 (N_982,N_757,N_99);
or U983 (N_983,N_799,N_583);
xnor U984 (N_984,N_645,N_270);
nand U985 (N_985,N_611,In_126);
and U986 (N_986,In_503,N_796);
nand U987 (N_987,In_604,In_1190);
xnor U988 (N_988,N_23,N_642);
and U989 (N_989,In_1124,N_784);
and U990 (N_990,In_402,N_719);
nand U991 (N_991,N_603,In_704);
and U992 (N_992,N_36,N_314);
and U993 (N_993,N_268,In_549);
nand U994 (N_994,N_559,N_542);
xor U995 (N_995,N_744,N_544);
xor U996 (N_996,N_261,N_655);
or U997 (N_997,N_57,In_28);
nor U998 (N_998,In_1105,N_771);
nand U999 (N_999,N_256,N_85);
xnor U1000 (N_1000,N_699,In_265);
and U1001 (N_1001,N_242,In_480);
xnor U1002 (N_1002,N_61,N_928);
or U1003 (N_1003,In_1488,N_834);
nand U1004 (N_1004,In_1394,N_647);
or U1005 (N_1005,N_470,N_962);
nor U1006 (N_1006,N_468,N_963);
nor U1007 (N_1007,N_915,N_989);
and U1008 (N_1008,N_918,In_438);
nand U1009 (N_1009,N_880,N_948);
xnor U1010 (N_1010,N_725,N_887);
nand U1011 (N_1011,N_420,N_158);
xnor U1012 (N_1012,In_1481,N_728);
xnor U1013 (N_1013,N_739,N_810);
xnor U1014 (N_1014,In_1416,In_449);
xnor U1015 (N_1015,N_965,N_500);
nand U1016 (N_1016,N_332,N_303);
nor U1017 (N_1017,N_78,In_4);
and U1018 (N_1018,N_852,N_415);
nor U1019 (N_1019,In_1249,N_823);
or U1020 (N_1020,N_295,In_481);
xnor U1021 (N_1021,N_480,N_847);
nor U1022 (N_1022,N_809,N_203);
xnor U1023 (N_1023,N_970,N_981);
xnor U1024 (N_1024,N_824,N_612);
and U1025 (N_1025,N_748,N_856);
and U1026 (N_1026,N_850,N_985);
nor U1027 (N_1027,N_844,N_613);
and U1028 (N_1028,N_459,N_465);
nand U1029 (N_1029,In_1428,N_979);
and U1030 (N_1030,N_738,N_949);
xnor U1031 (N_1031,N_714,N_652);
xor U1032 (N_1032,N_947,N_43);
xor U1033 (N_1033,N_833,N_791);
and U1034 (N_1034,In_1156,N_939);
nand U1035 (N_1035,N_175,N_879);
or U1036 (N_1036,N_924,N_688);
xor U1037 (N_1037,N_575,N_749);
xor U1038 (N_1038,N_300,N_654);
or U1039 (N_1039,N_828,N_730);
nor U1040 (N_1040,N_990,N_901);
nor U1041 (N_1041,In_677,N_600);
xor U1042 (N_1042,N_869,N_639);
xor U1043 (N_1043,N_316,N_995);
nand U1044 (N_1044,In_695,In_1476);
xnor U1045 (N_1045,N_395,N_845);
nand U1046 (N_1046,N_294,N_836);
and U1047 (N_1047,N_853,In_974);
xor U1048 (N_1048,N_877,N_721);
nand U1049 (N_1049,N_882,N_899);
nand U1050 (N_1050,In_826,N_960);
or U1051 (N_1051,N_641,N_665);
or U1052 (N_1052,In_846,In_1180);
nor U1053 (N_1053,N_803,In_315);
nand U1054 (N_1054,N_902,N_863);
nor U1055 (N_1055,N_591,N_954);
or U1056 (N_1056,N_374,N_886);
and U1057 (N_1057,N_994,N_894);
nor U1058 (N_1058,In_1168,In_329);
or U1059 (N_1059,In_298,N_826);
xnor U1060 (N_1060,N_711,N_820);
xor U1061 (N_1061,N_46,N_905);
nand U1062 (N_1062,N_561,In_810);
xnor U1063 (N_1063,N_585,In_21);
and U1064 (N_1064,In_43,N_545);
xor U1065 (N_1065,N_760,In_169);
or U1066 (N_1066,N_792,N_490);
or U1067 (N_1067,In_1454,N_167);
nor U1068 (N_1068,N_726,N_839);
nor U1069 (N_1069,N_783,N_419);
or U1070 (N_1070,N_933,N_858);
xnor U1071 (N_1071,In_623,N_983);
nand U1072 (N_1072,N_364,In_710);
nor U1073 (N_1073,N_773,In_274);
nor U1074 (N_1074,N_483,N_132);
xnor U1075 (N_1075,N_789,N_309);
nor U1076 (N_1076,N_822,N_945);
xor U1077 (N_1077,In_1363,N_896);
nand U1078 (N_1078,N_756,N_346);
xnor U1079 (N_1079,In_717,N_815);
and U1080 (N_1080,N_919,N_988);
and U1081 (N_1081,N_838,N_888);
xor U1082 (N_1082,N_944,N_842);
nand U1083 (N_1083,N_602,N_306);
and U1084 (N_1084,In_891,N_549);
and U1085 (N_1085,N_325,N_615);
nor U1086 (N_1086,N_959,In_913);
and U1087 (N_1087,N_651,N_925);
nor U1088 (N_1088,N_546,N_964);
nor U1089 (N_1089,N_957,In_228);
and U1090 (N_1090,In_348,N_977);
or U1091 (N_1091,In_1227,N_837);
or U1092 (N_1092,In_1069,N_255);
nand U1093 (N_1093,N_911,N_998);
nand U1094 (N_1094,N_808,In_14);
nand U1095 (N_1095,In_120,In_439);
nand U1096 (N_1096,N_804,In_578);
or U1097 (N_1097,N_570,N_566);
xor U1098 (N_1098,N_126,N_746);
nand U1099 (N_1099,N_971,N_599);
and U1100 (N_1100,In_1471,N_868);
xor U1101 (N_1101,N_448,N_875);
or U1102 (N_1102,N_638,In_754);
or U1103 (N_1103,N_155,N_449);
xor U1104 (N_1104,N_862,In_1312);
nand U1105 (N_1105,N_390,N_790);
and U1106 (N_1106,N_920,N_581);
nand U1107 (N_1107,N_788,N_953);
nor U1108 (N_1108,N_700,In_110);
nand U1109 (N_1109,N_740,N_742);
nand U1110 (N_1110,In_344,N_625);
xnor U1111 (N_1111,N_892,In_1027);
nor U1112 (N_1112,In_533,In_723);
and U1113 (N_1113,N_840,N_881);
nand U1114 (N_1114,N_975,N_614);
nand U1115 (N_1115,N_707,N_767);
nor U1116 (N_1116,N_696,In_1217);
nand U1117 (N_1117,N_101,N_593);
nor U1118 (N_1118,N_903,In_588);
nand U1119 (N_1119,N_955,N_966);
or U1120 (N_1120,N_499,N_564);
nor U1121 (N_1121,N_424,In_752);
or U1122 (N_1122,N_898,N_846);
and U1123 (N_1123,N_978,N_951);
or U1124 (N_1124,In_415,In_1425);
or U1125 (N_1125,N_934,In_874);
or U1126 (N_1126,N_793,In_320);
and U1127 (N_1127,N_624,In_1207);
nor U1128 (N_1128,N_864,N_241);
and U1129 (N_1129,In_93,N_359);
or U1130 (N_1130,In_1203,N_404);
nor U1131 (N_1131,In_1478,N_676);
nor U1132 (N_1132,N_932,N_857);
nor U1133 (N_1133,In_739,N_440);
nor U1134 (N_1134,In_786,N_849);
and U1135 (N_1135,N_946,N_814);
nand U1136 (N_1136,N_113,N_200);
nand U1137 (N_1137,N_950,N_872);
nor U1138 (N_1138,N_569,N_138);
or U1139 (N_1139,N_452,In_139);
nand U1140 (N_1140,N_355,N_941);
nor U1141 (N_1141,In_868,In_463);
nand U1142 (N_1142,N_692,N_670);
nor U1143 (N_1143,N_907,N_818);
or U1144 (N_1144,In_1283,In_1268);
or U1145 (N_1145,N_106,N_938);
and U1146 (N_1146,N_874,N_835);
nand U1147 (N_1147,In_1043,N_461);
nand U1148 (N_1148,N_610,N_967);
nor U1149 (N_1149,In_1319,N_636);
or U1150 (N_1150,N_821,N_806);
or U1151 (N_1151,N_800,N_668);
nand U1152 (N_1152,N_891,N_782);
or U1153 (N_1153,In_36,N_969);
xnor U1154 (N_1154,N_634,N_579);
xnor U1155 (N_1155,In_719,N_916);
nand U1156 (N_1156,N_871,N_761);
nand U1157 (N_1157,In_703,N_403);
xor U1158 (N_1158,N_235,N_972);
nor U1159 (N_1159,N_604,N_958);
xor U1160 (N_1160,N_693,N_999);
nor U1161 (N_1161,N_626,N_399);
and U1162 (N_1162,N_536,N_878);
nand U1163 (N_1163,N_568,N_408);
nor U1164 (N_1164,N_866,In_196);
nor U1165 (N_1165,N_628,N_706);
nor U1166 (N_1166,N_710,N_952);
xnor U1167 (N_1167,In_1364,N_930);
nand U1168 (N_1168,N_801,N_535);
nand U1169 (N_1169,N_884,N_272);
nor U1170 (N_1170,N_588,N_596);
or U1171 (N_1171,N_457,N_675);
xnor U1172 (N_1172,N_984,N_917);
and U1173 (N_1173,N_770,N_910);
nand U1174 (N_1174,N_313,N_745);
xor U1175 (N_1175,N_883,N_997);
and U1176 (N_1176,In_983,N_841);
nor U1177 (N_1177,N_914,N_695);
nand U1178 (N_1178,N_870,In_1401);
xor U1179 (N_1179,N_900,In_989);
nand U1180 (N_1180,In_861,In_959);
or U1181 (N_1181,N_993,N_674);
nand U1182 (N_1182,In_127,N_619);
xor U1183 (N_1183,N_943,N_825);
nand U1184 (N_1184,N_805,In_443);
xor U1185 (N_1185,N_227,N_992);
and U1186 (N_1186,N_854,N_548);
nand U1187 (N_1187,N_478,N_435);
xnor U1188 (N_1188,N_860,In_718);
and U1189 (N_1189,N_661,N_733);
nor U1190 (N_1190,N_913,N_921);
and U1191 (N_1191,N_908,N_644);
and U1192 (N_1192,N_937,N_518);
nand U1193 (N_1193,N_996,In_470);
xnor U1194 (N_1194,In_1046,N_922);
or U1195 (N_1195,N_987,N_893);
xnor U1196 (N_1196,N_974,In_856);
nand U1197 (N_1197,N_673,N_889);
xor U1198 (N_1198,N_867,In_267);
and U1199 (N_1199,N_859,N_816);
nor U1200 (N_1200,N_1084,N_885);
xnor U1201 (N_1201,N_1132,N_1077);
nand U1202 (N_1202,N_807,N_679);
xnor U1203 (N_1203,N_890,N_1064);
xor U1204 (N_1204,N_530,N_1180);
xnor U1205 (N_1205,N_1004,N_1195);
xor U1206 (N_1206,N_1027,N_1140);
xor U1207 (N_1207,N_450,N_1094);
nand U1208 (N_1208,N_865,N_1146);
nor U1209 (N_1209,N_1069,N_1193);
or U1210 (N_1210,N_712,N_961);
and U1211 (N_1211,N_1163,N_629);
nor U1212 (N_1212,N_1013,N_923);
and U1213 (N_1213,N_1028,N_1192);
nand U1214 (N_1214,N_114,N_1179);
nand U1215 (N_1215,N_317,N_1014);
nor U1216 (N_1216,N_640,N_1174);
or U1217 (N_1217,N_1153,N_1187);
and U1218 (N_1218,N_697,In_626);
nand U1219 (N_1219,N_1092,N_1020);
xor U1220 (N_1220,N_1051,In_670);
and U1221 (N_1221,N_1111,N_1196);
and U1222 (N_1222,N_1058,N_1042);
nand U1223 (N_1223,In_451,N_474);
xor U1224 (N_1224,N_1168,In_1443);
xnor U1225 (N_1225,N_1190,N_1106);
nand U1226 (N_1226,N_1115,In_1280);
and U1227 (N_1227,N_1155,N_1026);
xnor U1228 (N_1228,N_1120,N_982);
or U1229 (N_1229,N_494,N_686);
and U1230 (N_1230,N_1088,N_1109);
or U1231 (N_1231,N_1105,N_1172);
and U1232 (N_1232,N_1113,N_1049);
nor U1233 (N_1233,N_1082,In_1261);
xor U1234 (N_1234,N_1183,N_1171);
and U1235 (N_1235,N_1127,In_711);
nor U1236 (N_1236,N_129,N_1039);
nand U1237 (N_1237,N_1100,N_228);
or U1238 (N_1238,N_1054,N_1009);
nand U1239 (N_1239,N_1018,N_1142);
and U1240 (N_1240,N_1099,N_1175);
nor U1241 (N_1241,N_811,N_1037);
and U1242 (N_1242,N_1083,N_1101);
nand U1243 (N_1243,N_787,N_986);
xor U1244 (N_1244,N_1011,N_1046);
and U1245 (N_1245,N_717,N_1110);
xor U1246 (N_1246,N_1118,N_1126);
xnor U1247 (N_1247,N_1145,N_1103);
or U1248 (N_1248,N_617,N_897);
or U1249 (N_1249,N_1061,N_1074);
nor U1250 (N_1250,N_750,N_1116);
nand U1251 (N_1251,N_605,N_968);
nor U1252 (N_1252,N_1107,N_1073);
nor U1253 (N_1253,N_1031,N_1038);
or U1254 (N_1254,N_1029,N_1005);
nand U1255 (N_1255,N_876,N_1068);
xnor U1256 (N_1256,N_1067,N_980);
xnor U1257 (N_1257,N_633,N_1102);
nand U1258 (N_1258,N_906,N_1041);
or U1259 (N_1259,N_1161,N_1090);
nor U1260 (N_1260,N_931,N_1040);
xor U1261 (N_1261,N_1149,In_1383);
or U1262 (N_1262,N_1000,N_1125);
nand U1263 (N_1263,N_1169,N_926);
nor U1264 (N_1264,N_1122,N_705);
nor U1265 (N_1265,N_935,N_1060);
nand U1266 (N_1266,N_832,N_1010);
nor U1267 (N_1267,N_843,N_630);
or U1268 (N_1268,N_1093,N_1108);
and U1269 (N_1269,N_1012,N_1136);
xnor U1270 (N_1270,N_572,N_1144);
nor U1271 (N_1271,N_1056,In_1438);
nor U1272 (N_1272,N_1159,N_1006);
or U1273 (N_1273,N_1089,N_827);
nand U1274 (N_1274,N_895,N_1057);
and U1275 (N_1275,N_976,N_1199);
xor U1276 (N_1276,In_851,N_1166);
or U1277 (N_1277,N_1071,N_747);
nand U1278 (N_1278,N_1164,N_848);
or U1279 (N_1279,N_1138,N_1112);
nand U1280 (N_1280,N_909,N_1019);
xor U1281 (N_1281,N_1165,N_1022);
xor U1282 (N_1282,N_1008,N_829);
xor U1283 (N_1283,N_1157,In_474);
nor U1284 (N_1284,N_1121,N_831);
nor U1285 (N_1285,N_812,N_1095);
xor U1286 (N_1286,N_1130,N_1160);
nand U1287 (N_1287,N_1197,N_1024);
or U1288 (N_1288,N_1189,N_498);
nor U1289 (N_1289,N_1177,N_1081);
xnor U1290 (N_1290,N_1025,N_819);
or U1291 (N_1291,N_1085,N_813);
xnor U1292 (N_1292,N_1035,N_1182);
xor U1293 (N_1293,N_873,N_1032);
nor U1294 (N_1294,N_1079,N_1052);
nor U1295 (N_1295,N_1181,N_1135);
nand U1296 (N_1296,N_991,N_1170);
nor U1297 (N_1297,N_1185,N_1087);
xor U1298 (N_1298,N_1198,N_1123);
nand U1299 (N_1299,N_1133,N_1045);
or U1300 (N_1300,N_1131,N_1129);
nor U1301 (N_1301,N_279,N_4);
xor U1302 (N_1302,N_1188,N_580);
xor U1303 (N_1303,N_1023,N_1176);
nand U1304 (N_1304,N_1044,N_1075);
and U1305 (N_1305,N_327,N_1086);
nand U1306 (N_1306,N_936,N_1065);
nand U1307 (N_1307,N_632,N_817);
nand U1308 (N_1308,N_1017,N_1173);
and U1309 (N_1309,N_1141,N_1194);
nor U1310 (N_1310,N_1021,N_956);
nor U1311 (N_1311,N_1097,N_1154);
nand U1312 (N_1312,N_1156,N_1147);
xnor U1313 (N_1313,N_1139,N_904);
or U1314 (N_1314,N_1062,N_1002);
or U1315 (N_1315,N_1191,N_649);
or U1316 (N_1316,N_942,In_808);
xnor U1317 (N_1317,N_406,N_1080);
nand U1318 (N_1318,N_1119,N_1137);
nand U1319 (N_1319,N_1063,N_1117);
nor U1320 (N_1320,N_927,N_1036);
nand U1321 (N_1321,N_1134,N_1076);
xnor U1322 (N_1322,N_861,N_855);
xor U1323 (N_1323,N_1151,N_704);
nand U1324 (N_1324,N_1184,N_1048);
and U1325 (N_1325,N_1124,N_1098);
nor U1326 (N_1326,N_929,N_973);
and U1327 (N_1327,N_1186,N_1178);
nand U1328 (N_1328,N_1043,N_851);
nand U1329 (N_1329,N_1162,N_1070);
and U1330 (N_1330,N_1015,N_141);
nand U1331 (N_1331,N_830,N_1053);
xor U1332 (N_1332,N_1050,N_1158);
xor U1333 (N_1333,N_1096,In_777);
nor U1334 (N_1334,N_1001,N_1150);
nor U1335 (N_1335,N_1030,N_1114);
and U1336 (N_1336,N_683,N_912);
nor U1337 (N_1337,N_1047,N_1003);
and U1338 (N_1338,N_940,N_1033);
nor U1339 (N_1339,N_1055,N_1091);
xnor U1340 (N_1340,N_802,N_1059);
or U1341 (N_1341,N_607,N_1148);
nand U1342 (N_1342,N_464,N_1152);
nor U1343 (N_1343,N_1078,N_1016);
nand U1344 (N_1344,N_1034,N_1143);
or U1345 (N_1345,N_1066,N_1167);
or U1346 (N_1346,In_10,N_1072);
or U1347 (N_1347,N_1128,N_1007);
nand U1348 (N_1348,N_1104,N_684);
nor U1349 (N_1349,In_637,N_606);
or U1350 (N_1350,N_1093,N_940);
nand U1351 (N_1351,N_876,N_1144);
or U1352 (N_1352,N_1019,N_897);
nor U1353 (N_1353,N_1130,N_1103);
and U1354 (N_1354,N_750,N_1179);
nor U1355 (N_1355,N_980,N_942);
nand U1356 (N_1356,N_1167,N_530);
or U1357 (N_1357,N_1001,N_1132);
nor U1358 (N_1358,N_1145,In_1261);
or U1359 (N_1359,N_712,N_1169);
and U1360 (N_1360,N_830,N_829);
and U1361 (N_1361,N_1093,N_1048);
nand U1362 (N_1362,N_1112,N_787);
nor U1363 (N_1363,N_697,N_1163);
or U1364 (N_1364,N_1170,N_1050);
and U1365 (N_1365,N_807,N_1004);
xor U1366 (N_1366,N_1193,N_861);
or U1367 (N_1367,N_1130,N_1023);
nand U1368 (N_1368,N_811,N_1187);
or U1369 (N_1369,N_927,N_1039);
or U1370 (N_1370,N_929,N_1094);
nand U1371 (N_1371,N_1102,N_942);
nand U1372 (N_1372,N_1021,N_141);
xnor U1373 (N_1373,N_982,N_1065);
nor U1374 (N_1374,N_1017,N_1045);
nor U1375 (N_1375,N_1164,N_1089);
or U1376 (N_1376,In_711,N_895);
nor U1377 (N_1377,N_1186,N_1021);
xnor U1378 (N_1378,N_1091,N_865);
xor U1379 (N_1379,N_1123,In_451);
xor U1380 (N_1380,N_1097,N_1080);
xnor U1381 (N_1381,In_670,N_935);
nand U1382 (N_1382,N_1085,N_1182);
xnor U1383 (N_1383,N_1030,In_808);
nand U1384 (N_1384,N_926,N_1165);
nand U1385 (N_1385,N_1118,N_1057);
or U1386 (N_1386,N_1198,N_1142);
nand U1387 (N_1387,N_1141,N_1123);
nor U1388 (N_1388,N_1109,N_1128);
nand U1389 (N_1389,N_843,N_1132);
and U1390 (N_1390,N_1072,N_1077);
xor U1391 (N_1391,N_1165,N_1093);
or U1392 (N_1392,N_633,N_1063);
nand U1393 (N_1393,N_1079,N_1105);
and U1394 (N_1394,N_530,N_787);
nand U1395 (N_1395,N_606,N_865);
nor U1396 (N_1396,N_1098,N_474);
nor U1397 (N_1397,In_474,N_1071);
nor U1398 (N_1398,N_1158,N_1020);
and U1399 (N_1399,N_1126,N_1129);
and U1400 (N_1400,N_1333,N_1334);
nor U1401 (N_1401,N_1279,N_1288);
nor U1402 (N_1402,N_1370,N_1209);
nand U1403 (N_1403,N_1391,N_1332);
xnor U1404 (N_1404,N_1392,N_1290);
nor U1405 (N_1405,N_1267,N_1344);
xor U1406 (N_1406,N_1379,N_1331);
nand U1407 (N_1407,N_1305,N_1256);
or U1408 (N_1408,N_1346,N_1356);
or U1409 (N_1409,N_1335,N_1214);
nand U1410 (N_1410,N_1295,N_1327);
xor U1411 (N_1411,N_1311,N_1272);
nand U1412 (N_1412,N_1397,N_1235);
nor U1413 (N_1413,N_1200,N_1342);
xor U1414 (N_1414,N_1247,N_1358);
xor U1415 (N_1415,N_1243,N_1225);
xnor U1416 (N_1416,N_1321,N_1329);
xor U1417 (N_1417,N_1398,N_1315);
nand U1418 (N_1418,N_1385,N_1278);
nand U1419 (N_1419,N_1367,N_1314);
nor U1420 (N_1420,N_1280,N_1396);
nand U1421 (N_1421,N_1368,N_1387);
nor U1422 (N_1422,N_1258,N_1263);
or U1423 (N_1423,N_1282,N_1325);
xor U1424 (N_1424,N_1217,N_1303);
nor U1425 (N_1425,N_1343,N_1328);
or U1426 (N_1426,N_1299,N_1259);
nor U1427 (N_1427,N_1202,N_1205);
and U1428 (N_1428,N_1316,N_1366);
and U1429 (N_1429,N_1248,N_1307);
or U1430 (N_1430,N_1241,N_1322);
xnor U1431 (N_1431,N_1292,N_1380);
nor U1432 (N_1432,N_1394,N_1340);
or U1433 (N_1433,N_1291,N_1339);
or U1434 (N_1434,N_1276,N_1338);
xor U1435 (N_1435,N_1306,N_1395);
xor U1436 (N_1436,N_1260,N_1281);
nand U1437 (N_1437,N_1312,N_1257);
xor U1438 (N_1438,N_1360,N_1294);
xnor U1439 (N_1439,N_1262,N_1233);
nand U1440 (N_1440,N_1353,N_1313);
nor U1441 (N_1441,N_1374,N_1249);
xor U1442 (N_1442,N_1293,N_1219);
and U1443 (N_1443,N_1271,N_1376);
xnor U1444 (N_1444,N_1347,N_1245);
nor U1445 (N_1445,N_1389,N_1352);
nor U1446 (N_1446,N_1213,N_1246);
nand U1447 (N_1447,N_1264,N_1227);
xor U1448 (N_1448,N_1359,N_1240);
and U1449 (N_1449,N_1230,N_1345);
nor U1450 (N_1450,N_1222,N_1285);
nor U1451 (N_1451,N_1355,N_1289);
or U1452 (N_1452,N_1323,N_1218);
nor U1453 (N_1453,N_1393,N_1348);
or U1454 (N_1454,N_1296,N_1317);
nand U1455 (N_1455,N_1275,N_1369);
nor U1456 (N_1456,N_1212,N_1269);
and U1457 (N_1457,N_1228,N_1224);
or U1458 (N_1458,N_1372,N_1261);
or U1459 (N_1459,N_1204,N_1252);
nand U1460 (N_1460,N_1373,N_1211);
nor U1461 (N_1461,N_1324,N_1283);
and U1462 (N_1462,N_1242,N_1377);
and U1463 (N_1463,N_1320,N_1255);
and U1464 (N_1464,N_1251,N_1201);
nor U1465 (N_1465,N_1337,N_1234);
or U1466 (N_1466,N_1206,N_1383);
xor U1467 (N_1467,N_1253,N_1351);
xnor U1468 (N_1468,N_1286,N_1302);
or U1469 (N_1469,N_1208,N_1236);
nor U1470 (N_1470,N_1326,N_1203);
xnor U1471 (N_1471,N_1309,N_1378);
nand U1472 (N_1472,N_1371,N_1221);
or U1473 (N_1473,N_1277,N_1254);
or U1474 (N_1474,N_1297,N_1266);
xor U1475 (N_1475,N_1300,N_1388);
xnor U1476 (N_1476,N_1232,N_1231);
nor U1477 (N_1477,N_1220,N_1363);
nand U1478 (N_1478,N_1284,N_1386);
or U1479 (N_1479,N_1298,N_1229);
nand U1480 (N_1480,N_1287,N_1226);
nand U1481 (N_1481,N_1223,N_1349);
nor U1482 (N_1482,N_1365,N_1207);
nand U1483 (N_1483,N_1310,N_1308);
nor U1484 (N_1484,N_1354,N_1330);
and U1485 (N_1485,N_1274,N_1270);
nand U1486 (N_1486,N_1361,N_1215);
nor U1487 (N_1487,N_1357,N_1216);
nand U1488 (N_1488,N_1341,N_1210);
xnor U1489 (N_1489,N_1265,N_1238);
and U1490 (N_1490,N_1301,N_1381);
or U1491 (N_1491,N_1364,N_1239);
xor U1492 (N_1492,N_1390,N_1336);
xnor U1493 (N_1493,N_1384,N_1350);
nand U1494 (N_1494,N_1250,N_1382);
or U1495 (N_1495,N_1304,N_1244);
and U1496 (N_1496,N_1319,N_1237);
or U1497 (N_1497,N_1362,N_1399);
xnor U1498 (N_1498,N_1375,N_1318);
or U1499 (N_1499,N_1268,N_1273);
nor U1500 (N_1500,N_1273,N_1347);
nor U1501 (N_1501,N_1258,N_1287);
xor U1502 (N_1502,N_1319,N_1261);
xor U1503 (N_1503,N_1282,N_1338);
nand U1504 (N_1504,N_1216,N_1280);
nand U1505 (N_1505,N_1355,N_1332);
and U1506 (N_1506,N_1260,N_1346);
nand U1507 (N_1507,N_1308,N_1393);
nand U1508 (N_1508,N_1205,N_1260);
and U1509 (N_1509,N_1321,N_1394);
nor U1510 (N_1510,N_1365,N_1370);
nand U1511 (N_1511,N_1323,N_1260);
nand U1512 (N_1512,N_1343,N_1210);
xnor U1513 (N_1513,N_1310,N_1347);
xnor U1514 (N_1514,N_1352,N_1207);
nand U1515 (N_1515,N_1250,N_1295);
nor U1516 (N_1516,N_1280,N_1249);
and U1517 (N_1517,N_1218,N_1376);
or U1518 (N_1518,N_1317,N_1343);
or U1519 (N_1519,N_1203,N_1271);
xnor U1520 (N_1520,N_1219,N_1226);
and U1521 (N_1521,N_1292,N_1367);
nand U1522 (N_1522,N_1286,N_1246);
and U1523 (N_1523,N_1306,N_1230);
nand U1524 (N_1524,N_1376,N_1204);
xor U1525 (N_1525,N_1283,N_1352);
xnor U1526 (N_1526,N_1337,N_1348);
nor U1527 (N_1527,N_1224,N_1207);
or U1528 (N_1528,N_1240,N_1322);
or U1529 (N_1529,N_1218,N_1209);
xor U1530 (N_1530,N_1388,N_1276);
and U1531 (N_1531,N_1311,N_1266);
and U1532 (N_1532,N_1336,N_1262);
nor U1533 (N_1533,N_1218,N_1242);
nor U1534 (N_1534,N_1258,N_1299);
and U1535 (N_1535,N_1308,N_1219);
nor U1536 (N_1536,N_1290,N_1393);
and U1537 (N_1537,N_1384,N_1223);
nor U1538 (N_1538,N_1223,N_1237);
and U1539 (N_1539,N_1227,N_1259);
and U1540 (N_1540,N_1204,N_1209);
nand U1541 (N_1541,N_1346,N_1285);
nor U1542 (N_1542,N_1321,N_1380);
nor U1543 (N_1543,N_1254,N_1214);
nor U1544 (N_1544,N_1310,N_1298);
nand U1545 (N_1545,N_1355,N_1249);
xnor U1546 (N_1546,N_1266,N_1298);
and U1547 (N_1547,N_1288,N_1383);
nor U1548 (N_1548,N_1335,N_1341);
xor U1549 (N_1549,N_1275,N_1263);
or U1550 (N_1550,N_1390,N_1341);
or U1551 (N_1551,N_1321,N_1393);
or U1552 (N_1552,N_1324,N_1365);
and U1553 (N_1553,N_1322,N_1306);
nand U1554 (N_1554,N_1210,N_1233);
xnor U1555 (N_1555,N_1346,N_1251);
and U1556 (N_1556,N_1369,N_1376);
nor U1557 (N_1557,N_1285,N_1326);
and U1558 (N_1558,N_1316,N_1396);
xnor U1559 (N_1559,N_1346,N_1244);
nand U1560 (N_1560,N_1234,N_1269);
xor U1561 (N_1561,N_1253,N_1393);
and U1562 (N_1562,N_1277,N_1347);
xnor U1563 (N_1563,N_1328,N_1226);
or U1564 (N_1564,N_1336,N_1216);
nor U1565 (N_1565,N_1271,N_1393);
and U1566 (N_1566,N_1257,N_1370);
or U1567 (N_1567,N_1228,N_1212);
nor U1568 (N_1568,N_1219,N_1207);
xor U1569 (N_1569,N_1313,N_1305);
nor U1570 (N_1570,N_1391,N_1337);
and U1571 (N_1571,N_1231,N_1335);
xor U1572 (N_1572,N_1270,N_1376);
xor U1573 (N_1573,N_1291,N_1299);
nor U1574 (N_1574,N_1293,N_1394);
or U1575 (N_1575,N_1389,N_1368);
and U1576 (N_1576,N_1390,N_1215);
and U1577 (N_1577,N_1341,N_1354);
xnor U1578 (N_1578,N_1370,N_1307);
nand U1579 (N_1579,N_1361,N_1246);
xnor U1580 (N_1580,N_1299,N_1379);
xor U1581 (N_1581,N_1283,N_1305);
nand U1582 (N_1582,N_1339,N_1392);
nor U1583 (N_1583,N_1266,N_1308);
and U1584 (N_1584,N_1368,N_1373);
xor U1585 (N_1585,N_1227,N_1350);
and U1586 (N_1586,N_1240,N_1320);
or U1587 (N_1587,N_1334,N_1317);
or U1588 (N_1588,N_1251,N_1359);
and U1589 (N_1589,N_1305,N_1381);
or U1590 (N_1590,N_1304,N_1236);
xor U1591 (N_1591,N_1388,N_1367);
xnor U1592 (N_1592,N_1384,N_1394);
nand U1593 (N_1593,N_1240,N_1222);
nor U1594 (N_1594,N_1323,N_1311);
and U1595 (N_1595,N_1363,N_1280);
nand U1596 (N_1596,N_1239,N_1363);
or U1597 (N_1597,N_1222,N_1372);
nand U1598 (N_1598,N_1300,N_1391);
nor U1599 (N_1599,N_1335,N_1201);
xnor U1600 (N_1600,N_1489,N_1544);
or U1601 (N_1601,N_1532,N_1491);
nor U1602 (N_1602,N_1446,N_1498);
xnor U1603 (N_1603,N_1499,N_1512);
nor U1604 (N_1604,N_1471,N_1466);
xor U1605 (N_1605,N_1570,N_1460);
or U1606 (N_1606,N_1463,N_1447);
xor U1607 (N_1607,N_1482,N_1445);
or U1608 (N_1608,N_1502,N_1540);
or U1609 (N_1609,N_1516,N_1587);
or U1610 (N_1610,N_1593,N_1479);
xor U1611 (N_1611,N_1421,N_1592);
xnor U1612 (N_1612,N_1572,N_1550);
nor U1613 (N_1613,N_1530,N_1406);
xor U1614 (N_1614,N_1432,N_1433);
or U1615 (N_1615,N_1443,N_1563);
nand U1616 (N_1616,N_1430,N_1477);
or U1617 (N_1617,N_1413,N_1545);
xor U1618 (N_1618,N_1454,N_1425);
nor U1619 (N_1619,N_1458,N_1495);
or U1620 (N_1620,N_1555,N_1528);
nand U1621 (N_1621,N_1529,N_1537);
nand U1622 (N_1622,N_1574,N_1598);
nand U1623 (N_1623,N_1575,N_1594);
or U1624 (N_1624,N_1401,N_1405);
and U1625 (N_1625,N_1467,N_1581);
nand U1626 (N_1626,N_1493,N_1452);
nor U1627 (N_1627,N_1553,N_1449);
nor U1628 (N_1628,N_1585,N_1588);
and U1629 (N_1629,N_1514,N_1518);
and U1630 (N_1630,N_1408,N_1486);
xor U1631 (N_1631,N_1539,N_1461);
and U1632 (N_1632,N_1577,N_1507);
and U1633 (N_1633,N_1474,N_1591);
xor U1634 (N_1634,N_1549,N_1568);
nor U1635 (N_1635,N_1462,N_1451);
xnor U1636 (N_1636,N_1464,N_1571);
nand U1637 (N_1637,N_1519,N_1557);
and U1638 (N_1638,N_1534,N_1582);
and U1639 (N_1639,N_1481,N_1586);
and U1640 (N_1640,N_1526,N_1543);
nor U1641 (N_1641,N_1513,N_1459);
nand U1642 (N_1642,N_1444,N_1475);
xnor U1643 (N_1643,N_1522,N_1567);
or U1644 (N_1644,N_1435,N_1485);
nor U1645 (N_1645,N_1440,N_1455);
xnor U1646 (N_1646,N_1415,N_1448);
nand U1647 (N_1647,N_1465,N_1450);
nand U1648 (N_1648,N_1584,N_1510);
xor U1649 (N_1649,N_1535,N_1580);
nand U1650 (N_1650,N_1473,N_1525);
and U1651 (N_1651,N_1480,N_1517);
xor U1652 (N_1652,N_1578,N_1402);
or U1653 (N_1653,N_1441,N_1538);
nand U1654 (N_1654,N_1558,N_1494);
nor U1655 (N_1655,N_1503,N_1416);
nor U1656 (N_1656,N_1547,N_1428);
nor U1657 (N_1657,N_1566,N_1434);
or U1658 (N_1658,N_1599,N_1497);
nor U1659 (N_1659,N_1411,N_1515);
xnor U1660 (N_1660,N_1403,N_1478);
or U1661 (N_1661,N_1409,N_1490);
nor U1662 (N_1662,N_1492,N_1483);
and U1663 (N_1663,N_1583,N_1419);
xnor U1664 (N_1664,N_1590,N_1436);
and U1665 (N_1665,N_1410,N_1596);
nor U1666 (N_1666,N_1511,N_1505);
and U1667 (N_1667,N_1442,N_1429);
and U1668 (N_1668,N_1438,N_1509);
nor U1669 (N_1669,N_1439,N_1521);
or U1670 (N_1670,N_1595,N_1597);
nor U1671 (N_1671,N_1542,N_1564);
nor U1672 (N_1672,N_1551,N_1536);
and U1673 (N_1673,N_1569,N_1424);
xor U1674 (N_1674,N_1559,N_1422);
xor U1675 (N_1675,N_1476,N_1456);
or U1676 (N_1676,N_1423,N_1457);
and U1677 (N_1677,N_1579,N_1420);
xnor U1678 (N_1678,N_1520,N_1418);
nand U1679 (N_1679,N_1453,N_1506);
nor U1680 (N_1680,N_1508,N_1533);
and U1681 (N_1681,N_1414,N_1484);
and U1682 (N_1682,N_1400,N_1576);
nor U1683 (N_1683,N_1427,N_1417);
nor U1684 (N_1684,N_1488,N_1500);
and U1685 (N_1685,N_1556,N_1496);
nor U1686 (N_1686,N_1426,N_1589);
xor U1687 (N_1687,N_1541,N_1548);
nand U1688 (N_1688,N_1573,N_1437);
or U1689 (N_1689,N_1501,N_1472);
xor U1690 (N_1690,N_1469,N_1504);
and U1691 (N_1691,N_1431,N_1546);
or U1692 (N_1692,N_1552,N_1523);
nor U1693 (N_1693,N_1527,N_1524);
nand U1694 (N_1694,N_1531,N_1407);
and U1695 (N_1695,N_1561,N_1412);
nor U1696 (N_1696,N_1562,N_1468);
xnor U1697 (N_1697,N_1470,N_1554);
nand U1698 (N_1698,N_1487,N_1560);
nand U1699 (N_1699,N_1565,N_1404);
nand U1700 (N_1700,N_1423,N_1589);
and U1701 (N_1701,N_1442,N_1555);
nand U1702 (N_1702,N_1463,N_1553);
xor U1703 (N_1703,N_1453,N_1500);
xnor U1704 (N_1704,N_1496,N_1579);
nand U1705 (N_1705,N_1538,N_1492);
nor U1706 (N_1706,N_1439,N_1418);
or U1707 (N_1707,N_1540,N_1503);
and U1708 (N_1708,N_1437,N_1572);
nor U1709 (N_1709,N_1411,N_1486);
and U1710 (N_1710,N_1437,N_1432);
nor U1711 (N_1711,N_1441,N_1517);
nor U1712 (N_1712,N_1580,N_1499);
and U1713 (N_1713,N_1423,N_1432);
and U1714 (N_1714,N_1468,N_1575);
xnor U1715 (N_1715,N_1419,N_1529);
or U1716 (N_1716,N_1434,N_1541);
and U1717 (N_1717,N_1415,N_1453);
or U1718 (N_1718,N_1561,N_1592);
xnor U1719 (N_1719,N_1538,N_1411);
nand U1720 (N_1720,N_1475,N_1468);
nand U1721 (N_1721,N_1514,N_1571);
or U1722 (N_1722,N_1457,N_1524);
and U1723 (N_1723,N_1596,N_1563);
nand U1724 (N_1724,N_1597,N_1505);
xnor U1725 (N_1725,N_1428,N_1432);
or U1726 (N_1726,N_1419,N_1494);
and U1727 (N_1727,N_1552,N_1508);
and U1728 (N_1728,N_1581,N_1587);
xor U1729 (N_1729,N_1404,N_1524);
xor U1730 (N_1730,N_1537,N_1473);
nor U1731 (N_1731,N_1465,N_1484);
nor U1732 (N_1732,N_1432,N_1477);
nand U1733 (N_1733,N_1417,N_1509);
nor U1734 (N_1734,N_1409,N_1446);
or U1735 (N_1735,N_1527,N_1557);
nand U1736 (N_1736,N_1533,N_1581);
and U1737 (N_1737,N_1516,N_1554);
xor U1738 (N_1738,N_1525,N_1485);
or U1739 (N_1739,N_1411,N_1415);
nor U1740 (N_1740,N_1466,N_1486);
and U1741 (N_1741,N_1458,N_1566);
or U1742 (N_1742,N_1496,N_1596);
xor U1743 (N_1743,N_1508,N_1440);
or U1744 (N_1744,N_1590,N_1461);
nand U1745 (N_1745,N_1590,N_1526);
nand U1746 (N_1746,N_1410,N_1547);
xnor U1747 (N_1747,N_1595,N_1570);
nor U1748 (N_1748,N_1535,N_1482);
xor U1749 (N_1749,N_1429,N_1417);
nand U1750 (N_1750,N_1585,N_1535);
or U1751 (N_1751,N_1495,N_1549);
nand U1752 (N_1752,N_1517,N_1576);
nor U1753 (N_1753,N_1473,N_1506);
nand U1754 (N_1754,N_1546,N_1597);
nor U1755 (N_1755,N_1594,N_1527);
nand U1756 (N_1756,N_1558,N_1442);
and U1757 (N_1757,N_1499,N_1524);
nand U1758 (N_1758,N_1447,N_1512);
nand U1759 (N_1759,N_1489,N_1407);
nor U1760 (N_1760,N_1527,N_1455);
xor U1761 (N_1761,N_1532,N_1511);
xnor U1762 (N_1762,N_1490,N_1588);
or U1763 (N_1763,N_1526,N_1413);
nor U1764 (N_1764,N_1410,N_1406);
xnor U1765 (N_1765,N_1495,N_1574);
nand U1766 (N_1766,N_1507,N_1500);
and U1767 (N_1767,N_1581,N_1460);
or U1768 (N_1768,N_1407,N_1594);
nand U1769 (N_1769,N_1496,N_1527);
nand U1770 (N_1770,N_1491,N_1485);
xor U1771 (N_1771,N_1575,N_1464);
or U1772 (N_1772,N_1515,N_1464);
nor U1773 (N_1773,N_1499,N_1433);
or U1774 (N_1774,N_1456,N_1489);
nor U1775 (N_1775,N_1453,N_1459);
nand U1776 (N_1776,N_1411,N_1490);
and U1777 (N_1777,N_1550,N_1500);
nor U1778 (N_1778,N_1464,N_1536);
and U1779 (N_1779,N_1405,N_1513);
and U1780 (N_1780,N_1594,N_1416);
and U1781 (N_1781,N_1516,N_1579);
or U1782 (N_1782,N_1538,N_1552);
or U1783 (N_1783,N_1416,N_1575);
nor U1784 (N_1784,N_1423,N_1456);
nand U1785 (N_1785,N_1591,N_1598);
nand U1786 (N_1786,N_1585,N_1598);
nor U1787 (N_1787,N_1473,N_1499);
nand U1788 (N_1788,N_1544,N_1534);
nand U1789 (N_1789,N_1442,N_1591);
or U1790 (N_1790,N_1506,N_1499);
xnor U1791 (N_1791,N_1476,N_1408);
xnor U1792 (N_1792,N_1509,N_1520);
and U1793 (N_1793,N_1525,N_1455);
nor U1794 (N_1794,N_1595,N_1574);
xnor U1795 (N_1795,N_1440,N_1575);
xor U1796 (N_1796,N_1497,N_1504);
or U1797 (N_1797,N_1573,N_1508);
nand U1798 (N_1798,N_1403,N_1424);
nor U1799 (N_1799,N_1489,N_1581);
xnor U1800 (N_1800,N_1788,N_1658);
nand U1801 (N_1801,N_1621,N_1672);
nor U1802 (N_1802,N_1663,N_1636);
and U1803 (N_1803,N_1684,N_1790);
xnor U1804 (N_1804,N_1757,N_1784);
nand U1805 (N_1805,N_1720,N_1601);
and U1806 (N_1806,N_1727,N_1606);
nand U1807 (N_1807,N_1722,N_1662);
nand U1808 (N_1808,N_1660,N_1744);
xnor U1809 (N_1809,N_1779,N_1705);
nand U1810 (N_1810,N_1768,N_1664);
xor U1811 (N_1811,N_1773,N_1690);
xnor U1812 (N_1812,N_1761,N_1716);
nor U1813 (N_1813,N_1692,N_1751);
xor U1814 (N_1814,N_1627,N_1702);
and U1815 (N_1815,N_1798,N_1670);
xor U1816 (N_1816,N_1615,N_1654);
or U1817 (N_1817,N_1721,N_1776);
nand U1818 (N_1818,N_1647,N_1715);
xnor U1819 (N_1819,N_1703,N_1674);
nand U1820 (N_1820,N_1603,N_1725);
or U1821 (N_1821,N_1632,N_1626);
nand U1822 (N_1822,N_1650,N_1764);
nor U1823 (N_1823,N_1657,N_1762);
or U1824 (N_1824,N_1668,N_1750);
nand U1825 (N_1825,N_1775,N_1707);
nand U1826 (N_1826,N_1619,N_1719);
nor U1827 (N_1827,N_1700,N_1602);
or U1828 (N_1828,N_1780,N_1641);
and U1829 (N_1829,N_1679,N_1754);
nor U1830 (N_1830,N_1649,N_1613);
xnor U1831 (N_1831,N_1617,N_1782);
nor U1832 (N_1832,N_1749,N_1781);
xor U1833 (N_1833,N_1624,N_1607);
nor U1834 (N_1834,N_1767,N_1753);
or U1835 (N_1835,N_1659,N_1785);
or U1836 (N_1836,N_1651,N_1644);
or U1837 (N_1837,N_1665,N_1708);
nand U1838 (N_1838,N_1673,N_1728);
and U1839 (N_1839,N_1612,N_1697);
and U1840 (N_1840,N_1709,N_1730);
and U1841 (N_1841,N_1683,N_1699);
and U1842 (N_1842,N_1706,N_1710);
nor U1843 (N_1843,N_1772,N_1676);
nor U1844 (N_1844,N_1666,N_1633);
xnor U1845 (N_1845,N_1731,N_1678);
or U1846 (N_1846,N_1696,N_1743);
and U1847 (N_1847,N_1777,N_1738);
xor U1848 (N_1848,N_1799,N_1765);
or U1849 (N_1849,N_1638,N_1656);
nor U1850 (N_1850,N_1688,N_1723);
xnor U1851 (N_1851,N_1763,N_1685);
and U1852 (N_1852,N_1600,N_1667);
nor U1853 (N_1853,N_1620,N_1682);
xnor U1854 (N_1854,N_1616,N_1655);
nand U1855 (N_1855,N_1739,N_1746);
and U1856 (N_1856,N_1693,N_1695);
or U1857 (N_1857,N_1628,N_1604);
nor U1858 (N_1858,N_1736,N_1745);
and U1859 (N_1859,N_1766,N_1791);
or U1860 (N_1860,N_1786,N_1689);
and U1861 (N_1861,N_1712,N_1759);
or U1862 (N_1862,N_1635,N_1642);
nand U1863 (N_1863,N_1783,N_1758);
or U1864 (N_1864,N_1681,N_1748);
nor U1865 (N_1865,N_1741,N_1614);
and U1866 (N_1866,N_1629,N_1717);
nand U1867 (N_1867,N_1724,N_1769);
nand U1868 (N_1868,N_1609,N_1634);
or U1869 (N_1869,N_1778,N_1646);
nor U1870 (N_1870,N_1735,N_1729);
or U1871 (N_1871,N_1752,N_1680);
or U1872 (N_1872,N_1795,N_1793);
and U1873 (N_1873,N_1610,N_1698);
and U1874 (N_1874,N_1733,N_1755);
and U1875 (N_1875,N_1605,N_1675);
nand U1876 (N_1876,N_1630,N_1797);
nor U1877 (N_1877,N_1608,N_1623);
xor U1878 (N_1878,N_1639,N_1794);
and U1879 (N_1879,N_1653,N_1669);
nor U1880 (N_1880,N_1711,N_1770);
and U1881 (N_1881,N_1789,N_1637);
xor U1882 (N_1882,N_1796,N_1652);
nor U1883 (N_1883,N_1640,N_1691);
nand U1884 (N_1884,N_1687,N_1694);
or U1885 (N_1885,N_1726,N_1771);
xnor U1886 (N_1886,N_1734,N_1618);
nand U1887 (N_1887,N_1737,N_1714);
and U1888 (N_1888,N_1787,N_1774);
and U1889 (N_1889,N_1740,N_1732);
nor U1890 (N_1890,N_1713,N_1671);
nor U1891 (N_1891,N_1661,N_1622);
or U1892 (N_1892,N_1648,N_1747);
nor U1893 (N_1893,N_1631,N_1704);
and U1894 (N_1894,N_1686,N_1718);
xor U1895 (N_1895,N_1677,N_1701);
nor U1896 (N_1896,N_1742,N_1643);
xnor U1897 (N_1897,N_1792,N_1756);
nor U1898 (N_1898,N_1760,N_1625);
and U1899 (N_1899,N_1645,N_1611);
nor U1900 (N_1900,N_1773,N_1625);
and U1901 (N_1901,N_1781,N_1777);
and U1902 (N_1902,N_1738,N_1629);
xnor U1903 (N_1903,N_1787,N_1702);
nor U1904 (N_1904,N_1747,N_1759);
or U1905 (N_1905,N_1660,N_1616);
and U1906 (N_1906,N_1752,N_1672);
xnor U1907 (N_1907,N_1752,N_1614);
or U1908 (N_1908,N_1603,N_1753);
and U1909 (N_1909,N_1775,N_1774);
nand U1910 (N_1910,N_1740,N_1625);
nor U1911 (N_1911,N_1728,N_1770);
nor U1912 (N_1912,N_1712,N_1741);
or U1913 (N_1913,N_1603,N_1640);
and U1914 (N_1914,N_1793,N_1627);
or U1915 (N_1915,N_1794,N_1710);
nand U1916 (N_1916,N_1611,N_1788);
nand U1917 (N_1917,N_1667,N_1790);
xnor U1918 (N_1918,N_1626,N_1645);
nor U1919 (N_1919,N_1761,N_1616);
and U1920 (N_1920,N_1701,N_1679);
xor U1921 (N_1921,N_1608,N_1660);
nand U1922 (N_1922,N_1729,N_1632);
and U1923 (N_1923,N_1767,N_1685);
xor U1924 (N_1924,N_1686,N_1689);
nand U1925 (N_1925,N_1794,N_1627);
nand U1926 (N_1926,N_1733,N_1619);
nor U1927 (N_1927,N_1799,N_1749);
or U1928 (N_1928,N_1787,N_1691);
xor U1929 (N_1929,N_1767,N_1605);
or U1930 (N_1930,N_1754,N_1738);
and U1931 (N_1931,N_1688,N_1613);
xor U1932 (N_1932,N_1704,N_1700);
nand U1933 (N_1933,N_1671,N_1744);
nor U1934 (N_1934,N_1671,N_1712);
nor U1935 (N_1935,N_1699,N_1736);
or U1936 (N_1936,N_1627,N_1694);
xor U1937 (N_1937,N_1751,N_1647);
and U1938 (N_1938,N_1771,N_1700);
nor U1939 (N_1939,N_1607,N_1658);
nor U1940 (N_1940,N_1636,N_1772);
and U1941 (N_1941,N_1723,N_1691);
nand U1942 (N_1942,N_1732,N_1687);
xnor U1943 (N_1943,N_1792,N_1622);
or U1944 (N_1944,N_1715,N_1640);
nor U1945 (N_1945,N_1791,N_1677);
nor U1946 (N_1946,N_1643,N_1656);
nand U1947 (N_1947,N_1700,N_1754);
or U1948 (N_1948,N_1656,N_1714);
xnor U1949 (N_1949,N_1763,N_1737);
xor U1950 (N_1950,N_1605,N_1657);
and U1951 (N_1951,N_1623,N_1668);
xor U1952 (N_1952,N_1725,N_1774);
and U1953 (N_1953,N_1640,N_1738);
and U1954 (N_1954,N_1767,N_1765);
and U1955 (N_1955,N_1709,N_1737);
nand U1956 (N_1956,N_1761,N_1684);
xor U1957 (N_1957,N_1646,N_1686);
xnor U1958 (N_1958,N_1691,N_1722);
and U1959 (N_1959,N_1744,N_1699);
nor U1960 (N_1960,N_1676,N_1763);
nand U1961 (N_1961,N_1758,N_1652);
nand U1962 (N_1962,N_1791,N_1753);
nand U1963 (N_1963,N_1629,N_1701);
xor U1964 (N_1964,N_1685,N_1641);
xnor U1965 (N_1965,N_1629,N_1687);
xnor U1966 (N_1966,N_1701,N_1654);
nand U1967 (N_1967,N_1728,N_1749);
and U1968 (N_1968,N_1632,N_1609);
xor U1969 (N_1969,N_1795,N_1750);
and U1970 (N_1970,N_1666,N_1630);
and U1971 (N_1971,N_1767,N_1692);
nand U1972 (N_1972,N_1767,N_1650);
or U1973 (N_1973,N_1685,N_1635);
nand U1974 (N_1974,N_1649,N_1642);
nand U1975 (N_1975,N_1708,N_1685);
or U1976 (N_1976,N_1736,N_1613);
or U1977 (N_1977,N_1601,N_1731);
xor U1978 (N_1978,N_1729,N_1744);
xnor U1979 (N_1979,N_1607,N_1700);
nand U1980 (N_1980,N_1798,N_1736);
nor U1981 (N_1981,N_1703,N_1774);
and U1982 (N_1982,N_1776,N_1620);
or U1983 (N_1983,N_1614,N_1745);
or U1984 (N_1984,N_1789,N_1780);
and U1985 (N_1985,N_1637,N_1762);
xnor U1986 (N_1986,N_1641,N_1682);
and U1987 (N_1987,N_1682,N_1707);
nand U1988 (N_1988,N_1694,N_1771);
nand U1989 (N_1989,N_1720,N_1678);
xnor U1990 (N_1990,N_1704,N_1723);
nor U1991 (N_1991,N_1741,N_1750);
xnor U1992 (N_1992,N_1655,N_1639);
xnor U1993 (N_1993,N_1784,N_1684);
and U1994 (N_1994,N_1679,N_1619);
or U1995 (N_1995,N_1603,N_1644);
nor U1996 (N_1996,N_1709,N_1633);
xor U1997 (N_1997,N_1744,N_1779);
xor U1998 (N_1998,N_1665,N_1778);
nor U1999 (N_1999,N_1676,N_1741);
or U2000 (N_2000,N_1815,N_1800);
and U2001 (N_2001,N_1942,N_1953);
xor U2002 (N_2002,N_1929,N_1838);
or U2003 (N_2003,N_1978,N_1911);
or U2004 (N_2004,N_1835,N_1857);
and U2005 (N_2005,N_1892,N_1991);
or U2006 (N_2006,N_1941,N_1869);
or U2007 (N_2007,N_1845,N_1971);
and U2008 (N_2008,N_1844,N_1822);
xnor U2009 (N_2009,N_1957,N_1837);
or U2010 (N_2010,N_1908,N_1875);
nor U2011 (N_2011,N_1823,N_1950);
or U2012 (N_2012,N_1810,N_1930);
xor U2013 (N_2013,N_1905,N_1829);
or U2014 (N_2014,N_1945,N_1910);
xor U2015 (N_2015,N_1856,N_1985);
nor U2016 (N_2016,N_1917,N_1867);
and U2017 (N_2017,N_1820,N_1847);
nand U2018 (N_2018,N_1934,N_1851);
nand U2019 (N_2019,N_1955,N_1956);
nand U2020 (N_2020,N_1962,N_1988);
xor U2021 (N_2021,N_1969,N_1889);
nor U2022 (N_2022,N_1992,N_1984);
nand U2023 (N_2023,N_1968,N_1965);
nor U2024 (N_2024,N_1814,N_1949);
and U2025 (N_2025,N_1891,N_1848);
nand U2026 (N_2026,N_1938,N_1860);
nor U2027 (N_2027,N_1913,N_1931);
or U2028 (N_2028,N_1927,N_1979);
nand U2029 (N_2029,N_1983,N_1817);
and U2030 (N_2030,N_1887,N_1987);
nor U2031 (N_2031,N_1967,N_1808);
nor U2032 (N_2032,N_1964,N_1895);
and U2033 (N_2033,N_1853,N_1998);
nand U2034 (N_2034,N_1854,N_1870);
nor U2035 (N_2035,N_1813,N_1958);
nor U2036 (N_2036,N_1970,N_1852);
nand U2037 (N_2037,N_1874,N_1846);
xnor U2038 (N_2038,N_1919,N_1937);
xor U2039 (N_2039,N_1882,N_1995);
xnor U2040 (N_2040,N_1818,N_1805);
nor U2041 (N_2041,N_1948,N_1943);
nor U2042 (N_2042,N_1916,N_1861);
or U2043 (N_2043,N_1824,N_1862);
or U2044 (N_2044,N_1932,N_1909);
nor U2045 (N_2045,N_1906,N_1939);
and U2046 (N_2046,N_1816,N_1963);
or U2047 (N_2047,N_1825,N_1961);
nand U2048 (N_2048,N_1947,N_1855);
or U2049 (N_2049,N_1986,N_1878);
and U2050 (N_2050,N_1974,N_1936);
or U2051 (N_2051,N_1952,N_1876);
or U2052 (N_2052,N_1868,N_1993);
xnor U2053 (N_2053,N_1806,N_1996);
xnor U2054 (N_2054,N_1951,N_1833);
xnor U2055 (N_2055,N_1839,N_1826);
or U2056 (N_2056,N_1954,N_1920);
and U2057 (N_2057,N_1894,N_1897);
nor U2058 (N_2058,N_1831,N_1828);
nand U2059 (N_2059,N_1914,N_1802);
xor U2060 (N_2060,N_1830,N_1903);
nand U2061 (N_2061,N_1863,N_1886);
or U2062 (N_2062,N_1900,N_1821);
and U2063 (N_2063,N_1843,N_1858);
nand U2064 (N_2064,N_1926,N_1866);
nand U2065 (N_2065,N_1977,N_1980);
nor U2066 (N_2066,N_1881,N_1827);
nand U2067 (N_2067,N_1896,N_1975);
or U2068 (N_2068,N_1901,N_1994);
nor U2069 (N_2069,N_1966,N_1890);
or U2070 (N_2070,N_1864,N_1976);
nor U2071 (N_2071,N_1877,N_1884);
nor U2072 (N_2072,N_1918,N_1925);
and U2073 (N_2073,N_1849,N_1834);
or U2074 (N_2074,N_1946,N_1928);
xor U2075 (N_2075,N_1923,N_1997);
or U2076 (N_2076,N_1842,N_1915);
nand U2077 (N_2077,N_1811,N_1999);
xor U2078 (N_2078,N_1819,N_1883);
nor U2079 (N_2079,N_1907,N_1804);
xnor U2080 (N_2080,N_1888,N_1836);
nor U2081 (N_2081,N_1933,N_1865);
and U2082 (N_2082,N_1924,N_1960);
xnor U2083 (N_2083,N_1850,N_1879);
xor U2084 (N_2084,N_1940,N_1801);
nand U2085 (N_2085,N_1880,N_1899);
xor U2086 (N_2086,N_1972,N_1944);
and U2087 (N_2087,N_1872,N_1840);
nand U2088 (N_2088,N_1859,N_1922);
xor U2089 (N_2089,N_1902,N_1959);
nor U2090 (N_2090,N_1871,N_1893);
nor U2091 (N_2091,N_1873,N_1912);
or U2092 (N_2092,N_1803,N_1904);
nor U2093 (N_2093,N_1921,N_1841);
nand U2094 (N_2094,N_1973,N_1809);
nor U2095 (N_2095,N_1812,N_1990);
and U2096 (N_2096,N_1982,N_1935);
xor U2097 (N_2097,N_1981,N_1885);
or U2098 (N_2098,N_1807,N_1898);
or U2099 (N_2099,N_1832,N_1989);
nor U2100 (N_2100,N_1993,N_1893);
xnor U2101 (N_2101,N_1913,N_1878);
and U2102 (N_2102,N_1966,N_1864);
nor U2103 (N_2103,N_1859,N_1817);
nand U2104 (N_2104,N_1972,N_1849);
nor U2105 (N_2105,N_1953,N_1937);
nor U2106 (N_2106,N_1887,N_1992);
nor U2107 (N_2107,N_1864,N_1988);
xnor U2108 (N_2108,N_1829,N_1964);
or U2109 (N_2109,N_1847,N_1840);
xnor U2110 (N_2110,N_1926,N_1932);
nand U2111 (N_2111,N_1934,N_1832);
nor U2112 (N_2112,N_1988,N_1821);
xor U2113 (N_2113,N_1995,N_1998);
or U2114 (N_2114,N_1852,N_1811);
or U2115 (N_2115,N_1847,N_1915);
and U2116 (N_2116,N_1937,N_1895);
and U2117 (N_2117,N_1992,N_1947);
nor U2118 (N_2118,N_1885,N_1999);
xor U2119 (N_2119,N_1820,N_1995);
or U2120 (N_2120,N_1843,N_1989);
nand U2121 (N_2121,N_1947,N_1921);
nor U2122 (N_2122,N_1991,N_1968);
and U2123 (N_2123,N_1854,N_1881);
and U2124 (N_2124,N_1876,N_1842);
nand U2125 (N_2125,N_1909,N_1867);
or U2126 (N_2126,N_1882,N_1852);
or U2127 (N_2127,N_1919,N_1941);
xnor U2128 (N_2128,N_1988,N_1803);
and U2129 (N_2129,N_1822,N_1953);
and U2130 (N_2130,N_1992,N_1996);
or U2131 (N_2131,N_1889,N_1954);
and U2132 (N_2132,N_1801,N_1824);
or U2133 (N_2133,N_1849,N_1879);
xor U2134 (N_2134,N_1964,N_1974);
xor U2135 (N_2135,N_1859,N_1926);
or U2136 (N_2136,N_1876,N_1990);
and U2137 (N_2137,N_1993,N_1992);
nor U2138 (N_2138,N_1851,N_1870);
and U2139 (N_2139,N_1829,N_1873);
nand U2140 (N_2140,N_1942,N_1801);
and U2141 (N_2141,N_1825,N_1856);
nor U2142 (N_2142,N_1935,N_1807);
nand U2143 (N_2143,N_1809,N_1874);
and U2144 (N_2144,N_1889,N_1806);
or U2145 (N_2145,N_1828,N_1942);
and U2146 (N_2146,N_1806,N_1991);
or U2147 (N_2147,N_1888,N_1875);
and U2148 (N_2148,N_1802,N_1976);
and U2149 (N_2149,N_1827,N_1880);
nor U2150 (N_2150,N_1953,N_1876);
and U2151 (N_2151,N_1833,N_1960);
or U2152 (N_2152,N_1980,N_1823);
nor U2153 (N_2153,N_1813,N_1806);
nor U2154 (N_2154,N_1963,N_1988);
nand U2155 (N_2155,N_1947,N_1807);
nor U2156 (N_2156,N_1914,N_1992);
xor U2157 (N_2157,N_1984,N_1949);
xor U2158 (N_2158,N_1935,N_1955);
nor U2159 (N_2159,N_1888,N_1827);
nor U2160 (N_2160,N_1832,N_1869);
xor U2161 (N_2161,N_1954,N_1859);
and U2162 (N_2162,N_1979,N_1997);
and U2163 (N_2163,N_1813,N_1938);
nand U2164 (N_2164,N_1855,N_1930);
nand U2165 (N_2165,N_1900,N_1802);
nor U2166 (N_2166,N_1873,N_1830);
xnor U2167 (N_2167,N_1934,N_1830);
nor U2168 (N_2168,N_1912,N_1901);
nand U2169 (N_2169,N_1969,N_1966);
nor U2170 (N_2170,N_1867,N_1837);
and U2171 (N_2171,N_1892,N_1815);
or U2172 (N_2172,N_1956,N_1816);
nand U2173 (N_2173,N_1889,N_1922);
xor U2174 (N_2174,N_1954,N_1816);
or U2175 (N_2175,N_1845,N_1835);
nor U2176 (N_2176,N_1982,N_1836);
and U2177 (N_2177,N_1919,N_1902);
nor U2178 (N_2178,N_1847,N_1833);
nand U2179 (N_2179,N_1995,N_1993);
xor U2180 (N_2180,N_1935,N_1920);
nand U2181 (N_2181,N_1860,N_1855);
nand U2182 (N_2182,N_1982,N_1918);
or U2183 (N_2183,N_1976,N_1869);
xor U2184 (N_2184,N_1812,N_1807);
or U2185 (N_2185,N_1894,N_1827);
xnor U2186 (N_2186,N_1974,N_1820);
nor U2187 (N_2187,N_1864,N_1813);
and U2188 (N_2188,N_1958,N_1957);
xor U2189 (N_2189,N_1969,N_1821);
xor U2190 (N_2190,N_1881,N_1842);
nor U2191 (N_2191,N_1955,N_1927);
or U2192 (N_2192,N_1853,N_1840);
nor U2193 (N_2193,N_1856,N_1946);
nor U2194 (N_2194,N_1848,N_1874);
nand U2195 (N_2195,N_1817,N_1993);
or U2196 (N_2196,N_1985,N_1955);
nor U2197 (N_2197,N_1895,N_1871);
and U2198 (N_2198,N_1995,N_1915);
or U2199 (N_2199,N_1830,N_1966);
nand U2200 (N_2200,N_2060,N_2170);
nand U2201 (N_2201,N_2125,N_2191);
nor U2202 (N_2202,N_2019,N_2114);
and U2203 (N_2203,N_2068,N_2065);
nor U2204 (N_2204,N_2129,N_2111);
or U2205 (N_2205,N_2102,N_2087);
xnor U2206 (N_2206,N_2091,N_2122);
nor U2207 (N_2207,N_2023,N_2185);
xnor U2208 (N_2208,N_2014,N_2131);
xnor U2209 (N_2209,N_2105,N_2006);
and U2210 (N_2210,N_2187,N_2186);
nand U2211 (N_2211,N_2184,N_2126);
nand U2212 (N_2212,N_2045,N_2034);
and U2213 (N_2213,N_2152,N_2144);
xor U2214 (N_2214,N_2029,N_2199);
and U2215 (N_2215,N_2047,N_2067);
nand U2216 (N_2216,N_2176,N_2048);
nor U2217 (N_2217,N_2095,N_2033);
or U2218 (N_2218,N_2072,N_2017);
nor U2219 (N_2219,N_2112,N_2054);
nand U2220 (N_2220,N_2062,N_2008);
or U2221 (N_2221,N_2197,N_2077);
xor U2222 (N_2222,N_2026,N_2093);
or U2223 (N_2223,N_2041,N_2022);
and U2224 (N_2224,N_2084,N_2110);
xor U2225 (N_2225,N_2178,N_2027);
xnor U2226 (N_2226,N_2043,N_2113);
and U2227 (N_2227,N_2037,N_2153);
and U2228 (N_2228,N_2150,N_2073);
and U2229 (N_2229,N_2015,N_2128);
nor U2230 (N_2230,N_2013,N_2012);
nor U2231 (N_2231,N_2075,N_2154);
or U2232 (N_2232,N_2036,N_2116);
or U2233 (N_2233,N_2143,N_2040);
nor U2234 (N_2234,N_2192,N_2009);
xnor U2235 (N_2235,N_2133,N_2140);
and U2236 (N_2236,N_2139,N_2002);
or U2237 (N_2237,N_2051,N_2085);
or U2238 (N_2238,N_2127,N_2123);
nand U2239 (N_2239,N_2094,N_2064);
nor U2240 (N_2240,N_2195,N_2030);
and U2241 (N_2241,N_2179,N_2104);
or U2242 (N_2242,N_2096,N_2171);
xor U2243 (N_2243,N_2103,N_2115);
nor U2244 (N_2244,N_2039,N_2046);
nand U2245 (N_2245,N_2149,N_2090);
nor U2246 (N_2246,N_2099,N_2003);
xor U2247 (N_2247,N_2145,N_2000);
nand U2248 (N_2248,N_2194,N_2098);
or U2249 (N_2249,N_2097,N_2025);
and U2250 (N_2250,N_2190,N_2196);
and U2251 (N_2251,N_2169,N_2052);
nor U2252 (N_2252,N_2038,N_2167);
and U2253 (N_2253,N_2193,N_2120);
nand U2254 (N_2254,N_2181,N_2134);
and U2255 (N_2255,N_2079,N_2172);
nand U2256 (N_2256,N_2004,N_2141);
nand U2257 (N_2257,N_2146,N_2021);
nand U2258 (N_2258,N_2118,N_2078);
or U2259 (N_2259,N_2159,N_2157);
and U2260 (N_2260,N_2138,N_2020);
nor U2261 (N_2261,N_2081,N_2010);
nand U2262 (N_2262,N_2106,N_2056);
xnor U2263 (N_2263,N_2100,N_2147);
xor U2264 (N_2264,N_2024,N_2173);
or U2265 (N_2265,N_2166,N_2182);
and U2266 (N_2266,N_2151,N_2080);
nor U2267 (N_2267,N_2053,N_2124);
and U2268 (N_2268,N_2001,N_2121);
xnor U2269 (N_2269,N_2028,N_2155);
or U2270 (N_2270,N_2183,N_2088);
and U2271 (N_2271,N_2031,N_2198);
nor U2272 (N_2272,N_2175,N_2160);
and U2273 (N_2273,N_2109,N_2092);
and U2274 (N_2274,N_2162,N_2188);
xnor U2275 (N_2275,N_2074,N_2089);
or U2276 (N_2276,N_2108,N_2082);
xnor U2277 (N_2277,N_2163,N_2158);
and U2278 (N_2278,N_2135,N_2032);
and U2279 (N_2279,N_2035,N_2107);
nand U2280 (N_2280,N_2165,N_2189);
nand U2281 (N_2281,N_2117,N_2063);
xnor U2282 (N_2282,N_2119,N_2142);
nand U2283 (N_2283,N_2076,N_2058);
xor U2284 (N_2284,N_2070,N_2018);
xnor U2285 (N_2285,N_2177,N_2050);
nand U2286 (N_2286,N_2016,N_2137);
and U2287 (N_2287,N_2005,N_2061);
xnor U2288 (N_2288,N_2174,N_2180);
or U2289 (N_2289,N_2044,N_2101);
nor U2290 (N_2290,N_2161,N_2066);
nor U2291 (N_2291,N_2057,N_2164);
and U2292 (N_2292,N_2007,N_2156);
and U2293 (N_2293,N_2168,N_2011);
and U2294 (N_2294,N_2059,N_2132);
nor U2295 (N_2295,N_2086,N_2049);
nor U2296 (N_2296,N_2083,N_2148);
and U2297 (N_2297,N_2042,N_2055);
nand U2298 (N_2298,N_2130,N_2136);
nor U2299 (N_2299,N_2071,N_2069);
and U2300 (N_2300,N_2122,N_2053);
nor U2301 (N_2301,N_2016,N_2099);
or U2302 (N_2302,N_2120,N_2032);
nand U2303 (N_2303,N_2167,N_2017);
nand U2304 (N_2304,N_2101,N_2172);
xnor U2305 (N_2305,N_2115,N_2170);
nand U2306 (N_2306,N_2091,N_2098);
nand U2307 (N_2307,N_2128,N_2073);
nor U2308 (N_2308,N_2027,N_2014);
and U2309 (N_2309,N_2112,N_2145);
nor U2310 (N_2310,N_2167,N_2112);
and U2311 (N_2311,N_2049,N_2172);
nand U2312 (N_2312,N_2175,N_2025);
nor U2313 (N_2313,N_2173,N_2029);
or U2314 (N_2314,N_2102,N_2017);
xnor U2315 (N_2315,N_2143,N_2088);
and U2316 (N_2316,N_2044,N_2012);
nor U2317 (N_2317,N_2161,N_2080);
or U2318 (N_2318,N_2123,N_2105);
nand U2319 (N_2319,N_2141,N_2187);
and U2320 (N_2320,N_2023,N_2140);
xor U2321 (N_2321,N_2164,N_2114);
and U2322 (N_2322,N_2023,N_2181);
nor U2323 (N_2323,N_2024,N_2062);
and U2324 (N_2324,N_2171,N_2170);
nand U2325 (N_2325,N_2008,N_2136);
nand U2326 (N_2326,N_2042,N_2003);
xor U2327 (N_2327,N_2195,N_2094);
nor U2328 (N_2328,N_2046,N_2187);
xor U2329 (N_2329,N_2127,N_2153);
nand U2330 (N_2330,N_2024,N_2055);
nor U2331 (N_2331,N_2057,N_2030);
nor U2332 (N_2332,N_2164,N_2193);
and U2333 (N_2333,N_2155,N_2174);
xnor U2334 (N_2334,N_2109,N_2091);
or U2335 (N_2335,N_2018,N_2001);
nor U2336 (N_2336,N_2171,N_2150);
and U2337 (N_2337,N_2177,N_2039);
and U2338 (N_2338,N_2178,N_2136);
or U2339 (N_2339,N_2027,N_2184);
or U2340 (N_2340,N_2079,N_2112);
nor U2341 (N_2341,N_2098,N_2018);
and U2342 (N_2342,N_2055,N_2035);
xnor U2343 (N_2343,N_2136,N_2106);
nand U2344 (N_2344,N_2089,N_2192);
nor U2345 (N_2345,N_2107,N_2120);
and U2346 (N_2346,N_2043,N_2027);
nor U2347 (N_2347,N_2083,N_2014);
and U2348 (N_2348,N_2108,N_2153);
and U2349 (N_2349,N_2092,N_2172);
or U2350 (N_2350,N_2103,N_2122);
nand U2351 (N_2351,N_2069,N_2060);
nor U2352 (N_2352,N_2055,N_2090);
xor U2353 (N_2353,N_2095,N_2026);
xnor U2354 (N_2354,N_2085,N_2001);
xnor U2355 (N_2355,N_2057,N_2185);
xnor U2356 (N_2356,N_2047,N_2165);
or U2357 (N_2357,N_2127,N_2033);
and U2358 (N_2358,N_2121,N_2131);
xor U2359 (N_2359,N_2156,N_2053);
nand U2360 (N_2360,N_2176,N_2059);
nand U2361 (N_2361,N_2180,N_2003);
nand U2362 (N_2362,N_2154,N_2150);
xnor U2363 (N_2363,N_2077,N_2083);
nor U2364 (N_2364,N_2057,N_2097);
or U2365 (N_2365,N_2176,N_2181);
nand U2366 (N_2366,N_2038,N_2109);
or U2367 (N_2367,N_2102,N_2046);
xor U2368 (N_2368,N_2058,N_2175);
nor U2369 (N_2369,N_2006,N_2190);
nor U2370 (N_2370,N_2136,N_2015);
xnor U2371 (N_2371,N_2125,N_2054);
or U2372 (N_2372,N_2062,N_2114);
nand U2373 (N_2373,N_2053,N_2128);
nand U2374 (N_2374,N_2078,N_2197);
or U2375 (N_2375,N_2045,N_2031);
nor U2376 (N_2376,N_2055,N_2153);
and U2377 (N_2377,N_2105,N_2155);
or U2378 (N_2378,N_2161,N_2046);
nor U2379 (N_2379,N_2018,N_2111);
nor U2380 (N_2380,N_2142,N_2029);
nor U2381 (N_2381,N_2150,N_2046);
nand U2382 (N_2382,N_2090,N_2010);
nand U2383 (N_2383,N_2077,N_2137);
nor U2384 (N_2384,N_2084,N_2005);
nand U2385 (N_2385,N_2183,N_2136);
nand U2386 (N_2386,N_2054,N_2009);
xnor U2387 (N_2387,N_2178,N_2081);
or U2388 (N_2388,N_2059,N_2102);
nand U2389 (N_2389,N_2059,N_2172);
or U2390 (N_2390,N_2070,N_2159);
xnor U2391 (N_2391,N_2121,N_2137);
xor U2392 (N_2392,N_2152,N_2185);
nand U2393 (N_2393,N_2080,N_2046);
nor U2394 (N_2394,N_2161,N_2101);
nand U2395 (N_2395,N_2086,N_2029);
or U2396 (N_2396,N_2139,N_2054);
xnor U2397 (N_2397,N_2139,N_2070);
or U2398 (N_2398,N_2017,N_2158);
xor U2399 (N_2399,N_2151,N_2030);
nor U2400 (N_2400,N_2291,N_2353);
nor U2401 (N_2401,N_2399,N_2221);
or U2402 (N_2402,N_2352,N_2285);
or U2403 (N_2403,N_2335,N_2385);
nor U2404 (N_2404,N_2307,N_2290);
xor U2405 (N_2405,N_2276,N_2311);
xor U2406 (N_2406,N_2280,N_2329);
xor U2407 (N_2407,N_2318,N_2238);
nor U2408 (N_2408,N_2343,N_2295);
xor U2409 (N_2409,N_2231,N_2259);
or U2410 (N_2410,N_2227,N_2356);
and U2411 (N_2411,N_2225,N_2355);
and U2412 (N_2412,N_2371,N_2250);
xor U2413 (N_2413,N_2289,N_2233);
and U2414 (N_2414,N_2330,N_2296);
and U2415 (N_2415,N_2292,N_2388);
or U2416 (N_2416,N_2218,N_2387);
nand U2417 (N_2417,N_2297,N_2316);
and U2418 (N_2418,N_2398,N_2306);
nor U2419 (N_2419,N_2246,N_2300);
and U2420 (N_2420,N_2337,N_2308);
nand U2421 (N_2421,N_2245,N_2315);
or U2422 (N_2422,N_2380,N_2286);
xor U2423 (N_2423,N_2362,N_2274);
nand U2424 (N_2424,N_2224,N_2229);
nor U2425 (N_2425,N_2322,N_2202);
nor U2426 (N_2426,N_2217,N_2317);
xnor U2427 (N_2427,N_2288,N_2379);
and U2428 (N_2428,N_2234,N_2277);
xnor U2429 (N_2429,N_2204,N_2220);
and U2430 (N_2430,N_2369,N_2340);
nor U2431 (N_2431,N_2255,N_2214);
and U2432 (N_2432,N_2282,N_2293);
xor U2433 (N_2433,N_2346,N_2382);
nor U2434 (N_2434,N_2391,N_2240);
nor U2435 (N_2435,N_2358,N_2305);
and U2436 (N_2436,N_2310,N_2396);
nand U2437 (N_2437,N_2203,N_2251);
nand U2438 (N_2438,N_2215,N_2390);
xor U2439 (N_2439,N_2332,N_2339);
or U2440 (N_2440,N_2256,N_2260);
or U2441 (N_2441,N_2367,N_2205);
xor U2442 (N_2442,N_2287,N_2360);
and U2443 (N_2443,N_2394,N_2375);
or U2444 (N_2444,N_2264,N_2275);
xor U2445 (N_2445,N_2248,N_2208);
and U2446 (N_2446,N_2323,N_2365);
and U2447 (N_2447,N_2266,N_2303);
nand U2448 (N_2448,N_2376,N_2359);
xnor U2449 (N_2449,N_2232,N_2269);
nor U2450 (N_2450,N_2368,N_2386);
nor U2451 (N_2451,N_2347,N_2393);
or U2452 (N_2452,N_2209,N_2370);
nor U2453 (N_2453,N_2263,N_2210);
and U2454 (N_2454,N_2216,N_2324);
nor U2455 (N_2455,N_2331,N_2254);
nand U2456 (N_2456,N_2281,N_2392);
nand U2457 (N_2457,N_2261,N_2364);
nand U2458 (N_2458,N_2273,N_2294);
xor U2459 (N_2459,N_2201,N_2314);
and U2460 (N_2460,N_2284,N_2241);
nand U2461 (N_2461,N_2350,N_2239);
xor U2462 (N_2462,N_2207,N_2372);
xnor U2463 (N_2463,N_2351,N_2298);
nor U2464 (N_2464,N_2278,N_2279);
nand U2465 (N_2465,N_2389,N_2328);
xnor U2466 (N_2466,N_2338,N_2252);
xnor U2467 (N_2467,N_2253,N_2336);
xnor U2468 (N_2468,N_2223,N_2377);
or U2469 (N_2469,N_2244,N_2272);
nand U2470 (N_2470,N_2247,N_2395);
nand U2471 (N_2471,N_2258,N_2299);
or U2472 (N_2472,N_2257,N_2378);
nand U2473 (N_2473,N_2366,N_2230);
nor U2474 (N_2474,N_2267,N_2304);
nor U2475 (N_2475,N_2262,N_2236);
nor U2476 (N_2476,N_2243,N_2219);
nand U2477 (N_2477,N_2271,N_2349);
and U2478 (N_2478,N_2342,N_2222);
nor U2479 (N_2479,N_2320,N_2235);
and U2480 (N_2480,N_2348,N_2334);
nand U2481 (N_2481,N_2374,N_2361);
or U2482 (N_2482,N_2200,N_2249);
xor U2483 (N_2483,N_2344,N_2268);
and U2484 (N_2484,N_2265,N_2345);
nor U2485 (N_2485,N_2206,N_2363);
nand U2486 (N_2486,N_2270,N_2326);
or U2487 (N_2487,N_2397,N_2384);
nand U2488 (N_2488,N_2325,N_2321);
nand U2489 (N_2489,N_2213,N_2228);
xor U2490 (N_2490,N_2301,N_2211);
xnor U2491 (N_2491,N_2226,N_2309);
nor U2492 (N_2492,N_2373,N_2354);
or U2493 (N_2493,N_2242,N_2357);
xor U2494 (N_2494,N_2302,N_2341);
or U2495 (N_2495,N_2212,N_2237);
and U2496 (N_2496,N_2283,N_2313);
nor U2497 (N_2497,N_2327,N_2312);
or U2498 (N_2498,N_2319,N_2383);
xor U2499 (N_2499,N_2333,N_2381);
or U2500 (N_2500,N_2300,N_2276);
and U2501 (N_2501,N_2208,N_2291);
or U2502 (N_2502,N_2358,N_2357);
and U2503 (N_2503,N_2378,N_2236);
nand U2504 (N_2504,N_2234,N_2359);
or U2505 (N_2505,N_2330,N_2354);
xor U2506 (N_2506,N_2263,N_2385);
nor U2507 (N_2507,N_2277,N_2266);
nor U2508 (N_2508,N_2358,N_2267);
and U2509 (N_2509,N_2333,N_2358);
and U2510 (N_2510,N_2378,N_2318);
nand U2511 (N_2511,N_2252,N_2329);
nor U2512 (N_2512,N_2321,N_2201);
and U2513 (N_2513,N_2384,N_2371);
nand U2514 (N_2514,N_2318,N_2213);
and U2515 (N_2515,N_2395,N_2260);
xnor U2516 (N_2516,N_2317,N_2228);
nand U2517 (N_2517,N_2304,N_2264);
nand U2518 (N_2518,N_2369,N_2268);
nor U2519 (N_2519,N_2332,N_2335);
nor U2520 (N_2520,N_2235,N_2321);
nand U2521 (N_2521,N_2238,N_2206);
nor U2522 (N_2522,N_2252,N_2242);
nand U2523 (N_2523,N_2303,N_2321);
xnor U2524 (N_2524,N_2395,N_2239);
and U2525 (N_2525,N_2244,N_2346);
or U2526 (N_2526,N_2277,N_2206);
nand U2527 (N_2527,N_2250,N_2376);
xnor U2528 (N_2528,N_2290,N_2361);
nand U2529 (N_2529,N_2374,N_2313);
nor U2530 (N_2530,N_2246,N_2291);
and U2531 (N_2531,N_2222,N_2247);
and U2532 (N_2532,N_2226,N_2356);
and U2533 (N_2533,N_2392,N_2249);
or U2534 (N_2534,N_2211,N_2309);
nand U2535 (N_2535,N_2317,N_2235);
xnor U2536 (N_2536,N_2206,N_2205);
and U2537 (N_2537,N_2367,N_2249);
nand U2538 (N_2538,N_2297,N_2389);
nand U2539 (N_2539,N_2290,N_2215);
or U2540 (N_2540,N_2277,N_2264);
nor U2541 (N_2541,N_2228,N_2376);
xor U2542 (N_2542,N_2201,N_2399);
nor U2543 (N_2543,N_2297,N_2295);
and U2544 (N_2544,N_2246,N_2239);
or U2545 (N_2545,N_2268,N_2334);
xnor U2546 (N_2546,N_2361,N_2210);
xnor U2547 (N_2547,N_2294,N_2343);
and U2548 (N_2548,N_2219,N_2256);
and U2549 (N_2549,N_2231,N_2257);
nand U2550 (N_2550,N_2233,N_2257);
xnor U2551 (N_2551,N_2362,N_2366);
xor U2552 (N_2552,N_2280,N_2370);
xor U2553 (N_2553,N_2349,N_2293);
or U2554 (N_2554,N_2296,N_2336);
or U2555 (N_2555,N_2254,N_2389);
nand U2556 (N_2556,N_2241,N_2206);
xor U2557 (N_2557,N_2255,N_2352);
nor U2558 (N_2558,N_2372,N_2310);
nor U2559 (N_2559,N_2392,N_2336);
xnor U2560 (N_2560,N_2309,N_2312);
xnor U2561 (N_2561,N_2364,N_2385);
or U2562 (N_2562,N_2225,N_2345);
nor U2563 (N_2563,N_2224,N_2255);
nand U2564 (N_2564,N_2378,N_2395);
xor U2565 (N_2565,N_2207,N_2275);
and U2566 (N_2566,N_2286,N_2336);
and U2567 (N_2567,N_2387,N_2343);
nand U2568 (N_2568,N_2315,N_2308);
or U2569 (N_2569,N_2345,N_2254);
nand U2570 (N_2570,N_2361,N_2254);
nand U2571 (N_2571,N_2333,N_2344);
nand U2572 (N_2572,N_2369,N_2230);
xnor U2573 (N_2573,N_2340,N_2302);
or U2574 (N_2574,N_2234,N_2301);
nor U2575 (N_2575,N_2361,N_2368);
nand U2576 (N_2576,N_2314,N_2361);
or U2577 (N_2577,N_2384,N_2202);
nor U2578 (N_2578,N_2335,N_2379);
nor U2579 (N_2579,N_2378,N_2297);
xor U2580 (N_2580,N_2353,N_2380);
and U2581 (N_2581,N_2331,N_2322);
nand U2582 (N_2582,N_2347,N_2203);
or U2583 (N_2583,N_2398,N_2357);
xnor U2584 (N_2584,N_2361,N_2335);
and U2585 (N_2585,N_2288,N_2247);
nand U2586 (N_2586,N_2279,N_2201);
xor U2587 (N_2587,N_2366,N_2257);
and U2588 (N_2588,N_2343,N_2325);
and U2589 (N_2589,N_2351,N_2270);
and U2590 (N_2590,N_2294,N_2235);
nand U2591 (N_2591,N_2267,N_2343);
and U2592 (N_2592,N_2245,N_2371);
and U2593 (N_2593,N_2344,N_2231);
xnor U2594 (N_2594,N_2349,N_2212);
or U2595 (N_2595,N_2225,N_2271);
and U2596 (N_2596,N_2258,N_2260);
and U2597 (N_2597,N_2262,N_2284);
xnor U2598 (N_2598,N_2244,N_2371);
and U2599 (N_2599,N_2226,N_2264);
xor U2600 (N_2600,N_2569,N_2402);
xor U2601 (N_2601,N_2422,N_2455);
nor U2602 (N_2602,N_2410,N_2409);
or U2603 (N_2603,N_2585,N_2574);
or U2604 (N_2604,N_2513,N_2519);
nand U2605 (N_2605,N_2440,N_2419);
nand U2606 (N_2606,N_2545,N_2454);
nor U2607 (N_2607,N_2507,N_2515);
xnor U2608 (N_2608,N_2433,N_2496);
xnor U2609 (N_2609,N_2497,N_2491);
and U2610 (N_2610,N_2473,N_2528);
and U2611 (N_2611,N_2427,N_2561);
nand U2612 (N_2612,N_2598,N_2508);
nor U2613 (N_2613,N_2577,N_2538);
or U2614 (N_2614,N_2488,N_2583);
and U2615 (N_2615,N_2543,N_2570);
nand U2616 (N_2616,N_2460,N_2542);
xnor U2617 (N_2617,N_2479,N_2533);
nor U2618 (N_2618,N_2465,N_2550);
nand U2619 (N_2619,N_2459,N_2596);
nand U2620 (N_2620,N_2551,N_2430);
or U2621 (N_2621,N_2527,N_2595);
nand U2622 (N_2622,N_2597,N_2504);
nand U2623 (N_2623,N_2462,N_2571);
nor U2624 (N_2624,N_2444,N_2493);
nand U2625 (N_2625,N_2498,N_2431);
nand U2626 (N_2626,N_2437,N_2441);
nor U2627 (N_2627,N_2403,N_2565);
nor U2628 (N_2628,N_2576,N_2438);
or U2629 (N_2629,N_2499,N_2526);
and U2630 (N_2630,N_2572,N_2552);
and U2631 (N_2631,N_2503,N_2413);
nand U2632 (N_2632,N_2566,N_2476);
nor U2633 (N_2633,N_2531,N_2467);
nor U2634 (N_2634,N_2408,N_2546);
xor U2635 (N_2635,N_2406,N_2429);
nor U2636 (N_2636,N_2450,N_2478);
or U2637 (N_2637,N_2564,N_2494);
or U2638 (N_2638,N_2401,N_2553);
xnor U2639 (N_2639,N_2523,N_2540);
nand U2640 (N_2640,N_2575,N_2547);
and U2641 (N_2641,N_2416,N_2525);
nor U2642 (N_2642,N_2421,N_2567);
and U2643 (N_2643,N_2581,N_2502);
nand U2644 (N_2644,N_2529,N_2517);
and U2645 (N_2645,N_2534,N_2555);
nand U2646 (N_2646,N_2461,N_2489);
or U2647 (N_2647,N_2510,N_2469);
nor U2648 (N_2648,N_2474,N_2592);
xor U2649 (N_2649,N_2434,N_2480);
xnor U2650 (N_2650,N_2580,N_2447);
nor U2651 (N_2651,N_2557,N_2400);
nor U2652 (N_2652,N_2405,N_2544);
xnor U2653 (N_2653,N_2562,N_2559);
nor U2654 (N_2654,N_2456,N_2448);
nor U2655 (N_2655,N_2500,N_2594);
xor U2656 (N_2656,N_2495,N_2404);
xor U2657 (N_2657,N_2483,N_2536);
and U2658 (N_2658,N_2591,N_2463);
and U2659 (N_2659,N_2418,N_2482);
nor U2660 (N_2660,N_2541,N_2518);
xnor U2661 (N_2661,N_2587,N_2573);
nand U2662 (N_2662,N_2490,N_2520);
xor U2663 (N_2663,N_2516,N_2423);
nor U2664 (N_2664,N_2442,N_2466);
or U2665 (N_2665,N_2586,N_2578);
nand U2666 (N_2666,N_2558,N_2506);
xnor U2667 (N_2667,N_2445,N_2439);
xor U2668 (N_2668,N_2548,N_2472);
nor U2669 (N_2669,N_2484,N_2537);
or U2670 (N_2670,N_2556,N_2424);
nor U2671 (N_2671,N_2511,N_2464);
xor U2672 (N_2672,N_2446,N_2492);
nor U2673 (N_2673,N_2563,N_2414);
or U2674 (N_2674,N_2486,N_2425);
nand U2675 (N_2675,N_2449,N_2443);
nor U2676 (N_2676,N_2452,N_2530);
nor U2677 (N_2677,N_2432,N_2549);
or U2678 (N_2678,N_2568,N_2477);
and U2679 (N_2679,N_2589,N_2599);
xnor U2680 (N_2680,N_2417,N_2487);
or U2681 (N_2681,N_2453,N_2522);
nand U2682 (N_2682,N_2512,N_2539);
and U2683 (N_2683,N_2524,N_2588);
nor U2684 (N_2684,N_2593,N_2435);
nand U2685 (N_2685,N_2535,N_2590);
nor U2686 (N_2686,N_2436,N_2582);
or U2687 (N_2687,N_2415,N_2501);
nor U2688 (N_2688,N_2584,N_2407);
nand U2689 (N_2689,N_2560,N_2509);
xnor U2690 (N_2690,N_2505,N_2412);
xor U2691 (N_2691,N_2521,N_2451);
nor U2692 (N_2692,N_2471,N_2420);
xor U2693 (N_2693,N_2485,N_2470);
or U2694 (N_2694,N_2468,N_2475);
nor U2695 (N_2695,N_2426,N_2428);
xnor U2696 (N_2696,N_2481,N_2411);
nor U2697 (N_2697,N_2458,N_2579);
xnor U2698 (N_2698,N_2532,N_2554);
and U2699 (N_2699,N_2514,N_2457);
nor U2700 (N_2700,N_2597,N_2554);
and U2701 (N_2701,N_2599,N_2469);
nand U2702 (N_2702,N_2595,N_2479);
nor U2703 (N_2703,N_2408,N_2499);
nand U2704 (N_2704,N_2559,N_2514);
and U2705 (N_2705,N_2539,N_2567);
nor U2706 (N_2706,N_2482,N_2423);
or U2707 (N_2707,N_2559,N_2586);
nor U2708 (N_2708,N_2506,N_2510);
nor U2709 (N_2709,N_2488,N_2402);
nor U2710 (N_2710,N_2480,N_2462);
or U2711 (N_2711,N_2552,N_2438);
and U2712 (N_2712,N_2590,N_2573);
xor U2713 (N_2713,N_2452,N_2524);
and U2714 (N_2714,N_2546,N_2423);
nand U2715 (N_2715,N_2570,N_2587);
nor U2716 (N_2716,N_2402,N_2452);
nor U2717 (N_2717,N_2416,N_2421);
nand U2718 (N_2718,N_2562,N_2405);
nand U2719 (N_2719,N_2597,N_2595);
nor U2720 (N_2720,N_2588,N_2530);
and U2721 (N_2721,N_2575,N_2503);
nor U2722 (N_2722,N_2558,N_2427);
xor U2723 (N_2723,N_2574,N_2427);
xnor U2724 (N_2724,N_2429,N_2508);
and U2725 (N_2725,N_2486,N_2448);
or U2726 (N_2726,N_2534,N_2578);
or U2727 (N_2727,N_2572,N_2592);
nand U2728 (N_2728,N_2522,N_2558);
and U2729 (N_2729,N_2407,N_2488);
xor U2730 (N_2730,N_2551,N_2543);
nor U2731 (N_2731,N_2405,N_2437);
and U2732 (N_2732,N_2529,N_2535);
nor U2733 (N_2733,N_2449,N_2577);
or U2734 (N_2734,N_2581,N_2488);
and U2735 (N_2735,N_2407,N_2400);
xnor U2736 (N_2736,N_2503,N_2406);
xor U2737 (N_2737,N_2555,N_2592);
nor U2738 (N_2738,N_2598,N_2500);
nand U2739 (N_2739,N_2576,N_2567);
nor U2740 (N_2740,N_2476,N_2597);
and U2741 (N_2741,N_2486,N_2506);
xor U2742 (N_2742,N_2535,N_2490);
nor U2743 (N_2743,N_2414,N_2559);
or U2744 (N_2744,N_2535,N_2557);
nand U2745 (N_2745,N_2505,N_2413);
xnor U2746 (N_2746,N_2429,N_2438);
or U2747 (N_2747,N_2403,N_2560);
xor U2748 (N_2748,N_2506,N_2552);
or U2749 (N_2749,N_2424,N_2443);
xnor U2750 (N_2750,N_2554,N_2424);
nor U2751 (N_2751,N_2564,N_2583);
and U2752 (N_2752,N_2548,N_2563);
nor U2753 (N_2753,N_2514,N_2543);
nand U2754 (N_2754,N_2467,N_2496);
or U2755 (N_2755,N_2410,N_2568);
xor U2756 (N_2756,N_2554,N_2596);
or U2757 (N_2757,N_2558,N_2560);
nor U2758 (N_2758,N_2400,N_2517);
nor U2759 (N_2759,N_2494,N_2515);
xnor U2760 (N_2760,N_2529,N_2462);
and U2761 (N_2761,N_2415,N_2570);
xnor U2762 (N_2762,N_2427,N_2422);
nor U2763 (N_2763,N_2475,N_2524);
or U2764 (N_2764,N_2502,N_2410);
or U2765 (N_2765,N_2475,N_2503);
xor U2766 (N_2766,N_2581,N_2553);
and U2767 (N_2767,N_2513,N_2447);
nand U2768 (N_2768,N_2558,N_2426);
and U2769 (N_2769,N_2501,N_2541);
nand U2770 (N_2770,N_2461,N_2431);
nand U2771 (N_2771,N_2586,N_2447);
or U2772 (N_2772,N_2445,N_2437);
nor U2773 (N_2773,N_2493,N_2514);
or U2774 (N_2774,N_2461,N_2575);
or U2775 (N_2775,N_2582,N_2487);
and U2776 (N_2776,N_2553,N_2491);
nor U2777 (N_2777,N_2536,N_2527);
nand U2778 (N_2778,N_2564,N_2535);
and U2779 (N_2779,N_2466,N_2511);
nand U2780 (N_2780,N_2465,N_2538);
nand U2781 (N_2781,N_2581,N_2461);
or U2782 (N_2782,N_2420,N_2489);
or U2783 (N_2783,N_2431,N_2483);
xor U2784 (N_2784,N_2425,N_2469);
nand U2785 (N_2785,N_2503,N_2534);
and U2786 (N_2786,N_2421,N_2594);
xor U2787 (N_2787,N_2433,N_2536);
xor U2788 (N_2788,N_2516,N_2417);
or U2789 (N_2789,N_2452,N_2406);
nor U2790 (N_2790,N_2498,N_2591);
xnor U2791 (N_2791,N_2451,N_2546);
xor U2792 (N_2792,N_2525,N_2427);
and U2793 (N_2793,N_2402,N_2458);
and U2794 (N_2794,N_2475,N_2579);
nand U2795 (N_2795,N_2423,N_2594);
nand U2796 (N_2796,N_2557,N_2485);
or U2797 (N_2797,N_2568,N_2522);
xnor U2798 (N_2798,N_2410,N_2564);
xor U2799 (N_2799,N_2415,N_2432);
and U2800 (N_2800,N_2697,N_2620);
nor U2801 (N_2801,N_2645,N_2778);
or U2802 (N_2802,N_2707,N_2703);
nor U2803 (N_2803,N_2619,N_2750);
or U2804 (N_2804,N_2797,N_2781);
nor U2805 (N_2805,N_2798,N_2749);
nand U2806 (N_2806,N_2603,N_2639);
or U2807 (N_2807,N_2660,N_2640);
nor U2808 (N_2808,N_2729,N_2723);
and U2809 (N_2809,N_2653,N_2602);
and U2810 (N_2810,N_2732,N_2679);
and U2811 (N_2811,N_2699,N_2644);
nor U2812 (N_2812,N_2740,N_2706);
and U2813 (N_2813,N_2783,N_2688);
and U2814 (N_2814,N_2685,N_2704);
or U2815 (N_2815,N_2659,N_2700);
nor U2816 (N_2816,N_2759,N_2677);
nand U2817 (N_2817,N_2730,N_2634);
xor U2818 (N_2818,N_2655,N_2651);
nor U2819 (N_2819,N_2607,N_2770);
nor U2820 (N_2820,N_2686,N_2771);
and U2821 (N_2821,N_2622,N_2752);
xnor U2822 (N_2822,N_2772,N_2613);
or U2823 (N_2823,N_2769,N_2625);
or U2824 (N_2824,N_2755,N_2667);
xor U2825 (N_2825,N_2689,N_2608);
xor U2826 (N_2826,N_2629,N_2780);
xor U2827 (N_2827,N_2606,N_2741);
nand U2828 (N_2828,N_2726,N_2669);
or U2829 (N_2829,N_2784,N_2616);
xnor U2830 (N_2830,N_2761,N_2692);
nand U2831 (N_2831,N_2674,N_2649);
or U2832 (N_2832,N_2657,N_2654);
xnor U2833 (N_2833,N_2736,N_2615);
or U2834 (N_2834,N_2714,N_2733);
xor U2835 (N_2835,N_2662,N_2623);
nand U2836 (N_2836,N_2696,N_2748);
nor U2837 (N_2837,N_2746,N_2643);
nor U2838 (N_2838,N_2787,N_2676);
nor U2839 (N_2839,N_2624,N_2682);
and U2840 (N_2840,N_2604,N_2789);
or U2841 (N_2841,N_2790,N_2713);
and U2842 (N_2842,N_2742,N_2743);
and U2843 (N_2843,N_2665,N_2648);
nor U2844 (N_2844,N_2701,N_2747);
nor U2845 (N_2845,N_2767,N_2627);
or U2846 (N_2846,N_2652,N_2765);
and U2847 (N_2847,N_2666,N_2776);
or U2848 (N_2848,N_2661,N_2728);
or U2849 (N_2849,N_2788,N_2664);
and U2850 (N_2850,N_2785,N_2690);
xnor U2851 (N_2851,N_2756,N_2668);
or U2852 (N_2852,N_2610,N_2710);
xor U2853 (N_2853,N_2601,N_2777);
and U2854 (N_2854,N_2646,N_2737);
and U2855 (N_2855,N_2628,N_2631);
nand U2856 (N_2856,N_2751,N_2632);
nand U2857 (N_2857,N_2609,N_2734);
nand U2858 (N_2858,N_2708,N_2678);
nand U2859 (N_2859,N_2712,N_2744);
or U2860 (N_2860,N_2672,N_2757);
nor U2861 (N_2861,N_2630,N_2638);
nor U2862 (N_2862,N_2663,N_2735);
nand U2863 (N_2863,N_2731,N_2719);
and U2864 (N_2864,N_2725,N_2611);
nand U2865 (N_2865,N_2766,N_2775);
nor U2866 (N_2866,N_2758,N_2702);
xnor U2867 (N_2867,N_2779,N_2684);
nand U2868 (N_2868,N_2683,N_2739);
xnor U2869 (N_2869,N_2791,N_2637);
xor U2870 (N_2870,N_2760,N_2642);
nor U2871 (N_2871,N_2773,N_2786);
nand U2872 (N_2872,N_2799,N_2633);
nand U2873 (N_2873,N_2794,N_2796);
nor U2874 (N_2874,N_2754,N_2641);
or U2875 (N_2875,N_2720,N_2636);
nand U2876 (N_2876,N_2715,N_2671);
nor U2877 (N_2877,N_2738,N_2753);
and U2878 (N_2878,N_2763,N_2670);
nand U2879 (N_2879,N_2681,N_2656);
xor U2880 (N_2880,N_2617,N_2721);
nor U2881 (N_2881,N_2768,N_2614);
nor U2882 (N_2882,N_2793,N_2722);
nor U2883 (N_2883,N_2698,N_2717);
or U2884 (N_2884,N_2605,N_2673);
or U2885 (N_2885,N_2618,N_2716);
and U2886 (N_2886,N_2774,N_2795);
and U2887 (N_2887,N_2680,N_2705);
or U2888 (N_2888,N_2724,N_2694);
and U2889 (N_2889,N_2792,N_2675);
nor U2890 (N_2890,N_2687,N_2693);
and U2891 (N_2891,N_2626,N_2635);
nand U2892 (N_2892,N_2718,N_2745);
and U2893 (N_2893,N_2600,N_2709);
nand U2894 (N_2894,N_2621,N_2691);
xor U2895 (N_2895,N_2658,N_2762);
xnor U2896 (N_2896,N_2764,N_2647);
or U2897 (N_2897,N_2711,N_2612);
and U2898 (N_2898,N_2695,N_2782);
xnor U2899 (N_2899,N_2650,N_2727);
and U2900 (N_2900,N_2758,N_2730);
nand U2901 (N_2901,N_2790,N_2697);
nor U2902 (N_2902,N_2698,N_2666);
xor U2903 (N_2903,N_2714,N_2792);
or U2904 (N_2904,N_2645,N_2624);
nor U2905 (N_2905,N_2767,N_2744);
nand U2906 (N_2906,N_2721,N_2722);
xor U2907 (N_2907,N_2733,N_2784);
and U2908 (N_2908,N_2738,N_2662);
xnor U2909 (N_2909,N_2710,N_2688);
xor U2910 (N_2910,N_2619,N_2672);
xnor U2911 (N_2911,N_2751,N_2675);
and U2912 (N_2912,N_2600,N_2691);
nor U2913 (N_2913,N_2727,N_2612);
xnor U2914 (N_2914,N_2621,N_2778);
nor U2915 (N_2915,N_2668,N_2714);
nand U2916 (N_2916,N_2706,N_2690);
nand U2917 (N_2917,N_2674,N_2729);
nand U2918 (N_2918,N_2788,N_2676);
and U2919 (N_2919,N_2734,N_2754);
nand U2920 (N_2920,N_2772,N_2627);
xor U2921 (N_2921,N_2624,N_2683);
xor U2922 (N_2922,N_2742,N_2747);
or U2923 (N_2923,N_2683,N_2723);
and U2924 (N_2924,N_2632,N_2629);
xor U2925 (N_2925,N_2734,N_2689);
nand U2926 (N_2926,N_2670,N_2710);
or U2927 (N_2927,N_2641,N_2688);
xnor U2928 (N_2928,N_2653,N_2629);
nor U2929 (N_2929,N_2696,N_2767);
or U2930 (N_2930,N_2601,N_2780);
nand U2931 (N_2931,N_2600,N_2605);
nand U2932 (N_2932,N_2749,N_2716);
and U2933 (N_2933,N_2741,N_2789);
nor U2934 (N_2934,N_2627,N_2705);
nor U2935 (N_2935,N_2704,N_2775);
nand U2936 (N_2936,N_2611,N_2616);
xor U2937 (N_2937,N_2715,N_2626);
nand U2938 (N_2938,N_2736,N_2766);
nand U2939 (N_2939,N_2684,N_2704);
nor U2940 (N_2940,N_2644,N_2795);
nor U2941 (N_2941,N_2637,N_2789);
and U2942 (N_2942,N_2760,N_2723);
xnor U2943 (N_2943,N_2629,N_2720);
nand U2944 (N_2944,N_2749,N_2795);
xnor U2945 (N_2945,N_2772,N_2615);
nand U2946 (N_2946,N_2767,N_2676);
and U2947 (N_2947,N_2777,N_2638);
or U2948 (N_2948,N_2776,N_2604);
or U2949 (N_2949,N_2675,N_2776);
and U2950 (N_2950,N_2721,N_2601);
or U2951 (N_2951,N_2653,N_2799);
nand U2952 (N_2952,N_2617,N_2682);
or U2953 (N_2953,N_2640,N_2623);
nor U2954 (N_2954,N_2669,N_2661);
xnor U2955 (N_2955,N_2784,N_2698);
and U2956 (N_2956,N_2616,N_2607);
xor U2957 (N_2957,N_2721,N_2647);
nand U2958 (N_2958,N_2711,N_2776);
nor U2959 (N_2959,N_2755,N_2688);
or U2960 (N_2960,N_2699,N_2701);
nand U2961 (N_2961,N_2733,N_2676);
or U2962 (N_2962,N_2757,N_2707);
xnor U2963 (N_2963,N_2682,N_2797);
and U2964 (N_2964,N_2765,N_2714);
nor U2965 (N_2965,N_2671,N_2713);
nor U2966 (N_2966,N_2668,N_2789);
and U2967 (N_2967,N_2634,N_2708);
nand U2968 (N_2968,N_2718,N_2603);
nor U2969 (N_2969,N_2692,N_2765);
nand U2970 (N_2970,N_2736,N_2630);
and U2971 (N_2971,N_2700,N_2761);
nor U2972 (N_2972,N_2652,N_2602);
or U2973 (N_2973,N_2623,N_2742);
nand U2974 (N_2974,N_2669,N_2609);
nor U2975 (N_2975,N_2794,N_2614);
or U2976 (N_2976,N_2776,N_2714);
and U2977 (N_2977,N_2635,N_2649);
xor U2978 (N_2978,N_2717,N_2624);
nand U2979 (N_2979,N_2611,N_2652);
xor U2980 (N_2980,N_2676,N_2664);
xor U2981 (N_2981,N_2740,N_2773);
xnor U2982 (N_2982,N_2660,N_2669);
nor U2983 (N_2983,N_2731,N_2627);
or U2984 (N_2984,N_2722,N_2685);
and U2985 (N_2985,N_2683,N_2657);
nor U2986 (N_2986,N_2787,N_2655);
nor U2987 (N_2987,N_2763,N_2690);
or U2988 (N_2988,N_2652,N_2692);
or U2989 (N_2989,N_2796,N_2629);
nor U2990 (N_2990,N_2683,N_2764);
or U2991 (N_2991,N_2620,N_2704);
and U2992 (N_2992,N_2732,N_2609);
nor U2993 (N_2993,N_2725,N_2786);
and U2994 (N_2994,N_2683,N_2702);
nand U2995 (N_2995,N_2695,N_2662);
or U2996 (N_2996,N_2734,N_2634);
nor U2997 (N_2997,N_2690,N_2618);
nand U2998 (N_2998,N_2660,N_2780);
xor U2999 (N_2999,N_2779,N_2740);
and U3000 (N_3000,N_2862,N_2847);
or U3001 (N_3001,N_2982,N_2864);
xnor U3002 (N_3002,N_2907,N_2899);
nor U3003 (N_3003,N_2969,N_2916);
or U3004 (N_3004,N_2889,N_2875);
nor U3005 (N_3005,N_2854,N_2941);
nor U3006 (N_3006,N_2930,N_2966);
nor U3007 (N_3007,N_2936,N_2809);
nor U3008 (N_3008,N_2852,N_2984);
nand U3009 (N_3009,N_2857,N_2812);
nor U3010 (N_3010,N_2995,N_2900);
or U3011 (N_3011,N_2841,N_2863);
and U3012 (N_3012,N_2992,N_2981);
nand U3013 (N_3013,N_2877,N_2979);
nor U3014 (N_3014,N_2903,N_2914);
or U3015 (N_3015,N_2853,N_2950);
and U3016 (N_3016,N_2834,N_2839);
xor U3017 (N_3017,N_2837,N_2865);
or U3018 (N_3018,N_2893,N_2949);
xnor U3019 (N_3019,N_2895,N_2927);
xor U3020 (N_3020,N_2817,N_2998);
nand U3021 (N_3021,N_2832,N_2994);
xnor U3022 (N_3022,N_2858,N_2810);
xor U3023 (N_3023,N_2974,N_2882);
nor U3024 (N_3024,N_2823,N_2821);
and U3025 (N_3025,N_2831,N_2924);
and U3026 (N_3026,N_2801,N_2824);
nand U3027 (N_3027,N_2961,N_2991);
and U3028 (N_3028,N_2946,N_2956);
or U3029 (N_3029,N_2990,N_2978);
nand U3030 (N_3030,N_2897,N_2977);
xnor U3031 (N_3031,N_2973,N_2892);
or U3032 (N_3032,N_2953,N_2993);
or U3033 (N_3033,N_2828,N_2942);
nor U3034 (N_3034,N_2806,N_2879);
nand U3035 (N_3035,N_2909,N_2846);
or U3036 (N_3036,N_2898,N_2962);
or U3037 (N_3037,N_2968,N_2957);
nor U3038 (N_3038,N_2825,N_2922);
xor U3039 (N_3039,N_2869,N_2970);
xnor U3040 (N_3040,N_2840,N_2844);
nand U3041 (N_3041,N_2999,N_2965);
or U3042 (N_3042,N_2880,N_2881);
nand U3043 (N_3043,N_2934,N_2971);
nor U3044 (N_3044,N_2835,N_2803);
and U3045 (N_3045,N_2931,N_2805);
nand U3046 (N_3046,N_2985,N_2887);
xor U3047 (N_3047,N_2883,N_2925);
nand U3048 (N_3048,N_2986,N_2976);
xor U3049 (N_3049,N_2822,N_2983);
and U3050 (N_3050,N_2943,N_2814);
xor U3051 (N_3051,N_2911,N_2912);
xnor U3052 (N_3052,N_2947,N_2815);
or U3053 (N_3053,N_2891,N_2819);
nand U3054 (N_3054,N_2827,N_2804);
xor U3055 (N_3055,N_2873,N_2800);
or U3056 (N_3056,N_2894,N_2807);
nor U3057 (N_3057,N_2921,N_2820);
xor U3058 (N_3058,N_2871,N_2996);
xnor U3059 (N_3059,N_2902,N_2851);
or U3060 (N_3060,N_2888,N_2808);
and U3061 (N_3061,N_2843,N_2967);
xor U3062 (N_3062,N_2945,N_2849);
and U3063 (N_3063,N_2811,N_2972);
xnor U3064 (N_3064,N_2884,N_2935);
nor U3065 (N_3065,N_2955,N_2818);
xor U3066 (N_3066,N_2830,N_2833);
or U3067 (N_3067,N_2829,N_2944);
and U3068 (N_3068,N_2954,N_2845);
or U3069 (N_3069,N_2826,N_2868);
and U3070 (N_3070,N_2980,N_2908);
and U3071 (N_3071,N_2987,N_2948);
nand U3072 (N_3072,N_2813,N_2910);
or U3073 (N_3073,N_2913,N_2964);
xor U3074 (N_3074,N_2896,N_2940);
and U3075 (N_3075,N_2861,N_2850);
and U3076 (N_3076,N_2885,N_2918);
and U3077 (N_3077,N_2917,N_2960);
and U3078 (N_3078,N_2859,N_2848);
or U3079 (N_3079,N_2929,N_2951);
nor U3080 (N_3080,N_2802,N_2963);
or U3081 (N_3081,N_2952,N_2938);
nor U3082 (N_3082,N_2906,N_2939);
or U3083 (N_3083,N_2915,N_2923);
nor U3084 (N_3084,N_2997,N_2933);
xnor U3085 (N_3085,N_2816,N_2860);
nor U3086 (N_3086,N_2904,N_2937);
xnor U3087 (N_3087,N_2872,N_2928);
xnor U3088 (N_3088,N_2901,N_2920);
xnor U3089 (N_3089,N_2842,N_2874);
nand U3090 (N_3090,N_2856,N_2836);
xor U3091 (N_3091,N_2919,N_2905);
nor U3092 (N_3092,N_2878,N_2975);
nand U3093 (N_3093,N_2959,N_2989);
or U3094 (N_3094,N_2932,N_2958);
nand U3095 (N_3095,N_2876,N_2838);
and U3096 (N_3096,N_2926,N_2890);
xnor U3097 (N_3097,N_2886,N_2867);
xor U3098 (N_3098,N_2870,N_2988);
nand U3099 (N_3099,N_2866,N_2855);
nand U3100 (N_3100,N_2824,N_2931);
and U3101 (N_3101,N_2903,N_2806);
and U3102 (N_3102,N_2803,N_2944);
nor U3103 (N_3103,N_2902,N_2907);
and U3104 (N_3104,N_2821,N_2978);
xor U3105 (N_3105,N_2922,N_2832);
or U3106 (N_3106,N_2865,N_2905);
or U3107 (N_3107,N_2859,N_2815);
and U3108 (N_3108,N_2826,N_2805);
xor U3109 (N_3109,N_2935,N_2995);
or U3110 (N_3110,N_2997,N_2923);
or U3111 (N_3111,N_2875,N_2979);
xnor U3112 (N_3112,N_2895,N_2922);
nand U3113 (N_3113,N_2917,N_2943);
and U3114 (N_3114,N_2929,N_2849);
nor U3115 (N_3115,N_2924,N_2992);
nand U3116 (N_3116,N_2862,N_2879);
xnor U3117 (N_3117,N_2979,N_2923);
and U3118 (N_3118,N_2868,N_2853);
and U3119 (N_3119,N_2870,N_2849);
nor U3120 (N_3120,N_2843,N_2821);
nand U3121 (N_3121,N_2853,N_2838);
or U3122 (N_3122,N_2958,N_2957);
xor U3123 (N_3123,N_2800,N_2870);
xnor U3124 (N_3124,N_2923,N_2870);
or U3125 (N_3125,N_2831,N_2835);
xnor U3126 (N_3126,N_2921,N_2804);
nor U3127 (N_3127,N_2961,N_2901);
nand U3128 (N_3128,N_2947,N_2922);
and U3129 (N_3129,N_2818,N_2959);
and U3130 (N_3130,N_2803,N_2914);
xnor U3131 (N_3131,N_2831,N_2832);
or U3132 (N_3132,N_2950,N_2829);
xor U3133 (N_3133,N_2942,N_2995);
xor U3134 (N_3134,N_2907,N_2965);
nand U3135 (N_3135,N_2927,N_2891);
nor U3136 (N_3136,N_2803,N_2856);
and U3137 (N_3137,N_2849,N_2999);
nand U3138 (N_3138,N_2995,N_2845);
or U3139 (N_3139,N_2948,N_2829);
or U3140 (N_3140,N_2868,N_2967);
xnor U3141 (N_3141,N_2918,N_2984);
or U3142 (N_3142,N_2925,N_2870);
nor U3143 (N_3143,N_2937,N_2967);
nand U3144 (N_3144,N_2818,N_2923);
or U3145 (N_3145,N_2899,N_2807);
nor U3146 (N_3146,N_2999,N_2923);
xnor U3147 (N_3147,N_2891,N_2898);
xor U3148 (N_3148,N_2958,N_2896);
nand U3149 (N_3149,N_2820,N_2917);
nand U3150 (N_3150,N_2819,N_2826);
nand U3151 (N_3151,N_2907,N_2838);
or U3152 (N_3152,N_2963,N_2810);
xor U3153 (N_3153,N_2816,N_2899);
nand U3154 (N_3154,N_2946,N_2906);
and U3155 (N_3155,N_2979,N_2950);
xnor U3156 (N_3156,N_2873,N_2899);
or U3157 (N_3157,N_2997,N_2971);
xnor U3158 (N_3158,N_2891,N_2822);
xor U3159 (N_3159,N_2856,N_2913);
and U3160 (N_3160,N_2851,N_2837);
nand U3161 (N_3161,N_2829,N_2919);
and U3162 (N_3162,N_2842,N_2891);
or U3163 (N_3163,N_2845,N_2959);
xor U3164 (N_3164,N_2980,N_2949);
xnor U3165 (N_3165,N_2925,N_2988);
and U3166 (N_3166,N_2812,N_2803);
xor U3167 (N_3167,N_2982,N_2827);
xor U3168 (N_3168,N_2830,N_2902);
and U3169 (N_3169,N_2849,N_2820);
nand U3170 (N_3170,N_2886,N_2865);
xnor U3171 (N_3171,N_2801,N_2880);
and U3172 (N_3172,N_2977,N_2835);
or U3173 (N_3173,N_2955,N_2904);
nand U3174 (N_3174,N_2834,N_2918);
or U3175 (N_3175,N_2908,N_2892);
nand U3176 (N_3176,N_2974,N_2993);
xnor U3177 (N_3177,N_2887,N_2804);
or U3178 (N_3178,N_2811,N_2884);
nor U3179 (N_3179,N_2910,N_2939);
xor U3180 (N_3180,N_2967,N_2997);
nand U3181 (N_3181,N_2893,N_2969);
nor U3182 (N_3182,N_2853,N_2922);
xnor U3183 (N_3183,N_2924,N_2995);
and U3184 (N_3184,N_2845,N_2946);
nor U3185 (N_3185,N_2879,N_2946);
xnor U3186 (N_3186,N_2863,N_2908);
nor U3187 (N_3187,N_2853,N_2921);
and U3188 (N_3188,N_2904,N_2918);
nor U3189 (N_3189,N_2858,N_2812);
nor U3190 (N_3190,N_2823,N_2955);
or U3191 (N_3191,N_2821,N_2828);
and U3192 (N_3192,N_2960,N_2901);
xor U3193 (N_3193,N_2869,N_2905);
xnor U3194 (N_3194,N_2958,N_2951);
or U3195 (N_3195,N_2865,N_2964);
nand U3196 (N_3196,N_2890,N_2931);
nand U3197 (N_3197,N_2834,N_2931);
xor U3198 (N_3198,N_2993,N_2969);
and U3199 (N_3199,N_2830,N_2952);
or U3200 (N_3200,N_3118,N_3113);
xor U3201 (N_3201,N_3196,N_3128);
xnor U3202 (N_3202,N_3062,N_3142);
xnor U3203 (N_3203,N_3042,N_3159);
nor U3204 (N_3204,N_3052,N_3071);
or U3205 (N_3205,N_3134,N_3067);
and U3206 (N_3206,N_3168,N_3189);
nor U3207 (N_3207,N_3083,N_3172);
nand U3208 (N_3208,N_3043,N_3064);
xnor U3209 (N_3209,N_3199,N_3176);
and U3210 (N_3210,N_3038,N_3029);
nor U3211 (N_3211,N_3000,N_3102);
nor U3212 (N_3212,N_3175,N_3161);
xor U3213 (N_3213,N_3023,N_3088);
nand U3214 (N_3214,N_3021,N_3166);
nor U3215 (N_3215,N_3077,N_3003);
nand U3216 (N_3216,N_3146,N_3024);
or U3217 (N_3217,N_3135,N_3066);
and U3218 (N_3218,N_3080,N_3092);
and U3219 (N_3219,N_3170,N_3155);
nand U3220 (N_3220,N_3111,N_3049);
nor U3221 (N_3221,N_3085,N_3075);
or U3222 (N_3222,N_3163,N_3122);
or U3223 (N_3223,N_3059,N_3120);
nor U3224 (N_3224,N_3013,N_3078);
or U3225 (N_3225,N_3103,N_3138);
nand U3226 (N_3226,N_3002,N_3136);
and U3227 (N_3227,N_3018,N_3139);
and U3228 (N_3228,N_3114,N_3150);
xnor U3229 (N_3229,N_3022,N_3145);
nand U3230 (N_3230,N_3179,N_3006);
nor U3231 (N_3231,N_3094,N_3091);
nor U3232 (N_3232,N_3053,N_3044);
nand U3233 (N_3233,N_3182,N_3147);
or U3234 (N_3234,N_3143,N_3194);
or U3235 (N_3235,N_3164,N_3084);
or U3236 (N_3236,N_3187,N_3151);
nor U3237 (N_3237,N_3169,N_3031);
xor U3238 (N_3238,N_3190,N_3156);
nand U3239 (N_3239,N_3070,N_3109);
nand U3240 (N_3240,N_3068,N_3061);
nor U3241 (N_3241,N_3121,N_3093);
or U3242 (N_3242,N_3015,N_3106);
or U3243 (N_3243,N_3027,N_3055);
xor U3244 (N_3244,N_3115,N_3101);
nand U3245 (N_3245,N_3017,N_3158);
or U3246 (N_3246,N_3045,N_3020);
nor U3247 (N_3247,N_3099,N_3195);
nand U3248 (N_3248,N_3047,N_3191);
or U3249 (N_3249,N_3127,N_3110);
xnor U3250 (N_3250,N_3041,N_3048);
nor U3251 (N_3251,N_3119,N_3073);
nand U3252 (N_3252,N_3181,N_3039);
or U3253 (N_3253,N_3098,N_3050);
xnor U3254 (N_3254,N_3025,N_3171);
xnor U3255 (N_3255,N_3090,N_3037);
xnor U3256 (N_3256,N_3019,N_3148);
or U3257 (N_3257,N_3034,N_3058);
nand U3258 (N_3258,N_3131,N_3167);
or U3259 (N_3259,N_3186,N_3086);
xnor U3260 (N_3260,N_3087,N_3079);
nand U3261 (N_3261,N_3112,N_3157);
xor U3262 (N_3262,N_3005,N_3116);
or U3263 (N_3263,N_3007,N_3117);
nand U3264 (N_3264,N_3160,N_3030);
and U3265 (N_3265,N_3174,N_3123);
or U3266 (N_3266,N_3100,N_3065);
nor U3267 (N_3267,N_3096,N_3081);
nand U3268 (N_3268,N_3082,N_3057);
and U3269 (N_3269,N_3153,N_3033);
and U3270 (N_3270,N_3028,N_3183);
nor U3271 (N_3271,N_3012,N_3076);
nand U3272 (N_3272,N_3188,N_3063);
xor U3273 (N_3273,N_3180,N_3072);
nor U3274 (N_3274,N_3152,N_3124);
or U3275 (N_3275,N_3011,N_3089);
nand U3276 (N_3276,N_3016,N_3040);
nor U3277 (N_3277,N_3173,N_3095);
nand U3278 (N_3278,N_3074,N_3130);
nor U3279 (N_3279,N_3032,N_3008);
xor U3280 (N_3280,N_3178,N_3144);
and U3281 (N_3281,N_3184,N_3141);
nor U3282 (N_3282,N_3009,N_3140);
or U3283 (N_3283,N_3132,N_3197);
nand U3284 (N_3284,N_3108,N_3104);
and U3285 (N_3285,N_3105,N_3154);
nor U3286 (N_3286,N_3193,N_3046);
nor U3287 (N_3287,N_3001,N_3026);
xor U3288 (N_3288,N_3097,N_3014);
and U3289 (N_3289,N_3069,N_3056);
or U3290 (N_3290,N_3149,N_3060);
or U3291 (N_3291,N_3137,N_3133);
xor U3292 (N_3292,N_3107,N_3010);
or U3293 (N_3293,N_3051,N_3035);
xor U3294 (N_3294,N_3165,N_3125);
nor U3295 (N_3295,N_3177,N_3162);
nand U3296 (N_3296,N_3126,N_3054);
and U3297 (N_3297,N_3185,N_3192);
nor U3298 (N_3298,N_3004,N_3036);
xnor U3299 (N_3299,N_3129,N_3198);
and U3300 (N_3300,N_3006,N_3050);
xnor U3301 (N_3301,N_3045,N_3115);
xnor U3302 (N_3302,N_3005,N_3044);
xnor U3303 (N_3303,N_3157,N_3171);
or U3304 (N_3304,N_3067,N_3193);
xnor U3305 (N_3305,N_3038,N_3009);
and U3306 (N_3306,N_3188,N_3141);
xnor U3307 (N_3307,N_3084,N_3199);
nand U3308 (N_3308,N_3020,N_3196);
and U3309 (N_3309,N_3087,N_3195);
nor U3310 (N_3310,N_3005,N_3084);
nor U3311 (N_3311,N_3046,N_3144);
and U3312 (N_3312,N_3025,N_3132);
xnor U3313 (N_3313,N_3032,N_3079);
or U3314 (N_3314,N_3100,N_3036);
or U3315 (N_3315,N_3184,N_3114);
nor U3316 (N_3316,N_3150,N_3070);
or U3317 (N_3317,N_3063,N_3154);
xnor U3318 (N_3318,N_3061,N_3132);
xor U3319 (N_3319,N_3140,N_3132);
and U3320 (N_3320,N_3077,N_3107);
nor U3321 (N_3321,N_3063,N_3155);
nand U3322 (N_3322,N_3099,N_3165);
nand U3323 (N_3323,N_3186,N_3085);
and U3324 (N_3324,N_3146,N_3084);
nor U3325 (N_3325,N_3051,N_3144);
nand U3326 (N_3326,N_3100,N_3150);
nor U3327 (N_3327,N_3107,N_3012);
nand U3328 (N_3328,N_3127,N_3089);
or U3329 (N_3329,N_3062,N_3053);
and U3330 (N_3330,N_3059,N_3195);
nor U3331 (N_3331,N_3152,N_3084);
nor U3332 (N_3332,N_3073,N_3019);
xor U3333 (N_3333,N_3112,N_3146);
or U3334 (N_3334,N_3107,N_3184);
and U3335 (N_3335,N_3197,N_3039);
or U3336 (N_3336,N_3099,N_3158);
nor U3337 (N_3337,N_3083,N_3038);
xnor U3338 (N_3338,N_3001,N_3164);
and U3339 (N_3339,N_3014,N_3126);
xor U3340 (N_3340,N_3126,N_3068);
or U3341 (N_3341,N_3117,N_3011);
and U3342 (N_3342,N_3162,N_3103);
nor U3343 (N_3343,N_3175,N_3060);
and U3344 (N_3344,N_3046,N_3082);
nand U3345 (N_3345,N_3044,N_3022);
xnor U3346 (N_3346,N_3169,N_3154);
nand U3347 (N_3347,N_3059,N_3165);
or U3348 (N_3348,N_3115,N_3137);
and U3349 (N_3349,N_3109,N_3066);
or U3350 (N_3350,N_3106,N_3131);
or U3351 (N_3351,N_3166,N_3108);
nor U3352 (N_3352,N_3162,N_3148);
and U3353 (N_3353,N_3100,N_3051);
and U3354 (N_3354,N_3184,N_3051);
or U3355 (N_3355,N_3137,N_3152);
and U3356 (N_3356,N_3165,N_3148);
or U3357 (N_3357,N_3136,N_3063);
xnor U3358 (N_3358,N_3064,N_3118);
or U3359 (N_3359,N_3126,N_3038);
and U3360 (N_3360,N_3061,N_3198);
and U3361 (N_3361,N_3073,N_3148);
xnor U3362 (N_3362,N_3009,N_3118);
or U3363 (N_3363,N_3105,N_3074);
nand U3364 (N_3364,N_3103,N_3196);
nand U3365 (N_3365,N_3071,N_3191);
or U3366 (N_3366,N_3152,N_3191);
nand U3367 (N_3367,N_3180,N_3011);
or U3368 (N_3368,N_3173,N_3099);
nand U3369 (N_3369,N_3038,N_3078);
or U3370 (N_3370,N_3033,N_3090);
nor U3371 (N_3371,N_3155,N_3120);
nand U3372 (N_3372,N_3133,N_3047);
or U3373 (N_3373,N_3065,N_3119);
nand U3374 (N_3374,N_3193,N_3168);
nor U3375 (N_3375,N_3069,N_3007);
and U3376 (N_3376,N_3107,N_3147);
nand U3377 (N_3377,N_3116,N_3110);
and U3378 (N_3378,N_3173,N_3102);
xor U3379 (N_3379,N_3096,N_3055);
nor U3380 (N_3380,N_3011,N_3058);
nor U3381 (N_3381,N_3184,N_3059);
or U3382 (N_3382,N_3018,N_3193);
nand U3383 (N_3383,N_3085,N_3153);
nand U3384 (N_3384,N_3126,N_3063);
xnor U3385 (N_3385,N_3196,N_3028);
xor U3386 (N_3386,N_3141,N_3154);
or U3387 (N_3387,N_3146,N_3171);
and U3388 (N_3388,N_3172,N_3192);
nand U3389 (N_3389,N_3173,N_3020);
or U3390 (N_3390,N_3143,N_3153);
xor U3391 (N_3391,N_3189,N_3103);
and U3392 (N_3392,N_3021,N_3004);
nor U3393 (N_3393,N_3172,N_3035);
or U3394 (N_3394,N_3047,N_3144);
xnor U3395 (N_3395,N_3155,N_3050);
xor U3396 (N_3396,N_3070,N_3069);
and U3397 (N_3397,N_3094,N_3098);
or U3398 (N_3398,N_3074,N_3187);
xnor U3399 (N_3399,N_3073,N_3129);
xnor U3400 (N_3400,N_3286,N_3315);
nand U3401 (N_3401,N_3269,N_3242);
or U3402 (N_3402,N_3399,N_3338);
nor U3403 (N_3403,N_3296,N_3310);
and U3404 (N_3404,N_3256,N_3380);
and U3405 (N_3405,N_3249,N_3347);
and U3406 (N_3406,N_3308,N_3307);
xor U3407 (N_3407,N_3370,N_3209);
or U3408 (N_3408,N_3212,N_3213);
or U3409 (N_3409,N_3265,N_3351);
nand U3410 (N_3410,N_3288,N_3263);
nand U3411 (N_3411,N_3394,N_3301);
and U3412 (N_3412,N_3348,N_3357);
or U3413 (N_3413,N_3246,N_3396);
xnor U3414 (N_3414,N_3368,N_3322);
and U3415 (N_3415,N_3208,N_3233);
xor U3416 (N_3416,N_3339,N_3312);
and U3417 (N_3417,N_3287,N_3290);
xor U3418 (N_3418,N_3217,N_3354);
xnor U3419 (N_3419,N_3214,N_3275);
xnor U3420 (N_3420,N_3273,N_3359);
nor U3421 (N_3421,N_3237,N_3364);
and U3422 (N_3422,N_3373,N_3341);
and U3423 (N_3423,N_3393,N_3205);
or U3424 (N_3424,N_3227,N_3344);
and U3425 (N_3425,N_3385,N_3231);
or U3426 (N_3426,N_3384,N_3277);
and U3427 (N_3427,N_3362,N_3320);
xnor U3428 (N_3428,N_3335,N_3395);
or U3429 (N_3429,N_3306,N_3252);
nand U3430 (N_3430,N_3352,N_3244);
nand U3431 (N_3431,N_3309,N_3271);
xor U3432 (N_3432,N_3215,N_3374);
nand U3433 (N_3433,N_3378,N_3391);
and U3434 (N_3434,N_3363,N_3200);
and U3435 (N_3435,N_3302,N_3334);
and U3436 (N_3436,N_3280,N_3257);
or U3437 (N_3437,N_3366,N_3201);
xnor U3438 (N_3438,N_3248,N_3336);
and U3439 (N_3439,N_3379,N_3323);
xor U3440 (N_3440,N_3311,N_3260);
xnor U3441 (N_3441,N_3207,N_3204);
nand U3442 (N_3442,N_3369,N_3324);
and U3443 (N_3443,N_3304,N_3313);
xor U3444 (N_3444,N_3397,N_3356);
xnor U3445 (N_3445,N_3232,N_3388);
or U3446 (N_3446,N_3264,N_3314);
nand U3447 (N_3447,N_3222,N_3330);
or U3448 (N_3448,N_3353,N_3235);
xor U3449 (N_3449,N_3345,N_3291);
nand U3450 (N_3450,N_3333,N_3389);
nor U3451 (N_3451,N_3375,N_3343);
nand U3452 (N_3452,N_3272,N_3262);
or U3453 (N_3453,N_3350,N_3250);
xnor U3454 (N_3454,N_3387,N_3298);
nand U3455 (N_3455,N_3266,N_3274);
xnor U3456 (N_3456,N_3225,N_3285);
or U3457 (N_3457,N_3216,N_3376);
and U3458 (N_3458,N_3261,N_3211);
xor U3459 (N_3459,N_3329,N_3293);
and U3460 (N_3460,N_3342,N_3316);
nor U3461 (N_3461,N_3331,N_3245);
and U3462 (N_3462,N_3294,N_3360);
nand U3463 (N_3463,N_3367,N_3327);
and U3464 (N_3464,N_3390,N_3337);
nor U3465 (N_3465,N_3238,N_3254);
and U3466 (N_3466,N_3382,N_3383);
xor U3467 (N_3467,N_3258,N_3267);
and U3468 (N_3468,N_3318,N_3228);
nand U3469 (N_3469,N_3317,N_3203);
or U3470 (N_3470,N_3305,N_3239);
nor U3471 (N_3471,N_3281,N_3319);
xnor U3472 (N_3472,N_3240,N_3210);
and U3473 (N_3473,N_3372,N_3295);
nand U3474 (N_3474,N_3303,N_3278);
nor U3475 (N_3475,N_3300,N_3355);
xnor U3476 (N_3476,N_3365,N_3224);
xnor U3477 (N_3477,N_3268,N_3234);
or U3478 (N_3478,N_3292,N_3381);
nand U3479 (N_3479,N_3230,N_3202);
xnor U3480 (N_3480,N_3223,N_3229);
and U3481 (N_3481,N_3251,N_3346);
and U3482 (N_3482,N_3253,N_3332);
nor U3483 (N_3483,N_3386,N_3326);
nand U3484 (N_3484,N_3398,N_3371);
and U3485 (N_3485,N_3321,N_3297);
or U3486 (N_3486,N_3236,N_3325);
nand U3487 (N_3487,N_3279,N_3241);
or U3488 (N_3488,N_3218,N_3340);
nor U3489 (N_3489,N_3358,N_3206);
xnor U3490 (N_3490,N_3377,N_3349);
nor U3491 (N_3491,N_3221,N_3247);
and U3492 (N_3492,N_3284,N_3289);
nor U3493 (N_3493,N_3243,N_3361);
xnor U3494 (N_3494,N_3283,N_3328);
nor U3495 (N_3495,N_3276,N_3270);
nor U3496 (N_3496,N_3255,N_3219);
xor U3497 (N_3497,N_3220,N_3392);
nand U3498 (N_3498,N_3299,N_3259);
and U3499 (N_3499,N_3226,N_3282);
or U3500 (N_3500,N_3345,N_3344);
and U3501 (N_3501,N_3245,N_3309);
xnor U3502 (N_3502,N_3235,N_3286);
and U3503 (N_3503,N_3376,N_3379);
or U3504 (N_3504,N_3277,N_3264);
or U3505 (N_3505,N_3349,N_3339);
or U3506 (N_3506,N_3371,N_3240);
nor U3507 (N_3507,N_3274,N_3350);
and U3508 (N_3508,N_3217,N_3346);
or U3509 (N_3509,N_3342,N_3257);
or U3510 (N_3510,N_3206,N_3393);
or U3511 (N_3511,N_3260,N_3246);
or U3512 (N_3512,N_3258,N_3282);
or U3513 (N_3513,N_3220,N_3329);
and U3514 (N_3514,N_3390,N_3316);
nand U3515 (N_3515,N_3352,N_3267);
nand U3516 (N_3516,N_3341,N_3309);
or U3517 (N_3517,N_3235,N_3292);
nand U3518 (N_3518,N_3258,N_3200);
and U3519 (N_3519,N_3358,N_3309);
nor U3520 (N_3520,N_3328,N_3269);
nand U3521 (N_3521,N_3381,N_3303);
nand U3522 (N_3522,N_3238,N_3291);
nor U3523 (N_3523,N_3240,N_3258);
or U3524 (N_3524,N_3293,N_3305);
xnor U3525 (N_3525,N_3369,N_3309);
nor U3526 (N_3526,N_3259,N_3380);
xnor U3527 (N_3527,N_3251,N_3351);
nor U3528 (N_3528,N_3236,N_3289);
xnor U3529 (N_3529,N_3296,N_3230);
nor U3530 (N_3530,N_3389,N_3356);
and U3531 (N_3531,N_3209,N_3389);
nand U3532 (N_3532,N_3231,N_3283);
and U3533 (N_3533,N_3248,N_3358);
nor U3534 (N_3534,N_3250,N_3295);
nand U3535 (N_3535,N_3395,N_3330);
xnor U3536 (N_3536,N_3338,N_3351);
or U3537 (N_3537,N_3223,N_3241);
xor U3538 (N_3538,N_3279,N_3301);
nand U3539 (N_3539,N_3343,N_3304);
and U3540 (N_3540,N_3371,N_3354);
and U3541 (N_3541,N_3291,N_3381);
or U3542 (N_3542,N_3393,N_3328);
nand U3543 (N_3543,N_3233,N_3207);
or U3544 (N_3544,N_3255,N_3261);
nor U3545 (N_3545,N_3337,N_3286);
nand U3546 (N_3546,N_3398,N_3271);
nand U3547 (N_3547,N_3253,N_3255);
or U3548 (N_3548,N_3243,N_3213);
or U3549 (N_3549,N_3292,N_3361);
xnor U3550 (N_3550,N_3382,N_3204);
xor U3551 (N_3551,N_3227,N_3266);
xnor U3552 (N_3552,N_3209,N_3335);
and U3553 (N_3553,N_3393,N_3371);
nand U3554 (N_3554,N_3308,N_3360);
nand U3555 (N_3555,N_3219,N_3201);
nand U3556 (N_3556,N_3226,N_3394);
or U3557 (N_3557,N_3202,N_3258);
nand U3558 (N_3558,N_3358,N_3267);
xnor U3559 (N_3559,N_3242,N_3280);
and U3560 (N_3560,N_3389,N_3235);
nor U3561 (N_3561,N_3231,N_3343);
and U3562 (N_3562,N_3209,N_3374);
nor U3563 (N_3563,N_3320,N_3339);
xor U3564 (N_3564,N_3336,N_3294);
or U3565 (N_3565,N_3229,N_3205);
and U3566 (N_3566,N_3283,N_3269);
or U3567 (N_3567,N_3200,N_3356);
and U3568 (N_3568,N_3295,N_3270);
nor U3569 (N_3569,N_3356,N_3281);
and U3570 (N_3570,N_3288,N_3353);
or U3571 (N_3571,N_3372,N_3291);
xnor U3572 (N_3572,N_3286,N_3375);
and U3573 (N_3573,N_3364,N_3304);
nor U3574 (N_3574,N_3362,N_3281);
xor U3575 (N_3575,N_3286,N_3277);
xor U3576 (N_3576,N_3381,N_3398);
and U3577 (N_3577,N_3352,N_3280);
or U3578 (N_3578,N_3312,N_3259);
nand U3579 (N_3579,N_3226,N_3272);
and U3580 (N_3580,N_3325,N_3374);
nand U3581 (N_3581,N_3393,N_3311);
nand U3582 (N_3582,N_3272,N_3386);
nand U3583 (N_3583,N_3315,N_3363);
nor U3584 (N_3584,N_3235,N_3349);
or U3585 (N_3585,N_3227,N_3385);
nor U3586 (N_3586,N_3259,N_3382);
nor U3587 (N_3587,N_3316,N_3221);
and U3588 (N_3588,N_3277,N_3205);
nor U3589 (N_3589,N_3362,N_3213);
nand U3590 (N_3590,N_3362,N_3325);
xnor U3591 (N_3591,N_3215,N_3217);
nand U3592 (N_3592,N_3381,N_3250);
xnor U3593 (N_3593,N_3242,N_3344);
xnor U3594 (N_3594,N_3244,N_3315);
nand U3595 (N_3595,N_3240,N_3205);
nor U3596 (N_3596,N_3266,N_3390);
xor U3597 (N_3597,N_3277,N_3351);
or U3598 (N_3598,N_3311,N_3357);
or U3599 (N_3599,N_3321,N_3244);
and U3600 (N_3600,N_3424,N_3469);
or U3601 (N_3601,N_3530,N_3406);
nand U3602 (N_3602,N_3589,N_3426);
xor U3603 (N_3603,N_3546,N_3563);
nor U3604 (N_3604,N_3445,N_3591);
or U3605 (N_3605,N_3483,N_3521);
nand U3606 (N_3606,N_3553,N_3438);
nor U3607 (N_3607,N_3537,N_3423);
or U3608 (N_3608,N_3544,N_3517);
xor U3609 (N_3609,N_3543,N_3568);
xor U3610 (N_3610,N_3479,N_3585);
xnor U3611 (N_3611,N_3562,N_3583);
nor U3612 (N_3612,N_3566,N_3598);
nor U3613 (N_3613,N_3453,N_3448);
nand U3614 (N_3614,N_3579,N_3417);
and U3615 (N_3615,N_3405,N_3597);
or U3616 (N_3616,N_3470,N_3547);
and U3617 (N_3617,N_3408,N_3475);
nand U3618 (N_3618,N_3581,N_3454);
or U3619 (N_3619,N_3441,N_3430);
nand U3620 (N_3620,N_3588,N_3552);
or U3621 (N_3621,N_3526,N_3594);
xnor U3622 (N_3622,N_3497,N_3542);
and U3623 (N_3623,N_3564,N_3422);
or U3624 (N_3624,N_3490,N_3431);
and U3625 (N_3625,N_3559,N_3550);
nand U3626 (N_3626,N_3502,N_3403);
or U3627 (N_3627,N_3481,N_3493);
or U3628 (N_3628,N_3414,N_3458);
nor U3629 (N_3629,N_3539,N_3501);
and U3630 (N_3630,N_3512,N_3467);
nor U3631 (N_3631,N_3465,N_3450);
and U3632 (N_3632,N_3531,N_3511);
nor U3633 (N_3633,N_3404,N_3482);
and U3634 (N_3634,N_3571,N_3477);
nor U3635 (N_3635,N_3527,N_3570);
nand U3636 (N_3636,N_3491,N_3495);
nand U3637 (N_3637,N_3519,N_3525);
or U3638 (N_3638,N_3560,N_3508);
or U3639 (N_3639,N_3593,N_3449);
and U3640 (N_3640,N_3576,N_3522);
or U3641 (N_3641,N_3435,N_3433);
nand U3642 (N_3642,N_3509,N_3541);
xnor U3643 (N_3643,N_3504,N_3462);
nor U3644 (N_3644,N_3557,N_3599);
or U3645 (N_3645,N_3584,N_3529);
nand U3646 (N_3646,N_3567,N_3487);
nor U3647 (N_3647,N_3503,N_3443);
nand U3648 (N_3648,N_3460,N_3586);
nand U3649 (N_3649,N_3459,N_3569);
xor U3650 (N_3650,N_3551,N_3442);
or U3651 (N_3651,N_3484,N_3596);
and U3652 (N_3652,N_3420,N_3440);
or U3653 (N_3653,N_3498,N_3480);
nand U3654 (N_3654,N_3510,N_3488);
nor U3655 (N_3655,N_3437,N_3486);
and U3656 (N_3656,N_3520,N_3523);
or U3657 (N_3657,N_3573,N_3436);
nor U3658 (N_3658,N_3565,N_3500);
nor U3659 (N_3659,N_3411,N_3474);
nand U3660 (N_3660,N_3413,N_3492);
nand U3661 (N_3661,N_3540,N_3515);
nand U3662 (N_3662,N_3548,N_3428);
xor U3663 (N_3663,N_3402,N_3507);
nand U3664 (N_3664,N_3572,N_3578);
nor U3665 (N_3665,N_3561,N_3485);
nand U3666 (N_3666,N_3466,N_3472);
and U3667 (N_3667,N_3577,N_3451);
nand U3668 (N_3668,N_3429,N_3452);
nand U3669 (N_3669,N_3457,N_3401);
xnor U3670 (N_3670,N_3456,N_3524);
or U3671 (N_3671,N_3421,N_3532);
nand U3672 (N_3672,N_3463,N_3516);
and U3673 (N_3673,N_3439,N_3549);
xnor U3674 (N_3674,N_3494,N_3415);
nand U3675 (N_3675,N_3446,N_3535);
nor U3676 (N_3676,N_3434,N_3528);
nand U3677 (N_3677,N_3574,N_3410);
and U3678 (N_3678,N_3538,N_3400);
nor U3679 (N_3679,N_3556,N_3505);
and U3680 (N_3680,N_3447,N_3514);
and U3681 (N_3681,N_3444,N_3473);
xor U3682 (N_3682,N_3464,N_3555);
or U3683 (N_3683,N_3427,N_3582);
or U3684 (N_3684,N_3496,N_3506);
xnor U3685 (N_3685,N_3558,N_3412);
or U3686 (N_3686,N_3418,N_3536);
xnor U3687 (N_3687,N_3409,N_3432);
nand U3688 (N_3688,N_3461,N_3476);
nor U3689 (N_3689,N_3554,N_3590);
xnor U3690 (N_3690,N_3489,N_3534);
xnor U3691 (N_3691,N_3575,N_3587);
nand U3692 (N_3692,N_3419,N_3545);
nor U3693 (N_3693,N_3468,N_3580);
nor U3694 (N_3694,N_3455,N_3425);
nor U3695 (N_3695,N_3407,N_3513);
nand U3696 (N_3696,N_3471,N_3592);
or U3697 (N_3697,N_3416,N_3478);
xor U3698 (N_3698,N_3533,N_3499);
nand U3699 (N_3699,N_3518,N_3595);
nand U3700 (N_3700,N_3462,N_3511);
xor U3701 (N_3701,N_3467,N_3432);
or U3702 (N_3702,N_3445,N_3402);
xor U3703 (N_3703,N_3498,N_3561);
or U3704 (N_3704,N_3459,N_3559);
xnor U3705 (N_3705,N_3412,N_3484);
or U3706 (N_3706,N_3563,N_3527);
xnor U3707 (N_3707,N_3441,N_3499);
nor U3708 (N_3708,N_3578,N_3512);
nand U3709 (N_3709,N_3470,N_3437);
nor U3710 (N_3710,N_3580,N_3426);
or U3711 (N_3711,N_3421,N_3503);
nand U3712 (N_3712,N_3522,N_3536);
nand U3713 (N_3713,N_3537,N_3480);
nor U3714 (N_3714,N_3401,N_3498);
and U3715 (N_3715,N_3534,N_3493);
nor U3716 (N_3716,N_3455,N_3597);
or U3717 (N_3717,N_3489,N_3567);
nand U3718 (N_3718,N_3566,N_3525);
nor U3719 (N_3719,N_3477,N_3595);
nand U3720 (N_3720,N_3504,N_3461);
nand U3721 (N_3721,N_3543,N_3552);
xor U3722 (N_3722,N_3448,N_3530);
nand U3723 (N_3723,N_3436,N_3437);
xor U3724 (N_3724,N_3462,N_3408);
nand U3725 (N_3725,N_3476,N_3542);
or U3726 (N_3726,N_3537,N_3584);
nor U3727 (N_3727,N_3585,N_3507);
and U3728 (N_3728,N_3426,N_3409);
nor U3729 (N_3729,N_3449,N_3581);
xor U3730 (N_3730,N_3503,N_3582);
and U3731 (N_3731,N_3400,N_3410);
or U3732 (N_3732,N_3543,N_3420);
nor U3733 (N_3733,N_3593,N_3474);
and U3734 (N_3734,N_3599,N_3438);
nand U3735 (N_3735,N_3493,N_3589);
nand U3736 (N_3736,N_3401,N_3486);
or U3737 (N_3737,N_3539,N_3425);
or U3738 (N_3738,N_3571,N_3576);
xnor U3739 (N_3739,N_3539,N_3594);
or U3740 (N_3740,N_3425,N_3432);
xor U3741 (N_3741,N_3561,N_3441);
nand U3742 (N_3742,N_3469,N_3482);
and U3743 (N_3743,N_3563,N_3555);
or U3744 (N_3744,N_3454,N_3504);
xnor U3745 (N_3745,N_3477,N_3549);
nor U3746 (N_3746,N_3473,N_3558);
or U3747 (N_3747,N_3561,N_3565);
or U3748 (N_3748,N_3534,N_3555);
and U3749 (N_3749,N_3498,N_3487);
xnor U3750 (N_3750,N_3467,N_3568);
nor U3751 (N_3751,N_3571,N_3586);
and U3752 (N_3752,N_3428,N_3480);
nor U3753 (N_3753,N_3498,N_3461);
nor U3754 (N_3754,N_3546,N_3451);
nor U3755 (N_3755,N_3504,N_3464);
nor U3756 (N_3756,N_3511,N_3494);
and U3757 (N_3757,N_3432,N_3584);
and U3758 (N_3758,N_3491,N_3543);
nand U3759 (N_3759,N_3532,N_3408);
or U3760 (N_3760,N_3569,N_3535);
nor U3761 (N_3761,N_3592,N_3586);
nand U3762 (N_3762,N_3470,N_3555);
or U3763 (N_3763,N_3438,N_3459);
nor U3764 (N_3764,N_3469,N_3452);
nand U3765 (N_3765,N_3517,N_3453);
and U3766 (N_3766,N_3415,N_3504);
and U3767 (N_3767,N_3407,N_3541);
or U3768 (N_3768,N_3546,N_3426);
or U3769 (N_3769,N_3476,N_3420);
nor U3770 (N_3770,N_3573,N_3535);
nor U3771 (N_3771,N_3484,N_3400);
xnor U3772 (N_3772,N_3436,N_3465);
xnor U3773 (N_3773,N_3596,N_3419);
or U3774 (N_3774,N_3557,N_3476);
nor U3775 (N_3775,N_3503,N_3548);
nor U3776 (N_3776,N_3447,N_3566);
xor U3777 (N_3777,N_3475,N_3445);
xnor U3778 (N_3778,N_3486,N_3482);
or U3779 (N_3779,N_3419,N_3400);
nor U3780 (N_3780,N_3452,N_3578);
nand U3781 (N_3781,N_3486,N_3544);
nand U3782 (N_3782,N_3544,N_3548);
nand U3783 (N_3783,N_3424,N_3439);
or U3784 (N_3784,N_3413,N_3426);
and U3785 (N_3785,N_3419,N_3557);
nand U3786 (N_3786,N_3588,N_3443);
and U3787 (N_3787,N_3438,N_3433);
nand U3788 (N_3788,N_3595,N_3479);
and U3789 (N_3789,N_3573,N_3442);
xnor U3790 (N_3790,N_3468,N_3446);
and U3791 (N_3791,N_3488,N_3587);
xnor U3792 (N_3792,N_3517,N_3438);
nand U3793 (N_3793,N_3551,N_3439);
nand U3794 (N_3794,N_3435,N_3431);
nand U3795 (N_3795,N_3558,N_3502);
and U3796 (N_3796,N_3503,N_3527);
nor U3797 (N_3797,N_3568,N_3464);
nor U3798 (N_3798,N_3518,N_3507);
nand U3799 (N_3799,N_3537,N_3495);
or U3800 (N_3800,N_3768,N_3749);
nor U3801 (N_3801,N_3604,N_3715);
nand U3802 (N_3802,N_3607,N_3634);
and U3803 (N_3803,N_3698,N_3627);
or U3804 (N_3804,N_3603,N_3663);
nor U3805 (N_3805,N_3703,N_3655);
and U3806 (N_3806,N_3732,N_3696);
nor U3807 (N_3807,N_3741,N_3693);
xor U3808 (N_3808,N_3700,N_3637);
or U3809 (N_3809,N_3785,N_3714);
and U3810 (N_3810,N_3636,N_3738);
and U3811 (N_3811,N_3769,N_3601);
nand U3812 (N_3812,N_3695,N_3684);
nor U3813 (N_3813,N_3620,N_3667);
nand U3814 (N_3814,N_3639,N_3721);
nor U3815 (N_3815,N_3600,N_3681);
nand U3816 (N_3816,N_3730,N_3668);
and U3817 (N_3817,N_3635,N_3725);
or U3818 (N_3818,N_3756,N_3778);
xor U3819 (N_3819,N_3746,N_3711);
xor U3820 (N_3820,N_3617,N_3680);
and U3821 (N_3821,N_3774,N_3657);
xor U3822 (N_3822,N_3767,N_3609);
nand U3823 (N_3823,N_3632,N_3688);
nor U3824 (N_3824,N_3709,N_3705);
or U3825 (N_3825,N_3618,N_3679);
and U3826 (N_3826,N_3704,N_3644);
and U3827 (N_3827,N_3777,N_3613);
or U3828 (N_3828,N_3716,N_3640);
and U3829 (N_3829,N_3788,N_3702);
or U3830 (N_3830,N_3687,N_3792);
nand U3831 (N_3831,N_3628,N_3674);
nor U3832 (N_3832,N_3676,N_3795);
and U3833 (N_3833,N_3659,N_3762);
nor U3834 (N_3834,N_3685,N_3648);
nand U3835 (N_3835,N_3727,N_3699);
or U3836 (N_3836,N_3694,N_3686);
or U3837 (N_3837,N_3625,N_3775);
nor U3838 (N_3838,N_3757,N_3656);
xor U3839 (N_3839,N_3758,N_3755);
nor U3840 (N_3840,N_3610,N_3664);
or U3841 (N_3841,N_3643,N_3759);
and U3842 (N_3842,N_3733,N_3739);
and U3843 (N_3843,N_3649,N_3658);
or U3844 (N_3844,N_3707,N_3682);
nor U3845 (N_3845,N_3708,N_3740);
and U3846 (N_3846,N_3671,N_3623);
nor U3847 (N_3847,N_3771,N_3787);
or U3848 (N_3848,N_3670,N_3605);
xnor U3849 (N_3849,N_3798,N_3719);
or U3850 (N_3850,N_3744,N_3742);
or U3851 (N_3851,N_3784,N_3776);
nor U3852 (N_3852,N_3647,N_3736);
nor U3853 (N_3853,N_3669,N_3765);
or U3854 (N_3854,N_3629,N_3726);
xnor U3855 (N_3855,N_3691,N_3672);
and U3856 (N_3856,N_3723,N_3772);
xor U3857 (N_3857,N_3764,N_3683);
xnor U3858 (N_3858,N_3645,N_3677);
or U3859 (N_3859,N_3633,N_3641);
nand U3860 (N_3860,N_3750,N_3616);
nor U3861 (N_3861,N_3763,N_3630);
or U3862 (N_3862,N_3783,N_3794);
nand U3863 (N_3863,N_3780,N_3608);
or U3864 (N_3864,N_3761,N_3754);
or U3865 (N_3865,N_3747,N_3712);
or U3866 (N_3866,N_3722,N_3770);
xnor U3867 (N_3867,N_3697,N_3622);
or U3868 (N_3868,N_3766,N_3642);
and U3869 (N_3869,N_3734,N_3638);
xnor U3870 (N_3870,N_3673,N_3621);
xnor U3871 (N_3871,N_3602,N_3678);
and U3872 (N_3872,N_3729,N_3753);
and U3873 (N_3873,N_3713,N_3654);
and U3874 (N_3874,N_3790,N_3720);
xnor U3875 (N_3875,N_3631,N_3653);
nor U3876 (N_3876,N_3748,N_3760);
nand U3877 (N_3877,N_3710,N_3796);
nor U3878 (N_3878,N_3717,N_3665);
xor U3879 (N_3879,N_3799,N_3662);
and U3880 (N_3880,N_3735,N_3619);
xnor U3881 (N_3881,N_3652,N_3782);
xnor U3882 (N_3882,N_3615,N_3706);
nand U3883 (N_3883,N_3661,N_3612);
or U3884 (N_3884,N_3660,N_3773);
nand U3885 (N_3885,N_3737,N_3724);
nor U3886 (N_3886,N_3690,N_3745);
xor U3887 (N_3887,N_3779,N_3666);
nor U3888 (N_3888,N_3797,N_3651);
xnor U3889 (N_3889,N_3611,N_3701);
nor U3890 (N_3890,N_3791,N_3752);
nand U3891 (N_3891,N_3751,N_3626);
nand U3892 (N_3892,N_3781,N_3731);
xnor U3893 (N_3893,N_3689,N_3718);
nand U3894 (N_3894,N_3692,N_3606);
xor U3895 (N_3895,N_3786,N_3624);
nand U3896 (N_3896,N_3793,N_3743);
xnor U3897 (N_3897,N_3650,N_3728);
nor U3898 (N_3898,N_3789,N_3646);
xor U3899 (N_3899,N_3675,N_3614);
or U3900 (N_3900,N_3647,N_3737);
or U3901 (N_3901,N_3693,N_3623);
and U3902 (N_3902,N_3643,N_3686);
nand U3903 (N_3903,N_3691,N_3724);
nor U3904 (N_3904,N_3762,N_3677);
or U3905 (N_3905,N_3768,N_3626);
nor U3906 (N_3906,N_3642,N_3776);
xor U3907 (N_3907,N_3629,N_3699);
xor U3908 (N_3908,N_3693,N_3709);
or U3909 (N_3909,N_3781,N_3611);
nor U3910 (N_3910,N_3704,N_3696);
xnor U3911 (N_3911,N_3797,N_3699);
xnor U3912 (N_3912,N_3723,N_3696);
or U3913 (N_3913,N_3704,N_3693);
xnor U3914 (N_3914,N_3769,N_3699);
nor U3915 (N_3915,N_3696,N_3671);
nand U3916 (N_3916,N_3613,N_3795);
or U3917 (N_3917,N_3708,N_3709);
and U3918 (N_3918,N_3699,N_3622);
nand U3919 (N_3919,N_3672,N_3632);
nand U3920 (N_3920,N_3626,N_3649);
xnor U3921 (N_3921,N_3652,N_3762);
and U3922 (N_3922,N_3778,N_3727);
nand U3923 (N_3923,N_3611,N_3712);
xnor U3924 (N_3924,N_3654,N_3746);
and U3925 (N_3925,N_3692,N_3635);
and U3926 (N_3926,N_3787,N_3690);
xnor U3927 (N_3927,N_3757,N_3786);
nand U3928 (N_3928,N_3653,N_3620);
nand U3929 (N_3929,N_3619,N_3742);
nand U3930 (N_3930,N_3627,N_3734);
and U3931 (N_3931,N_3628,N_3615);
nand U3932 (N_3932,N_3703,N_3709);
and U3933 (N_3933,N_3720,N_3608);
xor U3934 (N_3934,N_3702,N_3768);
and U3935 (N_3935,N_3699,N_3603);
nor U3936 (N_3936,N_3665,N_3678);
and U3937 (N_3937,N_3730,N_3765);
and U3938 (N_3938,N_3660,N_3643);
and U3939 (N_3939,N_3786,N_3770);
and U3940 (N_3940,N_3728,N_3755);
xnor U3941 (N_3941,N_3772,N_3638);
xor U3942 (N_3942,N_3736,N_3632);
or U3943 (N_3943,N_3603,N_3784);
or U3944 (N_3944,N_3623,N_3733);
or U3945 (N_3945,N_3728,N_3746);
xor U3946 (N_3946,N_3629,N_3755);
nand U3947 (N_3947,N_3669,N_3740);
or U3948 (N_3948,N_3614,N_3779);
or U3949 (N_3949,N_3746,N_3762);
and U3950 (N_3950,N_3687,N_3630);
nor U3951 (N_3951,N_3799,N_3753);
xor U3952 (N_3952,N_3672,N_3627);
xnor U3953 (N_3953,N_3681,N_3684);
or U3954 (N_3954,N_3722,N_3669);
xor U3955 (N_3955,N_3600,N_3753);
or U3956 (N_3956,N_3617,N_3774);
or U3957 (N_3957,N_3786,N_3691);
xnor U3958 (N_3958,N_3602,N_3715);
nor U3959 (N_3959,N_3770,N_3724);
nand U3960 (N_3960,N_3796,N_3700);
or U3961 (N_3961,N_3601,N_3782);
xor U3962 (N_3962,N_3672,N_3676);
and U3963 (N_3963,N_3718,N_3701);
nand U3964 (N_3964,N_3666,N_3724);
and U3965 (N_3965,N_3749,N_3684);
xor U3966 (N_3966,N_3776,N_3648);
and U3967 (N_3967,N_3735,N_3795);
xor U3968 (N_3968,N_3655,N_3751);
or U3969 (N_3969,N_3783,N_3695);
or U3970 (N_3970,N_3655,N_3700);
nor U3971 (N_3971,N_3663,N_3785);
and U3972 (N_3972,N_3707,N_3768);
and U3973 (N_3973,N_3779,N_3623);
nand U3974 (N_3974,N_3647,N_3654);
nand U3975 (N_3975,N_3612,N_3794);
or U3976 (N_3976,N_3750,N_3625);
nor U3977 (N_3977,N_3689,N_3613);
nand U3978 (N_3978,N_3702,N_3670);
nor U3979 (N_3979,N_3685,N_3703);
nand U3980 (N_3980,N_3722,N_3789);
xor U3981 (N_3981,N_3681,N_3677);
xor U3982 (N_3982,N_3642,N_3758);
and U3983 (N_3983,N_3744,N_3729);
nor U3984 (N_3984,N_3634,N_3790);
xnor U3985 (N_3985,N_3652,N_3678);
or U3986 (N_3986,N_3706,N_3665);
xor U3987 (N_3987,N_3674,N_3705);
xnor U3988 (N_3988,N_3701,N_3726);
nand U3989 (N_3989,N_3770,N_3753);
xnor U3990 (N_3990,N_3780,N_3631);
and U3991 (N_3991,N_3620,N_3753);
nand U3992 (N_3992,N_3637,N_3723);
xor U3993 (N_3993,N_3656,N_3749);
or U3994 (N_3994,N_3747,N_3693);
nor U3995 (N_3995,N_3606,N_3771);
or U3996 (N_3996,N_3780,N_3726);
nand U3997 (N_3997,N_3631,N_3674);
xnor U3998 (N_3998,N_3674,N_3647);
or U3999 (N_3999,N_3753,N_3739);
or U4000 (N_4000,N_3937,N_3924);
nor U4001 (N_4001,N_3877,N_3868);
xor U4002 (N_4002,N_3839,N_3825);
and U4003 (N_4003,N_3837,N_3899);
or U4004 (N_4004,N_3863,N_3938);
and U4005 (N_4005,N_3923,N_3889);
nor U4006 (N_4006,N_3892,N_3961);
nor U4007 (N_4007,N_3830,N_3955);
xor U4008 (N_4008,N_3990,N_3968);
and U4009 (N_4009,N_3921,N_3823);
and U4010 (N_4010,N_3907,N_3959);
and U4011 (N_4011,N_3926,N_3940);
nor U4012 (N_4012,N_3887,N_3883);
nand U4013 (N_4013,N_3953,N_3972);
or U4014 (N_4014,N_3956,N_3919);
or U4015 (N_4015,N_3845,N_3808);
nand U4016 (N_4016,N_3894,N_3895);
nor U4017 (N_4017,N_3901,N_3958);
xnor U4018 (N_4018,N_3971,N_3866);
and U4019 (N_4019,N_3975,N_3912);
and U4020 (N_4020,N_3976,N_3950);
and U4021 (N_4021,N_3900,N_3902);
or U4022 (N_4022,N_3982,N_3852);
xor U4023 (N_4023,N_3985,N_3980);
and U4024 (N_4024,N_3934,N_3947);
nand U4025 (N_4025,N_3893,N_3915);
and U4026 (N_4026,N_3995,N_3939);
or U4027 (N_4027,N_3865,N_3843);
nand U4028 (N_4028,N_3917,N_3842);
or U4029 (N_4029,N_3810,N_3989);
and U4030 (N_4030,N_3898,N_3993);
nor U4031 (N_4031,N_3960,N_3874);
nor U4032 (N_4032,N_3831,N_3964);
nor U4033 (N_4033,N_3962,N_3970);
xnor U4034 (N_4034,N_3858,N_3954);
xnor U4035 (N_4035,N_3822,N_3983);
xnor U4036 (N_4036,N_3946,N_3813);
nor U4037 (N_4037,N_3996,N_3911);
and U4038 (N_4038,N_3806,N_3826);
nor U4039 (N_4039,N_3966,N_3849);
nand U4040 (N_4040,N_3903,N_3851);
and U4041 (N_4041,N_3832,N_3875);
or U4042 (N_4042,N_3999,N_3988);
nor U4043 (N_4043,N_3977,N_3978);
nor U4044 (N_4044,N_3871,N_3876);
or U4045 (N_4045,N_3801,N_3969);
xor U4046 (N_4046,N_3994,N_3827);
nor U4047 (N_4047,N_3909,N_3949);
nor U4048 (N_4048,N_3974,N_3981);
xor U4049 (N_4049,N_3848,N_3906);
nand U4050 (N_4050,N_3885,N_3836);
nand U4051 (N_4051,N_3884,N_3914);
or U4052 (N_4052,N_3847,N_3897);
or U4053 (N_4053,N_3805,N_3841);
nand U4054 (N_4054,N_3828,N_3821);
and U4055 (N_4055,N_3869,N_3824);
nor U4056 (N_4056,N_3834,N_3853);
and U4057 (N_4057,N_3931,N_3922);
nand U4058 (N_4058,N_3935,N_3920);
xnor U4059 (N_4059,N_3802,N_3862);
nor U4060 (N_4060,N_3927,N_3857);
xor U4061 (N_4061,N_3930,N_3973);
nand U4062 (N_4062,N_3818,N_3814);
nand U4063 (N_4063,N_3929,N_3979);
xnor U4064 (N_4064,N_3846,N_3859);
nand U4065 (N_4065,N_3856,N_3967);
nand U4066 (N_4066,N_3891,N_3942);
xor U4067 (N_4067,N_3844,N_3873);
or U4068 (N_4068,N_3888,N_3916);
nand U4069 (N_4069,N_3881,N_3872);
nor U4070 (N_4070,N_3833,N_3992);
nand U4071 (N_4071,N_3951,N_3804);
nand U4072 (N_4072,N_3997,N_3910);
xnor U4073 (N_4073,N_3936,N_3854);
nand U4074 (N_4074,N_3835,N_3944);
or U4075 (N_4075,N_3800,N_3918);
xor U4076 (N_4076,N_3945,N_3803);
xnor U4077 (N_4077,N_3840,N_3896);
nor U4078 (N_4078,N_3984,N_3890);
nor U4079 (N_4079,N_3807,N_3880);
or U4080 (N_4080,N_3998,N_3838);
nor U4081 (N_4081,N_3817,N_3867);
nand U4082 (N_4082,N_3886,N_3965);
or U4083 (N_4083,N_3908,N_3957);
and U4084 (N_4084,N_3882,N_3913);
or U4085 (N_4085,N_3948,N_3986);
or U4086 (N_4086,N_3819,N_3879);
nor U4087 (N_4087,N_3855,N_3928);
xnor U4088 (N_4088,N_3850,N_3815);
nor U4089 (N_4089,N_3809,N_3991);
and U4090 (N_4090,N_3860,N_3904);
or U4091 (N_4091,N_3952,N_3932);
nor U4092 (N_4092,N_3816,N_3861);
nand U4093 (N_4093,N_3987,N_3941);
xnor U4094 (N_4094,N_3864,N_3933);
nand U4095 (N_4095,N_3905,N_3820);
nand U4096 (N_4096,N_3943,N_3829);
or U4097 (N_4097,N_3870,N_3811);
nand U4098 (N_4098,N_3925,N_3812);
or U4099 (N_4099,N_3878,N_3963);
and U4100 (N_4100,N_3928,N_3986);
and U4101 (N_4101,N_3985,N_3839);
nand U4102 (N_4102,N_3977,N_3986);
nor U4103 (N_4103,N_3914,N_3841);
nand U4104 (N_4104,N_3989,N_3918);
or U4105 (N_4105,N_3842,N_3908);
nand U4106 (N_4106,N_3913,N_3838);
nor U4107 (N_4107,N_3859,N_3939);
nor U4108 (N_4108,N_3846,N_3809);
nand U4109 (N_4109,N_3954,N_3872);
or U4110 (N_4110,N_3923,N_3992);
or U4111 (N_4111,N_3931,N_3837);
xnor U4112 (N_4112,N_3954,N_3919);
xnor U4113 (N_4113,N_3812,N_3831);
and U4114 (N_4114,N_3966,N_3848);
and U4115 (N_4115,N_3811,N_3955);
or U4116 (N_4116,N_3831,N_3903);
and U4117 (N_4117,N_3888,N_3946);
and U4118 (N_4118,N_3827,N_3826);
and U4119 (N_4119,N_3823,N_3951);
or U4120 (N_4120,N_3871,N_3864);
nor U4121 (N_4121,N_3962,N_3830);
xnor U4122 (N_4122,N_3908,N_3925);
nand U4123 (N_4123,N_3834,N_3965);
nor U4124 (N_4124,N_3921,N_3953);
or U4125 (N_4125,N_3942,N_3935);
xnor U4126 (N_4126,N_3993,N_3859);
and U4127 (N_4127,N_3809,N_3821);
nand U4128 (N_4128,N_3860,N_3926);
nor U4129 (N_4129,N_3846,N_3901);
and U4130 (N_4130,N_3904,N_3864);
or U4131 (N_4131,N_3931,N_3831);
xnor U4132 (N_4132,N_3805,N_3826);
nand U4133 (N_4133,N_3857,N_3974);
or U4134 (N_4134,N_3840,N_3874);
or U4135 (N_4135,N_3924,N_3865);
or U4136 (N_4136,N_3899,N_3942);
xnor U4137 (N_4137,N_3904,N_3819);
xnor U4138 (N_4138,N_3837,N_3979);
nor U4139 (N_4139,N_3893,N_3874);
or U4140 (N_4140,N_3847,N_3808);
xnor U4141 (N_4141,N_3992,N_3977);
xor U4142 (N_4142,N_3838,N_3841);
nor U4143 (N_4143,N_3849,N_3958);
nor U4144 (N_4144,N_3895,N_3918);
xnor U4145 (N_4145,N_3966,N_3869);
xnor U4146 (N_4146,N_3866,N_3826);
nand U4147 (N_4147,N_3831,N_3982);
xnor U4148 (N_4148,N_3835,N_3837);
nand U4149 (N_4149,N_3937,N_3805);
xnor U4150 (N_4150,N_3985,N_3917);
and U4151 (N_4151,N_3993,N_3895);
or U4152 (N_4152,N_3840,N_3960);
xnor U4153 (N_4153,N_3855,N_3926);
or U4154 (N_4154,N_3889,N_3877);
nor U4155 (N_4155,N_3889,N_3811);
nor U4156 (N_4156,N_3906,N_3845);
and U4157 (N_4157,N_3912,N_3966);
xor U4158 (N_4158,N_3829,N_3916);
and U4159 (N_4159,N_3884,N_3821);
xnor U4160 (N_4160,N_3870,N_3812);
or U4161 (N_4161,N_3952,N_3837);
nor U4162 (N_4162,N_3853,N_3944);
nor U4163 (N_4163,N_3971,N_3815);
nand U4164 (N_4164,N_3891,N_3951);
nand U4165 (N_4165,N_3811,N_3892);
xnor U4166 (N_4166,N_3812,N_3988);
xnor U4167 (N_4167,N_3936,N_3888);
nor U4168 (N_4168,N_3923,N_3989);
nand U4169 (N_4169,N_3888,N_3933);
nand U4170 (N_4170,N_3818,N_3842);
and U4171 (N_4171,N_3973,N_3874);
nor U4172 (N_4172,N_3996,N_3803);
or U4173 (N_4173,N_3890,N_3968);
xor U4174 (N_4174,N_3948,N_3944);
xnor U4175 (N_4175,N_3905,N_3950);
or U4176 (N_4176,N_3946,N_3999);
xnor U4177 (N_4177,N_3924,N_3994);
or U4178 (N_4178,N_3979,N_3963);
or U4179 (N_4179,N_3947,N_3802);
nand U4180 (N_4180,N_3851,N_3929);
nand U4181 (N_4181,N_3847,N_3842);
or U4182 (N_4182,N_3909,N_3885);
xor U4183 (N_4183,N_3856,N_3961);
and U4184 (N_4184,N_3838,N_3844);
and U4185 (N_4185,N_3845,N_3819);
nand U4186 (N_4186,N_3897,N_3928);
nand U4187 (N_4187,N_3984,N_3987);
nand U4188 (N_4188,N_3983,N_3976);
or U4189 (N_4189,N_3983,N_3924);
nor U4190 (N_4190,N_3852,N_3908);
xor U4191 (N_4191,N_3812,N_3848);
xor U4192 (N_4192,N_3819,N_3936);
nand U4193 (N_4193,N_3856,N_3947);
nand U4194 (N_4194,N_3830,N_3983);
and U4195 (N_4195,N_3875,N_3882);
nor U4196 (N_4196,N_3844,N_3992);
nand U4197 (N_4197,N_3899,N_3916);
and U4198 (N_4198,N_3992,N_3830);
or U4199 (N_4199,N_3931,N_3957);
nor U4200 (N_4200,N_4051,N_4064);
xnor U4201 (N_4201,N_4158,N_4054);
nand U4202 (N_4202,N_4141,N_4165);
nor U4203 (N_4203,N_4090,N_4146);
nor U4204 (N_4204,N_4034,N_4110);
nor U4205 (N_4205,N_4143,N_4097);
xor U4206 (N_4206,N_4013,N_4018);
and U4207 (N_4207,N_4038,N_4198);
nand U4208 (N_4208,N_4063,N_4183);
nand U4209 (N_4209,N_4022,N_4071);
xor U4210 (N_4210,N_4060,N_4056);
or U4211 (N_4211,N_4148,N_4108);
nor U4212 (N_4212,N_4027,N_4138);
xor U4213 (N_4213,N_4073,N_4040);
or U4214 (N_4214,N_4029,N_4070);
nor U4215 (N_4215,N_4048,N_4014);
and U4216 (N_4216,N_4155,N_4190);
or U4217 (N_4217,N_4062,N_4150);
xnor U4218 (N_4218,N_4119,N_4001);
xor U4219 (N_4219,N_4164,N_4153);
and U4220 (N_4220,N_4095,N_4188);
nor U4221 (N_4221,N_4181,N_4159);
xor U4222 (N_4222,N_4160,N_4086);
nand U4223 (N_4223,N_4025,N_4006);
xor U4224 (N_4224,N_4145,N_4082);
or U4225 (N_4225,N_4170,N_4067);
xor U4226 (N_4226,N_4099,N_4123);
or U4227 (N_4227,N_4078,N_4179);
and U4228 (N_4228,N_4177,N_4065);
xnor U4229 (N_4229,N_4135,N_4031);
or U4230 (N_4230,N_4166,N_4028);
and U4231 (N_4231,N_4147,N_4168);
nor U4232 (N_4232,N_4017,N_4058);
xnor U4233 (N_4233,N_4186,N_4093);
and U4234 (N_4234,N_4121,N_4197);
xor U4235 (N_4235,N_4049,N_4050);
nand U4236 (N_4236,N_4039,N_4035);
or U4237 (N_4237,N_4075,N_4195);
xnor U4238 (N_4238,N_4107,N_4068);
xnor U4239 (N_4239,N_4003,N_4131);
and U4240 (N_4240,N_4194,N_4045);
nor U4241 (N_4241,N_4191,N_4047);
xor U4242 (N_4242,N_4057,N_4124);
nor U4243 (N_4243,N_4019,N_4113);
nor U4244 (N_4244,N_4088,N_4137);
and U4245 (N_4245,N_4136,N_4098);
or U4246 (N_4246,N_4008,N_4042);
nor U4247 (N_4247,N_4021,N_4127);
and U4248 (N_4248,N_4052,N_4061);
xnor U4249 (N_4249,N_4005,N_4076);
or U4250 (N_4250,N_4026,N_4010);
nand U4251 (N_4251,N_4122,N_4174);
nor U4252 (N_4252,N_4133,N_4116);
nor U4253 (N_4253,N_4103,N_4134);
nor U4254 (N_4254,N_4009,N_4101);
nor U4255 (N_4255,N_4172,N_4091);
or U4256 (N_4256,N_4030,N_4012);
and U4257 (N_4257,N_4140,N_4176);
or U4258 (N_4258,N_4059,N_4069);
and U4259 (N_4259,N_4036,N_4199);
nor U4260 (N_4260,N_4041,N_4139);
nand U4261 (N_4261,N_4094,N_4184);
and U4262 (N_4262,N_4055,N_4152);
and U4263 (N_4263,N_4015,N_4044);
xnor U4264 (N_4264,N_4096,N_4154);
nor U4265 (N_4265,N_4128,N_4157);
and U4266 (N_4266,N_4118,N_4196);
xor U4267 (N_4267,N_4161,N_4020);
nand U4268 (N_4268,N_4072,N_4081);
xor U4269 (N_4269,N_4193,N_4002);
or U4270 (N_4270,N_4112,N_4007);
or U4271 (N_4271,N_4085,N_4192);
nand U4272 (N_4272,N_4126,N_4114);
xnor U4273 (N_4273,N_4032,N_4173);
nor U4274 (N_4274,N_4079,N_4167);
and U4275 (N_4275,N_4084,N_4080);
nand U4276 (N_4276,N_4077,N_4089);
xor U4277 (N_4277,N_4149,N_4185);
and U4278 (N_4278,N_4132,N_4043);
xor U4279 (N_4279,N_4125,N_4033);
nand U4280 (N_4280,N_4180,N_4046);
nand U4281 (N_4281,N_4106,N_4023);
xnor U4282 (N_4282,N_4144,N_4066);
nand U4283 (N_4283,N_4162,N_4092);
xor U4284 (N_4284,N_4178,N_4104);
xor U4285 (N_4285,N_4142,N_4130);
xor U4286 (N_4286,N_4011,N_4000);
or U4287 (N_4287,N_4053,N_4151);
xnor U4288 (N_4288,N_4156,N_4182);
nand U4289 (N_4289,N_4115,N_4117);
nand U4290 (N_4290,N_4016,N_4109);
nor U4291 (N_4291,N_4187,N_4169);
nand U4292 (N_4292,N_4074,N_4024);
nand U4293 (N_4293,N_4163,N_4189);
xnor U4294 (N_4294,N_4129,N_4083);
and U4295 (N_4295,N_4087,N_4004);
xnor U4296 (N_4296,N_4175,N_4037);
and U4297 (N_4297,N_4102,N_4111);
or U4298 (N_4298,N_4171,N_4105);
nand U4299 (N_4299,N_4100,N_4120);
and U4300 (N_4300,N_4019,N_4173);
and U4301 (N_4301,N_4178,N_4049);
or U4302 (N_4302,N_4127,N_4065);
xor U4303 (N_4303,N_4015,N_4059);
nand U4304 (N_4304,N_4171,N_4009);
nor U4305 (N_4305,N_4054,N_4076);
and U4306 (N_4306,N_4168,N_4068);
nand U4307 (N_4307,N_4191,N_4083);
and U4308 (N_4308,N_4194,N_4171);
nor U4309 (N_4309,N_4117,N_4008);
nor U4310 (N_4310,N_4058,N_4177);
nand U4311 (N_4311,N_4109,N_4098);
xor U4312 (N_4312,N_4184,N_4161);
nor U4313 (N_4313,N_4129,N_4020);
nor U4314 (N_4314,N_4064,N_4048);
or U4315 (N_4315,N_4041,N_4123);
nor U4316 (N_4316,N_4005,N_4196);
nand U4317 (N_4317,N_4136,N_4052);
nor U4318 (N_4318,N_4031,N_4005);
and U4319 (N_4319,N_4063,N_4062);
or U4320 (N_4320,N_4062,N_4174);
nand U4321 (N_4321,N_4028,N_4120);
nor U4322 (N_4322,N_4037,N_4101);
or U4323 (N_4323,N_4198,N_4087);
nor U4324 (N_4324,N_4113,N_4053);
or U4325 (N_4325,N_4020,N_4000);
or U4326 (N_4326,N_4002,N_4169);
and U4327 (N_4327,N_4152,N_4147);
nor U4328 (N_4328,N_4144,N_4069);
or U4329 (N_4329,N_4064,N_4150);
nand U4330 (N_4330,N_4148,N_4028);
or U4331 (N_4331,N_4138,N_4071);
xor U4332 (N_4332,N_4115,N_4089);
xnor U4333 (N_4333,N_4178,N_4154);
xnor U4334 (N_4334,N_4049,N_4131);
nor U4335 (N_4335,N_4063,N_4114);
nand U4336 (N_4336,N_4081,N_4060);
or U4337 (N_4337,N_4134,N_4091);
nand U4338 (N_4338,N_4083,N_4095);
nand U4339 (N_4339,N_4039,N_4106);
and U4340 (N_4340,N_4083,N_4052);
or U4341 (N_4341,N_4154,N_4130);
nand U4342 (N_4342,N_4070,N_4004);
or U4343 (N_4343,N_4048,N_4198);
xor U4344 (N_4344,N_4044,N_4062);
and U4345 (N_4345,N_4121,N_4029);
nand U4346 (N_4346,N_4088,N_4193);
nand U4347 (N_4347,N_4151,N_4011);
nor U4348 (N_4348,N_4141,N_4006);
xor U4349 (N_4349,N_4129,N_4058);
and U4350 (N_4350,N_4072,N_4109);
or U4351 (N_4351,N_4006,N_4067);
and U4352 (N_4352,N_4056,N_4114);
and U4353 (N_4353,N_4107,N_4027);
nand U4354 (N_4354,N_4186,N_4027);
nand U4355 (N_4355,N_4106,N_4044);
and U4356 (N_4356,N_4143,N_4136);
and U4357 (N_4357,N_4179,N_4007);
and U4358 (N_4358,N_4093,N_4158);
xnor U4359 (N_4359,N_4072,N_4187);
or U4360 (N_4360,N_4009,N_4168);
nor U4361 (N_4361,N_4190,N_4122);
and U4362 (N_4362,N_4156,N_4173);
nand U4363 (N_4363,N_4175,N_4006);
and U4364 (N_4364,N_4199,N_4018);
nand U4365 (N_4365,N_4110,N_4000);
nor U4366 (N_4366,N_4152,N_4016);
and U4367 (N_4367,N_4062,N_4125);
nand U4368 (N_4368,N_4095,N_4013);
nand U4369 (N_4369,N_4110,N_4015);
or U4370 (N_4370,N_4090,N_4195);
xor U4371 (N_4371,N_4007,N_4003);
or U4372 (N_4372,N_4186,N_4196);
or U4373 (N_4373,N_4189,N_4020);
nand U4374 (N_4374,N_4121,N_4153);
nor U4375 (N_4375,N_4107,N_4023);
xnor U4376 (N_4376,N_4171,N_4112);
xnor U4377 (N_4377,N_4000,N_4079);
nor U4378 (N_4378,N_4185,N_4198);
nand U4379 (N_4379,N_4080,N_4175);
nor U4380 (N_4380,N_4025,N_4002);
or U4381 (N_4381,N_4140,N_4010);
nand U4382 (N_4382,N_4114,N_4187);
nand U4383 (N_4383,N_4064,N_4138);
nor U4384 (N_4384,N_4179,N_4088);
and U4385 (N_4385,N_4180,N_4112);
and U4386 (N_4386,N_4138,N_4004);
xnor U4387 (N_4387,N_4050,N_4019);
and U4388 (N_4388,N_4166,N_4050);
nor U4389 (N_4389,N_4094,N_4000);
nand U4390 (N_4390,N_4026,N_4141);
nand U4391 (N_4391,N_4021,N_4108);
or U4392 (N_4392,N_4032,N_4168);
xor U4393 (N_4393,N_4113,N_4052);
or U4394 (N_4394,N_4126,N_4000);
xor U4395 (N_4395,N_4064,N_4029);
xor U4396 (N_4396,N_4047,N_4034);
and U4397 (N_4397,N_4156,N_4071);
or U4398 (N_4398,N_4023,N_4112);
xor U4399 (N_4399,N_4172,N_4052);
and U4400 (N_4400,N_4271,N_4216);
and U4401 (N_4401,N_4385,N_4345);
nor U4402 (N_4402,N_4340,N_4373);
nor U4403 (N_4403,N_4256,N_4293);
nand U4404 (N_4404,N_4357,N_4275);
xnor U4405 (N_4405,N_4378,N_4233);
and U4406 (N_4406,N_4370,N_4208);
or U4407 (N_4407,N_4310,N_4243);
nand U4408 (N_4408,N_4297,N_4278);
xnor U4409 (N_4409,N_4258,N_4205);
and U4410 (N_4410,N_4354,N_4228);
and U4411 (N_4411,N_4361,N_4213);
and U4412 (N_4412,N_4245,N_4248);
xnor U4413 (N_4413,N_4394,N_4353);
or U4414 (N_4414,N_4236,N_4250);
xnor U4415 (N_4415,N_4298,N_4269);
nand U4416 (N_4416,N_4322,N_4240);
or U4417 (N_4417,N_4399,N_4239);
xor U4418 (N_4418,N_4319,N_4257);
xor U4419 (N_4419,N_4302,N_4382);
and U4420 (N_4420,N_4253,N_4315);
and U4421 (N_4421,N_4262,N_4277);
xnor U4422 (N_4422,N_4380,N_4324);
nor U4423 (N_4423,N_4366,N_4300);
nand U4424 (N_4424,N_4368,N_4396);
or U4425 (N_4425,N_4395,N_4251);
and U4426 (N_4426,N_4393,N_4291);
nand U4427 (N_4427,N_4342,N_4305);
and U4428 (N_4428,N_4321,N_4212);
xnor U4429 (N_4429,N_4325,N_4219);
xnor U4430 (N_4430,N_4323,N_4367);
or U4431 (N_4431,N_4358,N_4365);
or U4432 (N_4432,N_4204,N_4254);
or U4433 (N_4433,N_4333,N_4252);
nand U4434 (N_4434,N_4210,N_4225);
and U4435 (N_4435,N_4303,N_4286);
nand U4436 (N_4436,N_4279,N_4246);
nand U4437 (N_4437,N_4392,N_4281);
nor U4438 (N_4438,N_4390,N_4371);
or U4439 (N_4439,N_4384,N_4311);
and U4440 (N_4440,N_4288,N_4261);
nand U4441 (N_4441,N_4346,N_4338);
nand U4442 (N_4442,N_4347,N_4352);
nor U4443 (N_4443,N_4318,N_4267);
nor U4444 (N_4444,N_4360,N_4398);
or U4445 (N_4445,N_4270,N_4383);
xor U4446 (N_4446,N_4217,N_4372);
and U4447 (N_4447,N_4351,N_4274);
nor U4448 (N_4448,N_4388,N_4249);
xnor U4449 (N_4449,N_4335,N_4306);
or U4450 (N_4450,N_4307,N_4223);
nand U4451 (N_4451,N_4255,N_4266);
xnor U4452 (N_4452,N_4285,N_4214);
xor U4453 (N_4453,N_4389,N_4329);
xnor U4454 (N_4454,N_4218,N_4276);
xnor U4455 (N_4455,N_4247,N_4290);
and U4456 (N_4456,N_4200,N_4272);
nand U4457 (N_4457,N_4209,N_4317);
and U4458 (N_4458,N_4296,N_4259);
xnor U4459 (N_4459,N_4234,N_4341);
and U4460 (N_4460,N_4202,N_4232);
and U4461 (N_4461,N_4230,N_4226);
or U4462 (N_4462,N_4241,N_4364);
nor U4463 (N_4463,N_4397,N_4375);
and U4464 (N_4464,N_4203,N_4350);
nand U4465 (N_4465,N_4283,N_4244);
or U4466 (N_4466,N_4289,N_4391);
nor U4467 (N_4467,N_4299,N_4220);
nor U4468 (N_4468,N_4237,N_4224);
and U4469 (N_4469,N_4260,N_4374);
nand U4470 (N_4470,N_4238,N_4334);
xor U4471 (N_4471,N_4332,N_4330);
xnor U4472 (N_4472,N_4222,N_4328);
nor U4473 (N_4473,N_4320,N_4355);
and U4474 (N_4474,N_4284,N_4227);
nand U4475 (N_4475,N_4304,N_4242);
and U4476 (N_4476,N_4211,N_4343);
nand U4477 (N_4477,N_4386,N_4316);
nand U4478 (N_4478,N_4294,N_4265);
xor U4479 (N_4479,N_4356,N_4377);
nand U4480 (N_4480,N_4369,N_4313);
xnor U4481 (N_4481,N_4337,N_4349);
nand U4482 (N_4482,N_4339,N_4363);
and U4483 (N_4483,N_4379,N_4201);
nand U4484 (N_4484,N_4326,N_4359);
or U4485 (N_4485,N_4309,N_4327);
or U4486 (N_4486,N_4235,N_4344);
nand U4487 (N_4487,N_4264,N_4231);
nor U4488 (N_4488,N_4282,N_4295);
nor U4489 (N_4489,N_4348,N_4221);
or U4490 (N_4490,N_4312,N_4336);
nor U4491 (N_4491,N_4206,N_4263);
and U4492 (N_4492,N_4381,N_4207);
xnor U4493 (N_4493,N_4287,N_4280);
xor U4494 (N_4494,N_4387,N_4215);
or U4495 (N_4495,N_4301,N_4331);
nor U4496 (N_4496,N_4314,N_4273);
nor U4497 (N_4497,N_4308,N_4376);
nand U4498 (N_4498,N_4268,N_4362);
xor U4499 (N_4499,N_4292,N_4229);
nand U4500 (N_4500,N_4291,N_4378);
nand U4501 (N_4501,N_4229,N_4291);
nor U4502 (N_4502,N_4374,N_4243);
and U4503 (N_4503,N_4327,N_4352);
nand U4504 (N_4504,N_4369,N_4372);
or U4505 (N_4505,N_4341,N_4203);
or U4506 (N_4506,N_4388,N_4203);
and U4507 (N_4507,N_4390,N_4202);
and U4508 (N_4508,N_4288,N_4217);
xor U4509 (N_4509,N_4393,N_4396);
or U4510 (N_4510,N_4212,N_4334);
or U4511 (N_4511,N_4370,N_4223);
nor U4512 (N_4512,N_4373,N_4211);
and U4513 (N_4513,N_4366,N_4277);
nor U4514 (N_4514,N_4354,N_4308);
xnor U4515 (N_4515,N_4248,N_4329);
nand U4516 (N_4516,N_4301,N_4307);
nand U4517 (N_4517,N_4252,N_4253);
or U4518 (N_4518,N_4375,N_4313);
or U4519 (N_4519,N_4222,N_4253);
xnor U4520 (N_4520,N_4219,N_4368);
xor U4521 (N_4521,N_4343,N_4262);
and U4522 (N_4522,N_4258,N_4251);
nand U4523 (N_4523,N_4372,N_4221);
nand U4524 (N_4524,N_4396,N_4298);
or U4525 (N_4525,N_4243,N_4383);
and U4526 (N_4526,N_4357,N_4399);
or U4527 (N_4527,N_4330,N_4262);
nor U4528 (N_4528,N_4339,N_4248);
and U4529 (N_4529,N_4357,N_4304);
and U4530 (N_4530,N_4378,N_4369);
and U4531 (N_4531,N_4387,N_4384);
xnor U4532 (N_4532,N_4239,N_4305);
nand U4533 (N_4533,N_4313,N_4269);
xor U4534 (N_4534,N_4225,N_4306);
xnor U4535 (N_4535,N_4327,N_4272);
xnor U4536 (N_4536,N_4298,N_4259);
nor U4537 (N_4537,N_4266,N_4322);
nor U4538 (N_4538,N_4211,N_4200);
and U4539 (N_4539,N_4239,N_4225);
and U4540 (N_4540,N_4202,N_4308);
or U4541 (N_4541,N_4308,N_4384);
or U4542 (N_4542,N_4250,N_4269);
and U4543 (N_4543,N_4271,N_4251);
nand U4544 (N_4544,N_4323,N_4297);
or U4545 (N_4545,N_4388,N_4288);
and U4546 (N_4546,N_4324,N_4358);
and U4547 (N_4547,N_4383,N_4240);
and U4548 (N_4548,N_4237,N_4205);
or U4549 (N_4549,N_4328,N_4377);
nor U4550 (N_4550,N_4299,N_4283);
and U4551 (N_4551,N_4275,N_4267);
nand U4552 (N_4552,N_4244,N_4376);
nand U4553 (N_4553,N_4324,N_4276);
nand U4554 (N_4554,N_4254,N_4308);
nand U4555 (N_4555,N_4299,N_4201);
or U4556 (N_4556,N_4226,N_4216);
xnor U4557 (N_4557,N_4275,N_4307);
nand U4558 (N_4558,N_4391,N_4213);
nor U4559 (N_4559,N_4309,N_4343);
and U4560 (N_4560,N_4361,N_4220);
nand U4561 (N_4561,N_4329,N_4204);
nand U4562 (N_4562,N_4212,N_4265);
nor U4563 (N_4563,N_4309,N_4381);
and U4564 (N_4564,N_4276,N_4317);
or U4565 (N_4565,N_4292,N_4338);
nand U4566 (N_4566,N_4203,N_4342);
or U4567 (N_4567,N_4289,N_4218);
xnor U4568 (N_4568,N_4293,N_4225);
nand U4569 (N_4569,N_4270,N_4290);
nor U4570 (N_4570,N_4383,N_4307);
or U4571 (N_4571,N_4388,N_4284);
xnor U4572 (N_4572,N_4238,N_4306);
nor U4573 (N_4573,N_4284,N_4323);
nand U4574 (N_4574,N_4267,N_4311);
nor U4575 (N_4575,N_4200,N_4359);
nor U4576 (N_4576,N_4255,N_4279);
nor U4577 (N_4577,N_4387,N_4359);
xor U4578 (N_4578,N_4395,N_4228);
nor U4579 (N_4579,N_4270,N_4320);
nand U4580 (N_4580,N_4331,N_4375);
nor U4581 (N_4581,N_4356,N_4291);
or U4582 (N_4582,N_4394,N_4335);
nor U4583 (N_4583,N_4327,N_4368);
and U4584 (N_4584,N_4221,N_4313);
nand U4585 (N_4585,N_4272,N_4382);
nand U4586 (N_4586,N_4372,N_4345);
nor U4587 (N_4587,N_4257,N_4201);
xor U4588 (N_4588,N_4300,N_4365);
xnor U4589 (N_4589,N_4253,N_4273);
nor U4590 (N_4590,N_4341,N_4216);
and U4591 (N_4591,N_4217,N_4310);
nor U4592 (N_4592,N_4333,N_4335);
xor U4593 (N_4593,N_4349,N_4243);
and U4594 (N_4594,N_4265,N_4360);
or U4595 (N_4595,N_4246,N_4388);
or U4596 (N_4596,N_4224,N_4341);
and U4597 (N_4597,N_4321,N_4327);
xor U4598 (N_4598,N_4393,N_4280);
and U4599 (N_4599,N_4261,N_4347);
and U4600 (N_4600,N_4406,N_4563);
nand U4601 (N_4601,N_4560,N_4454);
and U4602 (N_4602,N_4511,N_4449);
and U4603 (N_4603,N_4523,N_4445);
nor U4604 (N_4604,N_4478,N_4405);
xnor U4605 (N_4605,N_4404,N_4517);
xor U4606 (N_4606,N_4474,N_4467);
nor U4607 (N_4607,N_4562,N_4420);
nor U4608 (N_4608,N_4479,N_4427);
and U4609 (N_4609,N_4520,N_4482);
and U4610 (N_4610,N_4400,N_4456);
or U4611 (N_4611,N_4576,N_4458);
nor U4612 (N_4612,N_4512,N_4413);
and U4613 (N_4613,N_4419,N_4531);
and U4614 (N_4614,N_4503,N_4481);
nand U4615 (N_4615,N_4446,N_4425);
and U4616 (N_4616,N_4428,N_4593);
or U4617 (N_4617,N_4586,N_4522);
nand U4618 (N_4618,N_4549,N_4496);
xor U4619 (N_4619,N_4514,N_4533);
nand U4620 (N_4620,N_4436,N_4554);
and U4621 (N_4621,N_4594,N_4537);
xnor U4622 (N_4622,N_4557,N_4455);
nor U4623 (N_4623,N_4439,N_4519);
xor U4624 (N_4624,N_4542,N_4410);
nand U4625 (N_4625,N_4421,N_4493);
nand U4626 (N_4626,N_4408,N_4566);
or U4627 (N_4627,N_4555,N_4444);
xnor U4628 (N_4628,N_4575,N_4460);
nor U4629 (N_4629,N_4561,N_4508);
xor U4630 (N_4630,N_4471,N_4585);
and U4631 (N_4631,N_4409,N_4590);
or U4632 (N_4632,N_4592,N_4556);
and U4633 (N_4633,N_4553,N_4491);
nor U4634 (N_4634,N_4495,N_4475);
or U4635 (N_4635,N_4476,N_4488);
or U4636 (N_4636,N_4498,N_4530);
and U4637 (N_4637,N_4581,N_4435);
nor U4638 (N_4638,N_4422,N_4415);
and U4639 (N_4639,N_4452,N_4483);
nor U4640 (N_4640,N_4538,N_4429);
nand U4641 (N_4641,N_4571,N_4525);
nor U4642 (N_4642,N_4426,N_4540);
xnor U4643 (N_4643,N_4587,N_4434);
nand U4644 (N_4644,N_4453,N_4521);
nor U4645 (N_4645,N_4490,N_4598);
and U4646 (N_4646,N_4595,N_4416);
xnor U4647 (N_4647,N_4582,N_4599);
or U4648 (N_4648,N_4507,N_4527);
xor U4649 (N_4649,N_4567,N_4448);
and U4650 (N_4650,N_4486,N_4532);
and U4651 (N_4651,N_4465,N_4545);
xor U4652 (N_4652,N_4552,N_4457);
nor U4653 (N_4653,N_4492,N_4461);
and U4654 (N_4654,N_4577,N_4580);
nor U4655 (N_4655,N_4513,N_4485);
and U4656 (N_4656,N_4499,N_4418);
nor U4657 (N_4657,N_4526,N_4588);
nor U4658 (N_4658,N_4430,N_4411);
nand U4659 (N_4659,N_4569,N_4472);
and U4660 (N_4660,N_4441,N_4468);
nand U4661 (N_4661,N_4583,N_4402);
nand U4662 (N_4662,N_4447,N_4509);
or U4663 (N_4663,N_4414,N_4559);
xnor U4664 (N_4664,N_4412,N_4546);
and U4665 (N_4665,N_4459,N_4529);
nor U4666 (N_4666,N_4502,N_4494);
and U4667 (N_4667,N_4535,N_4463);
or U4668 (N_4668,N_4423,N_4536);
or U4669 (N_4669,N_4548,N_4438);
xor U4670 (N_4670,N_4565,N_4489);
and U4671 (N_4671,N_4437,N_4544);
nand U4672 (N_4672,N_4477,N_4506);
or U4673 (N_4673,N_4473,N_4596);
and U4674 (N_4674,N_4505,N_4589);
and U4675 (N_4675,N_4487,N_4431);
and U4676 (N_4676,N_4510,N_4442);
and U4677 (N_4677,N_4504,N_4401);
and U4678 (N_4678,N_4464,N_4534);
and U4679 (N_4679,N_4558,N_4578);
and U4680 (N_4680,N_4572,N_4450);
and U4681 (N_4681,N_4497,N_4484);
nand U4682 (N_4682,N_4480,N_4524);
xor U4683 (N_4683,N_4451,N_4584);
nand U4684 (N_4684,N_4500,N_4501);
nor U4685 (N_4685,N_4433,N_4417);
and U4686 (N_4686,N_4403,N_4424);
nand U4687 (N_4687,N_4470,N_4570);
nand U4688 (N_4688,N_4550,N_4462);
nand U4689 (N_4689,N_4573,N_4516);
nor U4690 (N_4690,N_4528,N_4547);
nand U4691 (N_4691,N_4515,N_4518);
and U4692 (N_4692,N_4466,N_4564);
nand U4693 (N_4693,N_4543,N_4597);
and U4694 (N_4694,N_4551,N_4568);
and U4695 (N_4695,N_4440,N_4539);
and U4696 (N_4696,N_4574,N_4469);
nand U4697 (N_4697,N_4541,N_4432);
and U4698 (N_4698,N_4591,N_4443);
nor U4699 (N_4699,N_4579,N_4407);
or U4700 (N_4700,N_4440,N_4400);
nand U4701 (N_4701,N_4519,N_4445);
or U4702 (N_4702,N_4531,N_4597);
nand U4703 (N_4703,N_4574,N_4493);
nand U4704 (N_4704,N_4552,N_4582);
xnor U4705 (N_4705,N_4524,N_4543);
and U4706 (N_4706,N_4554,N_4593);
nand U4707 (N_4707,N_4545,N_4457);
xor U4708 (N_4708,N_4555,N_4524);
nor U4709 (N_4709,N_4427,N_4528);
nor U4710 (N_4710,N_4455,N_4579);
or U4711 (N_4711,N_4513,N_4491);
or U4712 (N_4712,N_4411,N_4536);
and U4713 (N_4713,N_4491,N_4454);
and U4714 (N_4714,N_4478,N_4468);
nor U4715 (N_4715,N_4562,N_4527);
nor U4716 (N_4716,N_4449,N_4519);
nand U4717 (N_4717,N_4407,N_4483);
xor U4718 (N_4718,N_4574,N_4482);
nor U4719 (N_4719,N_4562,N_4545);
or U4720 (N_4720,N_4495,N_4525);
nor U4721 (N_4721,N_4452,N_4411);
and U4722 (N_4722,N_4412,N_4544);
nand U4723 (N_4723,N_4518,N_4563);
nor U4724 (N_4724,N_4597,N_4569);
or U4725 (N_4725,N_4410,N_4434);
nor U4726 (N_4726,N_4408,N_4443);
nand U4727 (N_4727,N_4416,N_4543);
nand U4728 (N_4728,N_4498,N_4476);
xnor U4729 (N_4729,N_4552,N_4415);
and U4730 (N_4730,N_4563,N_4521);
or U4731 (N_4731,N_4545,N_4403);
and U4732 (N_4732,N_4507,N_4567);
and U4733 (N_4733,N_4435,N_4559);
nand U4734 (N_4734,N_4589,N_4438);
nand U4735 (N_4735,N_4499,N_4595);
nor U4736 (N_4736,N_4599,N_4597);
nand U4737 (N_4737,N_4545,N_4437);
or U4738 (N_4738,N_4543,N_4402);
or U4739 (N_4739,N_4566,N_4498);
xnor U4740 (N_4740,N_4509,N_4564);
nor U4741 (N_4741,N_4437,N_4424);
and U4742 (N_4742,N_4509,N_4414);
and U4743 (N_4743,N_4503,N_4457);
and U4744 (N_4744,N_4470,N_4434);
nor U4745 (N_4745,N_4584,N_4512);
and U4746 (N_4746,N_4566,N_4486);
or U4747 (N_4747,N_4467,N_4566);
or U4748 (N_4748,N_4549,N_4537);
and U4749 (N_4749,N_4436,N_4519);
nor U4750 (N_4750,N_4449,N_4538);
xor U4751 (N_4751,N_4575,N_4536);
xor U4752 (N_4752,N_4552,N_4496);
nor U4753 (N_4753,N_4435,N_4599);
nand U4754 (N_4754,N_4548,N_4413);
xor U4755 (N_4755,N_4545,N_4401);
nor U4756 (N_4756,N_4490,N_4502);
nand U4757 (N_4757,N_4437,N_4568);
nor U4758 (N_4758,N_4578,N_4597);
xor U4759 (N_4759,N_4439,N_4470);
xor U4760 (N_4760,N_4535,N_4465);
or U4761 (N_4761,N_4465,N_4482);
and U4762 (N_4762,N_4458,N_4444);
nor U4763 (N_4763,N_4479,N_4500);
or U4764 (N_4764,N_4413,N_4443);
xor U4765 (N_4765,N_4537,N_4530);
xnor U4766 (N_4766,N_4527,N_4422);
and U4767 (N_4767,N_4563,N_4552);
xor U4768 (N_4768,N_4584,N_4521);
xor U4769 (N_4769,N_4574,N_4529);
nor U4770 (N_4770,N_4403,N_4436);
nand U4771 (N_4771,N_4565,N_4561);
or U4772 (N_4772,N_4468,N_4544);
or U4773 (N_4773,N_4536,N_4485);
nand U4774 (N_4774,N_4426,N_4454);
and U4775 (N_4775,N_4426,N_4467);
and U4776 (N_4776,N_4427,N_4501);
nor U4777 (N_4777,N_4409,N_4416);
xor U4778 (N_4778,N_4557,N_4462);
nand U4779 (N_4779,N_4487,N_4458);
xnor U4780 (N_4780,N_4431,N_4490);
and U4781 (N_4781,N_4481,N_4489);
nor U4782 (N_4782,N_4409,N_4509);
and U4783 (N_4783,N_4523,N_4583);
xnor U4784 (N_4784,N_4587,N_4473);
and U4785 (N_4785,N_4570,N_4401);
nor U4786 (N_4786,N_4511,N_4510);
or U4787 (N_4787,N_4556,N_4475);
nor U4788 (N_4788,N_4447,N_4434);
xnor U4789 (N_4789,N_4492,N_4476);
xor U4790 (N_4790,N_4499,N_4566);
and U4791 (N_4791,N_4562,N_4492);
nor U4792 (N_4792,N_4585,N_4511);
and U4793 (N_4793,N_4586,N_4450);
or U4794 (N_4794,N_4583,N_4494);
xor U4795 (N_4795,N_4595,N_4548);
or U4796 (N_4796,N_4554,N_4456);
nand U4797 (N_4797,N_4541,N_4476);
xnor U4798 (N_4798,N_4446,N_4569);
nand U4799 (N_4799,N_4510,N_4556);
and U4800 (N_4800,N_4697,N_4688);
nand U4801 (N_4801,N_4728,N_4671);
nand U4802 (N_4802,N_4749,N_4785);
or U4803 (N_4803,N_4776,N_4730);
and U4804 (N_4804,N_4608,N_4726);
nand U4805 (N_4805,N_4631,N_4638);
nor U4806 (N_4806,N_4692,N_4680);
nor U4807 (N_4807,N_4780,N_4754);
or U4808 (N_4808,N_4629,N_4746);
nor U4809 (N_4809,N_4743,N_4771);
and U4810 (N_4810,N_4712,N_4691);
nor U4811 (N_4811,N_4601,N_4705);
or U4812 (N_4812,N_4700,N_4751);
and U4813 (N_4813,N_4741,N_4791);
xnor U4814 (N_4814,N_4663,N_4618);
nand U4815 (N_4815,N_4759,N_4625);
and U4816 (N_4816,N_4725,N_4717);
nor U4817 (N_4817,N_4645,N_4723);
nand U4818 (N_4818,N_4769,N_4687);
nand U4819 (N_4819,N_4610,N_4650);
xor U4820 (N_4820,N_4626,N_4753);
nand U4821 (N_4821,N_4799,N_4624);
or U4822 (N_4822,N_4774,N_4742);
xor U4823 (N_4823,N_4651,N_4659);
nor U4824 (N_4824,N_4768,N_4789);
nand U4825 (N_4825,N_4729,N_4731);
xor U4826 (N_4826,N_4744,N_4613);
or U4827 (N_4827,N_4736,N_4701);
or U4828 (N_4828,N_4648,N_4611);
and U4829 (N_4829,N_4739,N_4628);
and U4830 (N_4830,N_4672,N_4644);
and U4831 (N_4831,N_4636,N_4615);
nand U4832 (N_4832,N_4675,N_4747);
nor U4833 (N_4833,N_4679,N_4604);
or U4834 (N_4834,N_4661,N_4653);
and U4835 (N_4835,N_4662,N_4765);
nor U4836 (N_4836,N_4737,N_4766);
or U4837 (N_4837,N_4681,N_4665);
nand U4838 (N_4838,N_4654,N_4715);
or U4839 (N_4839,N_4640,N_4655);
nor U4840 (N_4840,N_4642,N_4673);
xnor U4841 (N_4841,N_4708,N_4770);
nor U4842 (N_4842,N_4732,N_4738);
xnor U4843 (N_4843,N_4707,N_4760);
and U4844 (N_4844,N_4616,N_4790);
nor U4845 (N_4845,N_4600,N_4699);
or U4846 (N_4846,N_4720,N_4632);
nand U4847 (N_4847,N_4722,N_4750);
nor U4848 (N_4848,N_4693,N_4762);
nand U4849 (N_4849,N_4639,N_4706);
and U4850 (N_4850,N_4676,N_4761);
or U4851 (N_4851,N_4781,N_4678);
xnor U4852 (N_4852,N_4779,N_4740);
xnor U4853 (N_4853,N_4714,N_4668);
or U4854 (N_4854,N_4764,N_4683);
or U4855 (N_4855,N_4758,N_4724);
or U4856 (N_4856,N_4657,N_4633);
xor U4857 (N_4857,N_4627,N_4694);
nand U4858 (N_4858,N_4710,N_4772);
nor U4859 (N_4859,N_4652,N_4656);
and U4860 (N_4860,N_4685,N_4614);
or U4861 (N_4861,N_4670,N_4703);
and U4862 (N_4862,N_4649,N_4718);
xnor U4863 (N_4863,N_4775,N_4612);
and U4864 (N_4864,N_4794,N_4621);
xnor U4865 (N_4865,N_4646,N_4788);
or U4866 (N_4866,N_4660,N_4745);
or U4867 (N_4867,N_4606,N_4734);
or U4868 (N_4868,N_4719,N_4696);
or U4869 (N_4869,N_4637,N_4634);
xnor U4870 (N_4870,N_4795,N_4698);
nor U4871 (N_4871,N_4686,N_4674);
nor U4872 (N_4872,N_4622,N_4617);
and U4873 (N_4873,N_4689,N_4793);
or U4874 (N_4874,N_4620,N_4778);
nand U4875 (N_4875,N_4666,N_4798);
and U4876 (N_4876,N_4786,N_4630);
nand U4877 (N_4877,N_4647,N_4603);
xor U4878 (N_4878,N_4641,N_4767);
nand U4879 (N_4879,N_4607,N_4635);
nand U4880 (N_4880,N_4784,N_4721);
or U4881 (N_4881,N_4755,N_4716);
and U4882 (N_4882,N_4727,N_4664);
nand U4883 (N_4883,N_4704,N_4602);
xnor U4884 (N_4884,N_4792,N_4609);
xnor U4885 (N_4885,N_4763,N_4684);
nor U4886 (N_4886,N_4619,N_4796);
and U4887 (N_4887,N_4643,N_4682);
nor U4888 (N_4888,N_4690,N_4777);
xor U4889 (N_4889,N_4773,N_4658);
or U4890 (N_4890,N_4733,N_4709);
and U4891 (N_4891,N_4757,N_4677);
nand U4892 (N_4892,N_4735,N_4711);
and U4893 (N_4893,N_4787,N_4702);
xor U4894 (N_4894,N_4797,N_4748);
xnor U4895 (N_4895,N_4605,N_4713);
nor U4896 (N_4896,N_4756,N_4669);
nor U4897 (N_4897,N_4667,N_4623);
nor U4898 (N_4898,N_4695,N_4752);
nor U4899 (N_4899,N_4782,N_4783);
or U4900 (N_4900,N_4767,N_4662);
and U4901 (N_4901,N_4658,N_4683);
nand U4902 (N_4902,N_4700,N_4672);
nand U4903 (N_4903,N_4660,N_4778);
or U4904 (N_4904,N_4611,N_4605);
nor U4905 (N_4905,N_4654,N_4618);
or U4906 (N_4906,N_4629,N_4663);
and U4907 (N_4907,N_4704,N_4616);
and U4908 (N_4908,N_4621,N_4763);
or U4909 (N_4909,N_4738,N_4691);
nor U4910 (N_4910,N_4721,N_4728);
nor U4911 (N_4911,N_4661,N_4659);
xor U4912 (N_4912,N_4648,N_4602);
or U4913 (N_4913,N_4735,N_4661);
nor U4914 (N_4914,N_4720,N_4645);
or U4915 (N_4915,N_4677,N_4649);
and U4916 (N_4916,N_4606,N_4723);
or U4917 (N_4917,N_4770,N_4790);
nor U4918 (N_4918,N_4686,N_4796);
nor U4919 (N_4919,N_4605,N_4650);
and U4920 (N_4920,N_4610,N_4749);
or U4921 (N_4921,N_4686,N_4780);
nor U4922 (N_4922,N_4630,N_4734);
or U4923 (N_4923,N_4642,N_4795);
nand U4924 (N_4924,N_4715,N_4716);
or U4925 (N_4925,N_4765,N_4627);
and U4926 (N_4926,N_4631,N_4633);
and U4927 (N_4927,N_4645,N_4722);
nand U4928 (N_4928,N_4630,N_4650);
xor U4929 (N_4929,N_4789,N_4748);
and U4930 (N_4930,N_4698,N_4674);
nand U4931 (N_4931,N_4683,N_4708);
or U4932 (N_4932,N_4781,N_4733);
nor U4933 (N_4933,N_4637,N_4703);
nor U4934 (N_4934,N_4662,N_4774);
nand U4935 (N_4935,N_4678,N_4789);
xnor U4936 (N_4936,N_4747,N_4698);
or U4937 (N_4937,N_4699,N_4660);
nor U4938 (N_4938,N_4640,N_4741);
nand U4939 (N_4939,N_4616,N_4614);
or U4940 (N_4940,N_4703,N_4649);
xnor U4941 (N_4941,N_4778,N_4738);
nor U4942 (N_4942,N_4776,N_4787);
nand U4943 (N_4943,N_4685,N_4768);
and U4944 (N_4944,N_4693,N_4741);
nor U4945 (N_4945,N_4751,N_4674);
nor U4946 (N_4946,N_4602,N_4696);
or U4947 (N_4947,N_4643,N_4606);
xor U4948 (N_4948,N_4603,N_4740);
nand U4949 (N_4949,N_4736,N_4713);
xnor U4950 (N_4950,N_4747,N_4633);
nor U4951 (N_4951,N_4633,N_4628);
nand U4952 (N_4952,N_4690,N_4614);
or U4953 (N_4953,N_4678,N_4600);
nor U4954 (N_4954,N_4657,N_4709);
and U4955 (N_4955,N_4797,N_4698);
and U4956 (N_4956,N_4605,N_4733);
nand U4957 (N_4957,N_4768,N_4653);
or U4958 (N_4958,N_4713,N_4677);
nand U4959 (N_4959,N_4789,N_4742);
xor U4960 (N_4960,N_4752,N_4633);
or U4961 (N_4961,N_4611,N_4731);
and U4962 (N_4962,N_4652,N_4600);
xnor U4963 (N_4963,N_4617,N_4738);
or U4964 (N_4964,N_4725,N_4653);
or U4965 (N_4965,N_4715,N_4660);
nor U4966 (N_4966,N_4651,N_4686);
xnor U4967 (N_4967,N_4745,N_4680);
and U4968 (N_4968,N_4695,N_4716);
or U4969 (N_4969,N_4795,N_4736);
and U4970 (N_4970,N_4719,N_4738);
nor U4971 (N_4971,N_4703,N_4699);
nand U4972 (N_4972,N_4668,N_4774);
and U4973 (N_4973,N_4782,N_4754);
nand U4974 (N_4974,N_4616,N_4620);
or U4975 (N_4975,N_4739,N_4713);
nand U4976 (N_4976,N_4792,N_4741);
and U4977 (N_4977,N_4797,N_4763);
or U4978 (N_4978,N_4688,N_4731);
nor U4979 (N_4979,N_4669,N_4622);
xnor U4980 (N_4980,N_4682,N_4766);
xnor U4981 (N_4981,N_4699,N_4792);
nand U4982 (N_4982,N_4772,N_4730);
xnor U4983 (N_4983,N_4637,N_4650);
nand U4984 (N_4984,N_4729,N_4634);
nor U4985 (N_4985,N_4645,N_4673);
nand U4986 (N_4986,N_4609,N_4614);
xnor U4987 (N_4987,N_4682,N_4741);
or U4988 (N_4988,N_4778,N_4748);
or U4989 (N_4989,N_4693,N_4606);
nor U4990 (N_4990,N_4636,N_4709);
or U4991 (N_4991,N_4679,N_4780);
or U4992 (N_4992,N_4709,N_4646);
nor U4993 (N_4993,N_4603,N_4668);
xor U4994 (N_4994,N_4684,N_4783);
nor U4995 (N_4995,N_4769,N_4637);
or U4996 (N_4996,N_4761,N_4673);
and U4997 (N_4997,N_4767,N_4778);
xnor U4998 (N_4998,N_4676,N_4623);
nor U4999 (N_4999,N_4783,N_4693);
nand U5000 (N_5000,N_4919,N_4869);
nor U5001 (N_5001,N_4997,N_4942);
and U5002 (N_5002,N_4828,N_4809);
nor U5003 (N_5003,N_4978,N_4885);
nor U5004 (N_5004,N_4975,N_4848);
and U5005 (N_5005,N_4909,N_4887);
or U5006 (N_5006,N_4812,N_4999);
and U5007 (N_5007,N_4871,N_4946);
and U5008 (N_5008,N_4807,N_4977);
and U5009 (N_5009,N_4853,N_4846);
xnor U5010 (N_5010,N_4882,N_4886);
nor U5011 (N_5011,N_4821,N_4910);
and U5012 (N_5012,N_4990,N_4966);
nand U5013 (N_5013,N_4849,N_4884);
and U5014 (N_5014,N_4923,N_4940);
nor U5015 (N_5015,N_4991,N_4870);
and U5016 (N_5016,N_4891,N_4862);
and U5017 (N_5017,N_4802,N_4931);
xor U5018 (N_5018,N_4974,N_4826);
or U5019 (N_5019,N_4947,N_4959);
nand U5020 (N_5020,N_4987,N_4850);
xnor U5021 (N_5021,N_4934,N_4903);
and U5022 (N_5022,N_4897,N_4936);
or U5023 (N_5023,N_4957,N_4958);
and U5024 (N_5024,N_4805,N_4803);
xor U5025 (N_5025,N_4981,N_4836);
nand U5026 (N_5026,N_4814,N_4833);
and U5027 (N_5027,N_4854,N_4816);
nand U5028 (N_5028,N_4955,N_4857);
nand U5029 (N_5029,N_4855,N_4835);
xor U5030 (N_5030,N_4939,N_4918);
nor U5031 (N_5031,N_4993,N_4844);
and U5032 (N_5032,N_4800,N_4830);
nand U5033 (N_5033,N_4874,N_4920);
nand U5034 (N_5034,N_4856,N_4900);
and U5035 (N_5035,N_4983,N_4930);
nor U5036 (N_5036,N_4824,N_4924);
or U5037 (N_5037,N_4944,N_4962);
and U5038 (N_5038,N_4861,N_4912);
or U5039 (N_5039,N_4817,N_4965);
and U5040 (N_5040,N_4894,N_4956);
nand U5041 (N_5041,N_4994,N_4938);
or U5042 (N_5042,N_4867,N_4852);
xor U5043 (N_5043,N_4928,N_4937);
or U5044 (N_5044,N_4951,N_4973);
nand U5045 (N_5045,N_4915,N_4960);
nand U5046 (N_5046,N_4950,N_4877);
or U5047 (N_5047,N_4980,N_4875);
xnor U5048 (N_5048,N_4841,N_4906);
nand U5049 (N_5049,N_4819,N_4898);
and U5050 (N_5050,N_4925,N_4829);
nand U5051 (N_5051,N_4893,N_4963);
nand U5052 (N_5052,N_4883,N_4842);
xor U5053 (N_5053,N_4995,N_4922);
nor U5054 (N_5054,N_4948,N_4851);
or U5055 (N_5055,N_4834,N_4899);
and U5056 (N_5056,N_4804,N_4982);
xnor U5057 (N_5057,N_4845,N_4902);
nand U5058 (N_5058,N_4970,N_4892);
and U5059 (N_5059,N_4913,N_4865);
and U5060 (N_5060,N_4878,N_4941);
nand U5061 (N_5061,N_4972,N_4864);
and U5062 (N_5062,N_4908,N_4801);
nand U5063 (N_5063,N_4843,N_4911);
xnor U5064 (N_5064,N_4866,N_4896);
nor U5065 (N_5065,N_4859,N_4811);
nor U5066 (N_5066,N_4823,N_4847);
or U5067 (N_5067,N_4929,N_4971);
nand U5068 (N_5068,N_4889,N_4901);
and U5069 (N_5069,N_4890,N_4808);
nor U5070 (N_5070,N_4917,N_4863);
nor U5071 (N_5071,N_4954,N_4822);
nand U5072 (N_5072,N_4933,N_4876);
nand U5073 (N_5073,N_4964,N_4907);
nand U5074 (N_5074,N_4888,N_4921);
xnor U5075 (N_5075,N_4806,N_4825);
and U5076 (N_5076,N_4953,N_4967);
xor U5077 (N_5077,N_4952,N_4820);
or U5078 (N_5078,N_4932,N_4813);
nor U5079 (N_5079,N_4989,N_4984);
or U5080 (N_5080,N_4992,N_4986);
nor U5081 (N_5081,N_4969,N_4914);
or U5082 (N_5082,N_4873,N_4839);
xnor U5083 (N_5083,N_4998,N_4927);
nand U5084 (N_5084,N_4880,N_4868);
nor U5085 (N_5085,N_4935,N_4815);
xnor U5086 (N_5086,N_4926,N_4943);
xor U5087 (N_5087,N_4985,N_4837);
or U5088 (N_5088,N_4976,N_4827);
nor U5089 (N_5089,N_4904,N_4949);
nor U5090 (N_5090,N_4945,N_4988);
or U5091 (N_5091,N_4832,N_4895);
and U5092 (N_5092,N_4881,N_4916);
or U5093 (N_5093,N_4831,N_4905);
nand U5094 (N_5094,N_4840,N_4996);
or U5095 (N_5095,N_4961,N_4838);
nand U5096 (N_5096,N_4879,N_4818);
xor U5097 (N_5097,N_4858,N_4810);
xor U5098 (N_5098,N_4860,N_4872);
and U5099 (N_5099,N_4979,N_4968);
nor U5100 (N_5100,N_4866,N_4922);
nor U5101 (N_5101,N_4934,N_4853);
or U5102 (N_5102,N_4826,N_4865);
nand U5103 (N_5103,N_4801,N_4999);
nor U5104 (N_5104,N_4995,N_4811);
xor U5105 (N_5105,N_4806,N_4854);
nor U5106 (N_5106,N_4811,N_4841);
nor U5107 (N_5107,N_4817,N_4885);
nand U5108 (N_5108,N_4937,N_4826);
and U5109 (N_5109,N_4823,N_4821);
xor U5110 (N_5110,N_4844,N_4841);
nor U5111 (N_5111,N_4892,N_4863);
and U5112 (N_5112,N_4924,N_4878);
and U5113 (N_5113,N_4891,N_4810);
and U5114 (N_5114,N_4984,N_4955);
and U5115 (N_5115,N_4986,N_4922);
nand U5116 (N_5116,N_4805,N_4962);
nand U5117 (N_5117,N_4836,N_4854);
nor U5118 (N_5118,N_4995,N_4831);
nand U5119 (N_5119,N_4903,N_4803);
nor U5120 (N_5120,N_4949,N_4950);
or U5121 (N_5121,N_4932,N_4962);
nand U5122 (N_5122,N_4999,N_4857);
xor U5123 (N_5123,N_4990,N_4956);
nor U5124 (N_5124,N_4996,N_4897);
or U5125 (N_5125,N_4933,N_4812);
nand U5126 (N_5126,N_4948,N_4938);
and U5127 (N_5127,N_4841,N_4897);
and U5128 (N_5128,N_4909,N_4962);
xnor U5129 (N_5129,N_4860,N_4985);
nor U5130 (N_5130,N_4866,N_4973);
nor U5131 (N_5131,N_4912,N_4830);
nor U5132 (N_5132,N_4916,N_4848);
nand U5133 (N_5133,N_4844,N_4963);
nor U5134 (N_5134,N_4859,N_4816);
xor U5135 (N_5135,N_4952,N_4973);
xnor U5136 (N_5136,N_4878,N_4930);
xor U5137 (N_5137,N_4882,N_4961);
nor U5138 (N_5138,N_4873,N_4899);
and U5139 (N_5139,N_4815,N_4880);
or U5140 (N_5140,N_4834,N_4877);
nand U5141 (N_5141,N_4830,N_4996);
and U5142 (N_5142,N_4993,N_4882);
nand U5143 (N_5143,N_4967,N_4889);
and U5144 (N_5144,N_4991,N_4921);
xnor U5145 (N_5145,N_4927,N_4871);
or U5146 (N_5146,N_4928,N_4939);
nor U5147 (N_5147,N_4829,N_4906);
nor U5148 (N_5148,N_4964,N_4801);
or U5149 (N_5149,N_4922,N_4902);
xnor U5150 (N_5150,N_4943,N_4993);
and U5151 (N_5151,N_4824,N_4861);
nand U5152 (N_5152,N_4897,N_4817);
nand U5153 (N_5153,N_4930,N_4836);
xor U5154 (N_5154,N_4935,N_4952);
and U5155 (N_5155,N_4883,N_4869);
nand U5156 (N_5156,N_4849,N_4906);
or U5157 (N_5157,N_4834,N_4964);
and U5158 (N_5158,N_4843,N_4960);
or U5159 (N_5159,N_4932,N_4886);
nand U5160 (N_5160,N_4840,N_4898);
or U5161 (N_5161,N_4918,N_4808);
or U5162 (N_5162,N_4965,N_4973);
and U5163 (N_5163,N_4894,N_4880);
nor U5164 (N_5164,N_4923,N_4952);
and U5165 (N_5165,N_4814,N_4907);
or U5166 (N_5166,N_4940,N_4917);
xor U5167 (N_5167,N_4887,N_4839);
or U5168 (N_5168,N_4904,N_4973);
or U5169 (N_5169,N_4947,N_4988);
xnor U5170 (N_5170,N_4959,N_4902);
and U5171 (N_5171,N_4928,N_4992);
xnor U5172 (N_5172,N_4910,N_4888);
and U5173 (N_5173,N_4875,N_4910);
xnor U5174 (N_5174,N_4847,N_4959);
nor U5175 (N_5175,N_4844,N_4905);
xor U5176 (N_5176,N_4828,N_4940);
and U5177 (N_5177,N_4959,N_4849);
nor U5178 (N_5178,N_4870,N_4915);
xnor U5179 (N_5179,N_4924,N_4998);
or U5180 (N_5180,N_4963,N_4978);
nor U5181 (N_5181,N_4803,N_4934);
xnor U5182 (N_5182,N_4887,N_4970);
and U5183 (N_5183,N_4946,N_4867);
and U5184 (N_5184,N_4800,N_4975);
or U5185 (N_5185,N_4822,N_4873);
nand U5186 (N_5186,N_4967,N_4810);
or U5187 (N_5187,N_4829,N_4822);
nor U5188 (N_5188,N_4838,N_4888);
and U5189 (N_5189,N_4974,N_4959);
and U5190 (N_5190,N_4880,N_4916);
nand U5191 (N_5191,N_4858,N_4975);
nor U5192 (N_5192,N_4832,N_4899);
and U5193 (N_5193,N_4956,N_4947);
nor U5194 (N_5194,N_4811,N_4838);
nor U5195 (N_5195,N_4995,N_4844);
nor U5196 (N_5196,N_4947,N_4968);
or U5197 (N_5197,N_4839,N_4978);
nor U5198 (N_5198,N_4879,N_4920);
or U5199 (N_5199,N_4858,N_4958);
xor U5200 (N_5200,N_5004,N_5049);
and U5201 (N_5201,N_5198,N_5027);
and U5202 (N_5202,N_5103,N_5006);
and U5203 (N_5203,N_5130,N_5119);
and U5204 (N_5204,N_5191,N_5142);
or U5205 (N_5205,N_5154,N_5120);
nor U5206 (N_5206,N_5044,N_5149);
nor U5207 (N_5207,N_5177,N_5180);
nor U5208 (N_5208,N_5188,N_5164);
xnor U5209 (N_5209,N_5094,N_5173);
xor U5210 (N_5210,N_5045,N_5152);
or U5211 (N_5211,N_5012,N_5139);
nor U5212 (N_5212,N_5126,N_5058);
nor U5213 (N_5213,N_5144,N_5076);
nor U5214 (N_5214,N_5023,N_5155);
nand U5215 (N_5215,N_5011,N_5035);
or U5216 (N_5216,N_5010,N_5143);
nor U5217 (N_5217,N_5092,N_5059);
nor U5218 (N_5218,N_5100,N_5088);
xor U5219 (N_5219,N_5079,N_5145);
and U5220 (N_5220,N_5042,N_5082);
xor U5221 (N_5221,N_5160,N_5156);
and U5222 (N_5222,N_5068,N_5161);
or U5223 (N_5223,N_5115,N_5029);
or U5224 (N_5224,N_5072,N_5026);
or U5225 (N_5225,N_5040,N_5159);
and U5226 (N_5226,N_5034,N_5195);
xor U5227 (N_5227,N_5112,N_5106);
or U5228 (N_5228,N_5007,N_5081);
nand U5229 (N_5229,N_5107,N_5056);
xor U5230 (N_5230,N_5157,N_5066);
nand U5231 (N_5231,N_5168,N_5001);
nand U5232 (N_5232,N_5124,N_5117);
nand U5233 (N_5233,N_5170,N_5002);
or U5234 (N_5234,N_5057,N_5074);
xnor U5235 (N_5235,N_5053,N_5038);
nand U5236 (N_5236,N_5105,N_5122);
xnor U5237 (N_5237,N_5102,N_5169);
nor U5238 (N_5238,N_5048,N_5151);
nor U5239 (N_5239,N_5129,N_5089);
and U5240 (N_5240,N_5118,N_5185);
xnor U5241 (N_5241,N_5025,N_5109);
xor U5242 (N_5242,N_5099,N_5189);
nor U5243 (N_5243,N_5197,N_5005);
nor U5244 (N_5244,N_5146,N_5033);
xor U5245 (N_5245,N_5186,N_5137);
or U5246 (N_5246,N_5178,N_5015);
xor U5247 (N_5247,N_5054,N_5070);
nor U5248 (N_5248,N_5047,N_5116);
nor U5249 (N_5249,N_5075,N_5014);
or U5250 (N_5250,N_5138,N_5181);
nor U5251 (N_5251,N_5016,N_5060);
nor U5252 (N_5252,N_5008,N_5064);
and U5253 (N_5253,N_5017,N_5046);
nand U5254 (N_5254,N_5135,N_5021);
xnor U5255 (N_5255,N_5093,N_5071);
or U5256 (N_5256,N_5020,N_5077);
nor U5257 (N_5257,N_5018,N_5073);
nor U5258 (N_5258,N_5065,N_5087);
xnor U5259 (N_5259,N_5184,N_5167);
nor U5260 (N_5260,N_5111,N_5132);
and U5261 (N_5261,N_5183,N_5104);
xnor U5262 (N_5262,N_5061,N_5078);
xnor U5263 (N_5263,N_5096,N_5091);
nor U5264 (N_5264,N_5192,N_5024);
nand U5265 (N_5265,N_5063,N_5147);
nor U5266 (N_5266,N_5069,N_5171);
xnor U5267 (N_5267,N_5086,N_5030);
xnor U5268 (N_5268,N_5028,N_5190);
nand U5269 (N_5269,N_5003,N_5113);
nor U5270 (N_5270,N_5141,N_5041);
or U5271 (N_5271,N_5085,N_5114);
and U5272 (N_5272,N_5127,N_5176);
nand U5273 (N_5273,N_5162,N_5163);
xor U5274 (N_5274,N_5019,N_5150);
nand U5275 (N_5275,N_5080,N_5052);
nand U5276 (N_5276,N_5037,N_5174);
xnor U5277 (N_5277,N_5062,N_5194);
nor U5278 (N_5278,N_5199,N_5187);
xnor U5279 (N_5279,N_5172,N_5051);
nor U5280 (N_5280,N_5136,N_5153);
xor U5281 (N_5281,N_5097,N_5165);
nor U5282 (N_5282,N_5140,N_5179);
nor U5283 (N_5283,N_5133,N_5083);
or U5284 (N_5284,N_5050,N_5110);
nor U5285 (N_5285,N_5108,N_5134);
xor U5286 (N_5286,N_5022,N_5193);
and U5287 (N_5287,N_5196,N_5121);
xor U5288 (N_5288,N_5101,N_5084);
and U5289 (N_5289,N_5067,N_5158);
xor U5290 (N_5290,N_5175,N_5095);
and U5291 (N_5291,N_5125,N_5039);
nor U5292 (N_5292,N_5090,N_5098);
and U5293 (N_5293,N_5031,N_5043);
and U5294 (N_5294,N_5148,N_5182);
xor U5295 (N_5295,N_5123,N_5000);
nor U5296 (N_5296,N_5009,N_5128);
nand U5297 (N_5297,N_5131,N_5036);
and U5298 (N_5298,N_5032,N_5166);
and U5299 (N_5299,N_5055,N_5013);
nor U5300 (N_5300,N_5187,N_5094);
nand U5301 (N_5301,N_5045,N_5151);
xnor U5302 (N_5302,N_5153,N_5008);
nand U5303 (N_5303,N_5082,N_5134);
and U5304 (N_5304,N_5174,N_5156);
and U5305 (N_5305,N_5092,N_5120);
xnor U5306 (N_5306,N_5061,N_5025);
xor U5307 (N_5307,N_5166,N_5043);
xnor U5308 (N_5308,N_5025,N_5191);
nor U5309 (N_5309,N_5093,N_5169);
nor U5310 (N_5310,N_5038,N_5089);
and U5311 (N_5311,N_5123,N_5026);
or U5312 (N_5312,N_5150,N_5107);
nand U5313 (N_5313,N_5166,N_5142);
xnor U5314 (N_5314,N_5127,N_5088);
nand U5315 (N_5315,N_5000,N_5144);
and U5316 (N_5316,N_5105,N_5119);
nor U5317 (N_5317,N_5153,N_5150);
or U5318 (N_5318,N_5003,N_5166);
or U5319 (N_5319,N_5001,N_5011);
nor U5320 (N_5320,N_5086,N_5099);
nor U5321 (N_5321,N_5096,N_5165);
nor U5322 (N_5322,N_5049,N_5008);
xor U5323 (N_5323,N_5082,N_5074);
nand U5324 (N_5324,N_5133,N_5080);
nor U5325 (N_5325,N_5152,N_5138);
xnor U5326 (N_5326,N_5153,N_5148);
or U5327 (N_5327,N_5003,N_5120);
nor U5328 (N_5328,N_5050,N_5004);
xnor U5329 (N_5329,N_5005,N_5155);
and U5330 (N_5330,N_5006,N_5197);
xnor U5331 (N_5331,N_5035,N_5097);
nor U5332 (N_5332,N_5101,N_5111);
nor U5333 (N_5333,N_5186,N_5055);
or U5334 (N_5334,N_5011,N_5039);
nor U5335 (N_5335,N_5139,N_5019);
or U5336 (N_5336,N_5193,N_5017);
or U5337 (N_5337,N_5074,N_5178);
or U5338 (N_5338,N_5181,N_5111);
or U5339 (N_5339,N_5085,N_5148);
nor U5340 (N_5340,N_5169,N_5056);
or U5341 (N_5341,N_5149,N_5074);
xor U5342 (N_5342,N_5082,N_5050);
and U5343 (N_5343,N_5019,N_5015);
or U5344 (N_5344,N_5094,N_5022);
nand U5345 (N_5345,N_5007,N_5168);
or U5346 (N_5346,N_5075,N_5016);
nor U5347 (N_5347,N_5186,N_5078);
nor U5348 (N_5348,N_5139,N_5178);
nor U5349 (N_5349,N_5177,N_5023);
and U5350 (N_5350,N_5022,N_5109);
nand U5351 (N_5351,N_5001,N_5193);
nor U5352 (N_5352,N_5117,N_5055);
nand U5353 (N_5353,N_5148,N_5140);
and U5354 (N_5354,N_5041,N_5026);
and U5355 (N_5355,N_5020,N_5125);
nand U5356 (N_5356,N_5146,N_5040);
nor U5357 (N_5357,N_5195,N_5179);
or U5358 (N_5358,N_5050,N_5182);
nand U5359 (N_5359,N_5074,N_5069);
or U5360 (N_5360,N_5086,N_5143);
nand U5361 (N_5361,N_5078,N_5085);
nand U5362 (N_5362,N_5176,N_5168);
nand U5363 (N_5363,N_5070,N_5161);
and U5364 (N_5364,N_5035,N_5079);
xnor U5365 (N_5365,N_5051,N_5063);
nor U5366 (N_5366,N_5073,N_5150);
and U5367 (N_5367,N_5079,N_5183);
nor U5368 (N_5368,N_5147,N_5022);
nand U5369 (N_5369,N_5116,N_5146);
xnor U5370 (N_5370,N_5030,N_5049);
or U5371 (N_5371,N_5183,N_5094);
nor U5372 (N_5372,N_5013,N_5146);
nor U5373 (N_5373,N_5064,N_5196);
xor U5374 (N_5374,N_5008,N_5074);
nand U5375 (N_5375,N_5149,N_5073);
and U5376 (N_5376,N_5169,N_5058);
or U5377 (N_5377,N_5081,N_5085);
nand U5378 (N_5378,N_5198,N_5055);
xnor U5379 (N_5379,N_5035,N_5163);
nand U5380 (N_5380,N_5152,N_5125);
nand U5381 (N_5381,N_5017,N_5124);
or U5382 (N_5382,N_5017,N_5106);
and U5383 (N_5383,N_5142,N_5160);
nor U5384 (N_5384,N_5035,N_5159);
and U5385 (N_5385,N_5104,N_5185);
nand U5386 (N_5386,N_5131,N_5076);
or U5387 (N_5387,N_5017,N_5026);
nor U5388 (N_5388,N_5130,N_5053);
xor U5389 (N_5389,N_5023,N_5070);
nor U5390 (N_5390,N_5116,N_5015);
nand U5391 (N_5391,N_5065,N_5059);
and U5392 (N_5392,N_5016,N_5174);
or U5393 (N_5393,N_5193,N_5150);
and U5394 (N_5394,N_5020,N_5101);
nor U5395 (N_5395,N_5055,N_5065);
nor U5396 (N_5396,N_5070,N_5132);
or U5397 (N_5397,N_5082,N_5193);
or U5398 (N_5398,N_5160,N_5118);
nor U5399 (N_5399,N_5025,N_5009);
xor U5400 (N_5400,N_5331,N_5217);
xor U5401 (N_5401,N_5255,N_5336);
and U5402 (N_5402,N_5385,N_5275);
xnor U5403 (N_5403,N_5349,N_5202);
or U5404 (N_5404,N_5313,N_5243);
xor U5405 (N_5405,N_5271,N_5329);
and U5406 (N_5406,N_5317,N_5338);
nand U5407 (N_5407,N_5264,N_5396);
and U5408 (N_5408,N_5382,N_5220);
and U5409 (N_5409,N_5263,N_5237);
and U5410 (N_5410,N_5397,N_5280);
nor U5411 (N_5411,N_5326,N_5210);
nor U5412 (N_5412,N_5303,N_5286);
or U5413 (N_5413,N_5290,N_5278);
nand U5414 (N_5414,N_5228,N_5344);
or U5415 (N_5415,N_5309,N_5352);
nand U5416 (N_5416,N_5376,N_5388);
or U5417 (N_5417,N_5249,N_5330);
or U5418 (N_5418,N_5318,N_5325);
or U5419 (N_5419,N_5253,N_5219);
and U5420 (N_5420,N_5339,N_5244);
nor U5421 (N_5421,N_5347,N_5387);
nand U5422 (N_5422,N_5372,N_5240);
and U5423 (N_5423,N_5308,N_5273);
xor U5424 (N_5424,N_5301,N_5306);
nor U5425 (N_5425,N_5322,N_5393);
xor U5426 (N_5426,N_5236,N_5356);
nand U5427 (N_5427,N_5213,N_5223);
and U5428 (N_5428,N_5248,N_5321);
and U5429 (N_5429,N_5204,N_5399);
xnor U5430 (N_5430,N_5239,N_5386);
or U5431 (N_5431,N_5283,N_5246);
and U5432 (N_5432,N_5231,N_5335);
xnor U5433 (N_5433,N_5390,N_5394);
nand U5434 (N_5434,N_5207,N_5353);
and U5435 (N_5435,N_5293,N_5320);
or U5436 (N_5436,N_5374,N_5368);
xnor U5437 (N_5437,N_5297,N_5222);
xor U5438 (N_5438,N_5341,N_5337);
and U5439 (N_5439,N_5367,N_5380);
and U5440 (N_5440,N_5365,N_5302);
nand U5441 (N_5441,N_5216,N_5312);
nor U5442 (N_5442,N_5235,N_5226);
or U5443 (N_5443,N_5241,N_5319);
xnor U5444 (N_5444,N_5373,N_5360);
nor U5445 (N_5445,N_5208,N_5245);
xor U5446 (N_5446,N_5268,N_5211);
nor U5447 (N_5447,N_5332,N_5295);
and U5448 (N_5448,N_5291,N_5389);
xor U5449 (N_5449,N_5259,N_5221);
nand U5450 (N_5450,N_5247,N_5257);
nand U5451 (N_5451,N_5392,N_5258);
xnor U5452 (N_5452,N_5272,N_5334);
and U5453 (N_5453,N_5375,N_5285);
nor U5454 (N_5454,N_5277,N_5311);
xor U5455 (N_5455,N_5296,N_5370);
xnor U5456 (N_5456,N_5215,N_5357);
or U5457 (N_5457,N_5232,N_5371);
xnor U5458 (N_5458,N_5307,N_5355);
or U5459 (N_5459,N_5284,N_5354);
nand U5460 (N_5460,N_5242,N_5267);
nor U5461 (N_5461,N_5252,N_5254);
nand U5462 (N_5462,N_5324,N_5261);
nand U5463 (N_5463,N_5340,N_5206);
nand U5464 (N_5464,N_5205,N_5304);
nor U5465 (N_5465,N_5310,N_5230);
nor U5466 (N_5466,N_5305,N_5315);
or U5467 (N_5467,N_5351,N_5209);
and U5468 (N_5468,N_5233,N_5381);
xnor U5469 (N_5469,N_5395,N_5391);
xnor U5470 (N_5470,N_5281,N_5377);
nor U5471 (N_5471,N_5250,N_5266);
xor U5472 (N_5472,N_5287,N_5270);
xor U5473 (N_5473,N_5214,N_5298);
xnor U5474 (N_5474,N_5260,N_5346);
and U5475 (N_5475,N_5225,N_5362);
xor U5476 (N_5476,N_5358,N_5279);
and U5477 (N_5477,N_5292,N_5369);
nor U5478 (N_5478,N_5363,N_5229);
and U5479 (N_5479,N_5359,N_5316);
xor U5480 (N_5480,N_5224,N_5276);
nand U5481 (N_5481,N_5348,N_5342);
nor U5482 (N_5482,N_5203,N_5345);
nand U5483 (N_5483,N_5384,N_5256);
or U5484 (N_5484,N_5333,N_5265);
xnor U5485 (N_5485,N_5282,N_5300);
nor U5486 (N_5486,N_5398,N_5227);
or U5487 (N_5487,N_5288,N_5274);
nand U5488 (N_5488,N_5294,N_5201);
and U5489 (N_5489,N_5200,N_5251);
xnor U5490 (N_5490,N_5323,N_5327);
nand U5491 (N_5491,N_5269,N_5378);
nor U5492 (N_5492,N_5262,N_5238);
or U5493 (N_5493,N_5366,N_5328);
nor U5494 (N_5494,N_5383,N_5314);
xnor U5495 (N_5495,N_5364,N_5361);
or U5496 (N_5496,N_5234,N_5299);
nand U5497 (N_5497,N_5289,N_5350);
nor U5498 (N_5498,N_5212,N_5218);
and U5499 (N_5499,N_5343,N_5379);
nor U5500 (N_5500,N_5260,N_5374);
or U5501 (N_5501,N_5239,N_5228);
nor U5502 (N_5502,N_5272,N_5211);
nand U5503 (N_5503,N_5352,N_5236);
nand U5504 (N_5504,N_5355,N_5200);
and U5505 (N_5505,N_5233,N_5218);
nor U5506 (N_5506,N_5301,N_5223);
nand U5507 (N_5507,N_5398,N_5243);
xnor U5508 (N_5508,N_5291,N_5358);
or U5509 (N_5509,N_5327,N_5217);
and U5510 (N_5510,N_5328,N_5277);
xnor U5511 (N_5511,N_5233,N_5223);
nand U5512 (N_5512,N_5229,N_5391);
nand U5513 (N_5513,N_5285,N_5342);
and U5514 (N_5514,N_5280,N_5360);
xnor U5515 (N_5515,N_5208,N_5298);
or U5516 (N_5516,N_5314,N_5280);
nor U5517 (N_5517,N_5270,N_5304);
nand U5518 (N_5518,N_5290,N_5284);
and U5519 (N_5519,N_5237,N_5334);
nor U5520 (N_5520,N_5216,N_5351);
xor U5521 (N_5521,N_5346,N_5247);
nand U5522 (N_5522,N_5206,N_5246);
and U5523 (N_5523,N_5208,N_5340);
nand U5524 (N_5524,N_5222,N_5255);
xor U5525 (N_5525,N_5369,N_5340);
or U5526 (N_5526,N_5361,N_5242);
and U5527 (N_5527,N_5366,N_5320);
and U5528 (N_5528,N_5323,N_5314);
or U5529 (N_5529,N_5203,N_5296);
or U5530 (N_5530,N_5272,N_5259);
nand U5531 (N_5531,N_5392,N_5389);
nand U5532 (N_5532,N_5298,N_5212);
nand U5533 (N_5533,N_5262,N_5244);
nand U5534 (N_5534,N_5201,N_5386);
nand U5535 (N_5535,N_5335,N_5274);
xnor U5536 (N_5536,N_5352,N_5319);
nor U5537 (N_5537,N_5334,N_5274);
and U5538 (N_5538,N_5344,N_5307);
and U5539 (N_5539,N_5363,N_5323);
and U5540 (N_5540,N_5240,N_5226);
xnor U5541 (N_5541,N_5226,N_5232);
or U5542 (N_5542,N_5276,N_5271);
xnor U5543 (N_5543,N_5348,N_5341);
xor U5544 (N_5544,N_5385,N_5220);
nor U5545 (N_5545,N_5217,N_5223);
and U5546 (N_5546,N_5297,N_5379);
xor U5547 (N_5547,N_5350,N_5294);
or U5548 (N_5548,N_5327,N_5306);
and U5549 (N_5549,N_5223,N_5369);
or U5550 (N_5550,N_5392,N_5380);
nor U5551 (N_5551,N_5352,N_5202);
or U5552 (N_5552,N_5201,N_5317);
nor U5553 (N_5553,N_5318,N_5315);
nor U5554 (N_5554,N_5272,N_5247);
nor U5555 (N_5555,N_5211,N_5365);
nand U5556 (N_5556,N_5368,N_5210);
or U5557 (N_5557,N_5211,N_5287);
and U5558 (N_5558,N_5319,N_5215);
nor U5559 (N_5559,N_5382,N_5285);
and U5560 (N_5560,N_5366,N_5236);
nand U5561 (N_5561,N_5231,N_5310);
nand U5562 (N_5562,N_5278,N_5374);
nor U5563 (N_5563,N_5398,N_5213);
xnor U5564 (N_5564,N_5394,N_5329);
nand U5565 (N_5565,N_5296,N_5386);
and U5566 (N_5566,N_5201,N_5336);
or U5567 (N_5567,N_5272,N_5386);
nand U5568 (N_5568,N_5378,N_5310);
or U5569 (N_5569,N_5319,N_5367);
and U5570 (N_5570,N_5299,N_5290);
nand U5571 (N_5571,N_5288,N_5340);
nor U5572 (N_5572,N_5364,N_5399);
xor U5573 (N_5573,N_5255,N_5308);
nand U5574 (N_5574,N_5322,N_5218);
nand U5575 (N_5575,N_5301,N_5226);
xnor U5576 (N_5576,N_5343,N_5387);
xor U5577 (N_5577,N_5226,N_5375);
and U5578 (N_5578,N_5338,N_5282);
xnor U5579 (N_5579,N_5383,N_5267);
nor U5580 (N_5580,N_5256,N_5348);
or U5581 (N_5581,N_5229,N_5372);
nand U5582 (N_5582,N_5378,N_5238);
xor U5583 (N_5583,N_5340,N_5308);
xnor U5584 (N_5584,N_5274,N_5325);
nand U5585 (N_5585,N_5356,N_5201);
nand U5586 (N_5586,N_5208,N_5389);
and U5587 (N_5587,N_5235,N_5309);
nor U5588 (N_5588,N_5380,N_5251);
nand U5589 (N_5589,N_5353,N_5289);
xnor U5590 (N_5590,N_5248,N_5282);
nor U5591 (N_5591,N_5322,N_5247);
nor U5592 (N_5592,N_5354,N_5359);
xor U5593 (N_5593,N_5344,N_5230);
nor U5594 (N_5594,N_5344,N_5396);
and U5595 (N_5595,N_5205,N_5347);
xor U5596 (N_5596,N_5344,N_5350);
or U5597 (N_5597,N_5369,N_5327);
or U5598 (N_5598,N_5206,N_5290);
nand U5599 (N_5599,N_5276,N_5372);
or U5600 (N_5600,N_5507,N_5453);
or U5601 (N_5601,N_5598,N_5491);
or U5602 (N_5602,N_5422,N_5436);
nor U5603 (N_5603,N_5532,N_5538);
nor U5604 (N_5604,N_5466,N_5499);
and U5605 (N_5605,N_5469,N_5533);
or U5606 (N_5606,N_5480,N_5597);
and U5607 (N_5607,N_5564,N_5400);
or U5608 (N_5608,N_5555,N_5575);
nor U5609 (N_5609,N_5461,N_5467);
or U5610 (N_5610,N_5582,N_5410);
nand U5611 (N_5611,N_5585,N_5589);
and U5612 (N_5612,N_5421,N_5593);
nor U5613 (N_5613,N_5528,N_5581);
and U5614 (N_5614,N_5441,N_5475);
nand U5615 (N_5615,N_5402,N_5500);
nor U5616 (N_5616,N_5526,N_5543);
xor U5617 (N_5617,N_5444,N_5541);
or U5618 (N_5618,N_5508,N_5463);
or U5619 (N_5619,N_5503,N_5470);
xnor U5620 (N_5620,N_5591,N_5485);
xnor U5621 (N_5621,N_5456,N_5445);
xnor U5622 (N_5622,N_5553,N_5434);
nand U5623 (N_5623,N_5449,N_5407);
nand U5624 (N_5624,N_5588,N_5476);
or U5625 (N_5625,N_5473,N_5529);
nand U5626 (N_5626,N_5552,N_5557);
nor U5627 (N_5627,N_5403,N_5540);
xnor U5628 (N_5628,N_5587,N_5450);
or U5629 (N_5629,N_5418,N_5559);
xor U5630 (N_5630,N_5596,N_5539);
and U5631 (N_5631,N_5415,N_5512);
nand U5632 (N_5632,N_5516,N_5545);
nand U5633 (N_5633,N_5416,N_5537);
and U5634 (N_5634,N_5405,N_5431);
xnor U5635 (N_5635,N_5519,N_5595);
and U5636 (N_5636,N_5464,N_5550);
or U5637 (N_5637,N_5566,N_5429);
xnor U5638 (N_5638,N_5574,N_5411);
and U5639 (N_5639,N_5440,N_5478);
nor U5640 (N_5640,N_5572,N_5556);
and U5641 (N_5641,N_5542,N_5447);
or U5642 (N_5642,N_5510,N_5413);
xor U5643 (N_5643,N_5535,N_5577);
and U5644 (N_5644,N_5497,N_5534);
nand U5645 (N_5645,N_5546,N_5462);
or U5646 (N_5646,N_5455,N_5571);
nor U5647 (N_5647,N_5511,N_5548);
nor U5648 (N_5648,N_5487,N_5570);
nor U5649 (N_5649,N_5412,N_5567);
and U5650 (N_5650,N_5496,N_5425);
xnor U5651 (N_5651,N_5518,N_5417);
nand U5652 (N_5652,N_5494,N_5408);
and U5653 (N_5653,N_5486,N_5439);
and U5654 (N_5654,N_5424,N_5560);
nand U5655 (N_5655,N_5515,N_5506);
nor U5656 (N_5656,N_5406,N_5452);
and U5657 (N_5657,N_5520,N_5472);
nand U5658 (N_5658,N_5594,N_5592);
nor U5659 (N_5659,N_5590,N_5427);
or U5660 (N_5660,N_5465,N_5525);
and U5661 (N_5661,N_5547,N_5471);
xor U5662 (N_5662,N_5523,N_5563);
nor U5663 (N_5663,N_5554,N_5583);
xnor U5664 (N_5664,N_5562,N_5514);
and U5665 (N_5665,N_5423,N_5432);
nand U5666 (N_5666,N_5544,N_5505);
xnor U5667 (N_5667,N_5568,N_5457);
nand U5668 (N_5668,N_5451,N_5443);
nor U5669 (N_5669,N_5458,N_5483);
nand U5670 (N_5670,N_5437,N_5504);
and U5671 (N_5671,N_5488,N_5414);
nand U5672 (N_5672,N_5409,N_5576);
xor U5673 (N_5673,N_5502,N_5565);
xnor U5674 (N_5674,N_5419,N_5580);
xor U5675 (N_5675,N_5561,N_5477);
xor U5676 (N_5676,N_5481,N_5448);
and U5677 (N_5677,N_5435,N_5549);
nand U5678 (N_5678,N_5558,N_5530);
xor U5679 (N_5679,N_5426,N_5482);
nand U5680 (N_5680,N_5438,N_5484);
xnor U5681 (N_5681,N_5586,N_5579);
xor U5682 (N_5682,N_5501,N_5513);
xor U5683 (N_5683,N_5527,N_5401);
nor U5684 (N_5684,N_5569,N_5430);
or U5685 (N_5685,N_5493,N_5433);
or U5686 (N_5686,N_5404,N_5536);
or U5687 (N_5687,N_5420,N_5442);
nand U5688 (N_5688,N_5517,N_5459);
nor U5689 (N_5689,N_5489,N_5468);
xor U5690 (N_5690,N_5495,N_5492);
xor U5691 (N_5691,N_5460,N_5521);
nor U5692 (N_5692,N_5551,N_5524);
xnor U5693 (N_5693,N_5474,N_5454);
nor U5694 (N_5694,N_5498,N_5599);
nor U5695 (N_5695,N_5509,N_5490);
or U5696 (N_5696,N_5578,N_5531);
xnor U5697 (N_5697,N_5428,N_5479);
xor U5698 (N_5698,N_5446,N_5584);
nand U5699 (N_5699,N_5522,N_5573);
or U5700 (N_5700,N_5471,N_5560);
or U5701 (N_5701,N_5458,N_5536);
or U5702 (N_5702,N_5444,N_5554);
nor U5703 (N_5703,N_5563,N_5540);
xor U5704 (N_5704,N_5542,N_5412);
xnor U5705 (N_5705,N_5565,N_5548);
and U5706 (N_5706,N_5411,N_5571);
xnor U5707 (N_5707,N_5592,N_5473);
nand U5708 (N_5708,N_5445,N_5401);
nor U5709 (N_5709,N_5445,N_5433);
xnor U5710 (N_5710,N_5578,N_5586);
nand U5711 (N_5711,N_5447,N_5585);
nor U5712 (N_5712,N_5594,N_5436);
nand U5713 (N_5713,N_5521,N_5420);
xnor U5714 (N_5714,N_5444,N_5480);
xnor U5715 (N_5715,N_5512,N_5476);
nor U5716 (N_5716,N_5591,N_5598);
nand U5717 (N_5717,N_5583,N_5502);
or U5718 (N_5718,N_5453,N_5557);
nor U5719 (N_5719,N_5541,N_5593);
nor U5720 (N_5720,N_5523,N_5491);
xnor U5721 (N_5721,N_5481,N_5549);
nand U5722 (N_5722,N_5460,N_5402);
and U5723 (N_5723,N_5413,N_5523);
nor U5724 (N_5724,N_5438,N_5580);
nor U5725 (N_5725,N_5480,N_5502);
nand U5726 (N_5726,N_5477,N_5426);
nand U5727 (N_5727,N_5552,N_5598);
and U5728 (N_5728,N_5568,N_5430);
nor U5729 (N_5729,N_5559,N_5582);
xnor U5730 (N_5730,N_5503,N_5428);
xnor U5731 (N_5731,N_5592,N_5430);
nand U5732 (N_5732,N_5565,N_5569);
or U5733 (N_5733,N_5594,N_5584);
xnor U5734 (N_5734,N_5551,N_5469);
nor U5735 (N_5735,N_5547,N_5506);
xnor U5736 (N_5736,N_5543,N_5556);
and U5737 (N_5737,N_5490,N_5568);
or U5738 (N_5738,N_5534,N_5459);
or U5739 (N_5739,N_5493,N_5568);
xnor U5740 (N_5740,N_5482,N_5464);
or U5741 (N_5741,N_5559,N_5566);
nor U5742 (N_5742,N_5437,N_5584);
xor U5743 (N_5743,N_5428,N_5520);
xnor U5744 (N_5744,N_5564,N_5539);
xor U5745 (N_5745,N_5510,N_5588);
and U5746 (N_5746,N_5564,N_5591);
nor U5747 (N_5747,N_5534,N_5557);
and U5748 (N_5748,N_5587,N_5445);
or U5749 (N_5749,N_5538,N_5442);
xnor U5750 (N_5750,N_5523,N_5415);
nand U5751 (N_5751,N_5423,N_5424);
xor U5752 (N_5752,N_5477,N_5410);
xor U5753 (N_5753,N_5438,N_5514);
nor U5754 (N_5754,N_5540,N_5454);
xor U5755 (N_5755,N_5472,N_5548);
and U5756 (N_5756,N_5546,N_5518);
or U5757 (N_5757,N_5580,N_5477);
or U5758 (N_5758,N_5506,N_5400);
xnor U5759 (N_5759,N_5544,N_5430);
xor U5760 (N_5760,N_5552,N_5415);
and U5761 (N_5761,N_5556,N_5510);
and U5762 (N_5762,N_5402,N_5422);
nor U5763 (N_5763,N_5571,N_5538);
xor U5764 (N_5764,N_5476,N_5418);
and U5765 (N_5765,N_5496,N_5540);
and U5766 (N_5766,N_5491,N_5562);
and U5767 (N_5767,N_5445,N_5493);
and U5768 (N_5768,N_5498,N_5470);
or U5769 (N_5769,N_5418,N_5469);
and U5770 (N_5770,N_5502,N_5596);
xor U5771 (N_5771,N_5469,N_5548);
and U5772 (N_5772,N_5580,N_5467);
xor U5773 (N_5773,N_5534,N_5568);
nand U5774 (N_5774,N_5557,N_5577);
nor U5775 (N_5775,N_5479,N_5531);
xnor U5776 (N_5776,N_5549,N_5536);
or U5777 (N_5777,N_5494,N_5540);
or U5778 (N_5778,N_5447,N_5473);
nand U5779 (N_5779,N_5578,N_5414);
and U5780 (N_5780,N_5537,N_5430);
and U5781 (N_5781,N_5466,N_5498);
nand U5782 (N_5782,N_5400,N_5544);
and U5783 (N_5783,N_5581,N_5566);
xor U5784 (N_5784,N_5589,N_5409);
nand U5785 (N_5785,N_5521,N_5471);
and U5786 (N_5786,N_5474,N_5584);
nor U5787 (N_5787,N_5436,N_5514);
xnor U5788 (N_5788,N_5582,N_5427);
or U5789 (N_5789,N_5435,N_5468);
xnor U5790 (N_5790,N_5580,N_5521);
and U5791 (N_5791,N_5531,N_5498);
or U5792 (N_5792,N_5595,N_5576);
nor U5793 (N_5793,N_5535,N_5597);
nor U5794 (N_5794,N_5479,N_5518);
nand U5795 (N_5795,N_5420,N_5507);
or U5796 (N_5796,N_5573,N_5455);
xnor U5797 (N_5797,N_5421,N_5484);
or U5798 (N_5798,N_5405,N_5529);
xor U5799 (N_5799,N_5405,N_5471);
nand U5800 (N_5800,N_5682,N_5769);
and U5801 (N_5801,N_5702,N_5652);
nor U5802 (N_5802,N_5725,N_5608);
and U5803 (N_5803,N_5627,N_5718);
and U5804 (N_5804,N_5756,N_5700);
nor U5805 (N_5805,N_5614,N_5721);
xor U5806 (N_5806,N_5602,N_5775);
and U5807 (N_5807,N_5643,N_5778);
or U5808 (N_5808,N_5696,N_5678);
nand U5809 (N_5809,N_5737,N_5656);
nand U5810 (N_5810,N_5748,N_5707);
or U5811 (N_5811,N_5600,N_5792);
nor U5812 (N_5812,N_5771,N_5704);
or U5813 (N_5813,N_5781,N_5716);
or U5814 (N_5814,N_5669,N_5697);
or U5815 (N_5815,N_5635,N_5606);
nor U5816 (N_5816,N_5670,N_5685);
nor U5817 (N_5817,N_5663,N_5710);
nor U5818 (N_5818,N_5651,N_5699);
and U5819 (N_5819,N_5615,N_5644);
nand U5820 (N_5820,N_5621,N_5717);
xor U5821 (N_5821,N_5705,N_5640);
xor U5822 (N_5822,N_5776,N_5610);
or U5823 (N_5823,N_5679,N_5609);
xnor U5824 (N_5824,N_5730,N_5754);
and U5825 (N_5825,N_5658,N_5783);
xor U5826 (N_5826,N_5750,N_5698);
and U5827 (N_5827,N_5795,N_5654);
nand U5828 (N_5828,N_5642,N_5623);
and U5829 (N_5829,N_5741,N_5787);
xnor U5830 (N_5830,N_5605,N_5745);
xnor U5831 (N_5831,N_5728,N_5601);
nor U5832 (N_5832,N_5770,N_5779);
nand U5833 (N_5833,N_5733,N_5645);
or U5834 (N_5834,N_5767,N_5744);
xnor U5835 (N_5835,N_5758,N_5726);
nor U5836 (N_5836,N_5793,N_5731);
nand U5837 (N_5837,N_5780,N_5641);
nand U5838 (N_5838,N_5631,N_5648);
or U5839 (N_5839,N_5701,N_5712);
xnor U5840 (N_5840,N_5613,N_5671);
nor U5841 (N_5841,N_5759,N_5666);
nand U5842 (N_5842,N_5788,N_5639);
xnor U5843 (N_5843,N_5743,N_5740);
nand U5844 (N_5844,N_5749,N_5739);
xor U5845 (N_5845,N_5636,N_5761);
xor U5846 (N_5846,N_5691,N_5607);
nand U5847 (N_5847,N_5680,N_5768);
xnor U5848 (N_5848,N_5791,N_5638);
nand U5849 (N_5849,N_5676,N_5664);
nand U5850 (N_5850,N_5729,N_5720);
or U5851 (N_5851,N_5634,N_5777);
and U5852 (N_5852,N_5647,N_5684);
nand U5853 (N_5853,N_5675,N_5687);
nor U5854 (N_5854,N_5611,N_5723);
nor U5855 (N_5855,N_5622,N_5624);
and U5856 (N_5856,N_5708,N_5694);
nor U5857 (N_5857,N_5766,N_5603);
and U5858 (N_5858,N_5774,N_5785);
nand U5859 (N_5859,N_5646,N_5796);
nand U5860 (N_5860,N_5747,N_5703);
nand U5861 (N_5861,N_5690,N_5667);
or U5862 (N_5862,N_5661,N_5757);
or U5863 (N_5863,N_5765,N_5753);
or U5864 (N_5864,N_5713,N_5668);
or U5865 (N_5865,N_5752,N_5604);
xnor U5866 (N_5866,N_5689,N_5715);
or U5867 (N_5867,N_5782,N_5673);
and U5868 (N_5868,N_5714,N_5738);
nor U5869 (N_5869,N_5786,N_5709);
nand U5870 (N_5870,N_5798,N_5612);
and U5871 (N_5871,N_5653,N_5706);
and U5872 (N_5872,N_5616,N_5626);
and U5873 (N_5873,N_5762,N_5732);
nor U5874 (N_5874,N_5736,N_5688);
nor U5875 (N_5875,N_5764,N_5784);
nand U5876 (N_5876,N_5649,N_5772);
nor U5877 (N_5877,N_5751,N_5677);
xnor U5878 (N_5878,N_5790,N_5693);
nor U5879 (N_5879,N_5794,N_5650);
or U5880 (N_5880,N_5799,N_5742);
and U5881 (N_5881,N_5657,N_5695);
nor U5882 (N_5882,N_5659,N_5630);
or U5883 (N_5883,N_5618,N_5672);
nand U5884 (N_5884,N_5625,N_5797);
xnor U5885 (N_5885,N_5619,N_5665);
and U5886 (N_5886,N_5746,N_5662);
nand U5887 (N_5887,N_5617,N_5789);
or U5888 (N_5888,N_5674,N_5719);
nand U5889 (N_5889,N_5722,N_5633);
nand U5890 (N_5890,N_5763,N_5760);
or U5891 (N_5891,N_5735,N_5655);
and U5892 (N_5892,N_5620,N_5660);
xnor U5893 (N_5893,N_5681,N_5711);
nand U5894 (N_5894,N_5724,N_5629);
xor U5895 (N_5895,N_5632,N_5692);
or U5896 (N_5896,N_5683,N_5637);
or U5897 (N_5897,N_5686,N_5755);
nand U5898 (N_5898,N_5734,N_5628);
or U5899 (N_5899,N_5773,N_5727);
or U5900 (N_5900,N_5628,N_5687);
xor U5901 (N_5901,N_5678,N_5679);
and U5902 (N_5902,N_5751,N_5641);
nand U5903 (N_5903,N_5759,N_5638);
and U5904 (N_5904,N_5727,N_5708);
nor U5905 (N_5905,N_5771,N_5622);
or U5906 (N_5906,N_5636,N_5781);
nor U5907 (N_5907,N_5658,N_5713);
nand U5908 (N_5908,N_5748,N_5678);
nand U5909 (N_5909,N_5650,N_5637);
xnor U5910 (N_5910,N_5697,N_5612);
nand U5911 (N_5911,N_5705,N_5697);
or U5912 (N_5912,N_5623,N_5799);
or U5913 (N_5913,N_5719,N_5730);
or U5914 (N_5914,N_5755,N_5720);
and U5915 (N_5915,N_5625,N_5725);
nand U5916 (N_5916,N_5777,N_5778);
nand U5917 (N_5917,N_5639,N_5745);
and U5918 (N_5918,N_5666,N_5662);
and U5919 (N_5919,N_5710,N_5610);
and U5920 (N_5920,N_5719,N_5668);
or U5921 (N_5921,N_5779,N_5797);
xor U5922 (N_5922,N_5640,N_5635);
and U5923 (N_5923,N_5612,N_5793);
nor U5924 (N_5924,N_5777,N_5723);
nor U5925 (N_5925,N_5649,N_5792);
xnor U5926 (N_5926,N_5600,N_5695);
nor U5927 (N_5927,N_5763,N_5694);
xnor U5928 (N_5928,N_5751,N_5709);
xnor U5929 (N_5929,N_5604,N_5783);
xor U5930 (N_5930,N_5677,N_5680);
nor U5931 (N_5931,N_5605,N_5699);
or U5932 (N_5932,N_5635,N_5739);
or U5933 (N_5933,N_5633,N_5739);
xnor U5934 (N_5934,N_5769,N_5633);
and U5935 (N_5935,N_5642,N_5775);
nor U5936 (N_5936,N_5668,N_5757);
xnor U5937 (N_5937,N_5774,N_5715);
xor U5938 (N_5938,N_5630,N_5618);
nor U5939 (N_5939,N_5757,N_5751);
or U5940 (N_5940,N_5768,N_5657);
xor U5941 (N_5941,N_5642,N_5624);
xor U5942 (N_5942,N_5725,N_5782);
nand U5943 (N_5943,N_5761,N_5632);
or U5944 (N_5944,N_5742,N_5788);
or U5945 (N_5945,N_5619,N_5741);
nor U5946 (N_5946,N_5724,N_5726);
and U5947 (N_5947,N_5713,N_5728);
xor U5948 (N_5948,N_5704,N_5786);
and U5949 (N_5949,N_5699,N_5786);
and U5950 (N_5950,N_5608,N_5627);
xor U5951 (N_5951,N_5738,N_5615);
and U5952 (N_5952,N_5613,N_5765);
or U5953 (N_5953,N_5640,N_5724);
nand U5954 (N_5954,N_5730,N_5695);
nor U5955 (N_5955,N_5725,N_5667);
nor U5956 (N_5956,N_5742,N_5720);
nor U5957 (N_5957,N_5700,N_5707);
and U5958 (N_5958,N_5643,N_5711);
and U5959 (N_5959,N_5645,N_5727);
nor U5960 (N_5960,N_5671,N_5698);
and U5961 (N_5961,N_5741,N_5700);
nand U5962 (N_5962,N_5757,N_5789);
nor U5963 (N_5963,N_5708,N_5763);
xnor U5964 (N_5964,N_5645,N_5760);
xor U5965 (N_5965,N_5769,N_5621);
or U5966 (N_5966,N_5629,N_5689);
nand U5967 (N_5967,N_5689,N_5650);
nand U5968 (N_5968,N_5681,N_5716);
nand U5969 (N_5969,N_5753,N_5740);
nor U5970 (N_5970,N_5684,N_5771);
and U5971 (N_5971,N_5638,N_5695);
or U5972 (N_5972,N_5601,N_5784);
nor U5973 (N_5973,N_5718,N_5743);
and U5974 (N_5974,N_5707,N_5611);
nor U5975 (N_5975,N_5649,N_5710);
and U5976 (N_5976,N_5764,N_5628);
xor U5977 (N_5977,N_5613,N_5609);
or U5978 (N_5978,N_5647,N_5765);
and U5979 (N_5979,N_5631,N_5621);
nor U5980 (N_5980,N_5614,N_5734);
nand U5981 (N_5981,N_5645,N_5770);
and U5982 (N_5982,N_5638,N_5679);
and U5983 (N_5983,N_5634,N_5783);
and U5984 (N_5984,N_5641,N_5691);
and U5985 (N_5985,N_5723,N_5693);
or U5986 (N_5986,N_5680,N_5736);
or U5987 (N_5987,N_5746,N_5643);
nor U5988 (N_5988,N_5768,N_5777);
nor U5989 (N_5989,N_5728,N_5721);
nor U5990 (N_5990,N_5671,N_5652);
xnor U5991 (N_5991,N_5687,N_5737);
nor U5992 (N_5992,N_5613,N_5652);
nor U5993 (N_5993,N_5634,N_5698);
or U5994 (N_5994,N_5603,N_5671);
nor U5995 (N_5995,N_5678,N_5765);
xnor U5996 (N_5996,N_5755,N_5708);
xor U5997 (N_5997,N_5746,N_5724);
or U5998 (N_5998,N_5654,N_5791);
nand U5999 (N_5999,N_5619,N_5659);
xor U6000 (N_6000,N_5901,N_5931);
or U6001 (N_6001,N_5966,N_5974);
nor U6002 (N_6002,N_5911,N_5873);
xnor U6003 (N_6003,N_5929,N_5861);
and U6004 (N_6004,N_5835,N_5961);
nand U6005 (N_6005,N_5882,N_5913);
nor U6006 (N_6006,N_5833,N_5991);
nand U6007 (N_6007,N_5904,N_5927);
xnor U6008 (N_6008,N_5868,N_5806);
nand U6009 (N_6009,N_5887,N_5936);
nand U6010 (N_6010,N_5972,N_5847);
or U6011 (N_6011,N_5969,N_5889);
xnor U6012 (N_6012,N_5981,N_5978);
xnor U6013 (N_6013,N_5864,N_5823);
or U6014 (N_6014,N_5937,N_5954);
xnor U6015 (N_6015,N_5973,N_5917);
or U6016 (N_6016,N_5941,N_5896);
nand U6017 (N_6017,N_5858,N_5879);
or U6018 (N_6018,N_5866,N_5884);
nor U6019 (N_6019,N_5870,N_5925);
and U6020 (N_6020,N_5935,N_5869);
xnor U6021 (N_6021,N_5877,N_5965);
nor U6022 (N_6022,N_5957,N_5989);
or U6023 (N_6023,N_5865,N_5907);
or U6024 (N_6024,N_5976,N_5942);
and U6025 (N_6025,N_5977,N_5983);
or U6026 (N_6026,N_5830,N_5909);
or U6027 (N_6027,N_5919,N_5953);
and U6028 (N_6028,N_5853,N_5891);
and U6029 (N_6029,N_5899,N_5923);
and U6030 (N_6030,N_5808,N_5962);
or U6031 (N_6031,N_5897,N_5926);
nor U6032 (N_6032,N_5824,N_5809);
xor U6033 (N_6033,N_5968,N_5843);
or U6034 (N_6034,N_5836,N_5996);
nand U6035 (N_6035,N_5920,N_5863);
nand U6036 (N_6036,N_5924,N_5805);
or U6037 (N_6037,N_5902,N_5859);
nor U6038 (N_6038,N_5854,N_5867);
nand U6039 (N_6039,N_5855,N_5905);
and U6040 (N_6040,N_5993,N_5827);
or U6041 (N_6041,N_5938,N_5908);
nand U6042 (N_6042,N_5826,N_5828);
and U6043 (N_6043,N_5992,N_5852);
or U6044 (N_6044,N_5940,N_5845);
nand U6045 (N_6045,N_5850,N_5818);
xor U6046 (N_6046,N_5947,N_5811);
nand U6047 (N_6047,N_5825,N_5817);
nor U6048 (N_6048,N_5822,N_5888);
and U6049 (N_6049,N_5987,N_5807);
nor U6050 (N_6050,N_5930,N_5800);
and U6051 (N_6051,N_5918,N_5939);
nand U6052 (N_6052,N_5975,N_5890);
and U6053 (N_6053,N_5886,N_5812);
xor U6054 (N_6054,N_5837,N_5943);
nor U6055 (N_6055,N_5846,N_5810);
xnor U6056 (N_6056,N_5821,N_5802);
nor U6057 (N_6057,N_5814,N_5893);
nor U6058 (N_6058,N_5838,N_5898);
and U6059 (N_6059,N_5958,N_5963);
nand U6060 (N_6060,N_5834,N_5892);
xnor U6061 (N_6061,N_5832,N_5831);
nand U6062 (N_6062,N_5880,N_5872);
xnor U6063 (N_6063,N_5995,N_5955);
or U6064 (N_6064,N_5813,N_5900);
and U6065 (N_6065,N_5860,N_5819);
or U6066 (N_6066,N_5928,N_5840);
or U6067 (N_6067,N_5945,N_5804);
or U6068 (N_6068,N_5980,N_5932);
nand U6069 (N_6069,N_5914,N_5871);
or U6070 (N_6070,N_5998,N_5959);
and U6071 (N_6071,N_5949,N_5964);
and U6072 (N_6072,N_5994,N_5952);
nor U6073 (N_6073,N_5849,N_5951);
nor U6074 (N_6074,N_5856,N_5956);
nand U6075 (N_6075,N_5982,N_5944);
nand U6076 (N_6076,N_5997,N_5874);
and U6077 (N_6077,N_5971,N_5946);
nor U6078 (N_6078,N_5803,N_5876);
and U6079 (N_6079,N_5921,N_5934);
and U6080 (N_6080,N_5844,N_5839);
and U6081 (N_6081,N_5990,N_5829);
nor U6082 (N_6082,N_5875,N_5967);
xnor U6083 (N_6083,N_5895,N_5894);
nor U6084 (N_6084,N_5885,N_5979);
nor U6085 (N_6085,N_5842,N_5820);
nand U6086 (N_6086,N_5857,N_5916);
or U6087 (N_6087,N_5933,N_5906);
nor U6088 (N_6088,N_5816,N_5848);
or U6089 (N_6089,N_5878,N_5851);
nor U6090 (N_6090,N_5986,N_5985);
and U6091 (N_6091,N_5984,N_5915);
or U6092 (N_6092,N_5815,N_5841);
nor U6093 (N_6093,N_5922,N_5883);
xor U6094 (N_6094,N_5903,N_5912);
and U6095 (N_6095,N_5960,N_5999);
xor U6096 (N_6096,N_5948,N_5988);
nand U6097 (N_6097,N_5950,N_5881);
or U6098 (N_6098,N_5910,N_5862);
nor U6099 (N_6099,N_5801,N_5970);
and U6100 (N_6100,N_5910,N_5926);
nand U6101 (N_6101,N_5938,N_5916);
xnor U6102 (N_6102,N_5854,N_5897);
and U6103 (N_6103,N_5861,N_5990);
or U6104 (N_6104,N_5875,N_5933);
and U6105 (N_6105,N_5811,N_5992);
xor U6106 (N_6106,N_5844,N_5914);
xor U6107 (N_6107,N_5937,N_5889);
or U6108 (N_6108,N_5930,N_5860);
xor U6109 (N_6109,N_5863,N_5874);
or U6110 (N_6110,N_5907,N_5806);
and U6111 (N_6111,N_5986,N_5992);
and U6112 (N_6112,N_5964,N_5835);
nand U6113 (N_6113,N_5904,N_5807);
and U6114 (N_6114,N_5824,N_5963);
and U6115 (N_6115,N_5850,N_5990);
or U6116 (N_6116,N_5913,N_5918);
nor U6117 (N_6117,N_5949,N_5839);
nand U6118 (N_6118,N_5810,N_5903);
or U6119 (N_6119,N_5983,N_5905);
nor U6120 (N_6120,N_5926,N_5835);
or U6121 (N_6121,N_5968,N_5878);
nand U6122 (N_6122,N_5801,N_5992);
and U6123 (N_6123,N_5845,N_5865);
or U6124 (N_6124,N_5904,N_5967);
nor U6125 (N_6125,N_5917,N_5808);
nor U6126 (N_6126,N_5923,N_5916);
nand U6127 (N_6127,N_5816,N_5823);
nor U6128 (N_6128,N_5887,N_5909);
nor U6129 (N_6129,N_5995,N_5834);
and U6130 (N_6130,N_5881,N_5872);
nor U6131 (N_6131,N_5808,N_5902);
xor U6132 (N_6132,N_5967,N_5861);
and U6133 (N_6133,N_5958,N_5981);
nand U6134 (N_6134,N_5971,N_5905);
nand U6135 (N_6135,N_5953,N_5883);
xnor U6136 (N_6136,N_5949,N_5881);
nor U6137 (N_6137,N_5939,N_5854);
or U6138 (N_6138,N_5944,N_5821);
and U6139 (N_6139,N_5843,N_5972);
xor U6140 (N_6140,N_5921,N_5808);
nand U6141 (N_6141,N_5977,N_5882);
and U6142 (N_6142,N_5809,N_5800);
and U6143 (N_6143,N_5986,N_5825);
and U6144 (N_6144,N_5925,N_5944);
nand U6145 (N_6145,N_5929,N_5872);
nand U6146 (N_6146,N_5941,N_5860);
xor U6147 (N_6147,N_5801,N_5877);
nor U6148 (N_6148,N_5908,N_5801);
nand U6149 (N_6149,N_5892,N_5937);
nand U6150 (N_6150,N_5865,N_5893);
or U6151 (N_6151,N_5978,N_5912);
and U6152 (N_6152,N_5903,N_5995);
and U6153 (N_6153,N_5989,N_5931);
or U6154 (N_6154,N_5899,N_5948);
nand U6155 (N_6155,N_5936,N_5925);
or U6156 (N_6156,N_5848,N_5972);
and U6157 (N_6157,N_5802,N_5990);
xnor U6158 (N_6158,N_5988,N_5917);
or U6159 (N_6159,N_5992,N_5993);
nand U6160 (N_6160,N_5887,N_5876);
or U6161 (N_6161,N_5970,N_5916);
nand U6162 (N_6162,N_5869,N_5962);
nor U6163 (N_6163,N_5988,N_5893);
or U6164 (N_6164,N_5864,N_5863);
nand U6165 (N_6165,N_5822,N_5831);
xnor U6166 (N_6166,N_5846,N_5891);
xnor U6167 (N_6167,N_5862,N_5900);
or U6168 (N_6168,N_5956,N_5836);
and U6169 (N_6169,N_5997,N_5983);
or U6170 (N_6170,N_5833,N_5954);
and U6171 (N_6171,N_5867,N_5912);
and U6172 (N_6172,N_5837,N_5900);
nor U6173 (N_6173,N_5854,N_5816);
nand U6174 (N_6174,N_5892,N_5822);
and U6175 (N_6175,N_5858,N_5940);
nor U6176 (N_6176,N_5898,N_5862);
nand U6177 (N_6177,N_5828,N_5839);
nand U6178 (N_6178,N_5800,N_5945);
and U6179 (N_6179,N_5871,N_5999);
and U6180 (N_6180,N_5934,N_5800);
nand U6181 (N_6181,N_5802,N_5967);
nand U6182 (N_6182,N_5828,N_5976);
nor U6183 (N_6183,N_5931,N_5812);
nand U6184 (N_6184,N_5815,N_5802);
nor U6185 (N_6185,N_5827,N_5972);
xnor U6186 (N_6186,N_5817,N_5947);
or U6187 (N_6187,N_5804,N_5911);
or U6188 (N_6188,N_5987,N_5912);
nor U6189 (N_6189,N_5883,N_5983);
nor U6190 (N_6190,N_5843,N_5947);
xor U6191 (N_6191,N_5832,N_5974);
nor U6192 (N_6192,N_5990,N_5816);
or U6193 (N_6193,N_5950,N_5816);
or U6194 (N_6194,N_5822,N_5823);
or U6195 (N_6195,N_5841,N_5990);
xor U6196 (N_6196,N_5971,N_5910);
nand U6197 (N_6197,N_5871,N_5837);
nand U6198 (N_6198,N_5887,N_5962);
or U6199 (N_6199,N_5984,N_5804);
nor U6200 (N_6200,N_6053,N_6184);
and U6201 (N_6201,N_6126,N_6006);
and U6202 (N_6202,N_6018,N_6056);
or U6203 (N_6203,N_6171,N_6091);
nand U6204 (N_6204,N_6048,N_6183);
or U6205 (N_6205,N_6119,N_6003);
xor U6206 (N_6206,N_6136,N_6108);
nor U6207 (N_6207,N_6031,N_6002);
and U6208 (N_6208,N_6137,N_6051);
xnor U6209 (N_6209,N_6081,N_6140);
nor U6210 (N_6210,N_6172,N_6030);
nand U6211 (N_6211,N_6079,N_6133);
nor U6212 (N_6212,N_6064,N_6050);
or U6213 (N_6213,N_6099,N_6161);
xnor U6214 (N_6214,N_6023,N_6042);
xor U6215 (N_6215,N_6092,N_6177);
xnor U6216 (N_6216,N_6004,N_6186);
or U6217 (N_6217,N_6089,N_6174);
xnor U6218 (N_6218,N_6038,N_6170);
or U6219 (N_6219,N_6077,N_6135);
nor U6220 (N_6220,N_6111,N_6168);
or U6221 (N_6221,N_6026,N_6090);
nor U6222 (N_6222,N_6097,N_6029);
nand U6223 (N_6223,N_6139,N_6132);
nor U6224 (N_6224,N_6117,N_6082);
xnor U6225 (N_6225,N_6134,N_6185);
and U6226 (N_6226,N_6063,N_6025);
xnor U6227 (N_6227,N_6076,N_6113);
or U6228 (N_6228,N_6046,N_6070);
nand U6229 (N_6229,N_6198,N_6193);
and U6230 (N_6230,N_6182,N_6014);
xnor U6231 (N_6231,N_6138,N_6028);
nand U6232 (N_6232,N_6034,N_6129);
and U6233 (N_6233,N_6098,N_6194);
and U6234 (N_6234,N_6153,N_6175);
nand U6235 (N_6235,N_6005,N_6061);
xnor U6236 (N_6236,N_6106,N_6187);
and U6237 (N_6237,N_6093,N_6158);
nand U6238 (N_6238,N_6104,N_6128);
nand U6239 (N_6239,N_6109,N_6159);
nor U6240 (N_6240,N_6027,N_6143);
or U6241 (N_6241,N_6007,N_6103);
nand U6242 (N_6242,N_6116,N_6197);
xor U6243 (N_6243,N_6024,N_6164);
or U6244 (N_6244,N_6039,N_6015);
xor U6245 (N_6245,N_6118,N_6189);
xnor U6246 (N_6246,N_6021,N_6037);
xnor U6247 (N_6247,N_6057,N_6012);
nand U6248 (N_6248,N_6072,N_6040);
or U6249 (N_6249,N_6087,N_6020);
nand U6250 (N_6250,N_6156,N_6120);
nor U6251 (N_6251,N_6150,N_6167);
xnor U6252 (N_6252,N_6062,N_6094);
xnor U6253 (N_6253,N_6009,N_6035);
nand U6254 (N_6254,N_6043,N_6149);
and U6255 (N_6255,N_6165,N_6065);
or U6256 (N_6256,N_6142,N_6122);
xnor U6257 (N_6257,N_6144,N_6086);
xnor U6258 (N_6258,N_6196,N_6127);
nand U6259 (N_6259,N_6071,N_6124);
or U6260 (N_6260,N_6083,N_6054);
and U6261 (N_6261,N_6017,N_6102);
and U6262 (N_6262,N_6188,N_6121);
nor U6263 (N_6263,N_6199,N_6178);
or U6264 (N_6264,N_6107,N_6131);
and U6265 (N_6265,N_6073,N_6075);
or U6266 (N_6266,N_6141,N_6096);
or U6267 (N_6267,N_6125,N_6151);
nor U6268 (N_6268,N_6045,N_6100);
nand U6269 (N_6269,N_6160,N_6080);
nor U6270 (N_6270,N_6154,N_6163);
nand U6271 (N_6271,N_6173,N_6032);
xnor U6272 (N_6272,N_6146,N_6105);
nand U6273 (N_6273,N_6145,N_6000);
and U6274 (N_6274,N_6008,N_6147);
or U6275 (N_6275,N_6180,N_6166);
or U6276 (N_6276,N_6049,N_6010);
xor U6277 (N_6277,N_6195,N_6190);
nand U6278 (N_6278,N_6036,N_6074);
nand U6279 (N_6279,N_6068,N_6066);
nand U6280 (N_6280,N_6157,N_6191);
or U6281 (N_6281,N_6192,N_6181);
nand U6282 (N_6282,N_6179,N_6041);
and U6283 (N_6283,N_6148,N_6176);
nor U6284 (N_6284,N_6085,N_6001);
xnor U6285 (N_6285,N_6011,N_6110);
or U6286 (N_6286,N_6016,N_6055);
nand U6287 (N_6287,N_6115,N_6152);
xnor U6288 (N_6288,N_6123,N_6013);
xnor U6289 (N_6289,N_6095,N_6130);
xnor U6290 (N_6290,N_6088,N_6047);
nand U6291 (N_6291,N_6162,N_6155);
xor U6292 (N_6292,N_6019,N_6069);
nor U6293 (N_6293,N_6058,N_6112);
nand U6294 (N_6294,N_6101,N_6114);
xnor U6295 (N_6295,N_6084,N_6052);
nand U6296 (N_6296,N_6044,N_6067);
xnor U6297 (N_6297,N_6022,N_6169);
xnor U6298 (N_6298,N_6059,N_6033);
nand U6299 (N_6299,N_6078,N_6060);
nand U6300 (N_6300,N_6076,N_6138);
nand U6301 (N_6301,N_6142,N_6160);
nor U6302 (N_6302,N_6040,N_6058);
or U6303 (N_6303,N_6193,N_6020);
or U6304 (N_6304,N_6164,N_6139);
and U6305 (N_6305,N_6126,N_6066);
xor U6306 (N_6306,N_6038,N_6025);
nor U6307 (N_6307,N_6148,N_6167);
or U6308 (N_6308,N_6199,N_6165);
and U6309 (N_6309,N_6128,N_6053);
nand U6310 (N_6310,N_6045,N_6187);
nor U6311 (N_6311,N_6175,N_6120);
or U6312 (N_6312,N_6077,N_6011);
xnor U6313 (N_6313,N_6192,N_6037);
or U6314 (N_6314,N_6148,N_6023);
nand U6315 (N_6315,N_6116,N_6013);
nand U6316 (N_6316,N_6174,N_6093);
nor U6317 (N_6317,N_6196,N_6195);
nor U6318 (N_6318,N_6124,N_6026);
xor U6319 (N_6319,N_6120,N_6003);
nor U6320 (N_6320,N_6012,N_6064);
nor U6321 (N_6321,N_6081,N_6040);
or U6322 (N_6322,N_6040,N_6005);
or U6323 (N_6323,N_6117,N_6109);
and U6324 (N_6324,N_6089,N_6027);
and U6325 (N_6325,N_6047,N_6181);
nand U6326 (N_6326,N_6139,N_6096);
and U6327 (N_6327,N_6165,N_6109);
and U6328 (N_6328,N_6010,N_6058);
and U6329 (N_6329,N_6198,N_6157);
and U6330 (N_6330,N_6011,N_6062);
or U6331 (N_6331,N_6049,N_6197);
nand U6332 (N_6332,N_6019,N_6107);
nand U6333 (N_6333,N_6146,N_6016);
nand U6334 (N_6334,N_6001,N_6186);
nand U6335 (N_6335,N_6112,N_6096);
xor U6336 (N_6336,N_6191,N_6020);
nor U6337 (N_6337,N_6124,N_6010);
nand U6338 (N_6338,N_6016,N_6113);
and U6339 (N_6339,N_6170,N_6174);
nand U6340 (N_6340,N_6024,N_6026);
nor U6341 (N_6341,N_6161,N_6046);
or U6342 (N_6342,N_6177,N_6062);
nand U6343 (N_6343,N_6043,N_6195);
nand U6344 (N_6344,N_6177,N_6168);
nand U6345 (N_6345,N_6183,N_6021);
xnor U6346 (N_6346,N_6043,N_6025);
nand U6347 (N_6347,N_6039,N_6124);
nand U6348 (N_6348,N_6019,N_6165);
xnor U6349 (N_6349,N_6100,N_6146);
and U6350 (N_6350,N_6189,N_6181);
or U6351 (N_6351,N_6176,N_6111);
and U6352 (N_6352,N_6104,N_6058);
xnor U6353 (N_6353,N_6142,N_6066);
nor U6354 (N_6354,N_6014,N_6194);
nand U6355 (N_6355,N_6057,N_6059);
or U6356 (N_6356,N_6191,N_6062);
xor U6357 (N_6357,N_6117,N_6065);
and U6358 (N_6358,N_6059,N_6090);
and U6359 (N_6359,N_6015,N_6094);
nor U6360 (N_6360,N_6126,N_6134);
or U6361 (N_6361,N_6187,N_6171);
nor U6362 (N_6362,N_6030,N_6193);
nand U6363 (N_6363,N_6165,N_6048);
or U6364 (N_6364,N_6157,N_6128);
nor U6365 (N_6365,N_6071,N_6084);
and U6366 (N_6366,N_6059,N_6010);
and U6367 (N_6367,N_6094,N_6111);
xnor U6368 (N_6368,N_6022,N_6162);
nor U6369 (N_6369,N_6163,N_6160);
nand U6370 (N_6370,N_6089,N_6135);
nand U6371 (N_6371,N_6105,N_6058);
or U6372 (N_6372,N_6189,N_6021);
nand U6373 (N_6373,N_6004,N_6108);
or U6374 (N_6374,N_6178,N_6089);
or U6375 (N_6375,N_6113,N_6047);
nor U6376 (N_6376,N_6041,N_6093);
or U6377 (N_6377,N_6053,N_6192);
nand U6378 (N_6378,N_6137,N_6022);
xor U6379 (N_6379,N_6005,N_6178);
nor U6380 (N_6380,N_6102,N_6012);
nor U6381 (N_6381,N_6196,N_6101);
nand U6382 (N_6382,N_6150,N_6023);
nand U6383 (N_6383,N_6109,N_6137);
and U6384 (N_6384,N_6174,N_6114);
nor U6385 (N_6385,N_6101,N_6124);
xor U6386 (N_6386,N_6087,N_6015);
or U6387 (N_6387,N_6077,N_6198);
nor U6388 (N_6388,N_6086,N_6096);
xnor U6389 (N_6389,N_6063,N_6170);
or U6390 (N_6390,N_6193,N_6035);
nand U6391 (N_6391,N_6038,N_6164);
and U6392 (N_6392,N_6011,N_6197);
or U6393 (N_6393,N_6198,N_6017);
nor U6394 (N_6394,N_6030,N_6165);
nand U6395 (N_6395,N_6038,N_6180);
or U6396 (N_6396,N_6193,N_6034);
nand U6397 (N_6397,N_6054,N_6112);
nand U6398 (N_6398,N_6131,N_6113);
xor U6399 (N_6399,N_6119,N_6125);
xnor U6400 (N_6400,N_6302,N_6261);
or U6401 (N_6401,N_6369,N_6202);
or U6402 (N_6402,N_6306,N_6255);
and U6403 (N_6403,N_6319,N_6381);
xor U6404 (N_6404,N_6392,N_6293);
and U6405 (N_6405,N_6216,N_6291);
and U6406 (N_6406,N_6226,N_6245);
and U6407 (N_6407,N_6361,N_6228);
or U6408 (N_6408,N_6259,N_6386);
and U6409 (N_6409,N_6263,N_6203);
or U6410 (N_6410,N_6320,N_6391);
or U6411 (N_6411,N_6348,N_6277);
or U6412 (N_6412,N_6266,N_6344);
nand U6413 (N_6413,N_6350,N_6242);
nand U6414 (N_6414,N_6214,N_6235);
nand U6415 (N_6415,N_6368,N_6327);
or U6416 (N_6416,N_6340,N_6229);
and U6417 (N_6417,N_6385,N_6333);
nor U6418 (N_6418,N_6337,N_6278);
and U6419 (N_6419,N_6231,N_6287);
xor U6420 (N_6420,N_6397,N_6311);
and U6421 (N_6421,N_6238,N_6268);
nand U6422 (N_6422,N_6281,N_6294);
or U6423 (N_6423,N_6222,N_6272);
xor U6424 (N_6424,N_6285,N_6209);
and U6425 (N_6425,N_6317,N_6328);
nand U6426 (N_6426,N_6276,N_6349);
and U6427 (N_6427,N_6233,N_6223);
nor U6428 (N_6428,N_6211,N_6345);
and U6429 (N_6429,N_6347,N_6398);
xnor U6430 (N_6430,N_6224,N_6356);
xnor U6431 (N_6431,N_6265,N_6352);
and U6432 (N_6432,N_6307,N_6256);
nand U6433 (N_6433,N_6269,N_6338);
nor U6434 (N_6434,N_6239,N_6325);
xnor U6435 (N_6435,N_6301,N_6336);
nand U6436 (N_6436,N_6341,N_6205);
xnor U6437 (N_6437,N_6243,N_6200);
xor U6438 (N_6438,N_6283,N_6364);
and U6439 (N_6439,N_6329,N_6219);
nand U6440 (N_6440,N_6258,N_6384);
and U6441 (N_6441,N_6217,N_6377);
nor U6442 (N_6442,N_6373,N_6279);
or U6443 (N_6443,N_6355,N_6395);
and U6444 (N_6444,N_6286,N_6370);
xnor U6445 (N_6445,N_6289,N_6305);
xor U6446 (N_6446,N_6346,N_6382);
nor U6447 (N_6447,N_6379,N_6322);
xnor U6448 (N_6448,N_6248,N_6383);
and U6449 (N_6449,N_6380,N_6339);
or U6450 (N_6450,N_6343,N_6376);
xor U6451 (N_6451,N_6378,N_6360);
or U6452 (N_6452,N_6252,N_6299);
xor U6453 (N_6453,N_6210,N_6247);
or U6454 (N_6454,N_6257,N_6253);
nand U6455 (N_6455,N_6246,N_6331);
and U6456 (N_6456,N_6249,N_6204);
xor U6457 (N_6457,N_6330,N_6351);
nor U6458 (N_6458,N_6357,N_6236);
and U6459 (N_6459,N_6365,N_6371);
nor U6460 (N_6460,N_6367,N_6375);
or U6461 (N_6461,N_6284,N_6334);
nand U6462 (N_6462,N_6318,N_6326);
xor U6463 (N_6463,N_6353,N_6300);
nand U6464 (N_6464,N_6332,N_6237);
nor U6465 (N_6465,N_6366,N_6267);
nand U6466 (N_6466,N_6354,N_6394);
and U6467 (N_6467,N_6264,N_6323);
nand U6468 (N_6468,N_6312,N_6359);
xnor U6469 (N_6469,N_6342,N_6251);
nand U6470 (N_6470,N_6372,N_6316);
xor U6471 (N_6471,N_6212,N_6273);
or U6472 (N_6472,N_6292,N_6315);
xnor U6473 (N_6473,N_6288,N_6215);
nor U6474 (N_6474,N_6389,N_6358);
nand U6475 (N_6475,N_6374,N_6262);
nand U6476 (N_6476,N_6310,N_6388);
or U6477 (N_6477,N_6321,N_6298);
and U6478 (N_6478,N_6390,N_6207);
xnor U6479 (N_6479,N_6201,N_6335);
and U6480 (N_6480,N_6206,N_6260);
xnor U6481 (N_6481,N_6297,N_6282);
nand U6482 (N_6482,N_6308,N_6314);
xor U6483 (N_6483,N_6254,N_6208);
nor U6484 (N_6484,N_6271,N_6244);
and U6485 (N_6485,N_6396,N_6303);
xor U6486 (N_6486,N_6240,N_6362);
and U6487 (N_6487,N_6280,N_6295);
nor U6488 (N_6488,N_6232,N_6220);
and U6489 (N_6489,N_6227,N_6221);
nand U6490 (N_6490,N_6309,N_6275);
nand U6491 (N_6491,N_6274,N_6324);
or U6492 (N_6492,N_6290,N_6241);
or U6493 (N_6493,N_6218,N_6387);
nand U6494 (N_6494,N_6363,N_6399);
xor U6495 (N_6495,N_6230,N_6296);
nor U6496 (N_6496,N_6393,N_6213);
nor U6497 (N_6497,N_6313,N_6250);
nor U6498 (N_6498,N_6304,N_6225);
xor U6499 (N_6499,N_6234,N_6270);
nand U6500 (N_6500,N_6321,N_6270);
nor U6501 (N_6501,N_6307,N_6346);
or U6502 (N_6502,N_6254,N_6222);
xnor U6503 (N_6503,N_6316,N_6391);
nor U6504 (N_6504,N_6347,N_6354);
xnor U6505 (N_6505,N_6373,N_6397);
and U6506 (N_6506,N_6281,N_6289);
and U6507 (N_6507,N_6288,N_6274);
and U6508 (N_6508,N_6239,N_6388);
xnor U6509 (N_6509,N_6360,N_6351);
nand U6510 (N_6510,N_6248,N_6313);
nand U6511 (N_6511,N_6305,N_6217);
nand U6512 (N_6512,N_6390,N_6238);
or U6513 (N_6513,N_6327,N_6282);
and U6514 (N_6514,N_6333,N_6276);
or U6515 (N_6515,N_6364,N_6230);
and U6516 (N_6516,N_6392,N_6251);
nor U6517 (N_6517,N_6280,N_6270);
or U6518 (N_6518,N_6379,N_6344);
nor U6519 (N_6519,N_6232,N_6240);
nor U6520 (N_6520,N_6348,N_6202);
nor U6521 (N_6521,N_6279,N_6359);
nor U6522 (N_6522,N_6362,N_6349);
and U6523 (N_6523,N_6291,N_6373);
nand U6524 (N_6524,N_6274,N_6229);
xnor U6525 (N_6525,N_6289,N_6359);
and U6526 (N_6526,N_6347,N_6240);
nand U6527 (N_6527,N_6286,N_6390);
nand U6528 (N_6528,N_6342,N_6289);
or U6529 (N_6529,N_6206,N_6387);
nor U6530 (N_6530,N_6239,N_6244);
or U6531 (N_6531,N_6311,N_6225);
and U6532 (N_6532,N_6342,N_6247);
or U6533 (N_6533,N_6380,N_6263);
xor U6534 (N_6534,N_6344,N_6372);
xor U6535 (N_6535,N_6316,N_6226);
nand U6536 (N_6536,N_6352,N_6306);
xnor U6537 (N_6537,N_6281,N_6362);
or U6538 (N_6538,N_6256,N_6203);
or U6539 (N_6539,N_6276,N_6208);
nand U6540 (N_6540,N_6308,N_6395);
or U6541 (N_6541,N_6277,N_6260);
nor U6542 (N_6542,N_6262,N_6289);
nand U6543 (N_6543,N_6294,N_6362);
nand U6544 (N_6544,N_6209,N_6224);
or U6545 (N_6545,N_6298,N_6344);
nand U6546 (N_6546,N_6390,N_6219);
and U6547 (N_6547,N_6223,N_6306);
nor U6548 (N_6548,N_6243,N_6363);
xnor U6549 (N_6549,N_6229,N_6368);
nand U6550 (N_6550,N_6219,N_6204);
nor U6551 (N_6551,N_6391,N_6259);
nand U6552 (N_6552,N_6214,N_6232);
xnor U6553 (N_6553,N_6347,N_6251);
and U6554 (N_6554,N_6259,N_6284);
nand U6555 (N_6555,N_6394,N_6280);
nand U6556 (N_6556,N_6332,N_6358);
nor U6557 (N_6557,N_6296,N_6308);
nand U6558 (N_6558,N_6389,N_6363);
nor U6559 (N_6559,N_6236,N_6284);
and U6560 (N_6560,N_6213,N_6370);
xnor U6561 (N_6561,N_6200,N_6210);
and U6562 (N_6562,N_6215,N_6341);
xnor U6563 (N_6563,N_6280,N_6252);
nor U6564 (N_6564,N_6288,N_6293);
xor U6565 (N_6565,N_6249,N_6228);
nand U6566 (N_6566,N_6246,N_6285);
or U6567 (N_6567,N_6325,N_6281);
or U6568 (N_6568,N_6236,N_6228);
nor U6569 (N_6569,N_6280,N_6291);
or U6570 (N_6570,N_6354,N_6211);
xnor U6571 (N_6571,N_6314,N_6347);
nor U6572 (N_6572,N_6298,N_6212);
nand U6573 (N_6573,N_6358,N_6307);
nand U6574 (N_6574,N_6344,N_6273);
xor U6575 (N_6575,N_6252,N_6327);
or U6576 (N_6576,N_6285,N_6328);
and U6577 (N_6577,N_6303,N_6288);
xor U6578 (N_6578,N_6340,N_6249);
and U6579 (N_6579,N_6372,N_6289);
or U6580 (N_6580,N_6236,N_6238);
xnor U6581 (N_6581,N_6239,N_6231);
or U6582 (N_6582,N_6243,N_6207);
or U6583 (N_6583,N_6242,N_6218);
nor U6584 (N_6584,N_6230,N_6382);
nor U6585 (N_6585,N_6213,N_6233);
or U6586 (N_6586,N_6321,N_6356);
or U6587 (N_6587,N_6376,N_6352);
xor U6588 (N_6588,N_6349,N_6317);
xnor U6589 (N_6589,N_6385,N_6387);
nand U6590 (N_6590,N_6278,N_6365);
xor U6591 (N_6591,N_6318,N_6327);
and U6592 (N_6592,N_6348,N_6278);
nor U6593 (N_6593,N_6386,N_6307);
xor U6594 (N_6594,N_6369,N_6300);
or U6595 (N_6595,N_6377,N_6308);
or U6596 (N_6596,N_6217,N_6380);
xnor U6597 (N_6597,N_6319,N_6397);
nand U6598 (N_6598,N_6231,N_6266);
xor U6599 (N_6599,N_6293,N_6249);
or U6600 (N_6600,N_6404,N_6422);
nor U6601 (N_6601,N_6455,N_6513);
xor U6602 (N_6602,N_6464,N_6421);
or U6603 (N_6603,N_6558,N_6461);
xor U6604 (N_6604,N_6599,N_6428);
or U6605 (N_6605,N_6526,N_6587);
or U6606 (N_6606,N_6485,N_6446);
and U6607 (N_6607,N_6423,N_6552);
or U6608 (N_6608,N_6566,N_6564);
or U6609 (N_6609,N_6524,N_6501);
nor U6610 (N_6610,N_6519,N_6570);
or U6611 (N_6611,N_6520,N_6580);
nor U6612 (N_6612,N_6578,N_6507);
xnor U6613 (N_6613,N_6518,N_6505);
xnor U6614 (N_6614,N_6545,N_6589);
or U6615 (N_6615,N_6453,N_6540);
xnor U6616 (N_6616,N_6563,N_6411);
and U6617 (N_6617,N_6441,N_6593);
and U6618 (N_6618,N_6476,N_6445);
or U6619 (N_6619,N_6527,N_6573);
xor U6620 (N_6620,N_6562,N_6546);
nor U6621 (N_6621,N_6510,N_6444);
nor U6622 (N_6622,N_6450,N_6429);
or U6623 (N_6623,N_6407,N_6438);
and U6624 (N_6624,N_6581,N_6584);
nand U6625 (N_6625,N_6521,N_6538);
xnor U6626 (N_6626,N_6537,N_6588);
nand U6627 (N_6627,N_6419,N_6596);
and U6628 (N_6628,N_6454,N_6557);
xor U6629 (N_6629,N_6437,N_6469);
and U6630 (N_6630,N_6582,N_6583);
nand U6631 (N_6631,N_6555,N_6416);
nand U6632 (N_6632,N_6418,N_6548);
and U6633 (N_6633,N_6488,N_6465);
or U6634 (N_6634,N_6515,N_6591);
xor U6635 (N_6635,N_6494,N_6479);
nor U6636 (N_6636,N_6535,N_6402);
nor U6637 (N_6637,N_6482,N_6542);
and U6638 (N_6638,N_6594,N_6511);
or U6639 (N_6639,N_6477,N_6449);
and U6640 (N_6640,N_6560,N_6539);
or U6641 (N_6641,N_6550,N_6514);
xnor U6642 (N_6642,N_6480,N_6487);
xor U6643 (N_6643,N_6575,N_6456);
nor U6644 (N_6644,N_6484,N_6447);
and U6645 (N_6645,N_6448,N_6413);
and U6646 (N_6646,N_6532,N_6400);
nor U6647 (N_6647,N_6457,N_6590);
or U6648 (N_6648,N_6597,N_6431);
or U6649 (N_6649,N_6585,N_6533);
nand U6650 (N_6650,N_6528,N_6424);
and U6651 (N_6651,N_6420,N_6565);
and U6652 (N_6652,N_6543,N_6414);
nor U6653 (N_6653,N_6579,N_6439);
nand U6654 (N_6654,N_6406,N_6486);
xnor U6655 (N_6655,N_6572,N_6576);
nor U6656 (N_6656,N_6569,N_6517);
nand U6657 (N_6657,N_6432,N_6561);
or U6658 (N_6658,N_6451,N_6408);
or U6659 (N_6659,N_6595,N_6525);
and U6660 (N_6660,N_6499,N_6458);
or U6661 (N_6661,N_6498,N_6551);
or U6662 (N_6662,N_6536,N_6491);
nor U6663 (N_6663,N_6412,N_6506);
and U6664 (N_6664,N_6567,N_6427);
and U6665 (N_6665,N_6497,N_6577);
nor U6666 (N_6666,N_6463,N_6553);
and U6667 (N_6667,N_6547,N_6592);
xnor U6668 (N_6668,N_6473,N_6534);
or U6669 (N_6669,N_6409,N_6509);
or U6670 (N_6670,N_6529,N_6544);
or U6671 (N_6671,N_6436,N_6568);
nor U6672 (N_6672,N_6433,N_6502);
nor U6673 (N_6673,N_6462,N_6493);
and U6674 (N_6674,N_6504,N_6522);
nand U6675 (N_6675,N_6405,N_6492);
nand U6676 (N_6676,N_6478,N_6495);
nand U6677 (N_6677,N_6426,N_6559);
nand U6678 (N_6678,N_6496,N_6417);
or U6679 (N_6679,N_6574,N_6470);
and U6680 (N_6680,N_6598,N_6467);
nor U6681 (N_6681,N_6500,N_6531);
nor U6682 (N_6682,N_6541,N_6466);
or U6683 (N_6683,N_6586,N_6523);
nor U6684 (N_6684,N_6483,N_6530);
and U6685 (N_6685,N_6512,N_6460);
xor U6686 (N_6686,N_6549,N_6442);
nor U6687 (N_6687,N_6440,N_6475);
or U6688 (N_6688,N_6452,N_6403);
or U6689 (N_6689,N_6489,N_6425);
or U6690 (N_6690,N_6508,N_6443);
or U6691 (N_6691,N_6481,N_6554);
nand U6692 (N_6692,N_6434,N_6503);
xnor U6693 (N_6693,N_6471,N_6430);
xnor U6694 (N_6694,N_6556,N_6468);
nor U6695 (N_6695,N_6401,N_6490);
and U6696 (N_6696,N_6415,N_6435);
nor U6697 (N_6697,N_6474,N_6571);
nor U6698 (N_6698,N_6516,N_6472);
nand U6699 (N_6699,N_6410,N_6459);
xor U6700 (N_6700,N_6578,N_6530);
and U6701 (N_6701,N_6488,N_6422);
nor U6702 (N_6702,N_6476,N_6541);
nand U6703 (N_6703,N_6468,N_6429);
xnor U6704 (N_6704,N_6567,N_6479);
xnor U6705 (N_6705,N_6433,N_6514);
nand U6706 (N_6706,N_6589,N_6500);
nand U6707 (N_6707,N_6565,N_6540);
or U6708 (N_6708,N_6446,N_6575);
xor U6709 (N_6709,N_6572,N_6497);
nand U6710 (N_6710,N_6491,N_6496);
and U6711 (N_6711,N_6581,N_6494);
nor U6712 (N_6712,N_6563,N_6526);
and U6713 (N_6713,N_6501,N_6529);
nor U6714 (N_6714,N_6478,N_6411);
and U6715 (N_6715,N_6516,N_6524);
or U6716 (N_6716,N_6404,N_6434);
or U6717 (N_6717,N_6434,N_6577);
or U6718 (N_6718,N_6530,N_6501);
or U6719 (N_6719,N_6547,N_6403);
nand U6720 (N_6720,N_6515,N_6578);
nor U6721 (N_6721,N_6567,N_6480);
nor U6722 (N_6722,N_6426,N_6415);
and U6723 (N_6723,N_6509,N_6444);
xnor U6724 (N_6724,N_6440,N_6466);
nor U6725 (N_6725,N_6505,N_6438);
or U6726 (N_6726,N_6473,N_6442);
and U6727 (N_6727,N_6502,N_6411);
nand U6728 (N_6728,N_6415,N_6424);
nand U6729 (N_6729,N_6502,N_6575);
nor U6730 (N_6730,N_6599,N_6455);
or U6731 (N_6731,N_6511,N_6451);
nor U6732 (N_6732,N_6480,N_6411);
and U6733 (N_6733,N_6404,N_6532);
xor U6734 (N_6734,N_6554,N_6589);
xnor U6735 (N_6735,N_6461,N_6503);
and U6736 (N_6736,N_6474,N_6461);
nand U6737 (N_6737,N_6543,N_6421);
and U6738 (N_6738,N_6545,N_6530);
or U6739 (N_6739,N_6421,N_6436);
xnor U6740 (N_6740,N_6504,N_6501);
xnor U6741 (N_6741,N_6436,N_6516);
nor U6742 (N_6742,N_6573,N_6555);
xnor U6743 (N_6743,N_6416,N_6544);
nand U6744 (N_6744,N_6494,N_6502);
and U6745 (N_6745,N_6433,N_6583);
nor U6746 (N_6746,N_6497,N_6592);
nor U6747 (N_6747,N_6538,N_6490);
nor U6748 (N_6748,N_6403,N_6542);
or U6749 (N_6749,N_6506,N_6527);
or U6750 (N_6750,N_6478,N_6497);
nand U6751 (N_6751,N_6503,N_6541);
xor U6752 (N_6752,N_6482,N_6486);
or U6753 (N_6753,N_6450,N_6575);
nand U6754 (N_6754,N_6417,N_6520);
xor U6755 (N_6755,N_6410,N_6463);
and U6756 (N_6756,N_6503,N_6425);
and U6757 (N_6757,N_6556,N_6492);
xor U6758 (N_6758,N_6470,N_6476);
nand U6759 (N_6759,N_6586,N_6560);
and U6760 (N_6760,N_6599,N_6574);
nor U6761 (N_6761,N_6533,N_6470);
xnor U6762 (N_6762,N_6532,N_6453);
nand U6763 (N_6763,N_6515,N_6498);
and U6764 (N_6764,N_6596,N_6496);
nor U6765 (N_6765,N_6505,N_6582);
nor U6766 (N_6766,N_6537,N_6517);
nand U6767 (N_6767,N_6468,N_6436);
or U6768 (N_6768,N_6572,N_6439);
nand U6769 (N_6769,N_6550,N_6499);
nor U6770 (N_6770,N_6411,N_6559);
nor U6771 (N_6771,N_6407,N_6531);
nor U6772 (N_6772,N_6517,N_6506);
and U6773 (N_6773,N_6495,N_6402);
and U6774 (N_6774,N_6569,N_6478);
nor U6775 (N_6775,N_6472,N_6524);
nor U6776 (N_6776,N_6501,N_6434);
nand U6777 (N_6777,N_6557,N_6555);
xnor U6778 (N_6778,N_6567,N_6413);
nor U6779 (N_6779,N_6529,N_6402);
and U6780 (N_6780,N_6578,N_6552);
nor U6781 (N_6781,N_6441,N_6479);
and U6782 (N_6782,N_6558,N_6416);
nor U6783 (N_6783,N_6442,N_6419);
and U6784 (N_6784,N_6538,N_6559);
nand U6785 (N_6785,N_6464,N_6578);
and U6786 (N_6786,N_6487,N_6516);
nor U6787 (N_6787,N_6426,N_6501);
or U6788 (N_6788,N_6439,N_6408);
nor U6789 (N_6789,N_6565,N_6474);
or U6790 (N_6790,N_6456,N_6570);
xor U6791 (N_6791,N_6444,N_6503);
or U6792 (N_6792,N_6536,N_6498);
xor U6793 (N_6793,N_6453,N_6580);
nor U6794 (N_6794,N_6492,N_6584);
or U6795 (N_6795,N_6435,N_6431);
xor U6796 (N_6796,N_6497,N_6540);
or U6797 (N_6797,N_6467,N_6474);
nand U6798 (N_6798,N_6445,N_6586);
and U6799 (N_6799,N_6447,N_6557);
and U6800 (N_6800,N_6736,N_6785);
nand U6801 (N_6801,N_6723,N_6759);
or U6802 (N_6802,N_6788,N_6644);
xnor U6803 (N_6803,N_6637,N_6728);
and U6804 (N_6804,N_6673,N_6621);
xnor U6805 (N_6805,N_6661,N_6604);
nor U6806 (N_6806,N_6707,N_6710);
xnor U6807 (N_6807,N_6787,N_6657);
nand U6808 (N_6808,N_6786,N_6625);
and U6809 (N_6809,N_6777,N_6682);
nand U6810 (N_6810,N_6658,N_6679);
xor U6811 (N_6811,N_6704,N_6750);
xnor U6812 (N_6812,N_6711,N_6762);
or U6813 (N_6813,N_6738,N_6702);
or U6814 (N_6814,N_6744,N_6634);
nand U6815 (N_6815,N_6698,N_6602);
nor U6816 (N_6816,N_6626,N_6789);
xnor U6817 (N_6817,N_6774,N_6678);
or U6818 (N_6818,N_6791,N_6615);
nand U6819 (N_6819,N_6645,N_6666);
xnor U6820 (N_6820,N_6616,N_6671);
nand U6821 (N_6821,N_6747,N_6717);
and U6822 (N_6822,N_6713,N_6798);
nand U6823 (N_6823,N_6724,N_6731);
nand U6824 (N_6824,N_6768,N_6726);
and U6825 (N_6825,N_6624,N_6674);
nand U6826 (N_6826,N_6638,N_6641);
nand U6827 (N_6827,N_6632,N_6633);
nand U6828 (N_6828,N_6772,N_6781);
xor U6829 (N_6829,N_6796,N_6683);
or U6830 (N_6830,N_6613,N_6716);
or U6831 (N_6831,N_6709,N_6623);
xnor U6832 (N_6832,N_6672,N_6687);
or U6833 (N_6833,N_6732,N_6600);
nand U6834 (N_6834,N_6648,N_6776);
nor U6835 (N_6835,N_6746,N_6756);
nand U6836 (N_6836,N_6601,N_6792);
or U6837 (N_6837,N_6618,N_6606);
nor U6838 (N_6838,N_6790,N_6783);
nor U6839 (N_6839,N_6700,N_6694);
nand U6840 (N_6840,N_6771,N_6640);
or U6841 (N_6841,N_6761,N_6733);
and U6842 (N_6842,N_6766,N_6688);
xor U6843 (N_6843,N_6603,N_6767);
and U6844 (N_6844,N_6764,N_6655);
nand U6845 (N_6845,N_6769,N_6742);
xnor U6846 (N_6846,N_6605,N_6718);
and U6847 (N_6847,N_6651,N_6743);
nand U6848 (N_6848,N_6730,N_6741);
xor U6849 (N_6849,N_6706,N_6660);
or U6850 (N_6850,N_6778,N_6721);
or U6851 (N_6851,N_6685,N_6753);
nor U6852 (N_6852,N_6740,N_6631);
nor U6853 (N_6853,N_6697,N_6754);
and U6854 (N_6854,N_6757,N_6681);
nor U6855 (N_6855,N_6650,N_6676);
and U6856 (N_6856,N_6663,N_6636);
and U6857 (N_6857,N_6779,N_6675);
or U6858 (N_6858,N_6691,N_6797);
nor U6859 (N_6859,N_6639,N_6654);
or U6860 (N_6860,N_6729,N_6611);
xnor U6861 (N_6861,N_6668,N_6782);
nor U6862 (N_6862,N_6799,N_6735);
or U6863 (N_6863,N_6622,N_6758);
nand U6864 (N_6864,N_6629,N_6749);
xnor U6865 (N_6865,N_6689,N_6794);
nor U6866 (N_6866,N_6748,N_6614);
or U6867 (N_6867,N_6627,N_6712);
nand U6868 (N_6868,N_6680,N_6699);
or U6869 (N_6869,N_6739,N_6703);
nand U6870 (N_6870,N_6701,N_6608);
and U6871 (N_6871,N_6630,N_6696);
xnor U6872 (N_6872,N_6734,N_6751);
and U6873 (N_6873,N_6773,N_6652);
nand U6874 (N_6874,N_6737,N_6607);
nand U6875 (N_6875,N_6642,N_6662);
xor U6876 (N_6876,N_6695,N_6690);
nand U6877 (N_6877,N_6635,N_6780);
nor U6878 (N_6878,N_6752,N_6727);
xor U6879 (N_6879,N_6745,N_6653);
xnor U6880 (N_6880,N_6692,N_6610);
or U6881 (N_6881,N_6719,N_6665);
or U6882 (N_6882,N_6659,N_6643);
xnor U6883 (N_6883,N_6609,N_6656);
or U6884 (N_6884,N_6722,N_6720);
nor U6885 (N_6885,N_6686,N_6670);
and U6886 (N_6886,N_6619,N_6684);
or U6887 (N_6887,N_6725,N_6693);
nand U6888 (N_6888,N_6628,N_6612);
nand U6889 (N_6889,N_6793,N_6763);
nor U6890 (N_6890,N_6617,N_6760);
or U6891 (N_6891,N_6677,N_6770);
nand U6892 (N_6892,N_6715,N_6667);
and U6893 (N_6893,N_6705,N_6775);
or U6894 (N_6894,N_6708,N_6755);
nor U6895 (N_6895,N_6669,N_6765);
or U6896 (N_6896,N_6649,N_6647);
xor U6897 (N_6897,N_6795,N_6664);
nor U6898 (N_6898,N_6646,N_6620);
nor U6899 (N_6899,N_6784,N_6714);
xor U6900 (N_6900,N_6610,N_6652);
nor U6901 (N_6901,N_6676,N_6679);
or U6902 (N_6902,N_6745,N_6622);
nand U6903 (N_6903,N_6774,N_6713);
xor U6904 (N_6904,N_6786,N_6692);
xor U6905 (N_6905,N_6664,N_6767);
and U6906 (N_6906,N_6774,N_6778);
xnor U6907 (N_6907,N_6767,N_6750);
or U6908 (N_6908,N_6627,N_6794);
and U6909 (N_6909,N_6656,N_6687);
nor U6910 (N_6910,N_6690,N_6793);
or U6911 (N_6911,N_6650,N_6671);
and U6912 (N_6912,N_6672,N_6623);
or U6913 (N_6913,N_6784,N_6742);
or U6914 (N_6914,N_6660,N_6778);
and U6915 (N_6915,N_6620,N_6653);
or U6916 (N_6916,N_6650,N_6605);
nand U6917 (N_6917,N_6720,N_6616);
nand U6918 (N_6918,N_6607,N_6634);
nand U6919 (N_6919,N_6691,N_6724);
xnor U6920 (N_6920,N_6689,N_6683);
nor U6921 (N_6921,N_6694,N_6716);
xor U6922 (N_6922,N_6773,N_6628);
nand U6923 (N_6923,N_6781,N_6718);
or U6924 (N_6924,N_6664,N_6641);
nand U6925 (N_6925,N_6676,N_6715);
and U6926 (N_6926,N_6702,N_6705);
or U6927 (N_6927,N_6716,N_6660);
xnor U6928 (N_6928,N_6747,N_6639);
nor U6929 (N_6929,N_6780,N_6624);
nand U6930 (N_6930,N_6722,N_6634);
xnor U6931 (N_6931,N_6725,N_6710);
and U6932 (N_6932,N_6673,N_6787);
xnor U6933 (N_6933,N_6647,N_6779);
nand U6934 (N_6934,N_6617,N_6651);
nand U6935 (N_6935,N_6720,N_6769);
nor U6936 (N_6936,N_6690,N_6722);
nand U6937 (N_6937,N_6794,N_6657);
or U6938 (N_6938,N_6618,N_6686);
and U6939 (N_6939,N_6796,N_6743);
nor U6940 (N_6940,N_6776,N_6678);
nor U6941 (N_6941,N_6674,N_6603);
or U6942 (N_6942,N_6717,N_6727);
nor U6943 (N_6943,N_6667,N_6642);
xor U6944 (N_6944,N_6733,N_6795);
or U6945 (N_6945,N_6759,N_6721);
or U6946 (N_6946,N_6774,N_6720);
and U6947 (N_6947,N_6749,N_6621);
nand U6948 (N_6948,N_6668,N_6772);
nor U6949 (N_6949,N_6770,N_6765);
xnor U6950 (N_6950,N_6658,N_6663);
and U6951 (N_6951,N_6708,N_6639);
nand U6952 (N_6952,N_6780,N_6798);
or U6953 (N_6953,N_6770,N_6685);
nor U6954 (N_6954,N_6610,N_6774);
and U6955 (N_6955,N_6778,N_6694);
nor U6956 (N_6956,N_6769,N_6680);
or U6957 (N_6957,N_6764,N_6688);
and U6958 (N_6958,N_6614,N_6644);
or U6959 (N_6959,N_6611,N_6761);
or U6960 (N_6960,N_6746,N_6634);
nor U6961 (N_6961,N_6734,N_6716);
xnor U6962 (N_6962,N_6724,N_6675);
nand U6963 (N_6963,N_6615,N_6770);
or U6964 (N_6964,N_6625,N_6733);
nor U6965 (N_6965,N_6721,N_6776);
xor U6966 (N_6966,N_6620,N_6675);
xor U6967 (N_6967,N_6620,N_6633);
and U6968 (N_6968,N_6771,N_6749);
nand U6969 (N_6969,N_6712,N_6777);
nand U6970 (N_6970,N_6747,N_6677);
and U6971 (N_6971,N_6773,N_6737);
nor U6972 (N_6972,N_6710,N_6709);
and U6973 (N_6973,N_6666,N_6670);
xor U6974 (N_6974,N_6609,N_6635);
or U6975 (N_6975,N_6615,N_6792);
nand U6976 (N_6976,N_6621,N_6743);
nor U6977 (N_6977,N_6752,N_6663);
and U6978 (N_6978,N_6673,N_6792);
or U6979 (N_6979,N_6796,N_6697);
and U6980 (N_6980,N_6603,N_6715);
and U6981 (N_6981,N_6704,N_6629);
or U6982 (N_6982,N_6606,N_6751);
or U6983 (N_6983,N_6624,N_6771);
nand U6984 (N_6984,N_6689,N_6751);
nand U6985 (N_6985,N_6737,N_6651);
nand U6986 (N_6986,N_6636,N_6778);
and U6987 (N_6987,N_6731,N_6696);
or U6988 (N_6988,N_6617,N_6678);
and U6989 (N_6989,N_6721,N_6670);
and U6990 (N_6990,N_6772,N_6673);
and U6991 (N_6991,N_6700,N_6780);
nand U6992 (N_6992,N_6692,N_6651);
nand U6993 (N_6993,N_6688,N_6713);
xnor U6994 (N_6994,N_6718,N_6608);
and U6995 (N_6995,N_6649,N_6729);
nand U6996 (N_6996,N_6609,N_6799);
xor U6997 (N_6997,N_6637,N_6618);
or U6998 (N_6998,N_6726,N_6760);
nor U6999 (N_6999,N_6770,N_6761);
nand U7000 (N_7000,N_6816,N_6917);
nor U7001 (N_7001,N_6983,N_6957);
nor U7002 (N_7002,N_6924,N_6901);
nor U7003 (N_7003,N_6960,N_6853);
and U7004 (N_7004,N_6992,N_6953);
xnor U7005 (N_7005,N_6881,N_6949);
nand U7006 (N_7006,N_6915,N_6877);
nor U7007 (N_7007,N_6996,N_6879);
or U7008 (N_7008,N_6878,N_6839);
nor U7009 (N_7009,N_6927,N_6951);
nand U7010 (N_7010,N_6805,N_6874);
and U7011 (N_7011,N_6926,N_6837);
and U7012 (N_7012,N_6928,N_6833);
nand U7013 (N_7013,N_6962,N_6929);
or U7014 (N_7014,N_6986,N_6967);
and U7015 (N_7015,N_6932,N_6891);
or U7016 (N_7016,N_6885,N_6834);
and U7017 (N_7017,N_6975,N_6889);
or U7018 (N_7018,N_6974,N_6899);
nor U7019 (N_7019,N_6843,N_6988);
nand U7020 (N_7020,N_6825,N_6981);
nor U7021 (N_7021,N_6813,N_6993);
nor U7022 (N_7022,N_6990,N_6835);
or U7023 (N_7023,N_6958,N_6872);
xor U7024 (N_7024,N_6982,N_6998);
nor U7025 (N_7025,N_6806,N_6888);
and U7026 (N_7026,N_6846,N_6875);
nor U7027 (N_7027,N_6954,N_6966);
xnor U7028 (N_7028,N_6883,N_6937);
or U7029 (N_7029,N_6934,N_6999);
or U7030 (N_7030,N_6922,N_6923);
nand U7031 (N_7031,N_6900,N_6817);
nand U7032 (N_7032,N_6855,N_6904);
xnor U7033 (N_7033,N_6867,N_6819);
xor U7034 (N_7034,N_6896,N_6925);
nand U7035 (N_7035,N_6845,N_6919);
and U7036 (N_7036,N_6947,N_6909);
nand U7037 (N_7037,N_6895,N_6822);
or U7038 (N_7038,N_6848,N_6858);
xnor U7039 (N_7039,N_6801,N_6898);
xor U7040 (N_7040,N_6841,N_6829);
nand U7041 (N_7041,N_6930,N_6871);
and U7042 (N_7042,N_6897,N_6980);
or U7043 (N_7043,N_6863,N_6994);
and U7044 (N_7044,N_6987,N_6820);
xnor U7045 (N_7045,N_6938,N_6976);
nand U7046 (N_7046,N_6936,N_6859);
and U7047 (N_7047,N_6800,N_6995);
or U7048 (N_7048,N_6977,N_6973);
and U7049 (N_7049,N_6946,N_6943);
or U7050 (N_7050,N_6824,N_6902);
nand U7051 (N_7051,N_6876,N_6997);
or U7052 (N_7052,N_6964,N_6942);
nand U7053 (N_7053,N_6840,N_6887);
xor U7054 (N_7054,N_6911,N_6920);
nand U7055 (N_7055,N_6865,N_6884);
nand U7056 (N_7056,N_6972,N_6940);
nand U7057 (N_7057,N_6826,N_6956);
nand U7058 (N_7058,N_6815,N_6886);
nor U7059 (N_7059,N_6894,N_6852);
or U7060 (N_7060,N_6844,N_6818);
or U7061 (N_7061,N_6868,N_6944);
nand U7062 (N_7062,N_6832,N_6941);
xnor U7063 (N_7063,N_6912,N_6913);
and U7064 (N_7064,N_6856,N_6882);
or U7065 (N_7065,N_6803,N_6918);
nand U7066 (N_7066,N_6810,N_6850);
xnor U7067 (N_7067,N_6893,N_6851);
nand U7068 (N_7068,N_6959,N_6984);
nand U7069 (N_7069,N_6823,N_6880);
or U7070 (N_7070,N_6860,N_6892);
or U7071 (N_7071,N_6989,N_6828);
and U7072 (N_7072,N_6866,N_6906);
nor U7073 (N_7073,N_6907,N_6939);
nor U7074 (N_7074,N_6804,N_6812);
or U7075 (N_7075,N_6808,N_6950);
nand U7076 (N_7076,N_6861,N_6945);
nor U7077 (N_7077,N_6979,N_6849);
nand U7078 (N_7078,N_6965,N_6821);
or U7079 (N_7079,N_6969,N_6802);
nand U7080 (N_7080,N_6914,N_6931);
nand U7081 (N_7081,N_6847,N_6910);
xor U7082 (N_7082,N_6814,N_6890);
and U7083 (N_7083,N_6862,N_6836);
and U7084 (N_7084,N_6827,N_6870);
or U7085 (N_7085,N_6916,N_6955);
nand U7086 (N_7086,N_6991,N_6831);
and U7087 (N_7087,N_6842,N_6807);
and U7088 (N_7088,N_6971,N_6978);
nand U7089 (N_7089,N_6921,N_6963);
nand U7090 (N_7090,N_6864,N_6811);
and U7091 (N_7091,N_6961,N_6869);
xnor U7092 (N_7092,N_6908,N_6948);
and U7093 (N_7093,N_6854,N_6903);
nand U7094 (N_7094,N_6933,N_6905);
and U7095 (N_7095,N_6838,N_6952);
or U7096 (N_7096,N_6830,N_6968);
or U7097 (N_7097,N_6809,N_6970);
or U7098 (N_7098,N_6935,N_6857);
nor U7099 (N_7099,N_6873,N_6985);
nor U7100 (N_7100,N_6937,N_6916);
nand U7101 (N_7101,N_6939,N_6910);
or U7102 (N_7102,N_6826,N_6970);
xor U7103 (N_7103,N_6975,N_6811);
nand U7104 (N_7104,N_6837,N_6924);
or U7105 (N_7105,N_6980,N_6810);
nand U7106 (N_7106,N_6845,N_6933);
or U7107 (N_7107,N_6912,N_6981);
and U7108 (N_7108,N_6989,N_6972);
and U7109 (N_7109,N_6865,N_6814);
or U7110 (N_7110,N_6870,N_6866);
nor U7111 (N_7111,N_6922,N_6828);
xor U7112 (N_7112,N_6824,N_6895);
xor U7113 (N_7113,N_6876,N_6848);
or U7114 (N_7114,N_6924,N_6964);
nand U7115 (N_7115,N_6853,N_6981);
or U7116 (N_7116,N_6860,N_6993);
nor U7117 (N_7117,N_6856,N_6877);
nand U7118 (N_7118,N_6994,N_6949);
nor U7119 (N_7119,N_6897,N_6866);
nor U7120 (N_7120,N_6982,N_6825);
and U7121 (N_7121,N_6903,N_6834);
nand U7122 (N_7122,N_6843,N_6835);
and U7123 (N_7123,N_6917,N_6873);
nand U7124 (N_7124,N_6815,N_6950);
or U7125 (N_7125,N_6926,N_6893);
and U7126 (N_7126,N_6845,N_6937);
and U7127 (N_7127,N_6881,N_6821);
or U7128 (N_7128,N_6870,N_6878);
nand U7129 (N_7129,N_6890,N_6801);
nor U7130 (N_7130,N_6838,N_6915);
or U7131 (N_7131,N_6836,N_6973);
and U7132 (N_7132,N_6966,N_6843);
nor U7133 (N_7133,N_6958,N_6818);
xor U7134 (N_7134,N_6815,N_6920);
xnor U7135 (N_7135,N_6810,N_6958);
nand U7136 (N_7136,N_6973,N_6868);
xnor U7137 (N_7137,N_6905,N_6918);
nand U7138 (N_7138,N_6850,N_6805);
xor U7139 (N_7139,N_6878,N_6837);
nor U7140 (N_7140,N_6855,N_6978);
xnor U7141 (N_7141,N_6992,N_6946);
nor U7142 (N_7142,N_6863,N_6981);
and U7143 (N_7143,N_6914,N_6980);
or U7144 (N_7144,N_6807,N_6912);
or U7145 (N_7145,N_6878,N_6825);
or U7146 (N_7146,N_6912,N_6971);
or U7147 (N_7147,N_6886,N_6999);
nand U7148 (N_7148,N_6826,N_6854);
nor U7149 (N_7149,N_6988,N_6900);
nand U7150 (N_7150,N_6891,N_6943);
xor U7151 (N_7151,N_6910,N_6804);
xor U7152 (N_7152,N_6904,N_6806);
nor U7153 (N_7153,N_6824,N_6868);
or U7154 (N_7154,N_6974,N_6822);
nor U7155 (N_7155,N_6952,N_6957);
nand U7156 (N_7156,N_6975,N_6852);
and U7157 (N_7157,N_6974,N_6939);
nand U7158 (N_7158,N_6896,N_6963);
or U7159 (N_7159,N_6893,N_6922);
nand U7160 (N_7160,N_6980,N_6902);
xor U7161 (N_7161,N_6955,N_6837);
and U7162 (N_7162,N_6998,N_6832);
nor U7163 (N_7163,N_6812,N_6911);
nand U7164 (N_7164,N_6899,N_6886);
or U7165 (N_7165,N_6990,N_6844);
or U7166 (N_7166,N_6893,N_6999);
or U7167 (N_7167,N_6992,N_6973);
or U7168 (N_7168,N_6847,N_6897);
or U7169 (N_7169,N_6833,N_6993);
and U7170 (N_7170,N_6817,N_6895);
nor U7171 (N_7171,N_6995,N_6943);
or U7172 (N_7172,N_6939,N_6854);
and U7173 (N_7173,N_6872,N_6856);
or U7174 (N_7174,N_6803,N_6970);
and U7175 (N_7175,N_6804,N_6871);
nand U7176 (N_7176,N_6802,N_6932);
or U7177 (N_7177,N_6928,N_6932);
or U7178 (N_7178,N_6887,N_6890);
nand U7179 (N_7179,N_6930,N_6881);
and U7180 (N_7180,N_6825,N_6999);
nor U7181 (N_7181,N_6878,N_6897);
or U7182 (N_7182,N_6995,N_6947);
nand U7183 (N_7183,N_6844,N_6921);
or U7184 (N_7184,N_6868,N_6981);
nand U7185 (N_7185,N_6924,N_6965);
or U7186 (N_7186,N_6815,N_6990);
or U7187 (N_7187,N_6843,N_6997);
nand U7188 (N_7188,N_6814,N_6887);
or U7189 (N_7189,N_6864,N_6826);
xnor U7190 (N_7190,N_6985,N_6955);
nor U7191 (N_7191,N_6805,N_6801);
nor U7192 (N_7192,N_6840,N_6940);
or U7193 (N_7193,N_6842,N_6891);
xor U7194 (N_7194,N_6903,N_6913);
or U7195 (N_7195,N_6919,N_6920);
or U7196 (N_7196,N_6983,N_6800);
nor U7197 (N_7197,N_6847,N_6830);
and U7198 (N_7198,N_6962,N_6815);
nor U7199 (N_7199,N_6953,N_6825);
nor U7200 (N_7200,N_7033,N_7094);
or U7201 (N_7201,N_7185,N_7087);
or U7202 (N_7202,N_7156,N_7066);
nor U7203 (N_7203,N_7139,N_7148);
and U7204 (N_7204,N_7021,N_7192);
and U7205 (N_7205,N_7197,N_7022);
or U7206 (N_7206,N_7183,N_7096);
and U7207 (N_7207,N_7101,N_7102);
nor U7208 (N_7208,N_7002,N_7157);
and U7209 (N_7209,N_7116,N_7098);
or U7210 (N_7210,N_7184,N_7137);
and U7211 (N_7211,N_7028,N_7029);
nand U7212 (N_7212,N_7046,N_7080);
nand U7213 (N_7213,N_7173,N_7127);
and U7214 (N_7214,N_7031,N_7054);
or U7215 (N_7215,N_7011,N_7120);
or U7216 (N_7216,N_7108,N_7032);
or U7217 (N_7217,N_7118,N_7194);
and U7218 (N_7218,N_7065,N_7167);
nand U7219 (N_7219,N_7111,N_7043);
nor U7220 (N_7220,N_7084,N_7082);
or U7221 (N_7221,N_7069,N_7129);
nor U7222 (N_7222,N_7126,N_7189);
nand U7223 (N_7223,N_7160,N_7188);
or U7224 (N_7224,N_7196,N_7091);
xnor U7225 (N_7225,N_7198,N_7124);
xor U7226 (N_7226,N_7180,N_7056);
nand U7227 (N_7227,N_7105,N_7007);
and U7228 (N_7228,N_7039,N_7141);
nand U7229 (N_7229,N_7068,N_7143);
nand U7230 (N_7230,N_7186,N_7109);
and U7231 (N_7231,N_7115,N_7131);
nand U7232 (N_7232,N_7057,N_7051);
xnor U7233 (N_7233,N_7153,N_7005);
nor U7234 (N_7234,N_7162,N_7117);
nand U7235 (N_7235,N_7138,N_7099);
or U7236 (N_7236,N_7178,N_7163);
xnor U7237 (N_7237,N_7086,N_7103);
xor U7238 (N_7238,N_7042,N_7061);
or U7239 (N_7239,N_7121,N_7154);
and U7240 (N_7240,N_7179,N_7037);
nand U7241 (N_7241,N_7158,N_7170);
and U7242 (N_7242,N_7172,N_7190);
nand U7243 (N_7243,N_7125,N_7164);
nor U7244 (N_7244,N_7052,N_7159);
nand U7245 (N_7245,N_7135,N_7067);
and U7246 (N_7246,N_7079,N_7191);
nand U7247 (N_7247,N_7095,N_7083);
nand U7248 (N_7248,N_7088,N_7044);
xor U7249 (N_7249,N_7050,N_7155);
nor U7250 (N_7250,N_7058,N_7055);
nor U7251 (N_7251,N_7015,N_7014);
and U7252 (N_7252,N_7006,N_7047);
or U7253 (N_7253,N_7074,N_7049);
nor U7254 (N_7254,N_7176,N_7133);
and U7255 (N_7255,N_7025,N_7149);
xnor U7256 (N_7256,N_7174,N_7182);
or U7257 (N_7257,N_7045,N_7070);
nor U7258 (N_7258,N_7062,N_7072);
or U7259 (N_7259,N_7195,N_7144);
or U7260 (N_7260,N_7181,N_7114);
xor U7261 (N_7261,N_7018,N_7128);
nor U7262 (N_7262,N_7009,N_7017);
nor U7263 (N_7263,N_7026,N_7175);
or U7264 (N_7264,N_7100,N_7150);
or U7265 (N_7265,N_7147,N_7110);
and U7266 (N_7266,N_7177,N_7187);
nor U7267 (N_7267,N_7053,N_7071);
nand U7268 (N_7268,N_7085,N_7059);
nand U7269 (N_7269,N_7089,N_7146);
or U7270 (N_7270,N_7168,N_7023);
xor U7271 (N_7271,N_7092,N_7004);
or U7272 (N_7272,N_7010,N_7123);
and U7273 (N_7273,N_7076,N_7152);
nand U7274 (N_7274,N_7064,N_7130);
xnor U7275 (N_7275,N_7078,N_7016);
nor U7276 (N_7276,N_7104,N_7112);
nand U7277 (N_7277,N_7134,N_7073);
or U7278 (N_7278,N_7161,N_7119);
or U7279 (N_7279,N_7034,N_7060);
nor U7280 (N_7280,N_7193,N_7035);
xor U7281 (N_7281,N_7113,N_7019);
nand U7282 (N_7282,N_7003,N_7166);
and U7283 (N_7283,N_7036,N_7077);
nor U7284 (N_7284,N_7107,N_7013);
and U7285 (N_7285,N_7106,N_7171);
and U7286 (N_7286,N_7008,N_7012);
or U7287 (N_7287,N_7075,N_7024);
nand U7288 (N_7288,N_7020,N_7040);
xor U7289 (N_7289,N_7169,N_7145);
and U7290 (N_7290,N_7199,N_7048);
xor U7291 (N_7291,N_7136,N_7000);
nor U7292 (N_7292,N_7041,N_7038);
or U7293 (N_7293,N_7001,N_7122);
nand U7294 (N_7294,N_7142,N_7165);
or U7295 (N_7295,N_7063,N_7030);
and U7296 (N_7296,N_7132,N_7027);
xnor U7297 (N_7297,N_7097,N_7140);
and U7298 (N_7298,N_7151,N_7081);
or U7299 (N_7299,N_7090,N_7093);
nor U7300 (N_7300,N_7116,N_7087);
xor U7301 (N_7301,N_7091,N_7125);
or U7302 (N_7302,N_7069,N_7117);
nand U7303 (N_7303,N_7077,N_7105);
nor U7304 (N_7304,N_7073,N_7043);
or U7305 (N_7305,N_7040,N_7039);
or U7306 (N_7306,N_7074,N_7183);
or U7307 (N_7307,N_7184,N_7069);
nor U7308 (N_7308,N_7089,N_7117);
or U7309 (N_7309,N_7088,N_7139);
nor U7310 (N_7310,N_7133,N_7171);
and U7311 (N_7311,N_7070,N_7178);
xnor U7312 (N_7312,N_7074,N_7195);
and U7313 (N_7313,N_7104,N_7053);
nor U7314 (N_7314,N_7132,N_7060);
nor U7315 (N_7315,N_7178,N_7005);
xor U7316 (N_7316,N_7142,N_7077);
or U7317 (N_7317,N_7105,N_7139);
nor U7318 (N_7318,N_7048,N_7099);
or U7319 (N_7319,N_7090,N_7086);
or U7320 (N_7320,N_7068,N_7073);
or U7321 (N_7321,N_7009,N_7092);
nand U7322 (N_7322,N_7010,N_7165);
xnor U7323 (N_7323,N_7101,N_7187);
nand U7324 (N_7324,N_7070,N_7094);
or U7325 (N_7325,N_7023,N_7066);
nand U7326 (N_7326,N_7016,N_7008);
xnor U7327 (N_7327,N_7088,N_7127);
nand U7328 (N_7328,N_7121,N_7148);
and U7329 (N_7329,N_7195,N_7100);
or U7330 (N_7330,N_7129,N_7163);
or U7331 (N_7331,N_7088,N_7199);
nand U7332 (N_7332,N_7153,N_7108);
nor U7333 (N_7333,N_7042,N_7070);
or U7334 (N_7334,N_7122,N_7176);
and U7335 (N_7335,N_7028,N_7121);
and U7336 (N_7336,N_7146,N_7027);
xnor U7337 (N_7337,N_7097,N_7083);
nor U7338 (N_7338,N_7165,N_7107);
xnor U7339 (N_7339,N_7068,N_7167);
nand U7340 (N_7340,N_7183,N_7124);
and U7341 (N_7341,N_7096,N_7141);
nand U7342 (N_7342,N_7059,N_7198);
or U7343 (N_7343,N_7187,N_7111);
xnor U7344 (N_7344,N_7154,N_7116);
xnor U7345 (N_7345,N_7050,N_7019);
xor U7346 (N_7346,N_7033,N_7129);
or U7347 (N_7347,N_7155,N_7031);
nand U7348 (N_7348,N_7087,N_7004);
and U7349 (N_7349,N_7043,N_7086);
and U7350 (N_7350,N_7154,N_7125);
nor U7351 (N_7351,N_7065,N_7057);
nand U7352 (N_7352,N_7154,N_7012);
and U7353 (N_7353,N_7146,N_7189);
xnor U7354 (N_7354,N_7045,N_7171);
or U7355 (N_7355,N_7139,N_7040);
nand U7356 (N_7356,N_7113,N_7198);
nor U7357 (N_7357,N_7023,N_7074);
nand U7358 (N_7358,N_7105,N_7078);
nand U7359 (N_7359,N_7086,N_7074);
or U7360 (N_7360,N_7116,N_7009);
or U7361 (N_7361,N_7159,N_7033);
xor U7362 (N_7362,N_7036,N_7057);
xnor U7363 (N_7363,N_7058,N_7197);
xor U7364 (N_7364,N_7078,N_7082);
xnor U7365 (N_7365,N_7017,N_7031);
xor U7366 (N_7366,N_7063,N_7041);
and U7367 (N_7367,N_7132,N_7176);
and U7368 (N_7368,N_7084,N_7064);
and U7369 (N_7369,N_7158,N_7133);
or U7370 (N_7370,N_7043,N_7137);
nor U7371 (N_7371,N_7018,N_7044);
or U7372 (N_7372,N_7121,N_7024);
nor U7373 (N_7373,N_7099,N_7093);
xnor U7374 (N_7374,N_7163,N_7066);
nand U7375 (N_7375,N_7181,N_7154);
xnor U7376 (N_7376,N_7194,N_7152);
nand U7377 (N_7377,N_7091,N_7105);
xnor U7378 (N_7378,N_7065,N_7075);
nor U7379 (N_7379,N_7182,N_7067);
nand U7380 (N_7380,N_7096,N_7090);
nand U7381 (N_7381,N_7116,N_7044);
nor U7382 (N_7382,N_7149,N_7054);
nand U7383 (N_7383,N_7091,N_7088);
and U7384 (N_7384,N_7147,N_7131);
xnor U7385 (N_7385,N_7145,N_7005);
or U7386 (N_7386,N_7112,N_7014);
nor U7387 (N_7387,N_7147,N_7093);
xnor U7388 (N_7388,N_7189,N_7041);
nand U7389 (N_7389,N_7197,N_7142);
nand U7390 (N_7390,N_7014,N_7154);
nand U7391 (N_7391,N_7060,N_7094);
nor U7392 (N_7392,N_7191,N_7050);
or U7393 (N_7393,N_7117,N_7191);
or U7394 (N_7394,N_7104,N_7077);
xor U7395 (N_7395,N_7022,N_7071);
and U7396 (N_7396,N_7127,N_7133);
xor U7397 (N_7397,N_7104,N_7010);
xor U7398 (N_7398,N_7040,N_7094);
xor U7399 (N_7399,N_7129,N_7138);
or U7400 (N_7400,N_7279,N_7308);
xnor U7401 (N_7401,N_7390,N_7310);
xnor U7402 (N_7402,N_7242,N_7385);
or U7403 (N_7403,N_7399,N_7296);
xor U7404 (N_7404,N_7374,N_7284);
or U7405 (N_7405,N_7249,N_7245);
nand U7406 (N_7406,N_7337,N_7392);
and U7407 (N_7407,N_7240,N_7262);
or U7408 (N_7408,N_7386,N_7257);
or U7409 (N_7409,N_7204,N_7342);
or U7410 (N_7410,N_7312,N_7301);
xnor U7411 (N_7411,N_7377,N_7320);
xnor U7412 (N_7412,N_7307,N_7291);
xor U7413 (N_7413,N_7295,N_7311);
or U7414 (N_7414,N_7230,N_7233);
and U7415 (N_7415,N_7238,N_7353);
xnor U7416 (N_7416,N_7354,N_7394);
nand U7417 (N_7417,N_7289,N_7209);
or U7418 (N_7418,N_7317,N_7272);
xor U7419 (N_7419,N_7280,N_7202);
xor U7420 (N_7420,N_7373,N_7397);
nand U7421 (N_7421,N_7314,N_7247);
or U7422 (N_7422,N_7277,N_7269);
nand U7423 (N_7423,N_7232,N_7243);
nor U7424 (N_7424,N_7225,N_7341);
nand U7425 (N_7425,N_7275,N_7328);
nand U7426 (N_7426,N_7207,N_7323);
and U7427 (N_7427,N_7234,N_7261);
nand U7428 (N_7428,N_7203,N_7200);
nor U7429 (N_7429,N_7357,N_7201);
or U7430 (N_7430,N_7366,N_7348);
xor U7431 (N_7431,N_7218,N_7299);
xnor U7432 (N_7432,N_7274,N_7302);
or U7433 (N_7433,N_7263,N_7321);
and U7434 (N_7434,N_7344,N_7375);
xnor U7435 (N_7435,N_7379,N_7268);
or U7436 (N_7436,N_7389,N_7343);
and U7437 (N_7437,N_7316,N_7333);
or U7438 (N_7438,N_7215,N_7309);
xnor U7439 (N_7439,N_7259,N_7294);
and U7440 (N_7440,N_7362,N_7332);
and U7441 (N_7441,N_7290,N_7278);
nand U7442 (N_7442,N_7255,N_7372);
nand U7443 (N_7443,N_7398,N_7300);
or U7444 (N_7444,N_7219,N_7382);
nand U7445 (N_7445,N_7387,N_7250);
and U7446 (N_7446,N_7254,N_7251);
or U7447 (N_7447,N_7271,N_7347);
or U7448 (N_7448,N_7383,N_7351);
or U7449 (N_7449,N_7287,N_7248);
nor U7450 (N_7450,N_7208,N_7298);
or U7451 (N_7451,N_7244,N_7346);
or U7452 (N_7452,N_7358,N_7330);
nand U7453 (N_7453,N_7396,N_7359);
and U7454 (N_7454,N_7303,N_7267);
nand U7455 (N_7455,N_7340,N_7239);
nand U7456 (N_7456,N_7292,N_7227);
and U7457 (N_7457,N_7378,N_7221);
and U7458 (N_7458,N_7253,N_7288);
or U7459 (N_7459,N_7276,N_7217);
xnor U7460 (N_7460,N_7325,N_7206);
nor U7461 (N_7461,N_7270,N_7356);
nand U7462 (N_7462,N_7322,N_7313);
xor U7463 (N_7463,N_7350,N_7380);
xnor U7464 (N_7464,N_7335,N_7282);
nor U7465 (N_7465,N_7327,N_7336);
nand U7466 (N_7466,N_7384,N_7319);
or U7467 (N_7467,N_7226,N_7283);
nand U7468 (N_7468,N_7318,N_7381);
or U7469 (N_7469,N_7220,N_7329);
or U7470 (N_7470,N_7315,N_7236);
or U7471 (N_7471,N_7212,N_7246);
and U7472 (N_7472,N_7228,N_7368);
or U7473 (N_7473,N_7252,N_7391);
or U7474 (N_7474,N_7393,N_7214);
and U7475 (N_7475,N_7334,N_7369);
and U7476 (N_7476,N_7370,N_7224);
and U7477 (N_7477,N_7205,N_7326);
and U7478 (N_7478,N_7361,N_7216);
or U7479 (N_7479,N_7258,N_7297);
xnor U7480 (N_7480,N_7305,N_7324);
nor U7481 (N_7481,N_7211,N_7213);
xnor U7482 (N_7482,N_7293,N_7363);
xor U7483 (N_7483,N_7229,N_7352);
nor U7484 (N_7484,N_7376,N_7281);
and U7485 (N_7485,N_7395,N_7285);
or U7486 (N_7486,N_7339,N_7364);
nor U7487 (N_7487,N_7265,N_7286);
nand U7488 (N_7488,N_7241,N_7360);
or U7489 (N_7489,N_7349,N_7365);
or U7490 (N_7490,N_7388,N_7367);
xor U7491 (N_7491,N_7266,N_7210);
and U7492 (N_7492,N_7264,N_7345);
nor U7493 (N_7493,N_7231,N_7273);
xnor U7494 (N_7494,N_7223,N_7222);
xnor U7495 (N_7495,N_7331,N_7371);
nand U7496 (N_7496,N_7355,N_7235);
nor U7497 (N_7497,N_7256,N_7338);
or U7498 (N_7498,N_7304,N_7237);
nand U7499 (N_7499,N_7260,N_7306);
or U7500 (N_7500,N_7343,N_7333);
nor U7501 (N_7501,N_7381,N_7316);
nor U7502 (N_7502,N_7356,N_7223);
and U7503 (N_7503,N_7226,N_7246);
nor U7504 (N_7504,N_7354,N_7317);
xor U7505 (N_7505,N_7326,N_7252);
or U7506 (N_7506,N_7363,N_7328);
or U7507 (N_7507,N_7344,N_7231);
nor U7508 (N_7508,N_7312,N_7254);
and U7509 (N_7509,N_7233,N_7277);
nand U7510 (N_7510,N_7207,N_7344);
nand U7511 (N_7511,N_7243,N_7366);
or U7512 (N_7512,N_7362,N_7394);
nor U7513 (N_7513,N_7390,N_7253);
xor U7514 (N_7514,N_7248,N_7206);
nand U7515 (N_7515,N_7346,N_7373);
and U7516 (N_7516,N_7274,N_7203);
xor U7517 (N_7517,N_7292,N_7382);
and U7518 (N_7518,N_7336,N_7221);
xor U7519 (N_7519,N_7265,N_7255);
nand U7520 (N_7520,N_7391,N_7247);
nand U7521 (N_7521,N_7256,N_7231);
nand U7522 (N_7522,N_7240,N_7349);
nor U7523 (N_7523,N_7281,N_7280);
xor U7524 (N_7524,N_7253,N_7297);
or U7525 (N_7525,N_7378,N_7286);
and U7526 (N_7526,N_7318,N_7287);
or U7527 (N_7527,N_7288,N_7348);
nand U7528 (N_7528,N_7341,N_7393);
nor U7529 (N_7529,N_7357,N_7390);
and U7530 (N_7530,N_7283,N_7218);
or U7531 (N_7531,N_7271,N_7213);
xor U7532 (N_7532,N_7260,N_7249);
xor U7533 (N_7533,N_7360,N_7218);
xnor U7534 (N_7534,N_7259,N_7322);
xnor U7535 (N_7535,N_7316,N_7265);
or U7536 (N_7536,N_7348,N_7305);
xor U7537 (N_7537,N_7230,N_7380);
xnor U7538 (N_7538,N_7242,N_7313);
nor U7539 (N_7539,N_7200,N_7267);
or U7540 (N_7540,N_7340,N_7367);
and U7541 (N_7541,N_7285,N_7265);
xnor U7542 (N_7542,N_7399,N_7235);
or U7543 (N_7543,N_7256,N_7354);
nor U7544 (N_7544,N_7356,N_7207);
xor U7545 (N_7545,N_7344,N_7268);
nand U7546 (N_7546,N_7369,N_7204);
nor U7547 (N_7547,N_7349,N_7201);
or U7548 (N_7548,N_7319,N_7313);
xor U7549 (N_7549,N_7393,N_7244);
or U7550 (N_7550,N_7200,N_7286);
xnor U7551 (N_7551,N_7283,N_7246);
nor U7552 (N_7552,N_7373,N_7214);
nor U7553 (N_7553,N_7357,N_7252);
xnor U7554 (N_7554,N_7357,N_7222);
and U7555 (N_7555,N_7262,N_7349);
nor U7556 (N_7556,N_7374,N_7354);
or U7557 (N_7557,N_7240,N_7201);
or U7558 (N_7558,N_7202,N_7206);
nand U7559 (N_7559,N_7358,N_7242);
xor U7560 (N_7560,N_7297,N_7359);
nand U7561 (N_7561,N_7272,N_7243);
nor U7562 (N_7562,N_7284,N_7370);
xnor U7563 (N_7563,N_7304,N_7289);
nor U7564 (N_7564,N_7299,N_7366);
and U7565 (N_7565,N_7223,N_7284);
nor U7566 (N_7566,N_7354,N_7388);
or U7567 (N_7567,N_7286,N_7356);
or U7568 (N_7568,N_7274,N_7282);
and U7569 (N_7569,N_7381,N_7285);
nand U7570 (N_7570,N_7395,N_7255);
or U7571 (N_7571,N_7346,N_7216);
nand U7572 (N_7572,N_7287,N_7208);
or U7573 (N_7573,N_7258,N_7200);
nand U7574 (N_7574,N_7202,N_7288);
or U7575 (N_7575,N_7232,N_7389);
nor U7576 (N_7576,N_7236,N_7277);
and U7577 (N_7577,N_7341,N_7336);
or U7578 (N_7578,N_7217,N_7201);
or U7579 (N_7579,N_7293,N_7367);
nor U7580 (N_7580,N_7247,N_7377);
or U7581 (N_7581,N_7324,N_7393);
or U7582 (N_7582,N_7332,N_7310);
xor U7583 (N_7583,N_7396,N_7341);
and U7584 (N_7584,N_7348,N_7397);
and U7585 (N_7585,N_7252,N_7313);
and U7586 (N_7586,N_7319,N_7245);
nor U7587 (N_7587,N_7251,N_7304);
nand U7588 (N_7588,N_7281,N_7303);
nand U7589 (N_7589,N_7233,N_7315);
and U7590 (N_7590,N_7205,N_7321);
nand U7591 (N_7591,N_7324,N_7208);
and U7592 (N_7592,N_7363,N_7289);
or U7593 (N_7593,N_7381,N_7249);
and U7594 (N_7594,N_7235,N_7284);
nand U7595 (N_7595,N_7387,N_7348);
nand U7596 (N_7596,N_7392,N_7213);
and U7597 (N_7597,N_7238,N_7276);
nor U7598 (N_7598,N_7280,N_7338);
or U7599 (N_7599,N_7294,N_7370);
nor U7600 (N_7600,N_7483,N_7587);
nand U7601 (N_7601,N_7570,N_7463);
and U7602 (N_7602,N_7573,N_7533);
and U7603 (N_7603,N_7491,N_7415);
and U7604 (N_7604,N_7543,N_7448);
or U7605 (N_7605,N_7468,N_7422);
nor U7606 (N_7606,N_7552,N_7523);
xnor U7607 (N_7607,N_7429,N_7576);
xor U7608 (N_7608,N_7556,N_7599);
or U7609 (N_7609,N_7484,N_7541);
nor U7610 (N_7610,N_7458,N_7549);
or U7611 (N_7611,N_7545,N_7544);
nand U7612 (N_7612,N_7527,N_7574);
or U7613 (N_7613,N_7504,N_7526);
or U7614 (N_7614,N_7461,N_7447);
xnor U7615 (N_7615,N_7404,N_7407);
or U7616 (N_7616,N_7542,N_7409);
nor U7617 (N_7617,N_7569,N_7412);
nor U7618 (N_7618,N_7450,N_7590);
nand U7619 (N_7619,N_7437,N_7440);
or U7620 (N_7620,N_7413,N_7402);
nand U7621 (N_7621,N_7558,N_7473);
nand U7622 (N_7622,N_7488,N_7567);
nand U7623 (N_7623,N_7411,N_7431);
nor U7624 (N_7624,N_7403,N_7535);
nand U7625 (N_7625,N_7454,N_7534);
nor U7626 (N_7626,N_7501,N_7439);
and U7627 (N_7627,N_7459,N_7503);
nor U7628 (N_7628,N_7594,N_7519);
xor U7629 (N_7629,N_7455,N_7562);
nor U7630 (N_7630,N_7490,N_7506);
xnor U7631 (N_7631,N_7497,N_7586);
nor U7632 (N_7632,N_7593,N_7554);
nand U7633 (N_7633,N_7456,N_7419);
nor U7634 (N_7634,N_7494,N_7584);
nand U7635 (N_7635,N_7598,N_7478);
or U7636 (N_7636,N_7482,N_7470);
or U7637 (N_7637,N_7565,N_7537);
xnor U7638 (N_7638,N_7445,N_7525);
nor U7639 (N_7639,N_7550,N_7515);
xnor U7640 (N_7640,N_7547,N_7592);
xor U7641 (N_7641,N_7514,N_7414);
nand U7642 (N_7642,N_7513,N_7528);
xnor U7643 (N_7643,N_7424,N_7571);
and U7644 (N_7644,N_7585,N_7559);
and U7645 (N_7645,N_7453,N_7441);
nor U7646 (N_7646,N_7405,N_7566);
nand U7647 (N_7647,N_7423,N_7564);
nor U7648 (N_7648,N_7492,N_7493);
nor U7649 (N_7649,N_7435,N_7444);
nor U7650 (N_7650,N_7553,N_7582);
and U7651 (N_7651,N_7575,N_7511);
nand U7652 (N_7652,N_7560,N_7507);
and U7653 (N_7653,N_7529,N_7426);
xor U7654 (N_7654,N_7597,N_7466);
nor U7655 (N_7655,N_7521,N_7464);
xor U7656 (N_7656,N_7406,N_7589);
or U7657 (N_7657,N_7578,N_7555);
nand U7658 (N_7658,N_7474,N_7475);
nand U7659 (N_7659,N_7516,N_7417);
and U7660 (N_7660,N_7479,N_7410);
or U7661 (N_7661,N_7530,N_7577);
nand U7662 (N_7662,N_7512,N_7522);
xnor U7663 (N_7663,N_7496,N_7532);
xor U7664 (N_7664,N_7443,N_7487);
and U7665 (N_7665,N_7536,N_7548);
nand U7666 (N_7666,N_7495,N_7452);
nand U7667 (N_7667,N_7517,N_7580);
and U7668 (N_7668,N_7457,N_7421);
nor U7669 (N_7669,N_7539,N_7510);
or U7670 (N_7670,N_7499,N_7416);
nand U7671 (N_7671,N_7408,N_7505);
xnor U7672 (N_7672,N_7442,N_7425);
or U7673 (N_7673,N_7438,N_7486);
nor U7674 (N_7674,N_7485,N_7401);
xnor U7675 (N_7675,N_7418,N_7476);
and U7676 (N_7676,N_7420,N_7508);
xnor U7677 (N_7677,N_7436,N_7561);
and U7678 (N_7678,N_7465,N_7462);
xor U7679 (N_7679,N_7531,N_7581);
xor U7680 (N_7680,N_7563,N_7432);
xnor U7681 (N_7681,N_7467,N_7524);
and U7682 (N_7682,N_7460,N_7557);
or U7683 (N_7683,N_7579,N_7400);
xor U7684 (N_7684,N_7433,N_7568);
nor U7685 (N_7685,N_7449,N_7588);
and U7686 (N_7686,N_7500,N_7518);
and U7687 (N_7687,N_7596,N_7430);
and U7688 (N_7688,N_7469,N_7471);
and U7689 (N_7689,N_7427,N_7509);
nand U7690 (N_7690,N_7446,N_7595);
and U7691 (N_7691,N_7502,N_7546);
xor U7692 (N_7692,N_7591,N_7538);
or U7693 (N_7693,N_7498,N_7489);
nand U7694 (N_7694,N_7540,N_7428);
nand U7695 (N_7695,N_7472,N_7583);
and U7696 (N_7696,N_7477,N_7520);
nor U7697 (N_7697,N_7481,N_7572);
nor U7698 (N_7698,N_7451,N_7551);
nand U7699 (N_7699,N_7434,N_7480);
nand U7700 (N_7700,N_7457,N_7598);
and U7701 (N_7701,N_7464,N_7442);
xor U7702 (N_7702,N_7463,N_7421);
or U7703 (N_7703,N_7573,N_7467);
nand U7704 (N_7704,N_7535,N_7467);
nor U7705 (N_7705,N_7522,N_7446);
and U7706 (N_7706,N_7547,N_7409);
nand U7707 (N_7707,N_7522,N_7572);
xnor U7708 (N_7708,N_7494,N_7577);
xor U7709 (N_7709,N_7492,N_7535);
and U7710 (N_7710,N_7583,N_7494);
nor U7711 (N_7711,N_7509,N_7481);
and U7712 (N_7712,N_7554,N_7535);
nor U7713 (N_7713,N_7535,N_7446);
xnor U7714 (N_7714,N_7439,N_7442);
nand U7715 (N_7715,N_7587,N_7562);
nor U7716 (N_7716,N_7459,N_7435);
xor U7717 (N_7717,N_7433,N_7522);
xnor U7718 (N_7718,N_7499,N_7443);
nand U7719 (N_7719,N_7445,N_7503);
and U7720 (N_7720,N_7494,N_7533);
or U7721 (N_7721,N_7501,N_7438);
and U7722 (N_7722,N_7454,N_7406);
nand U7723 (N_7723,N_7408,N_7429);
nand U7724 (N_7724,N_7432,N_7541);
or U7725 (N_7725,N_7545,N_7578);
nor U7726 (N_7726,N_7408,N_7580);
xor U7727 (N_7727,N_7400,N_7593);
nand U7728 (N_7728,N_7509,N_7573);
or U7729 (N_7729,N_7456,N_7500);
nor U7730 (N_7730,N_7418,N_7511);
nor U7731 (N_7731,N_7543,N_7557);
nor U7732 (N_7732,N_7591,N_7598);
xnor U7733 (N_7733,N_7413,N_7508);
xnor U7734 (N_7734,N_7411,N_7447);
or U7735 (N_7735,N_7519,N_7542);
and U7736 (N_7736,N_7593,N_7415);
or U7737 (N_7737,N_7462,N_7466);
or U7738 (N_7738,N_7447,N_7557);
or U7739 (N_7739,N_7537,N_7597);
nand U7740 (N_7740,N_7433,N_7593);
xnor U7741 (N_7741,N_7545,N_7527);
nor U7742 (N_7742,N_7464,N_7404);
nor U7743 (N_7743,N_7481,N_7409);
or U7744 (N_7744,N_7595,N_7444);
or U7745 (N_7745,N_7565,N_7517);
nand U7746 (N_7746,N_7575,N_7505);
or U7747 (N_7747,N_7548,N_7414);
xnor U7748 (N_7748,N_7515,N_7456);
nand U7749 (N_7749,N_7420,N_7576);
and U7750 (N_7750,N_7584,N_7526);
and U7751 (N_7751,N_7416,N_7570);
nand U7752 (N_7752,N_7554,N_7594);
or U7753 (N_7753,N_7599,N_7508);
nor U7754 (N_7754,N_7539,N_7562);
xnor U7755 (N_7755,N_7441,N_7494);
nand U7756 (N_7756,N_7594,N_7410);
and U7757 (N_7757,N_7443,N_7543);
xnor U7758 (N_7758,N_7536,N_7491);
xnor U7759 (N_7759,N_7555,N_7530);
and U7760 (N_7760,N_7465,N_7415);
nand U7761 (N_7761,N_7454,N_7419);
and U7762 (N_7762,N_7531,N_7572);
nor U7763 (N_7763,N_7522,N_7415);
nor U7764 (N_7764,N_7469,N_7449);
xnor U7765 (N_7765,N_7431,N_7522);
or U7766 (N_7766,N_7401,N_7457);
or U7767 (N_7767,N_7450,N_7406);
nand U7768 (N_7768,N_7469,N_7576);
or U7769 (N_7769,N_7439,N_7429);
nand U7770 (N_7770,N_7475,N_7445);
nor U7771 (N_7771,N_7484,N_7455);
or U7772 (N_7772,N_7593,N_7561);
nand U7773 (N_7773,N_7561,N_7478);
nor U7774 (N_7774,N_7479,N_7518);
nand U7775 (N_7775,N_7567,N_7458);
xor U7776 (N_7776,N_7592,N_7415);
xor U7777 (N_7777,N_7484,N_7578);
nand U7778 (N_7778,N_7555,N_7404);
or U7779 (N_7779,N_7551,N_7484);
or U7780 (N_7780,N_7445,N_7515);
nand U7781 (N_7781,N_7504,N_7535);
and U7782 (N_7782,N_7581,N_7587);
or U7783 (N_7783,N_7548,N_7500);
nor U7784 (N_7784,N_7599,N_7567);
xor U7785 (N_7785,N_7549,N_7572);
or U7786 (N_7786,N_7400,N_7426);
nor U7787 (N_7787,N_7545,N_7423);
nand U7788 (N_7788,N_7593,N_7450);
nand U7789 (N_7789,N_7481,N_7402);
or U7790 (N_7790,N_7502,N_7432);
or U7791 (N_7791,N_7439,N_7489);
nor U7792 (N_7792,N_7492,N_7440);
nor U7793 (N_7793,N_7447,N_7473);
nor U7794 (N_7794,N_7543,N_7470);
and U7795 (N_7795,N_7581,N_7572);
nor U7796 (N_7796,N_7508,N_7484);
xor U7797 (N_7797,N_7478,N_7557);
nand U7798 (N_7798,N_7526,N_7596);
nand U7799 (N_7799,N_7459,N_7558);
nor U7800 (N_7800,N_7747,N_7749);
or U7801 (N_7801,N_7645,N_7796);
nor U7802 (N_7802,N_7762,N_7672);
nand U7803 (N_7803,N_7681,N_7707);
xor U7804 (N_7804,N_7760,N_7612);
nand U7805 (N_7805,N_7710,N_7785);
xnor U7806 (N_7806,N_7642,N_7618);
and U7807 (N_7807,N_7669,N_7781);
xor U7808 (N_7808,N_7696,N_7697);
xor U7809 (N_7809,N_7630,N_7606);
nand U7810 (N_7810,N_7691,N_7634);
nand U7811 (N_7811,N_7671,N_7713);
and U7812 (N_7812,N_7718,N_7687);
nor U7813 (N_7813,N_7735,N_7779);
and U7814 (N_7814,N_7641,N_7680);
nor U7815 (N_7815,N_7695,N_7655);
or U7816 (N_7816,N_7614,N_7782);
or U7817 (N_7817,N_7776,N_7715);
or U7818 (N_7818,N_7616,N_7739);
and U7819 (N_7819,N_7602,N_7656);
nor U7820 (N_7820,N_7643,N_7704);
or U7821 (N_7821,N_7756,N_7682);
xnor U7822 (N_7822,N_7726,N_7702);
or U7823 (N_7823,N_7744,N_7733);
nor U7824 (N_7824,N_7665,N_7632);
xor U7825 (N_7825,N_7738,N_7627);
and U7826 (N_7826,N_7652,N_7668);
and U7827 (N_7827,N_7727,N_7651);
nor U7828 (N_7828,N_7629,N_7615);
nand U7829 (N_7829,N_7748,N_7678);
or U7830 (N_7830,N_7646,N_7676);
and U7831 (N_7831,N_7664,N_7663);
nor U7832 (N_7832,N_7732,N_7712);
nor U7833 (N_7833,N_7633,N_7777);
and U7834 (N_7834,N_7650,N_7638);
nor U7835 (N_7835,N_7609,N_7767);
and U7836 (N_7836,N_7684,N_7639);
or U7837 (N_7837,N_7689,N_7619);
nor U7838 (N_7838,N_7795,N_7750);
nand U7839 (N_7839,N_7716,N_7608);
nor U7840 (N_7840,N_7741,N_7620);
or U7841 (N_7841,N_7723,N_7765);
xnor U7842 (N_7842,N_7690,N_7783);
xnor U7843 (N_7843,N_7728,N_7610);
or U7844 (N_7844,N_7692,N_7754);
xnor U7845 (N_7845,N_7709,N_7662);
nand U7846 (N_7846,N_7628,N_7794);
nand U7847 (N_7847,N_7724,N_7657);
or U7848 (N_7848,N_7721,N_7667);
nand U7849 (N_7849,N_7771,N_7737);
nor U7850 (N_7850,N_7604,N_7694);
or U7851 (N_7851,N_7780,N_7648);
nor U7852 (N_7852,N_7775,N_7778);
nand U7853 (N_7853,N_7725,N_7736);
nor U7854 (N_7854,N_7635,N_7770);
nor U7855 (N_7855,N_7761,N_7623);
nand U7856 (N_7856,N_7729,N_7647);
xor U7857 (N_7857,N_7685,N_7603);
and U7858 (N_7858,N_7640,N_7799);
or U7859 (N_7859,N_7720,N_7746);
nor U7860 (N_7860,N_7637,N_7624);
and U7861 (N_7861,N_7757,N_7607);
and U7862 (N_7862,N_7714,N_7769);
nand U7863 (N_7863,N_7792,N_7742);
xnor U7864 (N_7864,N_7743,N_7772);
nor U7865 (N_7865,N_7740,N_7717);
nor U7866 (N_7866,N_7673,N_7791);
nor U7867 (N_7867,N_7631,N_7686);
nor U7868 (N_7868,N_7751,N_7730);
or U7869 (N_7869,N_7763,N_7753);
and U7870 (N_7870,N_7711,N_7764);
nand U7871 (N_7871,N_7659,N_7773);
nand U7872 (N_7872,N_7605,N_7788);
and U7873 (N_7873,N_7797,N_7679);
or U7874 (N_7874,N_7613,N_7699);
or U7875 (N_7875,N_7731,N_7706);
and U7876 (N_7876,N_7705,N_7752);
and U7877 (N_7877,N_7677,N_7768);
nand U7878 (N_7878,N_7674,N_7701);
nor U7879 (N_7879,N_7789,N_7719);
or U7880 (N_7880,N_7601,N_7621);
and U7881 (N_7881,N_7766,N_7653);
nand U7882 (N_7882,N_7658,N_7722);
and U7883 (N_7883,N_7622,N_7644);
xor U7884 (N_7884,N_7626,N_7600);
or U7885 (N_7885,N_7703,N_7611);
nand U7886 (N_7886,N_7675,N_7625);
xor U7887 (N_7887,N_7698,N_7693);
nor U7888 (N_7888,N_7787,N_7790);
nor U7889 (N_7889,N_7700,N_7758);
nor U7890 (N_7890,N_7708,N_7661);
or U7891 (N_7891,N_7666,N_7784);
nand U7892 (N_7892,N_7755,N_7649);
or U7893 (N_7893,N_7793,N_7774);
xnor U7894 (N_7894,N_7786,N_7745);
nand U7895 (N_7895,N_7660,N_7683);
nor U7896 (N_7896,N_7654,N_7734);
nor U7897 (N_7897,N_7688,N_7636);
nor U7898 (N_7898,N_7670,N_7759);
and U7899 (N_7899,N_7798,N_7617);
nor U7900 (N_7900,N_7765,N_7767);
and U7901 (N_7901,N_7608,N_7665);
nand U7902 (N_7902,N_7737,N_7708);
nand U7903 (N_7903,N_7695,N_7706);
and U7904 (N_7904,N_7712,N_7668);
nor U7905 (N_7905,N_7777,N_7787);
nand U7906 (N_7906,N_7715,N_7670);
xor U7907 (N_7907,N_7728,N_7791);
and U7908 (N_7908,N_7733,N_7616);
nor U7909 (N_7909,N_7658,N_7624);
and U7910 (N_7910,N_7712,N_7650);
nand U7911 (N_7911,N_7672,N_7620);
nand U7912 (N_7912,N_7756,N_7692);
or U7913 (N_7913,N_7666,N_7637);
xnor U7914 (N_7914,N_7718,N_7659);
and U7915 (N_7915,N_7715,N_7772);
nor U7916 (N_7916,N_7728,N_7660);
or U7917 (N_7917,N_7770,N_7725);
or U7918 (N_7918,N_7763,N_7610);
nor U7919 (N_7919,N_7685,N_7734);
nor U7920 (N_7920,N_7739,N_7755);
xnor U7921 (N_7921,N_7668,N_7682);
nor U7922 (N_7922,N_7624,N_7733);
and U7923 (N_7923,N_7637,N_7753);
and U7924 (N_7924,N_7647,N_7666);
nand U7925 (N_7925,N_7605,N_7643);
nor U7926 (N_7926,N_7732,N_7773);
xor U7927 (N_7927,N_7784,N_7735);
and U7928 (N_7928,N_7629,N_7775);
nor U7929 (N_7929,N_7642,N_7613);
nor U7930 (N_7930,N_7616,N_7603);
or U7931 (N_7931,N_7682,N_7700);
nand U7932 (N_7932,N_7793,N_7719);
and U7933 (N_7933,N_7790,N_7697);
nand U7934 (N_7934,N_7662,N_7698);
nor U7935 (N_7935,N_7655,N_7776);
nor U7936 (N_7936,N_7733,N_7675);
and U7937 (N_7937,N_7655,N_7787);
xnor U7938 (N_7938,N_7632,N_7757);
or U7939 (N_7939,N_7630,N_7770);
nand U7940 (N_7940,N_7681,N_7777);
or U7941 (N_7941,N_7694,N_7674);
nand U7942 (N_7942,N_7655,N_7798);
or U7943 (N_7943,N_7618,N_7612);
or U7944 (N_7944,N_7750,N_7712);
nand U7945 (N_7945,N_7678,N_7657);
or U7946 (N_7946,N_7659,N_7676);
xor U7947 (N_7947,N_7768,N_7702);
or U7948 (N_7948,N_7733,N_7734);
or U7949 (N_7949,N_7638,N_7718);
nand U7950 (N_7950,N_7773,N_7783);
xnor U7951 (N_7951,N_7741,N_7734);
nand U7952 (N_7952,N_7611,N_7780);
or U7953 (N_7953,N_7754,N_7718);
nand U7954 (N_7954,N_7600,N_7795);
and U7955 (N_7955,N_7650,N_7798);
nand U7956 (N_7956,N_7756,N_7745);
nand U7957 (N_7957,N_7762,N_7736);
nor U7958 (N_7958,N_7689,N_7707);
and U7959 (N_7959,N_7724,N_7660);
or U7960 (N_7960,N_7700,N_7710);
nor U7961 (N_7961,N_7708,N_7629);
nor U7962 (N_7962,N_7736,N_7657);
xor U7963 (N_7963,N_7622,N_7767);
or U7964 (N_7964,N_7718,N_7676);
nand U7965 (N_7965,N_7693,N_7681);
nor U7966 (N_7966,N_7786,N_7610);
nor U7967 (N_7967,N_7769,N_7605);
xnor U7968 (N_7968,N_7725,N_7735);
xnor U7969 (N_7969,N_7718,N_7796);
nand U7970 (N_7970,N_7760,N_7628);
xor U7971 (N_7971,N_7694,N_7631);
and U7972 (N_7972,N_7750,N_7691);
nor U7973 (N_7973,N_7748,N_7740);
nand U7974 (N_7974,N_7602,N_7661);
and U7975 (N_7975,N_7746,N_7721);
nand U7976 (N_7976,N_7642,N_7718);
nor U7977 (N_7977,N_7723,N_7629);
nand U7978 (N_7978,N_7792,N_7631);
and U7979 (N_7979,N_7698,N_7784);
and U7980 (N_7980,N_7664,N_7766);
and U7981 (N_7981,N_7654,N_7662);
or U7982 (N_7982,N_7719,N_7730);
nand U7983 (N_7983,N_7675,N_7640);
xor U7984 (N_7984,N_7644,N_7616);
and U7985 (N_7985,N_7603,N_7645);
nor U7986 (N_7986,N_7786,N_7775);
and U7987 (N_7987,N_7685,N_7666);
nor U7988 (N_7988,N_7742,N_7695);
nor U7989 (N_7989,N_7795,N_7722);
xnor U7990 (N_7990,N_7641,N_7612);
nand U7991 (N_7991,N_7781,N_7653);
nand U7992 (N_7992,N_7708,N_7743);
xnor U7993 (N_7993,N_7624,N_7638);
or U7994 (N_7994,N_7741,N_7630);
xor U7995 (N_7995,N_7749,N_7712);
and U7996 (N_7996,N_7641,N_7684);
nand U7997 (N_7997,N_7744,N_7653);
nand U7998 (N_7998,N_7690,N_7795);
nand U7999 (N_7999,N_7698,N_7786);
xor U8000 (N_8000,N_7948,N_7819);
xnor U8001 (N_8001,N_7915,N_7918);
nor U8002 (N_8002,N_7837,N_7891);
nor U8003 (N_8003,N_7929,N_7821);
nor U8004 (N_8004,N_7909,N_7825);
xnor U8005 (N_8005,N_7973,N_7840);
xor U8006 (N_8006,N_7863,N_7861);
or U8007 (N_8007,N_7830,N_7803);
nor U8008 (N_8008,N_7910,N_7903);
xnor U8009 (N_8009,N_7969,N_7848);
xor U8010 (N_8010,N_7913,N_7866);
or U8011 (N_8011,N_7995,N_7912);
or U8012 (N_8012,N_7914,N_7998);
nand U8013 (N_8013,N_7824,N_7854);
nor U8014 (N_8014,N_7972,N_7906);
or U8015 (N_8015,N_7942,N_7927);
xor U8016 (N_8016,N_7981,N_7957);
or U8017 (N_8017,N_7958,N_7931);
nor U8018 (N_8018,N_7908,N_7823);
nand U8019 (N_8019,N_7939,N_7999);
xnor U8020 (N_8020,N_7952,N_7932);
nand U8021 (N_8021,N_7874,N_7851);
nand U8022 (N_8022,N_7826,N_7916);
nor U8023 (N_8023,N_7983,N_7880);
nor U8024 (N_8024,N_7868,N_7871);
nor U8025 (N_8025,N_7835,N_7945);
xnor U8026 (N_8026,N_7977,N_7856);
nor U8027 (N_8027,N_7917,N_7971);
nor U8028 (N_8028,N_7941,N_7859);
and U8029 (N_8029,N_7831,N_7961);
nor U8030 (N_8030,N_7838,N_7934);
and U8031 (N_8031,N_7814,N_7959);
nand U8032 (N_8032,N_7907,N_7935);
nor U8033 (N_8033,N_7855,N_7895);
or U8034 (N_8034,N_7872,N_7889);
xor U8035 (N_8035,N_7944,N_7844);
or U8036 (N_8036,N_7853,N_7873);
nand U8037 (N_8037,N_7922,N_7923);
and U8038 (N_8038,N_7834,N_7994);
nand U8039 (N_8039,N_7996,N_7955);
nand U8040 (N_8040,N_7887,N_7810);
nor U8041 (N_8041,N_7888,N_7954);
or U8042 (N_8042,N_7806,N_7883);
or U8043 (N_8043,N_7841,N_7911);
and U8044 (N_8044,N_7839,N_7843);
or U8045 (N_8045,N_7886,N_7978);
and U8046 (N_8046,N_7898,N_7930);
and U8047 (N_8047,N_7811,N_7885);
nand U8048 (N_8048,N_7893,N_7882);
nand U8049 (N_8049,N_7997,N_7902);
and U8050 (N_8050,N_7860,N_7901);
or U8051 (N_8051,N_7986,N_7818);
nand U8052 (N_8052,N_7822,N_7966);
nand U8053 (N_8053,N_7991,N_7896);
nand U8054 (N_8054,N_7992,N_7867);
nor U8055 (N_8055,N_7805,N_7963);
xor U8056 (N_8056,N_7812,N_7970);
and U8057 (N_8057,N_7960,N_7985);
nor U8058 (N_8058,N_7864,N_7975);
nor U8059 (N_8059,N_7919,N_7881);
xor U8060 (N_8060,N_7925,N_7849);
and U8061 (N_8061,N_7968,N_7946);
and U8062 (N_8062,N_7802,N_7842);
or U8063 (N_8063,N_7890,N_7852);
xnor U8064 (N_8064,N_7984,N_7921);
or U8065 (N_8065,N_7979,N_7832);
or U8066 (N_8066,N_7982,N_7928);
xor U8067 (N_8067,N_7894,N_7878);
or U8068 (N_8068,N_7956,N_7884);
or U8069 (N_8069,N_7924,N_7950);
and U8070 (N_8070,N_7967,N_7857);
and U8071 (N_8071,N_7949,N_7804);
xnor U8072 (N_8072,N_7936,N_7808);
nand U8073 (N_8073,N_7836,N_7877);
nor U8074 (N_8074,N_7989,N_7827);
nor U8075 (N_8075,N_7899,N_7962);
nand U8076 (N_8076,N_7865,N_7829);
xnor U8077 (N_8077,N_7801,N_7879);
xnor U8078 (N_8078,N_7862,N_7870);
nor U8079 (N_8079,N_7875,N_7987);
nand U8080 (N_8080,N_7828,N_7892);
nor U8081 (N_8081,N_7807,N_7953);
nand U8082 (N_8082,N_7817,N_7974);
xor U8083 (N_8083,N_7816,N_7976);
nor U8084 (N_8084,N_7858,N_7951);
and U8085 (N_8085,N_7943,N_7937);
nand U8086 (N_8086,N_7933,N_7965);
or U8087 (N_8087,N_7940,N_7938);
xor U8088 (N_8088,N_7920,N_7850);
xor U8089 (N_8089,N_7993,N_7869);
xnor U8090 (N_8090,N_7897,N_7905);
and U8091 (N_8091,N_7990,N_7833);
xor U8092 (N_8092,N_7815,N_7876);
or U8093 (N_8093,N_7980,N_7900);
and U8094 (N_8094,N_7800,N_7846);
and U8095 (N_8095,N_7964,N_7926);
or U8096 (N_8096,N_7947,N_7847);
or U8097 (N_8097,N_7988,N_7845);
nand U8098 (N_8098,N_7809,N_7904);
and U8099 (N_8099,N_7813,N_7820);
nor U8100 (N_8100,N_7969,N_7965);
or U8101 (N_8101,N_7949,N_7983);
xnor U8102 (N_8102,N_7831,N_7860);
xnor U8103 (N_8103,N_7937,N_7986);
or U8104 (N_8104,N_7910,N_7936);
nand U8105 (N_8105,N_7937,N_7907);
and U8106 (N_8106,N_7846,N_7953);
nand U8107 (N_8107,N_7855,N_7961);
xnor U8108 (N_8108,N_7970,N_7960);
or U8109 (N_8109,N_7906,N_7823);
and U8110 (N_8110,N_7838,N_7885);
or U8111 (N_8111,N_7921,N_7885);
or U8112 (N_8112,N_7976,N_7928);
nor U8113 (N_8113,N_7838,N_7845);
or U8114 (N_8114,N_7856,N_7967);
xnor U8115 (N_8115,N_7840,N_7864);
nor U8116 (N_8116,N_7850,N_7962);
xnor U8117 (N_8117,N_7985,N_7841);
nor U8118 (N_8118,N_7869,N_7914);
and U8119 (N_8119,N_7831,N_7826);
xor U8120 (N_8120,N_7805,N_7894);
xor U8121 (N_8121,N_7971,N_7895);
nor U8122 (N_8122,N_7922,N_7976);
or U8123 (N_8123,N_7843,N_7818);
nand U8124 (N_8124,N_7800,N_7923);
nand U8125 (N_8125,N_7918,N_7851);
and U8126 (N_8126,N_7911,N_7957);
or U8127 (N_8127,N_7864,N_7836);
nand U8128 (N_8128,N_7954,N_7920);
nand U8129 (N_8129,N_7997,N_7852);
xor U8130 (N_8130,N_7941,N_7830);
and U8131 (N_8131,N_7860,N_7978);
or U8132 (N_8132,N_7818,N_7985);
xnor U8133 (N_8133,N_7823,N_7990);
or U8134 (N_8134,N_7922,N_7810);
nand U8135 (N_8135,N_7845,N_7990);
nand U8136 (N_8136,N_7907,N_7943);
or U8137 (N_8137,N_7972,N_7965);
and U8138 (N_8138,N_7830,N_7921);
and U8139 (N_8139,N_7974,N_7859);
or U8140 (N_8140,N_7922,N_7882);
and U8141 (N_8141,N_7884,N_7861);
nand U8142 (N_8142,N_7824,N_7972);
or U8143 (N_8143,N_7905,N_7826);
and U8144 (N_8144,N_7952,N_7974);
nand U8145 (N_8145,N_7964,N_7914);
xor U8146 (N_8146,N_7997,N_7803);
nor U8147 (N_8147,N_7940,N_7873);
nor U8148 (N_8148,N_7924,N_7839);
xnor U8149 (N_8149,N_7920,N_7962);
and U8150 (N_8150,N_7919,N_7874);
xor U8151 (N_8151,N_7837,N_7974);
nand U8152 (N_8152,N_7941,N_7946);
and U8153 (N_8153,N_7992,N_7934);
or U8154 (N_8154,N_7819,N_7989);
xor U8155 (N_8155,N_7985,N_7894);
nor U8156 (N_8156,N_7877,N_7912);
nand U8157 (N_8157,N_7981,N_7963);
or U8158 (N_8158,N_7995,N_7813);
or U8159 (N_8159,N_7926,N_7952);
or U8160 (N_8160,N_7878,N_7879);
or U8161 (N_8161,N_7849,N_7844);
nand U8162 (N_8162,N_7929,N_7970);
xor U8163 (N_8163,N_7872,N_7842);
and U8164 (N_8164,N_7890,N_7933);
or U8165 (N_8165,N_7909,N_7863);
nor U8166 (N_8166,N_7968,N_7986);
or U8167 (N_8167,N_7826,N_7833);
nor U8168 (N_8168,N_7902,N_7853);
nor U8169 (N_8169,N_7872,N_7849);
nor U8170 (N_8170,N_7818,N_7971);
nand U8171 (N_8171,N_7962,N_7829);
and U8172 (N_8172,N_7954,N_7866);
nor U8173 (N_8173,N_7806,N_7826);
nor U8174 (N_8174,N_7823,N_7842);
or U8175 (N_8175,N_7808,N_7982);
nand U8176 (N_8176,N_7807,N_7877);
or U8177 (N_8177,N_7946,N_7898);
nand U8178 (N_8178,N_7937,N_7985);
xor U8179 (N_8179,N_7870,N_7809);
xnor U8180 (N_8180,N_7949,N_7817);
xor U8181 (N_8181,N_7954,N_7941);
or U8182 (N_8182,N_7806,N_7831);
nand U8183 (N_8183,N_7844,N_7907);
or U8184 (N_8184,N_7800,N_7810);
nor U8185 (N_8185,N_7957,N_7985);
nand U8186 (N_8186,N_7946,N_7809);
and U8187 (N_8187,N_7985,N_7895);
xnor U8188 (N_8188,N_7971,N_7893);
nand U8189 (N_8189,N_7877,N_7921);
nand U8190 (N_8190,N_7996,N_7983);
or U8191 (N_8191,N_7814,N_7895);
nor U8192 (N_8192,N_7814,N_7853);
nand U8193 (N_8193,N_7939,N_7899);
nor U8194 (N_8194,N_7980,N_7992);
and U8195 (N_8195,N_7979,N_7950);
xor U8196 (N_8196,N_7963,N_7978);
xor U8197 (N_8197,N_7934,N_7998);
nor U8198 (N_8198,N_7897,N_7966);
or U8199 (N_8199,N_7900,N_7878);
and U8200 (N_8200,N_8145,N_8090);
and U8201 (N_8201,N_8189,N_8185);
and U8202 (N_8202,N_8110,N_8141);
nor U8203 (N_8203,N_8190,N_8142);
nand U8204 (N_8204,N_8046,N_8114);
nor U8205 (N_8205,N_8057,N_8162);
xnor U8206 (N_8206,N_8058,N_8135);
or U8207 (N_8207,N_8080,N_8188);
xnor U8208 (N_8208,N_8035,N_8075);
xnor U8209 (N_8209,N_8106,N_8086);
and U8210 (N_8210,N_8164,N_8175);
and U8211 (N_8211,N_8138,N_8006);
or U8212 (N_8212,N_8176,N_8115);
and U8213 (N_8213,N_8036,N_8137);
nor U8214 (N_8214,N_8128,N_8179);
xor U8215 (N_8215,N_8074,N_8082);
nand U8216 (N_8216,N_8043,N_8184);
nand U8217 (N_8217,N_8178,N_8024);
nand U8218 (N_8218,N_8194,N_8060);
and U8219 (N_8219,N_8026,N_8186);
or U8220 (N_8220,N_8119,N_8032);
nand U8221 (N_8221,N_8061,N_8102);
xor U8222 (N_8222,N_8149,N_8052);
xnor U8223 (N_8223,N_8008,N_8195);
nand U8224 (N_8224,N_8017,N_8103);
nand U8225 (N_8225,N_8156,N_8023);
nand U8226 (N_8226,N_8171,N_8177);
and U8227 (N_8227,N_8012,N_8019);
nor U8228 (N_8228,N_8199,N_8126);
nand U8229 (N_8229,N_8042,N_8161);
nand U8230 (N_8230,N_8187,N_8085);
nand U8231 (N_8231,N_8091,N_8140);
nand U8232 (N_8232,N_8084,N_8097);
nand U8233 (N_8233,N_8117,N_8100);
or U8234 (N_8234,N_8131,N_8143);
nand U8235 (N_8235,N_8116,N_8122);
and U8236 (N_8236,N_8007,N_8013);
nand U8237 (N_8237,N_8120,N_8112);
nor U8238 (N_8238,N_8144,N_8160);
nand U8239 (N_8239,N_8172,N_8173);
nor U8240 (N_8240,N_8051,N_8124);
or U8241 (N_8241,N_8053,N_8081);
or U8242 (N_8242,N_8147,N_8154);
nor U8243 (N_8243,N_8113,N_8004);
xor U8244 (N_8244,N_8015,N_8001);
nand U8245 (N_8245,N_8034,N_8041);
or U8246 (N_8246,N_8157,N_8105);
nand U8247 (N_8247,N_8093,N_8067);
nand U8248 (N_8248,N_8045,N_8155);
xor U8249 (N_8249,N_8159,N_8166);
xnor U8250 (N_8250,N_8072,N_8158);
nor U8251 (N_8251,N_8170,N_8066);
nand U8252 (N_8252,N_8014,N_8197);
nand U8253 (N_8253,N_8181,N_8063);
or U8254 (N_8254,N_8183,N_8054);
xor U8255 (N_8255,N_8064,N_8071);
or U8256 (N_8256,N_8139,N_8065);
or U8257 (N_8257,N_8022,N_8132);
nand U8258 (N_8258,N_8136,N_8068);
or U8259 (N_8259,N_8076,N_8088);
or U8260 (N_8260,N_8033,N_8109);
or U8261 (N_8261,N_8062,N_8020);
or U8262 (N_8262,N_8130,N_8069);
nor U8263 (N_8263,N_8168,N_8134);
or U8264 (N_8264,N_8005,N_8010);
xor U8265 (N_8265,N_8098,N_8125);
and U8266 (N_8266,N_8038,N_8002);
or U8267 (N_8267,N_8055,N_8031);
or U8268 (N_8268,N_8027,N_8167);
and U8269 (N_8269,N_8095,N_8087);
nand U8270 (N_8270,N_8030,N_8191);
nor U8271 (N_8271,N_8169,N_8083);
and U8272 (N_8272,N_8073,N_8044);
nand U8273 (N_8273,N_8040,N_8107);
xor U8274 (N_8274,N_8152,N_8011);
nand U8275 (N_8275,N_8099,N_8111);
nand U8276 (N_8276,N_8070,N_8000);
nand U8277 (N_8277,N_8079,N_8089);
or U8278 (N_8278,N_8193,N_8163);
and U8279 (N_8279,N_8092,N_8118);
or U8280 (N_8280,N_8133,N_8021);
and U8281 (N_8281,N_8146,N_8028);
or U8282 (N_8282,N_8094,N_8196);
or U8283 (N_8283,N_8148,N_8096);
nor U8284 (N_8284,N_8180,N_8037);
xor U8285 (N_8285,N_8025,N_8129);
and U8286 (N_8286,N_8047,N_8003);
xor U8287 (N_8287,N_8123,N_8150);
xnor U8288 (N_8288,N_8108,N_8059);
or U8289 (N_8289,N_8153,N_8121);
xor U8290 (N_8290,N_8165,N_8018);
xnor U8291 (N_8291,N_8174,N_8056);
nor U8292 (N_8292,N_8048,N_8049);
nor U8293 (N_8293,N_8104,N_8016);
and U8294 (N_8294,N_8078,N_8151);
or U8295 (N_8295,N_8127,N_8009);
xnor U8296 (N_8296,N_8050,N_8182);
nand U8297 (N_8297,N_8198,N_8192);
nor U8298 (N_8298,N_8101,N_8029);
nand U8299 (N_8299,N_8039,N_8077);
and U8300 (N_8300,N_8079,N_8132);
xnor U8301 (N_8301,N_8180,N_8089);
nor U8302 (N_8302,N_8082,N_8083);
and U8303 (N_8303,N_8047,N_8107);
xnor U8304 (N_8304,N_8056,N_8019);
or U8305 (N_8305,N_8108,N_8183);
and U8306 (N_8306,N_8021,N_8025);
nand U8307 (N_8307,N_8080,N_8008);
and U8308 (N_8308,N_8029,N_8144);
nand U8309 (N_8309,N_8004,N_8164);
nor U8310 (N_8310,N_8010,N_8045);
and U8311 (N_8311,N_8039,N_8170);
nand U8312 (N_8312,N_8086,N_8021);
nand U8313 (N_8313,N_8052,N_8154);
xor U8314 (N_8314,N_8153,N_8126);
or U8315 (N_8315,N_8071,N_8162);
and U8316 (N_8316,N_8031,N_8092);
and U8317 (N_8317,N_8083,N_8076);
xor U8318 (N_8318,N_8180,N_8072);
nand U8319 (N_8319,N_8046,N_8075);
or U8320 (N_8320,N_8141,N_8076);
nor U8321 (N_8321,N_8089,N_8183);
or U8322 (N_8322,N_8102,N_8118);
or U8323 (N_8323,N_8044,N_8095);
and U8324 (N_8324,N_8059,N_8080);
or U8325 (N_8325,N_8016,N_8145);
nor U8326 (N_8326,N_8120,N_8011);
and U8327 (N_8327,N_8193,N_8022);
xor U8328 (N_8328,N_8080,N_8051);
or U8329 (N_8329,N_8145,N_8005);
and U8330 (N_8330,N_8060,N_8077);
nor U8331 (N_8331,N_8033,N_8030);
nor U8332 (N_8332,N_8158,N_8052);
or U8333 (N_8333,N_8120,N_8134);
nand U8334 (N_8334,N_8005,N_8049);
nand U8335 (N_8335,N_8131,N_8053);
xnor U8336 (N_8336,N_8185,N_8033);
or U8337 (N_8337,N_8055,N_8113);
and U8338 (N_8338,N_8176,N_8000);
xnor U8339 (N_8339,N_8041,N_8021);
nand U8340 (N_8340,N_8175,N_8061);
and U8341 (N_8341,N_8040,N_8111);
nand U8342 (N_8342,N_8196,N_8088);
nor U8343 (N_8343,N_8157,N_8164);
or U8344 (N_8344,N_8001,N_8168);
xor U8345 (N_8345,N_8051,N_8116);
or U8346 (N_8346,N_8053,N_8174);
nor U8347 (N_8347,N_8098,N_8184);
and U8348 (N_8348,N_8189,N_8090);
or U8349 (N_8349,N_8114,N_8068);
or U8350 (N_8350,N_8068,N_8133);
and U8351 (N_8351,N_8161,N_8077);
or U8352 (N_8352,N_8135,N_8068);
and U8353 (N_8353,N_8155,N_8197);
xnor U8354 (N_8354,N_8081,N_8006);
nand U8355 (N_8355,N_8055,N_8077);
xor U8356 (N_8356,N_8172,N_8020);
and U8357 (N_8357,N_8072,N_8054);
nor U8358 (N_8358,N_8135,N_8094);
nor U8359 (N_8359,N_8156,N_8064);
xor U8360 (N_8360,N_8172,N_8001);
and U8361 (N_8361,N_8008,N_8194);
xnor U8362 (N_8362,N_8164,N_8029);
and U8363 (N_8363,N_8121,N_8114);
nor U8364 (N_8364,N_8014,N_8020);
xnor U8365 (N_8365,N_8195,N_8192);
or U8366 (N_8366,N_8095,N_8110);
or U8367 (N_8367,N_8172,N_8168);
xnor U8368 (N_8368,N_8199,N_8185);
xor U8369 (N_8369,N_8188,N_8085);
and U8370 (N_8370,N_8006,N_8164);
xnor U8371 (N_8371,N_8064,N_8181);
or U8372 (N_8372,N_8024,N_8086);
or U8373 (N_8373,N_8020,N_8029);
xor U8374 (N_8374,N_8097,N_8159);
xnor U8375 (N_8375,N_8011,N_8196);
or U8376 (N_8376,N_8048,N_8084);
xnor U8377 (N_8377,N_8091,N_8038);
and U8378 (N_8378,N_8087,N_8074);
nor U8379 (N_8379,N_8157,N_8112);
or U8380 (N_8380,N_8133,N_8152);
or U8381 (N_8381,N_8159,N_8000);
xnor U8382 (N_8382,N_8082,N_8193);
nor U8383 (N_8383,N_8016,N_8181);
or U8384 (N_8384,N_8182,N_8143);
xnor U8385 (N_8385,N_8051,N_8180);
xor U8386 (N_8386,N_8092,N_8008);
xnor U8387 (N_8387,N_8024,N_8018);
xor U8388 (N_8388,N_8002,N_8144);
nand U8389 (N_8389,N_8110,N_8111);
or U8390 (N_8390,N_8122,N_8051);
nand U8391 (N_8391,N_8051,N_8175);
or U8392 (N_8392,N_8157,N_8142);
nand U8393 (N_8393,N_8084,N_8043);
xnor U8394 (N_8394,N_8175,N_8082);
or U8395 (N_8395,N_8197,N_8150);
and U8396 (N_8396,N_8040,N_8150);
and U8397 (N_8397,N_8123,N_8122);
xnor U8398 (N_8398,N_8152,N_8039);
nor U8399 (N_8399,N_8193,N_8053);
nor U8400 (N_8400,N_8202,N_8220);
nor U8401 (N_8401,N_8230,N_8319);
nand U8402 (N_8402,N_8381,N_8373);
nand U8403 (N_8403,N_8379,N_8238);
and U8404 (N_8404,N_8310,N_8217);
xor U8405 (N_8405,N_8371,N_8313);
xnor U8406 (N_8406,N_8392,N_8352);
nand U8407 (N_8407,N_8272,N_8232);
nor U8408 (N_8408,N_8299,N_8209);
or U8409 (N_8409,N_8341,N_8262);
or U8410 (N_8410,N_8354,N_8334);
xor U8411 (N_8411,N_8276,N_8387);
or U8412 (N_8412,N_8203,N_8236);
or U8413 (N_8413,N_8256,N_8382);
xor U8414 (N_8414,N_8287,N_8370);
nand U8415 (N_8415,N_8211,N_8305);
xor U8416 (N_8416,N_8391,N_8216);
xnor U8417 (N_8417,N_8350,N_8246);
nand U8418 (N_8418,N_8268,N_8207);
and U8419 (N_8419,N_8286,N_8339);
nand U8420 (N_8420,N_8367,N_8386);
nor U8421 (N_8421,N_8285,N_8227);
and U8422 (N_8422,N_8320,N_8298);
nand U8423 (N_8423,N_8214,N_8250);
or U8424 (N_8424,N_8326,N_8377);
xnor U8425 (N_8425,N_8331,N_8342);
and U8426 (N_8426,N_8212,N_8266);
or U8427 (N_8427,N_8255,N_8210);
nand U8428 (N_8428,N_8237,N_8396);
or U8429 (N_8429,N_8308,N_8275);
nor U8430 (N_8430,N_8361,N_8395);
nand U8431 (N_8431,N_8380,N_8221);
xor U8432 (N_8432,N_8228,N_8300);
nand U8433 (N_8433,N_8355,N_8394);
or U8434 (N_8434,N_8316,N_8325);
nand U8435 (N_8435,N_8281,N_8399);
and U8436 (N_8436,N_8231,N_8271);
xnor U8437 (N_8437,N_8233,N_8208);
nor U8438 (N_8438,N_8296,N_8254);
or U8439 (N_8439,N_8234,N_8329);
and U8440 (N_8440,N_8259,N_8279);
nor U8441 (N_8441,N_8359,N_8364);
and U8442 (N_8442,N_8384,N_8332);
nor U8443 (N_8443,N_8274,N_8290);
and U8444 (N_8444,N_8390,N_8306);
nand U8445 (N_8445,N_8204,N_8337);
xnor U8446 (N_8446,N_8340,N_8249);
and U8447 (N_8447,N_8215,N_8330);
nand U8448 (N_8448,N_8303,N_8376);
nand U8449 (N_8449,N_8218,N_8369);
nor U8450 (N_8450,N_8283,N_8309);
nand U8451 (N_8451,N_8317,N_8294);
xnor U8452 (N_8452,N_8229,N_8366);
xor U8453 (N_8453,N_8240,N_8345);
nand U8454 (N_8454,N_8343,N_8318);
nor U8455 (N_8455,N_8239,N_8200);
nor U8456 (N_8456,N_8321,N_8213);
or U8457 (N_8457,N_8324,N_8327);
nor U8458 (N_8458,N_8224,N_8336);
or U8459 (N_8459,N_8263,N_8261);
nand U8460 (N_8460,N_8235,N_8292);
nand U8461 (N_8461,N_8226,N_8247);
or U8462 (N_8462,N_8280,N_8362);
xnor U8463 (N_8463,N_8270,N_8388);
nor U8464 (N_8464,N_8284,N_8314);
nand U8465 (N_8465,N_8248,N_8222);
or U8466 (N_8466,N_8273,N_8282);
nand U8467 (N_8467,N_8397,N_8257);
and U8468 (N_8468,N_8265,N_8244);
nor U8469 (N_8469,N_8347,N_8251);
and U8470 (N_8470,N_8378,N_8252);
xnor U8471 (N_8471,N_8335,N_8385);
xnor U8472 (N_8472,N_8242,N_8289);
nand U8473 (N_8473,N_8383,N_8302);
and U8474 (N_8474,N_8293,N_8368);
xnor U8475 (N_8475,N_8338,N_8398);
nand U8476 (N_8476,N_8219,N_8297);
xnor U8477 (N_8477,N_8225,N_8288);
or U8478 (N_8478,N_8357,N_8269);
xor U8479 (N_8479,N_8264,N_8328);
xnor U8480 (N_8480,N_8253,N_8349);
nand U8481 (N_8481,N_8333,N_8365);
nand U8482 (N_8482,N_8241,N_8277);
or U8483 (N_8483,N_8201,N_8356);
nand U8484 (N_8484,N_8351,N_8312);
nand U8485 (N_8485,N_8393,N_8243);
xor U8486 (N_8486,N_8348,N_8360);
and U8487 (N_8487,N_8375,N_8260);
xor U8488 (N_8488,N_8223,N_8315);
nor U8489 (N_8489,N_8267,N_8353);
or U8490 (N_8490,N_8206,N_8374);
or U8491 (N_8491,N_8291,N_8301);
xor U8492 (N_8492,N_8344,N_8363);
xnor U8493 (N_8493,N_8295,N_8278);
and U8494 (N_8494,N_8205,N_8258);
xor U8495 (N_8495,N_8346,N_8372);
nand U8496 (N_8496,N_8389,N_8307);
xnor U8497 (N_8497,N_8245,N_8304);
nand U8498 (N_8498,N_8323,N_8311);
and U8499 (N_8499,N_8322,N_8358);
or U8500 (N_8500,N_8330,N_8263);
nor U8501 (N_8501,N_8397,N_8207);
nand U8502 (N_8502,N_8333,N_8392);
xnor U8503 (N_8503,N_8336,N_8390);
and U8504 (N_8504,N_8245,N_8386);
xnor U8505 (N_8505,N_8332,N_8370);
nand U8506 (N_8506,N_8354,N_8394);
and U8507 (N_8507,N_8305,N_8209);
and U8508 (N_8508,N_8276,N_8277);
or U8509 (N_8509,N_8398,N_8213);
nand U8510 (N_8510,N_8314,N_8324);
xnor U8511 (N_8511,N_8305,N_8398);
or U8512 (N_8512,N_8262,N_8390);
nor U8513 (N_8513,N_8390,N_8236);
and U8514 (N_8514,N_8317,N_8310);
and U8515 (N_8515,N_8297,N_8379);
nor U8516 (N_8516,N_8219,N_8216);
nand U8517 (N_8517,N_8389,N_8298);
and U8518 (N_8518,N_8212,N_8358);
and U8519 (N_8519,N_8336,N_8298);
nand U8520 (N_8520,N_8371,N_8312);
and U8521 (N_8521,N_8303,N_8237);
nand U8522 (N_8522,N_8206,N_8300);
nand U8523 (N_8523,N_8330,N_8365);
nand U8524 (N_8524,N_8201,N_8221);
or U8525 (N_8525,N_8385,N_8325);
xnor U8526 (N_8526,N_8224,N_8209);
or U8527 (N_8527,N_8247,N_8331);
nor U8528 (N_8528,N_8247,N_8207);
or U8529 (N_8529,N_8389,N_8364);
nand U8530 (N_8530,N_8389,N_8371);
nand U8531 (N_8531,N_8396,N_8205);
or U8532 (N_8532,N_8282,N_8367);
nand U8533 (N_8533,N_8266,N_8346);
and U8534 (N_8534,N_8222,N_8357);
or U8535 (N_8535,N_8217,N_8246);
and U8536 (N_8536,N_8318,N_8319);
xnor U8537 (N_8537,N_8222,N_8263);
and U8538 (N_8538,N_8208,N_8388);
and U8539 (N_8539,N_8269,N_8288);
or U8540 (N_8540,N_8250,N_8312);
xnor U8541 (N_8541,N_8374,N_8276);
nor U8542 (N_8542,N_8213,N_8378);
xor U8543 (N_8543,N_8247,N_8254);
xnor U8544 (N_8544,N_8387,N_8240);
or U8545 (N_8545,N_8243,N_8239);
or U8546 (N_8546,N_8354,N_8231);
xnor U8547 (N_8547,N_8236,N_8254);
nand U8548 (N_8548,N_8382,N_8216);
and U8549 (N_8549,N_8328,N_8257);
or U8550 (N_8550,N_8326,N_8254);
and U8551 (N_8551,N_8392,N_8291);
nor U8552 (N_8552,N_8220,N_8237);
xnor U8553 (N_8553,N_8237,N_8233);
nor U8554 (N_8554,N_8358,N_8284);
or U8555 (N_8555,N_8324,N_8333);
nor U8556 (N_8556,N_8265,N_8295);
nand U8557 (N_8557,N_8316,N_8216);
nand U8558 (N_8558,N_8299,N_8378);
or U8559 (N_8559,N_8236,N_8320);
nand U8560 (N_8560,N_8344,N_8272);
or U8561 (N_8561,N_8318,N_8269);
or U8562 (N_8562,N_8239,N_8308);
nand U8563 (N_8563,N_8364,N_8355);
and U8564 (N_8564,N_8332,N_8380);
xor U8565 (N_8565,N_8226,N_8221);
nand U8566 (N_8566,N_8266,N_8222);
nor U8567 (N_8567,N_8307,N_8210);
or U8568 (N_8568,N_8282,N_8392);
xnor U8569 (N_8569,N_8204,N_8336);
or U8570 (N_8570,N_8315,N_8360);
nor U8571 (N_8571,N_8207,N_8224);
or U8572 (N_8572,N_8315,N_8303);
xnor U8573 (N_8573,N_8380,N_8212);
xnor U8574 (N_8574,N_8367,N_8378);
nand U8575 (N_8575,N_8235,N_8202);
or U8576 (N_8576,N_8257,N_8380);
and U8577 (N_8577,N_8232,N_8399);
and U8578 (N_8578,N_8225,N_8368);
nand U8579 (N_8579,N_8290,N_8395);
nor U8580 (N_8580,N_8269,N_8385);
nor U8581 (N_8581,N_8372,N_8339);
xor U8582 (N_8582,N_8262,N_8364);
or U8583 (N_8583,N_8349,N_8324);
and U8584 (N_8584,N_8257,N_8385);
or U8585 (N_8585,N_8315,N_8366);
xor U8586 (N_8586,N_8282,N_8358);
xnor U8587 (N_8587,N_8360,N_8237);
nor U8588 (N_8588,N_8321,N_8214);
nand U8589 (N_8589,N_8300,N_8288);
nor U8590 (N_8590,N_8275,N_8228);
nor U8591 (N_8591,N_8259,N_8272);
nand U8592 (N_8592,N_8244,N_8296);
and U8593 (N_8593,N_8308,N_8211);
nand U8594 (N_8594,N_8336,N_8235);
and U8595 (N_8595,N_8315,N_8350);
nand U8596 (N_8596,N_8355,N_8312);
nor U8597 (N_8597,N_8259,N_8398);
nand U8598 (N_8598,N_8378,N_8370);
xor U8599 (N_8599,N_8344,N_8324);
xor U8600 (N_8600,N_8449,N_8537);
xor U8601 (N_8601,N_8563,N_8544);
nand U8602 (N_8602,N_8463,N_8474);
or U8603 (N_8603,N_8491,N_8472);
nor U8604 (N_8604,N_8598,N_8405);
nand U8605 (N_8605,N_8541,N_8403);
and U8606 (N_8606,N_8477,N_8443);
nand U8607 (N_8607,N_8485,N_8513);
or U8608 (N_8608,N_8462,N_8557);
xnor U8609 (N_8609,N_8448,N_8464);
xor U8610 (N_8610,N_8421,N_8533);
xnor U8611 (N_8611,N_8407,N_8585);
nor U8612 (N_8612,N_8436,N_8590);
nor U8613 (N_8613,N_8439,N_8578);
nand U8614 (N_8614,N_8527,N_8434);
nor U8615 (N_8615,N_8592,N_8424);
nand U8616 (N_8616,N_8499,N_8521);
and U8617 (N_8617,N_8414,N_8471);
xnor U8618 (N_8618,N_8586,N_8510);
nor U8619 (N_8619,N_8495,N_8481);
and U8620 (N_8620,N_8401,N_8546);
nor U8621 (N_8621,N_8504,N_8498);
nor U8622 (N_8622,N_8516,N_8540);
and U8623 (N_8623,N_8451,N_8593);
and U8624 (N_8624,N_8589,N_8534);
or U8625 (N_8625,N_8475,N_8554);
nor U8626 (N_8626,N_8415,N_8497);
and U8627 (N_8627,N_8579,N_8509);
nand U8628 (N_8628,N_8572,N_8530);
or U8629 (N_8629,N_8418,N_8599);
and U8630 (N_8630,N_8549,N_8465);
and U8631 (N_8631,N_8416,N_8483);
nor U8632 (N_8632,N_8412,N_8550);
xnor U8633 (N_8633,N_8486,N_8553);
xor U8634 (N_8634,N_8571,N_8506);
nand U8635 (N_8635,N_8512,N_8558);
and U8636 (N_8636,N_8548,N_8400);
xnor U8637 (N_8637,N_8425,N_8520);
xor U8638 (N_8638,N_8411,N_8461);
or U8639 (N_8639,N_8567,N_8577);
nor U8640 (N_8640,N_8404,N_8431);
nor U8641 (N_8641,N_8423,N_8442);
nor U8642 (N_8642,N_8435,N_8438);
and U8643 (N_8643,N_8591,N_8417);
xnor U8644 (N_8644,N_8524,N_8496);
xnor U8645 (N_8645,N_8445,N_8538);
and U8646 (N_8646,N_8479,N_8539);
and U8647 (N_8647,N_8576,N_8455);
or U8648 (N_8648,N_8525,N_8594);
nor U8649 (N_8649,N_8532,N_8597);
nor U8650 (N_8650,N_8409,N_8573);
xor U8651 (N_8651,N_8467,N_8511);
nor U8652 (N_8652,N_8427,N_8518);
and U8653 (N_8653,N_8528,N_8494);
and U8654 (N_8654,N_8587,N_8480);
or U8655 (N_8655,N_8582,N_8531);
nand U8656 (N_8656,N_8559,N_8447);
and U8657 (N_8657,N_8476,N_8562);
xor U8658 (N_8658,N_8551,N_8454);
xnor U8659 (N_8659,N_8568,N_8545);
xor U8660 (N_8660,N_8478,N_8526);
nand U8661 (N_8661,N_8515,N_8453);
nand U8662 (N_8662,N_8542,N_8505);
and U8663 (N_8663,N_8446,N_8569);
xor U8664 (N_8664,N_8580,N_8536);
and U8665 (N_8665,N_8493,N_8519);
and U8666 (N_8666,N_8535,N_8584);
xnor U8667 (N_8667,N_8419,N_8420);
xor U8668 (N_8668,N_8469,N_8556);
xnor U8669 (N_8669,N_8408,N_8444);
or U8670 (N_8670,N_8508,N_8575);
xnor U8671 (N_8671,N_8432,N_8564);
nand U8672 (N_8672,N_8422,N_8523);
and U8673 (N_8673,N_8503,N_8402);
and U8674 (N_8674,N_8517,N_8566);
nand U8675 (N_8675,N_8560,N_8514);
nand U8676 (N_8676,N_8547,N_8596);
xor U8677 (N_8677,N_8492,N_8410);
and U8678 (N_8678,N_8489,N_8433);
xor U8679 (N_8679,N_8543,N_8522);
and U8680 (N_8680,N_8430,N_8529);
and U8681 (N_8681,N_8440,N_8502);
or U8682 (N_8682,N_8507,N_8488);
xor U8683 (N_8683,N_8470,N_8460);
nor U8684 (N_8684,N_8450,N_8441);
and U8685 (N_8685,N_8456,N_8482);
and U8686 (N_8686,N_8561,N_8459);
nor U8687 (N_8687,N_8452,N_8487);
xnor U8688 (N_8688,N_8581,N_8552);
or U8689 (N_8689,N_8565,N_8595);
nor U8690 (N_8690,N_8437,N_8466);
xor U8691 (N_8691,N_8473,N_8406);
nand U8692 (N_8692,N_8428,N_8457);
nand U8693 (N_8693,N_8458,N_8426);
or U8694 (N_8694,N_8429,N_8484);
nor U8695 (N_8695,N_8555,N_8413);
or U8696 (N_8696,N_8468,N_8490);
nor U8697 (N_8697,N_8583,N_8570);
and U8698 (N_8698,N_8588,N_8500);
nand U8699 (N_8699,N_8574,N_8501);
or U8700 (N_8700,N_8431,N_8545);
nand U8701 (N_8701,N_8410,N_8547);
or U8702 (N_8702,N_8400,N_8420);
or U8703 (N_8703,N_8576,N_8423);
and U8704 (N_8704,N_8423,N_8544);
nand U8705 (N_8705,N_8566,N_8484);
nand U8706 (N_8706,N_8492,N_8497);
xor U8707 (N_8707,N_8443,N_8560);
nand U8708 (N_8708,N_8405,N_8531);
xnor U8709 (N_8709,N_8518,N_8433);
or U8710 (N_8710,N_8534,N_8462);
or U8711 (N_8711,N_8444,N_8523);
xor U8712 (N_8712,N_8537,N_8574);
or U8713 (N_8713,N_8592,N_8529);
or U8714 (N_8714,N_8527,N_8472);
xnor U8715 (N_8715,N_8409,N_8442);
xnor U8716 (N_8716,N_8568,N_8488);
or U8717 (N_8717,N_8512,N_8514);
nor U8718 (N_8718,N_8558,N_8485);
nand U8719 (N_8719,N_8455,N_8531);
nand U8720 (N_8720,N_8453,N_8444);
and U8721 (N_8721,N_8464,N_8450);
and U8722 (N_8722,N_8550,N_8441);
xor U8723 (N_8723,N_8571,N_8555);
and U8724 (N_8724,N_8448,N_8528);
and U8725 (N_8725,N_8475,N_8543);
nor U8726 (N_8726,N_8438,N_8573);
nor U8727 (N_8727,N_8536,N_8526);
nand U8728 (N_8728,N_8559,N_8595);
nand U8729 (N_8729,N_8592,N_8508);
xnor U8730 (N_8730,N_8405,N_8513);
xnor U8731 (N_8731,N_8583,N_8415);
or U8732 (N_8732,N_8423,N_8477);
nand U8733 (N_8733,N_8599,N_8434);
xnor U8734 (N_8734,N_8520,N_8490);
xnor U8735 (N_8735,N_8451,N_8556);
or U8736 (N_8736,N_8554,N_8529);
and U8737 (N_8737,N_8415,N_8596);
nor U8738 (N_8738,N_8404,N_8552);
or U8739 (N_8739,N_8484,N_8446);
or U8740 (N_8740,N_8442,N_8507);
xnor U8741 (N_8741,N_8558,N_8591);
or U8742 (N_8742,N_8571,N_8589);
nand U8743 (N_8743,N_8470,N_8502);
or U8744 (N_8744,N_8569,N_8597);
nand U8745 (N_8745,N_8409,N_8580);
nor U8746 (N_8746,N_8483,N_8485);
and U8747 (N_8747,N_8470,N_8464);
and U8748 (N_8748,N_8514,N_8447);
or U8749 (N_8749,N_8597,N_8552);
or U8750 (N_8750,N_8546,N_8553);
xnor U8751 (N_8751,N_8464,N_8574);
and U8752 (N_8752,N_8556,N_8426);
xnor U8753 (N_8753,N_8501,N_8497);
or U8754 (N_8754,N_8527,N_8470);
nand U8755 (N_8755,N_8425,N_8426);
and U8756 (N_8756,N_8438,N_8491);
xnor U8757 (N_8757,N_8563,N_8472);
xnor U8758 (N_8758,N_8489,N_8421);
nor U8759 (N_8759,N_8450,N_8589);
nor U8760 (N_8760,N_8457,N_8449);
and U8761 (N_8761,N_8557,N_8532);
nor U8762 (N_8762,N_8533,N_8490);
nor U8763 (N_8763,N_8446,N_8429);
nand U8764 (N_8764,N_8401,N_8536);
nor U8765 (N_8765,N_8426,N_8519);
nand U8766 (N_8766,N_8586,N_8402);
and U8767 (N_8767,N_8467,N_8466);
and U8768 (N_8768,N_8415,N_8595);
xor U8769 (N_8769,N_8403,N_8525);
xor U8770 (N_8770,N_8546,N_8460);
nand U8771 (N_8771,N_8575,N_8490);
or U8772 (N_8772,N_8425,N_8472);
and U8773 (N_8773,N_8445,N_8454);
nor U8774 (N_8774,N_8459,N_8487);
xnor U8775 (N_8775,N_8519,N_8459);
or U8776 (N_8776,N_8433,N_8579);
xor U8777 (N_8777,N_8482,N_8426);
nand U8778 (N_8778,N_8567,N_8488);
nor U8779 (N_8779,N_8468,N_8578);
or U8780 (N_8780,N_8439,N_8553);
and U8781 (N_8781,N_8420,N_8414);
and U8782 (N_8782,N_8510,N_8487);
and U8783 (N_8783,N_8567,N_8445);
and U8784 (N_8784,N_8417,N_8463);
nor U8785 (N_8785,N_8463,N_8519);
nor U8786 (N_8786,N_8416,N_8584);
nand U8787 (N_8787,N_8495,N_8457);
xor U8788 (N_8788,N_8480,N_8463);
nand U8789 (N_8789,N_8550,N_8596);
nor U8790 (N_8790,N_8567,N_8452);
or U8791 (N_8791,N_8405,N_8484);
or U8792 (N_8792,N_8597,N_8484);
and U8793 (N_8793,N_8523,N_8476);
nor U8794 (N_8794,N_8563,N_8570);
nor U8795 (N_8795,N_8465,N_8408);
or U8796 (N_8796,N_8502,N_8507);
and U8797 (N_8797,N_8480,N_8482);
and U8798 (N_8798,N_8527,N_8496);
or U8799 (N_8799,N_8502,N_8416);
xor U8800 (N_8800,N_8729,N_8724);
or U8801 (N_8801,N_8646,N_8761);
nor U8802 (N_8802,N_8770,N_8749);
and U8803 (N_8803,N_8658,N_8720);
and U8804 (N_8804,N_8702,N_8689);
nand U8805 (N_8805,N_8779,N_8601);
or U8806 (N_8806,N_8675,N_8691);
and U8807 (N_8807,N_8630,N_8678);
nand U8808 (N_8808,N_8640,N_8748);
xor U8809 (N_8809,N_8672,N_8754);
or U8810 (N_8810,N_8617,N_8606);
or U8811 (N_8811,N_8653,N_8621);
xnor U8812 (N_8812,N_8768,N_8767);
and U8813 (N_8813,N_8627,N_8792);
nand U8814 (N_8814,N_8622,N_8741);
nand U8815 (N_8815,N_8695,N_8626);
nor U8816 (N_8816,N_8789,N_8759);
xor U8817 (N_8817,N_8777,N_8743);
xor U8818 (N_8818,N_8730,N_8760);
or U8819 (N_8819,N_8731,N_8620);
and U8820 (N_8820,N_8733,N_8603);
nand U8821 (N_8821,N_8788,N_8758);
nor U8822 (N_8822,N_8610,N_8794);
and U8823 (N_8823,N_8696,N_8736);
nand U8824 (N_8824,N_8655,N_8719);
nor U8825 (N_8825,N_8667,N_8780);
xor U8826 (N_8826,N_8709,N_8628);
or U8827 (N_8827,N_8739,N_8745);
and U8828 (N_8828,N_8668,N_8652);
xor U8829 (N_8829,N_8661,N_8649);
nor U8830 (N_8830,N_8732,N_8635);
nor U8831 (N_8831,N_8756,N_8664);
or U8832 (N_8832,N_8639,N_8642);
nor U8833 (N_8833,N_8692,N_8656);
nor U8834 (N_8834,N_8685,N_8778);
or U8835 (N_8835,N_8644,N_8711);
or U8836 (N_8836,N_8795,N_8633);
or U8837 (N_8837,N_8604,N_8747);
nand U8838 (N_8838,N_8742,N_8632);
xor U8839 (N_8839,N_8625,N_8699);
nor U8840 (N_8840,N_8682,N_8796);
xor U8841 (N_8841,N_8684,N_8722);
xnor U8842 (N_8842,N_8766,N_8707);
xor U8843 (N_8843,N_8671,N_8654);
and U8844 (N_8844,N_8703,N_8791);
xnor U8845 (N_8845,N_8771,N_8700);
or U8846 (N_8846,N_8614,N_8681);
nor U8847 (N_8847,N_8624,N_8753);
and U8848 (N_8848,N_8773,N_8734);
xnor U8849 (N_8849,N_8718,N_8677);
nand U8850 (N_8850,N_8615,N_8697);
or U8851 (N_8851,N_8715,N_8650);
or U8852 (N_8852,N_8755,N_8662);
xor U8853 (N_8853,N_8686,N_8623);
nor U8854 (N_8854,N_8751,N_8714);
or U8855 (N_8855,N_8793,N_8645);
nor U8856 (N_8856,N_8781,N_8643);
nor U8857 (N_8857,N_8612,N_8647);
and U8858 (N_8858,N_8680,N_8631);
or U8859 (N_8859,N_8634,N_8784);
nor U8860 (N_8860,N_8694,N_8663);
nand U8861 (N_8861,N_8616,N_8775);
or U8862 (N_8862,N_8673,N_8776);
xor U8863 (N_8863,N_8674,N_8648);
nor U8864 (N_8864,N_8727,N_8746);
xor U8865 (N_8865,N_8602,N_8688);
nand U8866 (N_8866,N_8701,N_8782);
and U8867 (N_8867,N_8659,N_8798);
and U8868 (N_8868,N_8799,N_8763);
nor U8869 (N_8869,N_8687,N_8619);
nand U8870 (N_8870,N_8641,N_8750);
nor U8871 (N_8871,N_8683,N_8726);
nand U8872 (N_8872,N_8636,N_8744);
and U8873 (N_8873,N_8721,N_8786);
and U8874 (N_8874,N_8651,N_8723);
nor U8875 (N_8875,N_8608,N_8629);
or U8876 (N_8876,N_8710,N_8607);
nor U8877 (N_8877,N_8660,N_8708);
nor U8878 (N_8878,N_8679,N_8609);
nor U8879 (N_8879,N_8665,N_8790);
xor U8880 (N_8880,N_8787,N_8728);
and U8881 (N_8881,N_8638,N_8600);
xnor U8882 (N_8882,N_8605,N_8785);
xnor U8883 (N_8883,N_8712,N_8690);
nor U8884 (N_8884,N_8657,N_8698);
nand U8885 (N_8885,N_8693,N_8737);
nand U8886 (N_8886,N_8705,N_8725);
and U8887 (N_8887,N_8713,N_8797);
nand U8888 (N_8888,N_8740,N_8669);
nor U8889 (N_8889,N_8611,N_8676);
nor U8890 (N_8890,N_8783,N_8765);
and U8891 (N_8891,N_8704,N_8772);
nand U8892 (N_8892,N_8774,N_8716);
and U8893 (N_8893,N_8618,N_8670);
or U8894 (N_8894,N_8738,N_8717);
xnor U8895 (N_8895,N_8769,N_8752);
xnor U8896 (N_8896,N_8706,N_8666);
nor U8897 (N_8897,N_8637,N_8764);
and U8898 (N_8898,N_8762,N_8613);
nand U8899 (N_8899,N_8757,N_8735);
nand U8900 (N_8900,N_8655,N_8637);
nor U8901 (N_8901,N_8742,N_8703);
or U8902 (N_8902,N_8692,N_8691);
or U8903 (N_8903,N_8732,N_8698);
or U8904 (N_8904,N_8751,N_8715);
xnor U8905 (N_8905,N_8679,N_8748);
nor U8906 (N_8906,N_8625,N_8623);
and U8907 (N_8907,N_8758,N_8625);
nand U8908 (N_8908,N_8660,N_8753);
xnor U8909 (N_8909,N_8698,N_8785);
xnor U8910 (N_8910,N_8719,N_8676);
nand U8911 (N_8911,N_8769,N_8764);
xor U8912 (N_8912,N_8619,N_8668);
and U8913 (N_8913,N_8656,N_8716);
and U8914 (N_8914,N_8742,N_8765);
nor U8915 (N_8915,N_8677,N_8728);
nor U8916 (N_8916,N_8674,N_8659);
nand U8917 (N_8917,N_8651,N_8643);
nor U8918 (N_8918,N_8733,N_8786);
nor U8919 (N_8919,N_8787,N_8618);
or U8920 (N_8920,N_8638,N_8679);
nand U8921 (N_8921,N_8753,N_8798);
nor U8922 (N_8922,N_8753,N_8728);
xnor U8923 (N_8923,N_8627,N_8793);
xnor U8924 (N_8924,N_8639,N_8748);
and U8925 (N_8925,N_8618,N_8727);
nand U8926 (N_8926,N_8752,N_8704);
nand U8927 (N_8927,N_8648,N_8739);
nand U8928 (N_8928,N_8772,N_8736);
nand U8929 (N_8929,N_8751,N_8707);
or U8930 (N_8930,N_8717,N_8688);
nand U8931 (N_8931,N_8623,N_8794);
and U8932 (N_8932,N_8661,N_8721);
xor U8933 (N_8933,N_8729,N_8799);
and U8934 (N_8934,N_8613,N_8726);
and U8935 (N_8935,N_8695,N_8718);
and U8936 (N_8936,N_8784,N_8653);
xor U8937 (N_8937,N_8635,N_8625);
and U8938 (N_8938,N_8645,N_8617);
xor U8939 (N_8939,N_8682,N_8726);
or U8940 (N_8940,N_8796,N_8633);
xnor U8941 (N_8941,N_8677,N_8768);
and U8942 (N_8942,N_8785,N_8760);
or U8943 (N_8943,N_8630,N_8600);
nor U8944 (N_8944,N_8673,N_8653);
and U8945 (N_8945,N_8676,N_8644);
nor U8946 (N_8946,N_8711,N_8681);
nand U8947 (N_8947,N_8658,N_8741);
or U8948 (N_8948,N_8722,N_8798);
and U8949 (N_8949,N_8698,N_8797);
or U8950 (N_8950,N_8753,N_8667);
or U8951 (N_8951,N_8651,N_8766);
xor U8952 (N_8952,N_8643,N_8735);
nand U8953 (N_8953,N_8710,N_8646);
nand U8954 (N_8954,N_8616,N_8714);
and U8955 (N_8955,N_8616,N_8622);
xnor U8956 (N_8956,N_8720,N_8796);
xor U8957 (N_8957,N_8682,N_8714);
or U8958 (N_8958,N_8659,N_8792);
xor U8959 (N_8959,N_8637,N_8716);
and U8960 (N_8960,N_8777,N_8660);
nor U8961 (N_8961,N_8656,N_8686);
or U8962 (N_8962,N_8627,N_8619);
or U8963 (N_8963,N_8617,N_8673);
or U8964 (N_8964,N_8737,N_8786);
nor U8965 (N_8965,N_8729,N_8707);
or U8966 (N_8966,N_8611,N_8720);
and U8967 (N_8967,N_8741,N_8797);
or U8968 (N_8968,N_8689,N_8746);
and U8969 (N_8969,N_8731,N_8756);
and U8970 (N_8970,N_8622,N_8723);
nand U8971 (N_8971,N_8749,N_8736);
xor U8972 (N_8972,N_8706,N_8764);
or U8973 (N_8973,N_8616,N_8617);
and U8974 (N_8974,N_8675,N_8771);
nand U8975 (N_8975,N_8780,N_8675);
xor U8976 (N_8976,N_8651,N_8797);
and U8977 (N_8977,N_8627,N_8701);
xnor U8978 (N_8978,N_8628,N_8781);
nor U8979 (N_8979,N_8734,N_8702);
and U8980 (N_8980,N_8700,N_8781);
nand U8981 (N_8981,N_8791,N_8748);
nor U8982 (N_8982,N_8729,N_8634);
nand U8983 (N_8983,N_8745,N_8614);
nand U8984 (N_8984,N_8797,N_8610);
nand U8985 (N_8985,N_8675,N_8781);
and U8986 (N_8986,N_8778,N_8656);
and U8987 (N_8987,N_8710,N_8724);
nand U8988 (N_8988,N_8736,N_8780);
xnor U8989 (N_8989,N_8621,N_8770);
or U8990 (N_8990,N_8771,N_8779);
nor U8991 (N_8991,N_8702,N_8660);
xor U8992 (N_8992,N_8739,N_8761);
nand U8993 (N_8993,N_8620,N_8652);
xnor U8994 (N_8994,N_8785,N_8771);
nand U8995 (N_8995,N_8769,N_8794);
or U8996 (N_8996,N_8692,N_8600);
and U8997 (N_8997,N_8626,N_8672);
xor U8998 (N_8998,N_8799,N_8792);
or U8999 (N_8999,N_8786,N_8634);
nor U9000 (N_9000,N_8847,N_8921);
nor U9001 (N_9001,N_8848,N_8970);
xnor U9002 (N_9002,N_8932,N_8808);
nand U9003 (N_9003,N_8923,N_8976);
and U9004 (N_9004,N_8925,N_8850);
nand U9005 (N_9005,N_8889,N_8826);
nor U9006 (N_9006,N_8959,N_8904);
nor U9007 (N_9007,N_8806,N_8844);
nor U9008 (N_9008,N_8836,N_8967);
nor U9009 (N_9009,N_8802,N_8998);
and U9010 (N_9010,N_8989,N_8810);
and U9011 (N_9011,N_8897,N_8930);
nor U9012 (N_9012,N_8949,N_8852);
xnor U9013 (N_9013,N_8879,N_8895);
or U9014 (N_9014,N_8829,N_8974);
or U9015 (N_9015,N_8940,N_8917);
or U9016 (N_9016,N_8894,N_8872);
xnor U9017 (N_9017,N_8864,N_8855);
xor U9018 (N_9018,N_8824,N_8909);
nor U9019 (N_9019,N_8863,N_8983);
nor U9020 (N_9020,N_8945,N_8985);
and U9021 (N_9021,N_8832,N_8920);
and U9022 (N_9022,N_8843,N_8980);
or U9023 (N_9023,N_8933,N_8992);
xor U9024 (N_9024,N_8885,N_8803);
nor U9025 (N_9025,N_8886,N_8859);
nand U9026 (N_9026,N_8825,N_8997);
nand U9027 (N_9027,N_8971,N_8951);
nor U9028 (N_9028,N_8965,N_8880);
and U9029 (N_9029,N_8961,N_8870);
and U9030 (N_9030,N_8849,N_8981);
or U9031 (N_9031,N_8883,N_8882);
and U9032 (N_9032,N_8984,N_8966);
or U9033 (N_9033,N_8939,N_8868);
and U9034 (N_9034,N_8922,N_8827);
nand U9035 (N_9035,N_8861,N_8887);
or U9036 (N_9036,N_8817,N_8948);
nor U9037 (N_9037,N_8898,N_8874);
xnor U9038 (N_9038,N_8986,N_8916);
and U9039 (N_9039,N_8968,N_8867);
or U9040 (N_9040,N_8934,N_8805);
nand U9041 (N_9041,N_8907,N_8891);
nand U9042 (N_9042,N_8900,N_8800);
nand U9043 (N_9043,N_8857,N_8801);
and U9044 (N_9044,N_8823,N_8990);
nor U9045 (N_9045,N_8941,N_8964);
and U9046 (N_9046,N_8838,N_8860);
nand U9047 (N_9047,N_8969,N_8875);
nand U9048 (N_9048,N_8912,N_8944);
and U9049 (N_9049,N_8809,N_8873);
xnor U9050 (N_9050,N_8896,N_8804);
xnor U9051 (N_9051,N_8999,N_8987);
nor U9052 (N_9052,N_8956,N_8845);
xnor U9053 (N_9053,N_8819,N_8881);
or U9054 (N_9054,N_8908,N_8988);
nor U9055 (N_9055,N_8869,N_8830);
nor U9056 (N_9056,N_8834,N_8991);
nor U9057 (N_9057,N_8935,N_8821);
nor U9058 (N_9058,N_8822,N_8831);
nor U9059 (N_9059,N_8856,N_8947);
and U9060 (N_9060,N_8840,N_8812);
or U9061 (N_9061,N_8913,N_8833);
and U9062 (N_9062,N_8929,N_8931);
xnor U9063 (N_9063,N_8910,N_8924);
xnor U9064 (N_9064,N_8942,N_8818);
nor U9065 (N_9065,N_8858,N_8938);
nand U9066 (N_9066,N_8807,N_8811);
xnor U9067 (N_9067,N_8978,N_8884);
xor U9068 (N_9068,N_8975,N_8973);
xnor U9069 (N_9069,N_8950,N_8958);
and U9070 (N_9070,N_8994,N_8837);
and U9071 (N_9071,N_8946,N_8816);
nand U9072 (N_9072,N_8926,N_8955);
or U9073 (N_9073,N_8936,N_8915);
and U9074 (N_9074,N_8846,N_8993);
nor U9075 (N_9075,N_8892,N_8841);
xor U9076 (N_9076,N_8851,N_8919);
xor U9077 (N_9077,N_8928,N_8862);
nor U9078 (N_9078,N_8839,N_8962);
nand U9079 (N_9079,N_8871,N_8960);
nand U9080 (N_9080,N_8828,N_8954);
xnor U9081 (N_9081,N_8963,N_8914);
or U9082 (N_9082,N_8905,N_8820);
nor U9083 (N_9083,N_8982,N_8927);
nand U9084 (N_9084,N_8815,N_8901);
nand U9085 (N_9085,N_8996,N_8813);
xor U9086 (N_9086,N_8903,N_8952);
nand U9087 (N_9087,N_8899,N_8814);
xnor U9088 (N_9088,N_8893,N_8906);
nand U9089 (N_9089,N_8877,N_8979);
nand U9090 (N_9090,N_8957,N_8876);
xnor U9091 (N_9091,N_8995,N_8854);
and U9092 (N_9092,N_8842,N_8977);
and U9093 (N_9093,N_8888,N_8918);
nand U9094 (N_9094,N_8902,N_8835);
or U9095 (N_9095,N_8890,N_8853);
or U9096 (N_9096,N_8911,N_8866);
nand U9097 (N_9097,N_8943,N_8953);
xnor U9098 (N_9098,N_8937,N_8865);
xnor U9099 (N_9099,N_8972,N_8878);
nor U9100 (N_9100,N_8873,N_8969);
xnor U9101 (N_9101,N_8971,N_8847);
nor U9102 (N_9102,N_8861,N_8809);
xor U9103 (N_9103,N_8825,N_8871);
and U9104 (N_9104,N_8965,N_8873);
xor U9105 (N_9105,N_8907,N_8839);
nor U9106 (N_9106,N_8989,N_8931);
or U9107 (N_9107,N_8840,N_8938);
or U9108 (N_9108,N_8967,N_8834);
or U9109 (N_9109,N_8998,N_8947);
or U9110 (N_9110,N_8866,N_8848);
xor U9111 (N_9111,N_8900,N_8824);
xnor U9112 (N_9112,N_8907,N_8979);
nor U9113 (N_9113,N_8997,N_8939);
nand U9114 (N_9114,N_8806,N_8903);
nor U9115 (N_9115,N_8875,N_8814);
or U9116 (N_9116,N_8828,N_8845);
nor U9117 (N_9117,N_8909,N_8963);
and U9118 (N_9118,N_8800,N_8995);
or U9119 (N_9119,N_8899,N_8994);
and U9120 (N_9120,N_8871,N_8989);
xnor U9121 (N_9121,N_8880,N_8951);
or U9122 (N_9122,N_8902,N_8842);
xnor U9123 (N_9123,N_8849,N_8967);
xor U9124 (N_9124,N_8955,N_8868);
or U9125 (N_9125,N_8896,N_8803);
or U9126 (N_9126,N_8863,N_8850);
xor U9127 (N_9127,N_8970,N_8836);
nand U9128 (N_9128,N_8915,N_8876);
and U9129 (N_9129,N_8866,N_8925);
xnor U9130 (N_9130,N_8878,N_8969);
xnor U9131 (N_9131,N_8933,N_8813);
and U9132 (N_9132,N_8915,N_8978);
nand U9133 (N_9133,N_8900,N_8870);
nand U9134 (N_9134,N_8899,N_8880);
or U9135 (N_9135,N_8931,N_8993);
or U9136 (N_9136,N_8942,N_8867);
or U9137 (N_9137,N_8972,N_8891);
nor U9138 (N_9138,N_8914,N_8977);
xor U9139 (N_9139,N_8895,N_8863);
xnor U9140 (N_9140,N_8811,N_8900);
nor U9141 (N_9141,N_8865,N_8969);
or U9142 (N_9142,N_8989,N_8968);
nand U9143 (N_9143,N_8977,N_8894);
nand U9144 (N_9144,N_8980,N_8878);
nand U9145 (N_9145,N_8999,N_8821);
xor U9146 (N_9146,N_8873,N_8879);
or U9147 (N_9147,N_8908,N_8812);
or U9148 (N_9148,N_8802,N_8848);
nand U9149 (N_9149,N_8813,N_8984);
nor U9150 (N_9150,N_8996,N_8993);
nor U9151 (N_9151,N_8860,N_8924);
and U9152 (N_9152,N_8945,N_8974);
xor U9153 (N_9153,N_8988,N_8873);
nand U9154 (N_9154,N_8972,N_8966);
xor U9155 (N_9155,N_8950,N_8879);
nor U9156 (N_9156,N_8889,N_8863);
nand U9157 (N_9157,N_8805,N_8801);
and U9158 (N_9158,N_8993,N_8860);
xor U9159 (N_9159,N_8936,N_8979);
nand U9160 (N_9160,N_8870,N_8907);
or U9161 (N_9161,N_8986,N_8891);
xor U9162 (N_9162,N_8895,N_8997);
nand U9163 (N_9163,N_8824,N_8826);
nand U9164 (N_9164,N_8936,N_8954);
or U9165 (N_9165,N_8825,N_8958);
nor U9166 (N_9166,N_8994,N_8855);
xnor U9167 (N_9167,N_8964,N_8874);
xor U9168 (N_9168,N_8902,N_8948);
nand U9169 (N_9169,N_8855,N_8967);
nor U9170 (N_9170,N_8902,N_8843);
nor U9171 (N_9171,N_8915,N_8863);
nand U9172 (N_9172,N_8867,N_8983);
or U9173 (N_9173,N_8955,N_8860);
nor U9174 (N_9174,N_8967,N_8828);
xnor U9175 (N_9175,N_8920,N_8928);
or U9176 (N_9176,N_8985,N_8843);
and U9177 (N_9177,N_8825,N_8992);
or U9178 (N_9178,N_8945,N_8833);
and U9179 (N_9179,N_8910,N_8959);
nand U9180 (N_9180,N_8872,N_8806);
xor U9181 (N_9181,N_8883,N_8816);
nor U9182 (N_9182,N_8848,N_8809);
or U9183 (N_9183,N_8872,N_8936);
or U9184 (N_9184,N_8879,N_8901);
xor U9185 (N_9185,N_8969,N_8908);
xor U9186 (N_9186,N_8986,N_8866);
or U9187 (N_9187,N_8888,N_8892);
nor U9188 (N_9188,N_8822,N_8918);
nand U9189 (N_9189,N_8941,N_8971);
or U9190 (N_9190,N_8816,N_8866);
or U9191 (N_9191,N_8834,N_8880);
nand U9192 (N_9192,N_8883,N_8877);
xor U9193 (N_9193,N_8970,N_8929);
and U9194 (N_9194,N_8959,N_8847);
nor U9195 (N_9195,N_8852,N_8919);
xnor U9196 (N_9196,N_8833,N_8884);
and U9197 (N_9197,N_8848,N_8820);
xnor U9198 (N_9198,N_8880,N_8836);
nor U9199 (N_9199,N_8800,N_8888);
or U9200 (N_9200,N_9111,N_9035);
nor U9201 (N_9201,N_9146,N_9046);
nand U9202 (N_9202,N_9010,N_9175);
or U9203 (N_9203,N_9026,N_9079);
and U9204 (N_9204,N_9130,N_9188);
xnor U9205 (N_9205,N_9198,N_9117);
xnor U9206 (N_9206,N_9122,N_9030);
nor U9207 (N_9207,N_9107,N_9167);
nand U9208 (N_9208,N_9006,N_9015);
and U9209 (N_9209,N_9177,N_9065);
or U9210 (N_9210,N_9016,N_9143);
and U9211 (N_9211,N_9038,N_9158);
and U9212 (N_9212,N_9072,N_9112);
nor U9213 (N_9213,N_9108,N_9005);
or U9214 (N_9214,N_9058,N_9151);
nor U9215 (N_9215,N_9159,N_9189);
nor U9216 (N_9216,N_9050,N_9136);
nand U9217 (N_9217,N_9084,N_9052);
nor U9218 (N_9218,N_9053,N_9094);
or U9219 (N_9219,N_9078,N_9027);
nor U9220 (N_9220,N_9020,N_9007);
nand U9221 (N_9221,N_9069,N_9056);
or U9222 (N_9222,N_9033,N_9067);
nand U9223 (N_9223,N_9100,N_9161);
nor U9224 (N_9224,N_9157,N_9063);
nand U9225 (N_9225,N_9002,N_9199);
and U9226 (N_9226,N_9077,N_9062);
nand U9227 (N_9227,N_9105,N_9021);
and U9228 (N_9228,N_9097,N_9170);
and U9229 (N_9229,N_9031,N_9145);
or U9230 (N_9230,N_9081,N_9193);
xor U9231 (N_9231,N_9116,N_9156);
or U9232 (N_9232,N_9150,N_9133);
xnor U9233 (N_9233,N_9048,N_9068);
nand U9234 (N_9234,N_9032,N_9028);
xnor U9235 (N_9235,N_9114,N_9120);
and U9236 (N_9236,N_9043,N_9162);
nand U9237 (N_9237,N_9142,N_9080);
xor U9238 (N_9238,N_9037,N_9009);
and U9239 (N_9239,N_9057,N_9029);
nor U9240 (N_9240,N_9051,N_9049);
and U9241 (N_9241,N_9082,N_9076);
nor U9242 (N_9242,N_9042,N_9168);
and U9243 (N_9243,N_9060,N_9041);
or U9244 (N_9244,N_9092,N_9164);
xor U9245 (N_9245,N_9018,N_9154);
nand U9246 (N_9246,N_9187,N_9004);
nor U9247 (N_9247,N_9001,N_9073);
or U9248 (N_9248,N_9194,N_9195);
nor U9249 (N_9249,N_9113,N_9163);
xor U9250 (N_9250,N_9135,N_9132);
xnor U9251 (N_9251,N_9129,N_9086);
nor U9252 (N_9252,N_9025,N_9017);
and U9253 (N_9253,N_9186,N_9012);
and U9254 (N_9254,N_9137,N_9153);
nand U9255 (N_9255,N_9166,N_9000);
or U9256 (N_9256,N_9138,N_9176);
or U9257 (N_9257,N_9139,N_9183);
xor U9258 (N_9258,N_9022,N_9179);
and U9259 (N_9259,N_9047,N_9197);
or U9260 (N_9260,N_9074,N_9174);
and U9261 (N_9261,N_9184,N_9045);
xor U9262 (N_9262,N_9095,N_9125);
and U9263 (N_9263,N_9134,N_9091);
or U9264 (N_9264,N_9126,N_9059);
and U9265 (N_9265,N_9109,N_9118);
nor U9266 (N_9266,N_9190,N_9101);
and U9267 (N_9267,N_9149,N_9011);
and U9268 (N_9268,N_9191,N_9013);
nor U9269 (N_9269,N_9093,N_9070);
nand U9270 (N_9270,N_9140,N_9155);
nor U9271 (N_9271,N_9128,N_9099);
nand U9272 (N_9272,N_9054,N_9061);
nor U9273 (N_9273,N_9055,N_9173);
xnor U9274 (N_9274,N_9127,N_9121);
nor U9275 (N_9275,N_9181,N_9090);
nand U9276 (N_9276,N_9180,N_9123);
xor U9277 (N_9277,N_9171,N_9066);
and U9278 (N_9278,N_9178,N_9110);
or U9279 (N_9279,N_9087,N_9044);
xor U9280 (N_9280,N_9003,N_9124);
nand U9281 (N_9281,N_9008,N_9071);
xor U9282 (N_9282,N_9147,N_9064);
nand U9283 (N_9283,N_9160,N_9075);
nor U9284 (N_9284,N_9119,N_9115);
or U9285 (N_9285,N_9019,N_9096);
or U9286 (N_9286,N_9040,N_9098);
nand U9287 (N_9287,N_9172,N_9034);
or U9288 (N_9288,N_9104,N_9036);
or U9289 (N_9289,N_9152,N_9106);
and U9290 (N_9290,N_9085,N_9182);
or U9291 (N_9291,N_9089,N_9102);
xnor U9292 (N_9292,N_9185,N_9144);
or U9293 (N_9293,N_9141,N_9148);
nor U9294 (N_9294,N_9131,N_9014);
xnor U9295 (N_9295,N_9023,N_9192);
nand U9296 (N_9296,N_9039,N_9165);
nand U9297 (N_9297,N_9103,N_9083);
or U9298 (N_9298,N_9196,N_9088);
or U9299 (N_9299,N_9169,N_9024);
and U9300 (N_9300,N_9138,N_9154);
nor U9301 (N_9301,N_9129,N_9182);
xnor U9302 (N_9302,N_9154,N_9056);
and U9303 (N_9303,N_9028,N_9163);
xor U9304 (N_9304,N_9161,N_9096);
or U9305 (N_9305,N_9130,N_9196);
xnor U9306 (N_9306,N_9026,N_9105);
nor U9307 (N_9307,N_9038,N_9118);
and U9308 (N_9308,N_9014,N_9010);
nor U9309 (N_9309,N_9094,N_9161);
xor U9310 (N_9310,N_9005,N_9160);
and U9311 (N_9311,N_9061,N_9069);
or U9312 (N_9312,N_9168,N_9112);
and U9313 (N_9313,N_9169,N_9121);
xor U9314 (N_9314,N_9111,N_9078);
or U9315 (N_9315,N_9116,N_9196);
xnor U9316 (N_9316,N_9190,N_9092);
and U9317 (N_9317,N_9124,N_9182);
or U9318 (N_9318,N_9008,N_9153);
nand U9319 (N_9319,N_9068,N_9023);
nor U9320 (N_9320,N_9175,N_9182);
nor U9321 (N_9321,N_9020,N_9174);
nor U9322 (N_9322,N_9081,N_9036);
and U9323 (N_9323,N_9021,N_9075);
nor U9324 (N_9324,N_9092,N_9172);
xor U9325 (N_9325,N_9140,N_9065);
or U9326 (N_9326,N_9095,N_9058);
nand U9327 (N_9327,N_9103,N_9175);
or U9328 (N_9328,N_9180,N_9041);
nor U9329 (N_9329,N_9072,N_9085);
or U9330 (N_9330,N_9126,N_9096);
xnor U9331 (N_9331,N_9092,N_9184);
nor U9332 (N_9332,N_9061,N_9041);
and U9333 (N_9333,N_9013,N_9059);
xnor U9334 (N_9334,N_9048,N_9045);
and U9335 (N_9335,N_9054,N_9136);
and U9336 (N_9336,N_9036,N_9009);
or U9337 (N_9337,N_9017,N_9164);
xor U9338 (N_9338,N_9099,N_9081);
nand U9339 (N_9339,N_9140,N_9107);
and U9340 (N_9340,N_9118,N_9128);
xor U9341 (N_9341,N_9162,N_9137);
xor U9342 (N_9342,N_9048,N_9158);
and U9343 (N_9343,N_9016,N_9199);
nand U9344 (N_9344,N_9163,N_9148);
and U9345 (N_9345,N_9027,N_9086);
xor U9346 (N_9346,N_9092,N_9020);
nand U9347 (N_9347,N_9078,N_9199);
xor U9348 (N_9348,N_9146,N_9000);
and U9349 (N_9349,N_9173,N_9003);
and U9350 (N_9350,N_9122,N_9079);
nand U9351 (N_9351,N_9082,N_9147);
nor U9352 (N_9352,N_9045,N_9039);
xor U9353 (N_9353,N_9129,N_9022);
and U9354 (N_9354,N_9091,N_9019);
nand U9355 (N_9355,N_9046,N_9029);
or U9356 (N_9356,N_9002,N_9161);
nand U9357 (N_9357,N_9177,N_9027);
and U9358 (N_9358,N_9149,N_9163);
nor U9359 (N_9359,N_9031,N_9158);
and U9360 (N_9360,N_9054,N_9069);
or U9361 (N_9361,N_9178,N_9005);
nor U9362 (N_9362,N_9189,N_9199);
or U9363 (N_9363,N_9005,N_9093);
or U9364 (N_9364,N_9122,N_9049);
and U9365 (N_9365,N_9128,N_9112);
and U9366 (N_9366,N_9049,N_9174);
nor U9367 (N_9367,N_9145,N_9186);
xor U9368 (N_9368,N_9084,N_9102);
or U9369 (N_9369,N_9093,N_9104);
or U9370 (N_9370,N_9104,N_9131);
and U9371 (N_9371,N_9130,N_9028);
or U9372 (N_9372,N_9161,N_9116);
and U9373 (N_9373,N_9066,N_9114);
nor U9374 (N_9374,N_9090,N_9131);
and U9375 (N_9375,N_9130,N_9119);
nor U9376 (N_9376,N_9037,N_9101);
nand U9377 (N_9377,N_9183,N_9135);
and U9378 (N_9378,N_9130,N_9070);
xor U9379 (N_9379,N_9096,N_9129);
xnor U9380 (N_9380,N_9067,N_9117);
xor U9381 (N_9381,N_9161,N_9049);
xnor U9382 (N_9382,N_9006,N_9152);
and U9383 (N_9383,N_9029,N_9189);
nand U9384 (N_9384,N_9091,N_9008);
nand U9385 (N_9385,N_9026,N_9140);
or U9386 (N_9386,N_9178,N_9025);
nor U9387 (N_9387,N_9045,N_9142);
nor U9388 (N_9388,N_9077,N_9130);
nand U9389 (N_9389,N_9100,N_9088);
xor U9390 (N_9390,N_9038,N_9101);
and U9391 (N_9391,N_9048,N_9059);
nor U9392 (N_9392,N_9049,N_9139);
and U9393 (N_9393,N_9062,N_9149);
nor U9394 (N_9394,N_9053,N_9114);
and U9395 (N_9395,N_9143,N_9051);
nand U9396 (N_9396,N_9128,N_9125);
nand U9397 (N_9397,N_9180,N_9174);
xor U9398 (N_9398,N_9118,N_9040);
xor U9399 (N_9399,N_9066,N_9194);
or U9400 (N_9400,N_9285,N_9304);
or U9401 (N_9401,N_9308,N_9368);
or U9402 (N_9402,N_9386,N_9217);
or U9403 (N_9403,N_9320,N_9378);
nor U9404 (N_9404,N_9249,N_9295);
or U9405 (N_9405,N_9351,N_9273);
xor U9406 (N_9406,N_9233,N_9352);
nand U9407 (N_9407,N_9325,N_9251);
nor U9408 (N_9408,N_9252,N_9293);
and U9409 (N_9409,N_9312,N_9228);
xnor U9410 (N_9410,N_9306,N_9318);
nand U9411 (N_9411,N_9324,N_9388);
or U9412 (N_9412,N_9399,N_9329);
and U9413 (N_9413,N_9341,N_9392);
and U9414 (N_9414,N_9391,N_9206);
xnor U9415 (N_9415,N_9362,N_9340);
or U9416 (N_9416,N_9245,N_9365);
xor U9417 (N_9417,N_9343,N_9334);
and U9418 (N_9418,N_9246,N_9240);
or U9419 (N_9419,N_9395,N_9214);
or U9420 (N_9420,N_9313,N_9323);
nand U9421 (N_9421,N_9357,N_9204);
xor U9422 (N_9422,N_9381,N_9363);
nand U9423 (N_9423,N_9230,N_9372);
xor U9424 (N_9424,N_9254,N_9268);
nand U9425 (N_9425,N_9266,N_9307);
and U9426 (N_9426,N_9263,N_9319);
and U9427 (N_9427,N_9342,N_9379);
nor U9428 (N_9428,N_9213,N_9278);
nand U9429 (N_9429,N_9385,N_9299);
nand U9430 (N_9430,N_9262,N_9396);
nand U9431 (N_9431,N_9229,N_9258);
and U9432 (N_9432,N_9239,N_9294);
nor U9433 (N_9433,N_9282,N_9305);
or U9434 (N_9434,N_9302,N_9301);
or U9435 (N_9435,N_9348,N_9375);
xor U9436 (N_9436,N_9234,N_9353);
xnor U9437 (N_9437,N_9280,N_9328);
or U9438 (N_9438,N_9330,N_9347);
and U9439 (N_9439,N_9267,N_9298);
nor U9440 (N_9440,N_9215,N_9284);
nand U9441 (N_9441,N_9290,N_9311);
nor U9442 (N_9442,N_9287,N_9384);
or U9443 (N_9443,N_9255,N_9270);
nor U9444 (N_9444,N_9200,N_9373);
and U9445 (N_9445,N_9380,N_9296);
xnor U9446 (N_9446,N_9383,N_9345);
nand U9447 (N_9447,N_9338,N_9344);
nand U9448 (N_9448,N_9390,N_9201);
xnor U9449 (N_9449,N_9369,N_9218);
or U9450 (N_9450,N_9377,N_9212);
or U9451 (N_9451,N_9269,N_9370);
nand U9452 (N_9452,N_9309,N_9253);
xnor U9453 (N_9453,N_9297,N_9326);
nand U9454 (N_9454,N_9300,N_9259);
or U9455 (N_9455,N_9367,N_9393);
nand U9456 (N_9456,N_9281,N_9241);
nand U9457 (N_9457,N_9376,N_9317);
nor U9458 (N_9458,N_9337,N_9339);
nor U9459 (N_9459,N_9315,N_9274);
nor U9460 (N_9460,N_9216,N_9226);
and U9461 (N_9461,N_9332,N_9333);
xnor U9462 (N_9462,N_9288,N_9321);
xnor U9463 (N_9463,N_9350,N_9277);
nor U9464 (N_9464,N_9220,N_9237);
or U9465 (N_9465,N_9310,N_9243);
and U9466 (N_9466,N_9371,N_9223);
or U9467 (N_9467,N_9208,N_9219);
xor U9468 (N_9468,N_9221,N_9257);
or U9469 (N_9469,N_9303,N_9236);
and U9470 (N_9470,N_9261,N_9210);
xor U9471 (N_9471,N_9366,N_9349);
or U9472 (N_9472,N_9209,N_9265);
and U9473 (N_9473,N_9331,N_9283);
nand U9474 (N_9474,N_9361,N_9389);
or U9475 (N_9475,N_9286,N_9256);
nor U9476 (N_9476,N_9211,N_9356);
xor U9477 (N_9477,N_9360,N_9275);
xnor U9478 (N_9478,N_9222,N_9358);
or U9479 (N_9479,N_9394,N_9354);
nand U9480 (N_9480,N_9387,N_9289);
or U9481 (N_9481,N_9398,N_9397);
nor U9482 (N_9482,N_9248,N_9202);
or U9483 (N_9483,N_9374,N_9272);
or U9484 (N_9484,N_9292,N_9224);
xnor U9485 (N_9485,N_9355,N_9244);
xor U9486 (N_9486,N_9247,N_9364);
nand U9487 (N_9487,N_9242,N_9382);
nand U9488 (N_9488,N_9316,N_9314);
or U9489 (N_9489,N_9276,N_9225);
xor U9490 (N_9490,N_9232,N_9336);
or U9491 (N_9491,N_9327,N_9279);
and U9492 (N_9492,N_9322,N_9205);
and U9493 (N_9493,N_9203,N_9207);
or U9494 (N_9494,N_9264,N_9250);
or U9495 (N_9495,N_9235,N_9231);
nand U9496 (N_9496,N_9271,N_9260);
and U9497 (N_9497,N_9291,N_9359);
nor U9498 (N_9498,N_9238,N_9227);
nand U9499 (N_9499,N_9335,N_9346);
nand U9500 (N_9500,N_9348,N_9374);
nand U9501 (N_9501,N_9343,N_9211);
nor U9502 (N_9502,N_9278,N_9205);
or U9503 (N_9503,N_9204,N_9222);
nand U9504 (N_9504,N_9298,N_9339);
or U9505 (N_9505,N_9291,N_9338);
xor U9506 (N_9506,N_9383,N_9232);
or U9507 (N_9507,N_9227,N_9259);
and U9508 (N_9508,N_9243,N_9370);
nor U9509 (N_9509,N_9295,N_9397);
nor U9510 (N_9510,N_9229,N_9268);
nand U9511 (N_9511,N_9325,N_9300);
and U9512 (N_9512,N_9220,N_9354);
and U9513 (N_9513,N_9248,N_9328);
nor U9514 (N_9514,N_9335,N_9244);
and U9515 (N_9515,N_9330,N_9268);
nand U9516 (N_9516,N_9378,N_9347);
nor U9517 (N_9517,N_9366,N_9388);
or U9518 (N_9518,N_9238,N_9293);
and U9519 (N_9519,N_9296,N_9322);
and U9520 (N_9520,N_9381,N_9340);
or U9521 (N_9521,N_9391,N_9304);
nor U9522 (N_9522,N_9384,N_9282);
or U9523 (N_9523,N_9281,N_9341);
xnor U9524 (N_9524,N_9380,N_9215);
nor U9525 (N_9525,N_9329,N_9245);
nand U9526 (N_9526,N_9240,N_9310);
nand U9527 (N_9527,N_9396,N_9334);
or U9528 (N_9528,N_9336,N_9317);
and U9529 (N_9529,N_9311,N_9223);
nor U9530 (N_9530,N_9383,N_9270);
nor U9531 (N_9531,N_9384,N_9342);
and U9532 (N_9532,N_9206,N_9362);
nor U9533 (N_9533,N_9244,N_9290);
xnor U9534 (N_9534,N_9280,N_9208);
and U9535 (N_9535,N_9364,N_9343);
or U9536 (N_9536,N_9251,N_9383);
nor U9537 (N_9537,N_9272,N_9257);
and U9538 (N_9538,N_9271,N_9303);
and U9539 (N_9539,N_9358,N_9202);
and U9540 (N_9540,N_9214,N_9288);
or U9541 (N_9541,N_9312,N_9382);
nand U9542 (N_9542,N_9251,N_9344);
and U9543 (N_9543,N_9247,N_9381);
nor U9544 (N_9544,N_9210,N_9393);
or U9545 (N_9545,N_9318,N_9280);
xnor U9546 (N_9546,N_9266,N_9231);
nor U9547 (N_9547,N_9284,N_9304);
xnor U9548 (N_9548,N_9326,N_9228);
or U9549 (N_9549,N_9389,N_9288);
xnor U9550 (N_9550,N_9318,N_9286);
and U9551 (N_9551,N_9254,N_9382);
nor U9552 (N_9552,N_9331,N_9341);
or U9553 (N_9553,N_9275,N_9230);
or U9554 (N_9554,N_9228,N_9388);
nor U9555 (N_9555,N_9314,N_9309);
and U9556 (N_9556,N_9320,N_9265);
and U9557 (N_9557,N_9272,N_9345);
xor U9558 (N_9558,N_9279,N_9253);
nor U9559 (N_9559,N_9397,N_9309);
xnor U9560 (N_9560,N_9383,N_9212);
xnor U9561 (N_9561,N_9291,N_9366);
xor U9562 (N_9562,N_9211,N_9267);
and U9563 (N_9563,N_9397,N_9292);
nand U9564 (N_9564,N_9272,N_9204);
nand U9565 (N_9565,N_9323,N_9308);
nand U9566 (N_9566,N_9312,N_9318);
and U9567 (N_9567,N_9389,N_9243);
xor U9568 (N_9568,N_9211,N_9277);
nand U9569 (N_9569,N_9271,N_9333);
xor U9570 (N_9570,N_9221,N_9235);
and U9571 (N_9571,N_9227,N_9340);
nand U9572 (N_9572,N_9213,N_9275);
xor U9573 (N_9573,N_9327,N_9346);
xor U9574 (N_9574,N_9347,N_9329);
nor U9575 (N_9575,N_9207,N_9266);
or U9576 (N_9576,N_9237,N_9255);
and U9577 (N_9577,N_9275,N_9302);
nand U9578 (N_9578,N_9212,N_9398);
and U9579 (N_9579,N_9208,N_9286);
nor U9580 (N_9580,N_9233,N_9298);
nand U9581 (N_9581,N_9237,N_9247);
nand U9582 (N_9582,N_9368,N_9355);
and U9583 (N_9583,N_9368,N_9200);
or U9584 (N_9584,N_9341,N_9333);
or U9585 (N_9585,N_9205,N_9282);
and U9586 (N_9586,N_9207,N_9311);
nand U9587 (N_9587,N_9362,N_9394);
or U9588 (N_9588,N_9203,N_9294);
nor U9589 (N_9589,N_9288,N_9374);
nand U9590 (N_9590,N_9366,N_9347);
nor U9591 (N_9591,N_9313,N_9350);
and U9592 (N_9592,N_9340,N_9248);
nor U9593 (N_9593,N_9252,N_9251);
nor U9594 (N_9594,N_9258,N_9206);
xnor U9595 (N_9595,N_9238,N_9298);
nand U9596 (N_9596,N_9206,N_9200);
xnor U9597 (N_9597,N_9345,N_9319);
or U9598 (N_9598,N_9336,N_9262);
nor U9599 (N_9599,N_9213,N_9250);
nor U9600 (N_9600,N_9500,N_9596);
nor U9601 (N_9601,N_9597,N_9423);
xnor U9602 (N_9602,N_9468,N_9572);
or U9603 (N_9603,N_9426,N_9485);
nor U9604 (N_9604,N_9408,N_9466);
or U9605 (N_9605,N_9402,N_9411);
xnor U9606 (N_9606,N_9440,N_9444);
xor U9607 (N_9607,N_9527,N_9507);
or U9608 (N_9608,N_9516,N_9593);
xnor U9609 (N_9609,N_9584,N_9587);
or U9610 (N_9610,N_9523,N_9538);
and U9611 (N_9611,N_9595,N_9479);
nor U9612 (N_9612,N_9472,N_9561);
and U9613 (N_9613,N_9471,N_9414);
or U9614 (N_9614,N_9429,N_9469);
and U9615 (N_9615,N_9412,N_9547);
nand U9616 (N_9616,N_9432,N_9544);
or U9617 (N_9617,N_9583,N_9409);
or U9618 (N_9618,N_9588,N_9499);
xnor U9619 (N_9619,N_9439,N_9501);
nor U9620 (N_9620,N_9589,N_9556);
and U9621 (N_9621,N_9450,N_9590);
xor U9622 (N_9622,N_9577,N_9515);
or U9623 (N_9623,N_9497,N_9415);
nor U9624 (N_9624,N_9449,N_9553);
nand U9625 (N_9625,N_9457,N_9484);
xnor U9626 (N_9626,N_9433,N_9420);
nand U9627 (N_9627,N_9416,N_9438);
nor U9628 (N_9628,N_9566,N_9579);
and U9629 (N_9629,N_9502,N_9585);
nand U9630 (N_9630,N_9534,N_9563);
nor U9631 (N_9631,N_9418,N_9529);
xnor U9632 (N_9632,N_9537,N_9506);
nand U9633 (N_9633,N_9511,N_9434);
nor U9634 (N_9634,N_9480,N_9552);
nor U9635 (N_9635,N_9573,N_9571);
and U9636 (N_9636,N_9526,N_9513);
or U9637 (N_9637,N_9521,N_9549);
xor U9638 (N_9638,N_9442,N_9568);
or U9639 (N_9639,N_9405,N_9427);
or U9640 (N_9640,N_9581,N_9532);
nand U9641 (N_9641,N_9461,N_9454);
or U9642 (N_9642,N_9483,N_9533);
nand U9643 (N_9643,N_9447,N_9536);
nand U9644 (N_9644,N_9465,N_9540);
or U9645 (N_9645,N_9522,N_9413);
or U9646 (N_9646,N_9504,N_9417);
nor U9647 (N_9647,N_9481,N_9452);
or U9648 (N_9648,N_9419,N_9524);
or U9649 (N_9649,N_9475,N_9464);
nor U9650 (N_9650,N_9594,N_9430);
and U9651 (N_9651,N_9512,N_9493);
xor U9652 (N_9652,N_9564,N_9559);
or U9653 (N_9653,N_9435,N_9558);
xor U9654 (N_9654,N_9598,N_9491);
nand U9655 (N_9655,N_9498,N_9467);
or U9656 (N_9656,N_9599,N_9539);
xor U9657 (N_9657,N_9489,N_9578);
or U9658 (N_9658,N_9428,N_9508);
and U9659 (N_9659,N_9463,N_9531);
nand U9660 (N_9660,N_9448,N_9407);
or U9661 (N_9661,N_9494,N_9477);
nand U9662 (N_9662,N_9586,N_9482);
and U9663 (N_9663,N_9410,N_9554);
nand U9664 (N_9664,N_9446,N_9459);
nor U9665 (N_9665,N_9495,N_9574);
xor U9666 (N_9666,N_9421,N_9528);
or U9667 (N_9667,N_9496,N_9505);
and U9668 (N_9668,N_9406,N_9514);
or U9669 (N_9669,N_9575,N_9555);
nor U9670 (N_9670,N_9422,N_9403);
nor U9671 (N_9671,N_9557,N_9548);
nand U9672 (N_9672,N_9488,N_9487);
xor U9673 (N_9673,N_9517,N_9530);
or U9674 (N_9674,N_9401,N_9567);
nand U9675 (N_9675,N_9455,N_9476);
and U9676 (N_9676,N_9492,N_9535);
nor U9677 (N_9677,N_9562,N_9570);
nor U9678 (N_9678,N_9509,N_9456);
or U9679 (N_9679,N_9543,N_9569);
or U9680 (N_9680,N_9443,N_9424);
nand U9681 (N_9681,N_9545,N_9404);
nand U9682 (N_9682,N_9591,N_9436);
nand U9683 (N_9683,N_9431,N_9550);
xnor U9684 (N_9684,N_9400,N_9474);
or U9685 (N_9685,N_9490,N_9510);
or U9686 (N_9686,N_9478,N_9541);
nor U9687 (N_9687,N_9565,N_9460);
nor U9688 (N_9688,N_9437,N_9453);
nor U9689 (N_9689,N_9525,N_9462);
and U9690 (N_9690,N_9441,N_9425);
xor U9691 (N_9691,N_9520,N_9560);
or U9692 (N_9692,N_9486,N_9592);
or U9693 (N_9693,N_9470,N_9451);
or U9694 (N_9694,N_9518,N_9542);
or U9695 (N_9695,N_9580,N_9546);
xnor U9696 (N_9696,N_9576,N_9582);
and U9697 (N_9697,N_9519,N_9551);
nand U9698 (N_9698,N_9445,N_9503);
nor U9699 (N_9699,N_9473,N_9458);
nand U9700 (N_9700,N_9425,N_9515);
or U9701 (N_9701,N_9514,N_9509);
xor U9702 (N_9702,N_9420,N_9424);
xor U9703 (N_9703,N_9441,N_9590);
and U9704 (N_9704,N_9568,N_9550);
nand U9705 (N_9705,N_9417,N_9409);
xor U9706 (N_9706,N_9469,N_9450);
and U9707 (N_9707,N_9515,N_9570);
nor U9708 (N_9708,N_9500,N_9432);
and U9709 (N_9709,N_9450,N_9428);
nand U9710 (N_9710,N_9461,N_9445);
nor U9711 (N_9711,N_9437,N_9510);
and U9712 (N_9712,N_9565,N_9438);
and U9713 (N_9713,N_9415,N_9528);
xnor U9714 (N_9714,N_9576,N_9598);
xnor U9715 (N_9715,N_9582,N_9588);
nor U9716 (N_9716,N_9461,N_9558);
and U9717 (N_9717,N_9570,N_9516);
xnor U9718 (N_9718,N_9522,N_9501);
nor U9719 (N_9719,N_9445,N_9405);
nor U9720 (N_9720,N_9461,N_9587);
xor U9721 (N_9721,N_9485,N_9542);
or U9722 (N_9722,N_9460,N_9470);
nand U9723 (N_9723,N_9585,N_9482);
and U9724 (N_9724,N_9433,N_9431);
and U9725 (N_9725,N_9542,N_9470);
xor U9726 (N_9726,N_9487,N_9508);
or U9727 (N_9727,N_9569,N_9514);
or U9728 (N_9728,N_9542,N_9581);
or U9729 (N_9729,N_9539,N_9575);
and U9730 (N_9730,N_9457,N_9492);
xor U9731 (N_9731,N_9492,N_9458);
nand U9732 (N_9732,N_9487,N_9481);
and U9733 (N_9733,N_9461,N_9583);
xnor U9734 (N_9734,N_9409,N_9451);
nand U9735 (N_9735,N_9587,N_9496);
xnor U9736 (N_9736,N_9549,N_9533);
xnor U9737 (N_9737,N_9496,N_9599);
nand U9738 (N_9738,N_9404,N_9533);
or U9739 (N_9739,N_9458,N_9512);
and U9740 (N_9740,N_9558,N_9513);
nand U9741 (N_9741,N_9478,N_9528);
nor U9742 (N_9742,N_9553,N_9596);
nand U9743 (N_9743,N_9526,N_9565);
nor U9744 (N_9744,N_9538,N_9415);
or U9745 (N_9745,N_9560,N_9590);
nor U9746 (N_9746,N_9415,N_9555);
xor U9747 (N_9747,N_9528,N_9498);
and U9748 (N_9748,N_9444,N_9584);
and U9749 (N_9749,N_9455,N_9410);
nor U9750 (N_9750,N_9491,N_9569);
xor U9751 (N_9751,N_9501,N_9568);
and U9752 (N_9752,N_9546,N_9596);
nor U9753 (N_9753,N_9413,N_9451);
nand U9754 (N_9754,N_9576,N_9546);
xor U9755 (N_9755,N_9526,N_9472);
nor U9756 (N_9756,N_9471,N_9428);
and U9757 (N_9757,N_9490,N_9574);
nor U9758 (N_9758,N_9401,N_9587);
xnor U9759 (N_9759,N_9529,N_9450);
nand U9760 (N_9760,N_9595,N_9418);
nand U9761 (N_9761,N_9472,N_9589);
and U9762 (N_9762,N_9581,N_9529);
nand U9763 (N_9763,N_9505,N_9544);
or U9764 (N_9764,N_9510,N_9406);
or U9765 (N_9765,N_9513,N_9410);
and U9766 (N_9766,N_9577,N_9574);
nand U9767 (N_9767,N_9471,N_9581);
nand U9768 (N_9768,N_9560,N_9577);
nor U9769 (N_9769,N_9562,N_9406);
xnor U9770 (N_9770,N_9470,N_9445);
nand U9771 (N_9771,N_9435,N_9475);
or U9772 (N_9772,N_9558,N_9503);
nor U9773 (N_9773,N_9446,N_9508);
xnor U9774 (N_9774,N_9507,N_9417);
nor U9775 (N_9775,N_9548,N_9571);
nand U9776 (N_9776,N_9574,N_9570);
and U9777 (N_9777,N_9499,N_9442);
xnor U9778 (N_9778,N_9462,N_9519);
and U9779 (N_9779,N_9512,N_9410);
or U9780 (N_9780,N_9503,N_9447);
and U9781 (N_9781,N_9529,N_9523);
nand U9782 (N_9782,N_9595,N_9494);
nand U9783 (N_9783,N_9523,N_9546);
xor U9784 (N_9784,N_9568,N_9562);
nor U9785 (N_9785,N_9428,N_9558);
and U9786 (N_9786,N_9551,N_9442);
or U9787 (N_9787,N_9474,N_9499);
nand U9788 (N_9788,N_9562,N_9531);
xnor U9789 (N_9789,N_9598,N_9561);
xor U9790 (N_9790,N_9498,N_9500);
nand U9791 (N_9791,N_9584,N_9571);
or U9792 (N_9792,N_9577,N_9537);
nor U9793 (N_9793,N_9421,N_9507);
xor U9794 (N_9794,N_9426,N_9459);
xnor U9795 (N_9795,N_9572,N_9583);
nor U9796 (N_9796,N_9596,N_9506);
or U9797 (N_9797,N_9448,N_9478);
xnor U9798 (N_9798,N_9535,N_9458);
nand U9799 (N_9799,N_9426,N_9452);
nor U9800 (N_9800,N_9695,N_9738);
and U9801 (N_9801,N_9788,N_9679);
and U9802 (N_9802,N_9605,N_9707);
nor U9803 (N_9803,N_9762,N_9630);
or U9804 (N_9804,N_9652,N_9631);
nor U9805 (N_9805,N_9799,N_9722);
xnor U9806 (N_9806,N_9608,N_9719);
xor U9807 (N_9807,N_9743,N_9637);
and U9808 (N_9808,N_9646,N_9639);
or U9809 (N_9809,N_9779,N_9622);
nand U9810 (N_9810,N_9697,N_9658);
nor U9811 (N_9811,N_9632,N_9665);
xor U9812 (N_9812,N_9663,N_9737);
xor U9813 (N_9813,N_9728,N_9681);
and U9814 (N_9814,N_9627,N_9619);
or U9815 (N_9815,N_9749,N_9772);
and U9816 (N_9816,N_9791,N_9671);
or U9817 (N_9817,N_9636,N_9773);
xor U9818 (N_9818,N_9684,N_9690);
and U9819 (N_9819,N_9763,N_9625);
nor U9820 (N_9820,N_9700,N_9698);
and U9821 (N_9821,N_9672,N_9611);
nand U9822 (N_9822,N_9733,N_9689);
nor U9823 (N_9823,N_9613,N_9668);
and U9824 (N_9824,N_9696,N_9606);
xnor U9825 (N_9825,N_9752,N_9640);
nand U9826 (N_9826,N_9699,N_9694);
or U9827 (N_9827,N_9651,N_9674);
nor U9828 (N_9828,N_9742,N_9648);
xnor U9829 (N_9829,N_9604,N_9601);
and U9830 (N_9830,N_9629,N_9670);
nand U9831 (N_9831,N_9621,N_9705);
and U9832 (N_9832,N_9778,N_9785);
or U9833 (N_9833,N_9677,N_9784);
xor U9834 (N_9834,N_9720,N_9615);
nand U9835 (N_9835,N_9740,N_9771);
nand U9836 (N_9836,N_9660,N_9715);
and U9837 (N_9837,N_9724,N_9798);
xnor U9838 (N_9838,N_9732,N_9711);
and U9839 (N_9839,N_9675,N_9747);
and U9840 (N_9840,N_9756,N_9692);
nor U9841 (N_9841,N_9612,N_9755);
nor U9842 (N_9842,N_9777,N_9664);
and U9843 (N_9843,N_9618,N_9610);
nor U9844 (N_9844,N_9769,N_9680);
nand U9845 (N_9845,N_9795,N_9662);
xnor U9846 (N_9846,N_9787,N_9653);
xnor U9847 (N_9847,N_9642,N_9641);
nor U9848 (N_9848,N_9725,N_9776);
nand U9849 (N_9849,N_9766,N_9765);
nand U9850 (N_9850,N_9710,N_9734);
or U9851 (N_9851,N_9770,N_9688);
xor U9852 (N_9852,N_9713,N_9757);
or U9853 (N_9853,N_9656,N_9667);
nor U9854 (N_9854,N_9716,N_9623);
nor U9855 (N_9855,N_9617,N_9761);
nand U9856 (N_9856,N_9616,N_9600);
or U9857 (N_9857,N_9794,N_9644);
or U9858 (N_9858,N_9714,N_9673);
xnor U9859 (N_9859,N_9659,N_9753);
and U9860 (N_9860,N_9635,N_9687);
xor U9861 (N_9861,N_9709,N_9796);
or U9862 (N_9862,N_9645,N_9745);
nor U9863 (N_9863,N_9751,N_9661);
and U9864 (N_9864,N_9614,N_9638);
nand U9865 (N_9865,N_9628,N_9774);
or U9866 (N_9866,N_9726,N_9634);
and U9867 (N_9867,N_9633,N_9767);
nor U9868 (N_9868,N_9704,N_9706);
or U9869 (N_9869,N_9786,N_9602);
and U9870 (N_9870,N_9702,N_9760);
nand U9871 (N_9871,N_9754,N_9708);
or U9872 (N_9872,N_9647,N_9654);
and U9873 (N_9873,N_9731,N_9683);
xor U9874 (N_9874,N_9603,N_9620);
or U9875 (N_9875,N_9729,N_9650);
nand U9876 (N_9876,N_9739,N_9775);
and U9877 (N_9877,N_9701,N_9741);
and U9878 (N_9878,N_9792,N_9721);
xor U9879 (N_9879,N_9759,N_9666);
nand U9880 (N_9880,N_9678,N_9693);
or U9881 (N_9881,N_9718,N_9768);
and U9882 (N_9882,N_9685,N_9780);
and U9883 (N_9883,N_9626,N_9797);
nand U9884 (N_9884,N_9758,N_9655);
nand U9885 (N_9885,N_9643,N_9691);
and U9886 (N_9886,N_9669,N_9723);
xnor U9887 (N_9887,N_9657,N_9746);
nand U9888 (N_9888,N_9735,N_9748);
or U9889 (N_9889,N_9789,N_9730);
nor U9890 (N_9890,N_9790,N_9712);
or U9891 (N_9891,N_9781,N_9607);
xor U9892 (N_9892,N_9744,N_9727);
or U9893 (N_9893,N_9682,N_9736);
or U9894 (N_9894,N_9783,N_9764);
nand U9895 (N_9895,N_9717,N_9703);
and U9896 (N_9896,N_9609,N_9624);
nor U9897 (N_9897,N_9750,N_9793);
nand U9898 (N_9898,N_9686,N_9782);
xnor U9899 (N_9899,N_9649,N_9676);
nor U9900 (N_9900,N_9674,N_9673);
nor U9901 (N_9901,N_9768,N_9616);
and U9902 (N_9902,N_9780,N_9617);
or U9903 (N_9903,N_9703,N_9720);
and U9904 (N_9904,N_9723,N_9786);
nor U9905 (N_9905,N_9673,N_9761);
nand U9906 (N_9906,N_9703,N_9755);
nor U9907 (N_9907,N_9789,N_9751);
nand U9908 (N_9908,N_9781,N_9700);
nor U9909 (N_9909,N_9698,N_9792);
and U9910 (N_9910,N_9626,N_9747);
nand U9911 (N_9911,N_9757,N_9641);
nand U9912 (N_9912,N_9723,N_9607);
xor U9913 (N_9913,N_9702,N_9686);
or U9914 (N_9914,N_9669,N_9649);
and U9915 (N_9915,N_9703,N_9708);
and U9916 (N_9916,N_9690,N_9617);
and U9917 (N_9917,N_9692,N_9688);
or U9918 (N_9918,N_9648,N_9665);
xnor U9919 (N_9919,N_9707,N_9718);
and U9920 (N_9920,N_9711,N_9699);
or U9921 (N_9921,N_9631,N_9716);
nand U9922 (N_9922,N_9647,N_9722);
nand U9923 (N_9923,N_9767,N_9628);
nor U9924 (N_9924,N_9777,N_9741);
and U9925 (N_9925,N_9763,N_9675);
xor U9926 (N_9926,N_9637,N_9747);
or U9927 (N_9927,N_9753,N_9647);
nor U9928 (N_9928,N_9657,N_9600);
and U9929 (N_9929,N_9748,N_9688);
nand U9930 (N_9930,N_9767,N_9789);
xnor U9931 (N_9931,N_9625,N_9721);
xnor U9932 (N_9932,N_9689,N_9699);
nand U9933 (N_9933,N_9706,N_9708);
xnor U9934 (N_9934,N_9664,N_9670);
xor U9935 (N_9935,N_9746,N_9630);
nor U9936 (N_9936,N_9609,N_9767);
nor U9937 (N_9937,N_9694,N_9706);
nor U9938 (N_9938,N_9787,N_9610);
and U9939 (N_9939,N_9729,N_9636);
nor U9940 (N_9940,N_9791,N_9717);
nor U9941 (N_9941,N_9750,N_9746);
nor U9942 (N_9942,N_9722,N_9604);
nor U9943 (N_9943,N_9632,N_9604);
nor U9944 (N_9944,N_9780,N_9638);
xor U9945 (N_9945,N_9617,N_9774);
and U9946 (N_9946,N_9754,N_9773);
nand U9947 (N_9947,N_9620,N_9702);
xnor U9948 (N_9948,N_9761,N_9689);
or U9949 (N_9949,N_9620,N_9716);
nor U9950 (N_9950,N_9651,N_9730);
xor U9951 (N_9951,N_9745,N_9692);
nand U9952 (N_9952,N_9681,N_9692);
or U9953 (N_9953,N_9625,N_9615);
nor U9954 (N_9954,N_9791,N_9693);
nor U9955 (N_9955,N_9770,N_9742);
xnor U9956 (N_9956,N_9627,N_9772);
xor U9957 (N_9957,N_9751,N_9612);
nand U9958 (N_9958,N_9703,N_9722);
and U9959 (N_9959,N_9717,N_9620);
nor U9960 (N_9960,N_9674,N_9777);
nor U9961 (N_9961,N_9703,N_9764);
nor U9962 (N_9962,N_9614,N_9784);
nand U9963 (N_9963,N_9709,N_9664);
xnor U9964 (N_9964,N_9734,N_9742);
or U9965 (N_9965,N_9703,N_9678);
nand U9966 (N_9966,N_9725,N_9744);
or U9967 (N_9967,N_9770,N_9722);
nor U9968 (N_9968,N_9693,N_9611);
xnor U9969 (N_9969,N_9731,N_9671);
and U9970 (N_9970,N_9734,N_9724);
xor U9971 (N_9971,N_9677,N_9710);
and U9972 (N_9972,N_9795,N_9642);
and U9973 (N_9973,N_9663,N_9608);
or U9974 (N_9974,N_9764,N_9650);
or U9975 (N_9975,N_9739,N_9776);
nor U9976 (N_9976,N_9722,N_9679);
xnor U9977 (N_9977,N_9632,N_9679);
xnor U9978 (N_9978,N_9701,N_9690);
nor U9979 (N_9979,N_9766,N_9725);
nor U9980 (N_9980,N_9685,N_9751);
nand U9981 (N_9981,N_9773,N_9701);
and U9982 (N_9982,N_9712,N_9679);
or U9983 (N_9983,N_9619,N_9721);
and U9984 (N_9984,N_9692,N_9797);
and U9985 (N_9985,N_9722,N_9619);
and U9986 (N_9986,N_9670,N_9644);
xor U9987 (N_9987,N_9644,N_9673);
nor U9988 (N_9988,N_9794,N_9603);
nand U9989 (N_9989,N_9680,N_9613);
nor U9990 (N_9990,N_9638,N_9756);
or U9991 (N_9991,N_9733,N_9714);
or U9992 (N_9992,N_9701,N_9672);
nand U9993 (N_9993,N_9780,N_9779);
and U9994 (N_9994,N_9788,N_9664);
nand U9995 (N_9995,N_9776,N_9688);
xnor U9996 (N_9996,N_9738,N_9705);
and U9997 (N_9997,N_9680,N_9686);
or U9998 (N_9998,N_9634,N_9676);
and U9999 (N_9999,N_9626,N_9632);
and U10000 (N_10000,N_9848,N_9851);
nor U10001 (N_10001,N_9979,N_9961);
nand U10002 (N_10002,N_9839,N_9958);
nand U10003 (N_10003,N_9951,N_9937);
xnor U10004 (N_10004,N_9941,N_9909);
and U10005 (N_10005,N_9931,N_9995);
and U10006 (N_10006,N_9802,N_9900);
and U10007 (N_10007,N_9868,N_9967);
xnor U10008 (N_10008,N_9946,N_9817);
xor U10009 (N_10009,N_9956,N_9996);
xor U10010 (N_10010,N_9828,N_9815);
xnor U10011 (N_10011,N_9975,N_9838);
nor U10012 (N_10012,N_9897,N_9891);
or U10013 (N_10013,N_9919,N_9861);
and U10014 (N_10014,N_9903,N_9883);
xnor U10015 (N_10015,N_9800,N_9843);
and U10016 (N_10016,N_9968,N_9882);
nor U10017 (N_10017,N_9904,N_9982);
and U10018 (N_10018,N_9929,N_9948);
or U10019 (N_10019,N_9927,N_9911);
xnor U10020 (N_10020,N_9879,N_9806);
and U10021 (N_10021,N_9976,N_9940);
nand U10022 (N_10022,N_9990,N_9847);
or U10023 (N_10023,N_9863,N_9952);
xnor U10024 (N_10024,N_9874,N_9998);
and U10025 (N_10025,N_9853,N_9965);
nand U10026 (N_10026,N_9824,N_9939);
nor U10027 (N_10027,N_9859,N_9814);
or U10028 (N_10028,N_9860,N_9962);
and U10029 (N_10029,N_9983,N_9978);
or U10030 (N_10030,N_9942,N_9905);
nor U10031 (N_10031,N_9811,N_9819);
or U10032 (N_10032,N_9857,N_9886);
nor U10033 (N_10033,N_9943,N_9888);
nand U10034 (N_10034,N_9823,N_9974);
and U10035 (N_10035,N_9841,N_9934);
nand U10036 (N_10036,N_9991,N_9833);
or U10037 (N_10037,N_9821,N_9932);
and U10038 (N_10038,N_9826,N_9960);
or U10039 (N_10039,N_9807,N_9878);
nor U10040 (N_10040,N_9953,N_9920);
and U10041 (N_10041,N_9969,N_9850);
or U10042 (N_10042,N_9987,N_9812);
nand U10043 (N_10043,N_9981,N_9926);
xnor U10044 (N_10044,N_9877,N_9816);
or U10045 (N_10045,N_9984,N_9836);
nor U10046 (N_10046,N_9892,N_9872);
nor U10047 (N_10047,N_9849,N_9894);
and U10048 (N_10048,N_9915,N_9936);
nor U10049 (N_10049,N_9906,N_9963);
and U10050 (N_10050,N_9856,N_9884);
xor U10051 (N_10051,N_9966,N_9930);
nor U10052 (N_10052,N_9852,N_9999);
xor U10053 (N_10053,N_9993,N_9858);
and U10054 (N_10054,N_9805,N_9801);
xnor U10055 (N_10055,N_9989,N_9855);
and U10056 (N_10056,N_9923,N_9908);
nand U10057 (N_10057,N_9870,N_9921);
nand U10058 (N_10058,N_9885,N_9820);
xnor U10059 (N_10059,N_9871,N_9970);
and U10060 (N_10060,N_9954,N_9804);
xor U10061 (N_10061,N_9898,N_9895);
nor U10062 (N_10062,N_9917,N_9980);
nand U10063 (N_10063,N_9947,N_9831);
and U10064 (N_10064,N_9832,N_9950);
or U10065 (N_10065,N_9822,N_9865);
nand U10066 (N_10066,N_9840,N_9835);
or U10067 (N_10067,N_9866,N_9876);
nor U10068 (N_10068,N_9869,N_9864);
and U10069 (N_10069,N_9867,N_9933);
or U10070 (N_10070,N_9837,N_9994);
nor U10071 (N_10071,N_9827,N_9829);
and U10072 (N_10072,N_9935,N_9834);
xor U10073 (N_10073,N_9809,N_9890);
and U10074 (N_10074,N_9972,N_9893);
or U10075 (N_10075,N_9887,N_9844);
xor U10076 (N_10076,N_9988,N_9964);
xnor U10077 (N_10077,N_9955,N_9924);
nor U10078 (N_10078,N_9825,N_9845);
and U10079 (N_10079,N_9875,N_9986);
nand U10080 (N_10080,N_9889,N_9912);
or U10081 (N_10081,N_9914,N_9902);
or U10082 (N_10082,N_9997,N_9818);
and U10083 (N_10083,N_9803,N_9813);
xor U10084 (N_10084,N_9973,N_9907);
or U10085 (N_10085,N_9810,N_9925);
nor U10086 (N_10086,N_9913,N_9842);
nand U10087 (N_10087,N_9910,N_9992);
and U10088 (N_10088,N_9945,N_9949);
xor U10089 (N_10089,N_9881,N_9880);
or U10090 (N_10090,N_9873,N_9918);
or U10091 (N_10091,N_9938,N_9830);
xnor U10092 (N_10092,N_9985,N_9928);
and U10093 (N_10093,N_9944,N_9899);
xor U10094 (N_10094,N_9922,N_9808);
or U10095 (N_10095,N_9896,N_9846);
and U10096 (N_10096,N_9971,N_9901);
nor U10097 (N_10097,N_9959,N_9854);
and U10098 (N_10098,N_9862,N_9977);
or U10099 (N_10099,N_9916,N_9957);
nand U10100 (N_10100,N_9948,N_9907);
xor U10101 (N_10101,N_9971,N_9853);
or U10102 (N_10102,N_9997,N_9971);
nand U10103 (N_10103,N_9826,N_9838);
and U10104 (N_10104,N_9836,N_9936);
and U10105 (N_10105,N_9834,N_9820);
nor U10106 (N_10106,N_9822,N_9885);
or U10107 (N_10107,N_9946,N_9997);
or U10108 (N_10108,N_9989,N_9959);
and U10109 (N_10109,N_9823,N_9990);
nor U10110 (N_10110,N_9850,N_9970);
or U10111 (N_10111,N_9986,N_9860);
and U10112 (N_10112,N_9988,N_9813);
nor U10113 (N_10113,N_9887,N_9842);
and U10114 (N_10114,N_9867,N_9911);
xor U10115 (N_10115,N_9971,N_9808);
or U10116 (N_10116,N_9840,N_9862);
and U10117 (N_10117,N_9868,N_9842);
xnor U10118 (N_10118,N_9948,N_9957);
nand U10119 (N_10119,N_9977,N_9912);
and U10120 (N_10120,N_9944,N_9966);
and U10121 (N_10121,N_9872,N_9950);
nor U10122 (N_10122,N_9980,N_9853);
xor U10123 (N_10123,N_9905,N_9944);
or U10124 (N_10124,N_9840,N_9856);
nand U10125 (N_10125,N_9923,N_9919);
or U10126 (N_10126,N_9999,N_9862);
or U10127 (N_10127,N_9996,N_9945);
and U10128 (N_10128,N_9964,N_9933);
and U10129 (N_10129,N_9944,N_9946);
nand U10130 (N_10130,N_9840,N_9866);
and U10131 (N_10131,N_9997,N_9894);
nand U10132 (N_10132,N_9951,N_9830);
xnor U10133 (N_10133,N_9997,N_9986);
or U10134 (N_10134,N_9956,N_9954);
or U10135 (N_10135,N_9871,N_9908);
nand U10136 (N_10136,N_9802,N_9941);
nand U10137 (N_10137,N_9874,N_9800);
and U10138 (N_10138,N_9916,N_9842);
and U10139 (N_10139,N_9861,N_9911);
xnor U10140 (N_10140,N_9805,N_9940);
xnor U10141 (N_10141,N_9973,N_9813);
or U10142 (N_10142,N_9975,N_9803);
or U10143 (N_10143,N_9887,N_9879);
nand U10144 (N_10144,N_9962,N_9872);
or U10145 (N_10145,N_9980,N_9876);
nand U10146 (N_10146,N_9804,N_9846);
nand U10147 (N_10147,N_9988,N_9809);
and U10148 (N_10148,N_9897,N_9940);
nand U10149 (N_10149,N_9926,N_9819);
or U10150 (N_10150,N_9831,N_9925);
and U10151 (N_10151,N_9915,N_9969);
or U10152 (N_10152,N_9944,N_9962);
nor U10153 (N_10153,N_9965,N_9910);
xor U10154 (N_10154,N_9966,N_9935);
nor U10155 (N_10155,N_9911,N_9906);
or U10156 (N_10156,N_9837,N_9995);
nor U10157 (N_10157,N_9847,N_9881);
nand U10158 (N_10158,N_9944,N_9970);
xor U10159 (N_10159,N_9978,N_9875);
and U10160 (N_10160,N_9866,N_9833);
nand U10161 (N_10161,N_9802,N_9834);
nor U10162 (N_10162,N_9983,N_9900);
nand U10163 (N_10163,N_9954,N_9968);
nand U10164 (N_10164,N_9800,N_9903);
xor U10165 (N_10165,N_9870,N_9881);
xnor U10166 (N_10166,N_9854,N_9836);
and U10167 (N_10167,N_9952,N_9819);
and U10168 (N_10168,N_9864,N_9803);
xnor U10169 (N_10169,N_9888,N_9850);
nor U10170 (N_10170,N_9869,N_9838);
nor U10171 (N_10171,N_9831,N_9913);
or U10172 (N_10172,N_9863,N_9866);
xnor U10173 (N_10173,N_9957,N_9904);
or U10174 (N_10174,N_9982,N_9847);
or U10175 (N_10175,N_9995,N_9994);
and U10176 (N_10176,N_9866,N_9917);
nor U10177 (N_10177,N_9932,N_9900);
xor U10178 (N_10178,N_9945,N_9988);
and U10179 (N_10179,N_9938,N_9969);
and U10180 (N_10180,N_9949,N_9833);
or U10181 (N_10181,N_9973,N_9989);
xnor U10182 (N_10182,N_9840,N_9996);
nor U10183 (N_10183,N_9898,N_9917);
nand U10184 (N_10184,N_9851,N_9882);
or U10185 (N_10185,N_9954,N_9906);
nor U10186 (N_10186,N_9976,N_9879);
and U10187 (N_10187,N_9803,N_9932);
and U10188 (N_10188,N_9878,N_9943);
nor U10189 (N_10189,N_9869,N_9986);
or U10190 (N_10190,N_9931,N_9980);
nand U10191 (N_10191,N_9854,N_9893);
nor U10192 (N_10192,N_9842,N_9909);
nand U10193 (N_10193,N_9826,N_9827);
xnor U10194 (N_10194,N_9840,N_9974);
nand U10195 (N_10195,N_9851,N_9891);
and U10196 (N_10196,N_9851,N_9900);
and U10197 (N_10197,N_9842,N_9911);
xor U10198 (N_10198,N_9942,N_9978);
xnor U10199 (N_10199,N_9961,N_9893);
and U10200 (N_10200,N_10029,N_10019);
or U10201 (N_10201,N_10152,N_10001);
or U10202 (N_10202,N_10113,N_10160);
or U10203 (N_10203,N_10101,N_10169);
nand U10204 (N_10204,N_10031,N_10150);
nor U10205 (N_10205,N_10181,N_10116);
and U10206 (N_10206,N_10036,N_10039);
nor U10207 (N_10207,N_10011,N_10143);
and U10208 (N_10208,N_10078,N_10096);
xor U10209 (N_10209,N_10115,N_10157);
nand U10210 (N_10210,N_10004,N_10089);
nand U10211 (N_10211,N_10154,N_10056);
nand U10212 (N_10212,N_10110,N_10174);
xor U10213 (N_10213,N_10091,N_10017);
nor U10214 (N_10214,N_10025,N_10087);
nor U10215 (N_10215,N_10075,N_10192);
nand U10216 (N_10216,N_10009,N_10074);
or U10217 (N_10217,N_10190,N_10142);
and U10218 (N_10218,N_10083,N_10197);
nor U10219 (N_10219,N_10045,N_10102);
or U10220 (N_10220,N_10023,N_10015);
and U10221 (N_10221,N_10038,N_10191);
nor U10222 (N_10222,N_10135,N_10063);
and U10223 (N_10223,N_10140,N_10168);
nand U10224 (N_10224,N_10007,N_10073);
nand U10225 (N_10225,N_10033,N_10139);
or U10226 (N_10226,N_10093,N_10059);
nand U10227 (N_10227,N_10165,N_10003);
nor U10228 (N_10228,N_10069,N_10054);
and U10229 (N_10229,N_10068,N_10111);
xor U10230 (N_10230,N_10043,N_10055);
nor U10231 (N_10231,N_10076,N_10121);
xnor U10232 (N_10232,N_10196,N_10052);
nand U10233 (N_10233,N_10133,N_10020);
xnor U10234 (N_10234,N_10049,N_10109);
nand U10235 (N_10235,N_10002,N_10030);
xnor U10236 (N_10236,N_10187,N_10067);
nand U10237 (N_10237,N_10041,N_10005);
or U10238 (N_10238,N_10097,N_10026);
nand U10239 (N_10239,N_10141,N_10148);
nand U10240 (N_10240,N_10125,N_10163);
nor U10241 (N_10241,N_10155,N_10183);
nand U10242 (N_10242,N_10048,N_10120);
nor U10243 (N_10243,N_10094,N_10162);
and U10244 (N_10244,N_10086,N_10161);
xor U10245 (N_10245,N_10062,N_10156);
nand U10246 (N_10246,N_10103,N_10095);
and U10247 (N_10247,N_10171,N_10064);
and U10248 (N_10248,N_10189,N_10081);
and U10249 (N_10249,N_10046,N_10184);
and U10250 (N_10250,N_10037,N_10061);
nand U10251 (N_10251,N_10159,N_10130);
nand U10252 (N_10252,N_10066,N_10199);
nand U10253 (N_10253,N_10153,N_10077);
nor U10254 (N_10254,N_10106,N_10042);
and U10255 (N_10255,N_10193,N_10058);
or U10256 (N_10256,N_10178,N_10166);
or U10257 (N_10257,N_10044,N_10092);
and U10258 (N_10258,N_10051,N_10008);
nor U10259 (N_10259,N_10176,N_10022);
xnor U10260 (N_10260,N_10100,N_10173);
xor U10261 (N_10261,N_10071,N_10194);
xor U10262 (N_10262,N_10104,N_10136);
nand U10263 (N_10263,N_10146,N_10032);
and U10264 (N_10264,N_10129,N_10172);
and U10265 (N_10265,N_10167,N_10127);
xnor U10266 (N_10266,N_10119,N_10118);
and U10267 (N_10267,N_10016,N_10158);
or U10268 (N_10268,N_10131,N_10014);
xor U10269 (N_10269,N_10035,N_10164);
and U10270 (N_10270,N_10132,N_10028);
xor U10271 (N_10271,N_10085,N_10185);
xor U10272 (N_10272,N_10182,N_10149);
nor U10273 (N_10273,N_10198,N_10122);
nand U10274 (N_10274,N_10180,N_10105);
or U10275 (N_10275,N_10053,N_10179);
nor U10276 (N_10276,N_10010,N_10088);
nand U10277 (N_10277,N_10040,N_10126);
or U10278 (N_10278,N_10112,N_10147);
nor U10279 (N_10279,N_10057,N_10072);
nor U10280 (N_10280,N_10188,N_10000);
or U10281 (N_10281,N_10034,N_10137);
and U10282 (N_10282,N_10027,N_10070);
xnor U10283 (N_10283,N_10013,N_10012);
nand U10284 (N_10284,N_10084,N_10128);
nand U10285 (N_10285,N_10175,N_10006);
and U10286 (N_10286,N_10079,N_10124);
nand U10287 (N_10287,N_10186,N_10145);
xnor U10288 (N_10288,N_10024,N_10090);
nor U10289 (N_10289,N_10134,N_10050);
or U10290 (N_10290,N_10098,N_10082);
xnor U10291 (N_10291,N_10047,N_10114);
or U10292 (N_10292,N_10021,N_10065);
or U10293 (N_10293,N_10138,N_10107);
and U10294 (N_10294,N_10195,N_10177);
xor U10295 (N_10295,N_10018,N_10151);
nand U10296 (N_10296,N_10080,N_10108);
and U10297 (N_10297,N_10117,N_10060);
or U10298 (N_10298,N_10099,N_10144);
nor U10299 (N_10299,N_10123,N_10170);
or U10300 (N_10300,N_10055,N_10102);
xor U10301 (N_10301,N_10049,N_10061);
or U10302 (N_10302,N_10057,N_10175);
xor U10303 (N_10303,N_10163,N_10095);
nand U10304 (N_10304,N_10005,N_10008);
nor U10305 (N_10305,N_10045,N_10161);
xnor U10306 (N_10306,N_10111,N_10199);
nand U10307 (N_10307,N_10165,N_10106);
nor U10308 (N_10308,N_10036,N_10011);
and U10309 (N_10309,N_10018,N_10063);
xor U10310 (N_10310,N_10129,N_10083);
nor U10311 (N_10311,N_10092,N_10161);
xnor U10312 (N_10312,N_10170,N_10178);
and U10313 (N_10313,N_10047,N_10112);
nand U10314 (N_10314,N_10106,N_10107);
nand U10315 (N_10315,N_10155,N_10044);
nor U10316 (N_10316,N_10141,N_10165);
or U10317 (N_10317,N_10141,N_10069);
xnor U10318 (N_10318,N_10129,N_10069);
nor U10319 (N_10319,N_10121,N_10168);
xnor U10320 (N_10320,N_10072,N_10089);
nor U10321 (N_10321,N_10147,N_10001);
nor U10322 (N_10322,N_10169,N_10172);
nor U10323 (N_10323,N_10088,N_10082);
or U10324 (N_10324,N_10122,N_10030);
nor U10325 (N_10325,N_10159,N_10050);
nand U10326 (N_10326,N_10161,N_10103);
or U10327 (N_10327,N_10194,N_10127);
nor U10328 (N_10328,N_10045,N_10090);
or U10329 (N_10329,N_10015,N_10126);
nor U10330 (N_10330,N_10146,N_10150);
and U10331 (N_10331,N_10010,N_10063);
nand U10332 (N_10332,N_10129,N_10106);
or U10333 (N_10333,N_10170,N_10074);
and U10334 (N_10334,N_10160,N_10135);
and U10335 (N_10335,N_10127,N_10107);
and U10336 (N_10336,N_10112,N_10129);
nor U10337 (N_10337,N_10103,N_10188);
and U10338 (N_10338,N_10168,N_10170);
and U10339 (N_10339,N_10145,N_10052);
nand U10340 (N_10340,N_10095,N_10075);
nand U10341 (N_10341,N_10058,N_10109);
or U10342 (N_10342,N_10049,N_10009);
or U10343 (N_10343,N_10163,N_10036);
nand U10344 (N_10344,N_10177,N_10178);
and U10345 (N_10345,N_10090,N_10159);
nand U10346 (N_10346,N_10042,N_10115);
nand U10347 (N_10347,N_10106,N_10099);
xor U10348 (N_10348,N_10139,N_10095);
or U10349 (N_10349,N_10087,N_10091);
nand U10350 (N_10350,N_10195,N_10073);
xor U10351 (N_10351,N_10190,N_10101);
nand U10352 (N_10352,N_10008,N_10193);
nand U10353 (N_10353,N_10102,N_10116);
and U10354 (N_10354,N_10158,N_10166);
xnor U10355 (N_10355,N_10149,N_10105);
nand U10356 (N_10356,N_10164,N_10139);
xnor U10357 (N_10357,N_10177,N_10149);
nand U10358 (N_10358,N_10166,N_10127);
or U10359 (N_10359,N_10018,N_10074);
xor U10360 (N_10360,N_10032,N_10003);
xor U10361 (N_10361,N_10158,N_10075);
nor U10362 (N_10362,N_10174,N_10191);
nor U10363 (N_10363,N_10139,N_10130);
or U10364 (N_10364,N_10106,N_10151);
nor U10365 (N_10365,N_10091,N_10178);
or U10366 (N_10366,N_10081,N_10158);
nor U10367 (N_10367,N_10116,N_10195);
or U10368 (N_10368,N_10061,N_10064);
or U10369 (N_10369,N_10078,N_10130);
nand U10370 (N_10370,N_10154,N_10050);
nand U10371 (N_10371,N_10127,N_10070);
nand U10372 (N_10372,N_10156,N_10021);
and U10373 (N_10373,N_10018,N_10078);
nor U10374 (N_10374,N_10039,N_10110);
nor U10375 (N_10375,N_10131,N_10101);
xnor U10376 (N_10376,N_10133,N_10196);
or U10377 (N_10377,N_10150,N_10139);
nand U10378 (N_10378,N_10035,N_10117);
and U10379 (N_10379,N_10024,N_10010);
or U10380 (N_10380,N_10160,N_10130);
or U10381 (N_10381,N_10009,N_10158);
nor U10382 (N_10382,N_10105,N_10116);
nor U10383 (N_10383,N_10131,N_10072);
xnor U10384 (N_10384,N_10157,N_10062);
nand U10385 (N_10385,N_10008,N_10167);
xor U10386 (N_10386,N_10167,N_10007);
nand U10387 (N_10387,N_10022,N_10089);
or U10388 (N_10388,N_10163,N_10126);
and U10389 (N_10389,N_10188,N_10192);
xor U10390 (N_10390,N_10044,N_10084);
nor U10391 (N_10391,N_10117,N_10194);
or U10392 (N_10392,N_10036,N_10133);
nand U10393 (N_10393,N_10139,N_10161);
nor U10394 (N_10394,N_10060,N_10097);
nor U10395 (N_10395,N_10114,N_10101);
nor U10396 (N_10396,N_10030,N_10028);
xnor U10397 (N_10397,N_10159,N_10074);
xnor U10398 (N_10398,N_10075,N_10064);
and U10399 (N_10399,N_10183,N_10158);
xnor U10400 (N_10400,N_10284,N_10257);
xor U10401 (N_10401,N_10322,N_10200);
or U10402 (N_10402,N_10357,N_10287);
xnor U10403 (N_10403,N_10214,N_10241);
nand U10404 (N_10404,N_10202,N_10304);
nand U10405 (N_10405,N_10333,N_10301);
and U10406 (N_10406,N_10283,N_10383);
and U10407 (N_10407,N_10290,N_10300);
or U10408 (N_10408,N_10204,N_10353);
nor U10409 (N_10409,N_10307,N_10350);
and U10410 (N_10410,N_10210,N_10240);
nor U10411 (N_10411,N_10340,N_10339);
nor U10412 (N_10412,N_10250,N_10334);
xnor U10413 (N_10413,N_10254,N_10272);
or U10414 (N_10414,N_10220,N_10323);
xor U10415 (N_10415,N_10309,N_10341);
nand U10416 (N_10416,N_10327,N_10310);
and U10417 (N_10417,N_10226,N_10303);
or U10418 (N_10418,N_10267,N_10361);
nor U10419 (N_10419,N_10381,N_10354);
nand U10420 (N_10420,N_10293,N_10286);
nor U10421 (N_10421,N_10319,N_10345);
and U10422 (N_10422,N_10230,N_10242);
or U10423 (N_10423,N_10203,N_10251);
nand U10424 (N_10424,N_10302,N_10281);
nor U10425 (N_10425,N_10325,N_10308);
nand U10426 (N_10426,N_10387,N_10278);
nand U10427 (N_10427,N_10374,N_10368);
xnor U10428 (N_10428,N_10270,N_10332);
nor U10429 (N_10429,N_10349,N_10365);
or U10430 (N_10430,N_10306,N_10318);
nand U10431 (N_10431,N_10206,N_10299);
xor U10432 (N_10432,N_10229,N_10385);
xnor U10433 (N_10433,N_10346,N_10363);
and U10434 (N_10434,N_10364,N_10377);
nor U10435 (N_10435,N_10276,N_10378);
or U10436 (N_10436,N_10295,N_10343);
xor U10437 (N_10437,N_10271,N_10273);
nor U10438 (N_10438,N_10296,N_10375);
and U10439 (N_10439,N_10369,N_10285);
xor U10440 (N_10440,N_10305,N_10320);
and U10441 (N_10441,N_10329,N_10233);
nand U10442 (N_10442,N_10397,N_10238);
and U10443 (N_10443,N_10314,N_10212);
or U10444 (N_10444,N_10260,N_10225);
nor U10445 (N_10445,N_10282,N_10298);
xnor U10446 (N_10446,N_10399,N_10382);
or U10447 (N_10447,N_10352,N_10342);
xor U10448 (N_10448,N_10224,N_10288);
and U10449 (N_10449,N_10360,N_10389);
xnor U10450 (N_10450,N_10324,N_10235);
and U10451 (N_10451,N_10213,N_10373);
or U10452 (N_10452,N_10231,N_10312);
or U10453 (N_10453,N_10264,N_10328);
nor U10454 (N_10454,N_10362,N_10217);
and U10455 (N_10455,N_10247,N_10266);
and U10456 (N_10456,N_10249,N_10253);
xor U10457 (N_10457,N_10274,N_10255);
xor U10458 (N_10458,N_10326,N_10236);
nand U10459 (N_10459,N_10315,N_10216);
nand U10460 (N_10460,N_10207,N_10379);
xor U10461 (N_10461,N_10338,N_10313);
nor U10462 (N_10462,N_10367,N_10258);
xor U10463 (N_10463,N_10297,N_10245);
nor U10464 (N_10464,N_10246,N_10205);
and U10465 (N_10465,N_10215,N_10259);
nor U10466 (N_10466,N_10321,N_10391);
nor U10467 (N_10467,N_10201,N_10330);
nor U10468 (N_10468,N_10371,N_10280);
and U10469 (N_10469,N_10372,N_10243);
nand U10470 (N_10470,N_10348,N_10252);
nor U10471 (N_10471,N_10393,N_10223);
nor U10472 (N_10472,N_10394,N_10395);
or U10473 (N_10473,N_10244,N_10316);
nand U10474 (N_10474,N_10358,N_10211);
xnor U10475 (N_10475,N_10292,N_10291);
and U10476 (N_10476,N_10265,N_10390);
nand U10477 (N_10477,N_10398,N_10208);
and U10478 (N_10478,N_10355,N_10222);
and U10479 (N_10479,N_10396,N_10237);
nor U10480 (N_10480,N_10344,N_10227);
nor U10481 (N_10481,N_10356,N_10277);
and U10482 (N_10482,N_10261,N_10269);
nor U10483 (N_10483,N_10386,N_10337);
nand U10484 (N_10484,N_10347,N_10275);
or U10485 (N_10485,N_10359,N_10221);
or U10486 (N_10486,N_10351,N_10331);
nand U10487 (N_10487,N_10218,N_10234);
or U10488 (N_10488,N_10239,N_10335);
and U10489 (N_10489,N_10392,N_10262);
or U10490 (N_10490,N_10209,N_10388);
nor U10491 (N_10491,N_10263,N_10228);
xor U10492 (N_10492,N_10219,N_10279);
and U10493 (N_10493,N_10268,N_10370);
and U10494 (N_10494,N_10336,N_10289);
xor U10495 (N_10495,N_10366,N_10311);
or U10496 (N_10496,N_10256,N_10384);
nand U10497 (N_10497,N_10380,N_10317);
xor U10498 (N_10498,N_10232,N_10294);
nor U10499 (N_10499,N_10248,N_10376);
xnor U10500 (N_10500,N_10390,N_10343);
nand U10501 (N_10501,N_10283,N_10302);
or U10502 (N_10502,N_10323,N_10372);
nand U10503 (N_10503,N_10268,N_10352);
and U10504 (N_10504,N_10397,N_10349);
nand U10505 (N_10505,N_10303,N_10240);
or U10506 (N_10506,N_10308,N_10248);
nor U10507 (N_10507,N_10259,N_10239);
and U10508 (N_10508,N_10366,N_10291);
nor U10509 (N_10509,N_10297,N_10329);
nand U10510 (N_10510,N_10209,N_10251);
nand U10511 (N_10511,N_10247,N_10290);
xor U10512 (N_10512,N_10232,N_10341);
and U10513 (N_10513,N_10303,N_10284);
or U10514 (N_10514,N_10324,N_10339);
nor U10515 (N_10515,N_10394,N_10286);
nor U10516 (N_10516,N_10253,N_10386);
or U10517 (N_10517,N_10369,N_10362);
xor U10518 (N_10518,N_10331,N_10332);
and U10519 (N_10519,N_10394,N_10282);
nand U10520 (N_10520,N_10288,N_10312);
nand U10521 (N_10521,N_10219,N_10202);
and U10522 (N_10522,N_10375,N_10396);
nor U10523 (N_10523,N_10262,N_10365);
nor U10524 (N_10524,N_10282,N_10284);
or U10525 (N_10525,N_10357,N_10231);
nor U10526 (N_10526,N_10266,N_10360);
nor U10527 (N_10527,N_10249,N_10262);
xor U10528 (N_10528,N_10248,N_10395);
or U10529 (N_10529,N_10386,N_10249);
nand U10530 (N_10530,N_10316,N_10212);
and U10531 (N_10531,N_10207,N_10314);
and U10532 (N_10532,N_10217,N_10355);
or U10533 (N_10533,N_10280,N_10266);
nor U10534 (N_10534,N_10395,N_10305);
nand U10535 (N_10535,N_10390,N_10361);
or U10536 (N_10536,N_10399,N_10250);
or U10537 (N_10537,N_10388,N_10287);
or U10538 (N_10538,N_10344,N_10331);
nand U10539 (N_10539,N_10353,N_10302);
nor U10540 (N_10540,N_10308,N_10212);
nand U10541 (N_10541,N_10375,N_10308);
or U10542 (N_10542,N_10251,N_10352);
and U10543 (N_10543,N_10323,N_10327);
and U10544 (N_10544,N_10346,N_10310);
and U10545 (N_10545,N_10368,N_10326);
xor U10546 (N_10546,N_10377,N_10246);
and U10547 (N_10547,N_10253,N_10323);
xor U10548 (N_10548,N_10319,N_10220);
and U10549 (N_10549,N_10381,N_10347);
and U10550 (N_10550,N_10320,N_10373);
and U10551 (N_10551,N_10252,N_10344);
xor U10552 (N_10552,N_10284,N_10398);
nor U10553 (N_10553,N_10276,N_10235);
nand U10554 (N_10554,N_10351,N_10342);
and U10555 (N_10555,N_10284,N_10313);
nor U10556 (N_10556,N_10374,N_10239);
nand U10557 (N_10557,N_10348,N_10220);
nand U10558 (N_10558,N_10350,N_10212);
and U10559 (N_10559,N_10363,N_10254);
xor U10560 (N_10560,N_10207,N_10248);
and U10561 (N_10561,N_10377,N_10210);
and U10562 (N_10562,N_10374,N_10371);
or U10563 (N_10563,N_10280,N_10224);
and U10564 (N_10564,N_10287,N_10281);
and U10565 (N_10565,N_10338,N_10394);
and U10566 (N_10566,N_10244,N_10287);
xnor U10567 (N_10567,N_10264,N_10396);
and U10568 (N_10568,N_10238,N_10213);
xor U10569 (N_10569,N_10250,N_10289);
nor U10570 (N_10570,N_10265,N_10343);
or U10571 (N_10571,N_10381,N_10337);
or U10572 (N_10572,N_10228,N_10237);
or U10573 (N_10573,N_10279,N_10205);
and U10574 (N_10574,N_10237,N_10224);
nor U10575 (N_10575,N_10243,N_10297);
and U10576 (N_10576,N_10246,N_10342);
nand U10577 (N_10577,N_10386,N_10309);
xnor U10578 (N_10578,N_10335,N_10330);
xnor U10579 (N_10579,N_10313,N_10227);
xnor U10580 (N_10580,N_10288,N_10270);
nand U10581 (N_10581,N_10284,N_10376);
or U10582 (N_10582,N_10303,N_10261);
and U10583 (N_10583,N_10217,N_10269);
or U10584 (N_10584,N_10357,N_10281);
nand U10585 (N_10585,N_10237,N_10318);
nor U10586 (N_10586,N_10228,N_10216);
nand U10587 (N_10587,N_10385,N_10329);
nand U10588 (N_10588,N_10254,N_10280);
nand U10589 (N_10589,N_10353,N_10362);
nand U10590 (N_10590,N_10324,N_10338);
nor U10591 (N_10591,N_10282,N_10346);
nand U10592 (N_10592,N_10209,N_10275);
nand U10593 (N_10593,N_10367,N_10397);
nand U10594 (N_10594,N_10267,N_10338);
nor U10595 (N_10595,N_10326,N_10384);
nand U10596 (N_10596,N_10369,N_10331);
and U10597 (N_10597,N_10277,N_10386);
or U10598 (N_10598,N_10329,N_10301);
xor U10599 (N_10599,N_10288,N_10242);
xor U10600 (N_10600,N_10590,N_10596);
nor U10601 (N_10601,N_10538,N_10479);
nand U10602 (N_10602,N_10437,N_10562);
and U10603 (N_10603,N_10540,N_10469);
or U10604 (N_10604,N_10447,N_10543);
nor U10605 (N_10605,N_10511,N_10411);
or U10606 (N_10606,N_10440,N_10442);
and U10607 (N_10607,N_10553,N_10552);
nor U10608 (N_10608,N_10555,N_10514);
and U10609 (N_10609,N_10412,N_10414);
xnor U10610 (N_10610,N_10512,N_10428);
nor U10611 (N_10611,N_10574,N_10401);
and U10612 (N_10612,N_10570,N_10505);
nand U10613 (N_10613,N_10436,N_10489);
nor U10614 (N_10614,N_10498,N_10467);
nand U10615 (N_10615,N_10485,N_10537);
or U10616 (N_10616,N_10515,N_10594);
or U10617 (N_10617,N_10441,N_10406);
xnor U10618 (N_10618,N_10519,N_10577);
nor U10619 (N_10619,N_10460,N_10400);
nand U10620 (N_10620,N_10420,N_10508);
and U10621 (N_10621,N_10539,N_10569);
nand U10622 (N_10622,N_10545,N_10458);
xor U10623 (N_10623,N_10421,N_10547);
nand U10624 (N_10624,N_10535,N_10587);
xnor U10625 (N_10625,N_10471,N_10430);
or U10626 (N_10626,N_10448,N_10528);
nor U10627 (N_10627,N_10483,N_10478);
or U10628 (N_10628,N_10408,N_10459);
nor U10629 (N_10629,N_10410,N_10455);
or U10630 (N_10630,N_10415,N_10571);
or U10631 (N_10631,N_10465,N_10523);
or U10632 (N_10632,N_10532,N_10588);
xor U10633 (N_10633,N_10426,N_10464);
or U10634 (N_10634,N_10443,N_10517);
and U10635 (N_10635,N_10524,N_10502);
xor U10636 (N_10636,N_10536,N_10579);
nor U10637 (N_10637,N_10595,N_10492);
and U10638 (N_10638,N_10445,N_10402);
nand U10639 (N_10639,N_10461,N_10446);
xor U10640 (N_10640,N_10586,N_10598);
xor U10641 (N_10641,N_10500,N_10534);
nand U10642 (N_10642,N_10513,N_10405);
and U10643 (N_10643,N_10476,N_10466);
xnor U10644 (N_10644,N_10403,N_10584);
or U10645 (N_10645,N_10418,N_10518);
xnor U10646 (N_10646,N_10533,N_10407);
or U10647 (N_10647,N_10488,N_10493);
or U10648 (N_10648,N_10435,N_10531);
xnor U10649 (N_10649,N_10453,N_10583);
nand U10650 (N_10650,N_10413,N_10472);
and U10651 (N_10651,N_10561,N_10578);
xnor U10652 (N_10652,N_10495,N_10544);
xor U10653 (N_10653,N_10449,N_10423);
or U10654 (N_10654,N_10431,N_10468);
nand U10655 (N_10655,N_10560,N_10462);
xnor U10656 (N_10656,N_10499,N_10593);
and U10657 (N_10657,N_10549,N_10557);
xor U10658 (N_10658,N_10509,N_10575);
nor U10659 (N_10659,N_10477,N_10527);
and U10660 (N_10660,N_10409,N_10529);
and U10661 (N_10661,N_10422,N_10456);
xor U10662 (N_10662,N_10482,N_10556);
xor U10663 (N_10663,N_10450,N_10567);
and U10664 (N_10664,N_10416,N_10580);
xor U10665 (N_10665,N_10541,N_10444);
nand U10666 (N_10666,N_10490,N_10568);
nor U10667 (N_10667,N_10592,N_10548);
or U10668 (N_10668,N_10457,N_10576);
and U10669 (N_10669,N_10530,N_10486);
xnor U10670 (N_10670,N_10566,N_10484);
nor U10671 (N_10671,N_10554,N_10516);
nand U10672 (N_10672,N_10597,N_10506);
and U10673 (N_10673,N_10551,N_10501);
or U10674 (N_10674,N_10487,N_10419);
or U10675 (N_10675,N_10404,N_10451);
or U10676 (N_10676,N_10454,N_10424);
nor U10677 (N_10677,N_10438,N_10542);
nor U10678 (N_10678,N_10546,N_10525);
xnor U10679 (N_10679,N_10522,N_10463);
nand U10680 (N_10680,N_10425,N_10475);
or U10681 (N_10681,N_10572,N_10497);
and U10682 (N_10682,N_10470,N_10550);
xnor U10683 (N_10683,N_10434,N_10474);
nor U10684 (N_10684,N_10581,N_10429);
nand U10685 (N_10685,N_10427,N_10564);
and U10686 (N_10686,N_10585,N_10481);
nand U10687 (N_10687,N_10494,N_10507);
nand U10688 (N_10688,N_10559,N_10432);
and U10689 (N_10689,N_10573,N_10417);
xor U10690 (N_10690,N_10565,N_10480);
or U10691 (N_10691,N_10563,N_10599);
nand U10692 (N_10692,N_10526,N_10503);
or U10693 (N_10693,N_10496,N_10433);
xor U10694 (N_10694,N_10520,N_10504);
or U10695 (N_10695,N_10439,N_10510);
and U10696 (N_10696,N_10591,N_10582);
nand U10697 (N_10697,N_10558,N_10473);
or U10698 (N_10698,N_10491,N_10589);
nand U10699 (N_10699,N_10521,N_10452);
or U10700 (N_10700,N_10400,N_10441);
and U10701 (N_10701,N_10579,N_10570);
nand U10702 (N_10702,N_10405,N_10521);
and U10703 (N_10703,N_10447,N_10418);
xnor U10704 (N_10704,N_10496,N_10532);
and U10705 (N_10705,N_10411,N_10569);
nor U10706 (N_10706,N_10594,N_10402);
nor U10707 (N_10707,N_10426,N_10547);
xnor U10708 (N_10708,N_10541,N_10408);
nor U10709 (N_10709,N_10425,N_10439);
nor U10710 (N_10710,N_10565,N_10530);
nor U10711 (N_10711,N_10474,N_10412);
nor U10712 (N_10712,N_10403,N_10575);
nor U10713 (N_10713,N_10485,N_10496);
or U10714 (N_10714,N_10556,N_10474);
and U10715 (N_10715,N_10529,N_10502);
nand U10716 (N_10716,N_10450,N_10404);
and U10717 (N_10717,N_10445,N_10574);
or U10718 (N_10718,N_10567,N_10492);
or U10719 (N_10719,N_10488,N_10468);
xor U10720 (N_10720,N_10453,N_10535);
xor U10721 (N_10721,N_10580,N_10477);
or U10722 (N_10722,N_10456,N_10419);
nand U10723 (N_10723,N_10557,N_10492);
or U10724 (N_10724,N_10561,N_10433);
or U10725 (N_10725,N_10453,N_10538);
and U10726 (N_10726,N_10498,N_10450);
and U10727 (N_10727,N_10457,N_10451);
nand U10728 (N_10728,N_10576,N_10536);
nand U10729 (N_10729,N_10455,N_10569);
nand U10730 (N_10730,N_10471,N_10461);
xnor U10731 (N_10731,N_10415,N_10508);
and U10732 (N_10732,N_10563,N_10504);
or U10733 (N_10733,N_10570,N_10434);
and U10734 (N_10734,N_10503,N_10426);
and U10735 (N_10735,N_10525,N_10579);
nor U10736 (N_10736,N_10465,N_10516);
xnor U10737 (N_10737,N_10408,N_10498);
and U10738 (N_10738,N_10546,N_10461);
and U10739 (N_10739,N_10582,N_10499);
or U10740 (N_10740,N_10410,N_10497);
nor U10741 (N_10741,N_10402,N_10438);
nand U10742 (N_10742,N_10453,N_10596);
nand U10743 (N_10743,N_10426,N_10570);
xnor U10744 (N_10744,N_10548,N_10405);
and U10745 (N_10745,N_10500,N_10445);
nor U10746 (N_10746,N_10543,N_10510);
or U10747 (N_10747,N_10482,N_10502);
or U10748 (N_10748,N_10446,N_10536);
or U10749 (N_10749,N_10507,N_10542);
nor U10750 (N_10750,N_10463,N_10419);
and U10751 (N_10751,N_10519,N_10551);
nand U10752 (N_10752,N_10457,N_10514);
nand U10753 (N_10753,N_10426,N_10596);
nor U10754 (N_10754,N_10439,N_10578);
and U10755 (N_10755,N_10506,N_10551);
or U10756 (N_10756,N_10516,N_10459);
and U10757 (N_10757,N_10493,N_10422);
nor U10758 (N_10758,N_10563,N_10492);
nor U10759 (N_10759,N_10532,N_10578);
or U10760 (N_10760,N_10578,N_10550);
nor U10761 (N_10761,N_10489,N_10427);
xnor U10762 (N_10762,N_10455,N_10599);
or U10763 (N_10763,N_10591,N_10448);
or U10764 (N_10764,N_10504,N_10429);
nand U10765 (N_10765,N_10581,N_10432);
and U10766 (N_10766,N_10496,N_10571);
and U10767 (N_10767,N_10544,N_10507);
and U10768 (N_10768,N_10517,N_10455);
xnor U10769 (N_10769,N_10520,N_10558);
and U10770 (N_10770,N_10574,N_10576);
nand U10771 (N_10771,N_10592,N_10436);
nand U10772 (N_10772,N_10418,N_10557);
nor U10773 (N_10773,N_10405,N_10452);
and U10774 (N_10774,N_10402,N_10449);
nor U10775 (N_10775,N_10528,N_10598);
nand U10776 (N_10776,N_10557,N_10536);
nand U10777 (N_10777,N_10508,N_10527);
or U10778 (N_10778,N_10403,N_10591);
and U10779 (N_10779,N_10544,N_10542);
or U10780 (N_10780,N_10551,N_10588);
or U10781 (N_10781,N_10473,N_10417);
or U10782 (N_10782,N_10430,N_10507);
nor U10783 (N_10783,N_10522,N_10438);
and U10784 (N_10784,N_10481,N_10459);
and U10785 (N_10785,N_10496,N_10443);
or U10786 (N_10786,N_10537,N_10553);
or U10787 (N_10787,N_10482,N_10571);
xnor U10788 (N_10788,N_10441,N_10456);
and U10789 (N_10789,N_10558,N_10580);
nand U10790 (N_10790,N_10535,N_10572);
nand U10791 (N_10791,N_10440,N_10534);
and U10792 (N_10792,N_10487,N_10443);
and U10793 (N_10793,N_10410,N_10420);
nand U10794 (N_10794,N_10536,N_10574);
xor U10795 (N_10795,N_10566,N_10402);
xor U10796 (N_10796,N_10574,N_10429);
and U10797 (N_10797,N_10434,N_10433);
xor U10798 (N_10798,N_10480,N_10441);
xor U10799 (N_10799,N_10483,N_10476);
or U10800 (N_10800,N_10750,N_10634);
and U10801 (N_10801,N_10680,N_10651);
or U10802 (N_10802,N_10757,N_10733);
nor U10803 (N_10803,N_10630,N_10642);
xor U10804 (N_10804,N_10646,N_10644);
xor U10805 (N_10805,N_10653,N_10782);
nor U10806 (N_10806,N_10743,N_10789);
nand U10807 (N_10807,N_10697,N_10768);
xor U10808 (N_10808,N_10712,N_10649);
xnor U10809 (N_10809,N_10640,N_10754);
or U10810 (N_10810,N_10667,N_10610);
nor U10811 (N_10811,N_10675,N_10766);
nand U10812 (N_10812,N_10702,N_10775);
nor U10813 (N_10813,N_10688,N_10723);
xor U10814 (N_10814,N_10730,N_10658);
nor U10815 (N_10815,N_10622,N_10607);
nor U10816 (N_10816,N_10618,N_10608);
xnor U10817 (N_10817,N_10660,N_10693);
nor U10818 (N_10818,N_10612,N_10710);
or U10819 (N_10819,N_10691,N_10665);
nor U10820 (N_10820,N_10701,N_10635);
nand U10821 (N_10821,N_10709,N_10783);
and U10822 (N_10822,N_10793,N_10695);
or U10823 (N_10823,N_10752,N_10699);
nor U10824 (N_10824,N_10639,N_10707);
or U10825 (N_10825,N_10767,N_10616);
or U10826 (N_10826,N_10677,N_10625);
nand U10827 (N_10827,N_10736,N_10760);
and U10828 (N_10828,N_10714,N_10601);
or U10829 (N_10829,N_10778,N_10737);
nand U10830 (N_10830,N_10643,N_10682);
nor U10831 (N_10831,N_10609,N_10777);
nor U10832 (N_10832,N_10759,N_10615);
xnor U10833 (N_10833,N_10711,N_10603);
xnor U10834 (N_10834,N_10698,N_10794);
or U10835 (N_10835,N_10687,N_10662);
nand U10836 (N_10836,N_10741,N_10788);
nor U10837 (N_10837,N_10694,N_10657);
and U10838 (N_10838,N_10786,N_10787);
and U10839 (N_10839,N_10755,N_10792);
nand U10840 (N_10840,N_10638,N_10706);
nand U10841 (N_10841,N_10721,N_10748);
xnor U10842 (N_10842,N_10773,N_10690);
and U10843 (N_10843,N_10746,N_10769);
nand U10844 (N_10844,N_10728,N_10774);
or U10845 (N_10845,N_10747,N_10600);
and U10846 (N_10846,N_10685,N_10670);
xnor U10847 (N_10847,N_10655,N_10664);
nand U10848 (N_10848,N_10744,N_10753);
or U10849 (N_10849,N_10708,N_10678);
or U10850 (N_10850,N_10795,N_10731);
xnor U10851 (N_10851,N_10717,N_10722);
or U10852 (N_10852,N_10732,N_10703);
or U10853 (N_10853,N_10790,N_10626);
or U10854 (N_10854,N_10617,N_10669);
and U10855 (N_10855,N_10636,N_10780);
and U10856 (N_10856,N_10650,N_10745);
xnor U10857 (N_10857,N_10656,N_10673);
nand U10858 (N_10858,N_10632,N_10645);
or U10859 (N_10859,N_10674,N_10686);
or U10860 (N_10860,N_10705,N_10765);
or U10861 (N_10861,N_10797,N_10604);
xnor U10862 (N_10862,N_10654,N_10627);
and U10863 (N_10863,N_10734,N_10629);
and U10864 (N_10864,N_10676,N_10666);
nor U10865 (N_10865,N_10772,N_10700);
xnor U10866 (N_10866,N_10623,N_10647);
xnor U10867 (N_10867,N_10692,N_10763);
xnor U10868 (N_10868,N_10724,N_10684);
nand U10869 (N_10869,N_10739,N_10671);
xnor U10870 (N_10870,N_10661,N_10738);
xor U10871 (N_10871,N_10624,N_10631);
xor U10872 (N_10872,N_10611,N_10672);
nand U10873 (N_10873,N_10796,N_10637);
and U10874 (N_10874,N_10663,N_10798);
and U10875 (N_10875,N_10781,N_10681);
xnor U10876 (N_10876,N_10761,N_10758);
and U10877 (N_10877,N_10770,N_10726);
xnor U10878 (N_10878,N_10771,N_10620);
or U10879 (N_10879,N_10784,N_10716);
xnor U10880 (N_10880,N_10641,N_10613);
xnor U10881 (N_10881,N_10619,N_10751);
nor U10882 (N_10882,N_10720,N_10735);
xor U10883 (N_10883,N_10648,N_10628);
or U10884 (N_10884,N_10742,N_10756);
or U10885 (N_10885,N_10762,N_10704);
xor U10886 (N_10886,N_10718,N_10779);
or U10887 (N_10887,N_10785,N_10729);
nand U10888 (N_10888,N_10715,N_10652);
or U10889 (N_10889,N_10776,N_10799);
or U10890 (N_10890,N_10679,N_10605);
nand U10891 (N_10891,N_10606,N_10740);
nand U10892 (N_10892,N_10668,N_10659);
and U10893 (N_10893,N_10749,N_10696);
or U10894 (N_10894,N_10602,N_10621);
xor U10895 (N_10895,N_10719,N_10791);
or U10896 (N_10896,N_10764,N_10683);
and U10897 (N_10897,N_10713,N_10727);
nor U10898 (N_10898,N_10633,N_10614);
nor U10899 (N_10899,N_10725,N_10689);
nand U10900 (N_10900,N_10631,N_10648);
and U10901 (N_10901,N_10633,N_10670);
and U10902 (N_10902,N_10660,N_10775);
nor U10903 (N_10903,N_10636,N_10723);
or U10904 (N_10904,N_10727,N_10631);
or U10905 (N_10905,N_10600,N_10776);
or U10906 (N_10906,N_10747,N_10776);
nand U10907 (N_10907,N_10725,N_10604);
nand U10908 (N_10908,N_10728,N_10799);
or U10909 (N_10909,N_10612,N_10665);
or U10910 (N_10910,N_10694,N_10754);
nor U10911 (N_10911,N_10723,N_10718);
nand U10912 (N_10912,N_10706,N_10679);
xnor U10913 (N_10913,N_10604,N_10751);
and U10914 (N_10914,N_10728,N_10652);
and U10915 (N_10915,N_10620,N_10694);
xnor U10916 (N_10916,N_10699,N_10795);
nor U10917 (N_10917,N_10717,N_10767);
or U10918 (N_10918,N_10773,N_10681);
nand U10919 (N_10919,N_10672,N_10669);
nand U10920 (N_10920,N_10733,N_10731);
and U10921 (N_10921,N_10706,N_10731);
xor U10922 (N_10922,N_10654,N_10622);
nor U10923 (N_10923,N_10770,N_10628);
xor U10924 (N_10924,N_10747,N_10635);
nor U10925 (N_10925,N_10754,N_10651);
xor U10926 (N_10926,N_10752,N_10758);
and U10927 (N_10927,N_10759,N_10770);
xnor U10928 (N_10928,N_10622,N_10739);
nand U10929 (N_10929,N_10787,N_10665);
and U10930 (N_10930,N_10790,N_10709);
xnor U10931 (N_10931,N_10669,N_10664);
nor U10932 (N_10932,N_10676,N_10790);
and U10933 (N_10933,N_10683,N_10626);
nand U10934 (N_10934,N_10607,N_10617);
or U10935 (N_10935,N_10742,N_10675);
xor U10936 (N_10936,N_10770,N_10657);
and U10937 (N_10937,N_10608,N_10657);
or U10938 (N_10938,N_10786,N_10629);
xor U10939 (N_10939,N_10710,N_10651);
or U10940 (N_10940,N_10781,N_10662);
nor U10941 (N_10941,N_10635,N_10704);
nor U10942 (N_10942,N_10675,N_10797);
xnor U10943 (N_10943,N_10746,N_10619);
or U10944 (N_10944,N_10647,N_10673);
nor U10945 (N_10945,N_10763,N_10789);
nand U10946 (N_10946,N_10735,N_10663);
or U10947 (N_10947,N_10747,N_10737);
nor U10948 (N_10948,N_10654,N_10650);
or U10949 (N_10949,N_10754,N_10799);
nor U10950 (N_10950,N_10670,N_10735);
nor U10951 (N_10951,N_10798,N_10708);
and U10952 (N_10952,N_10669,N_10760);
and U10953 (N_10953,N_10763,N_10786);
nor U10954 (N_10954,N_10660,N_10752);
xor U10955 (N_10955,N_10607,N_10787);
xor U10956 (N_10956,N_10741,N_10697);
nand U10957 (N_10957,N_10646,N_10695);
nor U10958 (N_10958,N_10631,N_10625);
or U10959 (N_10959,N_10776,N_10689);
or U10960 (N_10960,N_10673,N_10701);
xnor U10961 (N_10961,N_10756,N_10735);
nor U10962 (N_10962,N_10753,N_10719);
xor U10963 (N_10963,N_10711,N_10762);
and U10964 (N_10964,N_10720,N_10773);
nor U10965 (N_10965,N_10756,N_10644);
xor U10966 (N_10966,N_10794,N_10663);
nor U10967 (N_10967,N_10635,N_10763);
xnor U10968 (N_10968,N_10731,N_10798);
nor U10969 (N_10969,N_10625,N_10670);
xor U10970 (N_10970,N_10784,N_10739);
and U10971 (N_10971,N_10779,N_10770);
nor U10972 (N_10972,N_10616,N_10700);
xnor U10973 (N_10973,N_10612,N_10785);
xnor U10974 (N_10974,N_10772,N_10661);
nor U10975 (N_10975,N_10635,N_10620);
nor U10976 (N_10976,N_10706,N_10656);
nor U10977 (N_10977,N_10673,N_10687);
nand U10978 (N_10978,N_10686,N_10683);
nand U10979 (N_10979,N_10662,N_10771);
xnor U10980 (N_10980,N_10689,N_10656);
nand U10981 (N_10981,N_10708,N_10775);
and U10982 (N_10982,N_10739,N_10760);
nand U10983 (N_10983,N_10621,N_10795);
or U10984 (N_10984,N_10771,N_10764);
xor U10985 (N_10985,N_10637,N_10715);
nor U10986 (N_10986,N_10740,N_10795);
or U10987 (N_10987,N_10623,N_10654);
and U10988 (N_10988,N_10655,N_10637);
xor U10989 (N_10989,N_10680,N_10757);
or U10990 (N_10990,N_10664,N_10676);
nand U10991 (N_10991,N_10716,N_10606);
or U10992 (N_10992,N_10778,N_10711);
xor U10993 (N_10993,N_10663,N_10763);
nand U10994 (N_10994,N_10637,N_10723);
xor U10995 (N_10995,N_10607,N_10750);
nand U10996 (N_10996,N_10794,N_10659);
nand U10997 (N_10997,N_10774,N_10733);
nand U10998 (N_10998,N_10683,N_10608);
and U10999 (N_10999,N_10682,N_10646);
or U11000 (N_11000,N_10942,N_10840);
nand U11001 (N_11001,N_10988,N_10985);
and U11002 (N_11002,N_10885,N_10891);
nor U11003 (N_11003,N_10906,N_10995);
nor U11004 (N_11004,N_10990,N_10803);
xor U11005 (N_11005,N_10883,N_10954);
or U11006 (N_11006,N_10887,N_10959);
or U11007 (N_11007,N_10969,N_10882);
nor U11008 (N_11008,N_10869,N_10807);
xor U11009 (N_11009,N_10968,N_10813);
or U11010 (N_11010,N_10913,N_10839);
xnor U11011 (N_11011,N_10801,N_10831);
nand U11012 (N_11012,N_10931,N_10925);
or U11013 (N_11013,N_10978,N_10987);
or U11014 (N_11014,N_10937,N_10953);
or U11015 (N_11015,N_10889,N_10853);
and U11016 (N_11016,N_10993,N_10881);
xnor U11017 (N_11017,N_10974,N_10980);
xor U11018 (N_11018,N_10917,N_10911);
xnor U11019 (N_11019,N_10905,N_10809);
and U11020 (N_11020,N_10864,N_10874);
and U11021 (N_11021,N_10938,N_10894);
or U11022 (N_11022,N_10895,N_10847);
and U11023 (N_11023,N_10877,N_10863);
xor U11024 (N_11024,N_10902,N_10908);
nor U11025 (N_11025,N_10983,N_10947);
xor U11026 (N_11026,N_10836,N_10884);
nor U11027 (N_11027,N_10832,N_10926);
and U11028 (N_11028,N_10860,N_10868);
nor U11029 (N_11029,N_10818,N_10970);
or U11030 (N_11030,N_10935,N_10963);
and U11031 (N_11031,N_10967,N_10907);
nand U11032 (N_11032,N_10962,N_10867);
nor U11033 (N_11033,N_10823,N_10879);
or U11034 (N_11034,N_10956,N_10945);
nor U11035 (N_11035,N_10944,N_10950);
xor U11036 (N_11036,N_10830,N_10934);
or U11037 (N_11037,N_10851,N_10927);
or U11038 (N_11038,N_10897,N_10855);
or U11039 (N_11039,N_10859,N_10876);
xor U11040 (N_11040,N_10845,N_10930);
nand U11041 (N_11041,N_10837,N_10824);
xor U11042 (N_11042,N_10841,N_10834);
or U11043 (N_11043,N_10920,N_10866);
and U11044 (N_11044,N_10914,N_10886);
nor U11045 (N_11045,N_10904,N_10829);
nor U11046 (N_11046,N_10804,N_10862);
or U11047 (N_11047,N_10856,N_10826);
xnor U11048 (N_11048,N_10939,N_10910);
xor U11049 (N_11049,N_10828,N_10981);
and U11050 (N_11050,N_10991,N_10909);
and U11051 (N_11051,N_10900,N_10903);
and U11052 (N_11052,N_10973,N_10833);
nand U11053 (N_11053,N_10992,N_10940);
nor U11054 (N_11054,N_10806,N_10957);
nand U11055 (N_11055,N_10918,N_10946);
nand U11056 (N_11056,N_10994,N_10848);
or U11057 (N_11057,N_10928,N_10805);
xnor U11058 (N_11058,N_10815,N_10960);
or U11059 (N_11059,N_10852,N_10901);
or U11060 (N_11060,N_10941,N_10989);
nor U11061 (N_11061,N_10955,N_10825);
or U11062 (N_11062,N_10929,N_10933);
nand U11063 (N_11063,N_10916,N_10923);
xor U11064 (N_11064,N_10893,N_10958);
or U11065 (N_11065,N_10854,N_10971);
nor U11066 (N_11066,N_10844,N_10948);
nor U11067 (N_11067,N_10984,N_10865);
xor U11068 (N_11068,N_10936,N_10975);
xnor U11069 (N_11069,N_10977,N_10814);
and U11070 (N_11070,N_10846,N_10820);
nor U11071 (N_11071,N_10808,N_10802);
xnor U11072 (N_11072,N_10878,N_10890);
nor U11073 (N_11073,N_10875,N_10966);
nand U11074 (N_11074,N_10811,N_10872);
and U11075 (N_11075,N_10861,N_10979);
or U11076 (N_11076,N_10800,N_10915);
nand U11077 (N_11077,N_10842,N_10998);
nand U11078 (N_11078,N_10965,N_10819);
and U11079 (N_11079,N_10817,N_10838);
or U11080 (N_11080,N_10982,N_10943);
nand U11081 (N_11081,N_10924,N_10986);
xnor U11082 (N_11082,N_10873,N_10888);
nand U11083 (N_11083,N_10972,N_10997);
and U11084 (N_11084,N_10849,N_10822);
nor U11085 (N_11085,N_10816,N_10961);
or U11086 (N_11086,N_10850,N_10899);
nand U11087 (N_11087,N_10919,N_10835);
or U11088 (N_11088,N_10952,N_10812);
nand U11089 (N_11089,N_10857,N_10810);
nand U11090 (N_11090,N_10843,N_10921);
nor U11091 (N_11091,N_10870,N_10896);
nand U11092 (N_11092,N_10880,N_10996);
nor U11093 (N_11093,N_10827,N_10871);
or U11094 (N_11094,N_10892,N_10912);
and U11095 (N_11095,N_10976,N_10922);
xnor U11096 (N_11096,N_10951,N_10898);
xor U11097 (N_11097,N_10858,N_10964);
xor U11098 (N_11098,N_10949,N_10932);
or U11099 (N_11099,N_10999,N_10821);
xor U11100 (N_11100,N_10925,N_10935);
or U11101 (N_11101,N_10901,N_10929);
nor U11102 (N_11102,N_10840,N_10911);
nand U11103 (N_11103,N_10819,N_10851);
nand U11104 (N_11104,N_10837,N_10808);
nand U11105 (N_11105,N_10909,N_10970);
or U11106 (N_11106,N_10986,N_10867);
or U11107 (N_11107,N_10807,N_10832);
nand U11108 (N_11108,N_10908,N_10854);
nand U11109 (N_11109,N_10939,N_10867);
nor U11110 (N_11110,N_10962,N_10919);
or U11111 (N_11111,N_10902,N_10859);
nand U11112 (N_11112,N_10904,N_10822);
nand U11113 (N_11113,N_10954,N_10834);
or U11114 (N_11114,N_10816,N_10904);
and U11115 (N_11115,N_10856,N_10864);
or U11116 (N_11116,N_10966,N_10965);
and U11117 (N_11117,N_10915,N_10981);
or U11118 (N_11118,N_10991,N_10992);
nor U11119 (N_11119,N_10876,N_10806);
or U11120 (N_11120,N_10902,N_10816);
and U11121 (N_11121,N_10957,N_10892);
nand U11122 (N_11122,N_10987,N_10855);
and U11123 (N_11123,N_10974,N_10897);
xnor U11124 (N_11124,N_10985,N_10867);
nor U11125 (N_11125,N_10894,N_10911);
xor U11126 (N_11126,N_10930,N_10876);
or U11127 (N_11127,N_10904,N_10925);
nor U11128 (N_11128,N_10969,N_10883);
or U11129 (N_11129,N_10906,N_10883);
and U11130 (N_11130,N_10821,N_10969);
nand U11131 (N_11131,N_10872,N_10806);
nand U11132 (N_11132,N_10905,N_10980);
nand U11133 (N_11133,N_10882,N_10880);
xnor U11134 (N_11134,N_10918,N_10904);
nor U11135 (N_11135,N_10878,N_10869);
and U11136 (N_11136,N_10989,N_10999);
nor U11137 (N_11137,N_10864,N_10954);
or U11138 (N_11138,N_10913,N_10957);
and U11139 (N_11139,N_10982,N_10868);
and U11140 (N_11140,N_10996,N_10934);
nand U11141 (N_11141,N_10920,N_10918);
xor U11142 (N_11142,N_10844,N_10914);
nand U11143 (N_11143,N_10963,N_10816);
nor U11144 (N_11144,N_10924,N_10999);
or U11145 (N_11145,N_10842,N_10962);
and U11146 (N_11146,N_10993,N_10899);
nor U11147 (N_11147,N_10981,N_10852);
nor U11148 (N_11148,N_10942,N_10993);
or U11149 (N_11149,N_10891,N_10941);
nand U11150 (N_11150,N_10885,N_10882);
nand U11151 (N_11151,N_10896,N_10952);
and U11152 (N_11152,N_10948,N_10969);
and U11153 (N_11153,N_10886,N_10973);
xor U11154 (N_11154,N_10896,N_10922);
xor U11155 (N_11155,N_10912,N_10824);
nand U11156 (N_11156,N_10997,N_10929);
or U11157 (N_11157,N_10801,N_10927);
and U11158 (N_11158,N_10862,N_10972);
xnor U11159 (N_11159,N_10867,N_10884);
or U11160 (N_11160,N_10957,N_10928);
nand U11161 (N_11161,N_10854,N_10912);
nor U11162 (N_11162,N_10965,N_10989);
nand U11163 (N_11163,N_10953,N_10871);
xnor U11164 (N_11164,N_10850,N_10806);
or U11165 (N_11165,N_10971,N_10943);
nor U11166 (N_11166,N_10908,N_10920);
xnor U11167 (N_11167,N_10935,N_10940);
or U11168 (N_11168,N_10929,N_10894);
nor U11169 (N_11169,N_10865,N_10922);
and U11170 (N_11170,N_10849,N_10974);
and U11171 (N_11171,N_10962,N_10988);
and U11172 (N_11172,N_10875,N_10990);
or U11173 (N_11173,N_10983,N_10938);
nand U11174 (N_11174,N_10969,N_10988);
nor U11175 (N_11175,N_10986,N_10978);
and U11176 (N_11176,N_10937,N_10979);
nand U11177 (N_11177,N_10933,N_10993);
xor U11178 (N_11178,N_10996,N_10977);
nand U11179 (N_11179,N_10887,N_10885);
nand U11180 (N_11180,N_10897,N_10996);
or U11181 (N_11181,N_10960,N_10912);
xor U11182 (N_11182,N_10935,N_10915);
xor U11183 (N_11183,N_10940,N_10900);
nor U11184 (N_11184,N_10833,N_10936);
nor U11185 (N_11185,N_10809,N_10978);
and U11186 (N_11186,N_10894,N_10941);
or U11187 (N_11187,N_10808,N_10992);
and U11188 (N_11188,N_10836,N_10903);
or U11189 (N_11189,N_10978,N_10933);
nand U11190 (N_11190,N_10858,N_10887);
or U11191 (N_11191,N_10948,N_10852);
and U11192 (N_11192,N_10853,N_10992);
nor U11193 (N_11193,N_10989,N_10908);
or U11194 (N_11194,N_10944,N_10877);
nor U11195 (N_11195,N_10829,N_10975);
or U11196 (N_11196,N_10955,N_10946);
or U11197 (N_11197,N_10844,N_10882);
nor U11198 (N_11198,N_10845,N_10882);
and U11199 (N_11199,N_10929,N_10906);
nor U11200 (N_11200,N_11077,N_11017);
or U11201 (N_11201,N_11071,N_11075);
nor U11202 (N_11202,N_11040,N_11147);
xor U11203 (N_11203,N_11100,N_11192);
xnor U11204 (N_11204,N_11012,N_11102);
or U11205 (N_11205,N_11157,N_11087);
nor U11206 (N_11206,N_11004,N_11171);
or U11207 (N_11207,N_11074,N_11042);
and U11208 (N_11208,N_11043,N_11088);
nand U11209 (N_11209,N_11132,N_11116);
and U11210 (N_11210,N_11140,N_11150);
or U11211 (N_11211,N_11118,N_11011);
nor U11212 (N_11212,N_11014,N_11135);
or U11213 (N_11213,N_11174,N_11162);
or U11214 (N_11214,N_11052,N_11110);
xor U11215 (N_11215,N_11041,N_11024);
or U11216 (N_11216,N_11115,N_11121);
nor U11217 (N_11217,N_11107,N_11096);
and U11218 (N_11218,N_11038,N_11058);
nand U11219 (N_11219,N_11154,N_11032);
xor U11220 (N_11220,N_11081,N_11172);
xor U11221 (N_11221,N_11060,N_11008);
or U11222 (N_11222,N_11046,N_11002);
or U11223 (N_11223,N_11062,N_11120);
nand U11224 (N_11224,N_11184,N_11051);
or U11225 (N_11225,N_11084,N_11175);
xor U11226 (N_11226,N_11159,N_11108);
and U11227 (N_11227,N_11180,N_11007);
and U11228 (N_11228,N_11029,N_11101);
nand U11229 (N_11229,N_11050,N_11057);
nor U11230 (N_11230,N_11182,N_11005);
nand U11231 (N_11231,N_11036,N_11146);
nor U11232 (N_11232,N_11085,N_11161);
nand U11233 (N_11233,N_11009,N_11033);
nand U11234 (N_11234,N_11073,N_11022);
nand U11235 (N_11235,N_11076,N_11148);
xor U11236 (N_11236,N_11056,N_11151);
or U11237 (N_11237,N_11082,N_11191);
nor U11238 (N_11238,N_11186,N_11019);
and U11239 (N_11239,N_11141,N_11138);
xor U11240 (N_11240,N_11093,N_11048);
or U11241 (N_11241,N_11189,N_11124);
and U11242 (N_11242,N_11103,N_11021);
xor U11243 (N_11243,N_11083,N_11168);
and U11244 (N_11244,N_11136,N_11063);
nand U11245 (N_11245,N_11128,N_11176);
or U11246 (N_11246,N_11045,N_11030);
or U11247 (N_11247,N_11034,N_11109);
nor U11248 (N_11248,N_11006,N_11086);
xor U11249 (N_11249,N_11031,N_11064);
xnor U11250 (N_11250,N_11122,N_11078);
nand U11251 (N_11251,N_11027,N_11061);
nand U11252 (N_11252,N_11054,N_11095);
nor U11253 (N_11253,N_11139,N_11163);
or U11254 (N_11254,N_11160,N_11145);
and U11255 (N_11255,N_11142,N_11114);
nand U11256 (N_11256,N_11018,N_11164);
and U11257 (N_11257,N_11090,N_11047);
xor U11258 (N_11258,N_11131,N_11133);
nand U11259 (N_11259,N_11105,N_11013);
nand U11260 (N_11260,N_11067,N_11069);
or U11261 (N_11261,N_11190,N_11039);
nor U11262 (N_11262,N_11188,N_11183);
nand U11263 (N_11263,N_11165,N_11106);
nand U11264 (N_11264,N_11097,N_11185);
and U11265 (N_11265,N_11198,N_11130);
or U11266 (N_11266,N_11049,N_11068);
and U11267 (N_11267,N_11196,N_11003);
xnor U11268 (N_11268,N_11035,N_11127);
xor U11269 (N_11269,N_11079,N_11028);
xor U11270 (N_11270,N_11166,N_11187);
and U11271 (N_11271,N_11153,N_11037);
nor U11272 (N_11272,N_11092,N_11156);
or U11273 (N_11273,N_11179,N_11044);
nand U11274 (N_11274,N_11020,N_11134);
nor U11275 (N_11275,N_11072,N_11113);
or U11276 (N_11276,N_11177,N_11023);
or U11277 (N_11277,N_11091,N_11119);
and U11278 (N_11278,N_11193,N_11066);
xor U11279 (N_11279,N_11111,N_11181);
and U11280 (N_11280,N_11155,N_11152);
nand U11281 (N_11281,N_11089,N_11197);
nor U11282 (N_11282,N_11195,N_11167);
xnor U11283 (N_11283,N_11173,N_11112);
nor U11284 (N_11284,N_11016,N_11123);
or U11285 (N_11285,N_11169,N_11000);
nand U11286 (N_11286,N_11158,N_11001);
nand U11287 (N_11287,N_11055,N_11010);
nand U11288 (N_11288,N_11117,N_11080);
nor U11289 (N_11289,N_11026,N_11094);
or U11290 (N_11290,N_11053,N_11065);
xnor U11291 (N_11291,N_11015,N_11070);
nor U11292 (N_11292,N_11125,N_11144);
nor U11293 (N_11293,N_11199,N_11143);
and U11294 (N_11294,N_11194,N_11098);
or U11295 (N_11295,N_11059,N_11149);
nor U11296 (N_11296,N_11137,N_11170);
xor U11297 (N_11297,N_11025,N_11104);
nor U11298 (N_11298,N_11126,N_11129);
nand U11299 (N_11299,N_11178,N_11099);
xnor U11300 (N_11300,N_11040,N_11001);
nand U11301 (N_11301,N_11072,N_11050);
or U11302 (N_11302,N_11183,N_11111);
xnor U11303 (N_11303,N_11079,N_11047);
or U11304 (N_11304,N_11162,N_11185);
nand U11305 (N_11305,N_11024,N_11178);
nand U11306 (N_11306,N_11062,N_11133);
nand U11307 (N_11307,N_11045,N_11106);
nor U11308 (N_11308,N_11131,N_11083);
nand U11309 (N_11309,N_11064,N_11137);
or U11310 (N_11310,N_11131,N_11119);
xnor U11311 (N_11311,N_11085,N_11078);
xor U11312 (N_11312,N_11067,N_11112);
or U11313 (N_11313,N_11144,N_11011);
nand U11314 (N_11314,N_11070,N_11054);
nand U11315 (N_11315,N_11139,N_11094);
and U11316 (N_11316,N_11002,N_11020);
nand U11317 (N_11317,N_11016,N_11089);
and U11318 (N_11318,N_11017,N_11121);
xor U11319 (N_11319,N_11131,N_11150);
xnor U11320 (N_11320,N_11056,N_11073);
and U11321 (N_11321,N_11122,N_11156);
and U11322 (N_11322,N_11090,N_11178);
or U11323 (N_11323,N_11119,N_11079);
and U11324 (N_11324,N_11081,N_11151);
and U11325 (N_11325,N_11079,N_11091);
xnor U11326 (N_11326,N_11145,N_11192);
nand U11327 (N_11327,N_11189,N_11115);
and U11328 (N_11328,N_11166,N_11188);
nor U11329 (N_11329,N_11031,N_11047);
nor U11330 (N_11330,N_11187,N_11061);
nor U11331 (N_11331,N_11106,N_11056);
or U11332 (N_11332,N_11123,N_11164);
nor U11333 (N_11333,N_11047,N_11088);
nand U11334 (N_11334,N_11170,N_11013);
xor U11335 (N_11335,N_11119,N_11059);
or U11336 (N_11336,N_11078,N_11028);
nor U11337 (N_11337,N_11004,N_11073);
nand U11338 (N_11338,N_11174,N_11199);
nor U11339 (N_11339,N_11071,N_11042);
and U11340 (N_11340,N_11025,N_11086);
nand U11341 (N_11341,N_11040,N_11153);
nand U11342 (N_11342,N_11091,N_11136);
or U11343 (N_11343,N_11118,N_11032);
or U11344 (N_11344,N_11110,N_11054);
nand U11345 (N_11345,N_11153,N_11021);
nor U11346 (N_11346,N_11107,N_11085);
and U11347 (N_11347,N_11046,N_11086);
nor U11348 (N_11348,N_11038,N_11191);
xnor U11349 (N_11349,N_11145,N_11043);
nand U11350 (N_11350,N_11039,N_11196);
or U11351 (N_11351,N_11102,N_11136);
or U11352 (N_11352,N_11169,N_11134);
or U11353 (N_11353,N_11126,N_11074);
xor U11354 (N_11354,N_11172,N_11178);
nand U11355 (N_11355,N_11033,N_11000);
and U11356 (N_11356,N_11198,N_11153);
nand U11357 (N_11357,N_11020,N_11080);
xnor U11358 (N_11358,N_11088,N_11159);
or U11359 (N_11359,N_11046,N_11178);
nand U11360 (N_11360,N_11110,N_11111);
and U11361 (N_11361,N_11136,N_11027);
nand U11362 (N_11362,N_11070,N_11100);
or U11363 (N_11363,N_11168,N_11072);
nand U11364 (N_11364,N_11182,N_11116);
and U11365 (N_11365,N_11188,N_11164);
nor U11366 (N_11366,N_11123,N_11192);
nor U11367 (N_11367,N_11058,N_11165);
or U11368 (N_11368,N_11169,N_11124);
and U11369 (N_11369,N_11116,N_11065);
and U11370 (N_11370,N_11014,N_11116);
nand U11371 (N_11371,N_11153,N_11043);
xor U11372 (N_11372,N_11130,N_11126);
or U11373 (N_11373,N_11125,N_11089);
nand U11374 (N_11374,N_11143,N_11054);
or U11375 (N_11375,N_11100,N_11193);
nor U11376 (N_11376,N_11106,N_11133);
nor U11377 (N_11377,N_11106,N_11178);
and U11378 (N_11378,N_11120,N_11052);
or U11379 (N_11379,N_11170,N_11157);
xnor U11380 (N_11380,N_11053,N_11133);
nor U11381 (N_11381,N_11157,N_11090);
or U11382 (N_11382,N_11145,N_11146);
and U11383 (N_11383,N_11041,N_11039);
and U11384 (N_11384,N_11096,N_11111);
or U11385 (N_11385,N_11114,N_11075);
or U11386 (N_11386,N_11121,N_11185);
xor U11387 (N_11387,N_11026,N_11030);
xor U11388 (N_11388,N_11177,N_11199);
xor U11389 (N_11389,N_11188,N_11179);
and U11390 (N_11390,N_11012,N_11115);
xor U11391 (N_11391,N_11003,N_11159);
and U11392 (N_11392,N_11005,N_11058);
or U11393 (N_11393,N_11060,N_11084);
and U11394 (N_11394,N_11073,N_11172);
xnor U11395 (N_11395,N_11083,N_11097);
nand U11396 (N_11396,N_11072,N_11037);
xor U11397 (N_11397,N_11087,N_11123);
xnor U11398 (N_11398,N_11146,N_11199);
and U11399 (N_11399,N_11184,N_11064);
nand U11400 (N_11400,N_11283,N_11224);
or U11401 (N_11401,N_11211,N_11366);
or U11402 (N_11402,N_11281,N_11206);
and U11403 (N_11403,N_11335,N_11361);
and U11404 (N_11404,N_11337,N_11261);
nand U11405 (N_11405,N_11230,N_11369);
nand U11406 (N_11406,N_11307,N_11324);
and U11407 (N_11407,N_11223,N_11385);
or U11408 (N_11408,N_11250,N_11227);
nand U11409 (N_11409,N_11263,N_11213);
or U11410 (N_11410,N_11380,N_11204);
or U11411 (N_11411,N_11296,N_11387);
nor U11412 (N_11412,N_11269,N_11378);
or U11413 (N_11413,N_11272,N_11254);
xor U11414 (N_11414,N_11236,N_11341);
or U11415 (N_11415,N_11200,N_11332);
nor U11416 (N_11416,N_11388,N_11358);
xor U11417 (N_11417,N_11363,N_11330);
or U11418 (N_11418,N_11339,N_11399);
or U11419 (N_11419,N_11310,N_11379);
nor U11420 (N_11420,N_11329,N_11390);
or U11421 (N_11421,N_11209,N_11267);
and U11422 (N_11422,N_11392,N_11262);
nand U11423 (N_11423,N_11303,N_11221);
nor U11424 (N_11424,N_11359,N_11278);
nand U11425 (N_11425,N_11293,N_11353);
xnor U11426 (N_11426,N_11247,N_11288);
nand U11427 (N_11427,N_11322,N_11289);
nor U11428 (N_11428,N_11285,N_11350);
xor U11429 (N_11429,N_11372,N_11314);
or U11430 (N_11430,N_11316,N_11232);
and U11431 (N_11431,N_11246,N_11234);
or U11432 (N_11432,N_11257,N_11377);
xor U11433 (N_11433,N_11391,N_11349);
nor U11434 (N_11434,N_11321,N_11365);
xnor U11435 (N_11435,N_11238,N_11331);
xnor U11436 (N_11436,N_11344,N_11343);
xor U11437 (N_11437,N_11231,N_11320);
nor U11438 (N_11438,N_11208,N_11277);
and U11439 (N_11439,N_11264,N_11352);
or U11440 (N_11440,N_11276,N_11300);
and U11441 (N_11441,N_11243,N_11371);
nor U11442 (N_11442,N_11367,N_11306);
or U11443 (N_11443,N_11203,N_11241);
or U11444 (N_11444,N_11364,N_11338);
or U11445 (N_11445,N_11218,N_11284);
nor U11446 (N_11446,N_11253,N_11282);
or U11447 (N_11447,N_11291,N_11205);
and U11448 (N_11448,N_11301,N_11327);
and U11449 (N_11449,N_11274,N_11345);
nor U11450 (N_11450,N_11245,N_11389);
xnor U11451 (N_11451,N_11315,N_11299);
xor U11452 (N_11452,N_11356,N_11207);
xnor U11453 (N_11453,N_11355,N_11212);
xnor U11454 (N_11454,N_11382,N_11240);
nand U11455 (N_11455,N_11297,N_11304);
and U11456 (N_11456,N_11248,N_11362);
and U11457 (N_11457,N_11239,N_11268);
nor U11458 (N_11458,N_11279,N_11287);
nand U11459 (N_11459,N_11266,N_11298);
and U11460 (N_11460,N_11309,N_11319);
xnor U11461 (N_11461,N_11244,N_11368);
nand U11462 (N_11462,N_11215,N_11271);
xor U11463 (N_11463,N_11233,N_11202);
nand U11464 (N_11464,N_11383,N_11348);
nor U11465 (N_11465,N_11290,N_11333);
and U11466 (N_11466,N_11351,N_11375);
and U11467 (N_11467,N_11242,N_11210);
nor U11468 (N_11468,N_11313,N_11373);
xor U11469 (N_11469,N_11258,N_11217);
nand U11470 (N_11470,N_11354,N_11325);
and U11471 (N_11471,N_11222,N_11374);
nor U11472 (N_11472,N_11398,N_11219);
nor U11473 (N_11473,N_11286,N_11295);
nand U11474 (N_11474,N_11384,N_11201);
xor U11475 (N_11475,N_11235,N_11357);
and U11476 (N_11476,N_11226,N_11256);
nand U11477 (N_11477,N_11305,N_11347);
nand U11478 (N_11478,N_11381,N_11397);
or U11479 (N_11479,N_11395,N_11249);
xnor U11480 (N_11480,N_11340,N_11370);
xor U11481 (N_11481,N_11334,N_11336);
xor U11482 (N_11482,N_11386,N_11273);
nand U11483 (N_11483,N_11312,N_11216);
xnor U11484 (N_11484,N_11323,N_11259);
nor U11485 (N_11485,N_11228,N_11237);
xor U11486 (N_11486,N_11292,N_11252);
nor U11487 (N_11487,N_11376,N_11396);
nor U11488 (N_11488,N_11393,N_11251);
and U11489 (N_11489,N_11275,N_11326);
or U11490 (N_11490,N_11265,N_11346);
nand U11491 (N_11491,N_11214,N_11311);
or U11492 (N_11492,N_11342,N_11280);
xor U11493 (N_11493,N_11255,N_11328);
nor U11494 (N_11494,N_11360,N_11318);
xor U11495 (N_11495,N_11302,N_11225);
or U11496 (N_11496,N_11394,N_11317);
and U11497 (N_11497,N_11308,N_11270);
and U11498 (N_11498,N_11229,N_11260);
nand U11499 (N_11499,N_11294,N_11220);
nand U11500 (N_11500,N_11229,N_11251);
and U11501 (N_11501,N_11350,N_11203);
nor U11502 (N_11502,N_11312,N_11345);
nor U11503 (N_11503,N_11318,N_11328);
nand U11504 (N_11504,N_11310,N_11264);
nor U11505 (N_11505,N_11339,N_11363);
and U11506 (N_11506,N_11368,N_11332);
xnor U11507 (N_11507,N_11359,N_11293);
and U11508 (N_11508,N_11236,N_11310);
xor U11509 (N_11509,N_11208,N_11370);
nand U11510 (N_11510,N_11313,N_11323);
nor U11511 (N_11511,N_11231,N_11333);
nand U11512 (N_11512,N_11302,N_11397);
nor U11513 (N_11513,N_11394,N_11298);
nand U11514 (N_11514,N_11271,N_11217);
xor U11515 (N_11515,N_11398,N_11259);
xnor U11516 (N_11516,N_11234,N_11204);
nand U11517 (N_11517,N_11254,N_11219);
nand U11518 (N_11518,N_11376,N_11321);
nand U11519 (N_11519,N_11357,N_11344);
nand U11520 (N_11520,N_11376,N_11245);
nand U11521 (N_11521,N_11342,N_11238);
nor U11522 (N_11522,N_11306,N_11387);
or U11523 (N_11523,N_11314,N_11339);
nor U11524 (N_11524,N_11317,N_11230);
xnor U11525 (N_11525,N_11359,N_11259);
nor U11526 (N_11526,N_11344,N_11354);
or U11527 (N_11527,N_11274,N_11206);
xnor U11528 (N_11528,N_11283,N_11271);
xor U11529 (N_11529,N_11237,N_11267);
or U11530 (N_11530,N_11237,N_11219);
or U11531 (N_11531,N_11365,N_11266);
and U11532 (N_11532,N_11284,N_11262);
and U11533 (N_11533,N_11379,N_11339);
nand U11534 (N_11534,N_11210,N_11232);
and U11535 (N_11535,N_11384,N_11302);
xor U11536 (N_11536,N_11381,N_11340);
or U11537 (N_11537,N_11257,N_11201);
nor U11538 (N_11538,N_11386,N_11224);
nor U11539 (N_11539,N_11331,N_11360);
nor U11540 (N_11540,N_11378,N_11351);
xnor U11541 (N_11541,N_11236,N_11354);
nor U11542 (N_11542,N_11295,N_11208);
nor U11543 (N_11543,N_11307,N_11238);
or U11544 (N_11544,N_11313,N_11240);
and U11545 (N_11545,N_11347,N_11329);
xor U11546 (N_11546,N_11311,N_11273);
xnor U11547 (N_11547,N_11368,N_11366);
and U11548 (N_11548,N_11257,N_11209);
nor U11549 (N_11549,N_11246,N_11382);
nor U11550 (N_11550,N_11209,N_11376);
or U11551 (N_11551,N_11244,N_11344);
nor U11552 (N_11552,N_11335,N_11233);
xnor U11553 (N_11553,N_11207,N_11292);
nor U11554 (N_11554,N_11383,N_11375);
xor U11555 (N_11555,N_11281,N_11364);
or U11556 (N_11556,N_11354,N_11326);
nor U11557 (N_11557,N_11265,N_11395);
nand U11558 (N_11558,N_11308,N_11326);
nand U11559 (N_11559,N_11364,N_11319);
nand U11560 (N_11560,N_11334,N_11262);
nor U11561 (N_11561,N_11329,N_11353);
xnor U11562 (N_11562,N_11273,N_11290);
nand U11563 (N_11563,N_11214,N_11376);
or U11564 (N_11564,N_11394,N_11249);
xnor U11565 (N_11565,N_11335,N_11268);
nand U11566 (N_11566,N_11232,N_11366);
nand U11567 (N_11567,N_11344,N_11330);
or U11568 (N_11568,N_11220,N_11203);
nor U11569 (N_11569,N_11240,N_11307);
nand U11570 (N_11570,N_11382,N_11363);
or U11571 (N_11571,N_11382,N_11356);
nor U11572 (N_11572,N_11371,N_11396);
nand U11573 (N_11573,N_11292,N_11389);
nand U11574 (N_11574,N_11314,N_11236);
nor U11575 (N_11575,N_11255,N_11340);
nor U11576 (N_11576,N_11314,N_11233);
or U11577 (N_11577,N_11314,N_11227);
nand U11578 (N_11578,N_11313,N_11220);
nor U11579 (N_11579,N_11216,N_11241);
nand U11580 (N_11580,N_11381,N_11290);
xnor U11581 (N_11581,N_11370,N_11312);
nand U11582 (N_11582,N_11303,N_11208);
xnor U11583 (N_11583,N_11323,N_11350);
nor U11584 (N_11584,N_11391,N_11370);
nor U11585 (N_11585,N_11263,N_11233);
xnor U11586 (N_11586,N_11395,N_11300);
nor U11587 (N_11587,N_11359,N_11343);
nand U11588 (N_11588,N_11367,N_11201);
or U11589 (N_11589,N_11364,N_11268);
xor U11590 (N_11590,N_11360,N_11342);
xnor U11591 (N_11591,N_11259,N_11279);
and U11592 (N_11592,N_11321,N_11231);
and U11593 (N_11593,N_11353,N_11295);
nand U11594 (N_11594,N_11291,N_11288);
and U11595 (N_11595,N_11385,N_11218);
or U11596 (N_11596,N_11267,N_11240);
xnor U11597 (N_11597,N_11341,N_11261);
xor U11598 (N_11598,N_11273,N_11285);
or U11599 (N_11599,N_11250,N_11390);
or U11600 (N_11600,N_11486,N_11452);
and U11601 (N_11601,N_11525,N_11589);
or U11602 (N_11602,N_11503,N_11562);
or U11603 (N_11603,N_11456,N_11464);
and U11604 (N_11604,N_11553,N_11442);
xnor U11605 (N_11605,N_11565,N_11413);
and U11606 (N_11606,N_11404,N_11446);
nand U11607 (N_11607,N_11536,N_11508);
nor U11608 (N_11608,N_11491,N_11585);
nor U11609 (N_11609,N_11535,N_11477);
or U11610 (N_11610,N_11445,N_11559);
nor U11611 (N_11611,N_11515,N_11432);
xnor U11612 (N_11612,N_11526,N_11557);
and U11613 (N_11613,N_11566,N_11554);
and U11614 (N_11614,N_11469,N_11529);
xor U11615 (N_11615,N_11523,N_11483);
xor U11616 (N_11616,N_11592,N_11509);
xnor U11617 (N_11617,N_11465,N_11517);
xnor U11618 (N_11618,N_11499,N_11466);
xnor U11619 (N_11619,N_11593,N_11458);
nand U11620 (N_11620,N_11484,N_11474);
xnor U11621 (N_11621,N_11551,N_11583);
nor U11622 (N_11622,N_11549,N_11462);
and U11623 (N_11623,N_11463,N_11577);
nor U11624 (N_11624,N_11560,N_11485);
or U11625 (N_11625,N_11473,N_11480);
and U11626 (N_11626,N_11451,N_11527);
nor U11627 (N_11627,N_11421,N_11402);
nor U11628 (N_11628,N_11435,N_11438);
xor U11629 (N_11629,N_11496,N_11580);
xnor U11630 (N_11630,N_11406,N_11574);
nor U11631 (N_11631,N_11428,N_11423);
or U11632 (N_11632,N_11403,N_11455);
and U11633 (N_11633,N_11556,N_11471);
or U11634 (N_11634,N_11461,N_11595);
nor U11635 (N_11635,N_11498,N_11575);
nor U11636 (N_11636,N_11460,N_11411);
and U11637 (N_11637,N_11573,N_11495);
or U11638 (N_11638,N_11558,N_11489);
nor U11639 (N_11639,N_11487,N_11599);
or U11640 (N_11640,N_11530,N_11409);
and U11641 (N_11641,N_11405,N_11548);
xnor U11642 (N_11642,N_11518,N_11492);
and U11643 (N_11643,N_11490,N_11581);
or U11644 (N_11644,N_11436,N_11415);
nor U11645 (N_11645,N_11454,N_11570);
nor U11646 (N_11646,N_11520,N_11513);
xor U11647 (N_11647,N_11430,N_11497);
and U11648 (N_11648,N_11552,N_11475);
nand U11649 (N_11649,N_11453,N_11420);
nand U11650 (N_11650,N_11450,N_11433);
xnor U11651 (N_11651,N_11537,N_11576);
xor U11652 (N_11652,N_11561,N_11505);
or U11653 (N_11653,N_11419,N_11596);
and U11654 (N_11654,N_11534,N_11544);
nor U11655 (N_11655,N_11532,N_11510);
or U11656 (N_11656,N_11417,N_11571);
nand U11657 (N_11657,N_11400,N_11493);
or U11658 (N_11658,N_11516,N_11564);
and U11659 (N_11659,N_11441,N_11478);
nand U11660 (N_11660,N_11457,N_11448);
nand U11661 (N_11661,N_11504,N_11408);
or U11662 (N_11662,N_11541,N_11437);
xnor U11663 (N_11663,N_11476,N_11422);
or U11664 (N_11664,N_11439,N_11587);
nand U11665 (N_11665,N_11590,N_11514);
nand U11666 (N_11666,N_11588,N_11444);
and U11667 (N_11667,N_11414,N_11598);
or U11668 (N_11668,N_11443,N_11416);
nor U11669 (N_11669,N_11494,N_11550);
and U11670 (N_11670,N_11568,N_11540);
nand U11671 (N_11671,N_11426,N_11528);
and U11672 (N_11672,N_11427,N_11470);
and U11673 (N_11673,N_11538,N_11511);
nand U11674 (N_11674,N_11500,N_11524);
and U11675 (N_11675,N_11545,N_11449);
nor U11676 (N_11676,N_11563,N_11488);
xor U11677 (N_11677,N_11542,N_11582);
nor U11678 (N_11678,N_11440,N_11539);
nand U11679 (N_11679,N_11555,N_11410);
nand U11680 (N_11680,N_11591,N_11401);
xor U11681 (N_11681,N_11481,N_11407);
xor U11682 (N_11682,N_11579,N_11418);
nor U11683 (N_11683,N_11546,N_11521);
or U11684 (N_11684,N_11425,N_11412);
nand U11685 (N_11685,N_11522,N_11472);
xor U11686 (N_11686,N_11431,N_11482);
and U11687 (N_11687,N_11429,N_11447);
and U11688 (N_11688,N_11468,N_11594);
nor U11689 (N_11689,N_11434,N_11467);
nand U11690 (N_11690,N_11501,N_11597);
or U11691 (N_11691,N_11507,N_11584);
xor U11692 (N_11692,N_11547,N_11586);
or U11693 (N_11693,N_11479,N_11572);
and U11694 (N_11694,N_11506,N_11459);
nand U11695 (N_11695,N_11519,N_11502);
nand U11696 (N_11696,N_11543,N_11531);
nor U11697 (N_11697,N_11424,N_11578);
nor U11698 (N_11698,N_11533,N_11567);
xnor U11699 (N_11699,N_11512,N_11569);
or U11700 (N_11700,N_11455,N_11423);
or U11701 (N_11701,N_11410,N_11444);
nor U11702 (N_11702,N_11571,N_11495);
nand U11703 (N_11703,N_11500,N_11468);
xor U11704 (N_11704,N_11520,N_11411);
and U11705 (N_11705,N_11452,N_11400);
and U11706 (N_11706,N_11465,N_11547);
or U11707 (N_11707,N_11599,N_11432);
xnor U11708 (N_11708,N_11442,N_11593);
and U11709 (N_11709,N_11569,N_11408);
nand U11710 (N_11710,N_11508,N_11557);
or U11711 (N_11711,N_11479,N_11499);
or U11712 (N_11712,N_11418,N_11416);
or U11713 (N_11713,N_11468,N_11510);
xnor U11714 (N_11714,N_11594,N_11438);
nor U11715 (N_11715,N_11492,N_11472);
or U11716 (N_11716,N_11409,N_11441);
and U11717 (N_11717,N_11441,N_11496);
or U11718 (N_11718,N_11492,N_11551);
xnor U11719 (N_11719,N_11428,N_11518);
and U11720 (N_11720,N_11412,N_11485);
and U11721 (N_11721,N_11528,N_11524);
and U11722 (N_11722,N_11523,N_11591);
xor U11723 (N_11723,N_11598,N_11463);
nand U11724 (N_11724,N_11448,N_11429);
nor U11725 (N_11725,N_11448,N_11581);
nand U11726 (N_11726,N_11431,N_11450);
nor U11727 (N_11727,N_11566,N_11505);
xnor U11728 (N_11728,N_11423,N_11403);
nor U11729 (N_11729,N_11515,N_11464);
and U11730 (N_11730,N_11423,N_11559);
or U11731 (N_11731,N_11565,N_11453);
and U11732 (N_11732,N_11551,N_11518);
and U11733 (N_11733,N_11550,N_11515);
or U11734 (N_11734,N_11420,N_11562);
or U11735 (N_11735,N_11439,N_11515);
nor U11736 (N_11736,N_11499,N_11500);
or U11737 (N_11737,N_11422,N_11415);
xnor U11738 (N_11738,N_11487,N_11581);
nor U11739 (N_11739,N_11495,N_11488);
and U11740 (N_11740,N_11572,N_11594);
nand U11741 (N_11741,N_11474,N_11557);
nand U11742 (N_11742,N_11492,N_11437);
nand U11743 (N_11743,N_11493,N_11473);
nand U11744 (N_11744,N_11471,N_11587);
xor U11745 (N_11745,N_11437,N_11408);
nand U11746 (N_11746,N_11525,N_11535);
nand U11747 (N_11747,N_11434,N_11448);
nor U11748 (N_11748,N_11510,N_11450);
xnor U11749 (N_11749,N_11537,N_11521);
and U11750 (N_11750,N_11402,N_11586);
nand U11751 (N_11751,N_11563,N_11484);
nor U11752 (N_11752,N_11436,N_11525);
and U11753 (N_11753,N_11433,N_11423);
nor U11754 (N_11754,N_11571,N_11400);
xnor U11755 (N_11755,N_11462,N_11491);
xor U11756 (N_11756,N_11481,N_11482);
nand U11757 (N_11757,N_11576,N_11517);
nand U11758 (N_11758,N_11412,N_11446);
nand U11759 (N_11759,N_11508,N_11516);
nand U11760 (N_11760,N_11481,N_11444);
xnor U11761 (N_11761,N_11559,N_11587);
nand U11762 (N_11762,N_11465,N_11482);
nor U11763 (N_11763,N_11409,N_11453);
nand U11764 (N_11764,N_11469,N_11537);
and U11765 (N_11765,N_11405,N_11528);
and U11766 (N_11766,N_11448,N_11404);
nor U11767 (N_11767,N_11455,N_11524);
nor U11768 (N_11768,N_11570,N_11485);
nand U11769 (N_11769,N_11594,N_11578);
nand U11770 (N_11770,N_11531,N_11432);
nand U11771 (N_11771,N_11528,N_11566);
and U11772 (N_11772,N_11591,N_11431);
nor U11773 (N_11773,N_11589,N_11541);
and U11774 (N_11774,N_11407,N_11410);
xnor U11775 (N_11775,N_11581,N_11497);
xor U11776 (N_11776,N_11565,N_11592);
nor U11777 (N_11777,N_11582,N_11497);
nand U11778 (N_11778,N_11562,N_11536);
xnor U11779 (N_11779,N_11587,N_11413);
or U11780 (N_11780,N_11495,N_11504);
or U11781 (N_11781,N_11407,N_11510);
and U11782 (N_11782,N_11434,N_11592);
nor U11783 (N_11783,N_11422,N_11506);
or U11784 (N_11784,N_11423,N_11421);
nand U11785 (N_11785,N_11408,N_11537);
xnor U11786 (N_11786,N_11547,N_11596);
and U11787 (N_11787,N_11428,N_11521);
and U11788 (N_11788,N_11422,N_11461);
nor U11789 (N_11789,N_11503,N_11505);
xnor U11790 (N_11790,N_11455,N_11486);
or U11791 (N_11791,N_11524,N_11503);
and U11792 (N_11792,N_11450,N_11439);
nand U11793 (N_11793,N_11538,N_11499);
nor U11794 (N_11794,N_11542,N_11455);
nor U11795 (N_11795,N_11550,N_11549);
xor U11796 (N_11796,N_11530,N_11440);
nor U11797 (N_11797,N_11570,N_11541);
or U11798 (N_11798,N_11464,N_11586);
nand U11799 (N_11799,N_11529,N_11563);
xnor U11800 (N_11800,N_11710,N_11702);
nand U11801 (N_11801,N_11632,N_11665);
or U11802 (N_11802,N_11703,N_11749);
xnor U11803 (N_11803,N_11671,N_11706);
and U11804 (N_11804,N_11789,N_11691);
xnor U11805 (N_11805,N_11794,N_11745);
nor U11806 (N_11806,N_11782,N_11799);
or U11807 (N_11807,N_11644,N_11692);
or U11808 (N_11808,N_11660,N_11781);
or U11809 (N_11809,N_11733,N_11776);
and U11810 (N_11810,N_11750,N_11677);
nor U11811 (N_11811,N_11653,N_11721);
nand U11812 (N_11812,N_11662,N_11641);
nor U11813 (N_11813,N_11747,N_11615);
or U11814 (N_11814,N_11609,N_11622);
or U11815 (N_11815,N_11725,N_11766);
xor U11816 (N_11816,N_11613,N_11631);
and U11817 (N_11817,N_11650,N_11748);
and U11818 (N_11818,N_11707,N_11648);
nor U11819 (N_11819,N_11605,N_11759);
nor U11820 (N_11820,N_11611,N_11729);
and U11821 (N_11821,N_11723,N_11656);
or U11822 (N_11822,N_11731,N_11639);
and U11823 (N_11823,N_11674,N_11714);
and U11824 (N_11824,N_11764,N_11682);
or U11825 (N_11825,N_11786,N_11783);
nor U11826 (N_11826,N_11607,N_11798);
nor U11827 (N_11827,N_11755,N_11791);
or U11828 (N_11828,N_11771,N_11664);
or U11829 (N_11829,N_11685,N_11636);
or U11830 (N_11830,N_11777,N_11601);
nand U11831 (N_11831,N_11753,N_11772);
xor U11832 (N_11832,N_11673,N_11757);
and U11833 (N_11833,N_11732,N_11667);
nor U11834 (N_11834,N_11630,N_11688);
or U11835 (N_11835,N_11720,N_11627);
nand U11836 (N_11836,N_11762,N_11704);
xor U11837 (N_11837,N_11687,N_11659);
nand U11838 (N_11838,N_11719,N_11694);
or U11839 (N_11839,N_11634,N_11790);
and U11840 (N_11840,N_11726,N_11724);
nor U11841 (N_11841,N_11796,N_11779);
nand U11842 (N_11842,N_11713,N_11633);
nand U11843 (N_11843,N_11684,N_11795);
nand U11844 (N_11844,N_11763,N_11666);
or U11845 (N_11845,N_11775,N_11623);
nand U11846 (N_11846,N_11708,N_11770);
nor U11847 (N_11847,N_11744,N_11649);
nor U11848 (N_11848,N_11696,N_11742);
xor U11849 (N_11849,N_11716,N_11681);
nor U11850 (N_11850,N_11785,N_11758);
and U11851 (N_11851,N_11661,N_11701);
and U11852 (N_11852,N_11608,N_11709);
nand U11853 (N_11853,N_11743,N_11668);
or U11854 (N_11854,N_11693,N_11651);
nand U11855 (N_11855,N_11752,N_11730);
or U11856 (N_11856,N_11655,N_11679);
nor U11857 (N_11857,N_11676,N_11715);
xor U11858 (N_11858,N_11618,N_11635);
nor U11859 (N_11859,N_11740,N_11722);
or U11860 (N_11860,N_11683,N_11699);
nor U11861 (N_11861,N_11700,N_11769);
nand U11862 (N_11862,N_11695,N_11640);
xor U11863 (N_11863,N_11625,N_11784);
xnor U11864 (N_11864,N_11689,N_11738);
xor U11865 (N_11865,N_11626,N_11670);
and U11866 (N_11866,N_11754,N_11654);
nor U11867 (N_11867,N_11767,N_11765);
nor U11868 (N_11868,N_11669,N_11619);
and U11869 (N_11869,N_11672,N_11734);
nor U11870 (N_11870,N_11658,N_11652);
nand U11871 (N_11871,N_11774,N_11739);
xor U11872 (N_11872,N_11768,N_11761);
nand U11873 (N_11873,N_11647,N_11737);
nor U11874 (N_11874,N_11604,N_11600);
or U11875 (N_11875,N_11788,N_11690);
xnor U11876 (N_11876,N_11705,N_11686);
or U11877 (N_11877,N_11680,N_11675);
nor U11878 (N_11878,N_11746,N_11621);
and U11879 (N_11879,N_11778,N_11780);
xor U11880 (N_11880,N_11638,N_11663);
nand U11881 (N_11881,N_11606,N_11751);
nor U11882 (N_11882,N_11741,N_11678);
or U11883 (N_11883,N_11612,N_11712);
nor U11884 (N_11884,N_11717,N_11620);
and U11885 (N_11885,N_11616,N_11711);
xor U11886 (N_11886,N_11792,N_11787);
and U11887 (N_11887,N_11793,N_11642);
nand U11888 (N_11888,N_11645,N_11617);
or U11889 (N_11889,N_11728,N_11643);
xor U11890 (N_11890,N_11697,N_11614);
xor U11891 (N_11891,N_11698,N_11610);
xnor U11892 (N_11892,N_11624,N_11735);
or U11893 (N_11893,N_11628,N_11646);
or U11894 (N_11894,N_11773,N_11756);
xor U11895 (N_11895,N_11657,N_11736);
nor U11896 (N_11896,N_11797,N_11637);
and U11897 (N_11897,N_11602,N_11603);
nand U11898 (N_11898,N_11760,N_11727);
or U11899 (N_11899,N_11718,N_11629);
or U11900 (N_11900,N_11748,N_11638);
nor U11901 (N_11901,N_11717,N_11785);
xor U11902 (N_11902,N_11624,N_11601);
or U11903 (N_11903,N_11737,N_11761);
nor U11904 (N_11904,N_11636,N_11610);
and U11905 (N_11905,N_11761,N_11727);
and U11906 (N_11906,N_11725,N_11701);
nor U11907 (N_11907,N_11735,N_11614);
nand U11908 (N_11908,N_11754,N_11744);
xor U11909 (N_11909,N_11790,N_11678);
nor U11910 (N_11910,N_11709,N_11796);
xor U11911 (N_11911,N_11676,N_11777);
nor U11912 (N_11912,N_11798,N_11688);
nor U11913 (N_11913,N_11715,N_11798);
or U11914 (N_11914,N_11703,N_11638);
xor U11915 (N_11915,N_11674,N_11745);
and U11916 (N_11916,N_11682,N_11643);
or U11917 (N_11917,N_11712,N_11785);
and U11918 (N_11918,N_11619,N_11739);
xnor U11919 (N_11919,N_11679,N_11739);
nand U11920 (N_11920,N_11618,N_11782);
or U11921 (N_11921,N_11622,N_11761);
or U11922 (N_11922,N_11783,N_11757);
nand U11923 (N_11923,N_11690,N_11714);
or U11924 (N_11924,N_11752,N_11693);
and U11925 (N_11925,N_11753,N_11696);
nand U11926 (N_11926,N_11703,N_11620);
xnor U11927 (N_11927,N_11759,N_11671);
and U11928 (N_11928,N_11736,N_11785);
nor U11929 (N_11929,N_11797,N_11654);
nor U11930 (N_11930,N_11622,N_11769);
or U11931 (N_11931,N_11695,N_11691);
or U11932 (N_11932,N_11716,N_11684);
nand U11933 (N_11933,N_11617,N_11708);
or U11934 (N_11934,N_11608,N_11653);
xor U11935 (N_11935,N_11706,N_11697);
xor U11936 (N_11936,N_11679,N_11735);
xnor U11937 (N_11937,N_11641,N_11789);
nor U11938 (N_11938,N_11721,N_11608);
nand U11939 (N_11939,N_11749,N_11730);
and U11940 (N_11940,N_11658,N_11790);
nand U11941 (N_11941,N_11636,N_11698);
and U11942 (N_11942,N_11649,N_11747);
and U11943 (N_11943,N_11726,N_11693);
xor U11944 (N_11944,N_11717,N_11673);
or U11945 (N_11945,N_11730,N_11664);
or U11946 (N_11946,N_11649,N_11757);
xnor U11947 (N_11947,N_11795,N_11787);
xor U11948 (N_11948,N_11658,N_11630);
nand U11949 (N_11949,N_11631,N_11764);
and U11950 (N_11950,N_11676,N_11668);
xor U11951 (N_11951,N_11714,N_11788);
and U11952 (N_11952,N_11684,N_11660);
xnor U11953 (N_11953,N_11773,N_11693);
xnor U11954 (N_11954,N_11629,N_11712);
nor U11955 (N_11955,N_11608,N_11752);
and U11956 (N_11956,N_11681,N_11668);
xor U11957 (N_11957,N_11741,N_11731);
nor U11958 (N_11958,N_11783,N_11715);
xnor U11959 (N_11959,N_11612,N_11774);
and U11960 (N_11960,N_11650,N_11637);
xor U11961 (N_11961,N_11626,N_11777);
or U11962 (N_11962,N_11678,N_11739);
nand U11963 (N_11963,N_11798,N_11728);
nor U11964 (N_11964,N_11724,N_11686);
and U11965 (N_11965,N_11704,N_11622);
and U11966 (N_11966,N_11778,N_11747);
nor U11967 (N_11967,N_11657,N_11792);
nor U11968 (N_11968,N_11773,N_11683);
nand U11969 (N_11969,N_11754,N_11711);
nor U11970 (N_11970,N_11705,N_11791);
nand U11971 (N_11971,N_11686,N_11629);
nand U11972 (N_11972,N_11791,N_11635);
or U11973 (N_11973,N_11788,N_11711);
xor U11974 (N_11974,N_11635,N_11718);
nand U11975 (N_11975,N_11703,N_11760);
and U11976 (N_11976,N_11757,N_11660);
and U11977 (N_11977,N_11732,N_11797);
nand U11978 (N_11978,N_11760,N_11796);
nor U11979 (N_11979,N_11765,N_11697);
and U11980 (N_11980,N_11741,N_11632);
xor U11981 (N_11981,N_11651,N_11650);
nand U11982 (N_11982,N_11761,N_11641);
or U11983 (N_11983,N_11682,N_11705);
nor U11984 (N_11984,N_11680,N_11753);
and U11985 (N_11985,N_11722,N_11798);
and U11986 (N_11986,N_11739,N_11715);
xnor U11987 (N_11987,N_11713,N_11784);
and U11988 (N_11988,N_11620,N_11624);
xnor U11989 (N_11989,N_11657,N_11711);
nand U11990 (N_11990,N_11665,N_11608);
or U11991 (N_11991,N_11618,N_11644);
nand U11992 (N_11992,N_11749,N_11676);
or U11993 (N_11993,N_11710,N_11662);
or U11994 (N_11994,N_11656,N_11761);
nor U11995 (N_11995,N_11707,N_11617);
or U11996 (N_11996,N_11713,N_11708);
nand U11997 (N_11997,N_11634,N_11793);
nor U11998 (N_11998,N_11663,N_11797);
nand U11999 (N_11999,N_11691,N_11672);
xnor U12000 (N_12000,N_11948,N_11908);
xor U12001 (N_12001,N_11821,N_11828);
xnor U12002 (N_12002,N_11843,N_11886);
xor U12003 (N_12003,N_11909,N_11862);
nand U12004 (N_12004,N_11856,N_11876);
or U12005 (N_12005,N_11981,N_11975);
nor U12006 (N_12006,N_11953,N_11854);
nand U12007 (N_12007,N_11928,N_11964);
xor U12008 (N_12008,N_11824,N_11873);
and U12009 (N_12009,N_11939,N_11874);
nand U12010 (N_12010,N_11883,N_11809);
nor U12011 (N_12011,N_11857,N_11802);
nand U12012 (N_12012,N_11890,N_11838);
xnor U12013 (N_12013,N_11916,N_11870);
xnor U12014 (N_12014,N_11852,N_11917);
nand U12015 (N_12015,N_11910,N_11967);
nand U12016 (N_12016,N_11897,N_11957);
xor U12017 (N_12017,N_11947,N_11952);
xnor U12018 (N_12018,N_11884,N_11973);
and U12019 (N_12019,N_11819,N_11926);
nand U12020 (N_12020,N_11989,N_11920);
or U12021 (N_12021,N_11905,N_11841);
nand U12022 (N_12022,N_11823,N_11921);
or U12023 (N_12023,N_11861,N_11960);
nand U12024 (N_12024,N_11913,N_11895);
and U12025 (N_12025,N_11946,N_11842);
and U12026 (N_12026,N_11945,N_11914);
and U12027 (N_12027,N_11922,N_11980);
xor U12028 (N_12028,N_11845,N_11814);
nand U12029 (N_12029,N_11924,N_11871);
xor U12030 (N_12030,N_11984,N_11912);
or U12031 (N_12031,N_11877,N_11974);
nand U12032 (N_12032,N_11805,N_11806);
xor U12033 (N_12033,N_11990,N_11878);
and U12034 (N_12034,N_11970,N_11961);
nand U12035 (N_12035,N_11995,N_11977);
xor U12036 (N_12036,N_11804,N_11847);
xor U12037 (N_12037,N_11919,N_11860);
or U12038 (N_12038,N_11801,N_11903);
and U12039 (N_12039,N_11839,N_11867);
nand U12040 (N_12040,N_11971,N_11896);
or U12041 (N_12041,N_11965,N_11993);
nand U12042 (N_12042,N_11998,N_11994);
or U12043 (N_12043,N_11837,N_11825);
or U12044 (N_12044,N_11866,N_11858);
nand U12045 (N_12045,N_11979,N_11817);
nor U12046 (N_12046,N_11968,N_11830);
xnor U12047 (N_12047,N_11863,N_11906);
nor U12048 (N_12048,N_11935,N_11832);
and U12049 (N_12049,N_11963,N_11931);
and U12050 (N_12050,N_11966,N_11879);
or U12051 (N_12051,N_11950,N_11959);
and U12052 (N_12052,N_11923,N_11986);
nand U12053 (N_12053,N_11869,N_11846);
nand U12054 (N_12054,N_11851,N_11985);
and U12055 (N_12055,N_11996,N_11956);
nor U12056 (N_12056,N_11958,N_11900);
and U12057 (N_12057,N_11891,N_11901);
nand U12058 (N_12058,N_11987,N_11816);
or U12059 (N_12059,N_11999,N_11898);
nor U12060 (N_12060,N_11872,N_11937);
or U12061 (N_12061,N_11976,N_11833);
nor U12062 (N_12062,N_11962,N_11943);
and U12063 (N_12063,N_11865,N_11818);
xor U12064 (N_12064,N_11829,N_11992);
or U12065 (N_12065,N_11855,N_11954);
nor U12066 (N_12066,N_11822,N_11949);
xor U12067 (N_12067,N_11930,N_11820);
and U12068 (N_12068,N_11812,N_11978);
nor U12069 (N_12069,N_11835,N_11881);
nor U12070 (N_12070,N_11885,N_11827);
or U12071 (N_12071,N_11936,N_11888);
nand U12072 (N_12072,N_11868,N_11887);
or U12073 (N_12073,N_11918,N_11982);
or U12074 (N_12074,N_11848,N_11907);
xor U12075 (N_12075,N_11929,N_11859);
nor U12076 (N_12076,N_11988,N_11875);
nor U12077 (N_12077,N_11836,N_11997);
or U12078 (N_12078,N_11813,N_11850);
and U12079 (N_12079,N_11934,N_11944);
xor U12080 (N_12080,N_11800,N_11902);
or U12081 (N_12081,N_11882,N_11826);
and U12082 (N_12082,N_11938,N_11940);
xnor U12083 (N_12083,N_11941,N_11810);
and U12084 (N_12084,N_11894,N_11972);
nand U12085 (N_12085,N_11899,N_11925);
or U12086 (N_12086,N_11991,N_11849);
nor U12087 (N_12087,N_11933,N_11892);
nand U12088 (N_12088,N_11955,N_11911);
or U12089 (N_12089,N_11969,N_11904);
nor U12090 (N_12090,N_11932,N_11803);
or U12091 (N_12091,N_11915,N_11880);
xor U12092 (N_12092,N_11942,N_11864);
xor U12093 (N_12093,N_11831,N_11808);
nand U12094 (N_12094,N_11853,N_11811);
or U12095 (N_12095,N_11889,N_11844);
nand U12096 (N_12096,N_11983,N_11815);
or U12097 (N_12097,N_11893,N_11951);
nand U12098 (N_12098,N_11834,N_11807);
xnor U12099 (N_12099,N_11927,N_11840);
and U12100 (N_12100,N_11912,N_11888);
nor U12101 (N_12101,N_11887,N_11946);
nor U12102 (N_12102,N_11894,N_11866);
nand U12103 (N_12103,N_11956,N_11987);
nor U12104 (N_12104,N_11901,N_11908);
xor U12105 (N_12105,N_11854,N_11805);
nand U12106 (N_12106,N_11861,N_11826);
and U12107 (N_12107,N_11819,N_11905);
xor U12108 (N_12108,N_11899,N_11801);
nand U12109 (N_12109,N_11854,N_11913);
nand U12110 (N_12110,N_11852,N_11993);
and U12111 (N_12111,N_11900,N_11944);
xor U12112 (N_12112,N_11923,N_11870);
nor U12113 (N_12113,N_11865,N_11835);
nor U12114 (N_12114,N_11800,N_11972);
xnor U12115 (N_12115,N_11897,N_11898);
nor U12116 (N_12116,N_11929,N_11943);
nor U12117 (N_12117,N_11987,N_11979);
or U12118 (N_12118,N_11883,N_11869);
and U12119 (N_12119,N_11975,N_11952);
nand U12120 (N_12120,N_11897,N_11943);
or U12121 (N_12121,N_11804,N_11976);
and U12122 (N_12122,N_11831,N_11864);
or U12123 (N_12123,N_11996,N_11820);
nor U12124 (N_12124,N_11809,N_11970);
and U12125 (N_12125,N_11945,N_11985);
nand U12126 (N_12126,N_11831,N_11836);
nor U12127 (N_12127,N_11808,N_11800);
and U12128 (N_12128,N_11816,N_11812);
and U12129 (N_12129,N_11919,N_11924);
xor U12130 (N_12130,N_11970,N_11872);
or U12131 (N_12131,N_11918,N_11949);
and U12132 (N_12132,N_11883,N_11889);
nand U12133 (N_12133,N_11981,N_11983);
nand U12134 (N_12134,N_11852,N_11846);
nor U12135 (N_12135,N_11903,N_11847);
or U12136 (N_12136,N_11922,N_11828);
or U12137 (N_12137,N_11980,N_11873);
xor U12138 (N_12138,N_11970,N_11888);
xor U12139 (N_12139,N_11840,N_11888);
nor U12140 (N_12140,N_11927,N_11866);
nand U12141 (N_12141,N_11960,N_11865);
nor U12142 (N_12142,N_11837,N_11899);
xor U12143 (N_12143,N_11913,N_11847);
nand U12144 (N_12144,N_11850,N_11879);
xnor U12145 (N_12145,N_11987,N_11933);
or U12146 (N_12146,N_11984,N_11903);
nor U12147 (N_12147,N_11952,N_11936);
nand U12148 (N_12148,N_11924,N_11934);
nor U12149 (N_12149,N_11936,N_11978);
xor U12150 (N_12150,N_11815,N_11852);
and U12151 (N_12151,N_11890,N_11808);
nand U12152 (N_12152,N_11956,N_11935);
nand U12153 (N_12153,N_11844,N_11981);
and U12154 (N_12154,N_11918,N_11896);
nor U12155 (N_12155,N_11956,N_11818);
nand U12156 (N_12156,N_11833,N_11920);
or U12157 (N_12157,N_11802,N_11821);
and U12158 (N_12158,N_11844,N_11983);
and U12159 (N_12159,N_11892,N_11852);
nor U12160 (N_12160,N_11978,N_11940);
nor U12161 (N_12161,N_11978,N_11963);
xnor U12162 (N_12162,N_11984,N_11996);
nor U12163 (N_12163,N_11895,N_11882);
nor U12164 (N_12164,N_11930,N_11899);
or U12165 (N_12165,N_11962,N_11850);
or U12166 (N_12166,N_11980,N_11859);
xor U12167 (N_12167,N_11872,N_11871);
nand U12168 (N_12168,N_11898,N_11874);
xnor U12169 (N_12169,N_11875,N_11896);
or U12170 (N_12170,N_11870,N_11804);
nand U12171 (N_12171,N_11969,N_11975);
or U12172 (N_12172,N_11980,N_11890);
nor U12173 (N_12173,N_11913,N_11943);
nor U12174 (N_12174,N_11908,N_11997);
and U12175 (N_12175,N_11912,N_11829);
nand U12176 (N_12176,N_11924,N_11882);
nand U12177 (N_12177,N_11854,N_11905);
xnor U12178 (N_12178,N_11826,N_11995);
and U12179 (N_12179,N_11935,N_11892);
nand U12180 (N_12180,N_11827,N_11967);
xnor U12181 (N_12181,N_11923,N_11939);
nor U12182 (N_12182,N_11859,N_11893);
or U12183 (N_12183,N_11900,N_11927);
and U12184 (N_12184,N_11857,N_11910);
xor U12185 (N_12185,N_11909,N_11823);
or U12186 (N_12186,N_11869,N_11940);
and U12187 (N_12187,N_11833,N_11981);
or U12188 (N_12188,N_11865,N_11970);
xnor U12189 (N_12189,N_11956,N_11971);
nor U12190 (N_12190,N_11810,N_11853);
nand U12191 (N_12191,N_11947,N_11875);
or U12192 (N_12192,N_11917,N_11877);
and U12193 (N_12193,N_11940,N_11930);
or U12194 (N_12194,N_11862,N_11993);
and U12195 (N_12195,N_11958,N_11914);
or U12196 (N_12196,N_11885,N_11951);
or U12197 (N_12197,N_11875,N_11828);
or U12198 (N_12198,N_11826,N_11996);
xnor U12199 (N_12199,N_11909,N_11942);
and U12200 (N_12200,N_12137,N_12141);
nand U12201 (N_12201,N_12065,N_12153);
nor U12202 (N_12202,N_12096,N_12149);
and U12203 (N_12203,N_12112,N_12002);
nand U12204 (N_12204,N_12019,N_12157);
or U12205 (N_12205,N_12148,N_12068);
or U12206 (N_12206,N_12172,N_12115);
xnor U12207 (N_12207,N_12132,N_12134);
or U12208 (N_12208,N_12171,N_12143);
and U12209 (N_12209,N_12183,N_12080);
and U12210 (N_12210,N_12184,N_12135);
nand U12211 (N_12211,N_12175,N_12188);
xor U12212 (N_12212,N_12166,N_12165);
nand U12213 (N_12213,N_12042,N_12057);
nor U12214 (N_12214,N_12027,N_12178);
and U12215 (N_12215,N_12140,N_12063);
nor U12216 (N_12216,N_12170,N_12197);
and U12217 (N_12217,N_12189,N_12104);
xor U12218 (N_12218,N_12113,N_12014);
or U12219 (N_12219,N_12161,N_12168);
nor U12220 (N_12220,N_12029,N_12088);
and U12221 (N_12221,N_12047,N_12111);
or U12222 (N_12222,N_12128,N_12145);
nand U12223 (N_12223,N_12036,N_12018);
nand U12224 (N_12224,N_12163,N_12147);
xor U12225 (N_12225,N_12131,N_12092);
and U12226 (N_12226,N_12006,N_12154);
and U12227 (N_12227,N_12050,N_12001);
and U12228 (N_12228,N_12009,N_12110);
and U12229 (N_12229,N_12159,N_12011);
xor U12230 (N_12230,N_12117,N_12123);
nand U12231 (N_12231,N_12079,N_12031);
nand U12232 (N_12232,N_12054,N_12162);
nand U12233 (N_12233,N_12000,N_12102);
nor U12234 (N_12234,N_12194,N_12186);
xnor U12235 (N_12235,N_12138,N_12017);
or U12236 (N_12236,N_12158,N_12106);
or U12237 (N_12237,N_12059,N_12152);
nand U12238 (N_12238,N_12198,N_12037);
nand U12239 (N_12239,N_12090,N_12005);
nor U12240 (N_12240,N_12010,N_12173);
nor U12241 (N_12241,N_12073,N_12032);
and U12242 (N_12242,N_12087,N_12044);
and U12243 (N_12243,N_12192,N_12034);
or U12244 (N_12244,N_12139,N_12187);
xor U12245 (N_12245,N_12043,N_12176);
and U12246 (N_12246,N_12013,N_12093);
nor U12247 (N_12247,N_12064,N_12179);
nand U12248 (N_12248,N_12150,N_12026);
and U12249 (N_12249,N_12066,N_12038);
nand U12250 (N_12250,N_12193,N_12052);
nor U12251 (N_12251,N_12182,N_12012);
and U12252 (N_12252,N_12181,N_12056);
xor U12253 (N_12253,N_12133,N_12021);
nand U12254 (N_12254,N_12167,N_12062);
and U12255 (N_12255,N_12109,N_12028);
xnor U12256 (N_12256,N_12033,N_12097);
and U12257 (N_12257,N_12156,N_12122);
xor U12258 (N_12258,N_12164,N_12020);
or U12259 (N_12259,N_12146,N_12091);
nor U12260 (N_12260,N_12035,N_12169);
nand U12261 (N_12261,N_12070,N_12105);
nand U12262 (N_12262,N_12084,N_12119);
or U12263 (N_12263,N_12126,N_12040);
nor U12264 (N_12264,N_12185,N_12069);
xnor U12265 (N_12265,N_12078,N_12015);
nor U12266 (N_12266,N_12071,N_12108);
nand U12267 (N_12267,N_12196,N_12008);
and U12268 (N_12268,N_12082,N_12045);
or U12269 (N_12269,N_12025,N_12130);
xnor U12270 (N_12270,N_12101,N_12107);
xor U12271 (N_12271,N_12074,N_12076);
and U12272 (N_12272,N_12155,N_12058);
nand U12273 (N_12273,N_12003,N_12089);
xnor U12274 (N_12274,N_12121,N_12030);
xor U12275 (N_12275,N_12151,N_12072);
nor U12276 (N_12276,N_12125,N_12016);
nor U12277 (N_12277,N_12199,N_12127);
and U12278 (N_12278,N_12103,N_12048);
nor U12279 (N_12279,N_12142,N_12094);
xor U12280 (N_12280,N_12081,N_12041);
and U12281 (N_12281,N_12124,N_12023);
and U12282 (N_12282,N_12174,N_12051);
nand U12283 (N_12283,N_12116,N_12180);
and U12284 (N_12284,N_12067,N_12160);
xor U12285 (N_12285,N_12144,N_12095);
xor U12286 (N_12286,N_12129,N_12053);
nor U12287 (N_12287,N_12060,N_12098);
nand U12288 (N_12288,N_12024,N_12075);
and U12289 (N_12289,N_12114,N_12086);
nor U12290 (N_12290,N_12007,N_12195);
nor U12291 (N_12291,N_12004,N_12177);
xor U12292 (N_12292,N_12120,N_12055);
and U12293 (N_12293,N_12046,N_12190);
xnor U12294 (N_12294,N_12083,N_12022);
and U12295 (N_12295,N_12191,N_12100);
nand U12296 (N_12296,N_12136,N_12118);
or U12297 (N_12297,N_12061,N_12049);
xnor U12298 (N_12298,N_12099,N_12077);
xnor U12299 (N_12299,N_12085,N_12039);
nor U12300 (N_12300,N_12134,N_12109);
xnor U12301 (N_12301,N_12099,N_12056);
nand U12302 (N_12302,N_12131,N_12041);
xor U12303 (N_12303,N_12077,N_12085);
or U12304 (N_12304,N_12128,N_12180);
nand U12305 (N_12305,N_12126,N_12045);
and U12306 (N_12306,N_12092,N_12116);
or U12307 (N_12307,N_12065,N_12143);
nand U12308 (N_12308,N_12053,N_12083);
and U12309 (N_12309,N_12088,N_12035);
or U12310 (N_12310,N_12092,N_12122);
xor U12311 (N_12311,N_12115,N_12123);
xor U12312 (N_12312,N_12190,N_12176);
nand U12313 (N_12313,N_12088,N_12186);
and U12314 (N_12314,N_12001,N_12048);
nand U12315 (N_12315,N_12179,N_12079);
xor U12316 (N_12316,N_12105,N_12128);
nand U12317 (N_12317,N_12026,N_12014);
nor U12318 (N_12318,N_12006,N_12030);
and U12319 (N_12319,N_12122,N_12026);
nor U12320 (N_12320,N_12116,N_12089);
nor U12321 (N_12321,N_12114,N_12028);
nand U12322 (N_12322,N_12057,N_12005);
nand U12323 (N_12323,N_12018,N_12148);
xor U12324 (N_12324,N_12042,N_12049);
nand U12325 (N_12325,N_12036,N_12078);
xor U12326 (N_12326,N_12045,N_12084);
xnor U12327 (N_12327,N_12092,N_12115);
nor U12328 (N_12328,N_12001,N_12094);
and U12329 (N_12329,N_12096,N_12155);
xor U12330 (N_12330,N_12110,N_12081);
and U12331 (N_12331,N_12039,N_12090);
nand U12332 (N_12332,N_12027,N_12052);
nand U12333 (N_12333,N_12167,N_12188);
nor U12334 (N_12334,N_12173,N_12095);
or U12335 (N_12335,N_12104,N_12055);
xnor U12336 (N_12336,N_12026,N_12047);
nor U12337 (N_12337,N_12109,N_12165);
or U12338 (N_12338,N_12186,N_12005);
nand U12339 (N_12339,N_12033,N_12042);
or U12340 (N_12340,N_12033,N_12083);
nand U12341 (N_12341,N_12106,N_12167);
and U12342 (N_12342,N_12081,N_12150);
or U12343 (N_12343,N_12130,N_12062);
xnor U12344 (N_12344,N_12109,N_12143);
and U12345 (N_12345,N_12054,N_12003);
nor U12346 (N_12346,N_12055,N_12023);
xnor U12347 (N_12347,N_12164,N_12055);
nand U12348 (N_12348,N_12116,N_12187);
or U12349 (N_12349,N_12106,N_12066);
nor U12350 (N_12350,N_12070,N_12072);
and U12351 (N_12351,N_12053,N_12191);
xnor U12352 (N_12352,N_12130,N_12037);
nand U12353 (N_12353,N_12130,N_12147);
xnor U12354 (N_12354,N_12058,N_12012);
or U12355 (N_12355,N_12148,N_12008);
xnor U12356 (N_12356,N_12178,N_12041);
and U12357 (N_12357,N_12149,N_12107);
nor U12358 (N_12358,N_12094,N_12087);
and U12359 (N_12359,N_12044,N_12100);
and U12360 (N_12360,N_12012,N_12165);
and U12361 (N_12361,N_12048,N_12183);
nand U12362 (N_12362,N_12158,N_12022);
or U12363 (N_12363,N_12064,N_12007);
xnor U12364 (N_12364,N_12076,N_12049);
nand U12365 (N_12365,N_12051,N_12084);
nor U12366 (N_12366,N_12031,N_12058);
nor U12367 (N_12367,N_12180,N_12169);
nand U12368 (N_12368,N_12184,N_12140);
and U12369 (N_12369,N_12148,N_12043);
nand U12370 (N_12370,N_12011,N_12147);
nand U12371 (N_12371,N_12161,N_12040);
nor U12372 (N_12372,N_12073,N_12111);
nor U12373 (N_12373,N_12149,N_12041);
or U12374 (N_12374,N_12168,N_12123);
or U12375 (N_12375,N_12132,N_12073);
xor U12376 (N_12376,N_12061,N_12135);
or U12377 (N_12377,N_12041,N_12090);
nand U12378 (N_12378,N_12033,N_12098);
and U12379 (N_12379,N_12054,N_12031);
and U12380 (N_12380,N_12018,N_12187);
or U12381 (N_12381,N_12051,N_12004);
nor U12382 (N_12382,N_12092,N_12129);
and U12383 (N_12383,N_12073,N_12029);
xor U12384 (N_12384,N_12173,N_12088);
nor U12385 (N_12385,N_12087,N_12120);
nand U12386 (N_12386,N_12062,N_12079);
nand U12387 (N_12387,N_12129,N_12025);
or U12388 (N_12388,N_12091,N_12192);
xnor U12389 (N_12389,N_12102,N_12174);
nand U12390 (N_12390,N_12106,N_12121);
nand U12391 (N_12391,N_12005,N_12179);
nor U12392 (N_12392,N_12057,N_12038);
or U12393 (N_12393,N_12037,N_12196);
or U12394 (N_12394,N_12170,N_12066);
nor U12395 (N_12395,N_12033,N_12127);
nand U12396 (N_12396,N_12199,N_12036);
xor U12397 (N_12397,N_12171,N_12075);
or U12398 (N_12398,N_12079,N_12113);
xor U12399 (N_12399,N_12004,N_12010);
or U12400 (N_12400,N_12383,N_12293);
xor U12401 (N_12401,N_12256,N_12272);
and U12402 (N_12402,N_12262,N_12397);
or U12403 (N_12403,N_12322,N_12288);
nor U12404 (N_12404,N_12253,N_12235);
and U12405 (N_12405,N_12247,N_12213);
nand U12406 (N_12406,N_12274,N_12241);
and U12407 (N_12407,N_12231,N_12207);
and U12408 (N_12408,N_12346,N_12296);
xor U12409 (N_12409,N_12384,N_12280);
nand U12410 (N_12410,N_12363,N_12279);
or U12411 (N_12411,N_12350,N_12298);
xor U12412 (N_12412,N_12373,N_12237);
or U12413 (N_12413,N_12372,N_12277);
and U12414 (N_12414,N_12200,N_12378);
nor U12415 (N_12415,N_12357,N_12345);
nand U12416 (N_12416,N_12331,N_12368);
nand U12417 (N_12417,N_12206,N_12287);
nor U12418 (N_12418,N_12358,N_12223);
xor U12419 (N_12419,N_12324,N_12392);
and U12420 (N_12420,N_12220,N_12334);
and U12421 (N_12421,N_12219,N_12259);
and U12422 (N_12422,N_12362,N_12315);
nand U12423 (N_12423,N_12254,N_12236);
nor U12424 (N_12424,N_12240,N_12349);
and U12425 (N_12425,N_12308,N_12359);
xnor U12426 (N_12426,N_12330,N_12335);
or U12427 (N_12427,N_12264,N_12234);
xor U12428 (N_12428,N_12365,N_12270);
or U12429 (N_12429,N_12267,N_12367);
nor U12430 (N_12430,N_12297,N_12348);
nand U12431 (N_12431,N_12321,N_12281);
and U12432 (N_12432,N_12214,N_12306);
and U12433 (N_12433,N_12337,N_12381);
nor U12434 (N_12434,N_12309,N_12375);
and U12435 (N_12435,N_12300,N_12258);
xor U12436 (N_12436,N_12250,N_12252);
nor U12437 (N_12437,N_12283,N_12347);
nor U12438 (N_12438,N_12376,N_12261);
nand U12439 (N_12439,N_12313,N_12266);
nand U12440 (N_12440,N_12354,N_12394);
nand U12441 (N_12441,N_12380,N_12260);
xor U12442 (N_12442,N_12278,N_12202);
nand U12443 (N_12443,N_12232,N_12389);
xnor U12444 (N_12444,N_12239,N_12269);
or U12445 (N_12445,N_12336,N_12273);
and U12446 (N_12446,N_12326,N_12221);
xnor U12447 (N_12447,N_12325,N_12385);
nor U12448 (N_12448,N_12374,N_12341);
nand U12449 (N_12449,N_12311,N_12387);
nor U12450 (N_12450,N_12217,N_12371);
or U12451 (N_12451,N_12285,N_12303);
nor U12452 (N_12452,N_12360,N_12230);
or U12453 (N_12453,N_12343,N_12388);
nand U12454 (N_12454,N_12390,N_12314);
and U12455 (N_12455,N_12242,N_12344);
and U12456 (N_12456,N_12291,N_12265);
xnor U12457 (N_12457,N_12205,N_12275);
and U12458 (N_12458,N_12292,N_12332);
or U12459 (N_12459,N_12339,N_12227);
or U12460 (N_12460,N_12316,N_12209);
or U12461 (N_12461,N_12229,N_12386);
or U12462 (N_12462,N_12340,N_12244);
xor U12463 (N_12463,N_12201,N_12370);
nand U12464 (N_12464,N_12276,N_12204);
or U12465 (N_12465,N_12304,N_12249);
xor U12466 (N_12466,N_12268,N_12333);
and U12467 (N_12467,N_12355,N_12233);
nor U12468 (N_12468,N_12301,N_12224);
and U12469 (N_12469,N_12382,N_12302);
or U12470 (N_12470,N_12245,N_12319);
nor U12471 (N_12471,N_12212,N_12294);
or U12472 (N_12472,N_12218,N_12305);
nand U12473 (N_12473,N_12286,N_12395);
nor U12474 (N_12474,N_12352,N_12295);
or U12475 (N_12475,N_12312,N_12222);
nor U12476 (N_12476,N_12307,N_12328);
nand U12477 (N_12477,N_12255,N_12228);
nand U12478 (N_12478,N_12238,N_12377);
and U12479 (N_12479,N_12398,N_12353);
nor U12480 (N_12480,N_12393,N_12215);
nor U12481 (N_12481,N_12379,N_12211);
or U12482 (N_12482,N_12226,N_12290);
or U12483 (N_12483,N_12271,N_12338);
or U12484 (N_12484,N_12399,N_12327);
and U12485 (N_12485,N_12251,N_12310);
or U12486 (N_12486,N_12391,N_12329);
or U12487 (N_12487,N_12361,N_12225);
or U12488 (N_12488,N_12282,N_12320);
nand U12489 (N_12489,N_12284,N_12208);
xor U12490 (N_12490,N_12210,N_12356);
nor U12491 (N_12491,N_12342,N_12366);
xor U12492 (N_12492,N_12248,N_12364);
or U12493 (N_12493,N_12246,N_12243);
xnor U12494 (N_12494,N_12351,N_12299);
or U12495 (N_12495,N_12203,N_12289);
nand U12496 (N_12496,N_12318,N_12257);
nor U12497 (N_12497,N_12317,N_12369);
xnor U12498 (N_12498,N_12263,N_12323);
xor U12499 (N_12499,N_12396,N_12216);
nor U12500 (N_12500,N_12372,N_12269);
and U12501 (N_12501,N_12218,N_12269);
xor U12502 (N_12502,N_12362,N_12364);
xnor U12503 (N_12503,N_12251,N_12301);
xor U12504 (N_12504,N_12227,N_12398);
xor U12505 (N_12505,N_12232,N_12311);
xnor U12506 (N_12506,N_12382,N_12391);
nand U12507 (N_12507,N_12363,N_12372);
and U12508 (N_12508,N_12347,N_12397);
xnor U12509 (N_12509,N_12366,N_12285);
nand U12510 (N_12510,N_12348,N_12292);
nor U12511 (N_12511,N_12312,N_12321);
xnor U12512 (N_12512,N_12231,N_12302);
or U12513 (N_12513,N_12308,N_12378);
nand U12514 (N_12514,N_12365,N_12398);
and U12515 (N_12515,N_12298,N_12275);
nand U12516 (N_12516,N_12285,N_12291);
and U12517 (N_12517,N_12322,N_12289);
and U12518 (N_12518,N_12279,N_12217);
or U12519 (N_12519,N_12342,N_12225);
nor U12520 (N_12520,N_12269,N_12276);
nand U12521 (N_12521,N_12259,N_12276);
nand U12522 (N_12522,N_12357,N_12363);
xnor U12523 (N_12523,N_12334,N_12252);
nor U12524 (N_12524,N_12277,N_12214);
and U12525 (N_12525,N_12206,N_12249);
or U12526 (N_12526,N_12290,N_12246);
nand U12527 (N_12527,N_12285,N_12230);
and U12528 (N_12528,N_12320,N_12206);
nand U12529 (N_12529,N_12266,N_12304);
nor U12530 (N_12530,N_12251,N_12206);
nand U12531 (N_12531,N_12304,N_12260);
and U12532 (N_12532,N_12309,N_12215);
and U12533 (N_12533,N_12211,N_12382);
or U12534 (N_12534,N_12297,N_12264);
or U12535 (N_12535,N_12265,N_12252);
or U12536 (N_12536,N_12260,N_12233);
or U12537 (N_12537,N_12299,N_12288);
or U12538 (N_12538,N_12352,N_12313);
nand U12539 (N_12539,N_12301,N_12342);
nor U12540 (N_12540,N_12324,N_12293);
and U12541 (N_12541,N_12322,N_12248);
xnor U12542 (N_12542,N_12284,N_12219);
nand U12543 (N_12543,N_12376,N_12353);
nand U12544 (N_12544,N_12363,N_12355);
xnor U12545 (N_12545,N_12305,N_12302);
or U12546 (N_12546,N_12261,N_12229);
or U12547 (N_12547,N_12239,N_12363);
nor U12548 (N_12548,N_12328,N_12257);
nor U12549 (N_12549,N_12391,N_12306);
and U12550 (N_12550,N_12240,N_12314);
and U12551 (N_12551,N_12275,N_12379);
or U12552 (N_12552,N_12249,N_12254);
xor U12553 (N_12553,N_12283,N_12391);
nand U12554 (N_12554,N_12255,N_12367);
and U12555 (N_12555,N_12214,N_12338);
and U12556 (N_12556,N_12296,N_12343);
nor U12557 (N_12557,N_12369,N_12249);
nor U12558 (N_12558,N_12392,N_12225);
and U12559 (N_12559,N_12294,N_12325);
or U12560 (N_12560,N_12362,N_12280);
nand U12561 (N_12561,N_12329,N_12201);
and U12562 (N_12562,N_12227,N_12289);
or U12563 (N_12563,N_12228,N_12349);
nor U12564 (N_12564,N_12335,N_12394);
or U12565 (N_12565,N_12258,N_12259);
or U12566 (N_12566,N_12264,N_12395);
xnor U12567 (N_12567,N_12369,N_12285);
or U12568 (N_12568,N_12264,N_12337);
nor U12569 (N_12569,N_12279,N_12268);
or U12570 (N_12570,N_12317,N_12252);
xnor U12571 (N_12571,N_12253,N_12261);
nor U12572 (N_12572,N_12380,N_12318);
nand U12573 (N_12573,N_12230,N_12234);
and U12574 (N_12574,N_12224,N_12361);
or U12575 (N_12575,N_12365,N_12379);
xor U12576 (N_12576,N_12203,N_12211);
nor U12577 (N_12577,N_12312,N_12343);
xor U12578 (N_12578,N_12323,N_12293);
nand U12579 (N_12579,N_12255,N_12350);
or U12580 (N_12580,N_12286,N_12376);
nor U12581 (N_12581,N_12214,N_12360);
or U12582 (N_12582,N_12370,N_12244);
or U12583 (N_12583,N_12215,N_12220);
or U12584 (N_12584,N_12397,N_12209);
nor U12585 (N_12585,N_12339,N_12218);
and U12586 (N_12586,N_12297,N_12263);
or U12587 (N_12587,N_12295,N_12275);
xor U12588 (N_12588,N_12283,N_12296);
and U12589 (N_12589,N_12279,N_12264);
and U12590 (N_12590,N_12356,N_12361);
and U12591 (N_12591,N_12217,N_12285);
and U12592 (N_12592,N_12345,N_12298);
nor U12593 (N_12593,N_12395,N_12288);
nand U12594 (N_12594,N_12286,N_12213);
and U12595 (N_12595,N_12364,N_12261);
or U12596 (N_12596,N_12353,N_12234);
and U12597 (N_12597,N_12264,N_12208);
nand U12598 (N_12598,N_12362,N_12381);
xor U12599 (N_12599,N_12354,N_12346);
and U12600 (N_12600,N_12515,N_12555);
nand U12601 (N_12601,N_12469,N_12552);
xnor U12602 (N_12602,N_12586,N_12403);
xnor U12603 (N_12603,N_12446,N_12561);
nand U12604 (N_12604,N_12412,N_12413);
nor U12605 (N_12605,N_12548,N_12503);
or U12606 (N_12606,N_12571,N_12589);
or U12607 (N_12607,N_12463,N_12437);
or U12608 (N_12608,N_12583,N_12529);
or U12609 (N_12609,N_12535,N_12514);
nor U12610 (N_12610,N_12498,N_12579);
or U12611 (N_12611,N_12482,N_12542);
nand U12612 (N_12612,N_12546,N_12504);
nor U12613 (N_12613,N_12577,N_12499);
nand U12614 (N_12614,N_12440,N_12594);
nor U12615 (N_12615,N_12430,N_12418);
and U12616 (N_12616,N_12458,N_12592);
nand U12617 (N_12617,N_12435,N_12473);
and U12618 (N_12618,N_12584,N_12596);
or U12619 (N_12619,N_12461,N_12532);
nand U12620 (N_12620,N_12533,N_12509);
nor U12621 (N_12621,N_12474,N_12443);
xnor U12622 (N_12622,N_12526,N_12585);
nand U12623 (N_12623,N_12449,N_12534);
and U12624 (N_12624,N_12550,N_12408);
or U12625 (N_12625,N_12574,N_12481);
or U12626 (N_12626,N_12434,N_12530);
nand U12627 (N_12627,N_12576,N_12490);
and U12628 (N_12628,N_12562,N_12587);
and U12629 (N_12629,N_12554,N_12420);
xor U12630 (N_12630,N_12531,N_12497);
or U12631 (N_12631,N_12450,N_12580);
and U12632 (N_12632,N_12519,N_12537);
or U12633 (N_12633,N_12527,N_12484);
xor U12634 (N_12634,N_12563,N_12512);
nor U12635 (N_12635,N_12410,N_12540);
and U12636 (N_12636,N_12553,N_12453);
or U12637 (N_12637,N_12429,N_12451);
and U12638 (N_12638,N_12517,N_12457);
xor U12639 (N_12639,N_12578,N_12433);
nor U12640 (N_12640,N_12494,N_12505);
nand U12641 (N_12641,N_12559,N_12564);
xnor U12642 (N_12642,N_12456,N_12448);
nand U12643 (N_12643,N_12428,N_12572);
and U12644 (N_12644,N_12427,N_12471);
nand U12645 (N_12645,N_12582,N_12501);
nor U12646 (N_12646,N_12581,N_12478);
nand U12647 (N_12647,N_12496,N_12522);
or U12648 (N_12648,N_12447,N_12414);
and U12649 (N_12649,N_12558,N_12479);
nor U12650 (N_12650,N_12421,N_12441);
nor U12651 (N_12651,N_12470,N_12566);
nor U12652 (N_12652,N_12445,N_12400);
and U12653 (N_12653,N_12439,N_12464);
or U12654 (N_12654,N_12468,N_12426);
or U12655 (N_12655,N_12477,N_12513);
or U12656 (N_12656,N_12523,N_12568);
xnor U12657 (N_12657,N_12521,N_12415);
nor U12658 (N_12658,N_12569,N_12599);
xor U12659 (N_12659,N_12405,N_12539);
or U12660 (N_12660,N_12436,N_12573);
nand U12661 (N_12661,N_12422,N_12538);
xor U12662 (N_12662,N_12595,N_12485);
or U12663 (N_12663,N_12491,N_12570);
xnor U12664 (N_12664,N_12455,N_12544);
or U12665 (N_12665,N_12465,N_12502);
and U12666 (N_12666,N_12567,N_12402);
xor U12667 (N_12667,N_12590,N_12460);
xnor U12668 (N_12668,N_12475,N_12486);
and U12669 (N_12669,N_12493,N_12549);
or U12670 (N_12670,N_12432,N_12419);
nand U12671 (N_12671,N_12407,N_12506);
and U12672 (N_12672,N_12598,N_12597);
nand U12673 (N_12673,N_12588,N_12518);
and U12674 (N_12674,N_12454,N_12516);
or U12675 (N_12675,N_12560,N_12593);
xor U12676 (N_12676,N_12557,N_12528);
and U12677 (N_12677,N_12462,N_12466);
xnor U12678 (N_12678,N_12492,N_12565);
nand U12679 (N_12679,N_12423,N_12575);
or U12680 (N_12680,N_12547,N_12591);
nand U12681 (N_12681,N_12483,N_12404);
nand U12682 (N_12682,N_12543,N_12480);
and U12683 (N_12683,N_12545,N_12551);
nor U12684 (N_12684,N_12424,N_12476);
and U12685 (N_12685,N_12495,N_12507);
nand U12686 (N_12686,N_12467,N_12487);
and U12687 (N_12687,N_12411,N_12444);
nor U12688 (N_12688,N_12409,N_12511);
or U12689 (N_12689,N_12406,N_12500);
or U12690 (N_12690,N_12431,N_12541);
and U12691 (N_12691,N_12417,N_12556);
nor U12692 (N_12692,N_12520,N_12472);
xnor U12693 (N_12693,N_12452,N_12416);
xnor U12694 (N_12694,N_12442,N_12488);
xor U12695 (N_12695,N_12525,N_12508);
and U12696 (N_12696,N_12510,N_12536);
nor U12697 (N_12697,N_12489,N_12459);
nand U12698 (N_12698,N_12438,N_12401);
xor U12699 (N_12699,N_12524,N_12425);
or U12700 (N_12700,N_12477,N_12481);
and U12701 (N_12701,N_12430,N_12549);
xor U12702 (N_12702,N_12456,N_12454);
xor U12703 (N_12703,N_12567,N_12518);
or U12704 (N_12704,N_12493,N_12550);
and U12705 (N_12705,N_12498,N_12529);
nand U12706 (N_12706,N_12501,N_12566);
and U12707 (N_12707,N_12433,N_12553);
or U12708 (N_12708,N_12444,N_12453);
nor U12709 (N_12709,N_12460,N_12500);
or U12710 (N_12710,N_12466,N_12452);
xor U12711 (N_12711,N_12499,N_12592);
and U12712 (N_12712,N_12557,N_12521);
or U12713 (N_12713,N_12410,N_12463);
and U12714 (N_12714,N_12422,N_12511);
nand U12715 (N_12715,N_12410,N_12477);
xnor U12716 (N_12716,N_12437,N_12571);
nand U12717 (N_12717,N_12534,N_12487);
or U12718 (N_12718,N_12545,N_12436);
and U12719 (N_12719,N_12557,N_12437);
and U12720 (N_12720,N_12492,N_12570);
or U12721 (N_12721,N_12469,N_12403);
nand U12722 (N_12722,N_12497,N_12467);
and U12723 (N_12723,N_12429,N_12594);
and U12724 (N_12724,N_12407,N_12556);
nand U12725 (N_12725,N_12424,N_12530);
or U12726 (N_12726,N_12529,N_12413);
nor U12727 (N_12727,N_12556,N_12537);
and U12728 (N_12728,N_12568,N_12424);
nand U12729 (N_12729,N_12506,N_12519);
and U12730 (N_12730,N_12592,N_12474);
nand U12731 (N_12731,N_12469,N_12457);
and U12732 (N_12732,N_12515,N_12492);
xnor U12733 (N_12733,N_12593,N_12408);
nand U12734 (N_12734,N_12502,N_12558);
and U12735 (N_12735,N_12505,N_12417);
nor U12736 (N_12736,N_12480,N_12595);
xnor U12737 (N_12737,N_12430,N_12504);
xnor U12738 (N_12738,N_12548,N_12472);
nor U12739 (N_12739,N_12530,N_12507);
and U12740 (N_12740,N_12479,N_12550);
xnor U12741 (N_12741,N_12556,N_12476);
nand U12742 (N_12742,N_12542,N_12525);
or U12743 (N_12743,N_12504,N_12492);
nand U12744 (N_12744,N_12444,N_12537);
or U12745 (N_12745,N_12586,N_12555);
nor U12746 (N_12746,N_12580,N_12502);
and U12747 (N_12747,N_12456,N_12450);
or U12748 (N_12748,N_12579,N_12586);
or U12749 (N_12749,N_12430,N_12536);
nand U12750 (N_12750,N_12489,N_12527);
nand U12751 (N_12751,N_12594,N_12525);
nor U12752 (N_12752,N_12562,N_12531);
nand U12753 (N_12753,N_12443,N_12535);
nor U12754 (N_12754,N_12500,N_12499);
and U12755 (N_12755,N_12497,N_12452);
or U12756 (N_12756,N_12455,N_12524);
and U12757 (N_12757,N_12532,N_12587);
nor U12758 (N_12758,N_12477,N_12499);
and U12759 (N_12759,N_12493,N_12412);
xor U12760 (N_12760,N_12400,N_12451);
or U12761 (N_12761,N_12541,N_12592);
nand U12762 (N_12762,N_12511,N_12474);
or U12763 (N_12763,N_12419,N_12563);
nor U12764 (N_12764,N_12469,N_12598);
xor U12765 (N_12765,N_12555,N_12566);
xnor U12766 (N_12766,N_12405,N_12580);
and U12767 (N_12767,N_12536,N_12571);
nand U12768 (N_12768,N_12552,N_12567);
and U12769 (N_12769,N_12498,N_12575);
xnor U12770 (N_12770,N_12453,N_12438);
nand U12771 (N_12771,N_12560,N_12556);
or U12772 (N_12772,N_12426,N_12535);
xnor U12773 (N_12773,N_12528,N_12597);
and U12774 (N_12774,N_12424,N_12427);
or U12775 (N_12775,N_12481,N_12551);
and U12776 (N_12776,N_12475,N_12566);
and U12777 (N_12777,N_12560,N_12575);
xnor U12778 (N_12778,N_12464,N_12517);
nor U12779 (N_12779,N_12470,N_12415);
xnor U12780 (N_12780,N_12460,N_12490);
nand U12781 (N_12781,N_12598,N_12416);
nand U12782 (N_12782,N_12530,N_12486);
nor U12783 (N_12783,N_12477,N_12585);
and U12784 (N_12784,N_12506,N_12438);
and U12785 (N_12785,N_12575,N_12410);
xor U12786 (N_12786,N_12523,N_12593);
nand U12787 (N_12787,N_12596,N_12466);
nand U12788 (N_12788,N_12582,N_12485);
nand U12789 (N_12789,N_12496,N_12575);
or U12790 (N_12790,N_12534,N_12468);
xnor U12791 (N_12791,N_12409,N_12423);
nand U12792 (N_12792,N_12449,N_12458);
or U12793 (N_12793,N_12536,N_12532);
or U12794 (N_12794,N_12567,N_12599);
or U12795 (N_12795,N_12546,N_12492);
nand U12796 (N_12796,N_12449,N_12514);
nor U12797 (N_12797,N_12490,N_12488);
xor U12798 (N_12798,N_12573,N_12597);
nor U12799 (N_12799,N_12548,N_12443);
xor U12800 (N_12800,N_12664,N_12721);
nand U12801 (N_12801,N_12633,N_12706);
nor U12802 (N_12802,N_12611,N_12747);
and U12803 (N_12803,N_12768,N_12755);
or U12804 (N_12804,N_12651,N_12696);
nor U12805 (N_12805,N_12635,N_12794);
and U12806 (N_12806,N_12669,N_12629);
xor U12807 (N_12807,N_12738,N_12621);
nand U12808 (N_12808,N_12638,N_12766);
and U12809 (N_12809,N_12788,N_12695);
or U12810 (N_12810,N_12736,N_12751);
nand U12811 (N_12811,N_12607,N_12661);
or U12812 (N_12812,N_12620,N_12615);
xnor U12813 (N_12813,N_12626,N_12796);
xnor U12814 (N_12814,N_12682,N_12754);
xor U12815 (N_12815,N_12782,N_12717);
and U12816 (N_12816,N_12764,N_12731);
nor U12817 (N_12817,N_12627,N_12746);
nand U12818 (N_12818,N_12734,N_12618);
nor U12819 (N_12819,N_12634,N_12610);
and U12820 (N_12820,N_12771,N_12785);
nand U12821 (N_12821,N_12648,N_12623);
nand U12822 (N_12822,N_12761,N_12625);
xnor U12823 (N_12823,N_12719,N_12688);
nor U12824 (N_12824,N_12628,N_12658);
xnor U12825 (N_12825,N_12786,N_12767);
nand U12826 (N_12826,N_12645,N_12663);
nor U12827 (N_12827,N_12647,N_12740);
nor U12828 (N_12828,N_12653,N_12693);
or U12829 (N_12829,N_12703,N_12795);
nor U12830 (N_12830,N_12699,N_12713);
nor U12831 (N_12831,N_12685,N_12714);
and U12832 (N_12832,N_12781,N_12667);
or U12833 (N_12833,N_12650,N_12646);
nand U12834 (N_12834,N_12726,N_12660);
and U12835 (N_12835,N_12655,N_12614);
nand U12836 (N_12836,N_12622,N_12617);
nor U12837 (N_12837,N_12643,N_12665);
or U12838 (N_12838,N_12712,N_12636);
or U12839 (N_12839,N_12742,N_12798);
nor U12840 (N_12840,N_12637,N_12644);
xnor U12841 (N_12841,N_12765,N_12674);
nor U12842 (N_12842,N_12737,N_12739);
and U12843 (N_12843,N_12729,N_12715);
nand U12844 (N_12844,N_12612,N_12704);
and U12845 (N_12845,N_12631,N_12718);
and U12846 (N_12846,N_12709,N_12780);
xor U12847 (N_12847,N_12758,N_12642);
and U12848 (N_12848,N_12728,N_12750);
xnor U12849 (N_12849,N_12679,N_12748);
nand U12850 (N_12850,N_12694,N_12763);
xnor U12851 (N_12851,N_12797,N_12745);
xor U12852 (N_12852,N_12652,N_12753);
nor U12853 (N_12853,N_12600,N_12789);
or U12854 (N_12854,N_12659,N_12668);
xor U12855 (N_12855,N_12630,N_12662);
xnor U12856 (N_12856,N_12698,N_12707);
and U12857 (N_12857,N_12656,N_12670);
or U12858 (N_12858,N_12671,N_12723);
nand U12859 (N_12859,N_12735,N_12732);
or U12860 (N_12860,N_12601,N_12608);
nor U12861 (N_12861,N_12677,N_12790);
nand U12862 (N_12862,N_12609,N_12678);
nor U12863 (N_12863,N_12772,N_12720);
and U12864 (N_12864,N_12690,N_12716);
and U12865 (N_12865,N_12770,N_12701);
xor U12866 (N_12866,N_12779,N_12752);
nand U12867 (N_12867,N_12606,N_12641);
and U12868 (N_12868,N_12756,N_12792);
and U12869 (N_12869,N_12784,N_12775);
nand U12870 (N_12870,N_12692,N_12657);
nor U12871 (N_12871,N_12776,N_12743);
nand U12872 (N_12872,N_12705,N_12799);
xor U12873 (N_12873,N_12708,N_12639);
or U12874 (N_12874,N_12760,N_12759);
and U12875 (N_12875,N_12787,N_12686);
xor U12876 (N_12876,N_12683,N_12744);
xor U12877 (N_12877,N_12624,N_12680);
nand U12878 (N_12878,N_12681,N_12604);
or U12879 (N_12879,N_12778,N_12725);
xnor U12880 (N_12880,N_12672,N_12603);
and U12881 (N_12881,N_12673,N_12722);
or U12882 (N_12882,N_12793,N_12724);
or U12883 (N_12883,N_12602,N_12700);
nor U12884 (N_12884,N_12666,N_12791);
or U12885 (N_12885,N_12675,N_12741);
nor U12886 (N_12886,N_12684,N_12632);
nand U12887 (N_12887,N_12640,N_12727);
xor U12888 (N_12888,N_12711,N_12777);
and U12889 (N_12889,N_12783,N_12702);
and U12890 (N_12890,N_12605,N_12733);
nor U12891 (N_12891,N_12654,N_12773);
nand U12892 (N_12892,N_12769,N_12691);
xor U12893 (N_12893,N_12613,N_12619);
nand U12894 (N_12894,N_12710,N_12730);
or U12895 (N_12895,N_12616,N_12757);
xor U12896 (N_12896,N_12689,N_12676);
nand U12897 (N_12897,N_12649,N_12697);
nand U12898 (N_12898,N_12687,N_12749);
and U12899 (N_12899,N_12762,N_12774);
xor U12900 (N_12900,N_12661,N_12732);
and U12901 (N_12901,N_12797,N_12741);
nand U12902 (N_12902,N_12738,N_12688);
and U12903 (N_12903,N_12779,N_12797);
nor U12904 (N_12904,N_12703,N_12748);
or U12905 (N_12905,N_12690,N_12601);
or U12906 (N_12906,N_12697,N_12776);
or U12907 (N_12907,N_12789,N_12797);
and U12908 (N_12908,N_12698,N_12717);
nand U12909 (N_12909,N_12630,N_12798);
and U12910 (N_12910,N_12777,N_12685);
nand U12911 (N_12911,N_12709,N_12784);
nand U12912 (N_12912,N_12662,N_12651);
nor U12913 (N_12913,N_12786,N_12685);
xor U12914 (N_12914,N_12706,N_12675);
or U12915 (N_12915,N_12674,N_12613);
or U12916 (N_12916,N_12602,N_12647);
nor U12917 (N_12917,N_12764,N_12744);
nand U12918 (N_12918,N_12650,N_12658);
and U12919 (N_12919,N_12738,N_12660);
and U12920 (N_12920,N_12790,N_12606);
or U12921 (N_12921,N_12756,N_12709);
nor U12922 (N_12922,N_12778,N_12790);
and U12923 (N_12923,N_12708,N_12742);
xnor U12924 (N_12924,N_12689,N_12705);
nor U12925 (N_12925,N_12701,N_12620);
nand U12926 (N_12926,N_12696,N_12692);
nor U12927 (N_12927,N_12649,N_12791);
or U12928 (N_12928,N_12722,N_12714);
and U12929 (N_12929,N_12627,N_12779);
and U12930 (N_12930,N_12693,N_12781);
xor U12931 (N_12931,N_12659,N_12665);
or U12932 (N_12932,N_12653,N_12763);
or U12933 (N_12933,N_12636,N_12703);
xnor U12934 (N_12934,N_12642,N_12656);
nor U12935 (N_12935,N_12617,N_12639);
or U12936 (N_12936,N_12712,N_12702);
nand U12937 (N_12937,N_12620,N_12749);
xor U12938 (N_12938,N_12625,N_12737);
and U12939 (N_12939,N_12798,N_12786);
xor U12940 (N_12940,N_12735,N_12659);
xnor U12941 (N_12941,N_12768,N_12702);
or U12942 (N_12942,N_12688,N_12615);
and U12943 (N_12943,N_12738,N_12768);
and U12944 (N_12944,N_12665,N_12799);
and U12945 (N_12945,N_12751,N_12700);
and U12946 (N_12946,N_12792,N_12722);
nor U12947 (N_12947,N_12790,N_12678);
or U12948 (N_12948,N_12738,N_12758);
and U12949 (N_12949,N_12722,N_12609);
nand U12950 (N_12950,N_12757,N_12792);
nand U12951 (N_12951,N_12790,N_12769);
and U12952 (N_12952,N_12621,N_12707);
nand U12953 (N_12953,N_12760,N_12618);
nor U12954 (N_12954,N_12633,N_12798);
and U12955 (N_12955,N_12736,N_12792);
xnor U12956 (N_12956,N_12653,N_12682);
nand U12957 (N_12957,N_12731,N_12727);
or U12958 (N_12958,N_12657,N_12612);
nand U12959 (N_12959,N_12762,N_12637);
xnor U12960 (N_12960,N_12715,N_12753);
nand U12961 (N_12961,N_12606,N_12749);
xor U12962 (N_12962,N_12735,N_12771);
nand U12963 (N_12963,N_12758,N_12710);
or U12964 (N_12964,N_12679,N_12689);
nor U12965 (N_12965,N_12703,N_12625);
nand U12966 (N_12966,N_12704,N_12615);
xor U12967 (N_12967,N_12626,N_12640);
xor U12968 (N_12968,N_12772,N_12737);
nor U12969 (N_12969,N_12790,N_12785);
or U12970 (N_12970,N_12719,N_12687);
or U12971 (N_12971,N_12695,N_12759);
or U12972 (N_12972,N_12606,N_12780);
nor U12973 (N_12973,N_12675,N_12661);
and U12974 (N_12974,N_12727,N_12786);
or U12975 (N_12975,N_12613,N_12704);
nand U12976 (N_12976,N_12643,N_12659);
and U12977 (N_12977,N_12737,N_12776);
nand U12978 (N_12978,N_12716,N_12669);
or U12979 (N_12979,N_12673,N_12702);
xnor U12980 (N_12980,N_12723,N_12610);
nand U12981 (N_12981,N_12764,N_12758);
or U12982 (N_12982,N_12627,N_12789);
nor U12983 (N_12983,N_12695,N_12615);
nand U12984 (N_12984,N_12744,N_12737);
and U12985 (N_12985,N_12691,N_12711);
nand U12986 (N_12986,N_12629,N_12638);
or U12987 (N_12987,N_12752,N_12645);
xor U12988 (N_12988,N_12705,N_12620);
and U12989 (N_12989,N_12636,N_12650);
or U12990 (N_12990,N_12757,N_12648);
or U12991 (N_12991,N_12705,N_12758);
or U12992 (N_12992,N_12637,N_12607);
and U12993 (N_12993,N_12684,N_12756);
or U12994 (N_12994,N_12773,N_12675);
and U12995 (N_12995,N_12654,N_12612);
and U12996 (N_12996,N_12729,N_12766);
or U12997 (N_12997,N_12652,N_12655);
or U12998 (N_12998,N_12685,N_12752);
xnor U12999 (N_12999,N_12765,N_12680);
nand U13000 (N_13000,N_12866,N_12887);
or U13001 (N_13001,N_12920,N_12865);
or U13002 (N_13002,N_12925,N_12807);
xnor U13003 (N_13003,N_12882,N_12913);
or U13004 (N_13004,N_12822,N_12857);
nor U13005 (N_13005,N_12802,N_12935);
or U13006 (N_13006,N_12843,N_12858);
xnor U13007 (N_13007,N_12958,N_12812);
or U13008 (N_13008,N_12817,N_12934);
and U13009 (N_13009,N_12986,N_12830);
xnor U13010 (N_13010,N_12870,N_12828);
and U13011 (N_13011,N_12927,N_12991);
or U13012 (N_13012,N_12885,N_12914);
xnor U13013 (N_13013,N_12856,N_12979);
nor U13014 (N_13014,N_12988,N_12861);
nor U13015 (N_13015,N_12970,N_12845);
and U13016 (N_13016,N_12951,N_12944);
xnor U13017 (N_13017,N_12862,N_12909);
nand U13018 (N_13018,N_12829,N_12969);
xor U13019 (N_13019,N_12849,N_12893);
xor U13020 (N_13020,N_12808,N_12924);
nor U13021 (N_13021,N_12850,N_12959);
or U13022 (N_13022,N_12827,N_12846);
nor U13023 (N_13023,N_12881,N_12839);
nand U13024 (N_13024,N_12989,N_12886);
xor U13025 (N_13025,N_12968,N_12884);
nand U13026 (N_13026,N_12901,N_12900);
and U13027 (N_13027,N_12842,N_12872);
and U13028 (N_13028,N_12956,N_12910);
xor U13029 (N_13029,N_12998,N_12844);
xor U13030 (N_13030,N_12883,N_12985);
xnor U13031 (N_13031,N_12942,N_12929);
xor U13032 (N_13032,N_12869,N_12908);
nor U13033 (N_13033,N_12936,N_12810);
xnor U13034 (N_13034,N_12896,N_12904);
nand U13035 (N_13035,N_12868,N_12917);
nor U13036 (N_13036,N_12953,N_12938);
or U13037 (N_13037,N_12931,N_12863);
xor U13038 (N_13038,N_12820,N_12859);
and U13039 (N_13039,N_12852,N_12980);
nand U13040 (N_13040,N_12871,N_12873);
xnor U13041 (N_13041,N_12981,N_12889);
and U13042 (N_13042,N_12939,N_12945);
or U13043 (N_13043,N_12906,N_12918);
or U13044 (N_13044,N_12994,N_12964);
or U13045 (N_13045,N_12818,N_12947);
nor U13046 (N_13046,N_12905,N_12965);
xnor U13047 (N_13047,N_12974,N_12867);
or U13048 (N_13048,N_12853,N_12890);
nor U13049 (N_13049,N_12806,N_12875);
nand U13050 (N_13050,N_12847,N_12948);
or U13051 (N_13051,N_12813,N_12961);
xnor U13052 (N_13052,N_12874,N_12831);
xor U13053 (N_13053,N_12800,N_12815);
and U13054 (N_13054,N_12916,N_12876);
nand U13055 (N_13055,N_12878,N_12922);
nor U13056 (N_13056,N_12940,N_12814);
nor U13057 (N_13057,N_12950,N_12855);
xor U13058 (N_13058,N_12804,N_12946);
or U13059 (N_13059,N_12841,N_12836);
nor U13060 (N_13060,N_12962,N_12894);
xor U13061 (N_13061,N_12982,N_12803);
nand U13062 (N_13062,N_12915,N_12923);
and U13063 (N_13063,N_12903,N_12996);
nand U13064 (N_13064,N_12960,N_12811);
and U13065 (N_13065,N_12930,N_12877);
nand U13066 (N_13066,N_12943,N_12897);
or U13067 (N_13067,N_12933,N_12912);
nand U13068 (N_13068,N_12949,N_12921);
xnor U13069 (N_13069,N_12937,N_12834);
and U13070 (N_13070,N_12826,N_12983);
xnor U13071 (N_13071,N_12848,N_12963);
nand U13072 (N_13072,N_12824,N_12892);
xor U13073 (N_13073,N_12860,N_12854);
nor U13074 (N_13074,N_12957,N_12941);
xor U13075 (N_13075,N_12895,N_12809);
or U13076 (N_13076,N_12972,N_12999);
and U13077 (N_13077,N_12966,N_12902);
or U13078 (N_13078,N_12835,N_12891);
nor U13079 (N_13079,N_12978,N_12821);
xnor U13080 (N_13080,N_12823,N_12993);
nand U13081 (N_13081,N_12805,N_12967);
xnor U13082 (N_13082,N_12997,N_12840);
and U13083 (N_13083,N_12992,N_12880);
nor U13084 (N_13084,N_12911,N_12926);
xnor U13085 (N_13085,N_12975,N_12955);
nor U13086 (N_13086,N_12899,N_12816);
nor U13087 (N_13087,N_12952,N_12973);
xnor U13088 (N_13088,N_12990,N_12977);
nor U13089 (N_13089,N_12995,N_12838);
xnor U13090 (N_13090,N_12907,N_12928);
nor U13091 (N_13091,N_12976,N_12954);
and U13092 (N_13092,N_12833,N_12888);
xnor U13093 (N_13093,N_12984,N_12919);
and U13094 (N_13094,N_12832,N_12898);
and U13095 (N_13095,N_12932,N_12851);
xnor U13096 (N_13096,N_12879,N_12801);
or U13097 (N_13097,N_12987,N_12971);
nor U13098 (N_13098,N_12837,N_12825);
nand U13099 (N_13099,N_12864,N_12819);
and U13100 (N_13100,N_12834,N_12818);
nor U13101 (N_13101,N_12839,N_12880);
nand U13102 (N_13102,N_12873,N_12861);
or U13103 (N_13103,N_12894,N_12881);
nor U13104 (N_13104,N_12945,N_12838);
nand U13105 (N_13105,N_12822,N_12817);
nand U13106 (N_13106,N_12969,N_12857);
nand U13107 (N_13107,N_12980,N_12955);
nand U13108 (N_13108,N_12875,N_12993);
or U13109 (N_13109,N_12909,N_12994);
xor U13110 (N_13110,N_12872,N_12977);
and U13111 (N_13111,N_12900,N_12909);
xnor U13112 (N_13112,N_12833,N_12952);
nor U13113 (N_13113,N_12977,N_12861);
or U13114 (N_13114,N_12906,N_12967);
and U13115 (N_13115,N_12848,N_12899);
nand U13116 (N_13116,N_12918,N_12815);
nand U13117 (N_13117,N_12877,N_12851);
or U13118 (N_13118,N_12874,N_12917);
and U13119 (N_13119,N_12834,N_12892);
nor U13120 (N_13120,N_12913,N_12857);
and U13121 (N_13121,N_12979,N_12917);
and U13122 (N_13122,N_12963,N_12807);
or U13123 (N_13123,N_12808,N_12991);
xor U13124 (N_13124,N_12847,N_12926);
nor U13125 (N_13125,N_12887,N_12857);
xnor U13126 (N_13126,N_12830,N_12893);
nand U13127 (N_13127,N_12944,N_12985);
and U13128 (N_13128,N_12845,N_12870);
and U13129 (N_13129,N_12931,N_12872);
xor U13130 (N_13130,N_12973,N_12980);
nor U13131 (N_13131,N_12965,N_12882);
nor U13132 (N_13132,N_12851,N_12981);
or U13133 (N_13133,N_12844,N_12937);
xor U13134 (N_13134,N_12956,N_12859);
or U13135 (N_13135,N_12971,N_12888);
nand U13136 (N_13136,N_12872,N_12899);
and U13137 (N_13137,N_12878,N_12982);
xor U13138 (N_13138,N_12849,N_12958);
xnor U13139 (N_13139,N_12858,N_12804);
or U13140 (N_13140,N_12854,N_12963);
nand U13141 (N_13141,N_12841,N_12983);
xnor U13142 (N_13142,N_12876,N_12938);
nand U13143 (N_13143,N_12974,N_12862);
or U13144 (N_13144,N_12845,N_12813);
or U13145 (N_13145,N_12929,N_12875);
or U13146 (N_13146,N_12881,N_12869);
xnor U13147 (N_13147,N_12968,N_12907);
and U13148 (N_13148,N_12997,N_12814);
or U13149 (N_13149,N_12938,N_12825);
and U13150 (N_13150,N_12853,N_12829);
xor U13151 (N_13151,N_12859,N_12850);
nand U13152 (N_13152,N_12977,N_12959);
and U13153 (N_13153,N_12976,N_12807);
xor U13154 (N_13154,N_12849,N_12876);
nor U13155 (N_13155,N_12827,N_12917);
nor U13156 (N_13156,N_12804,N_12936);
nand U13157 (N_13157,N_12878,N_12834);
nor U13158 (N_13158,N_12872,N_12890);
nand U13159 (N_13159,N_12840,N_12982);
nand U13160 (N_13160,N_12811,N_12996);
xor U13161 (N_13161,N_12833,N_12945);
nor U13162 (N_13162,N_12949,N_12845);
xor U13163 (N_13163,N_12813,N_12952);
nand U13164 (N_13164,N_12818,N_12986);
nor U13165 (N_13165,N_12874,N_12842);
nor U13166 (N_13166,N_12921,N_12983);
nor U13167 (N_13167,N_12987,N_12957);
and U13168 (N_13168,N_12948,N_12818);
xnor U13169 (N_13169,N_12855,N_12853);
or U13170 (N_13170,N_12954,N_12833);
and U13171 (N_13171,N_12803,N_12969);
nand U13172 (N_13172,N_12915,N_12940);
or U13173 (N_13173,N_12807,N_12887);
or U13174 (N_13174,N_12826,N_12841);
or U13175 (N_13175,N_12957,N_12966);
and U13176 (N_13176,N_12869,N_12862);
or U13177 (N_13177,N_12895,N_12852);
or U13178 (N_13178,N_12895,N_12869);
nor U13179 (N_13179,N_12830,N_12940);
nor U13180 (N_13180,N_12852,N_12884);
nor U13181 (N_13181,N_12839,N_12917);
nor U13182 (N_13182,N_12880,N_12884);
xnor U13183 (N_13183,N_12935,N_12844);
nand U13184 (N_13184,N_12813,N_12979);
or U13185 (N_13185,N_12841,N_12892);
and U13186 (N_13186,N_12946,N_12927);
and U13187 (N_13187,N_12890,N_12843);
or U13188 (N_13188,N_12816,N_12938);
nand U13189 (N_13189,N_12920,N_12825);
xnor U13190 (N_13190,N_12823,N_12999);
and U13191 (N_13191,N_12804,N_12890);
and U13192 (N_13192,N_12838,N_12889);
nand U13193 (N_13193,N_12916,N_12894);
xnor U13194 (N_13194,N_12807,N_12927);
xnor U13195 (N_13195,N_12854,N_12876);
nand U13196 (N_13196,N_12897,N_12845);
and U13197 (N_13197,N_12816,N_12993);
nand U13198 (N_13198,N_12961,N_12924);
nor U13199 (N_13199,N_12886,N_12965);
nand U13200 (N_13200,N_13153,N_13045);
and U13201 (N_13201,N_13093,N_13151);
xor U13202 (N_13202,N_13092,N_13184);
or U13203 (N_13203,N_13021,N_13169);
nand U13204 (N_13204,N_13103,N_13076);
xnor U13205 (N_13205,N_13071,N_13055);
nand U13206 (N_13206,N_13126,N_13105);
or U13207 (N_13207,N_13161,N_13121);
nand U13208 (N_13208,N_13175,N_13008);
xnor U13209 (N_13209,N_13051,N_13172);
xnor U13210 (N_13210,N_13022,N_13028);
or U13211 (N_13211,N_13174,N_13159);
and U13212 (N_13212,N_13050,N_13111);
nand U13213 (N_13213,N_13043,N_13006);
xor U13214 (N_13214,N_13130,N_13143);
xnor U13215 (N_13215,N_13192,N_13033);
and U13216 (N_13216,N_13134,N_13181);
nand U13217 (N_13217,N_13041,N_13189);
nand U13218 (N_13218,N_13069,N_13199);
or U13219 (N_13219,N_13053,N_13019);
nand U13220 (N_13220,N_13039,N_13048);
xnor U13221 (N_13221,N_13080,N_13142);
xor U13222 (N_13222,N_13099,N_13162);
xnor U13223 (N_13223,N_13003,N_13074);
or U13224 (N_13224,N_13070,N_13165);
nand U13225 (N_13225,N_13179,N_13046);
xor U13226 (N_13226,N_13096,N_13187);
xor U13227 (N_13227,N_13110,N_13135);
nor U13228 (N_13228,N_13095,N_13060);
xnor U13229 (N_13229,N_13047,N_13035);
xnor U13230 (N_13230,N_13023,N_13198);
or U13231 (N_13231,N_13029,N_13073);
nor U13232 (N_13232,N_13145,N_13088);
nand U13233 (N_13233,N_13131,N_13078);
or U13234 (N_13234,N_13077,N_13156);
or U13235 (N_13235,N_13090,N_13166);
xnor U13236 (N_13236,N_13109,N_13018);
and U13237 (N_13237,N_13102,N_13177);
xnor U13238 (N_13238,N_13180,N_13101);
nor U13239 (N_13239,N_13042,N_13144);
nand U13240 (N_13240,N_13004,N_13157);
xnor U13241 (N_13241,N_13072,N_13167);
or U13242 (N_13242,N_13170,N_13122);
or U13243 (N_13243,N_13136,N_13016);
xnor U13244 (N_13244,N_13138,N_13061);
nor U13245 (N_13245,N_13067,N_13191);
or U13246 (N_13246,N_13062,N_13186);
nand U13247 (N_13247,N_13007,N_13085);
xnor U13248 (N_13248,N_13010,N_13112);
xor U13249 (N_13249,N_13097,N_13066);
and U13250 (N_13250,N_13098,N_13068);
or U13251 (N_13251,N_13148,N_13087);
nand U13252 (N_13252,N_13183,N_13012);
nor U13253 (N_13253,N_13123,N_13064);
nor U13254 (N_13254,N_13094,N_13149);
xor U13255 (N_13255,N_13147,N_13132);
and U13256 (N_13256,N_13027,N_13056);
nor U13257 (N_13257,N_13158,N_13196);
xnor U13258 (N_13258,N_13188,N_13049);
or U13259 (N_13259,N_13185,N_13163);
nand U13260 (N_13260,N_13089,N_13015);
nand U13261 (N_13261,N_13063,N_13057);
nand U13262 (N_13262,N_13036,N_13020);
xor U13263 (N_13263,N_13114,N_13178);
nor U13264 (N_13264,N_13024,N_13150);
nand U13265 (N_13265,N_13082,N_13037);
nor U13266 (N_13266,N_13083,N_13116);
or U13267 (N_13267,N_13002,N_13118);
nand U13268 (N_13268,N_13017,N_13030);
and U13269 (N_13269,N_13104,N_13164);
or U13270 (N_13270,N_13034,N_13173);
and U13271 (N_13271,N_13044,N_13058);
and U13272 (N_13272,N_13091,N_13154);
nor U13273 (N_13273,N_13107,N_13125);
and U13274 (N_13274,N_13059,N_13106);
xnor U13275 (N_13275,N_13026,N_13124);
and U13276 (N_13276,N_13075,N_13128);
nand U13277 (N_13277,N_13054,N_13160);
xor U13278 (N_13278,N_13137,N_13100);
and U13279 (N_13279,N_13079,N_13190);
nor U13280 (N_13280,N_13146,N_13168);
nor U13281 (N_13281,N_13171,N_13176);
or U13282 (N_13282,N_13113,N_13009);
or U13283 (N_13283,N_13140,N_13032);
and U13284 (N_13284,N_13013,N_13139);
nor U13285 (N_13285,N_13197,N_13084);
or U13286 (N_13286,N_13052,N_13001);
or U13287 (N_13287,N_13194,N_13193);
and U13288 (N_13288,N_13108,N_13115);
nor U13289 (N_13289,N_13127,N_13195);
nor U13290 (N_13290,N_13040,N_13065);
or U13291 (N_13291,N_13155,N_13086);
nand U13292 (N_13292,N_13129,N_13011);
and U13293 (N_13293,N_13133,N_13119);
or U13294 (N_13294,N_13152,N_13117);
and U13295 (N_13295,N_13038,N_13182);
or U13296 (N_13296,N_13031,N_13000);
xor U13297 (N_13297,N_13141,N_13014);
or U13298 (N_13298,N_13005,N_13025);
and U13299 (N_13299,N_13120,N_13081);
nor U13300 (N_13300,N_13037,N_13070);
nand U13301 (N_13301,N_13046,N_13075);
nor U13302 (N_13302,N_13187,N_13192);
nor U13303 (N_13303,N_13158,N_13178);
or U13304 (N_13304,N_13162,N_13041);
and U13305 (N_13305,N_13041,N_13028);
nor U13306 (N_13306,N_13145,N_13007);
and U13307 (N_13307,N_13154,N_13057);
and U13308 (N_13308,N_13143,N_13037);
nor U13309 (N_13309,N_13102,N_13123);
and U13310 (N_13310,N_13058,N_13155);
xnor U13311 (N_13311,N_13150,N_13124);
xnor U13312 (N_13312,N_13123,N_13098);
xor U13313 (N_13313,N_13126,N_13155);
xnor U13314 (N_13314,N_13168,N_13067);
or U13315 (N_13315,N_13008,N_13034);
or U13316 (N_13316,N_13061,N_13082);
xor U13317 (N_13317,N_13136,N_13188);
xor U13318 (N_13318,N_13122,N_13159);
and U13319 (N_13319,N_13070,N_13155);
xor U13320 (N_13320,N_13142,N_13131);
nor U13321 (N_13321,N_13018,N_13007);
or U13322 (N_13322,N_13135,N_13122);
nand U13323 (N_13323,N_13170,N_13097);
or U13324 (N_13324,N_13057,N_13029);
nor U13325 (N_13325,N_13007,N_13173);
nand U13326 (N_13326,N_13016,N_13010);
nor U13327 (N_13327,N_13017,N_13160);
and U13328 (N_13328,N_13130,N_13117);
xor U13329 (N_13329,N_13022,N_13123);
or U13330 (N_13330,N_13113,N_13004);
nor U13331 (N_13331,N_13052,N_13121);
nand U13332 (N_13332,N_13180,N_13008);
nor U13333 (N_13333,N_13055,N_13076);
nor U13334 (N_13334,N_13198,N_13095);
nand U13335 (N_13335,N_13184,N_13014);
or U13336 (N_13336,N_13089,N_13124);
and U13337 (N_13337,N_13066,N_13169);
xnor U13338 (N_13338,N_13032,N_13081);
nand U13339 (N_13339,N_13111,N_13087);
and U13340 (N_13340,N_13188,N_13097);
or U13341 (N_13341,N_13125,N_13084);
xnor U13342 (N_13342,N_13077,N_13018);
xor U13343 (N_13343,N_13139,N_13006);
and U13344 (N_13344,N_13040,N_13164);
or U13345 (N_13345,N_13131,N_13003);
or U13346 (N_13346,N_13095,N_13018);
nand U13347 (N_13347,N_13005,N_13039);
and U13348 (N_13348,N_13010,N_13158);
nor U13349 (N_13349,N_13077,N_13129);
or U13350 (N_13350,N_13129,N_13007);
or U13351 (N_13351,N_13158,N_13118);
and U13352 (N_13352,N_13076,N_13068);
nand U13353 (N_13353,N_13120,N_13052);
xor U13354 (N_13354,N_13184,N_13074);
and U13355 (N_13355,N_13184,N_13197);
nor U13356 (N_13356,N_13148,N_13104);
or U13357 (N_13357,N_13149,N_13000);
or U13358 (N_13358,N_13193,N_13182);
nor U13359 (N_13359,N_13012,N_13049);
nor U13360 (N_13360,N_13129,N_13168);
and U13361 (N_13361,N_13178,N_13171);
nor U13362 (N_13362,N_13155,N_13193);
nand U13363 (N_13363,N_13155,N_13001);
nor U13364 (N_13364,N_13105,N_13027);
nor U13365 (N_13365,N_13105,N_13065);
nor U13366 (N_13366,N_13176,N_13078);
nand U13367 (N_13367,N_13138,N_13115);
or U13368 (N_13368,N_13166,N_13065);
and U13369 (N_13369,N_13197,N_13026);
nand U13370 (N_13370,N_13173,N_13041);
xnor U13371 (N_13371,N_13109,N_13113);
or U13372 (N_13372,N_13198,N_13166);
xnor U13373 (N_13373,N_13175,N_13182);
xor U13374 (N_13374,N_13041,N_13072);
xor U13375 (N_13375,N_13107,N_13031);
and U13376 (N_13376,N_13170,N_13168);
or U13377 (N_13377,N_13020,N_13074);
and U13378 (N_13378,N_13071,N_13083);
nand U13379 (N_13379,N_13039,N_13070);
nand U13380 (N_13380,N_13029,N_13094);
and U13381 (N_13381,N_13009,N_13048);
or U13382 (N_13382,N_13161,N_13044);
nand U13383 (N_13383,N_13089,N_13197);
xor U13384 (N_13384,N_13074,N_13142);
or U13385 (N_13385,N_13182,N_13016);
and U13386 (N_13386,N_13024,N_13136);
xnor U13387 (N_13387,N_13024,N_13149);
or U13388 (N_13388,N_13021,N_13052);
nand U13389 (N_13389,N_13008,N_13142);
xnor U13390 (N_13390,N_13199,N_13098);
xor U13391 (N_13391,N_13036,N_13197);
and U13392 (N_13392,N_13178,N_13073);
nand U13393 (N_13393,N_13047,N_13188);
nor U13394 (N_13394,N_13156,N_13141);
xnor U13395 (N_13395,N_13091,N_13025);
nand U13396 (N_13396,N_13160,N_13037);
nor U13397 (N_13397,N_13062,N_13197);
nor U13398 (N_13398,N_13184,N_13076);
nor U13399 (N_13399,N_13020,N_13150);
xor U13400 (N_13400,N_13263,N_13387);
or U13401 (N_13401,N_13319,N_13378);
nor U13402 (N_13402,N_13362,N_13363);
nor U13403 (N_13403,N_13380,N_13222);
xor U13404 (N_13404,N_13262,N_13251);
xnor U13405 (N_13405,N_13257,N_13352);
nand U13406 (N_13406,N_13287,N_13364);
nor U13407 (N_13407,N_13342,N_13366);
xnor U13408 (N_13408,N_13269,N_13204);
and U13409 (N_13409,N_13312,N_13389);
xor U13410 (N_13410,N_13397,N_13235);
or U13411 (N_13411,N_13355,N_13255);
nand U13412 (N_13412,N_13246,N_13375);
nand U13413 (N_13413,N_13340,N_13323);
xnor U13414 (N_13414,N_13330,N_13327);
or U13415 (N_13415,N_13360,N_13325);
xnor U13416 (N_13416,N_13374,N_13245);
and U13417 (N_13417,N_13335,N_13234);
or U13418 (N_13418,N_13253,N_13357);
xor U13419 (N_13419,N_13259,N_13386);
and U13420 (N_13420,N_13280,N_13268);
nand U13421 (N_13421,N_13256,N_13293);
xor U13422 (N_13422,N_13314,N_13345);
xor U13423 (N_13423,N_13365,N_13379);
and U13424 (N_13424,N_13336,N_13205);
or U13425 (N_13425,N_13281,N_13200);
or U13426 (N_13426,N_13326,N_13244);
or U13427 (N_13427,N_13265,N_13332);
nand U13428 (N_13428,N_13271,N_13228);
nor U13429 (N_13429,N_13396,N_13288);
xor U13430 (N_13430,N_13213,N_13267);
and U13431 (N_13431,N_13347,N_13224);
nand U13432 (N_13432,N_13295,N_13368);
and U13433 (N_13433,N_13381,N_13308);
and U13434 (N_13434,N_13392,N_13286);
nand U13435 (N_13435,N_13320,N_13382);
nor U13436 (N_13436,N_13284,N_13359);
or U13437 (N_13437,N_13328,N_13261);
nor U13438 (N_13438,N_13220,N_13349);
and U13439 (N_13439,N_13338,N_13292);
xor U13440 (N_13440,N_13249,N_13348);
nor U13441 (N_13441,N_13217,N_13302);
xnor U13442 (N_13442,N_13232,N_13337);
nor U13443 (N_13443,N_13350,N_13305);
nand U13444 (N_13444,N_13260,N_13210);
nor U13445 (N_13445,N_13294,N_13277);
and U13446 (N_13446,N_13273,N_13208);
nor U13447 (N_13447,N_13377,N_13339);
or U13448 (N_13448,N_13231,N_13384);
or U13449 (N_13449,N_13229,N_13290);
or U13450 (N_13450,N_13300,N_13258);
nor U13451 (N_13451,N_13317,N_13206);
nor U13452 (N_13452,N_13272,N_13343);
and U13453 (N_13453,N_13236,N_13264);
and U13454 (N_13454,N_13225,N_13282);
or U13455 (N_13455,N_13369,N_13313);
nand U13456 (N_13456,N_13270,N_13278);
xnor U13457 (N_13457,N_13391,N_13331);
xor U13458 (N_13458,N_13209,N_13356);
or U13459 (N_13459,N_13315,N_13226);
xnor U13460 (N_13460,N_13247,N_13289);
or U13461 (N_13461,N_13285,N_13201);
nand U13462 (N_13462,N_13393,N_13341);
nand U13463 (N_13463,N_13301,N_13309);
and U13464 (N_13464,N_13283,N_13351);
xnor U13465 (N_13465,N_13321,N_13250);
and U13466 (N_13466,N_13371,N_13223);
xor U13467 (N_13467,N_13304,N_13346);
and U13468 (N_13468,N_13358,N_13388);
nor U13469 (N_13469,N_13334,N_13214);
xor U13470 (N_13470,N_13203,N_13344);
or U13471 (N_13471,N_13394,N_13227);
xnor U13472 (N_13472,N_13252,N_13310);
nor U13473 (N_13473,N_13212,N_13395);
or U13474 (N_13474,N_13298,N_13316);
xor U13475 (N_13475,N_13297,N_13275);
or U13476 (N_13476,N_13291,N_13221);
nand U13477 (N_13477,N_13324,N_13274);
xor U13478 (N_13478,N_13373,N_13353);
nand U13479 (N_13479,N_13202,N_13254);
or U13480 (N_13480,N_13299,N_13311);
and U13481 (N_13481,N_13329,N_13215);
or U13482 (N_13482,N_13239,N_13306);
or U13483 (N_13483,N_13207,N_13242);
nand U13484 (N_13484,N_13211,N_13279);
nor U13485 (N_13485,N_13376,N_13398);
xnor U13486 (N_13486,N_13390,N_13333);
xor U13487 (N_13487,N_13303,N_13399);
and U13488 (N_13488,N_13385,N_13216);
or U13489 (N_13489,N_13238,N_13248);
nor U13490 (N_13490,N_13361,N_13230);
and U13491 (N_13491,N_13243,N_13237);
nand U13492 (N_13492,N_13354,N_13276);
nand U13493 (N_13493,N_13233,N_13219);
nor U13494 (N_13494,N_13318,N_13370);
or U13495 (N_13495,N_13383,N_13372);
xnor U13496 (N_13496,N_13322,N_13307);
or U13497 (N_13497,N_13266,N_13367);
xor U13498 (N_13498,N_13218,N_13241);
xor U13499 (N_13499,N_13240,N_13296);
nand U13500 (N_13500,N_13265,N_13202);
nand U13501 (N_13501,N_13253,N_13378);
nand U13502 (N_13502,N_13372,N_13290);
xnor U13503 (N_13503,N_13394,N_13255);
nor U13504 (N_13504,N_13392,N_13343);
nand U13505 (N_13505,N_13325,N_13397);
and U13506 (N_13506,N_13380,N_13297);
nor U13507 (N_13507,N_13337,N_13328);
xor U13508 (N_13508,N_13211,N_13264);
nor U13509 (N_13509,N_13291,N_13290);
nand U13510 (N_13510,N_13361,N_13319);
nor U13511 (N_13511,N_13297,N_13388);
xor U13512 (N_13512,N_13274,N_13323);
and U13513 (N_13513,N_13377,N_13244);
and U13514 (N_13514,N_13285,N_13258);
nand U13515 (N_13515,N_13362,N_13270);
xor U13516 (N_13516,N_13254,N_13346);
nand U13517 (N_13517,N_13216,N_13208);
or U13518 (N_13518,N_13219,N_13235);
or U13519 (N_13519,N_13247,N_13321);
and U13520 (N_13520,N_13347,N_13266);
xor U13521 (N_13521,N_13298,N_13225);
and U13522 (N_13522,N_13337,N_13338);
and U13523 (N_13523,N_13243,N_13318);
nand U13524 (N_13524,N_13240,N_13336);
or U13525 (N_13525,N_13380,N_13291);
nor U13526 (N_13526,N_13297,N_13369);
and U13527 (N_13527,N_13362,N_13227);
nand U13528 (N_13528,N_13296,N_13274);
xnor U13529 (N_13529,N_13335,N_13253);
and U13530 (N_13530,N_13263,N_13221);
xor U13531 (N_13531,N_13307,N_13324);
and U13532 (N_13532,N_13378,N_13286);
and U13533 (N_13533,N_13271,N_13267);
and U13534 (N_13534,N_13362,N_13374);
nor U13535 (N_13535,N_13239,N_13366);
and U13536 (N_13536,N_13270,N_13352);
and U13537 (N_13537,N_13298,N_13244);
or U13538 (N_13538,N_13355,N_13389);
nand U13539 (N_13539,N_13204,N_13376);
nor U13540 (N_13540,N_13244,N_13367);
and U13541 (N_13541,N_13374,N_13256);
xnor U13542 (N_13542,N_13291,N_13236);
xor U13543 (N_13543,N_13343,N_13341);
and U13544 (N_13544,N_13283,N_13314);
nor U13545 (N_13545,N_13369,N_13359);
or U13546 (N_13546,N_13358,N_13367);
and U13547 (N_13547,N_13310,N_13315);
nand U13548 (N_13548,N_13332,N_13390);
nand U13549 (N_13549,N_13314,N_13219);
and U13550 (N_13550,N_13343,N_13399);
or U13551 (N_13551,N_13273,N_13343);
and U13552 (N_13552,N_13380,N_13235);
nand U13553 (N_13553,N_13205,N_13244);
nand U13554 (N_13554,N_13214,N_13388);
or U13555 (N_13555,N_13264,N_13262);
or U13556 (N_13556,N_13297,N_13323);
nand U13557 (N_13557,N_13279,N_13245);
nor U13558 (N_13558,N_13330,N_13394);
nor U13559 (N_13559,N_13201,N_13255);
nor U13560 (N_13560,N_13281,N_13305);
xor U13561 (N_13561,N_13358,N_13393);
nor U13562 (N_13562,N_13302,N_13316);
nand U13563 (N_13563,N_13346,N_13230);
and U13564 (N_13564,N_13283,N_13324);
and U13565 (N_13565,N_13283,N_13378);
nand U13566 (N_13566,N_13207,N_13302);
xor U13567 (N_13567,N_13234,N_13206);
or U13568 (N_13568,N_13364,N_13204);
xnor U13569 (N_13569,N_13283,N_13349);
nand U13570 (N_13570,N_13307,N_13229);
nand U13571 (N_13571,N_13253,N_13390);
xnor U13572 (N_13572,N_13376,N_13381);
xor U13573 (N_13573,N_13292,N_13283);
xnor U13574 (N_13574,N_13341,N_13240);
nor U13575 (N_13575,N_13307,N_13345);
nor U13576 (N_13576,N_13226,N_13245);
nand U13577 (N_13577,N_13212,N_13295);
nor U13578 (N_13578,N_13314,N_13386);
xnor U13579 (N_13579,N_13351,N_13252);
xnor U13580 (N_13580,N_13290,N_13227);
xor U13581 (N_13581,N_13359,N_13356);
xnor U13582 (N_13582,N_13257,N_13260);
and U13583 (N_13583,N_13369,N_13392);
xnor U13584 (N_13584,N_13203,N_13354);
nor U13585 (N_13585,N_13304,N_13311);
or U13586 (N_13586,N_13248,N_13314);
nor U13587 (N_13587,N_13359,N_13354);
nand U13588 (N_13588,N_13276,N_13291);
nand U13589 (N_13589,N_13344,N_13393);
nor U13590 (N_13590,N_13296,N_13267);
xor U13591 (N_13591,N_13391,N_13277);
or U13592 (N_13592,N_13317,N_13256);
nand U13593 (N_13593,N_13360,N_13296);
or U13594 (N_13594,N_13291,N_13344);
or U13595 (N_13595,N_13205,N_13316);
and U13596 (N_13596,N_13309,N_13246);
nand U13597 (N_13597,N_13398,N_13305);
nor U13598 (N_13598,N_13220,N_13334);
or U13599 (N_13599,N_13395,N_13390);
xnor U13600 (N_13600,N_13490,N_13485);
xnor U13601 (N_13601,N_13572,N_13592);
nand U13602 (N_13602,N_13440,N_13400);
nor U13603 (N_13603,N_13560,N_13570);
and U13604 (N_13604,N_13564,N_13503);
nand U13605 (N_13605,N_13526,N_13532);
or U13606 (N_13606,N_13553,N_13457);
nand U13607 (N_13607,N_13595,N_13416);
and U13608 (N_13608,N_13468,N_13434);
xor U13609 (N_13609,N_13475,N_13489);
xnor U13610 (N_13610,N_13427,N_13548);
nand U13611 (N_13611,N_13589,N_13533);
xor U13612 (N_13612,N_13537,N_13536);
nor U13613 (N_13613,N_13588,N_13497);
and U13614 (N_13614,N_13477,N_13576);
nor U13615 (N_13615,N_13422,N_13513);
nor U13616 (N_13616,N_13462,N_13574);
and U13617 (N_13617,N_13585,N_13445);
nor U13618 (N_13618,N_13478,N_13542);
xor U13619 (N_13619,N_13569,N_13586);
nand U13620 (N_13620,N_13549,N_13556);
nand U13621 (N_13621,N_13522,N_13410);
nand U13622 (N_13622,N_13500,N_13419);
and U13623 (N_13623,N_13438,N_13428);
nand U13624 (N_13624,N_13402,N_13568);
nor U13625 (N_13625,N_13412,N_13535);
or U13626 (N_13626,N_13442,N_13559);
and U13627 (N_13627,N_13429,N_13431);
or U13628 (N_13628,N_13470,N_13528);
and U13629 (N_13629,N_13437,N_13571);
nand U13630 (N_13630,N_13447,N_13448);
xor U13631 (N_13631,N_13558,N_13599);
or U13632 (N_13632,N_13492,N_13474);
or U13633 (N_13633,N_13488,N_13544);
and U13634 (N_13634,N_13481,N_13540);
and U13635 (N_13635,N_13552,N_13527);
and U13636 (N_13636,N_13543,N_13529);
and U13637 (N_13637,N_13405,N_13517);
or U13638 (N_13638,N_13596,N_13458);
nand U13639 (N_13639,N_13509,N_13487);
and U13640 (N_13640,N_13551,N_13463);
xor U13641 (N_13641,N_13515,N_13578);
xor U13642 (N_13642,N_13483,N_13584);
and U13643 (N_13643,N_13521,N_13464);
nand U13644 (N_13644,N_13461,N_13456);
and U13645 (N_13645,N_13441,N_13494);
or U13646 (N_13646,N_13491,N_13444);
xnor U13647 (N_13647,N_13591,N_13538);
nand U13648 (N_13648,N_13414,N_13415);
nor U13649 (N_13649,N_13547,N_13505);
nor U13650 (N_13650,N_13486,N_13580);
xor U13651 (N_13651,N_13453,N_13508);
xnor U13652 (N_13652,N_13484,N_13598);
and U13653 (N_13653,N_13546,N_13413);
and U13654 (N_13654,N_13401,N_13476);
nand U13655 (N_13655,N_13451,N_13561);
or U13656 (N_13656,N_13582,N_13480);
nand U13657 (N_13657,N_13421,N_13423);
nor U13658 (N_13658,N_13573,N_13449);
nor U13659 (N_13659,N_13443,N_13417);
nor U13660 (N_13660,N_13432,N_13408);
nand U13661 (N_13661,N_13499,N_13469);
xnor U13662 (N_13662,N_13436,N_13473);
or U13663 (N_13663,N_13563,N_13404);
nand U13664 (N_13664,N_13587,N_13541);
and U13665 (N_13665,N_13554,N_13518);
nand U13666 (N_13666,N_13465,N_13493);
nor U13667 (N_13667,N_13454,N_13459);
or U13668 (N_13668,N_13472,N_13594);
or U13669 (N_13669,N_13496,N_13575);
nand U13670 (N_13670,N_13426,N_13498);
and U13671 (N_13671,N_13501,N_13504);
and U13672 (N_13672,N_13420,N_13525);
xnor U13673 (N_13673,N_13524,N_13403);
nor U13674 (N_13674,N_13577,N_13507);
nand U13675 (N_13675,N_13450,N_13479);
or U13676 (N_13676,N_13516,N_13424);
xor U13677 (N_13677,N_13567,N_13466);
xor U13678 (N_13678,N_13531,N_13555);
or U13679 (N_13679,N_13520,N_13562);
xnor U13680 (N_13680,N_13467,N_13510);
xnor U13681 (N_13681,N_13455,N_13439);
nand U13682 (N_13682,N_13523,N_13593);
and U13683 (N_13683,N_13425,N_13579);
and U13684 (N_13684,N_13597,N_13506);
nand U13685 (N_13685,N_13435,N_13590);
nand U13686 (N_13686,N_13482,N_13512);
and U13687 (N_13687,N_13565,N_13583);
and U13688 (N_13688,N_13550,N_13495);
and U13689 (N_13689,N_13539,N_13519);
and U13690 (N_13690,N_13411,N_13530);
xor U13691 (N_13691,N_13452,N_13502);
nand U13692 (N_13692,N_13433,N_13446);
and U13693 (N_13693,N_13581,N_13407);
or U13694 (N_13694,N_13545,N_13418);
nand U13695 (N_13695,N_13566,N_13534);
or U13696 (N_13696,N_13406,N_13409);
xnor U13697 (N_13697,N_13514,N_13557);
and U13698 (N_13698,N_13511,N_13430);
and U13699 (N_13699,N_13460,N_13471);
nand U13700 (N_13700,N_13548,N_13510);
nand U13701 (N_13701,N_13428,N_13527);
nand U13702 (N_13702,N_13581,N_13481);
or U13703 (N_13703,N_13428,N_13419);
and U13704 (N_13704,N_13526,N_13412);
nand U13705 (N_13705,N_13549,N_13463);
nand U13706 (N_13706,N_13432,N_13414);
xor U13707 (N_13707,N_13494,N_13422);
nor U13708 (N_13708,N_13427,N_13518);
and U13709 (N_13709,N_13531,N_13456);
and U13710 (N_13710,N_13555,N_13556);
xor U13711 (N_13711,N_13484,N_13567);
and U13712 (N_13712,N_13451,N_13534);
nand U13713 (N_13713,N_13412,N_13476);
or U13714 (N_13714,N_13594,N_13488);
xnor U13715 (N_13715,N_13531,N_13458);
nand U13716 (N_13716,N_13548,N_13535);
nor U13717 (N_13717,N_13529,N_13468);
nand U13718 (N_13718,N_13456,N_13442);
or U13719 (N_13719,N_13484,N_13429);
nand U13720 (N_13720,N_13422,N_13520);
nand U13721 (N_13721,N_13571,N_13436);
nor U13722 (N_13722,N_13559,N_13594);
nor U13723 (N_13723,N_13520,N_13498);
nand U13724 (N_13724,N_13519,N_13594);
or U13725 (N_13725,N_13428,N_13422);
xor U13726 (N_13726,N_13400,N_13587);
nor U13727 (N_13727,N_13579,N_13444);
or U13728 (N_13728,N_13583,N_13499);
xor U13729 (N_13729,N_13417,N_13537);
and U13730 (N_13730,N_13484,N_13582);
nor U13731 (N_13731,N_13475,N_13403);
or U13732 (N_13732,N_13486,N_13442);
nand U13733 (N_13733,N_13406,N_13543);
and U13734 (N_13734,N_13413,N_13572);
nand U13735 (N_13735,N_13412,N_13513);
xor U13736 (N_13736,N_13483,N_13486);
or U13737 (N_13737,N_13589,N_13415);
and U13738 (N_13738,N_13554,N_13567);
nand U13739 (N_13739,N_13558,N_13566);
or U13740 (N_13740,N_13478,N_13544);
xnor U13741 (N_13741,N_13599,N_13424);
or U13742 (N_13742,N_13449,N_13438);
or U13743 (N_13743,N_13436,N_13581);
xor U13744 (N_13744,N_13456,N_13532);
nand U13745 (N_13745,N_13577,N_13553);
and U13746 (N_13746,N_13498,N_13583);
nor U13747 (N_13747,N_13447,N_13584);
or U13748 (N_13748,N_13554,N_13537);
or U13749 (N_13749,N_13421,N_13499);
nand U13750 (N_13750,N_13538,N_13459);
and U13751 (N_13751,N_13507,N_13518);
and U13752 (N_13752,N_13469,N_13536);
or U13753 (N_13753,N_13488,N_13464);
and U13754 (N_13754,N_13566,N_13543);
or U13755 (N_13755,N_13561,N_13448);
nor U13756 (N_13756,N_13456,N_13565);
nor U13757 (N_13757,N_13415,N_13465);
xnor U13758 (N_13758,N_13406,N_13423);
or U13759 (N_13759,N_13578,N_13513);
xor U13760 (N_13760,N_13581,N_13446);
and U13761 (N_13761,N_13478,N_13561);
nor U13762 (N_13762,N_13402,N_13508);
nor U13763 (N_13763,N_13462,N_13431);
nor U13764 (N_13764,N_13558,N_13586);
nor U13765 (N_13765,N_13444,N_13479);
nand U13766 (N_13766,N_13521,N_13411);
nor U13767 (N_13767,N_13512,N_13476);
or U13768 (N_13768,N_13482,N_13456);
nor U13769 (N_13769,N_13505,N_13551);
nor U13770 (N_13770,N_13428,N_13456);
or U13771 (N_13771,N_13511,N_13586);
nor U13772 (N_13772,N_13568,N_13416);
xor U13773 (N_13773,N_13564,N_13400);
or U13774 (N_13774,N_13550,N_13585);
nand U13775 (N_13775,N_13571,N_13585);
and U13776 (N_13776,N_13568,N_13555);
or U13777 (N_13777,N_13413,N_13405);
nand U13778 (N_13778,N_13551,N_13567);
and U13779 (N_13779,N_13428,N_13570);
xor U13780 (N_13780,N_13523,N_13572);
and U13781 (N_13781,N_13479,N_13552);
nand U13782 (N_13782,N_13480,N_13599);
and U13783 (N_13783,N_13566,N_13492);
or U13784 (N_13784,N_13544,N_13510);
or U13785 (N_13785,N_13588,N_13508);
or U13786 (N_13786,N_13489,N_13591);
and U13787 (N_13787,N_13595,N_13464);
nand U13788 (N_13788,N_13525,N_13459);
xor U13789 (N_13789,N_13576,N_13575);
nand U13790 (N_13790,N_13506,N_13521);
or U13791 (N_13791,N_13489,N_13452);
nand U13792 (N_13792,N_13411,N_13586);
nand U13793 (N_13793,N_13503,N_13485);
or U13794 (N_13794,N_13501,N_13502);
nor U13795 (N_13795,N_13452,N_13469);
or U13796 (N_13796,N_13540,N_13412);
or U13797 (N_13797,N_13512,N_13526);
nand U13798 (N_13798,N_13405,N_13522);
and U13799 (N_13799,N_13590,N_13514);
nor U13800 (N_13800,N_13790,N_13720);
nand U13801 (N_13801,N_13641,N_13614);
nor U13802 (N_13802,N_13677,N_13687);
nor U13803 (N_13803,N_13681,N_13606);
xnor U13804 (N_13804,N_13635,N_13650);
xnor U13805 (N_13805,N_13730,N_13691);
xnor U13806 (N_13806,N_13715,N_13658);
nand U13807 (N_13807,N_13620,N_13666);
nor U13808 (N_13808,N_13762,N_13798);
nand U13809 (N_13809,N_13741,N_13604);
nand U13810 (N_13810,N_13724,N_13622);
or U13811 (N_13811,N_13646,N_13752);
and U13812 (N_13812,N_13655,N_13678);
or U13813 (N_13813,N_13776,N_13638);
and U13814 (N_13814,N_13653,N_13686);
nor U13815 (N_13815,N_13605,N_13700);
xor U13816 (N_13816,N_13772,N_13656);
xnor U13817 (N_13817,N_13789,N_13795);
or U13818 (N_13818,N_13727,N_13777);
xor U13819 (N_13819,N_13703,N_13663);
and U13820 (N_13820,N_13702,N_13694);
xor U13821 (N_13821,N_13639,N_13749);
and U13822 (N_13822,N_13626,N_13657);
and U13823 (N_13823,N_13661,N_13654);
or U13824 (N_13824,N_13609,N_13721);
and U13825 (N_13825,N_13615,N_13644);
and U13826 (N_13826,N_13796,N_13685);
or U13827 (N_13827,N_13610,N_13698);
nand U13828 (N_13828,N_13643,N_13710);
nor U13829 (N_13829,N_13787,N_13695);
nor U13830 (N_13830,N_13769,N_13765);
or U13831 (N_13831,N_13679,N_13764);
nand U13832 (N_13832,N_13726,N_13770);
xor U13833 (N_13833,N_13775,N_13779);
nand U13834 (N_13834,N_13692,N_13759);
nor U13835 (N_13835,N_13688,N_13709);
nand U13836 (N_13836,N_13608,N_13744);
or U13837 (N_13837,N_13723,N_13766);
nand U13838 (N_13838,N_13725,N_13745);
nand U13839 (N_13839,N_13746,N_13781);
xnor U13840 (N_13840,N_13649,N_13793);
and U13841 (N_13841,N_13672,N_13637);
nor U13842 (N_13842,N_13755,N_13631);
or U13843 (N_13843,N_13717,N_13768);
or U13844 (N_13844,N_13645,N_13624);
nand U13845 (N_13845,N_13739,N_13734);
or U13846 (N_13846,N_13674,N_13716);
nor U13847 (N_13847,N_13712,N_13665);
and U13848 (N_13848,N_13785,N_13659);
or U13849 (N_13849,N_13611,N_13774);
nor U13850 (N_13850,N_13690,N_13636);
or U13851 (N_13851,N_13601,N_13680);
xnor U13852 (N_13852,N_13640,N_13751);
or U13853 (N_13853,N_13782,N_13621);
nand U13854 (N_13854,N_13760,N_13699);
or U13855 (N_13855,N_13705,N_13794);
and U13856 (N_13856,N_13667,N_13767);
nor U13857 (N_13857,N_13792,N_13756);
nand U13858 (N_13858,N_13761,N_13758);
and U13859 (N_13859,N_13728,N_13634);
nor U13860 (N_13860,N_13607,N_13706);
xnor U13861 (N_13861,N_13673,N_13708);
xnor U13862 (N_13862,N_13729,N_13733);
nand U13863 (N_13863,N_13757,N_13763);
xor U13864 (N_13864,N_13651,N_13754);
and U13865 (N_13865,N_13625,N_13753);
nor U13866 (N_13866,N_13786,N_13642);
or U13867 (N_13867,N_13740,N_13603);
and U13868 (N_13868,N_13684,N_13696);
or U13869 (N_13869,N_13662,N_13616);
nand U13870 (N_13870,N_13736,N_13675);
xnor U13871 (N_13871,N_13633,N_13683);
and U13872 (N_13872,N_13619,N_13647);
and U13873 (N_13873,N_13697,N_13784);
nand U13874 (N_13874,N_13718,N_13788);
and U13875 (N_13875,N_13618,N_13670);
nor U13876 (N_13876,N_13773,N_13738);
xor U13877 (N_13877,N_13799,N_13735);
nand U13878 (N_13878,N_13797,N_13693);
or U13879 (N_13879,N_13689,N_13630);
nand U13880 (N_13880,N_13748,N_13707);
xnor U13881 (N_13881,N_13676,N_13791);
nand U13882 (N_13882,N_13719,N_13771);
and U13883 (N_13883,N_13722,N_13743);
or U13884 (N_13884,N_13737,N_13742);
xnor U13885 (N_13885,N_13652,N_13783);
and U13886 (N_13886,N_13617,N_13731);
nor U13887 (N_13887,N_13623,N_13632);
or U13888 (N_13888,N_13732,N_13714);
nor U13889 (N_13889,N_13668,N_13648);
nand U13890 (N_13890,N_13612,N_13780);
nor U13891 (N_13891,N_13669,N_13704);
nor U13892 (N_13892,N_13602,N_13627);
or U13893 (N_13893,N_13713,N_13747);
and U13894 (N_13894,N_13628,N_13682);
xor U13895 (N_13895,N_13613,N_13664);
xor U13896 (N_13896,N_13701,N_13711);
and U13897 (N_13897,N_13671,N_13629);
or U13898 (N_13898,N_13778,N_13600);
xor U13899 (N_13899,N_13660,N_13750);
or U13900 (N_13900,N_13712,N_13737);
xnor U13901 (N_13901,N_13620,N_13710);
nor U13902 (N_13902,N_13780,N_13663);
or U13903 (N_13903,N_13746,N_13649);
and U13904 (N_13904,N_13712,N_13762);
or U13905 (N_13905,N_13684,N_13705);
or U13906 (N_13906,N_13745,N_13677);
nor U13907 (N_13907,N_13785,N_13758);
xor U13908 (N_13908,N_13635,N_13768);
nand U13909 (N_13909,N_13624,N_13718);
nand U13910 (N_13910,N_13674,N_13608);
nand U13911 (N_13911,N_13758,N_13798);
and U13912 (N_13912,N_13608,N_13630);
xnor U13913 (N_13913,N_13617,N_13771);
or U13914 (N_13914,N_13638,N_13782);
nor U13915 (N_13915,N_13655,N_13669);
and U13916 (N_13916,N_13786,N_13762);
xnor U13917 (N_13917,N_13652,N_13784);
nand U13918 (N_13918,N_13652,N_13600);
nor U13919 (N_13919,N_13647,N_13780);
or U13920 (N_13920,N_13620,N_13655);
or U13921 (N_13921,N_13660,N_13721);
and U13922 (N_13922,N_13634,N_13777);
nor U13923 (N_13923,N_13703,N_13687);
or U13924 (N_13924,N_13692,N_13730);
xor U13925 (N_13925,N_13639,N_13681);
or U13926 (N_13926,N_13622,N_13700);
and U13927 (N_13927,N_13635,N_13737);
nor U13928 (N_13928,N_13722,N_13667);
nand U13929 (N_13929,N_13608,N_13621);
and U13930 (N_13930,N_13775,N_13705);
nor U13931 (N_13931,N_13707,N_13670);
or U13932 (N_13932,N_13708,N_13624);
nand U13933 (N_13933,N_13680,N_13623);
nand U13934 (N_13934,N_13728,N_13720);
nand U13935 (N_13935,N_13649,N_13680);
nor U13936 (N_13936,N_13770,N_13616);
xor U13937 (N_13937,N_13631,N_13665);
nand U13938 (N_13938,N_13611,N_13622);
or U13939 (N_13939,N_13663,N_13611);
or U13940 (N_13940,N_13770,N_13684);
nor U13941 (N_13941,N_13782,N_13760);
or U13942 (N_13942,N_13627,N_13609);
xnor U13943 (N_13943,N_13755,N_13691);
xnor U13944 (N_13944,N_13651,N_13748);
nand U13945 (N_13945,N_13761,N_13655);
xnor U13946 (N_13946,N_13707,N_13661);
xor U13947 (N_13947,N_13682,N_13619);
and U13948 (N_13948,N_13693,N_13614);
nor U13949 (N_13949,N_13783,N_13727);
or U13950 (N_13950,N_13743,N_13666);
nor U13951 (N_13951,N_13761,N_13792);
nor U13952 (N_13952,N_13698,N_13717);
nor U13953 (N_13953,N_13704,N_13656);
xnor U13954 (N_13954,N_13743,N_13797);
nor U13955 (N_13955,N_13681,N_13657);
xnor U13956 (N_13956,N_13783,N_13738);
and U13957 (N_13957,N_13642,N_13756);
nand U13958 (N_13958,N_13739,N_13608);
nor U13959 (N_13959,N_13752,N_13643);
nor U13960 (N_13960,N_13723,N_13666);
xnor U13961 (N_13961,N_13710,N_13664);
and U13962 (N_13962,N_13742,N_13735);
nor U13963 (N_13963,N_13645,N_13633);
or U13964 (N_13964,N_13631,N_13781);
xor U13965 (N_13965,N_13711,N_13732);
and U13966 (N_13966,N_13757,N_13616);
and U13967 (N_13967,N_13658,N_13718);
xor U13968 (N_13968,N_13766,N_13620);
or U13969 (N_13969,N_13633,N_13638);
or U13970 (N_13970,N_13723,N_13798);
or U13971 (N_13971,N_13778,N_13656);
xnor U13972 (N_13972,N_13744,N_13680);
or U13973 (N_13973,N_13608,N_13668);
nand U13974 (N_13974,N_13628,N_13727);
xnor U13975 (N_13975,N_13626,N_13622);
nand U13976 (N_13976,N_13770,N_13745);
and U13977 (N_13977,N_13700,N_13635);
or U13978 (N_13978,N_13776,N_13607);
or U13979 (N_13979,N_13637,N_13706);
nand U13980 (N_13980,N_13614,N_13665);
or U13981 (N_13981,N_13758,N_13717);
and U13982 (N_13982,N_13705,N_13757);
nor U13983 (N_13983,N_13778,N_13744);
xor U13984 (N_13984,N_13660,N_13643);
or U13985 (N_13985,N_13723,N_13709);
xor U13986 (N_13986,N_13784,N_13798);
xnor U13987 (N_13987,N_13716,N_13647);
nor U13988 (N_13988,N_13768,N_13712);
and U13989 (N_13989,N_13642,N_13652);
nor U13990 (N_13990,N_13697,N_13769);
xnor U13991 (N_13991,N_13696,N_13669);
or U13992 (N_13992,N_13676,N_13760);
and U13993 (N_13993,N_13614,N_13791);
nor U13994 (N_13994,N_13785,N_13771);
xor U13995 (N_13995,N_13603,N_13751);
and U13996 (N_13996,N_13690,N_13649);
nor U13997 (N_13997,N_13618,N_13653);
or U13998 (N_13998,N_13651,N_13673);
or U13999 (N_13999,N_13751,N_13718);
xor U14000 (N_14000,N_13955,N_13994);
nand U14001 (N_14001,N_13917,N_13876);
or U14002 (N_14002,N_13993,N_13805);
nor U14003 (N_14003,N_13818,N_13830);
or U14004 (N_14004,N_13940,N_13868);
or U14005 (N_14005,N_13862,N_13922);
nand U14006 (N_14006,N_13971,N_13861);
xor U14007 (N_14007,N_13816,N_13803);
nand U14008 (N_14008,N_13867,N_13991);
nand U14009 (N_14009,N_13884,N_13938);
or U14010 (N_14010,N_13820,N_13918);
or U14011 (N_14011,N_13945,N_13964);
nor U14012 (N_14012,N_13927,N_13978);
xnor U14013 (N_14013,N_13970,N_13848);
nor U14014 (N_14014,N_13969,N_13972);
xnor U14015 (N_14015,N_13929,N_13941);
xnor U14016 (N_14016,N_13801,N_13845);
nor U14017 (N_14017,N_13959,N_13892);
xnor U14018 (N_14018,N_13921,N_13985);
nor U14019 (N_14019,N_13809,N_13881);
or U14020 (N_14020,N_13998,N_13897);
xor U14021 (N_14021,N_13873,N_13937);
or U14022 (N_14022,N_13857,N_13953);
nand U14023 (N_14023,N_13914,N_13939);
and U14024 (N_14024,N_13883,N_13996);
or U14025 (N_14025,N_13986,N_13808);
xnor U14026 (N_14026,N_13850,N_13880);
or U14027 (N_14027,N_13858,N_13979);
nor U14028 (N_14028,N_13948,N_13891);
nand U14029 (N_14029,N_13823,N_13981);
or U14030 (N_14030,N_13854,N_13901);
xor U14031 (N_14031,N_13821,N_13859);
xor U14032 (N_14032,N_13874,N_13842);
xnor U14033 (N_14033,N_13839,N_13961);
nand U14034 (N_14034,N_13912,N_13987);
xnor U14035 (N_14035,N_13844,N_13966);
nand U14036 (N_14036,N_13967,N_13957);
or U14037 (N_14037,N_13852,N_13944);
and U14038 (N_14038,N_13907,N_13846);
and U14039 (N_14039,N_13815,N_13942);
or U14040 (N_14040,N_13806,N_13962);
and U14041 (N_14041,N_13832,N_13887);
nor U14042 (N_14042,N_13824,N_13886);
xor U14043 (N_14043,N_13895,N_13877);
nand U14044 (N_14044,N_13995,N_13817);
or U14045 (N_14045,N_13870,N_13951);
nor U14046 (N_14046,N_13826,N_13829);
and U14047 (N_14047,N_13807,N_13980);
or U14048 (N_14048,N_13889,N_13843);
xnor U14049 (N_14049,N_13977,N_13952);
nand U14050 (N_14050,N_13804,N_13975);
and U14051 (N_14051,N_13838,N_13882);
or U14052 (N_14052,N_13903,N_13813);
and U14053 (N_14053,N_13812,N_13949);
nand U14054 (N_14054,N_13930,N_13871);
or U14055 (N_14055,N_13860,N_13849);
xnor U14056 (N_14056,N_13822,N_13866);
xor U14057 (N_14057,N_13934,N_13811);
xor U14058 (N_14058,N_13865,N_13932);
nand U14059 (N_14059,N_13896,N_13828);
and U14060 (N_14060,N_13974,N_13894);
xor U14061 (N_14061,N_13802,N_13847);
nor U14062 (N_14062,N_13915,N_13919);
or U14063 (N_14063,N_13827,N_13879);
and U14064 (N_14064,N_13968,N_13923);
nand U14065 (N_14065,N_13936,N_13837);
nand U14066 (N_14066,N_13810,N_13956);
and U14067 (N_14067,N_13913,N_13825);
nor U14068 (N_14068,N_13911,N_13988);
nor U14069 (N_14069,N_13946,N_13885);
xor U14070 (N_14070,N_13890,N_13954);
nand U14071 (N_14071,N_13872,N_13965);
xnor U14072 (N_14072,N_13836,N_13989);
nor U14073 (N_14073,N_13833,N_13910);
nor U14074 (N_14074,N_13931,N_13983);
and U14075 (N_14075,N_13899,N_13909);
and U14076 (N_14076,N_13943,N_13982);
xnor U14077 (N_14077,N_13841,N_13898);
or U14078 (N_14078,N_13875,N_13999);
xor U14079 (N_14079,N_13906,N_13947);
nor U14080 (N_14080,N_13904,N_13990);
or U14081 (N_14081,N_13976,N_13960);
nor U14082 (N_14082,N_13900,N_13851);
and U14083 (N_14083,N_13935,N_13834);
nand U14084 (N_14084,N_13997,N_13878);
nand U14085 (N_14085,N_13819,N_13925);
nor U14086 (N_14086,N_13908,N_13924);
nand U14087 (N_14087,N_13926,N_13863);
or U14088 (N_14088,N_13840,N_13864);
xnor U14089 (N_14089,N_13835,N_13855);
xor U14090 (N_14090,N_13831,N_13916);
nor U14091 (N_14091,N_13893,N_13928);
xnor U14092 (N_14092,N_13963,N_13888);
nand U14093 (N_14093,N_13853,N_13950);
nand U14094 (N_14094,N_13984,N_13800);
nor U14095 (N_14095,N_13992,N_13958);
or U14096 (N_14096,N_13856,N_13814);
nand U14097 (N_14097,N_13920,N_13869);
or U14098 (N_14098,N_13933,N_13905);
nand U14099 (N_14099,N_13973,N_13902);
or U14100 (N_14100,N_13810,N_13865);
nor U14101 (N_14101,N_13857,N_13883);
xnor U14102 (N_14102,N_13934,N_13868);
or U14103 (N_14103,N_13944,N_13835);
or U14104 (N_14104,N_13957,N_13800);
and U14105 (N_14105,N_13835,N_13800);
and U14106 (N_14106,N_13924,N_13917);
xnor U14107 (N_14107,N_13846,N_13871);
xnor U14108 (N_14108,N_13925,N_13982);
nor U14109 (N_14109,N_13813,N_13840);
nor U14110 (N_14110,N_13924,N_13843);
and U14111 (N_14111,N_13894,N_13969);
nor U14112 (N_14112,N_13952,N_13967);
nor U14113 (N_14113,N_13900,N_13846);
nor U14114 (N_14114,N_13898,N_13988);
nor U14115 (N_14115,N_13863,N_13885);
xor U14116 (N_14116,N_13847,N_13911);
nand U14117 (N_14117,N_13823,N_13841);
and U14118 (N_14118,N_13894,N_13983);
or U14119 (N_14119,N_13848,N_13959);
or U14120 (N_14120,N_13858,N_13883);
nor U14121 (N_14121,N_13806,N_13827);
and U14122 (N_14122,N_13885,N_13935);
xnor U14123 (N_14123,N_13989,N_13944);
or U14124 (N_14124,N_13890,N_13846);
nor U14125 (N_14125,N_13836,N_13985);
or U14126 (N_14126,N_13885,N_13920);
and U14127 (N_14127,N_13847,N_13905);
and U14128 (N_14128,N_13864,N_13832);
xor U14129 (N_14129,N_13983,N_13943);
nor U14130 (N_14130,N_13957,N_13876);
or U14131 (N_14131,N_13912,N_13989);
and U14132 (N_14132,N_13976,N_13989);
and U14133 (N_14133,N_13889,N_13808);
or U14134 (N_14134,N_13825,N_13802);
nand U14135 (N_14135,N_13802,N_13875);
or U14136 (N_14136,N_13885,N_13984);
xor U14137 (N_14137,N_13879,N_13838);
xor U14138 (N_14138,N_13988,N_13886);
nor U14139 (N_14139,N_13967,N_13827);
and U14140 (N_14140,N_13823,N_13893);
xnor U14141 (N_14141,N_13954,N_13862);
nand U14142 (N_14142,N_13845,N_13872);
xor U14143 (N_14143,N_13925,N_13949);
xnor U14144 (N_14144,N_13913,N_13855);
nand U14145 (N_14145,N_13869,N_13900);
nand U14146 (N_14146,N_13904,N_13868);
or U14147 (N_14147,N_13862,N_13848);
and U14148 (N_14148,N_13970,N_13914);
nor U14149 (N_14149,N_13892,N_13812);
or U14150 (N_14150,N_13875,N_13925);
or U14151 (N_14151,N_13874,N_13945);
or U14152 (N_14152,N_13822,N_13883);
nand U14153 (N_14153,N_13949,N_13883);
or U14154 (N_14154,N_13947,N_13824);
and U14155 (N_14155,N_13891,N_13833);
or U14156 (N_14156,N_13846,N_13984);
or U14157 (N_14157,N_13883,N_13809);
nand U14158 (N_14158,N_13906,N_13951);
nand U14159 (N_14159,N_13824,N_13924);
and U14160 (N_14160,N_13968,N_13977);
nor U14161 (N_14161,N_13864,N_13855);
nor U14162 (N_14162,N_13828,N_13972);
xnor U14163 (N_14163,N_13815,N_13877);
or U14164 (N_14164,N_13900,N_13994);
or U14165 (N_14165,N_13843,N_13931);
or U14166 (N_14166,N_13984,N_13829);
and U14167 (N_14167,N_13861,N_13941);
nand U14168 (N_14168,N_13975,N_13925);
nand U14169 (N_14169,N_13897,N_13921);
and U14170 (N_14170,N_13887,N_13976);
or U14171 (N_14171,N_13819,N_13874);
and U14172 (N_14172,N_13958,N_13892);
xor U14173 (N_14173,N_13873,N_13953);
nor U14174 (N_14174,N_13969,N_13929);
nand U14175 (N_14175,N_13936,N_13981);
xor U14176 (N_14176,N_13803,N_13936);
xnor U14177 (N_14177,N_13992,N_13861);
xnor U14178 (N_14178,N_13940,N_13824);
and U14179 (N_14179,N_13899,N_13926);
nand U14180 (N_14180,N_13961,N_13941);
or U14181 (N_14181,N_13890,N_13832);
or U14182 (N_14182,N_13835,N_13878);
and U14183 (N_14183,N_13918,N_13845);
or U14184 (N_14184,N_13908,N_13937);
and U14185 (N_14185,N_13958,N_13969);
and U14186 (N_14186,N_13909,N_13912);
xnor U14187 (N_14187,N_13884,N_13838);
and U14188 (N_14188,N_13987,N_13865);
nor U14189 (N_14189,N_13908,N_13948);
or U14190 (N_14190,N_13896,N_13885);
xnor U14191 (N_14191,N_13863,N_13946);
xor U14192 (N_14192,N_13937,N_13938);
nand U14193 (N_14193,N_13838,N_13934);
or U14194 (N_14194,N_13911,N_13863);
nor U14195 (N_14195,N_13929,N_13821);
or U14196 (N_14196,N_13924,N_13994);
xor U14197 (N_14197,N_13994,N_13977);
nand U14198 (N_14198,N_13896,N_13854);
or U14199 (N_14199,N_13856,N_13967);
or U14200 (N_14200,N_14035,N_14016);
xor U14201 (N_14201,N_14169,N_14181);
or U14202 (N_14202,N_14052,N_14094);
xor U14203 (N_14203,N_14160,N_14021);
or U14204 (N_14204,N_14147,N_14004);
nand U14205 (N_14205,N_14174,N_14034);
nor U14206 (N_14206,N_14099,N_14100);
xnor U14207 (N_14207,N_14042,N_14136);
nand U14208 (N_14208,N_14180,N_14003);
nor U14209 (N_14209,N_14159,N_14071);
and U14210 (N_14210,N_14111,N_14166);
nand U14211 (N_14211,N_14113,N_14010);
nor U14212 (N_14212,N_14092,N_14055);
or U14213 (N_14213,N_14152,N_14183);
and U14214 (N_14214,N_14109,N_14038);
and U14215 (N_14215,N_14137,N_14048);
and U14216 (N_14216,N_14050,N_14000);
nand U14217 (N_14217,N_14150,N_14128);
and U14218 (N_14218,N_14184,N_14197);
or U14219 (N_14219,N_14198,N_14008);
and U14220 (N_14220,N_14122,N_14025);
nor U14221 (N_14221,N_14193,N_14001);
or U14222 (N_14222,N_14154,N_14187);
and U14223 (N_14223,N_14095,N_14015);
nand U14224 (N_14224,N_14027,N_14081);
and U14225 (N_14225,N_14097,N_14143);
xnor U14226 (N_14226,N_14098,N_14108);
nand U14227 (N_14227,N_14129,N_14040);
nand U14228 (N_14228,N_14101,N_14170);
or U14229 (N_14229,N_14089,N_14120);
nor U14230 (N_14230,N_14104,N_14188);
and U14231 (N_14231,N_14033,N_14088);
xnor U14232 (N_14232,N_14086,N_14085);
or U14233 (N_14233,N_14141,N_14131);
or U14234 (N_14234,N_14106,N_14165);
xnor U14235 (N_14235,N_14047,N_14151);
and U14236 (N_14236,N_14041,N_14162);
xnor U14237 (N_14237,N_14102,N_14032);
xnor U14238 (N_14238,N_14069,N_14191);
or U14239 (N_14239,N_14103,N_14065);
nand U14240 (N_14240,N_14144,N_14167);
nor U14241 (N_14241,N_14118,N_14028);
or U14242 (N_14242,N_14133,N_14115);
or U14243 (N_14243,N_14186,N_14096);
nand U14244 (N_14244,N_14067,N_14145);
nor U14245 (N_14245,N_14070,N_14164);
nand U14246 (N_14246,N_14138,N_14139);
nor U14247 (N_14247,N_14177,N_14124);
and U14248 (N_14248,N_14084,N_14037);
xor U14249 (N_14249,N_14049,N_14132);
or U14250 (N_14250,N_14146,N_14107);
nor U14251 (N_14251,N_14013,N_14182);
or U14252 (N_14252,N_14073,N_14026);
nand U14253 (N_14253,N_14022,N_14168);
xor U14254 (N_14254,N_14024,N_14017);
xnor U14255 (N_14255,N_14123,N_14056);
or U14256 (N_14256,N_14005,N_14199);
xnor U14257 (N_14257,N_14019,N_14029);
nor U14258 (N_14258,N_14135,N_14121);
and U14259 (N_14259,N_14061,N_14030);
xnor U14260 (N_14260,N_14007,N_14062);
nand U14261 (N_14261,N_14006,N_14023);
nor U14262 (N_14262,N_14196,N_14105);
xor U14263 (N_14263,N_14114,N_14173);
xnor U14264 (N_14264,N_14077,N_14045);
xor U14265 (N_14265,N_14155,N_14063);
nor U14266 (N_14266,N_14059,N_14074);
or U14267 (N_14267,N_14011,N_14009);
and U14268 (N_14268,N_14171,N_14161);
nand U14269 (N_14269,N_14014,N_14082);
xnor U14270 (N_14270,N_14153,N_14054);
and U14271 (N_14271,N_14051,N_14090);
and U14272 (N_14272,N_14190,N_14116);
nand U14273 (N_14273,N_14148,N_14179);
xnor U14274 (N_14274,N_14158,N_14057);
and U14275 (N_14275,N_14046,N_14080);
or U14276 (N_14276,N_14189,N_14087);
nand U14277 (N_14277,N_14119,N_14036);
and U14278 (N_14278,N_14002,N_14110);
xnor U14279 (N_14279,N_14068,N_14093);
nor U14280 (N_14280,N_14163,N_14142);
nand U14281 (N_14281,N_14156,N_14018);
and U14282 (N_14282,N_14172,N_14012);
or U14283 (N_14283,N_14064,N_14112);
xor U14284 (N_14284,N_14140,N_14117);
xnor U14285 (N_14285,N_14178,N_14149);
nand U14286 (N_14286,N_14130,N_14134);
or U14287 (N_14287,N_14066,N_14058);
nor U14288 (N_14288,N_14091,N_14185);
xnor U14289 (N_14289,N_14039,N_14079);
and U14290 (N_14290,N_14127,N_14020);
nor U14291 (N_14291,N_14075,N_14157);
and U14292 (N_14292,N_14076,N_14125);
nor U14293 (N_14293,N_14194,N_14043);
nand U14294 (N_14294,N_14031,N_14126);
xor U14295 (N_14295,N_14060,N_14175);
or U14296 (N_14296,N_14083,N_14053);
nand U14297 (N_14297,N_14192,N_14044);
xor U14298 (N_14298,N_14072,N_14078);
xor U14299 (N_14299,N_14195,N_14176);
or U14300 (N_14300,N_14014,N_14026);
nor U14301 (N_14301,N_14116,N_14086);
nor U14302 (N_14302,N_14027,N_14151);
and U14303 (N_14303,N_14024,N_14004);
or U14304 (N_14304,N_14127,N_14024);
xor U14305 (N_14305,N_14180,N_14132);
nor U14306 (N_14306,N_14179,N_14121);
nor U14307 (N_14307,N_14173,N_14004);
and U14308 (N_14308,N_14075,N_14048);
nand U14309 (N_14309,N_14135,N_14095);
or U14310 (N_14310,N_14040,N_14116);
or U14311 (N_14311,N_14188,N_14031);
xor U14312 (N_14312,N_14125,N_14194);
and U14313 (N_14313,N_14098,N_14189);
nor U14314 (N_14314,N_14095,N_14124);
and U14315 (N_14315,N_14012,N_14126);
or U14316 (N_14316,N_14136,N_14157);
nor U14317 (N_14317,N_14075,N_14074);
and U14318 (N_14318,N_14033,N_14179);
or U14319 (N_14319,N_14090,N_14093);
or U14320 (N_14320,N_14032,N_14007);
and U14321 (N_14321,N_14002,N_14127);
or U14322 (N_14322,N_14106,N_14075);
xor U14323 (N_14323,N_14102,N_14167);
xnor U14324 (N_14324,N_14143,N_14119);
nand U14325 (N_14325,N_14097,N_14063);
xnor U14326 (N_14326,N_14132,N_14102);
and U14327 (N_14327,N_14170,N_14167);
nand U14328 (N_14328,N_14090,N_14165);
xor U14329 (N_14329,N_14064,N_14137);
and U14330 (N_14330,N_14056,N_14101);
nor U14331 (N_14331,N_14165,N_14042);
nor U14332 (N_14332,N_14166,N_14042);
and U14333 (N_14333,N_14188,N_14128);
or U14334 (N_14334,N_14136,N_14097);
or U14335 (N_14335,N_14052,N_14169);
or U14336 (N_14336,N_14115,N_14130);
and U14337 (N_14337,N_14118,N_14083);
and U14338 (N_14338,N_14043,N_14124);
or U14339 (N_14339,N_14088,N_14147);
xor U14340 (N_14340,N_14018,N_14135);
xnor U14341 (N_14341,N_14111,N_14155);
xnor U14342 (N_14342,N_14159,N_14052);
nand U14343 (N_14343,N_14040,N_14109);
or U14344 (N_14344,N_14136,N_14140);
nor U14345 (N_14345,N_14018,N_14112);
or U14346 (N_14346,N_14003,N_14076);
nand U14347 (N_14347,N_14040,N_14147);
or U14348 (N_14348,N_14159,N_14024);
nand U14349 (N_14349,N_14021,N_14051);
and U14350 (N_14350,N_14045,N_14195);
or U14351 (N_14351,N_14114,N_14166);
and U14352 (N_14352,N_14076,N_14173);
nand U14353 (N_14353,N_14078,N_14142);
and U14354 (N_14354,N_14113,N_14026);
nor U14355 (N_14355,N_14104,N_14047);
nor U14356 (N_14356,N_14170,N_14131);
xnor U14357 (N_14357,N_14155,N_14043);
xor U14358 (N_14358,N_14124,N_14126);
nand U14359 (N_14359,N_14045,N_14196);
or U14360 (N_14360,N_14160,N_14108);
xnor U14361 (N_14361,N_14037,N_14108);
and U14362 (N_14362,N_14080,N_14174);
nor U14363 (N_14363,N_14042,N_14058);
nand U14364 (N_14364,N_14146,N_14065);
xor U14365 (N_14365,N_14138,N_14013);
xnor U14366 (N_14366,N_14165,N_14044);
nand U14367 (N_14367,N_14193,N_14084);
nor U14368 (N_14368,N_14064,N_14020);
nand U14369 (N_14369,N_14110,N_14148);
nand U14370 (N_14370,N_14114,N_14175);
xor U14371 (N_14371,N_14142,N_14173);
nor U14372 (N_14372,N_14075,N_14022);
nand U14373 (N_14373,N_14061,N_14057);
nor U14374 (N_14374,N_14089,N_14158);
and U14375 (N_14375,N_14047,N_14027);
nand U14376 (N_14376,N_14058,N_14030);
and U14377 (N_14377,N_14044,N_14161);
and U14378 (N_14378,N_14189,N_14164);
nor U14379 (N_14379,N_14179,N_14070);
nor U14380 (N_14380,N_14171,N_14087);
xor U14381 (N_14381,N_14129,N_14060);
nor U14382 (N_14382,N_14154,N_14113);
xnor U14383 (N_14383,N_14042,N_14145);
and U14384 (N_14384,N_14129,N_14143);
nor U14385 (N_14385,N_14024,N_14026);
or U14386 (N_14386,N_14189,N_14044);
and U14387 (N_14387,N_14172,N_14184);
or U14388 (N_14388,N_14089,N_14176);
nand U14389 (N_14389,N_14127,N_14164);
and U14390 (N_14390,N_14157,N_14199);
nand U14391 (N_14391,N_14060,N_14165);
and U14392 (N_14392,N_14173,N_14015);
and U14393 (N_14393,N_14132,N_14020);
xor U14394 (N_14394,N_14044,N_14054);
nand U14395 (N_14395,N_14190,N_14021);
xor U14396 (N_14396,N_14124,N_14117);
xnor U14397 (N_14397,N_14196,N_14094);
nand U14398 (N_14398,N_14170,N_14102);
nand U14399 (N_14399,N_14009,N_14099);
or U14400 (N_14400,N_14290,N_14385);
nand U14401 (N_14401,N_14336,N_14393);
or U14402 (N_14402,N_14370,N_14398);
nor U14403 (N_14403,N_14272,N_14225);
nand U14404 (N_14404,N_14217,N_14263);
and U14405 (N_14405,N_14269,N_14325);
xor U14406 (N_14406,N_14208,N_14399);
and U14407 (N_14407,N_14229,N_14331);
or U14408 (N_14408,N_14308,N_14227);
nand U14409 (N_14409,N_14338,N_14224);
or U14410 (N_14410,N_14340,N_14353);
xnor U14411 (N_14411,N_14260,N_14324);
or U14412 (N_14412,N_14350,N_14288);
nor U14413 (N_14413,N_14293,N_14275);
nor U14414 (N_14414,N_14396,N_14239);
and U14415 (N_14415,N_14366,N_14262);
xor U14416 (N_14416,N_14264,N_14332);
nor U14417 (N_14417,N_14236,N_14228);
nor U14418 (N_14418,N_14382,N_14352);
xnor U14419 (N_14419,N_14377,N_14360);
or U14420 (N_14420,N_14329,N_14361);
xor U14421 (N_14421,N_14287,N_14267);
nand U14422 (N_14422,N_14218,N_14342);
xnor U14423 (N_14423,N_14254,N_14315);
or U14424 (N_14424,N_14278,N_14364);
xor U14425 (N_14425,N_14304,N_14265);
nor U14426 (N_14426,N_14257,N_14251);
nor U14427 (N_14427,N_14241,N_14335);
nand U14428 (N_14428,N_14246,N_14348);
or U14429 (N_14429,N_14291,N_14367);
nand U14430 (N_14430,N_14245,N_14298);
nand U14431 (N_14431,N_14242,N_14253);
and U14432 (N_14432,N_14322,N_14333);
nor U14433 (N_14433,N_14365,N_14334);
nor U14434 (N_14434,N_14318,N_14320);
nor U14435 (N_14435,N_14213,N_14294);
xor U14436 (N_14436,N_14295,N_14258);
and U14437 (N_14437,N_14378,N_14391);
xnor U14438 (N_14438,N_14221,N_14238);
and U14439 (N_14439,N_14319,N_14379);
and U14440 (N_14440,N_14235,N_14248);
nor U14441 (N_14441,N_14255,N_14326);
nand U14442 (N_14442,N_14214,N_14202);
and U14443 (N_14443,N_14299,N_14273);
xor U14444 (N_14444,N_14369,N_14292);
xor U14445 (N_14445,N_14330,N_14357);
or U14446 (N_14446,N_14201,N_14368);
nand U14447 (N_14447,N_14309,N_14277);
nor U14448 (N_14448,N_14388,N_14233);
xnor U14449 (N_14449,N_14394,N_14343);
or U14450 (N_14450,N_14328,N_14302);
nand U14451 (N_14451,N_14215,N_14280);
xor U14452 (N_14452,N_14210,N_14313);
or U14453 (N_14453,N_14395,N_14211);
and U14454 (N_14454,N_14386,N_14301);
nor U14455 (N_14455,N_14212,N_14223);
nand U14456 (N_14456,N_14373,N_14363);
or U14457 (N_14457,N_14384,N_14270);
nor U14458 (N_14458,N_14339,N_14204);
nand U14459 (N_14459,N_14314,N_14234);
nor U14460 (N_14460,N_14206,N_14383);
nor U14461 (N_14461,N_14256,N_14200);
xor U14462 (N_14462,N_14327,N_14347);
or U14463 (N_14463,N_14219,N_14250);
and U14464 (N_14464,N_14349,N_14226);
nor U14465 (N_14465,N_14306,N_14310);
or U14466 (N_14466,N_14230,N_14266);
xnor U14467 (N_14467,N_14220,N_14297);
and U14468 (N_14468,N_14358,N_14305);
nand U14469 (N_14469,N_14323,N_14243);
nand U14470 (N_14470,N_14397,N_14286);
xnor U14471 (N_14471,N_14282,N_14312);
or U14472 (N_14472,N_14244,N_14261);
and U14473 (N_14473,N_14346,N_14271);
xor U14474 (N_14474,N_14247,N_14351);
xor U14475 (N_14475,N_14372,N_14259);
xnor U14476 (N_14476,N_14311,N_14289);
nor U14477 (N_14477,N_14205,N_14307);
nand U14478 (N_14478,N_14240,N_14276);
xor U14479 (N_14479,N_14317,N_14376);
and U14480 (N_14480,N_14231,N_14216);
and U14481 (N_14481,N_14296,N_14249);
nor U14482 (N_14482,N_14389,N_14232);
nor U14483 (N_14483,N_14316,N_14283);
or U14484 (N_14484,N_14355,N_14209);
xor U14485 (N_14485,N_14359,N_14321);
nand U14486 (N_14486,N_14285,N_14207);
or U14487 (N_14487,N_14237,N_14274);
xnor U14488 (N_14488,N_14380,N_14268);
nand U14489 (N_14489,N_14300,N_14279);
or U14490 (N_14490,N_14281,N_14341);
xor U14491 (N_14491,N_14381,N_14344);
xnor U14492 (N_14492,N_14362,N_14356);
or U14493 (N_14493,N_14371,N_14390);
nor U14494 (N_14494,N_14303,N_14337);
or U14495 (N_14495,N_14374,N_14222);
and U14496 (N_14496,N_14392,N_14252);
nor U14497 (N_14497,N_14375,N_14345);
xnor U14498 (N_14498,N_14387,N_14284);
nor U14499 (N_14499,N_14354,N_14203);
and U14500 (N_14500,N_14253,N_14352);
or U14501 (N_14501,N_14292,N_14220);
xor U14502 (N_14502,N_14389,N_14314);
xor U14503 (N_14503,N_14221,N_14302);
nand U14504 (N_14504,N_14257,N_14234);
nand U14505 (N_14505,N_14375,N_14381);
xnor U14506 (N_14506,N_14219,N_14282);
nand U14507 (N_14507,N_14368,N_14278);
nor U14508 (N_14508,N_14320,N_14331);
nand U14509 (N_14509,N_14320,N_14204);
or U14510 (N_14510,N_14297,N_14398);
nor U14511 (N_14511,N_14339,N_14255);
and U14512 (N_14512,N_14292,N_14276);
xor U14513 (N_14513,N_14324,N_14243);
and U14514 (N_14514,N_14248,N_14254);
nand U14515 (N_14515,N_14314,N_14270);
nor U14516 (N_14516,N_14226,N_14279);
nor U14517 (N_14517,N_14247,N_14312);
nor U14518 (N_14518,N_14344,N_14238);
nor U14519 (N_14519,N_14384,N_14329);
xnor U14520 (N_14520,N_14269,N_14365);
or U14521 (N_14521,N_14313,N_14301);
and U14522 (N_14522,N_14326,N_14293);
nand U14523 (N_14523,N_14314,N_14332);
nand U14524 (N_14524,N_14312,N_14205);
or U14525 (N_14525,N_14201,N_14309);
or U14526 (N_14526,N_14364,N_14379);
nand U14527 (N_14527,N_14285,N_14312);
nor U14528 (N_14528,N_14226,N_14254);
xor U14529 (N_14529,N_14361,N_14259);
nand U14530 (N_14530,N_14291,N_14362);
or U14531 (N_14531,N_14397,N_14259);
nor U14532 (N_14532,N_14252,N_14309);
nand U14533 (N_14533,N_14302,N_14231);
xnor U14534 (N_14534,N_14251,N_14243);
and U14535 (N_14535,N_14310,N_14336);
nor U14536 (N_14536,N_14314,N_14213);
or U14537 (N_14537,N_14276,N_14311);
or U14538 (N_14538,N_14287,N_14222);
nand U14539 (N_14539,N_14313,N_14212);
and U14540 (N_14540,N_14240,N_14212);
or U14541 (N_14541,N_14220,N_14202);
and U14542 (N_14542,N_14210,N_14331);
nor U14543 (N_14543,N_14393,N_14246);
xnor U14544 (N_14544,N_14350,N_14248);
and U14545 (N_14545,N_14317,N_14394);
nor U14546 (N_14546,N_14339,N_14347);
or U14547 (N_14547,N_14299,N_14308);
nand U14548 (N_14548,N_14285,N_14228);
nor U14549 (N_14549,N_14259,N_14235);
nor U14550 (N_14550,N_14283,N_14279);
and U14551 (N_14551,N_14389,N_14399);
xnor U14552 (N_14552,N_14336,N_14212);
nand U14553 (N_14553,N_14231,N_14298);
and U14554 (N_14554,N_14223,N_14292);
or U14555 (N_14555,N_14320,N_14398);
nand U14556 (N_14556,N_14214,N_14290);
xnor U14557 (N_14557,N_14291,N_14278);
xor U14558 (N_14558,N_14299,N_14356);
nor U14559 (N_14559,N_14308,N_14370);
and U14560 (N_14560,N_14230,N_14264);
or U14561 (N_14561,N_14347,N_14306);
and U14562 (N_14562,N_14221,N_14366);
or U14563 (N_14563,N_14296,N_14374);
nand U14564 (N_14564,N_14290,N_14367);
nor U14565 (N_14565,N_14336,N_14296);
nor U14566 (N_14566,N_14389,N_14243);
and U14567 (N_14567,N_14279,N_14381);
and U14568 (N_14568,N_14200,N_14299);
or U14569 (N_14569,N_14261,N_14386);
or U14570 (N_14570,N_14273,N_14207);
nand U14571 (N_14571,N_14348,N_14290);
or U14572 (N_14572,N_14214,N_14295);
xor U14573 (N_14573,N_14304,N_14201);
xor U14574 (N_14574,N_14249,N_14290);
nand U14575 (N_14575,N_14280,N_14307);
nor U14576 (N_14576,N_14223,N_14377);
nor U14577 (N_14577,N_14365,N_14294);
or U14578 (N_14578,N_14202,N_14200);
nor U14579 (N_14579,N_14302,N_14217);
or U14580 (N_14580,N_14330,N_14210);
and U14581 (N_14581,N_14262,N_14252);
nand U14582 (N_14582,N_14317,N_14255);
and U14583 (N_14583,N_14354,N_14391);
nand U14584 (N_14584,N_14301,N_14305);
nand U14585 (N_14585,N_14260,N_14242);
xnor U14586 (N_14586,N_14292,N_14205);
xor U14587 (N_14587,N_14395,N_14330);
nor U14588 (N_14588,N_14279,N_14332);
and U14589 (N_14589,N_14229,N_14294);
xnor U14590 (N_14590,N_14396,N_14308);
nand U14591 (N_14591,N_14311,N_14339);
or U14592 (N_14592,N_14275,N_14364);
and U14593 (N_14593,N_14280,N_14389);
nand U14594 (N_14594,N_14390,N_14271);
or U14595 (N_14595,N_14399,N_14348);
xor U14596 (N_14596,N_14266,N_14371);
nor U14597 (N_14597,N_14347,N_14246);
nor U14598 (N_14598,N_14373,N_14266);
nor U14599 (N_14599,N_14314,N_14285);
nand U14600 (N_14600,N_14593,N_14414);
nor U14601 (N_14601,N_14521,N_14508);
and U14602 (N_14602,N_14408,N_14570);
nor U14603 (N_14603,N_14440,N_14525);
nand U14604 (N_14604,N_14428,N_14492);
and U14605 (N_14605,N_14595,N_14491);
or U14606 (N_14606,N_14445,N_14466);
or U14607 (N_14607,N_14452,N_14441);
nand U14608 (N_14608,N_14544,N_14415);
nor U14609 (N_14609,N_14580,N_14547);
and U14610 (N_14610,N_14473,N_14465);
xnor U14611 (N_14611,N_14574,N_14454);
xor U14612 (N_14612,N_14424,N_14541);
nor U14613 (N_14613,N_14436,N_14406);
or U14614 (N_14614,N_14497,N_14499);
nand U14615 (N_14615,N_14462,N_14519);
xor U14616 (N_14616,N_14579,N_14439);
nor U14617 (N_14617,N_14422,N_14582);
nand U14618 (N_14618,N_14450,N_14448);
xnor U14619 (N_14619,N_14405,N_14548);
nor U14620 (N_14620,N_14420,N_14494);
nor U14621 (N_14621,N_14487,N_14526);
nor U14622 (N_14622,N_14576,N_14589);
or U14623 (N_14623,N_14455,N_14587);
or U14624 (N_14624,N_14426,N_14460);
nor U14625 (N_14625,N_14532,N_14483);
nor U14626 (N_14626,N_14482,N_14443);
nand U14627 (N_14627,N_14520,N_14588);
or U14628 (N_14628,N_14403,N_14554);
or U14629 (N_14629,N_14513,N_14597);
and U14630 (N_14630,N_14527,N_14502);
nand U14631 (N_14631,N_14505,N_14596);
nor U14632 (N_14632,N_14584,N_14484);
or U14633 (N_14633,N_14549,N_14506);
nand U14634 (N_14634,N_14552,N_14471);
xnor U14635 (N_14635,N_14540,N_14529);
and U14636 (N_14636,N_14539,N_14546);
nor U14637 (N_14637,N_14429,N_14567);
and U14638 (N_14638,N_14457,N_14488);
xnor U14639 (N_14639,N_14495,N_14478);
nor U14640 (N_14640,N_14500,N_14432);
nand U14641 (N_14641,N_14559,N_14400);
or U14642 (N_14642,N_14572,N_14485);
xnor U14643 (N_14643,N_14578,N_14461);
xnor U14644 (N_14644,N_14516,N_14474);
or U14645 (N_14645,N_14594,N_14528);
xnor U14646 (N_14646,N_14509,N_14560);
xnor U14647 (N_14647,N_14561,N_14583);
and U14648 (N_14648,N_14517,N_14430);
and U14649 (N_14649,N_14537,N_14458);
and U14650 (N_14650,N_14586,N_14413);
nand U14651 (N_14651,N_14453,N_14467);
nand U14652 (N_14652,N_14425,N_14514);
xor U14653 (N_14653,N_14459,N_14456);
xor U14654 (N_14654,N_14418,N_14469);
or U14655 (N_14655,N_14598,N_14522);
nand U14656 (N_14656,N_14433,N_14565);
xnor U14657 (N_14657,N_14417,N_14447);
or U14658 (N_14658,N_14479,N_14401);
nand U14659 (N_14659,N_14563,N_14558);
or U14660 (N_14660,N_14562,N_14496);
and U14661 (N_14661,N_14511,N_14556);
xnor U14662 (N_14662,N_14435,N_14470);
or U14663 (N_14663,N_14569,N_14530);
xnor U14664 (N_14664,N_14551,N_14490);
or U14665 (N_14665,N_14591,N_14468);
and U14666 (N_14666,N_14427,N_14524);
nand U14667 (N_14667,N_14477,N_14486);
or U14668 (N_14668,N_14411,N_14564);
and U14669 (N_14669,N_14599,N_14409);
nand U14670 (N_14670,N_14523,N_14553);
nand U14671 (N_14671,N_14498,N_14538);
and U14672 (N_14672,N_14407,N_14442);
nand U14673 (N_14673,N_14416,N_14568);
or U14674 (N_14674,N_14449,N_14423);
nand U14675 (N_14675,N_14481,N_14592);
and U14676 (N_14676,N_14404,N_14590);
nand U14677 (N_14677,N_14534,N_14419);
nor U14678 (N_14678,N_14504,N_14555);
and U14679 (N_14679,N_14431,N_14402);
xor U14680 (N_14680,N_14573,N_14575);
and U14681 (N_14681,N_14434,N_14451);
nor U14682 (N_14682,N_14476,N_14444);
and U14683 (N_14683,N_14437,N_14577);
nor U14684 (N_14684,N_14421,N_14533);
xor U14685 (N_14685,N_14472,N_14493);
xnor U14686 (N_14686,N_14501,N_14531);
xnor U14687 (N_14687,N_14446,N_14412);
nor U14688 (N_14688,N_14581,N_14510);
xor U14689 (N_14689,N_14543,N_14585);
and U14690 (N_14690,N_14475,N_14535);
or U14691 (N_14691,N_14550,N_14463);
xnor U14692 (N_14692,N_14507,N_14542);
nand U14693 (N_14693,N_14545,N_14566);
xnor U14694 (N_14694,N_14464,N_14410);
or U14695 (N_14695,N_14512,N_14480);
nor U14696 (N_14696,N_14518,N_14489);
nand U14697 (N_14697,N_14515,N_14503);
nor U14698 (N_14698,N_14438,N_14557);
and U14699 (N_14699,N_14571,N_14536);
nand U14700 (N_14700,N_14589,N_14567);
nor U14701 (N_14701,N_14561,N_14459);
nand U14702 (N_14702,N_14459,N_14594);
xnor U14703 (N_14703,N_14557,N_14537);
and U14704 (N_14704,N_14462,N_14497);
and U14705 (N_14705,N_14455,N_14431);
or U14706 (N_14706,N_14545,N_14425);
nor U14707 (N_14707,N_14550,N_14578);
xnor U14708 (N_14708,N_14434,N_14588);
and U14709 (N_14709,N_14422,N_14550);
xor U14710 (N_14710,N_14582,N_14522);
nor U14711 (N_14711,N_14461,N_14435);
nand U14712 (N_14712,N_14458,N_14552);
xor U14713 (N_14713,N_14544,N_14481);
nor U14714 (N_14714,N_14420,N_14422);
nor U14715 (N_14715,N_14456,N_14592);
xor U14716 (N_14716,N_14444,N_14553);
nand U14717 (N_14717,N_14541,N_14561);
or U14718 (N_14718,N_14427,N_14567);
or U14719 (N_14719,N_14594,N_14560);
xor U14720 (N_14720,N_14421,N_14597);
and U14721 (N_14721,N_14430,N_14560);
nor U14722 (N_14722,N_14485,N_14438);
nand U14723 (N_14723,N_14457,N_14478);
xor U14724 (N_14724,N_14593,N_14554);
nor U14725 (N_14725,N_14440,N_14490);
xnor U14726 (N_14726,N_14542,N_14419);
xnor U14727 (N_14727,N_14526,N_14559);
and U14728 (N_14728,N_14480,N_14569);
nor U14729 (N_14729,N_14436,N_14442);
nor U14730 (N_14730,N_14411,N_14493);
nor U14731 (N_14731,N_14565,N_14524);
and U14732 (N_14732,N_14402,N_14416);
xnor U14733 (N_14733,N_14541,N_14570);
xor U14734 (N_14734,N_14536,N_14413);
xnor U14735 (N_14735,N_14574,N_14486);
or U14736 (N_14736,N_14503,N_14443);
and U14737 (N_14737,N_14593,N_14422);
nor U14738 (N_14738,N_14590,N_14573);
nor U14739 (N_14739,N_14433,N_14474);
xnor U14740 (N_14740,N_14502,N_14556);
xnor U14741 (N_14741,N_14570,N_14426);
and U14742 (N_14742,N_14420,N_14510);
xnor U14743 (N_14743,N_14408,N_14518);
and U14744 (N_14744,N_14416,N_14410);
nand U14745 (N_14745,N_14452,N_14440);
and U14746 (N_14746,N_14501,N_14511);
xor U14747 (N_14747,N_14554,N_14458);
nor U14748 (N_14748,N_14540,N_14517);
nor U14749 (N_14749,N_14562,N_14435);
xnor U14750 (N_14750,N_14500,N_14536);
nand U14751 (N_14751,N_14418,N_14452);
nand U14752 (N_14752,N_14446,N_14494);
nor U14753 (N_14753,N_14592,N_14563);
nand U14754 (N_14754,N_14557,N_14479);
and U14755 (N_14755,N_14577,N_14403);
xnor U14756 (N_14756,N_14429,N_14500);
and U14757 (N_14757,N_14597,N_14512);
xor U14758 (N_14758,N_14430,N_14400);
nand U14759 (N_14759,N_14515,N_14500);
and U14760 (N_14760,N_14400,N_14539);
nor U14761 (N_14761,N_14461,N_14579);
nor U14762 (N_14762,N_14513,N_14507);
nand U14763 (N_14763,N_14538,N_14450);
xnor U14764 (N_14764,N_14523,N_14504);
or U14765 (N_14765,N_14581,N_14578);
xnor U14766 (N_14766,N_14548,N_14462);
and U14767 (N_14767,N_14408,N_14403);
and U14768 (N_14768,N_14507,N_14502);
and U14769 (N_14769,N_14455,N_14568);
nand U14770 (N_14770,N_14589,N_14596);
or U14771 (N_14771,N_14592,N_14492);
nand U14772 (N_14772,N_14422,N_14584);
xnor U14773 (N_14773,N_14564,N_14591);
and U14774 (N_14774,N_14549,N_14427);
xnor U14775 (N_14775,N_14428,N_14461);
nor U14776 (N_14776,N_14444,N_14526);
or U14777 (N_14777,N_14558,N_14422);
or U14778 (N_14778,N_14410,N_14499);
xor U14779 (N_14779,N_14500,N_14482);
nor U14780 (N_14780,N_14448,N_14462);
nand U14781 (N_14781,N_14496,N_14560);
nand U14782 (N_14782,N_14527,N_14594);
or U14783 (N_14783,N_14412,N_14535);
xnor U14784 (N_14784,N_14405,N_14516);
or U14785 (N_14785,N_14427,N_14544);
nand U14786 (N_14786,N_14545,N_14540);
and U14787 (N_14787,N_14548,N_14586);
nor U14788 (N_14788,N_14432,N_14465);
or U14789 (N_14789,N_14497,N_14474);
nand U14790 (N_14790,N_14406,N_14482);
nand U14791 (N_14791,N_14524,N_14528);
and U14792 (N_14792,N_14468,N_14545);
nor U14793 (N_14793,N_14457,N_14480);
xor U14794 (N_14794,N_14459,N_14457);
nand U14795 (N_14795,N_14517,N_14442);
or U14796 (N_14796,N_14579,N_14423);
and U14797 (N_14797,N_14499,N_14409);
xor U14798 (N_14798,N_14479,N_14485);
and U14799 (N_14799,N_14523,N_14581);
xnor U14800 (N_14800,N_14760,N_14757);
nand U14801 (N_14801,N_14776,N_14603);
or U14802 (N_14802,N_14629,N_14720);
or U14803 (N_14803,N_14735,N_14739);
and U14804 (N_14804,N_14785,N_14786);
nand U14805 (N_14805,N_14714,N_14729);
and U14806 (N_14806,N_14653,N_14655);
or U14807 (N_14807,N_14665,N_14634);
nand U14808 (N_14808,N_14719,N_14738);
nand U14809 (N_14809,N_14633,N_14777);
nand U14810 (N_14810,N_14605,N_14784);
or U14811 (N_14811,N_14708,N_14660);
or U14812 (N_14812,N_14702,N_14610);
nor U14813 (N_14813,N_14798,N_14624);
or U14814 (N_14814,N_14763,N_14761);
or U14815 (N_14815,N_14758,N_14669);
xnor U14816 (N_14816,N_14601,N_14794);
nand U14817 (N_14817,N_14713,N_14766);
nand U14818 (N_14818,N_14716,N_14694);
nand U14819 (N_14819,N_14604,N_14769);
or U14820 (N_14820,N_14683,N_14700);
or U14821 (N_14821,N_14728,N_14613);
or U14822 (N_14822,N_14682,N_14746);
nor U14823 (N_14823,N_14767,N_14711);
nand U14824 (N_14824,N_14636,N_14718);
nor U14825 (N_14825,N_14638,N_14644);
nand U14826 (N_14826,N_14755,N_14759);
or U14827 (N_14827,N_14619,N_14648);
or U14828 (N_14828,N_14689,N_14622);
xor U14829 (N_14829,N_14670,N_14751);
and U14830 (N_14830,N_14641,N_14775);
nand U14831 (N_14831,N_14764,N_14657);
xor U14832 (N_14832,N_14771,N_14640);
nand U14833 (N_14833,N_14611,N_14687);
or U14834 (N_14834,N_14673,N_14676);
xor U14835 (N_14835,N_14632,N_14768);
nor U14836 (N_14836,N_14789,N_14612);
nor U14837 (N_14837,N_14618,N_14787);
and U14838 (N_14838,N_14736,N_14664);
and U14839 (N_14839,N_14643,N_14639);
and U14840 (N_14840,N_14697,N_14795);
nand U14841 (N_14841,N_14745,N_14692);
nor U14842 (N_14842,N_14730,N_14698);
nor U14843 (N_14843,N_14696,N_14725);
nand U14844 (N_14844,N_14734,N_14796);
nand U14845 (N_14845,N_14765,N_14754);
xor U14846 (N_14846,N_14674,N_14680);
and U14847 (N_14847,N_14741,N_14793);
nand U14848 (N_14848,N_14712,N_14790);
and U14849 (N_14849,N_14727,N_14753);
or U14850 (N_14850,N_14666,N_14651);
or U14851 (N_14851,N_14607,N_14600);
nand U14852 (N_14852,N_14617,N_14609);
nor U14853 (N_14853,N_14656,N_14688);
or U14854 (N_14854,N_14742,N_14752);
and U14855 (N_14855,N_14645,N_14606);
nor U14856 (N_14856,N_14732,N_14770);
or U14857 (N_14857,N_14627,N_14699);
nor U14858 (N_14858,N_14748,N_14743);
nand U14859 (N_14859,N_14704,N_14630);
xor U14860 (N_14860,N_14717,N_14783);
or U14861 (N_14861,N_14625,N_14620);
nor U14862 (N_14862,N_14749,N_14703);
nand U14863 (N_14863,N_14671,N_14709);
xnor U14864 (N_14864,N_14681,N_14686);
xnor U14865 (N_14865,N_14721,N_14726);
or U14866 (N_14866,N_14724,N_14637);
nor U14867 (N_14867,N_14661,N_14668);
nor U14868 (N_14868,N_14691,N_14649);
and U14869 (N_14869,N_14706,N_14685);
or U14870 (N_14870,N_14792,N_14733);
nor U14871 (N_14871,N_14652,N_14667);
or U14872 (N_14872,N_14722,N_14780);
nand U14873 (N_14873,N_14690,N_14756);
or U14874 (N_14874,N_14679,N_14662);
xor U14875 (N_14875,N_14762,N_14705);
or U14876 (N_14876,N_14797,N_14778);
and U14877 (N_14877,N_14635,N_14663);
xnor U14878 (N_14878,N_14658,N_14715);
nor U14879 (N_14879,N_14740,N_14747);
xnor U14880 (N_14880,N_14701,N_14650);
nand U14881 (N_14881,N_14621,N_14646);
or U14882 (N_14882,N_14750,N_14731);
nand U14883 (N_14883,N_14602,N_14772);
or U14884 (N_14884,N_14773,N_14737);
and U14885 (N_14885,N_14675,N_14782);
nor U14886 (N_14886,N_14781,N_14774);
or U14887 (N_14887,N_14626,N_14799);
and U14888 (N_14888,N_14677,N_14693);
xor U14889 (N_14889,N_14628,N_14744);
nand U14890 (N_14890,N_14647,N_14779);
nor U14891 (N_14891,N_14723,N_14614);
xor U14892 (N_14892,N_14654,N_14672);
nor U14893 (N_14893,N_14642,N_14678);
xor U14894 (N_14894,N_14616,N_14623);
or U14895 (N_14895,N_14608,N_14788);
xor U14896 (N_14896,N_14631,N_14684);
nor U14897 (N_14897,N_14791,N_14695);
or U14898 (N_14898,N_14707,N_14710);
nor U14899 (N_14899,N_14615,N_14659);
nand U14900 (N_14900,N_14747,N_14721);
nand U14901 (N_14901,N_14757,N_14785);
xnor U14902 (N_14902,N_14774,N_14762);
xor U14903 (N_14903,N_14706,N_14686);
nand U14904 (N_14904,N_14790,N_14738);
nand U14905 (N_14905,N_14761,N_14795);
nor U14906 (N_14906,N_14669,N_14696);
and U14907 (N_14907,N_14776,N_14621);
or U14908 (N_14908,N_14782,N_14603);
and U14909 (N_14909,N_14771,N_14649);
and U14910 (N_14910,N_14633,N_14689);
and U14911 (N_14911,N_14729,N_14643);
nor U14912 (N_14912,N_14697,N_14621);
nor U14913 (N_14913,N_14641,N_14732);
or U14914 (N_14914,N_14742,N_14700);
nand U14915 (N_14915,N_14623,N_14728);
and U14916 (N_14916,N_14786,N_14716);
nand U14917 (N_14917,N_14674,N_14682);
nand U14918 (N_14918,N_14669,N_14742);
nor U14919 (N_14919,N_14686,N_14754);
and U14920 (N_14920,N_14680,N_14725);
nor U14921 (N_14921,N_14684,N_14788);
nor U14922 (N_14922,N_14746,N_14646);
and U14923 (N_14923,N_14609,N_14758);
nor U14924 (N_14924,N_14738,N_14636);
nand U14925 (N_14925,N_14619,N_14660);
or U14926 (N_14926,N_14777,N_14658);
or U14927 (N_14927,N_14790,N_14700);
nor U14928 (N_14928,N_14757,N_14754);
xor U14929 (N_14929,N_14725,N_14701);
or U14930 (N_14930,N_14630,N_14779);
and U14931 (N_14931,N_14720,N_14662);
nor U14932 (N_14932,N_14734,N_14711);
xor U14933 (N_14933,N_14722,N_14625);
xor U14934 (N_14934,N_14615,N_14654);
and U14935 (N_14935,N_14617,N_14727);
xnor U14936 (N_14936,N_14757,N_14746);
nand U14937 (N_14937,N_14603,N_14671);
and U14938 (N_14938,N_14738,N_14616);
nor U14939 (N_14939,N_14675,N_14688);
or U14940 (N_14940,N_14677,N_14618);
nand U14941 (N_14941,N_14711,N_14663);
nand U14942 (N_14942,N_14637,N_14642);
or U14943 (N_14943,N_14741,N_14692);
or U14944 (N_14944,N_14727,N_14749);
xnor U14945 (N_14945,N_14755,N_14722);
nor U14946 (N_14946,N_14707,N_14671);
or U14947 (N_14947,N_14742,N_14711);
xor U14948 (N_14948,N_14777,N_14698);
and U14949 (N_14949,N_14616,N_14673);
nand U14950 (N_14950,N_14671,N_14789);
nand U14951 (N_14951,N_14779,N_14758);
and U14952 (N_14952,N_14680,N_14749);
and U14953 (N_14953,N_14771,N_14634);
or U14954 (N_14954,N_14665,N_14711);
or U14955 (N_14955,N_14613,N_14687);
nand U14956 (N_14956,N_14744,N_14622);
and U14957 (N_14957,N_14668,N_14792);
nand U14958 (N_14958,N_14746,N_14689);
xor U14959 (N_14959,N_14781,N_14621);
nor U14960 (N_14960,N_14775,N_14664);
xnor U14961 (N_14961,N_14608,N_14696);
nor U14962 (N_14962,N_14622,N_14752);
or U14963 (N_14963,N_14734,N_14607);
nand U14964 (N_14964,N_14731,N_14692);
xnor U14965 (N_14965,N_14650,N_14753);
xor U14966 (N_14966,N_14743,N_14608);
xnor U14967 (N_14967,N_14758,N_14718);
xor U14968 (N_14968,N_14744,N_14684);
nand U14969 (N_14969,N_14668,N_14634);
and U14970 (N_14970,N_14715,N_14711);
or U14971 (N_14971,N_14631,N_14794);
xor U14972 (N_14972,N_14731,N_14672);
xnor U14973 (N_14973,N_14615,N_14717);
xor U14974 (N_14974,N_14673,N_14728);
and U14975 (N_14975,N_14675,N_14670);
nor U14976 (N_14976,N_14705,N_14720);
nor U14977 (N_14977,N_14759,N_14646);
nor U14978 (N_14978,N_14676,N_14785);
nor U14979 (N_14979,N_14793,N_14704);
nand U14980 (N_14980,N_14722,N_14621);
and U14981 (N_14981,N_14672,N_14779);
nand U14982 (N_14982,N_14700,N_14783);
xnor U14983 (N_14983,N_14721,N_14724);
nand U14984 (N_14984,N_14625,N_14697);
and U14985 (N_14985,N_14767,N_14695);
nand U14986 (N_14986,N_14773,N_14633);
and U14987 (N_14987,N_14773,N_14625);
or U14988 (N_14988,N_14737,N_14682);
or U14989 (N_14989,N_14718,N_14618);
and U14990 (N_14990,N_14618,N_14771);
or U14991 (N_14991,N_14705,N_14710);
and U14992 (N_14992,N_14772,N_14652);
or U14993 (N_14993,N_14616,N_14798);
and U14994 (N_14994,N_14616,N_14615);
nor U14995 (N_14995,N_14719,N_14654);
xor U14996 (N_14996,N_14660,N_14662);
nand U14997 (N_14997,N_14706,N_14772);
nor U14998 (N_14998,N_14787,N_14619);
or U14999 (N_14999,N_14661,N_14726);
or UO_0 (O_0,N_14950,N_14850);
or UO_1 (O_1,N_14890,N_14999);
xor UO_2 (O_2,N_14897,N_14823);
or UO_3 (O_3,N_14900,N_14936);
nor UO_4 (O_4,N_14948,N_14860);
or UO_5 (O_5,N_14800,N_14868);
xor UO_6 (O_6,N_14966,N_14894);
nor UO_7 (O_7,N_14967,N_14920);
nand UO_8 (O_8,N_14903,N_14910);
or UO_9 (O_9,N_14992,N_14921);
xnor UO_10 (O_10,N_14986,N_14886);
or UO_11 (O_11,N_14958,N_14954);
nor UO_12 (O_12,N_14902,N_14807);
or UO_13 (O_13,N_14804,N_14895);
nor UO_14 (O_14,N_14934,N_14856);
and UO_15 (O_15,N_14922,N_14857);
nor UO_16 (O_16,N_14928,N_14829);
nand UO_17 (O_17,N_14970,N_14963);
nand UO_18 (O_18,N_14861,N_14912);
or UO_19 (O_19,N_14849,N_14991);
and UO_20 (O_20,N_14837,N_14848);
nor UO_21 (O_21,N_14913,N_14918);
or UO_22 (O_22,N_14879,N_14956);
nor UO_23 (O_23,N_14867,N_14833);
and UO_24 (O_24,N_14998,N_14854);
or UO_25 (O_25,N_14847,N_14845);
nand UO_26 (O_26,N_14990,N_14989);
xor UO_27 (O_27,N_14814,N_14806);
xor UO_28 (O_28,N_14839,N_14947);
nor UO_29 (O_29,N_14938,N_14840);
xor UO_30 (O_30,N_14881,N_14968);
and UO_31 (O_31,N_14965,N_14935);
nor UO_32 (O_32,N_14870,N_14831);
or UO_33 (O_33,N_14960,N_14826);
and UO_34 (O_34,N_14951,N_14923);
nor UO_35 (O_35,N_14914,N_14863);
nand UO_36 (O_36,N_14891,N_14859);
nand UO_37 (O_37,N_14997,N_14802);
or UO_38 (O_38,N_14993,N_14979);
xnor UO_39 (O_39,N_14876,N_14952);
nor UO_40 (O_40,N_14904,N_14941);
and UO_41 (O_41,N_14866,N_14961);
nand UO_42 (O_42,N_14855,N_14893);
xor UO_43 (O_43,N_14909,N_14946);
and UO_44 (O_44,N_14932,N_14919);
and UO_45 (O_45,N_14907,N_14885);
xor UO_46 (O_46,N_14996,N_14982);
nor UO_47 (O_47,N_14901,N_14882);
or UO_48 (O_48,N_14873,N_14905);
xnor UO_49 (O_49,N_14875,N_14842);
or UO_50 (O_50,N_14944,N_14887);
nand UO_51 (O_51,N_14988,N_14892);
or UO_52 (O_52,N_14824,N_14813);
or UO_53 (O_53,N_14976,N_14884);
xor UO_54 (O_54,N_14811,N_14880);
nand UO_55 (O_55,N_14836,N_14975);
xor UO_56 (O_56,N_14931,N_14815);
nand UO_57 (O_57,N_14862,N_14852);
xnor UO_58 (O_58,N_14908,N_14825);
nand UO_59 (O_59,N_14980,N_14983);
nor UO_60 (O_60,N_14858,N_14955);
xnor UO_61 (O_61,N_14853,N_14805);
nand UO_62 (O_62,N_14851,N_14820);
and UO_63 (O_63,N_14973,N_14865);
nand UO_64 (O_64,N_14822,N_14972);
and UO_65 (O_65,N_14816,N_14844);
or UO_66 (O_66,N_14911,N_14981);
nor UO_67 (O_67,N_14917,N_14942);
or UO_68 (O_68,N_14812,N_14835);
xor UO_69 (O_69,N_14937,N_14828);
or UO_70 (O_70,N_14916,N_14803);
nor UO_71 (O_71,N_14953,N_14930);
xnor UO_72 (O_72,N_14838,N_14864);
xnor UO_73 (O_73,N_14985,N_14957);
nand UO_74 (O_74,N_14809,N_14821);
or UO_75 (O_75,N_14810,N_14871);
or UO_76 (O_76,N_14827,N_14888);
and UO_77 (O_77,N_14977,N_14915);
and UO_78 (O_78,N_14933,N_14995);
nand UO_79 (O_79,N_14924,N_14818);
nor UO_80 (O_80,N_14878,N_14830);
or UO_81 (O_81,N_14883,N_14846);
nand UO_82 (O_82,N_14945,N_14971);
xnor UO_83 (O_83,N_14899,N_14987);
xnor UO_84 (O_84,N_14808,N_14974);
nor UO_85 (O_85,N_14925,N_14877);
xor UO_86 (O_86,N_14969,N_14926);
nor UO_87 (O_87,N_14943,N_14939);
and UO_88 (O_88,N_14889,N_14841);
and UO_89 (O_89,N_14832,N_14872);
nand UO_90 (O_90,N_14964,N_14959);
or UO_91 (O_91,N_14869,N_14874);
xor UO_92 (O_92,N_14929,N_14819);
or UO_93 (O_93,N_14896,N_14949);
and UO_94 (O_94,N_14962,N_14801);
nor UO_95 (O_95,N_14898,N_14927);
nand UO_96 (O_96,N_14817,N_14940);
nand UO_97 (O_97,N_14843,N_14984);
nand UO_98 (O_98,N_14994,N_14834);
nand UO_99 (O_99,N_14906,N_14978);
xor UO_100 (O_100,N_14840,N_14853);
nand UO_101 (O_101,N_14975,N_14927);
xor UO_102 (O_102,N_14815,N_14915);
xnor UO_103 (O_103,N_14803,N_14918);
nand UO_104 (O_104,N_14867,N_14882);
xor UO_105 (O_105,N_14827,N_14802);
or UO_106 (O_106,N_14863,N_14958);
and UO_107 (O_107,N_14987,N_14935);
nand UO_108 (O_108,N_14953,N_14916);
or UO_109 (O_109,N_14938,N_14965);
or UO_110 (O_110,N_14997,N_14901);
nor UO_111 (O_111,N_14996,N_14902);
nor UO_112 (O_112,N_14810,N_14953);
nand UO_113 (O_113,N_14890,N_14937);
nand UO_114 (O_114,N_14879,N_14814);
or UO_115 (O_115,N_14942,N_14830);
or UO_116 (O_116,N_14951,N_14852);
or UO_117 (O_117,N_14804,N_14915);
nand UO_118 (O_118,N_14896,N_14820);
nor UO_119 (O_119,N_14997,N_14932);
nor UO_120 (O_120,N_14982,N_14814);
nor UO_121 (O_121,N_14880,N_14872);
xnor UO_122 (O_122,N_14825,N_14893);
or UO_123 (O_123,N_14899,N_14921);
or UO_124 (O_124,N_14884,N_14912);
xor UO_125 (O_125,N_14938,N_14873);
nand UO_126 (O_126,N_14933,N_14811);
or UO_127 (O_127,N_14818,N_14856);
xnor UO_128 (O_128,N_14958,N_14857);
nand UO_129 (O_129,N_14835,N_14981);
xor UO_130 (O_130,N_14906,N_14841);
or UO_131 (O_131,N_14810,N_14891);
and UO_132 (O_132,N_14907,N_14866);
nand UO_133 (O_133,N_14868,N_14801);
or UO_134 (O_134,N_14873,N_14872);
nand UO_135 (O_135,N_14855,N_14849);
nand UO_136 (O_136,N_14965,N_14876);
nor UO_137 (O_137,N_14844,N_14951);
or UO_138 (O_138,N_14800,N_14866);
xnor UO_139 (O_139,N_14889,N_14986);
and UO_140 (O_140,N_14960,N_14949);
or UO_141 (O_141,N_14860,N_14982);
nor UO_142 (O_142,N_14986,N_14908);
or UO_143 (O_143,N_14916,N_14996);
nand UO_144 (O_144,N_14862,N_14954);
nand UO_145 (O_145,N_14932,N_14938);
nor UO_146 (O_146,N_14948,N_14966);
nand UO_147 (O_147,N_14931,N_14950);
nand UO_148 (O_148,N_14874,N_14877);
nand UO_149 (O_149,N_14961,N_14892);
xor UO_150 (O_150,N_14978,N_14809);
nor UO_151 (O_151,N_14883,N_14924);
and UO_152 (O_152,N_14949,N_14976);
nor UO_153 (O_153,N_14863,N_14934);
and UO_154 (O_154,N_14947,N_14997);
or UO_155 (O_155,N_14905,N_14997);
or UO_156 (O_156,N_14856,N_14841);
or UO_157 (O_157,N_14908,N_14841);
xnor UO_158 (O_158,N_14912,N_14980);
and UO_159 (O_159,N_14809,N_14813);
nand UO_160 (O_160,N_14950,N_14938);
nand UO_161 (O_161,N_14976,N_14930);
nor UO_162 (O_162,N_14977,N_14897);
and UO_163 (O_163,N_14846,N_14984);
nor UO_164 (O_164,N_14953,N_14909);
and UO_165 (O_165,N_14855,N_14986);
and UO_166 (O_166,N_14872,N_14982);
and UO_167 (O_167,N_14812,N_14984);
xor UO_168 (O_168,N_14867,N_14919);
nand UO_169 (O_169,N_14836,N_14866);
and UO_170 (O_170,N_14809,N_14911);
nand UO_171 (O_171,N_14814,N_14802);
nor UO_172 (O_172,N_14997,N_14972);
or UO_173 (O_173,N_14827,N_14826);
xnor UO_174 (O_174,N_14972,N_14995);
nor UO_175 (O_175,N_14850,N_14806);
and UO_176 (O_176,N_14902,N_14961);
or UO_177 (O_177,N_14878,N_14863);
nor UO_178 (O_178,N_14898,N_14973);
xor UO_179 (O_179,N_14817,N_14801);
nor UO_180 (O_180,N_14885,N_14948);
and UO_181 (O_181,N_14869,N_14837);
nand UO_182 (O_182,N_14818,N_14960);
nand UO_183 (O_183,N_14963,N_14896);
nand UO_184 (O_184,N_14853,N_14966);
xnor UO_185 (O_185,N_14969,N_14824);
and UO_186 (O_186,N_14864,N_14969);
nor UO_187 (O_187,N_14886,N_14927);
nand UO_188 (O_188,N_14843,N_14937);
nand UO_189 (O_189,N_14834,N_14887);
or UO_190 (O_190,N_14990,N_14839);
or UO_191 (O_191,N_14896,N_14816);
xor UO_192 (O_192,N_14830,N_14828);
nand UO_193 (O_193,N_14902,N_14871);
nand UO_194 (O_194,N_14832,N_14901);
or UO_195 (O_195,N_14935,N_14802);
nor UO_196 (O_196,N_14865,N_14800);
nor UO_197 (O_197,N_14809,N_14849);
nand UO_198 (O_198,N_14952,N_14893);
or UO_199 (O_199,N_14907,N_14913);
or UO_200 (O_200,N_14849,N_14847);
or UO_201 (O_201,N_14921,N_14861);
and UO_202 (O_202,N_14976,N_14810);
nand UO_203 (O_203,N_14988,N_14971);
and UO_204 (O_204,N_14933,N_14945);
nor UO_205 (O_205,N_14896,N_14959);
xor UO_206 (O_206,N_14927,N_14909);
nand UO_207 (O_207,N_14873,N_14899);
xor UO_208 (O_208,N_14859,N_14857);
and UO_209 (O_209,N_14986,N_14858);
nor UO_210 (O_210,N_14822,N_14930);
nand UO_211 (O_211,N_14947,N_14883);
xnor UO_212 (O_212,N_14869,N_14884);
and UO_213 (O_213,N_14822,N_14827);
nor UO_214 (O_214,N_14891,N_14861);
nor UO_215 (O_215,N_14883,N_14973);
nand UO_216 (O_216,N_14891,N_14870);
and UO_217 (O_217,N_14998,N_14996);
and UO_218 (O_218,N_14861,N_14808);
nor UO_219 (O_219,N_14863,N_14822);
and UO_220 (O_220,N_14890,N_14936);
and UO_221 (O_221,N_14824,N_14965);
nand UO_222 (O_222,N_14821,N_14810);
or UO_223 (O_223,N_14912,N_14817);
nor UO_224 (O_224,N_14852,N_14985);
nand UO_225 (O_225,N_14962,N_14907);
or UO_226 (O_226,N_14934,N_14956);
and UO_227 (O_227,N_14841,N_14836);
nand UO_228 (O_228,N_14984,N_14968);
nand UO_229 (O_229,N_14845,N_14832);
xnor UO_230 (O_230,N_14995,N_14941);
nor UO_231 (O_231,N_14836,N_14994);
xor UO_232 (O_232,N_14805,N_14847);
xnor UO_233 (O_233,N_14811,N_14949);
or UO_234 (O_234,N_14943,N_14876);
xnor UO_235 (O_235,N_14926,N_14925);
nand UO_236 (O_236,N_14949,N_14898);
nand UO_237 (O_237,N_14804,N_14878);
and UO_238 (O_238,N_14838,N_14975);
nor UO_239 (O_239,N_14826,N_14808);
nor UO_240 (O_240,N_14864,N_14977);
or UO_241 (O_241,N_14993,N_14888);
nor UO_242 (O_242,N_14902,N_14959);
nand UO_243 (O_243,N_14888,N_14979);
or UO_244 (O_244,N_14872,N_14898);
nor UO_245 (O_245,N_14939,N_14991);
nand UO_246 (O_246,N_14924,N_14852);
or UO_247 (O_247,N_14811,N_14938);
nand UO_248 (O_248,N_14964,N_14836);
and UO_249 (O_249,N_14908,N_14901);
nand UO_250 (O_250,N_14949,N_14966);
nand UO_251 (O_251,N_14845,N_14927);
and UO_252 (O_252,N_14950,N_14860);
xor UO_253 (O_253,N_14889,N_14899);
and UO_254 (O_254,N_14918,N_14962);
xnor UO_255 (O_255,N_14948,N_14808);
xnor UO_256 (O_256,N_14894,N_14999);
xor UO_257 (O_257,N_14907,N_14808);
nand UO_258 (O_258,N_14922,N_14935);
xnor UO_259 (O_259,N_14853,N_14886);
and UO_260 (O_260,N_14864,N_14816);
or UO_261 (O_261,N_14834,N_14830);
or UO_262 (O_262,N_14977,N_14816);
or UO_263 (O_263,N_14964,N_14854);
or UO_264 (O_264,N_14975,N_14935);
xnor UO_265 (O_265,N_14905,N_14927);
xnor UO_266 (O_266,N_14952,N_14967);
and UO_267 (O_267,N_14863,N_14933);
or UO_268 (O_268,N_14849,N_14846);
xor UO_269 (O_269,N_14847,N_14873);
and UO_270 (O_270,N_14894,N_14857);
or UO_271 (O_271,N_14924,N_14869);
nand UO_272 (O_272,N_14821,N_14865);
or UO_273 (O_273,N_14811,N_14984);
nand UO_274 (O_274,N_14986,N_14950);
or UO_275 (O_275,N_14865,N_14953);
xor UO_276 (O_276,N_14965,N_14897);
nor UO_277 (O_277,N_14966,N_14898);
and UO_278 (O_278,N_14981,N_14832);
nor UO_279 (O_279,N_14804,N_14824);
xor UO_280 (O_280,N_14954,N_14973);
and UO_281 (O_281,N_14926,N_14867);
or UO_282 (O_282,N_14968,N_14827);
nand UO_283 (O_283,N_14916,N_14906);
and UO_284 (O_284,N_14835,N_14972);
nand UO_285 (O_285,N_14904,N_14857);
nand UO_286 (O_286,N_14846,N_14848);
or UO_287 (O_287,N_14879,N_14815);
and UO_288 (O_288,N_14944,N_14828);
nand UO_289 (O_289,N_14895,N_14982);
and UO_290 (O_290,N_14985,N_14861);
and UO_291 (O_291,N_14853,N_14947);
and UO_292 (O_292,N_14833,N_14935);
nand UO_293 (O_293,N_14963,N_14952);
xnor UO_294 (O_294,N_14949,N_14934);
or UO_295 (O_295,N_14928,N_14855);
and UO_296 (O_296,N_14985,N_14869);
xor UO_297 (O_297,N_14845,N_14980);
xor UO_298 (O_298,N_14906,N_14890);
and UO_299 (O_299,N_14876,N_14823);
xnor UO_300 (O_300,N_14985,N_14848);
or UO_301 (O_301,N_14851,N_14821);
nor UO_302 (O_302,N_14946,N_14837);
or UO_303 (O_303,N_14934,N_14946);
and UO_304 (O_304,N_14847,N_14904);
xor UO_305 (O_305,N_14955,N_14908);
and UO_306 (O_306,N_14831,N_14826);
nor UO_307 (O_307,N_14924,N_14955);
or UO_308 (O_308,N_14952,N_14869);
or UO_309 (O_309,N_14936,N_14977);
and UO_310 (O_310,N_14826,N_14830);
and UO_311 (O_311,N_14896,N_14994);
xnor UO_312 (O_312,N_14824,N_14822);
nand UO_313 (O_313,N_14914,N_14881);
nor UO_314 (O_314,N_14864,N_14988);
and UO_315 (O_315,N_14950,N_14911);
or UO_316 (O_316,N_14959,N_14840);
nand UO_317 (O_317,N_14876,N_14839);
nor UO_318 (O_318,N_14853,N_14999);
xnor UO_319 (O_319,N_14872,N_14907);
nand UO_320 (O_320,N_14996,N_14967);
nand UO_321 (O_321,N_14850,N_14866);
nand UO_322 (O_322,N_14832,N_14950);
nand UO_323 (O_323,N_14883,N_14826);
xor UO_324 (O_324,N_14969,N_14992);
and UO_325 (O_325,N_14815,N_14941);
or UO_326 (O_326,N_14935,N_14840);
nor UO_327 (O_327,N_14929,N_14995);
xnor UO_328 (O_328,N_14889,N_14974);
or UO_329 (O_329,N_14814,N_14997);
xor UO_330 (O_330,N_14836,N_14962);
and UO_331 (O_331,N_14883,N_14874);
nor UO_332 (O_332,N_14818,N_14833);
nand UO_333 (O_333,N_14828,N_14807);
and UO_334 (O_334,N_14869,N_14878);
and UO_335 (O_335,N_14810,N_14986);
nor UO_336 (O_336,N_14847,N_14994);
and UO_337 (O_337,N_14981,N_14861);
nand UO_338 (O_338,N_14854,N_14890);
xnor UO_339 (O_339,N_14987,N_14855);
xnor UO_340 (O_340,N_14953,N_14954);
or UO_341 (O_341,N_14822,N_14995);
and UO_342 (O_342,N_14838,N_14966);
xnor UO_343 (O_343,N_14908,N_14889);
xnor UO_344 (O_344,N_14930,N_14857);
or UO_345 (O_345,N_14902,N_14814);
or UO_346 (O_346,N_14971,N_14875);
nor UO_347 (O_347,N_14976,N_14925);
nor UO_348 (O_348,N_14879,N_14840);
nand UO_349 (O_349,N_14970,N_14897);
and UO_350 (O_350,N_14832,N_14874);
and UO_351 (O_351,N_14882,N_14994);
or UO_352 (O_352,N_14962,N_14975);
xor UO_353 (O_353,N_14975,N_14834);
and UO_354 (O_354,N_14902,N_14972);
and UO_355 (O_355,N_14974,N_14932);
and UO_356 (O_356,N_14865,N_14956);
or UO_357 (O_357,N_14855,N_14898);
xor UO_358 (O_358,N_14863,N_14998);
or UO_359 (O_359,N_14830,N_14820);
and UO_360 (O_360,N_14816,N_14813);
nand UO_361 (O_361,N_14966,N_14854);
nor UO_362 (O_362,N_14825,N_14993);
xor UO_363 (O_363,N_14992,N_14918);
nor UO_364 (O_364,N_14965,N_14941);
nor UO_365 (O_365,N_14840,N_14895);
and UO_366 (O_366,N_14834,N_14845);
and UO_367 (O_367,N_14981,N_14956);
nand UO_368 (O_368,N_14850,N_14851);
and UO_369 (O_369,N_14912,N_14969);
nor UO_370 (O_370,N_14952,N_14961);
xnor UO_371 (O_371,N_14809,N_14822);
and UO_372 (O_372,N_14910,N_14939);
nor UO_373 (O_373,N_14886,N_14835);
or UO_374 (O_374,N_14853,N_14986);
nand UO_375 (O_375,N_14803,N_14924);
xnor UO_376 (O_376,N_14801,N_14970);
nand UO_377 (O_377,N_14987,N_14891);
and UO_378 (O_378,N_14905,N_14914);
and UO_379 (O_379,N_14905,N_14910);
xnor UO_380 (O_380,N_14961,N_14980);
nand UO_381 (O_381,N_14985,N_14819);
xor UO_382 (O_382,N_14860,N_14915);
xnor UO_383 (O_383,N_14889,N_14882);
or UO_384 (O_384,N_14872,N_14986);
nor UO_385 (O_385,N_14815,N_14823);
or UO_386 (O_386,N_14929,N_14963);
or UO_387 (O_387,N_14873,N_14984);
xnor UO_388 (O_388,N_14941,N_14927);
and UO_389 (O_389,N_14912,N_14977);
xor UO_390 (O_390,N_14818,N_14898);
or UO_391 (O_391,N_14848,N_14902);
and UO_392 (O_392,N_14872,N_14848);
nand UO_393 (O_393,N_14899,N_14823);
xnor UO_394 (O_394,N_14805,N_14967);
or UO_395 (O_395,N_14881,N_14947);
and UO_396 (O_396,N_14805,N_14893);
nand UO_397 (O_397,N_14862,N_14919);
xor UO_398 (O_398,N_14873,N_14928);
or UO_399 (O_399,N_14803,N_14814);
and UO_400 (O_400,N_14862,N_14933);
or UO_401 (O_401,N_14970,N_14888);
nand UO_402 (O_402,N_14926,N_14902);
xnor UO_403 (O_403,N_14800,N_14883);
nor UO_404 (O_404,N_14922,N_14978);
xnor UO_405 (O_405,N_14861,N_14924);
or UO_406 (O_406,N_14815,N_14839);
or UO_407 (O_407,N_14881,N_14926);
nor UO_408 (O_408,N_14851,N_14990);
and UO_409 (O_409,N_14906,N_14965);
xnor UO_410 (O_410,N_14929,N_14837);
nor UO_411 (O_411,N_14845,N_14984);
nand UO_412 (O_412,N_14902,N_14843);
xnor UO_413 (O_413,N_14938,N_14897);
nand UO_414 (O_414,N_14836,N_14861);
or UO_415 (O_415,N_14873,N_14940);
or UO_416 (O_416,N_14802,N_14812);
or UO_417 (O_417,N_14991,N_14814);
nor UO_418 (O_418,N_14875,N_14810);
xnor UO_419 (O_419,N_14823,N_14906);
xnor UO_420 (O_420,N_14916,N_14833);
xor UO_421 (O_421,N_14978,N_14895);
or UO_422 (O_422,N_14856,N_14809);
and UO_423 (O_423,N_14959,N_14807);
xor UO_424 (O_424,N_14888,N_14938);
or UO_425 (O_425,N_14874,N_14984);
or UO_426 (O_426,N_14925,N_14812);
nor UO_427 (O_427,N_14917,N_14927);
nor UO_428 (O_428,N_14812,N_14880);
xnor UO_429 (O_429,N_14933,N_14962);
or UO_430 (O_430,N_14849,N_14972);
xor UO_431 (O_431,N_14861,N_14810);
xor UO_432 (O_432,N_14963,N_14851);
or UO_433 (O_433,N_14880,N_14851);
and UO_434 (O_434,N_14896,N_14901);
nor UO_435 (O_435,N_14986,N_14965);
xnor UO_436 (O_436,N_14889,N_14956);
nor UO_437 (O_437,N_14942,N_14841);
xnor UO_438 (O_438,N_14968,N_14991);
and UO_439 (O_439,N_14977,N_14945);
nand UO_440 (O_440,N_14910,N_14908);
nand UO_441 (O_441,N_14853,N_14837);
and UO_442 (O_442,N_14841,N_14838);
or UO_443 (O_443,N_14951,N_14800);
and UO_444 (O_444,N_14965,N_14853);
xor UO_445 (O_445,N_14969,N_14808);
or UO_446 (O_446,N_14949,N_14965);
nor UO_447 (O_447,N_14991,N_14857);
or UO_448 (O_448,N_14808,N_14968);
nor UO_449 (O_449,N_14816,N_14972);
or UO_450 (O_450,N_14866,N_14871);
or UO_451 (O_451,N_14908,N_14876);
nor UO_452 (O_452,N_14964,N_14987);
xnor UO_453 (O_453,N_14896,N_14928);
or UO_454 (O_454,N_14819,N_14972);
nor UO_455 (O_455,N_14822,N_14910);
nand UO_456 (O_456,N_14834,N_14933);
and UO_457 (O_457,N_14835,N_14934);
xnor UO_458 (O_458,N_14938,N_14853);
or UO_459 (O_459,N_14878,N_14948);
nor UO_460 (O_460,N_14831,N_14883);
nor UO_461 (O_461,N_14816,N_14853);
and UO_462 (O_462,N_14910,N_14885);
or UO_463 (O_463,N_14985,N_14916);
and UO_464 (O_464,N_14882,N_14938);
and UO_465 (O_465,N_14953,N_14920);
and UO_466 (O_466,N_14822,N_14803);
and UO_467 (O_467,N_14819,N_14943);
nand UO_468 (O_468,N_14853,N_14818);
and UO_469 (O_469,N_14914,N_14992);
or UO_470 (O_470,N_14938,N_14855);
nand UO_471 (O_471,N_14969,N_14996);
nand UO_472 (O_472,N_14858,N_14920);
or UO_473 (O_473,N_14877,N_14804);
nand UO_474 (O_474,N_14888,N_14889);
nor UO_475 (O_475,N_14896,N_14827);
nor UO_476 (O_476,N_14958,N_14987);
nand UO_477 (O_477,N_14806,N_14820);
xnor UO_478 (O_478,N_14840,N_14915);
nor UO_479 (O_479,N_14885,N_14950);
nand UO_480 (O_480,N_14817,N_14984);
or UO_481 (O_481,N_14966,N_14981);
xnor UO_482 (O_482,N_14907,N_14915);
nand UO_483 (O_483,N_14929,N_14836);
nor UO_484 (O_484,N_14985,N_14979);
nand UO_485 (O_485,N_14905,N_14969);
nand UO_486 (O_486,N_14954,N_14812);
xnor UO_487 (O_487,N_14926,N_14976);
or UO_488 (O_488,N_14950,N_14887);
and UO_489 (O_489,N_14959,N_14898);
or UO_490 (O_490,N_14880,N_14813);
xnor UO_491 (O_491,N_14891,N_14926);
and UO_492 (O_492,N_14894,N_14905);
nor UO_493 (O_493,N_14936,N_14815);
xnor UO_494 (O_494,N_14853,N_14990);
and UO_495 (O_495,N_14863,N_14823);
or UO_496 (O_496,N_14890,N_14951);
or UO_497 (O_497,N_14873,N_14808);
xor UO_498 (O_498,N_14835,N_14990);
or UO_499 (O_499,N_14955,N_14915);
or UO_500 (O_500,N_14824,N_14835);
xnor UO_501 (O_501,N_14906,N_14932);
nand UO_502 (O_502,N_14843,N_14893);
nand UO_503 (O_503,N_14905,N_14987);
xnor UO_504 (O_504,N_14960,N_14915);
nand UO_505 (O_505,N_14980,N_14917);
and UO_506 (O_506,N_14802,N_14923);
xnor UO_507 (O_507,N_14921,N_14805);
xnor UO_508 (O_508,N_14937,N_14932);
or UO_509 (O_509,N_14897,N_14822);
nor UO_510 (O_510,N_14857,N_14969);
xor UO_511 (O_511,N_14831,N_14966);
and UO_512 (O_512,N_14841,N_14879);
and UO_513 (O_513,N_14941,N_14997);
nand UO_514 (O_514,N_14842,N_14883);
xor UO_515 (O_515,N_14958,N_14901);
xnor UO_516 (O_516,N_14882,N_14861);
or UO_517 (O_517,N_14855,N_14958);
or UO_518 (O_518,N_14831,N_14901);
nor UO_519 (O_519,N_14968,N_14896);
xor UO_520 (O_520,N_14910,N_14803);
xnor UO_521 (O_521,N_14984,N_14852);
nand UO_522 (O_522,N_14944,N_14928);
xor UO_523 (O_523,N_14852,N_14949);
xor UO_524 (O_524,N_14895,N_14990);
and UO_525 (O_525,N_14990,N_14898);
nand UO_526 (O_526,N_14971,N_14807);
nor UO_527 (O_527,N_14876,N_14859);
or UO_528 (O_528,N_14980,N_14815);
nand UO_529 (O_529,N_14908,N_14821);
and UO_530 (O_530,N_14826,N_14882);
xnor UO_531 (O_531,N_14806,N_14934);
nand UO_532 (O_532,N_14964,N_14809);
xnor UO_533 (O_533,N_14835,N_14863);
and UO_534 (O_534,N_14878,N_14929);
nand UO_535 (O_535,N_14932,N_14980);
or UO_536 (O_536,N_14952,N_14864);
or UO_537 (O_537,N_14971,N_14846);
nor UO_538 (O_538,N_14811,N_14899);
nor UO_539 (O_539,N_14872,N_14853);
nor UO_540 (O_540,N_14887,N_14960);
and UO_541 (O_541,N_14901,N_14981);
nand UO_542 (O_542,N_14962,N_14854);
nand UO_543 (O_543,N_14834,N_14839);
or UO_544 (O_544,N_14863,N_14950);
nand UO_545 (O_545,N_14951,N_14924);
xnor UO_546 (O_546,N_14801,N_14847);
and UO_547 (O_547,N_14982,N_14947);
xnor UO_548 (O_548,N_14839,N_14855);
nor UO_549 (O_549,N_14987,N_14971);
nor UO_550 (O_550,N_14930,N_14882);
nand UO_551 (O_551,N_14934,N_14987);
or UO_552 (O_552,N_14890,N_14845);
xor UO_553 (O_553,N_14966,N_14807);
nor UO_554 (O_554,N_14856,N_14954);
or UO_555 (O_555,N_14817,N_14909);
xnor UO_556 (O_556,N_14848,N_14949);
nand UO_557 (O_557,N_14965,N_14998);
nand UO_558 (O_558,N_14958,N_14916);
or UO_559 (O_559,N_14920,N_14941);
xor UO_560 (O_560,N_14923,N_14887);
xor UO_561 (O_561,N_14877,N_14969);
nor UO_562 (O_562,N_14810,N_14908);
xnor UO_563 (O_563,N_14991,N_14981);
xnor UO_564 (O_564,N_14972,N_14987);
xnor UO_565 (O_565,N_14958,N_14995);
nand UO_566 (O_566,N_14890,N_14994);
nand UO_567 (O_567,N_14849,N_14802);
nor UO_568 (O_568,N_14903,N_14813);
xnor UO_569 (O_569,N_14829,N_14827);
nor UO_570 (O_570,N_14843,N_14924);
nor UO_571 (O_571,N_14820,N_14863);
nor UO_572 (O_572,N_14966,N_14982);
xor UO_573 (O_573,N_14938,N_14994);
and UO_574 (O_574,N_14911,N_14873);
nand UO_575 (O_575,N_14918,N_14818);
or UO_576 (O_576,N_14949,N_14939);
nor UO_577 (O_577,N_14820,N_14842);
nand UO_578 (O_578,N_14805,N_14868);
and UO_579 (O_579,N_14934,N_14801);
nand UO_580 (O_580,N_14991,N_14872);
or UO_581 (O_581,N_14986,N_14885);
nand UO_582 (O_582,N_14879,N_14898);
or UO_583 (O_583,N_14811,N_14943);
and UO_584 (O_584,N_14882,N_14879);
nor UO_585 (O_585,N_14986,N_14846);
nor UO_586 (O_586,N_14826,N_14838);
or UO_587 (O_587,N_14889,N_14876);
and UO_588 (O_588,N_14809,N_14819);
xnor UO_589 (O_589,N_14863,N_14980);
and UO_590 (O_590,N_14858,N_14939);
xor UO_591 (O_591,N_14982,N_14805);
nand UO_592 (O_592,N_14864,N_14915);
nor UO_593 (O_593,N_14903,N_14876);
and UO_594 (O_594,N_14839,N_14915);
or UO_595 (O_595,N_14900,N_14978);
nor UO_596 (O_596,N_14848,N_14833);
nand UO_597 (O_597,N_14879,N_14987);
nand UO_598 (O_598,N_14877,N_14880);
and UO_599 (O_599,N_14965,N_14901);
nand UO_600 (O_600,N_14969,N_14844);
nand UO_601 (O_601,N_14918,N_14946);
and UO_602 (O_602,N_14999,N_14870);
nand UO_603 (O_603,N_14963,N_14886);
and UO_604 (O_604,N_14807,N_14939);
and UO_605 (O_605,N_14923,N_14903);
nand UO_606 (O_606,N_14828,N_14963);
nand UO_607 (O_607,N_14981,N_14934);
nand UO_608 (O_608,N_14858,N_14875);
or UO_609 (O_609,N_14920,N_14971);
nor UO_610 (O_610,N_14897,N_14811);
nand UO_611 (O_611,N_14875,N_14853);
nand UO_612 (O_612,N_14850,N_14904);
nor UO_613 (O_613,N_14866,N_14851);
and UO_614 (O_614,N_14996,N_14828);
nor UO_615 (O_615,N_14991,N_14811);
xnor UO_616 (O_616,N_14923,N_14904);
nor UO_617 (O_617,N_14830,N_14951);
nand UO_618 (O_618,N_14874,N_14811);
or UO_619 (O_619,N_14934,N_14999);
xor UO_620 (O_620,N_14945,N_14860);
xnor UO_621 (O_621,N_14868,N_14995);
and UO_622 (O_622,N_14844,N_14839);
or UO_623 (O_623,N_14968,N_14962);
xor UO_624 (O_624,N_14976,N_14977);
xnor UO_625 (O_625,N_14830,N_14967);
nor UO_626 (O_626,N_14956,N_14996);
xnor UO_627 (O_627,N_14867,N_14913);
nand UO_628 (O_628,N_14845,N_14930);
nor UO_629 (O_629,N_14999,N_14962);
or UO_630 (O_630,N_14844,N_14824);
nor UO_631 (O_631,N_14987,N_14901);
xnor UO_632 (O_632,N_14915,N_14996);
nor UO_633 (O_633,N_14912,N_14921);
or UO_634 (O_634,N_14814,N_14848);
nor UO_635 (O_635,N_14830,N_14831);
nand UO_636 (O_636,N_14896,N_14942);
and UO_637 (O_637,N_14802,N_14937);
nor UO_638 (O_638,N_14954,N_14944);
nor UO_639 (O_639,N_14801,N_14983);
and UO_640 (O_640,N_14923,N_14885);
nand UO_641 (O_641,N_14977,N_14810);
xnor UO_642 (O_642,N_14829,N_14953);
or UO_643 (O_643,N_14895,N_14926);
nand UO_644 (O_644,N_14800,N_14813);
or UO_645 (O_645,N_14856,N_14998);
and UO_646 (O_646,N_14949,N_14955);
nor UO_647 (O_647,N_14845,N_14830);
nor UO_648 (O_648,N_14987,N_14867);
xnor UO_649 (O_649,N_14806,N_14993);
nor UO_650 (O_650,N_14839,N_14898);
nand UO_651 (O_651,N_14826,N_14972);
nand UO_652 (O_652,N_14874,N_14865);
nor UO_653 (O_653,N_14820,N_14977);
and UO_654 (O_654,N_14890,N_14971);
and UO_655 (O_655,N_14982,N_14884);
xor UO_656 (O_656,N_14811,N_14891);
xor UO_657 (O_657,N_14878,N_14887);
xnor UO_658 (O_658,N_14862,N_14840);
nand UO_659 (O_659,N_14980,N_14832);
nand UO_660 (O_660,N_14801,N_14921);
xnor UO_661 (O_661,N_14828,N_14858);
or UO_662 (O_662,N_14803,N_14900);
xor UO_663 (O_663,N_14979,N_14893);
and UO_664 (O_664,N_14843,N_14950);
xnor UO_665 (O_665,N_14960,N_14845);
nand UO_666 (O_666,N_14833,N_14987);
nand UO_667 (O_667,N_14993,N_14977);
nor UO_668 (O_668,N_14872,N_14928);
xnor UO_669 (O_669,N_14896,N_14937);
nand UO_670 (O_670,N_14910,N_14999);
xnor UO_671 (O_671,N_14908,N_14983);
or UO_672 (O_672,N_14898,N_14922);
nand UO_673 (O_673,N_14828,N_14847);
nand UO_674 (O_674,N_14880,N_14889);
nor UO_675 (O_675,N_14890,N_14924);
and UO_676 (O_676,N_14901,N_14998);
nor UO_677 (O_677,N_14884,N_14904);
nor UO_678 (O_678,N_14823,N_14891);
nor UO_679 (O_679,N_14891,N_14865);
and UO_680 (O_680,N_14875,N_14872);
and UO_681 (O_681,N_14808,N_14944);
nor UO_682 (O_682,N_14832,N_14922);
nand UO_683 (O_683,N_14867,N_14897);
or UO_684 (O_684,N_14952,N_14994);
nand UO_685 (O_685,N_14965,N_14991);
nand UO_686 (O_686,N_14812,N_14846);
nand UO_687 (O_687,N_14964,N_14831);
xor UO_688 (O_688,N_14852,N_14810);
and UO_689 (O_689,N_14987,N_14853);
and UO_690 (O_690,N_14961,N_14948);
or UO_691 (O_691,N_14873,N_14939);
and UO_692 (O_692,N_14853,N_14934);
nor UO_693 (O_693,N_14858,N_14806);
and UO_694 (O_694,N_14982,N_14961);
nor UO_695 (O_695,N_14991,N_14830);
and UO_696 (O_696,N_14810,N_14867);
or UO_697 (O_697,N_14849,N_14807);
or UO_698 (O_698,N_14879,N_14899);
nor UO_699 (O_699,N_14925,N_14890);
nor UO_700 (O_700,N_14957,N_14914);
xnor UO_701 (O_701,N_14916,N_14881);
and UO_702 (O_702,N_14946,N_14916);
nor UO_703 (O_703,N_14927,N_14831);
and UO_704 (O_704,N_14878,N_14816);
and UO_705 (O_705,N_14822,N_14997);
or UO_706 (O_706,N_14836,N_14933);
and UO_707 (O_707,N_14889,N_14895);
nor UO_708 (O_708,N_14998,N_14920);
nor UO_709 (O_709,N_14994,N_14965);
nand UO_710 (O_710,N_14878,N_14916);
xor UO_711 (O_711,N_14890,N_14911);
nor UO_712 (O_712,N_14918,N_14955);
or UO_713 (O_713,N_14858,N_14929);
nor UO_714 (O_714,N_14936,N_14970);
or UO_715 (O_715,N_14821,N_14950);
and UO_716 (O_716,N_14929,N_14911);
and UO_717 (O_717,N_14806,N_14855);
xnor UO_718 (O_718,N_14864,N_14844);
or UO_719 (O_719,N_14933,N_14914);
or UO_720 (O_720,N_14801,N_14829);
xor UO_721 (O_721,N_14983,N_14949);
xnor UO_722 (O_722,N_14825,N_14883);
and UO_723 (O_723,N_14920,N_14823);
nand UO_724 (O_724,N_14928,N_14977);
nand UO_725 (O_725,N_14869,N_14956);
nand UO_726 (O_726,N_14908,N_14934);
nand UO_727 (O_727,N_14918,N_14807);
xnor UO_728 (O_728,N_14859,N_14995);
nor UO_729 (O_729,N_14851,N_14809);
xor UO_730 (O_730,N_14997,N_14864);
nand UO_731 (O_731,N_14800,N_14895);
nor UO_732 (O_732,N_14970,N_14885);
nand UO_733 (O_733,N_14976,N_14857);
nand UO_734 (O_734,N_14891,N_14995);
nor UO_735 (O_735,N_14991,N_14848);
or UO_736 (O_736,N_14957,N_14818);
xnor UO_737 (O_737,N_14976,N_14989);
or UO_738 (O_738,N_14904,N_14887);
xor UO_739 (O_739,N_14920,N_14960);
nor UO_740 (O_740,N_14808,N_14823);
xnor UO_741 (O_741,N_14847,N_14915);
xnor UO_742 (O_742,N_14801,N_14886);
and UO_743 (O_743,N_14962,N_14921);
and UO_744 (O_744,N_14857,N_14944);
nor UO_745 (O_745,N_14840,N_14804);
xor UO_746 (O_746,N_14958,N_14889);
or UO_747 (O_747,N_14914,N_14842);
and UO_748 (O_748,N_14913,N_14892);
and UO_749 (O_749,N_14958,N_14850);
and UO_750 (O_750,N_14870,N_14826);
or UO_751 (O_751,N_14968,N_14895);
and UO_752 (O_752,N_14964,N_14843);
nor UO_753 (O_753,N_14842,N_14904);
xor UO_754 (O_754,N_14969,N_14893);
xnor UO_755 (O_755,N_14818,N_14997);
or UO_756 (O_756,N_14821,N_14850);
xor UO_757 (O_757,N_14837,N_14893);
nand UO_758 (O_758,N_14849,N_14993);
nand UO_759 (O_759,N_14878,N_14921);
xnor UO_760 (O_760,N_14938,N_14914);
and UO_761 (O_761,N_14975,N_14933);
and UO_762 (O_762,N_14834,N_14897);
xnor UO_763 (O_763,N_14926,N_14955);
nand UO_764 (O_764,N_14954,N_14878);
or UO_765 (O_765,N_14818,N_14843);
and UO_766 (O_766,N_14802,N_14906);
xnor UO_767 (O_767,N_14862,N_14903);
nor UO_768 (O_768,N_14936,N_14842);
and UO_769 (O_769,N_14897,N_14801);
nor UO_770 (O_770,N_14804,N_14913);
xnor UO_771 (O_771,N_14957,N_14912);
nand UO_772 (O_772,N_14970,N_14931);
xor UO_773 (O_773,N_14843,N_14943);
or UO_774 (O_774,N_14975,N_14810);
and UO_775 (O_775,N_14992,N_14919);
nand UO_776 (O_776,N_14809,N_14854);
and UO_777 (O_777,N_14884,N_14890);
nor UO_778 (O_778,N_14940,N_14932);
or UO_779 (O_779,N_14876,N_14874);
xor UO_780 (O_780,N_14801,N_14926);
xnor UO_781 (O_781,N_14810,N_14995);
xnor UO_782 (O_782,N_14935,N_14998);
xnor UO_783 (O_783,N_14934,N_14848);
nor UO_784 (O_784,N_14980,N_14843);
nand UO_785 (O_785,N_14873,N_14935);
xnor UO_786 (O_786,N_14812,N_14961);
xnor UO_787 (O_787,N_14944,N_14826);
nor UO_788 (O_788,N_14834,N_14976);
xor UO_789 (O_789,N_14965,N_14981);
xnor UO_790 (O_790,N_14919,N_14804);
nand UO_791 (O_791,N_14836,N_14849);
or UO_792 (O_792,N_14819,N_14823);
xor UO_793 (O_793,N_14836,N_14999);
nand UO_794 (O_794,N_14838,N_14960);
and UO_795 (O_795,N_14920,N_14850);
nor UO_796 (O_796,N_14970,N_14945);
nand UO_797 (O_797,N_14982,N_14951);
and UO_798 (O_798,N_14924,N_14948);
nand UO_799 (O_799,N_14975,N_14873);
xor UO_800 (O_800,N_14951,N_14968);
or UO_801 (O_801,N_14927,N_14916);
nand UO_802 (O_802,N_14863,N_14860);
xnor UO_803 (O_803,N_14877,N_14967);
nor UO_804 (O_804,N_14947,N_14856);
nor UO_805 (O_805,N_14899,N_14862);
or UO_806 (O_806,N_14923,N_14944);
nor UO_807 (O_807,N_14949,N_14891);
nand UO_808 (O_808,N_14852,N_14994);
nor UO_809 (O_809,N_14837,N_14950);
xnor UO_810 (O_810,N_14823,N_14803);
xor UO_811 (O_811,N_14854,N_14992);
nand UO_812 (O_812,N_14993,N_14814);
and UO_813 (O_813,N_14984,N_14921);
nor UO_814 (O_814,N_14942,N_14801);
and UO_815 (O_815,N_14841,N_14984);
nor UO_816 (O_816,N_14903,N_14824);
and UO_817 (O_817,N_14994,N_14924);
nand UO_818 (O_818,N_14969,N_14882);
nand UO_819 (O_819,N_14884,N_14899);
nor UO_820 (O_820,N_14901,N_14806);
or UO_821 (O_821,N_14986,N_14888);
nor UO_822 (O_822,N_14914,N_14805);
nor UO_823 (O_823,N_14970,N_14990);
or UO_824 (O_824,N_14860,N_14819);
or UO_825 (O_825,N_14968,N_14986);
and UO_826 (O_826,N_14894,N_14914);
or UO_827 (O_827,N_14846,N_14815);
nor UO_828 (O_828,N_14833,N_14983);
nor UO_829 (O_829,N_14821,N_14884);
xnor UO_830 (O_830,N_14866,N_14957);
or UO_831 (O_831,N_14847,N_14817);
and UO_832 (O_832,N_14856,N_14847);
nor UO_833 (O_833,N_14987,N_14810);
nand UO_834 (O_834,N_14908,N_14951);
nor UO_835 (O_835,N_14982,N_14911);
or UO_836 (O_836,N_14854,N_14870);
nor UO_837 (O_837,N_14879,N_14930);
xor UO_838 (O_838,N_14956,N_14894);
nand UO_839 (O_839,N_14811,N_14849);
nor UO_840 (O_840,N_14957,N_14868);
nor UO_841 (O_841,N_14898,N_14935);
nor UO_842 (O_842,N_14812,N_14931);
and UO_843 (O_843,N_14978,N_14944);
xnor UO_844 (O_844,N_14832,N_14804);
xor UO_845 (O_845,N_14834,N_14863);
nor UO_846 (O_846,N_14816,N_14996);
nor UO_847 (O_847,N_14997,N_14847);
nor UO_848 (O_848,N_14854,N_14875);
nor UO_849 (O_849,N_14969,N_14876);
xnor UO_850 (O_850,N_14914,N_14954);
xor UO_851 (O_851,N_14830,N_14842);
and UO_852 (O_852,N_14963,N_14943);
or UO_853 (O_853,N_14925,N_14948);
xnor UO_854 (O_854,N_14956,N_14837);
or UO_855 (O_855,N_14862,N_14858);
xor UO_856 (O_856,N_14859,N_14838);
xnor UO_857 (O_857,N_14977,N_14971);
nand UO_858 (O_858,N_14926,N_14871);
and UO_859 (O_859,N_14992,N_14859);
or UO_860 (O_860,N_14803,N_14968);
or UO_861 (O_861,N_14847,N_14924);
nand UO_862 (O_862,N_14913,N_14908);
nor UO_863 (O_863,N_14960,N_14867);
nand UO_864 (O_864,N_14966,N_14990);
nand UO_865 (O_865,N_14888,N_14944);
xnor UO_866 (O_866,N_14855,N_14876);
xnor UO_867 (O_867,N_14923,N_14913);
nand UO_868 (O_868,N_14979,N_14871);
xor UO_869 (O_869,N_14997,N_14815);
nand UO_870 (O_870,N_14941,N_14946);
nor UO_871 (O_871,N_14991,N_14945);
xnor UO_872 (O_872,N_14936,N_14840);
or UO_873 (O_873,N_14955,N_14866);
nor UO_874 (O_874,N_14934,N_14914);
and UO_875 (O_875,N_14969,N_14858);
and UO_876 (O_876,N_14994,N_14968);
xor UO_877 (O_877,N_14852,N_14952);
nor UO_878 (O_878,N_14986,N_14961);
xor UO_879 (O_879,N_14865,N_14849);
nand UO_880 (O_880,N_14827,N_14949);
xnor UO_881 (O_881,N_14869,N_14959);
nand UO_882 (O_882,N_14847,N_14907);
and UO_883 (O_883,N_14922,N_14970);
and UO_884 (O_884,N_14952,N_14854);
nand UO_885 (O_885,N_14800,N_14879);
xor UO_886 (O_886,N_14915,N_14843);
or UO_887 (O_887,N_14833,N_14865);
and UO_888 (O_888,N_14977,N_14979);
xor UO_889 (O_889,N_14903,N_14881);
and UO_890 (O_890,N_14801,N_14979);
nor UO_891 (O_891,N_14803,N_14805);
xnor UO_892 (O_892,N_14915,N_14822);
xnor UO_893 (O_893,N_14890,N_14806);
nor UO_894 (O_894,N_14990,N_14861);
or UO_895 (O_895,N_14952,N_14937);
and UO_896 (O_896,N_14928,N_14959);
nor UO_897 (O_897,N_14827,N_14824);
nor UO_898 (O_898,N_14809,N_14940);
nor UO_899 (O_899,N_14960,N_14981);
xnor UO_900 (O_900,N_14826,N_14920);
or UO_901 (O_901,N_14841,N_14917);
and UO_902 (O_902,N_14974,N_14947);
nand UO_903 (O_903,N_14830,N_14953);
and UO_904 (O_904,N_14922,N_14950);
nand UO_905 (O_905,N_14972,N_14868);
xor UO_906 (O_906,N_14822,N_14914);
nand UO_907 (O_907,N_14961,N_14914);
xnor UO_908 (O_908,N_14831,N_14983);
or UO_909 (O_909,N_14975,N_14896);
and UO_910 (O_910,N_14850,N_14849);
nor UO_911 (O_911,N_14859,N_14839);
nand UO_912 (O_912,N_14939,N_14915);
and UO_913 (O_913,N_14864,N_14884);
and UO_914 (O_914,N_14854,N_14948);
and UO_915 (O_915,N_14847,N_14851);
and UO_916 (O_916,N_14933,N_14973);
nand UO_917 (O_917,N_14951,N_14839);
nand UO_918 (O_918,N_14969,N_14956);
and UO_919 (O_919,N_14807,N_14816);
nand UO_920 (O_920,N_14867,N_14974);
nor UO_921 (O_921,N_14968,N_14911);
or UO_922 (O_922,N_14847,N_14819);
and UO_923 (O_923,N_14862,N_14843);
and UO_924 (O_924,N_14842,N_14986);
xor UO_925 (O_925,N_14851,N_14917);
and UO_926 (O_926,N_14809,N_14987);
or UO_927 (O_927,N_14821,N_14817);
or UO_928 (O_928,N_14880,N_14916);
nor UO_929 (O_929,N_14821,N_14940);
and UO_930 (O_930,N_14850,N_14819);
xnor UO_931 (O_931,N_14831,N_14955);
nand UO_932 (O_932,N_14933,N_14832);
nor UO_933 (O_933,N_14929,N_14943);
nand UO_934 (O_934,N_14844,N_14986);
nor UO_935 (O_935,N_14810,N_14830);
nor UO_936 (O_936,N_14900,N_14850);
nand UO_937 (O_937,N_14950,N_14848);
xnor UO_938 (O_938,N_14941,N_14883);
and UO_939 (O_939,N_14937,N_14821);
and UO_940 (O_940,N_14843,N_14812);
or UO_941 (O_941,N_14961,N_14951);
nor UO_942 (O_942,N_14941,N_14893);
xor UO_943 (O_943,N_14864,N_14840);
nor UO_944 (O_944,N_14988,N_14976);
nor UO_945 (O_945,N_14864,N_14849);
nand UO_946 (O_946,N_14804,N_14810);
or UO_947 (O_947,N_14841,N_14887);
and UO_948 (O_948,N_14951,N_14948);
and UO_949 (O_949,N_14923,N_14950);
or UO_950 (O_950,N_14855,N_14841);
nor UO_951 (O_951,N_14936,N_14895);
nand UO_952 (O_952,N_14814,N_14862);
nor UO_953 (O_953,N_14884,N_14805);
or UO_954 (O_954,N_14815,N_14876);
nor UO_955 (O_955,N_14934,N_14913);
and UO_956 (O_956,N_14971,N_14836);
or UO_957 (O_957,N_14804,N_14860);
xor UO_958 (O_958,N_14944,N_14853);
nor UO_959 (O_959,N_14903,N_14820);
nor UO_960 (O_960,N_14877,N_14896);
and UO_961 (O_961,N_14912,N_14897);
nor UO_962 (O_962,N_14834,N_14956);
nor UO_963 (O_963,N_14809,N_14806);
nand UO_964 (O_964,N_14906,N_14966);
nor UO_965 (O_965,N_14810,N_14970);
xnor UO_966 (O_966,N_14902,N_14941);
and UO_967 (O_967,N_14808,N_14928);
and UO_968 (O_968,N_14838,N_14845);
nor UO_969 (O_969,N_14995,N_14961);
or UO_970 (O_970,N_14962,N_14956);
and UO_971 (O_971,N_14881,N_14889);
nor UO_972 (O_972,N_14972,N_14978);
or UO_973 (O_973,N_14805,N_14975);
xnor UO_974 (O_974,N_14986,N_14880);
or UO_975 (O_975,N_14842,N_14809);
or UO_976 (O_976,N_14976,N_14948);
or UO_977 (O_977,N_14912,N_14859);
or UO_978 (O_978,N_14988,N_14839);
nor UO_979 (O_979,N_14970,N_14915);
nand UO_980 (O_980,N_14935,N_14915);
and UO_981 (O_981,N_14830,N_14970);
xnor UO_982 (O_982,N_14839,N_14926);
or UO_983 (O_983,N_14850,N_14909);
nor UO_984 (O_984,N_14946,N_14857);
xnor UO_985 (O_985,N_14897,N_14993);
nand UO_986 (O_986,N_14973,N_14949);
nand UO_987 (O_987,N_14895,N_14942);
nand UO_988 (O_988,N_14811,N_14869);
xor UO_989 (O_989,N_14864,N_14929);
xor UO_990 (O_990,N_14903,N_14938);
xnor UO_991 (O_991,N_14917,N_14957);
xor UO_992 (O_992,N_14918,N_14849);
or UO_993 (O_993,N_14984,N_14833);
nor UO_994 (O_994,N_14803,N_14876);
nor UO_995 (O_995,N_14998,N_14916);
xnor UO_996 (O_996,N_14887,N_14969);
xor UO_997 (O_997,N_14835,N_14823);
nand UO_998 (O_998,N_14925,N_14874);
nor UO_999 (O_999,N_14997,N_14877);
or UO_1000 (O_1000,N_14959,N_14974);
xnor UO_1001 (O_1001,N_14963,N_14881);
nand UO_1002 (O_1002,N_14890,N_14966);
or UO_1003 (O_1003,N_14910,N_14859);
or UO_1004 (O_1004,N_14885,N_14890);
nor UO_1005 (O_1005,N_14966,N_14934);
nand UO_1006 (O_1006,N_14852,N_14847);
or UO_1007 (O_1007,N_14883,N_14928);
or UO_1008 (O_1008,N_14887,N_14824);
or UO_1009 (O_1009,N_14816,N_14987);
and UO_1010 (O_1010,N_14903,N_14889);
nand UO_1011 (O_1011,N_14990,N_14886);
nor UO_1012 (O_1012,N_14960,N_14907);
xnor UO_1013 (O_1013,N_14975,N_14931);
or UO_1014 (O_1014,N_14805,N_14901);
nand UO_1015 (O_1015,N_14909,N_14936);
or UO_1016 (O_1016,N_14987,N_14969);
nor UO_1017 (O_1017,N_14867,N_14914);
xor UO_1018 (O_1018,N_14965,N_14850);
nand UO_1019 (O_1019,N_14934,N_14828);
nor UO_1020 (O_1020,N_14979,N_14972);
nor UO_1021 (O_1021,N_14946,N_14884);
nand UO_1022 (O_1022,N_14979,N_14828);
nor UO_1023 (O_1023,N_14865,N_14823);
nand UO_1024 (O_1024,N_14884,N_14966);
nor UO_1025 (O_1025,N_14909,N_14803);
xor UO_1026 (O_1026,N_14940,N_14947);
or UO_1027 (O_1027,N_14853,N_14923);
xor UO_1028 (O_1028,N_14824,N_14864);
or UO_1029 (O_1029,N_14946,N_14891);
nor UO_1030 (O_1030,N_14921,N_14955);
nand UO_1031 (O_1031,N_14833,N_14845);
or UO_1032 (O_1032,N_14936,N_14859);
nor UO_1033 (O_1033,N_14934,N_14939);
xnor UO_1034 (O_1034,N_14846,N_14959);
nor UO_1035 (O_1035,N_14935,N_14991);
xor UO_1036 (O_1036,N_14928,N_14800);
nand UO_1037 (O_1037,N_14953,N_14861);
nor UO_1038 (O_1038,N_14971,N_14869);
or UO_1039 (O_1039,N_14994,N_14984);
nand UO_1040 (O_1040,N_14941,N_14981);
and UO_1041 (O_1041,N_14816,N_14883);
nor UO_1042 (O_1042,N_14954,N_14870);
or UO_1043 (O_1043,N_14981,N_14883);
nor UO_1044 (O_1044,N_14839,N_14944);
xnor UO_1045 (O_1045,N_14831,N_14832);
and UO_1046 (O_1046,N_14887,N_14889);
nor UO_1047 (O_1047,N_14886,N_14877);
nand UO_1048 (O_1048,N_14809,N_14992);
and UO_1049 (O_1049,N_14942,N_14836);
and UO_1050 (O_1050,N_14941,N_14938);
or UO_1051 (O_1051,N_14956,N_14877);
nand UO_1052 (O_1052,N_14861,N_14809);
xor UO_1053 (O_1053,N_14972,N_14908);
or UO_1054 (O_1054,N_14925,N_14840);
and UO_1055 (O_1055,N_14916,N_14855);
and UO_1056 (O_1056,N_14827,N_14954);
nand UO_1057 (O_1057,N_14990,N_14806);
or UO_1058 (O_1058,N_14986,N_14818);
nor UO_1059 (O_1059,N_14892,N_14953);
or UO_1060 (O_1060,N_14800,N_14899);
xor UO_1061 (O_1061,N_14833,N_14997);
nor UO_1062 (O_1062,N_14901,N_14962);
nor UO_1063 (O_1063,N_14909,N_14808);
xnor UO_1064 (O_1064,N_14807,N_14968);
xnor UO_1065 (O_1065,N_14887,N_14909);
and UO_1066 (O_1066,N_14852,N_14805);
nor UO_1067 (O_1067,N_14879,N_14834);
or UO_1068 (O_1068,N_14972,N_14881);
nor UO_1069 (O_1069,N_14969,N_14899);
and UO_1070 (O_1070,N_14953,N_14964);
nor UO_1071 (O_1071,N_14960,N_14993);
nand UO_1072 (O_1072,N_14914,N_14953);
nor UO_1073 (O_1073,N_14984,N_14827);
and UO_1074 (O_1074,N_14942,N_14929);
nand UO_1075 (O_1075,N_14825,N_14841);
and UO_1076 (O_1076,N_14937,N_14922);
or UO_1077 (O_1077,N_14808,N_14913);
or UO_1078 (O_1078,N_14994,N_14998);
or UO_1079 (O_1079,N_14908,N_14978);
or UO_1080 (O_1080,N_14822,N_14843);
or UO_1081 (O_1081,N_14931,N_14800);
nand UO_1082 (O_1082,N_14883,N_14863);
or UO_1083 (O_1083,N_14937,N_14984);
or UO_1084 (O_1084,N_14851,N_14834);
nand UO_1085 (O_1085,N_14894,N_14845);
and UO_1086 (O_1086,N_14868,N_14909);
xnor UO_1087 (O_1087,N_14939,N_14968);
xnor UO_1088 (O_1088,N_14953,N_14893);
or UO_1089 (O_1089,N_14974,N_14895);
and UO_1090 (O_1090,N_14937,N_14851);
xnor UO_1091 (O_1091,N_14830,N_14862);
and UO_1092 (O_1092,N_14946,N_14953);
or UO_1093 (O_1093,N_14837,N_14991);
nand UO_1094 (O_1094,N_14804,N_14870);
or UO_1095 (O_1095,N_14860,N_14864);
nor UO_1096 (O_1096,N_14943,N_14842);
and UO_1097 (O_1097,N_14807,N_14850);
nor UO_1098 (O_1098,N_14930,N_14941);
nor UO_1099 (O_1099,N_14902,N_14862);
and UO_1100 (O_1100,N_14947,N_14813);
and UO_1101 (O_1101,N_14868,N_14996);
nor UO_1102 (O_1102,N_14830,N_14867);
nand UO_1103 (O_1103,N_14849,N_14986);
nor UO_1104 (O_1104,N_14866,N_14999);
xor UO_1105 (O_1105,N_14927,N_14900);
nand UO_1106 (O_1106,N_14972,N_14964);
or UO_1107 (O_1107,N_14809,N_14880);
or UO_1108 (O_1108,N_14935,N_14807);
nand UO_1109 (O_1109,N_14901,N_14975);
xnor UO_1110 (O_1110,N_14861,N_14846);
nor UO_1111 (O_1111,N_14976,N_14960);
nor UO_1112 (O_1112,N_14976,N_14908);
and UO_1113 (O_1113,N_14851,N_14979);
and UO_1114 (O_1114,N_14926,N_14815);
xnor UO_1115 (O_1115,N_14859,N_14980);
and UO_1116 (O_1116,N_14965,N_14912);
and UO_1117 (O_1117,N_14853,N_14828);
nand UO_1118 (O_1118,N_14847,N_14938);
and UO_1119 (O_1119,N_14826,N_14843);
nor UO_1120 (O_1120,N_14996,N_14992);
nand UO_1121 (O_1121,N_14900,N_14888);
nand UO_1122 (O_1122,N_14803,N_14819);
nand UO_1123 (O_1123,N_14946,N_14804);
nand UO_1124 (O_1124,N_14958,N_14832);
and UO_1125 (O_1125,N_14839,N_14838);
and UO_1126 (O_1126,N_14842,N_14920);
xor UO_1127 (O_1127,N_14917,N_14939);
and UO_1128 (O_1128,N_14969,N_14973);
nor UO_1129 (O_1129,N_14992,N_14838);
nor UO_1130 (O_1130,N_14831,N_14957);
nor UO_1131 (O_1131,N_14912,N_14951);
and UO_1132 (O_1132,N_14959,N_14809);
nand UO_1133 (O_1133,N_14907,N_14992);
nand UO_1134 (O_1134,N_14820,N_14948);
and UO_1135 (O_1135,N_14835,N_14884);
and UO_1136 (O_1136,N_14956,N_14895);
nand UO_1137 (O_1137,N_14846,N_14864);
xor UO_1138 (O_1138,N_14802,N_14919);
xnor UO_1139 (O_1139,N_14961,N_14803);
and UO_1140 (O_1140,N_14913,N_14822);
and UO_1141 (O_1141,N_14885,N_14844);
or UO_1142 (O_1142,N_14912,N_14928);
or UO_1143 (O_1143,N_14832,N_14976);
and UO_1144 (O_1144,N_14844,N_14979);
and UO_1145 (O_1145,N_14834,N_14872);
and UO_1146 (O_1146,N_14827,N_14933);
nand UO_1147 (O_1147,N_14955,N_14986);
nor UO_1148 (O_1148,N_14877,N_14840);
or UO_1149 (O_1149,N_14919,N_14989);
xor UO_1150 (O_1150,N_14875,N_14908);
and UO_1151 (O_1151,N_14918,N_14996);
nor UO_1152 (O_1152,N_14825,N_14875);
nand UO_1153 (O_1153,N_14892,N_14911);
or UO_1154 (O_1154,N_14983,N_14860);
or UO_1155 (O_1155,N_14825,N_14896);
nor UO_1156 (O_1156,N_14828,N_14891);
and UO_1157 (O_1157,N_14894,N_14852);
xor UO_1158 (O_1158,N_14916,N_14965);
nor UO_1159 (O_1159,N_14882,N_14838);
or UO_1160 (O_1160,N_14908,N_14970);
or UO_1161 (O_1161,N_14948,N_14893);
xor UO_1162 (O_1162,N_14937,N_14948);
nand UO_1163 (O_1163,N_14999,N_14863);
or UO_1164 (O_1164,N_14990,N_14998);
nor UO_1165 (O_1165,N_14985,N_14880);
and UO_1166 (O_1166,N_14854,N_14926);
xor UO_1167 (O_1167,N_14905,N_14830);
nor UO_1168 (O_1168,N_14802,N_14960);
xnor UO_1169 (O_1169,N_14954,N_14963);
nand UO_1170 (O_1170,N_14812,N_14967);
nand UO_1171 (O_1171,N_14994,N_14899);
xnor UO_1172 (O_1172,N_14972,N_14898);
nand UO_1173 (O_1173,N_14898,N_14967);
nand UO_1174 (O_1174,N_14878,N_14848);
or UO_1175 (O_1175,N_14943,N_14957);
nand UO_1176 (O_1176,N_14982,N_14844);
nand UO_1177 (O_1177,N_14808,N_14834);
xnor UO_1178 (O_1178,N_14843,N_14867);
xnor UO_1179 (O_1179,N_14966,N_14804);
and UO_1180 (O_1180,N_14881,N_14978);
nor UO_1181 (O_1181,N_14896,N_14831);
nand UO_1182 (O_1182,N_14849,N_14980);
xor UO_1183 (O_1183,N_14983,N_14872);
xor UO_1184 (O_1184,N_14973,N_14892);
nand UO_1185 (O_1185,N_14827,N_14913);
xnor UO_1186 (O_1186,N_14906,N_14950);
xnor UO_1187 (O_1187,N_14940,N_14816);
nand UO_1188 (O_1188,N_14852,N_14953);
nand UO_1189 (O_1189,N_14995,N_14980);
and UO_1190 (O_1190,N_14881,N_14887);
xnor UO_1191 (O_1191,N_14925,N_14801);
and UO_1192 (O_1192,N_14934,N_14957);
nor UO_1193 (O_1193,N_14936,N_14875);
nand UO_1194 (O_1194,N_14931,N_14821);
nand UO_1195 (O_1195,N_14839,N_14843);
or UO_1196 (O_1196,N_14971,N_14870);
nor UO_1197 (O_1197,N_14992,N_14932);
xor UO_1198 (O_1198,N_14978,N_14837);
nor UO_1199 (O_1199,N_14857,N_14943);
nand UO_1200 (O_1200,N_14859,N_14944);
or UO_1201 (O_1201,N_14806,N_14945);
nand UO_1202 (O_1202,N_14926,N_14948);
nor UO_1203 (O_1203,N_14859,N_14933);
or UO_1204 (O_1204,N_14980,N_14973);
xor UO_1205 (O_1205,N_14887,N_14865);
and UO_1206 (O_1206,N_14845,N_14934);
nor UO_1207 (O_1207,N_14925,N_14852);
xnor UO_1208 (O_1208,N_14894,N_14983);
xnor UO_1209 (O_1209,N_14827,N_14941);
xor UO_1210 (O_1210,N_14876,N_14991);
and UO_1211 (O_1211,N_14978,N_14952);
or UO_1212 (O_1212,N_14900,N_14989);
or UO_1213 (O_1213,N_14922,N_14838);
nand UO_1214 (O_1214,N_14870,N_14990);
nand UO_1215 (O_1215,N_14881,N_14830);
and UO_1216 (O_1216,N_14924,N_14983);
xor UO_1217 (O_1217,N_14897,N_14981);
xor UO_1218 (O_1218,N_14846,N_14911);
nor UO_1219 (O_1219,N_14989,N_14899);
xnor UO_1220 (O_1220,N_14921,N_14895);
and UO_1221 (O_1221,N_14924,N_14953);
or UO_1222 (O_1222,N_14883,N_14823);
xnor UO_1223 (O_1223,N_14934,N_14971);
and UO_1224 (O_1224,N_14895,N_14845);
nor UO_1225 (O_1225,N_14952,N_14988);
or UO_1226 (O_1226,N_14870,N_14969);
nand UO_1227 (O_1227,N_14899,N_14816);
or UO_1228 (O_1228,N_14985,N_14983);
or UO_1229 (O_1229,N_14935,N_14801);
or UO_1230 (O_1230,N_14861,N_14994);
nand UO_1231 (O_1231,N_14913,N_14912);
nand UO_1232 (O_1232,N_14999,N_14937);
or UO_1233 (O_1233,N_14833,N_14831);
nand UO_1234 (O_1234,N_14874,N_14957);
and UO_1235 (O_1235,N_14856,N_14958);
or UO_1236 (O_1236,N_14950,N_14984);
xnor UO_1237 (O_1237,N_14880,N_14849);
or UO_1238 (O_1238,N_14814,N_14995);
and UO_1239 (O_1239,N_14960,N_14900);
nor UO_1240 (O_1240,N_14999,N_14977);
nand UO_1241 (O_1241,N_14895,N_14951);
nor UO_1242 (O_1242,N_14898,N_14894);
xnor UO_1243 (O_1243,N_14957,N_14902);
and UO_1244 (O_1244,N_14843,N_14906);
and UO_1245 (O_1245,N_14813,N_14815);
or UO_1246 (O_1246,N_14885,N_14866);
and UO_1247 (O_1247,N_14822,N_14850);
or UO_1248 (O_1248,N_14863,N_14929);
or UO_1249 (O_1249,N_14956,N_14929);
or UO_1250 (O_1250,N_14815,N_14886);
or UO_1251 (O_1251,N_14938,N_14973);
nand UO_1252 (O_1252,N_14912,N_14890);
xnor UO_1253 (O_1253,N_14942,N_14858);
xnor UO_1254 (O_1254,N_14971,N_14964);
nor UO_1255 (O_1255,N_14886,N_14897);
nand UO_1256 (O_1256,N_14896,N_14969);
and UO_1257 (O_1257,N_14805,N_14883);
or UO_1258 (O_1258,N_14824,N_14831);
xor UO_1259 (O_1259,N_14981,N_14840);
nor UO_1260 (O_1260,N_14870,N_14911);
or UO_1261 (O_1261,N_14800,N_14848);
nor UO_1262 (O_1262,N_14895,N_14965);
xor UO_1263 (O_1263,N_14955,N_14846);
or UO_1264 (O_1264,N_14852,N_14876);
or UO_1265 (O_1265,N_14899,N_14964);
or UO_1266 (O_1266,N_14816,N_14989);
and UO_1267 (O_1267,N_14937,N_14966);
nor UO_1268 (O_1268,N_14870,N_14936);
and UO_1269 (O_1269,N_14869,N_14875);
and UO_1270 (O_1270,N_14835,N_14922);
or UO_1271 (O_1271,N_14894,N_14882);
nor UO_1272 (O_1272,N_14900,N_14828);
and UO_1273 (O_1273,N_14997,N_14983);
nand UO_1274 (O_1274,N_14904,N_14952);
nor UO_1275 (O_1275,N_14843,N_14870);
xnor UO_1276 (O_1276,N_14910,N_14845);
or UO_1277 (O_1277,N_14913,N_14919);
xor UO_1278 (O_1278,N_14817,N_14873);
and UO_1279 (O_1279,N_14913,N_14824);
or UO_1280 (O_1280,N_14874,N_14857);
nor UO_1281 (O_1281,N_14913,N_14970);
or UO_1282 (O_1282,N_14890,N_14997);
and UO_1283 (O_1283,N_14928,N_14950);
xor UO_1284 (O_1284,N_14906,N_14962);
or UO_1285 (O_1285,N_14836,N_14956);
or UO_1286 (O_1286,N_14968,N_14805);
nor UO_1287 (O_1287,N_14814,N_14900);
or UO_1288 (O_1288,N_14832,N_14817);
xnor UO_1289 (O_1289,N_14990,N_14993);
or UO_1290 (O_1290,N_14973,N_14905);
and UO_1291 (O_1291,N_14936,N_14805);
and UO_1292 (O_1292,N_14805,N_14951);
xnor UO_1293 (O_1293,N_14904,N_14801);
or UO_1294 (O_1294,N_14972,N_14875);
nand UO_1295 (O_1295,N_14890,N_14905);
xnor UO_1296 (O_1296,N_14821,N_14945);
xor UO_1297 (O_1297,N_14868,N_14827);
nand UO_1298 (O_1298,N_14858,N_14879);
nor UO_1299 (O_1299,N_14890,N_14996);
nor UO_1300 (O_1300,N_14808,N_14825);
nand UO_1301 (O_1301,N_14958,N_14830);
nor UO_1302 (O_1302,N_14852,N_14921);
xnor UO_1303 (O_1303,N_14868,N_14839);
and UO_1304 (O_1304,N_14969,N_14924);
xnor UO_1305 (O_1305,N_14955,N_14984);
nand UO_1306 (O_1306,N_14950,N_14976);
nor UO_1307 (O_1307,N_14834,N_14949);
nor UO_1308 (O_1308,N_14850,N_14944);
nand UO_1309 (O_1309,N_14854,N_14997);
nor UO_1310 (O_1310,N_14940,N_14976);
or UO_1311 (O_1311,N_14872,N_14847);
nand UO_1312 (O_1312,N_14920,N_14990);
nor UO_1313 (O_1313,N_14956,N_14857);
nor UO_1314 (O_1314,N_14921,N_14964);
xnor UO_1315 (O_1315,N_14929,N_14967);
nor UO_1316 (O_1316,N_14926,N_14863);
nor UO_1317 (O_1317,N_14988,N_14880);
nor UO_1318 (O_1318,N_14878,N_14936);
xnor UO_1319 (O_1319,N_14910,N_14834);
and UO_1320 (O_1320,N_14902,N_14914);
and UO_1321 (O_1321,N_14964,N_14934);
or UO_1322 (O_1322,N_14885,N_14963);
nor UO_1323 (O_1323,N_14845,N_14919);
or UO_1324 (O_1324,N_14884,N_14810);
nand UO_1325 (O_1325,N_14805,N_14937);
xor UO_1326 (O_1326,N_14804,N_14956);
and UO_1327 (O_1327,N_14872,N_14822);
and UO_1328 (O_1328,N_14803,N_14890);
and UO_1329 (O_1329,N_14958,N_14913);
and UO_1330 (O_1330,N_14898,N_14890);
nand UO_1331 (O_1331,N_14896,N_14826);
and UO_1332 (O_1332,N_14852,N_14958);
nand UO_1333 (O_1333,N_14948,N_14868);
and UO_1334 (O_1334,N_14945,N_14872);
xnor UO_1335 (O_1335,N_14943,N_14918);
and UO_1336 (O_1336,N_14865,N_14894);
xor UO_1337 (O_1337,N_14908,N_14826);
and UO_1338 (O_1338,N_14855,N_14925);
xnor UO_1339 (O_1339,N_14981,N_14954);
and UO_1340 (O_1340,N_14892,N_14807);
and UO_1341 (O_1341,N_14889,N_14914);
xnor UO_1342 (O_1342,N_14807,N_14948);
and UO_1343 (O_1343,N_14926,N_14924);
nand UO_1344 (O_1344,N_14975,N_14961);
xnor UO_1345 (O_1345,N_14829,N_14846);
and UO_1346 (O_1346,N_14891,N_14892);
xnor UO_1347 (O_1347,N_14817,N_14822);
or UO_1348 (O_1348,N_14929,N_14902);
or UO_1349 (O_1349,N_14866,N_14982);
nand UO_1350 (O_1350,N_14860,N_14977);
xnor UO_1351 (O_1351,N_14959,N_14859);
xor UO_1352 (O_1352,N_14886,N_14843);
nand UO_1353 (O_1353,N_14905,N_14883);
nand UO_1354 (O_1354,N_14901,N_14863);
xnor UO_1355 (O_1355,N_14993,N_14823);
nor UO_1356 (O_1356,N_14869,N_14922);
or UO_1357 (O_1357,N_14932,N_14854);
xor UO_1358 (O_1358,N_14913,N_14988);
xor UO_1359 (O_1359,N_14890,N_14840);
or UO_1360 (O_1360,N_14822,N_14857);
or UO_1361 (O_1361,N_14801,N_14955);
xor UO_1362 (O_1362,N_14873,N_14988);
and UO_1363 (O_1363,N_14979,N_14956);
xnor UO_1364 (O_1364,N_14925,N_14913);
nand UO_1365 (O_1365,N_14861,N_14825);
or UO_1366 (O_1366,N_14851,N_14999);
or UO_1367 (O_1367,N_14917,N_14894);
and UO_1368 (O_1368,N_14952,N_14968);
nor UO_1369 (O_1369,N_14937,N_14941);
and UO_1370 (O_1370,N_14888,N_14852);
nor UO_1371 (O_1371,N_14929,N_14880);
nand UO_1372 (O_1372,N_14897,N_14998);
or UO_1373 (O_1373,N_14933,N_14894);
and UO_1374 (O_1374,N_14885,N_14911);
nand UO_1375 (O_1375,N_14880,N_14917);
or UO_1376 (O_1376,N_14888,N_14958);
nor UO_1377 (O_1377,N_14866,N_14962);
or UO_1378 (O_1378,N_14970,N_14808);
nor UO_1379 (O_1379,N_14916,N_14892);
xnor UO_1380 (O_1380,N_14952,N_14995);
nor UO_1381 (O_1381,N_14900,N_14845);
xor UO_1382 (O_1382,N_14954,N_14903);
or UO_1383 (O_1383,N_14996,N_14988);
and UO_1384 (O_1384,N_14921,N_14869);
or UO_1385 (O_1385,N_14831,N_14944);
and UO_1386 (O_1386,N_14919,N_14929);
or UO_1387 (O_1387,N_14871,N_14962);
nand UO_1388 (O_1388,N_14845,N_14871);
nand UO_1389 (O_1389,N_14996,N_14833);
nand UO_1390 (O_1390,N_14953,N_14833);
xor UO_1391 (O_1391,N_14986,N_14816);
or UO_1392 (O_1392,N_14870,N_14885);
nand UO_1393 (O_1393,N_14995,N_14816);
or UO_1394 (O_1394,N_14979,N_14835);
and UO_1395 (O_1395,N_14870,N_14996);
and UO_1396 (O_1396,N_14879,N_14957);
nor UO_1397 (O_1397,N_14896,N_14982);
xnor UO_1398 (O_1398,N_14949,N_14905);
nand UO_1399 (O_1399,N_14814,N_14858);
nor UO_1400 (O_1400,N_14895,N_14870);
nand UO_1401 (O_1401,N_14809,N_14921);
or UO_1402 (O_1402,N_14868,N_14896);
xnor UO_1403 (O_1403,N_14831,N_14806);
or UO_1404 (O_1404,N_14836,N_14865);
and UO_1405 (O_1405,N_14967,N_14846);
nor UO_1406 (O_1406,N_14897,N_14873);
nor UO_1407 (O_1407,N_14805,N_14909);
nand UO_1408 (O_1408,N_14885,N_14957);
nand UO_1409 (O_1409,N_14823,N_14978);
and UO_1410 (O_1410,N_14874,N_14926);
nand UO_1411 (O_1411,N_14910,N_14998);
nand UO_1412 (O_1412,N_14830,N_14994);
nor UO_1413 (O_1413,N_14801,N_14929);
xor UO_1414 (O_1414,N_14831,N_14980);
xnor UO_1415 (O_1415,N_14970,N_14892);
and UO_1416 (O_1416,N_14969,N_14981);
and UO_1417 (O_1417,N_14994,N_14874);
xnor UO_1418 (O_1418,N_14820,N_14996);
or UO_1419 (O_1419,N_14975,N_14868);
and UO_1420 (O_1420,N_14814,N_14932);
and UO_1421 (O_1421,N_14999,N_14833);
and UO_1422 (O_1422,N_14836,N_14966);
nand UO_1423 (O_1423,N_14973,N_14839);
or UO_1424 (O_1424,N_14800,N_14995);
nor UO_1425 (O_1425,N_14895,N_14817);
or UO_1426 (O_1426,N_14904,N_14848);
nand UO_1427 (O_1427,N_14843,N_14934);
nand UO_1428 (O_1428,N_14962,N_14830);
xnor UO_1429 (O_1429,N_14900,N_14984);
and UO_1430 (O_1430,N_14814,N_14935);
nand UO_1431 (O_1431,N_14956,N_14994);
xnor UO_1432 (O_1432,N_14952,N_14801);
or UO_1433 (O_1433,N_14917,N_14951);
nand UO_1434 (O_1434,N_14999,N_14840);
xor UO_1435 (O_1435,N_14915,N_14889);
nand UO_1436 (O_1436,N_14905,N_14993);
xor UO_1437 (O_1437,N_14813,N_14834);
nor UO_1438 (O_1438,N_14862,N_14927);
nor UO_1439 (O_1439,N_14934,N_14884);
xor UO_1440 (O_1440,N_14823,N_14869);
xor UO_1441 (O_1441,N_14892,N_14968);
and UO_1442 (O_1442,N_14805,N_14973);
or UO_1443 (O_1443,N_14933,N_14930);
xnor UO_1444 (O_1444,N_14870,N_14818);
xnor UO_1445 (O_1445,N_14840,N_14849);
or UO_1446 (O_1446,N_14903,N_14961);
xor UO_1447 (O_1447,N_14961,N_14857);
xnor UO_1448 (O_1448,N_14849,N_14928);
nand UO_1449 (O_1449,N_14832,N_14807);
xnor UO_1450 (O_1450,N_14959,N_14901);
nor UO_1451 (O_1451,N_14984,N_14946);
or UO_1452 (O_1452,N_14884,N_14958);
or UO_1453 (O_1453,N_14807,N_14998);
nor UO_1454 (O_1454,N_14920,N_14913);
or UO_1455 (O_1455,N_14823,N_14988);
nor UO_1456 (O_1456,N_14835,N_14876);
nand UO_1457 (O_1457,N_14991,N_14964);
nand UO_1458 (O_1458,N_14927,N_14867);
xor UO_1459 (O_1459,N_14940,N_14911);
xor UO_1460 (O_1460,N_14982,N_14883);
nand UO_1461 (O_1461,N_14889,N_14906);
and UO_1462 (O_1462,N_14817,N_14833);
or UO_1463 (O_1463,N_14818,N_14950);
or UO_1464 (O_1464,N_14800,N_14982);
and UO_1465 (O_1465,N_14969,N_14971);
or UO_1466 (O_1466,N_14992,N_14885);
xnor UO_1467 (O_1467,N_14955,N_14995);
nand UO_1468 (O_1468,N_14854,N_14858);
nor UO_1469 (O_1469,N_14916,N_14823);
nand UO_1470 (O_1470,N_14933,N_14815);
xnor UO_1471 (O_1471,N_14877,N_14818);
xnor UO_1472 (O_1472,N_14994,N_14964);
nand UO_1473 (O_1473,N_14982,N_14802);
nand UO_1474 (O_1474,N_14824,N_14863);
nor UO_1475 (O_1475,N_14802,N_14962);
or UO_1476 (O_1476,N_14980,N_14959);
xor UO_1477 (O_1477,N_14805,N_14810);
nand UO_1478 (O_1478,N_14811,N_14867);
nor UO_1479 (O_1479,N_14838,N_14987);
xnor UO_1480 (O_1480,N_14818,N_14917);
or UO_1481 (O_1481,N_14846,N_14957);
nand UO_1482 (O_1482,N_14924,N_14946);
nand UO_1483 (O_1483,N_14961,N_14863);
nand UO_1484 (O_1484,N_14996,N_14824);
or UO_1485 (O_1485,N_14948,N_14975);
or UO_1486 (O_1486,N_14841,N_14965);
xor UO_1487 (O_1487,N_14913,N_14893);
xnor UO_1488 (O_1488,N_14978,N_14811);
nor UO_1489 (O_1489,N_14864,N_14802);
and UO_1490 (O_1490,N_14992,N_14972);
and UO_1491 (O_1491,N_14932,N_14948);
and UO_1492 (O_1492,N_14862,N_14881);
and UO_1493 (O_1493,N_14896,N_14844);
and UO_1494 (O_1494,N_14805,N_14899);
nor UO_1495 (O_1495,N_14938,N_14931);
or UO_1496 (O_1496,N_14863,N_14877);
or UO_1497 (O_1497,N_14953,N_14927);
and UO_1498 (O_1498,N_14925,N_14841);
xnor UO_1499 (O_1499,N_14971,N_14938);
and UO_1500 (O_1500,N_14908,N_14859);
nor UO_1501 (O_1501,N_14938,N_14879);
or UO_1502 (O_1502,N_14825,N_14959);
or UO_1503 (O_1503,N_14816,N_14847);
and UO_1504 (O_1504,N_14802,N_14878);
nand UO_1505 (O_1505,N_14833,N_14851);
nor UO_1506 (O_1506,N_14907,N_14850);
and UO_1507 (O_1507,N_14980,N_14882);
nand UO_1508 (O_1508,N_14999,N_14869);
xnor UO_1509 (O_1509,N_14801,N_14914);
and UO_1510 (O_1510,N_14983,N_14828);
nor UO_1511 (O_1511,N_14862,N_14953);
and UO_1512 (O_1512,N_14926,N_14917);
xor UO_1513 (O_1513,N_14957,N_14892);
or UO_1514 (O_1514,N_14987,N_14943);
or UO_1515 (O_1515,N_14802,N_14940);
and UO_1516 (O_1516,N_14842,N_14838);
and UO_1517 (O_1517,N_14861,N_14819);
and UO_1518 (O_1518,N_14901,N_14935);
xnor UO_1519 (O_1519,N_14885,N_14966);
xnor UO_1520 (O_1520,N_14925,N_14816);
and UO_1521 (O_1521,N_14886,N_14865);
and UO_1522 (O_1522,N_14882,N_14911);
nor UO_1523 (O_1523,N_14954,N_14925);
nand UO_1524 (O_1524,N_14932,N_14869);
nor UO_1525 (O_1525,N_14858,N_14982);
nor UO_1526 (O_1526,N_14903,N_14894);
or UO_1527 (O_1527,N_14967,N_14989);
xor UO_1528 (O_1528,N_14803,N_14998);
nand UO_1529 (O_1529,N_14992,N_14928);
nor UO_1530 (O_1530,N_14942,N_14872);
nand UO_1531 (O_1531,N_14973,N_14808);
and UO_1532 (O_1532,N_14870,N_14888);
nor UO_1533 (O_1533,N_14914,N_14839);
or UO_1534 (O_1534,N_14938,N_14870);
nand UO_1535 (O_1535,N_14880,N_14907);
xor UO_1536 (O_1536,N_14912,N_14881);
and UO_1537 (O_1537,N_14920,N_14817);
xor UO_1538 (O_1538,N_14997,N_14977);
or UO_1539 (O_1539,N_14993,N_14866);
or UO_1540 (O_1540,N_14930,N_14850);
nor UO_1541 (O_1541,N_14807,N_14984);
or UO_1542 (O_1542,N_14919,N_14950);
nor UO_1543 (O_1543,N_14875,N_14963);
and UO_1544 (O_1544,N_14946,N_14834);
nand UO_1545 (O_1545,N_14907,N_14938);
nand UO_1546 (O_1546,N_14996,N_14928);
xnor UO_1547 (O_1547,N_14866,N_14938);
or UO_1548 (O_1548,N_14938,N_14923);
nand UO_1549 (O_1549,N_14900,N_14836);
nand UO_1550 (O_1550,N_14882,N_14944);
and UO_1551 (O_1551,N_14928,N_14937);
or UO_1552 (O_1552,N_14942,N_14833);
or UO_1553 (O_1553,N_14890,N_14967);
xor UO_1554 (O_1554,N_14980,N_14885);
nand UO_1555 (O_1555,N_14835,N_14935);
and UO_1556 (O_1556,N_14825,N_14815);
and UO_1557 (O_1557,N_14883,N_14945);
xnor UO_1558 (O_1558,N_14973,N_14844);
or UO_1559 (O_1559,N_14816,N_14931);
and UO_1560 (O_1560,N_14911,N_14902);
or UO_1561 (O_1561,N_14805,N_14841);
nor UO_1562 (O_1562,N_14816,N_14846);
xnor UO_1563 (O_1563,N_14885,N_14803);
xnor UO_1564 (O_1564,N_14822,N_14964);
or UO_1565 (O_1565,N_14877,N_14940);
or UO_1566 (O_1566,N_14980,N_14964);
xnor UO_1567 (O_1567,N_14901,N_14913);
or UO_1568 (O_1568,N_14891,N_14901);
nand UO_1569 (O_1569,N_14911,N_14901);
and UO_1570 (O_1570,N_14849,N_14985);
or UO_1571 (O_1571,N_14930,N_14985);
nor UO_1572 (O_1572,N_14846,N_14916);
nand UO_1573 (O_1573,N_14970,N_14807);
or UO_1574 (O_1574,N_14958,N_14885);
and UO_1575 (O_1575,N_14913,N_14801);
or UO_1576 (O_1576,N_14959,N_14908);
nand UO_1577 (O_1577,N_14851,N_14898);
and UO_1578 (O_1578,N_14893,N_14908);
nand UO_1579 (O_1579,N_14861,N_14919);
xor UO_1580 (O_1580,N_14869,N_14982);
or UO_1581 (O_1581,N_14935,N_14961);
and UO_1582 (O_1582,N_14878,N_14922);
or UO_1583 (O_1583,N_14827,N_14971);
or UO_1584 (O_1584,N_14992,N_14955);
nand UO_1585 (O_1585,N_14976,N_14997);
nor UO_1586 (O_1586,N_14841,N_14913);
xor UO_1587 (O_1587,N_14841,N_14808);
nor UO_1588 (O_1588,N_14852,N_14819);
nand UO_1589 (O_1589,N_14954,N_14879);
xnor UO_1590 (O_1590,N_14811,N_14822);
or UO_1591 (O_1591,N_14902,N_14907);
or UO_1592 (O_1592,N_14887,N_14970);
nor UO_1593 (O_1593,N_14860,N_14850);
or UO_1594 (O_1594,N_14917,N_14953);
nor UO_1595 (O_1595,N_14846,N_14802);
and UO_1596 (O_1596,N_14904,N_14812);
and UO_1597 (O_1597,N_14917,N_14950);
nor UO_1598 (O_1598,N_14931,N_14911);
xor UO_1599 (O_1599,N_14834,N_14998);
and UO_1600 (O_1600,N_14859,N_14977);
or UO_1601 (O_1601,N_14968,N_14975);
xnor UO_1602 (O_1602,N_14927,N_14887);
nor UO_1603 (O_1603,N_14832,N_14939);
nand UO_1604 (O_1604,N_14977,N_14805);
nor UO_1605 (O_1605,N_14824,N_14868);
nand UO_1606 (O_1606,N_14869,N_14816);
xnor UO_1607 (O_1607,N_14901,N_14977);
or UO_1608 (O_1608,N_14807,N_14858);
and UO_1609 (O_1609,N_14904,N_14983);
nand UO_1610 (O_1610,N_14991,N_14898);
nor UO_1611 (O_1611,N_14985,N_14806);
nor UO_1612 (O_1612,N_14910,N_14917);
or UO_1613 (O_1613,N_14838,N_14951);
xor UO_1614 (O_1614,N_14957,N_14898);
xor UO_1615 (O_1615,N_14922,N_14979);
nor UO_1616 (O_1616,N_14968,N_14893);
or UO_1617 (O_1617,N_14897,N_14942);
and UO_1618 (O_1618,N_14871,N_14991);
xnor UO_1619 (O_1619,N_14958,N_14985);
xnor UO_1620 (O_1620,N_14852,N_14863);
or UO_1621 (O_1621,N_14866,N_14830);
nand UO_1622 (O_1622,N_14865,N_14970);
or UO_1623 (O_1623,N_14913,N_14851);
or UO_1624 (O_1624,N_14819,N_14912);
xor UO_1625 (O_1625,N_14803,N_14880);
nand UO_1626 (O_1626,N_14985,N_14945);
and UO_1627 (O_1627,N_14969,N_14921);
nand UO_1628 (O_1628,N_14969,N_14978);
and UO_1629 (O_1629,N_14801,N_14821);
and UO_1630 (O_1630,N_14906,N_14817);
nand UO_1631 (O_1631,N_14901,N_14917);
or UO_1632 (O_1632,N_14973,N_14962);
nor UO_1633 (O_1633,N_14945,N_14931);
nand UO_1634 (O_1634,N_14868,N_14934);
nand UO_1635 (O_1635,N_14862,N_14891);
nand UO_1636 (O_1636,N_14979,N_14827);
or UO_1637 (O_1637,N_14840,N_14928);
and UO_1638 (O_1638,N_14931,N_14936);
nand UO_1639 (O_1639,N_14924,N_14903);
or UO_1640 (O_1640,N_14981,N_14875);
and UO_1641 (O_1641,N_14841,N_14822);
or UO_1642 (O_1642,N_14926,N_14860);
nand UO_1643 (O_1643,N_14819,N_14874);
or UO_1644 (O_1644,N_14806,N_14826);
and UO_1645 (O_1645,N_14886,N_14999);
xor UO_1646 (O_1646,N_14887,N_14884);
nor UO_1647 (O_1647,N_14821,N_14807);
xnor UO_1648 (O_1648,N_14836,N_14905);
and UO_1649 (O_1649,N_14932,N_14858);
and UO_1650 (O_1650,N_14869,N_14911);
and UO_1651 (O_1651,N_14826,N_14913);
nor UO_1652 (O_1652,N_14830,N_14839);
and UO_1653 (O_1653,N_14875,N_14864);
xor UO_1654 (O_1654,N_14883,N_14996);
nor UO_1655 (O_1655,N_14985,N_14851);
nor UO_1656 (O_1656,N_14894,N_14906);
xor UO_1657 (O_1657,N_14810,N_14844);
xor UO_1658 (O_1658,N_14860,N_14966);
and UO_1659 (O_1659,N_14812,N_14944);
nand UO_1660 (O_1660,N_14939,N_14960);
nor UO_1661 (O_1661,N_14883,N_14828);
nand UO_1662 (O_1662,N_14847,N_14936);
nand UO_1663 (O_1663,N_14810,N_14979);
and UO_1664 (O_1664,N_14926,N_14819);
xnor UO_1665 (O_1665,N_14918,N_14981);
and UO_1666 (O_1666,N_14895,N_14810);
xnor UO_1667 (O_1667,N_14829,N_14951);
or UO_1668 (O_1668,N_14860,N_14942);
nor UO_1669 (O_1669,N_14939,N_14977);
and UO_1670 (O_1670,N_14849,N_14890);
or UO_1671 (O_1671,N_14921,N_14904);
and UO_1672 (O_1672,N_14988,N_14835);
or UO_1673 (O_1673,N_14825,N_14802);
xnor UO_1674 (O_1674,N_14909,N_14835);
and UO_1675 (O_1675,N_14963,N_14833);
nand UO_1676 (O_1676,N_14839,N_14961);
and UO_1677 (O_1677,N_14883,N_14892);
nor UO_1678 (O_1678,N_14807,N_14860);
and UO_1679 (O_1679,N_14856,N_14866);
or UO_1680 (O_1680,N_14976,N_14964);
or UO_1681 (O_1681,N_14825,N_14981);
or UO_1682 (O_1682,N_14826,N_14924);
xor UO_1683 (O_1683,N_14968,N_14934);
nor UO_1684 (O_1684,N_14887,N_14880);
and UO_1685 (O_1685,N_14946,N_14957);
nor UO_1686 (O_1686,N_14936,N_14906);
and UO_1687 (O_1687,N_14830,N_14854);
nand UO_1688 (O_1688,N_14993,N_14821);
or UO_1689 (O_1689,N_14931,N_14860);
xor UO_1690 (O_1690,N_14978,N_14812);
and UO_1691 (O_1691,N_14928,N_14864);
and UO_1692 (O_1692,N_14864,N_14880);
xnor UO_1693 (O_1693,N_14941,N_14967);
or UO_1694 (O_1694,N_14917,N_14816);
or UO_1695 (O_1695,N_14959,N_14925);
nor UO_1696 (O_1696,N_14928,N_14886);
xor UO_1697 (O_1697,N_14844,N_14847);
and UO_1698 (O_1698,N_14879,N_14941);
and UO_1699 (O_1699,N_14822,N_14844);
or UO_1700 (O_1700,N_14853,N_14949);
nand UO_1701 (O_1701,N_14980,N_14855);
or UO_1702 (O_1702,N_14988,N_14938);
and UO_1703 (O_1703,N_14885,N_14920);
nand UO_1704 (O_1704,N_14931,N_14978);
or UO_1705 (O_1705,N_14802,N_14933);
or UO_1706 (O_1706,N_14876,N_14984);
nor UO_1707 (O_1707,N_14876,N_14940);
nand UO_1708 (O_1708,N_14971,N_14867);
nor UO_1709 (O_1709,N_14863,N_14939);
and UO_1710 (O_1710,N_14834,N_14848);
nand UO_1711 (O_1711,N_14930,N_14961);
and UO_1712 (O_1712,N_14948,N_14967);
xor UO_1713 (O_1713,N_14870,N_14841);
nor UO_1714 (O_1714,N_14980,N_14984);
xor UO_1715 (O_1715,N_14973,N_14982);
and UO_1716 (O_1716,N_14840,N_14841);
nor UO_1717 (O_1717,N_14967,N_14872);
nor UO_1718 (O_1718,N_14865,N_14985);
nand UO_1719 (O_1719,N_14981,N_14888);
xnor UO_1720 (O_1720,N_14817,N_14825);
and UO_1721 (O_1721,N_14910,N_14897);
and UO_1722 (O_1722,N_14832,N_14823);
nand UO_1723 (O_1723,N_14905,N_14904);
nor UO_1724 (O_1724,N_14903,N_14915);
nand UO_1725 (O_1725,N_14944,N_14929);
nor UO_1726 (O_1726,N_14838,N_14989);
or UO_1727 (O_1727,N_14913,N_14955);
nor UO_1728 (O_1728,N_14905,N_14868);
or UO_1729 (O_1729,N_14929,N_14991);
xnor UO_1730 (O_1730,N_14912,N_14988);
xor UO_1731 (O_1731,N_14805,N_14897);
xnor UO_1732 (O_1732,N_14883,N_14933);
and UO_1733 (O_1733,N_14829,N_14883);
nand UO_1734 (O_1734,N_14991,N_14971);
nor UO_1735 (O_1735,N_14830,N_14822);
xnor UO_1736 (O_1736,N_14862,N_14813);
nand UO_1737 (O_1737,N_14886,N_14917);
nor UO_1738 (O_1738,N_14849,N_14978);
nand UO_1739 (O_1739,N_14865,N_14892);
and UO_1740 (O_1740,N_14986,N_14835);
and UO_1741 (O_1741,N_14976,N_14889);
nor UO_1742 (O_1742,N_14867,N_14828);
xor UO_1743 (O_1743,N_14986,N_14859);
nor UO_1744 (O_1744,N_14855,N_14934);
and UO_1745 (O_1745,N_14827,N_14849);
xor UO_1746 (O_1746,N_14995,N_14883);
nor UO_1747 (O_1747,N_14847,N_14955);
nor UO_1748 (O_1748,N_14903,N_14804);
xnor UO_1749 (O_1749,N_14955,N_14827);
and UO_1750 (O_1750,N_14997,N_14817);
or UO_1751 (O_1751,N_14840,N_14880);
nand UO_1752 (O_1752,N_14986,N_14870);
or UO_1753 (O_1753,N_14994,N_14849);
and UO_1754 (O_1754,N_14834,N_14900);
nor UO_1755 (O_1755,N_14884,N_14990);
and UO_1756 (O_1756,N_14989,N_14934);
nand UO_1757 (O_1757,N_14873,N_14995);
or UO_1758 (O_1758,N_14916,N_14839);
xnor UO_1759 (O_1759,N_14838,N_14924);
xnor UO_1760 (O_1760,N_14985,N_14873);
and UO_1761 (O_1761,N_14958,N_14926);
nand UO_1762 (O_1762,N_14832,N_14932);
nor UO_1763 (O_1763,N_14809,N_14811);
or UO_1764 (O_1764,N_14906,N_14828);
xor UO_1765 (O_1765,N_14808,N_14915);
and UO_1766 (O_1766,N_14953,N_14841);
or UO_1767 (O_1767,N_14925,N_14965);
xor UO_1768 (O_1768,N_14952,N_14998);
nand UO_1769 (O_1769,N_14846,N_14822);
or UO_1770 (O_1770,N_14803,N_14873);
nor UO_1771 (O_1771,N_14802,N_14983);
xnor UO_1772 (O_1772,N_14950,N_14909);
nand UO_1773 (O_1773,N_14887,N_14952);
nand UO_1774 (O_1774,N_14840,N_14867);
nor UO_1775 (O_1775,N_14843,N_14834);
nor UO_1776 (O_1776,N_14805,N_14985);
nor UO_1777 (O_1777,N_14897,N_14915);
nand UO_1778 (O_1778,N_14900,N_14974);
nand UO_1779 (O_1779,N_14824,N_14838);
nor UO_1780 (O_1780,N_14954,N_14880);
xor UO_1781 (O_1781,N_14932,N_14964);
nand UO_1782 (O_1782,N_14867,N_14819);
or UO_1783 (O_1783,N_14853,N_14841);
nand UO_1784 (O_1784,N_14964,N_14877);
nand UO_1785 (O_1785,N_14853,N_14843);
xor UO_1786 (O_1786,N_14952,N_14885);
nor UO_1787 (O_1787,N_14897,N_14828);
xor UO_1788 (O_1788,N_14890,N_14913);
or UO_1789 (O_1789,N_14966,N_14882);
nor UO_1790 (O_1790,N_14844,N_14811);
nor UO_1791 (O_1791,N_14839,N_14929);
or UO_1792 (O_1792,N_14823,N_14904);
and UO_1793 (O_1793,N_14998,N_14880);
nand UO_1794 (O_1794,N_14825,N_14831);
nand UO_1795 (O_1795,N_14918,N_14877);
nand UO_1796 (O_1796,N_14876,N_14866);
and UO_1797 (O_1797,N_14918,N_14953);
xor UO_1798 (O_1798,N_14825,N_14923);
or UO_1799 (O_1799,N_14915,N_14829);
xnor UO_1800 (O_1800,N_14828,N_14820);
nor UO_1801 (O_1801,N_14881,N_14905);
xor UO_1802 (O_1802,N_14957,N_14958);
and UO_1803 (O_1803,N_14951,N_14928);
or UO_1804 (O_1804,N_14865,N_14972);
or UO_1805 (O_1805,N_14980,N_14931);
nor UO_1806 (O_1806,N_14850,N_14910);
or UO_1807 (O_1807,N_14921,N_14820);
xnor UO_1808 (O_1808,N_14999,N_14822);
xnor UO_1809 (O_1809,N_14973,N_14840);
nand UO_1810 (O_1810,N_14918,N_14914);
nand UO_1811 (O_1811,N_14807,N_14803);
or UO_1812 (O_1812,N_14949,N_14990);
nand UO_1813 (O_1813,N_14979,N_14915);
nor UO_1814 (O_1814,N_14813,N_14876);
and UO_1815 (O_1815,N_14932,N_14803);
nand UO_1816 (O_1816,N_14868,N_14990);
nor UO_1817 (O_1817,N_14830,N_14915);
nor UO_1818 (O_1818,N_14954,N_14923);
or UO_1819 (O_1819,N_14863,N_14913);
nor UO_1820 (O_1820,N_14871,N_14803);
xnor UO_1821 (O_1821,N_14966,N_14931);
or UO_1822 (O_1822,N_14949,N_14862);
xor UO_1823 (O_1823,N_14948,N_14819);
nor UO_1824 (O_1824,N_14903,N_14995);
nor UO_1825 (O_1825,N_14878,N_14877);
or UO_1826 (O_1826,N_14895,N_14904);
and UO_1827 (O_1827,N_14825,N_14854);
nand UO_1828 (O_1828,N_14851,N_14914);
nand UO_1829 (O_1829,N_14826,N_14914);
xor UO_1830 (O_1830,N_14950,N_14927);
nor UO_1831 (O_1831,N_14976,N_14975);
nand UO_1832 (O_1832,N_14927,N_14948);
xnor UO_1833 (O_1833,N_14893,N_14885);
and UO_1834 (O_1834,N_14948,N_14958);
xor UO_1835 (O_1835,N_14873,N_14820);
nand UO_1836 (O_1836,N_14971,N_14868);
nand UO_1837 (O_1837,N_14829,N_14811);
xor UO_1838 (O_1838,N_14872,N_14831);
nand UO_1839 (O_1839,N_14968,N_14914);
and UO_1840 (O_1840,N_14844,N_14831);
or UO_1841 (O_1841,N_14873,N_14851);
xnor UO_1842 (O_1842,N_14944,N_14834);
xnor UO_1843 (O_1843,N_14980,N_14899);
nand UO_1844 (O_1844,N_14894,N_14823);
nor UO_1845 (O_1845,N_14920,N_14853);
xnor UO_1846 (O_1846,N_14928,N_14978);
and UO_1847 (O_1847,N_14880,N_14821);
and UO_1848 (O_1848,N_14978,N_14887);
and UO_1849 (O_1849,N_14945,N_14839);
or UO_1850 (O_1850,N_14973,N_14820);
and UO_1851 (O_1851,N_14942,N_14884);
nor UO_1852 (O_1852,N_14919,N_14938);
and UO_1853 (O_1853,N_14889,N_14941);
or UO_1854 (O_1854,N_14855,N_14902);
nor UO_1855 (O_1855,N_14878,N_14935);
or UO_1856 (O_1856,N_14962,N_14819);
and UO_1857 (O_1857,N_14916,N_14913);
or UO_1858 (O_1858,N_14944,N_14919);
nand UO_1859 (O_1859,N_14947,N_14932);
nand UO_1860 (O_1860,N_14870,N_14842);
nand UO_1861 (O_1861,N_14812,N_14893);
xor UO_1862 (O_1862,N_14829,N_14803);
nand UO_1863 (O_1863,N_14834,N_14966);
xor UO_1864 (O_1864,N_14993,N_14948);
nor UO_1865 (O_1865,N_14896,N_14870);
or UO_1866 (O_1866,N_14854,N_14823);
nor UO_1867 (O_1867,N_14815,N_14870);
and UO_1868 (O_1868,N_14944,N_14925);
nor UO_1869 (O_1869,N_14907,N_14980);
nor UO_1870 (O_1870,N_14948,N_14880);
xor UO_1871 (O_1871,N_14936,N_14883);
nor UO_1872 (O_1872,N_14937,N_14995);
xnor UO_1873 (O_1873,N_14950,N_14820);
or UO_1874 (O_1874,N_14937,N_14987);
xor UO_1875 (O_1875,N_14966,N_14954);
and UO_1876 (O_1876,N_14920,N_14942);
and UO_1877 (O_1877,N_14904,N_14981);
nor UO_1878 (O_1878,N_14884,N_14807);
nand UO_1879 (O_1879,N_14944,N_14996);
nand UO_1880 (O_1880,N_14997,N_14933);
nor UO_1881 (O_1881,N_14961,N_14976);
and UO_1882 (O_1882,N_14874,N_14983);
xnor UO_1883 (O_1883,N_14915,N_14987);
nand UO_1884 (O_1884,N_14883,N_14866);
or UO_1885 (O_1885,N_14803,N_14867);
nor UO_1886 (O_1886,N_14865,N_14863);
or UO_1887 (O_1887,N_14943,N_14802);
or UO_1888 (O_1888,N_14873,N_14929);
nand UO_1889 (O_1889,N_14831,N_14837);
nand UO_1890 (O_1890,N_14875,N_14910);
nand UO_1891 (O_1891,N_14905,N_14884);
nand UO_1892 (O_1892,N_14879,N_14819);
or UO_1893 (O_1893,N_14870,N_14893);
or UO_1894 (O_1894,N_14990,N_14881);
or UO_1895 (O_1895,N_14945,N_14941);
or UO_1896 (O_1896,N_14836,N_14889);
nor UO_1897 (O_1897,N_14988,N_14877);
xor UO_1898 (O_1898,N_14964,N_14958);
and UO_1899 (O_1899,N_14849,N_14979);
or UO_1900 (O_1900,N_14883,N_14864);
nor UO_1901 (O_1901,N_14982,N_14946);
xnor UO_1902 (O_1902,N_14943,N_14949);
and UO_1903 (O_1903,N_14832,N_14903);
or UO_1904 (O_1904,N_14972,N_14903);
nor UO_1905 (O_1905,N_14800,N_14888);
or UO_1906 (O_1906,N_14899,N_14953);
nand UO_1907 (O_1907,N_14831,N_14851);
xor UO_1908 (O_1908,N_14838,N_14934);
or UO_1909 (O_1909,N_14961,N_14974);
nand UO_1910 (O_1910,N_14867,N_14994);
nor UO_1911 (O_1911,N_14806,N_14848);
xor UO_1912 (O_1912,N_14903,N_14859);
or UO_1913 (O_1913,N_14927,N_14998);
nor UO_1914 (O_1914,N_14869,N_14822);
nand UO_1915 (O_1915,N_14870,N_14814);
or UO_1916 (O_1916,N_14825,N_14906);
and UO_1917 (O_1917,N_14918,N_14906);
or UO_1918 (O_1918,N_14879,N_14910);
or UO_1919 (O_1919,N_14850,N_14915);
and UO_1920 (O_1920,N_14888,N_14861);
nand UO_1921 (O_1921,N_14939,N_14850);
nor UO_1922 (O_1922,N_14986,N_14824);
nand UO_1923 (O_1923,N_14930,N_14979);
nor UO_1924 (O_1924,N_14985,N_14933);
nand UO_1925 (O_1925,N_14997,N_14830);
and UO_1926 (O_1926,N_14954,N_14851);
nor UO_1927 (O_1927,N_14809,N_14957);
and UO_1928 (O_1928,N_14803,N_14934);
and UO_1929 (O_1929,N_14992,N_14956);
xor UO_1930 (O_1930,N_14929,N_14865);
and UO_1931 (O_1931,N_14980,N_14921);
and UO_1932 (O_1932,N_14928,N_14930);
nand UO_1933 (O_1933,N_14922,N_14890);
nor UO_1934 (O_1934,N_14950,N_14974);
or UO_1935 (O_1935,N_14819,N_14944);
or UO_1936 (O_1936,N_14994,N_14872);
xnor UO_1937 (O_1937,N_14954,N_14876);
nor UO_1938 (O_1938,N_14881,N_14996);
nor UO_1939 (O_1939,N_14901,N_14934);
nor UO_1940 (O_1940,N_14988,N_14904);
or UO_1941 (O_1941,N_14961,N_14911);
and UO_1942 (O_1942,N_14806,N_14861);
nand UO_1943 (O_1943,N_14945,N_14831);
or UO_1944 (O_1944,N_14910,N_14890);
and UO_1945 (O_1945,N_14957,N_14847);
nor UO_1946 (O_1946,N_14877,N_14965);
xor UO_1947 (O_1947,N_14827,N_14935);
nor UO_1948 (O_1948,N_14866,N_14994);
xor UO_1949 (O_1949,N_14865,N_14939);
or UO_1950 (O_1950,N_14928,N_14816);
xnor UO_1951 (O_1951,N_14884,N_14832);
xor UO_1952 (O_1952,N_14924,N_14892);
and UO_1953 (O_1953,N_14989,N_14940);
or UO_1954 (O_1954,N_14926,N_14823);
xor UO_1955 (O_1955,N_14801,N_14992);
and UO_1956 (O_1956,N_14831,N_14835);
or UO_1957 (O_1957,N_14862,N_14808);
xor UO_1958 (O_1958,N_14953,N_14905);
and UO_1959 (O_1959,N_14807,N_14855);
nor UO_1960 (O_1960,N_14819,N_14987);
and UO_1961 (O_1961,N_14824,N_14893);
or UO_1962 (O_1962,N_14942,N_14901);
or UO_1963 (O_1963,N_14961,N_14925);
nor UO_1964 (O_1964,N_14940,N_14920);
xnor UO_1965 (O_1965,N_14984,N_14924);
nor UO_1966 (O_1966,N_14911,N_14925);
xor UO_1967 (O_1967,N_14996,N_14891);
nand UO_1968 (O_1968,N_14882,N_14885);
and UO_1969 (O_1969,N_14819,N_14824);
nand UO_1970 (O_1970,N_14812,N_14971);
xor UO_1971 (O_1971,N_14931,N_14987);
or UO_1972 (O_1972,N_14861,N_14813);
nand UO_1973 (O_1973,N_14966,N_14863);
xor UO_1974 (O_1974,N_14990,N_14837);
xor UO_1975 (O_1975,N_14886,N_14913);
nand UO_1976 (O_1976,N_14876,N_14871);
xor UO_1977 (O_1977,N_14815,N_14822);
xor UO_1978 (O_1978,N_14882,N_14920);
xor UO_1979 (O_1979,N_14818,N_14992);
and UO_1980 (O_1980,N_14846,N_14825);
or UO_1981 (O_1981,N_14834,N_14955);
xor UO_1982 (O_1982,N_14907,N_14924);
nor UO_1983 (O_1983,N_14934,N_14859);
nand UO_1984 (O_1984,N_14902,N_14990);
xnor UO_1985 (O_1985,N_14867,N_14801);
nor UO_1986 (O_1986,N_14912,N_14898);
nor UO_1987 (O_1987,N_14886,N_14870);
xor UO_1988 (O_1988,N_14859,N_14970);
nor UO_1989 (O_1989,N_14955,N_14923);
nor UO_1990 (O_1990,N_14828,N_14850);
nor UO_1991 (O_1991,N_14933,N_14998);
and UO_1992 (O_1992,N_14974,N_14976);
nor UO_1993 (O_1993,N_14826,N_14887);
xnor UO_1994 (O_1994,N_14897,N_14885);
nor UO_1995 (O_1995,N_14855,N_14880);
nor UO_1996 (O_1996,N_14801,N_14813);
xor UO_1997 (O_1997,N_14976,N_14991);
nand UO_1998 (O_1998,N_14835,N_14896);
nand UO_1999 (O_1999,N_14815,N_14853);
endmodule