module basic_3000_30000_3500_5_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_1734,In_143);
and U1 (N_1,In_154,In_1614);
nand U2 (N_2,In_1357,In_673);
xor U3 (N_3,In_613,In_2142);
and U4 (N_4,In_724,In_2315);
and U5 (N_5,In_815,In_2076);
nand U6 (N_6,In_245,In_2166);
and U7 (N_7,In_2106,In_2017);
or U8 (N_8,In_2697,In_78);
and U9 (N_9,In_2080,In_284);
nor U10 (N_10,In_763,In_1186);
nand U11 (N_11,In_2370,In_972);
nand U12 (N_12,In_2626,In_1711);
xnor U13 (N_13,In_865,In_2871);
and U14 (N_14,In_988,In_781);
nand U15 (N_15,In_1178,In_1298);
and U16 (N_16,In_2783,In_380);
nand U17 (N_17,In_2174,In_2978);
nor U18 (N_18,In_1330,In_2171);
and U19 (N_19,In_1954,In_877);
xnor U20 (N_20,In_417,In_158);
and U21 (N_21,In_180,In_99);
nand U22 (N_22,In_49,In_1724);
or U23 (N_23,In_429,In_23);
and U24 (N_24,In_1796,In_1717);
nand U25 (N_25,In_2696,In_2599);
and U26 (N_26,In_1538,In_2642);
or U27 (N_27,In_1755,In_2348);
or U28 (N_28,In_309,In_1608);
and U29 (N_29,In_490,In_1226);
or U30 (N_30,In_226,In_1552);
nand U31 (N_31,In_2590,In_293);
nor U32 (N_32,In_1514,In_460);
nand U33 (N_33,In_2369,In_616);
or U34 (N_34,In_2896,In_466);
nor U35 (N_35,In_1183,In_1117);
nand U36 (N_36,In_1038,In_2732);
nor U37 (N_37,In_981,In_2655);
xor U38 (N_38,In_1697,In_710);
and U39 (N_39,In_777,In_268);
or U40 (N_40,In_2149,In_1780);
nor U41 (N_41,In_1750,In_393);
nand U42 (N_42,In_2193,In_517);
nand U43 (N_43,In_2200,In_739);
and U44 (N_44,In_1549,In_1285);
nor U45 (N_45,In_141,In_975);
and U46 (N_46,In_125,In_1221);
and U47 (N_47,In_2102,In_2976);
xor U48 (N_48,In_1544,In_1385);
nand U49 (N_49,In_1577,In_1134);
or U50 (N_50,In_1363,In_906);
nand U51 (N_51,In_939,In_2298);
xor U52 (N_52,In_2961,In_860);
or U53 (N_53,In_1191,In_2343);
nand U54 (N_54,In_964,In_2859);
nor U55 (N_55,In_2714,In_894);
and U56 (N_56,In_1065,In_822);
xnor U57 (N_57,In_1873,In_2529);
and U58 (N_58,In_1599,In_1881);
nand U59 (N_59,In_2033,In_1740);
or U60 (N_60,In_2353,In_238);
nor U61 (N_61,In_1885,In_1259);
or U62 (N_62,In_2734,In_152);
xnor U63 (N_63,In_1797,In_2205);
or U64 (N_64,In_2606,In_830);
xnor U65 (N_65,In_884,In_1895);
or U66 (N_66,In_473,In_139);
or U67 (N_67,In_1069,In_2693);
or U68 (N_68,In_2989,In_1580);
xnor U69 (N_69,In_1723,In_1371);
or U70 (N_70,In_1367,In_2746);
xor U71 (N_71,In_113,In_2145);
xor U72 (N_72,In_151,In_2761);
nand U73 (N_73,In_2889,In_2270);
nand U74 (N_74,In_730,In_1477);
xnor U75 (N_75,In_1961,In_991);
nor U76 (N_76,In_2810,In_2706);
and U77 (N_77,In_622,In_2891);
nor U78 (N_78,In_553,In_1142);
nand U79 (N_79,In_270,In_169);
and U80 (N_80,In_802,In_1389);
xnor U81 (N_81,In_2533,In_493);
or U82 (N_82,In_838,In_544);
or U83 (N_83,In_2070,In_2436);
and U84 (N_84,In_2757,In_161);
and U85 (N_85,In_1453,In_2640);
or U86 (N_86,In_1773,In_1659);
xnor U87 (N_87,In_587,In_664);
nor U88 (N_88,In_891,In_29);
xnor U89 (N_89,In_1391,In_127);
nor U90 (N_90,In_1665,In_1624);
xor U91 (N_91,In_661,In_997);
nand U92 (N_92,In_2024,In_2897);
and U93 (N_93,In_829,In_1039);
and U94 (N_94,In_649,In_131);
nor U95 (N_95,In_532,In_2739);
xor U96 (N_96,In_1052,In_1027);
nor U97 (N_97,In_2015,In_2493);
xor U98 (N_98,In_1297,In_538);
nand U99 (N_99,In_346,In_465);
nor U100 (N_100,In_1299,In_1806);
and U101 (N_101,In_2737,In_1700);
and U102 (N_102,In_1026,In_2705);
nand U103 (N_103,In_770,In_966);
nand U104 (N_104,In_1889,In_1855);
or U105 (N_105,In_1013,In_419);
or U106 (N_106,In_976,In_344);
or U107 (N_107,In_1025,In_1958);
nand U108 (N_108,In_1653,In_1572);
nand U109 (N_109,In_2484,In_2302);
and U110 (N_110,In_381,In_1946);
and U111 (N_111,In_2090,In_1318);
and U112 (N_112,In_2314,In_2750);
or U113 (N_113,In_1319,In_2621);
xor U114 (N_114,In_2821,In_1105);
and U115 (N_115,In_88,In_1609);
xnor U116 (N_116,In_2403,In_2176);
and U117 (N_117,In_1392,In_513);
nor U118 (N_118,In_2313,In_2502);
nand U119 (N_119,In_2797,In_391);
nand U120 (N_120,In_2569,In_2341);
nor U121 (N_121,In_700,In_787);
or U122 (N_122,In_1587,In_2733);
nand U123 (N_123,In_2584,In_2300);
xor U124 (N_124,In_1625,In_520);
or U125 (N_125,In_2084,In_2187);
xnor U126 (N_126,In_1422,In_842);
xor U127 (N_127,In_1686,In_507);
xnor U128 (N_128,In_157,In_2636);
nor U129 (N_129,In_1467,In_747);
nand U130 (N_130,In_2937,In_2306);
or U131 (N_131,In_2855,In_349);
and U132 (N_132,In_1277,In_1059);
nand U133 (N_133,In_1411,In_1045);
or U134 (N_134,In_1541,In_1209);
and U135 (N_135,In_2656,In_212);
xor U136 (N_136,In_1671,In_1485);
or U137 (N_137,In_825,In_1111);
and U138 (N_138,In_1462,In_1000);
nor U139 (N_139,In_383,In_1339);
nor U140 (N_140,In_2127,In_742);
nand U141 (N_141,In_1014,In_2620);
nand U142 (N_142,In_633,In_2443);
xnor U143 (N_143,In_1581,In_2267);
or U144 (N_144,In_2924,In_2181);
or U145 (N_145,In_2688,In_364);
nor U146 (N_146,In_215,In_2373);
nor U147 (N_147,In_118,In_2602);
nand U148 (N_148,In_2472,In_1839);
and U149 (N_149,In_47,In_2483);
nor U150 (N_150,In_200,In_969);
xor U151 (N_151,In_1658,In_679);
xnor U152 (N_152,In_279,In_1493);
xor U153 (N_153,In_436,In_2492);
nand U154 (N_154,In_467,In_1057);
nand U155 (N_155,In_1271,In_1560);
nor U156 (N_156,In_1822,In_2622);
nand U157 (N_157,In_691,In_2180);
xnor U158 (N_158,In_2985,In_2049);
and U159 (N_159,In_2239,In_2144);
or U160 (N_160,In_222,In_1669);
and U161 (N_161,In_2233,In_1368);
or U162 (N_162,In_2241,In_1239);
nand U163 (N_163,In_808,In_1325);
nor U164 (N_164,In_1850,In_863);
nor U165 (N_165,In_290,In_937);
nand U166 (N_166,In_1730,In_2653);
nand U167 (N_167,In_2922,In_993);
or U168 (N_168,In_2381,In_2154);
and U169 (N_169,In_1116,In_1691);
nand U170 (N_170,In_2147,In_2574);
nand U171 (N_171,In_923,In_2929);
and U172 (N_172,In_2872,In_271);
nor U173 (N_173,In_2765,In_2422);
and U174 (N_174,In_67,In_1611);
and U175 (N_175,In_930,In_892);
or U176 (N_176,In_1964,In_2069);
nand U177 (N_177,In_322,In_1425);
or U178 (N_178,In_168,In_1194);
nand U179 (N_179,In_2707,In_2695);
nor U180 (N_180,In_2034,In_2344);
and U181 (N_181,In_2044,In_1820);
and U182 (N_182,In_1531,In_1306);
nor U183 (N_183,In_2444,In_1491);
and U184 (N_184,In_1103,In_1991);
nor U185 (N_185,In_2384,In_2950);
and U186 (N_186,In_371,In_1787);
nand U187 (N_187,In_504,In_713);
and U188 (N_188,In_1720,In_35);
and U189 (N_189,In_1504,In_382);
or U190 (N_190,In_2579,In_1547);
xnor U191 (N_191,In_90,In_2236);
or U192 (N_192,In_1989,In_2984);
and U193 (N_193,In_2235,In_1509);
and U194 (N_194,In_2994,In_2775);
or U195 (N_195,In_515,In_1451);
nor U196 (N_196,In_1551,In_1423);
nor U197 (N_197,In_1350,In_254);
nor U198 (N_198,In_185,In_1561);
or U199 (N_199,In_1250,In_1144);
xor U200 (N_200,In_859,In_2611);
and U201 (N_201,In_2108,In_1594);
and U202 (N_202,In_1415,In_395);
and U203 (N_203,In_1395,In_117);
or U204 (N_204,In_778,In_2466);
and U205 (N_205,In_1706,In_1699);
xor U206 (N_206,In_2433,In_1182);
nand U207 (N_207,In_999,In_1534);
xnor U208 (N_208,In_1129,In_2223);
xnor U209 (N_209,In_1761,In_1905);
nor U210 (N_210,In_1124,In_288);
nor U211 (N_211,In_1163,In_2956);
nor U212 (N_212,In_1113,In_1323);
and U213 (N_213,In_75,In_1987);
or U214 (N_214,In_2694,In_2575);
and U215 (N_215,In_1344,In_2587);
nand U216 (N_216,In_2375,In_1083);
nor U217 (N_217,In_1651,In_2368);
and U218 (N_218,In_2639,In_2346);
and U219 (N_219,In_281,In_0);
xor U220 (N_220,In_2046,In_935);
nand U221 (N_221,In_2586,In_170);
or U222 (N_222,In_1386,In_1212);
and U223 (N_223,In_1604,In_588);
and U224 (N_224,In_2992,In_363);
nor U225 (N_225,In_1909,In_632);
and U226 (N_226,In_1364,In_2197);
xor U227 (N_227,In_1102,In_480);
and U228 (N_228,In_1936,In_2411);
or U229 (N_229,In_2280,In_568);
and U230 (N_230,In_2162,In_1630);
and U231 (N_231,In_235,In_2323);
and U232 (N_232,In_489,In_2850);
nor U233 (N_233,In_130,In_1655);
and U234 (N_234,In_1536,In_2613);
or U235 (N_235,In_2552,In_1864);
xnor U236 (N_236,In_1836,In_2505);
nor U237 (N_237,In_2204,In_2629);
nand U238 (N_238,In_1372,In_602);
or U239 (N_239,In_1061,In_1390);
nand U240 (N_240,In_2150,In_1605);
xor U241 (N_241,In_74,In_1060);
nor U242 (N_242,In_1921,In_1986);
nand U243 (N_243,In_873,In_1776);
xnor U244 (N_244,In_753,In_427);
or U245 (N_245,In_1104,In_1248);
nor U246 (N_246,In_654,In_2951);
nor U247 (N_247,In_338,In_2271);
nand U248 (N_248,In_1128,In_627);
nand U249 (N_249,In_64,In_87);
or U250 (N_250,In_2349,In_1701);
and U251 (N_251,In_2207,In_1698);
nor U252 (N_252,In_1644,In_1400);
or U253 (N_253,In_2703,In_2038);
nor U254 (N_254,In_2843,In_2192);
or U255 (N_255,In_2806,In_2066);
or U256 (N_256,In_2648,In_618);
nand U257 (N_257,In_1783,In_1089);
nand U258 (N_258,In_453,In_2234);
or U259 (N_259,In_2059,In_85);
and U260 (N_260,In_2926,In_18);
and U261 (N_261,In_324,In_1728);
nand U262 (N_262,In_1643,In_2727);
nor U263 (N_263,In_2345,In_2949);
or U264 (N_264,In_2633,In_58);
nor U265 (N_265,In_1088,In_2331);
or U266 (N_266,In_2525,In_596);
nor U267 (N_267,In_2374,In_2141);
or U268 (N_268,In_2818,In_1677);
and U269 (N_269,In_2460,In_2933);
or U270 (N_270,In_631,In_1276);
nor U271 (N_271,In_225,In_949);
and U272 (N_272,In_2216,In_2161);
xor U273 (N_273,In_1165,In_2588);
xor U274 (N_274,In_876,In_598);
nor U275 (N_275,In_2284,In_2258);
xnor U276 (N_276,In_2538,In_2519);
xnor U277 (N_277,In_2486,In_2152);
xor U278 (N_278,In_172,In_38);
and U279 (N_279,In_784,In_1374);
xnor U280 (N_280,In_16,In_2837);
xnor U281 (N_281,In_249,In_2925);
xnor U282 (N_282,In_1281,In_86);
nand U283 (N_283,In_2095,In_1465);
or U284 (N_284,In_2708,In_1583);
or U285 (N_285,In_2857,In_1064);
and U286 (N_286,In_2036,In_379);
or U287 (N_287,In_576,In_672);
xnor U288 (N_288,In_670,In_252);
and U289 (N_289,In_500,In_2467);
nand U290 (N_290,In_1931,In_1246);
nor U291 (N_291,In_1661,In_1775);
nor U292 (N_292,In_2893,In_2308);
nand U293 (N_293,In_2347,In_1859);
nand U294 (N_294,In_1084,In_183);
nor U295 (N_295,In_901,In_703);
xnor U296 (N_296,In_2082,In_2330);
nor U297 (N_297,In_2395,In_893);
nor U298 (N_298,In_1854,In_1469);
or U299 (N_299,In_1406,In_1336);
nand U300 (N_300,In_297,In_1741);
nand U301 (N_301,In_2900,In_1497);
nand U302 (N_302,In_96,In_1366);
xor U303 (N_303,In_1672,In_209);
and U304 (N_304,In_1004,In_913);
or U305 (N_305,In_2825,In_1204);
or U306 (N_306,In_2337,In_370);
and U307 (N_307,In_927,In_2740);
nor U308 (N_308,In_1159,In_1891);
nor U309 (N_309,In_2698,In_606);
nand U310 (N_310,In_1109,In_1795);
and U311 (N_311,In_1307,In_316);
or U312 (N_312,In_1179,In_1982);
xor U313 (N_313,In_1526,In_779);
nand U314 (N_314,In_932,In_1066);
nor U315 (N_315,In_1043,In_793);
xor U316 (N_316,In_2332,In_1751);
and U317 (N_317,In_193,In_1589);
nor U318 (N_318,In_174,In_856);
and U319 (N_319,In_1825,In_601);
and U320 (N_320,In_1505,In_2260);
and U321 (N_321,In_1768,In_2682);
nor U322 (N_322,In_1649,In_1716);
nor U323 (N_323,In_61,In_1757);
or U324 (N_324,In_2317,In_1499);
nand U325 (N_325,In_599,In_1475);
xor U326 (N_326,In_1814,In_2838);
xnor U327 (N_327,In_503,In_237);
xnor U328 (N_328,In_496,In_529);
xnor U329 (N_329,In_1238,In_2126);
and U330 (N_330,In_2400,In_2730);
nand U331 (N_331,In_228,In_628);
and U332 (N_332,In_2990,In_2385);
and U333 (N_333,In_315,In_229);
nand U334 (N_334,In_1115,In_548);
or U335 (N_335,In_399,In_800);
xnor U336 (N_336,In_2352,In_1100);
nand U337 (N_337,In_2183,In_2670);
and U338 (N_338,In_552,In_1362);
or U339 (N_339,In_2995,In_2229);
xnor U340 (N_340,In_509,In_2652);
or U341 (N_341,In_1040,In_786);
nand U342 (N_342,In_1253,In_1222);
nor U343 (N_343,In_2096,In_1590);
xnor U344 (N_344,In_2848,In_1567);
xor U345 (N_345,In_2173,In_746);
and U346 (N_346,In_2829,In_744);
or U347 (N_347,In_1992,In_1145);
nand U348 (N_348,In_2041,In_2383);
nor U349 (N_349,In_928,In_1606);
or U350 (N_350,In_2788,In_1180);
or U351 (N_351,In_2953,In_1463);
xnor U352 (N_352,In_512,In_216);
and U353 (N_353,In_2558,In_1602);
nor U354 (N_354,In_253,In_723);
nand U355 (N_355,In_2111,In_2190);
xor U356 (N_356,In_1715,In_709);
nor U357 (N_357,In_2282,In_2310);
xor U358 (N_358,In_1530,In_2364);
nand U359 (N_359,In_1947,In_2269);
and U360 (N_360,In_1130,In_374);
and U361 (N_361,In_667,In_1024);
xnor U362 (N_362,In_103,In_1945);
nand U363 (N_363,In_1804,In_2491);
nand U364 (N_364,In_1305,In_948);
nand U365 (N_365,In_2944,In_129);
or U366 (N_366,In_2219,In_402);
or U367 (N_367,In_2971,In_905);
or U368 (N_368,In_2918,In_1170);
nor U369 (N_369,In_2378,In_2701);
nor U370 (N_370,In_1403,In_824);
nor U371 (N_371,In_2307,In_1232);
xnor U372 (N_372,In_2334,In_708);
nand U373 (N_373,In_1634,In_1472);
xnor U374 (N_374,In_2093,In_11);
nand U375 (N_375,In_2203,In_921);
nand U376 (N_376,In_806,In_1245);
nand U377 (N_377,In_745,In_401);
and U378 (N_378,In_2661,In_1553);
nand U379 (N_379,In_1459,In_2517);
and U380 (N_380,In_1094,In_2465);
or U381 (N_381,In_1431,In_2665);
xor U382 (N_382,In_2932,In_790);
or U383 (N_383,In_2781,In_275);
and U384 (N_384,In_411,In_1304);
xor U385 (N_385,In_21,In_1763);
nand U386 (N_386,In_2225,In_2780);
and U387 (N_387,In_2342,In_261);
xnor U388 (N_388,In_2565,In_2202);
nand U389 (N_389,In_2631,In_2055);
nor U390 (N_390,In_725,In_2299);
nand U391 (N_391,In_1028,In_2787);
or U392 (N_392,In_2774,In_2582);
or U393 (N_393,In_1901,In_721);
nor U394 (N_394,In_1402,In_2014);
or U395 (N_395,In_95,In_2265);
or U396 (N_396,In_2451,In_239);
nor U397 (N_397,In_2035,In_428);
xnor U398 (N_398,In_1164,In_2886);
nor U399 (N_399,In_1171,In_313);
xor U400 (N_400,In_1597,In_1545);
or U401 (N_401,In_2720,In_2304);
nand U402 (N_402,In_128,In_2715);
and U403 (N_403,In_1108,In_1537);
or U404 (N_404,In_1973,In_37);
and U405 (N_405,In_1237,In_486);
and U406 (N_406,In_276,In_1788);
nand U407 (N_407,In_651,In_1527);
or U408 (N_408,In_2567,In_1569);
nand U409 (N_409,In_1484,In_1160);
or U410 (N_410,In_760,In_983);
xor U411 (N_411,In_488,In_2755);
xor U412 (N_412,In_1879,In_219);
xor U413 (N_413,In_1338,In_2853);
and U414 (N_414,In_1049,In_1322);
xnor U415 (N_415,In_116,In_2133);
xor U416 (N_416,In_541,In_2407);
or U417 (N_417,In_1247,In_1202);
xor U418 (N_418,In_765,In_280);
nor U419 (N_419,In_1360,In_2598);
nand U420 (N_420,In_823,In_1923);
and U421 (N_421,In_456,In_1161);
or U422 (N_422,In_1007,In_1878);
nand U423 (N_423,In_2075,In_2297);
nor U424 (N_424,In_312,In_2120);
nor U425 (N_425,In_1439,In_1990);
nor U426 (N_426,In_491,In_2541);
nand U427 (N_427,In_984,In_333);
or U428 (N_428,In_1495,In_1019);
or U429 (N_429,In_1511,In_821);
or U430 (N_430,In_1072,In_2641);
nand U431 (N_431,In_484,In_2293);
and U432 (N_432,In_2646,In_2228);
or U433 (N_433,In_2431,In_1994);
nand U434 (N_434,In_1983,In_2420);
or U435 (N_435,In_858,In_1261);
xnor U436 (N_436,In_1888,In_307);
and U437 (N_437,In_140,In_1264);
nor U438 (N_438,In_2842,In_2296);
xor U439 (N_439,In_1224,In_2288);
or U440 (N_440,In_2717,In_2356);
nor U441 (N_441,In_586,In_1967);
xor U442 (N_442,In_846,In_2500);
and U443 (N_443,In_2912,In_973);
and U444 (N_444,In_1413,In_1009);
or U445 (N_445,In_866,In_1834);
nand U446 (N_446,In_81,In_1846);
or U447 (N_447,In_1693,In_2930);
or U448 (N_448,In_1290,In_164);
nand U449 (N_449,In_2585,In_1582);
nand U450 (N_450,In_1151,In_2092);
nor U451 (N_451,In_389,In_1195);
and U452 (N_452,In_2559,In_1107);
nor U453 (N_453,In_224,In_2894);
and U454 (N_454,In_2191,In_817);
and U455 (N_455,In_2058,In_1613);
nand U456 (N_456,In_899,In_39);
xor U457 (N_457,In_89,In_916);
or U458 (N_458,In_2964,In_968);
or U459 (N_459,In_1914,In_471);
nand U460 (N_460,In_1865,In_2328);
xor U461 (N_461,In_2913,In_2001);
or U462 (N_462,In_1317,In_2179);
or U463 (N_463,In_111,In_347);
nor U464 (N_464,In_1926,In_740);
or U465 (N_465,In_1566,In_1791);
and U466 (N_466,In_2089,In_595);
or U467 (N_467,In_1263,In_688);
nand U468 (N_468,In_2372,In_1838);
and U469 (N_469,In_1205,In_1880);
nor U470 (N_470,In_2594,In_296);
or U471 (N_471,In_2634,In_295);
or U472 (N_472,In_1042,In_625);
and U473 (N_473,In_241,In_54);
or U474 (N_474,In_2283,In_551);
xor U475 (N_475,In_1727,In_286);
xor U476 (N_476,In_878,In_1764);
and U477 (N_477,In_2657,In_1162);
and U478 (N_478,In_845,In_867);
or U479 (N_479,In_52,In_2865);
nor U480 (N_480,In_2019,In_1922);
and U481 (N_481,In_2266,In_1192);
or U482 (N_482,In_1736,In_2454);
xor U483 (N_483,In_1588,In_326);
xnor U484 (N_484,In_2844,In_1435);
and U485 (N_485,In_2387,In_1296);
and U486 (N_486,In_208,In_2521);
and U487 (N_487,In_2716,In_1749);
and U488 (N_488,In_2851,In_1240);
nor U489 (N_489,In_1352,In_2819);
nor U490 (N_490,In_2278,In_1707);
xnor U491 (N_491,In_794,In_1507);
or U492 (N_492,In_1396,In_1220);
or U493 (N_493,In_962,In_378);
and U494 (N_494,In_2286,In_273);
xor U495 (N_495,In_1705,In_2908);
nor U496 (N_496,In_868,In_9);
nand U497 (N_497,In_2498,In_2263);
nor U498 (N_498,In_423,In_1678);
and U499 (N_499,In_850,In_283);
nor U500 (N_500,In_2881,In_1355);
nor U501 (N_501,In_2380,In_361);
and U502 (N_502,In_2290,In_1458);
nor U503 (N_503,In_652,In_535);
and U504 (N_504,In_2856,In_1617);
nor U505 (N_505,In_2247,In_629);
or U506 (N_506,In_2792,In_248);
nor U507 (N_507,In_1255,In_348);
or U508 (N_508,In_681,In_619);
xor U509 (N_509,In_1486,In_1976);
nor U510 (N_510,In_108,In_656);
and U511 (N_511,In_883,In_2097);
nand U512 (N_512,In_1652,In_1139);
xnor U513 (N_513,In_126,In_2532);
nand U514 (N_514,In_15,In_2866);
nand U515 (N_515,In_34,In_2244);
nor U516 (N_516,In_1710,In_310);
or U517 (N_517,In_2899,In_2595);
and U518 (N_518,In_2610,In_2005);
or U519 (N_519,In_704,In_2416);
and U520 (N_520,In_1970,In_958);
and U521 (N_521,In_2068,In_1067);
xor U522 (N_522,In_1433,In_2604);
nand U523 (N_523,In_2251,In_1384);
nand U524 (N_524,In_365,In_826);
nand U525 (N_525,In_1558,In_2736);
or U526 (N_526,In_2042,In_1616);
nand U527 (N_527,In_1133,In_2404);
xor U528 (N_528,In_2421,In_2554);
nor U529 (N_529,In_1863,In_1030);
or U530 (N_530,In_944,In_2849);
xnor U531 (N_531,In_2966,In_2794);
nand U532 (N_532,In_1470,In_2677);
or U533 (N_533,In_274,In_2581);
nor U534 (N_534,In_2531,In_2281);
nor U535 (N_535,In_2450,In_676);
nand U536 (N_536,In_2801,In_481);
or U537 (N_537,In_617,In_2608);
xor U538 (N_538,In_63,In_2875);
and U539 (N_539,In_1852,In_580);
xor U540 (N_540,In_615,In_257);
xor U541 (N_541,In_1610,In_1326);
nand U542 (N_542,In_440,In_2895);
nand U543 (N_543,In_2000,In_2238);
or U544 (N_544,In_1550,In_243);
and U545 (N_545,In_2743,In_1965);
nor U546 (N_546,In_592,In_1944);
xnor U547 (N_547,In_2603,In_2940);
or U548 (N_548,In_1432,In_2366);
nand U549 (N_549,In_2528,In_1904);
nor U550 (N_550,In_2045,In_841);
or U551 (N_551,In_2729,In_2430);
or U552 (N_552,In_2030,In_2563);
nand U553 (N_553,In_812,In_1301);
or U554 (N_554,In_839,In_1910);
nand U555 (N_555,In_1951,In_2578);
xnor U556 (N_556,In_398,In_1011);
and U557 (N_557,In_2556,In_737);
nor U558 (N_558,In_521,In_2685);
nand U559 (N_559,In_2259,In_265);
xor U560 (N_560,In_1770,In_2536);
nor U561 (N_561,In_1099,In_356);
and U562 (N_562,In_1,In_149);
and U563 (N_563,In_630,In_31);
nand U564 (N_564,In_678,In_2607);
nand U565 (N_565,In_2333,In_518);
and U566 (N_566,In_819,In_769);
and U567 (N_567,In_2305,In_1473);
xor U568 (N_568,In_1682,In_115);
nand U569 (N_569,In_2083,In_1618);
or U570 (N_570,In_2128,In_420);
and U571 (N_571,In_1450,In_2250);
or U572 (N_572,In_2675,In_1681);
or U573 (N_573,In_2210,In_2906);
nand U574 (N_574,In_2021,In_918);
nand U575 (N_575,In_2398,In_441);
nor U576 (N_576,In_1157,In_526);
and U577 (N_577,In_358,In_795);
xnor U578 (N_578,In_2485,In_1466);
xnor U579 (N_579,In_530,In_264);
xnor U580 (N_580,In_776,In_773);
and U581 (N_581,In_3,In_614);
xnor U582 (N_582,In_1310,In_221);
nor U583 (N_583,In_1327,In_2619);
nor U584 (N_584,In_566,In_202);
or U585 (N_585,In_19,In_1862);
nand U586 (N_586,In_2911,In_2742);
or U587 (N_587,In_1794,In_2338);
or U588 (N_588,In_2617,In_1977);
or U589 (N_589,In_100,In_2934);
nor U590 (N_590,In_1078,In_611);
nand U591 (N_591,In_121,In_2800);
nor U592 (N_592,In_2119,In_2509);
or U593 (N_593,In_693,In_1427);
or U594 (N_594,In_2987,In_83);
and U595 (N_595,In_53,In_259);
and U596 (N_596,In_455,In_1956);
xor U597 (N_597,In_1335,In_2980);
nor U598 (N_598,In_2923,In_22);
or U599 (N_599,In_181,In_1314);
xor U600 (N_600,In_1844,In_1426);
nand U601 (N_601,In_926,In_743);
nand U602 (N_602,In_1437,In_1942);
xnor U603 (N_603,In_1037,In_1792);
nor U604 (N_604,In_1382,In_1405);
and U605 (N_605,In_1900,In_2751);
or U606 (N_606,In_2319,In_2516);
or U607 (N_607,In_1207,In_1571);
or U608 (N_608,In_1490,In_938);
nor U609 (N_609,In_20,In_422);
nand U610 (N_610,In_1288,In_2678);
nor U611 (N_611,In_2327,In_731);
nand U612 (N_612,In_1725,In_1647);
and U613 (N_613,In_1826,In_575);
xnor U614 (N_614,In_1809,In_1200);
nand U615 (N_615,In_2760,In_687);
or U616 (N_616,In_2294,In_56);
nor U617 (N_617,In_2452,In_2053);
or U618 (N_618,In_853,In_2429);
and U619 (N_619,In_772,In_2916);
and U620 (N_620,In_1801,In_2836);
nand U621 (N_621,In_2628,In_2996);
and U622 (N_622,In_766,In_946);
and U623 (N_623,In_1096,In_107);
xnor U624 (N_624,In_1920,In_2101);
and U625 (N_625,In_959,In_2960);
and U626 (N_626,In_1482,In_2943);
and U627 (N_627,In_1735,In_167);
xor U628 (N_628,In_2459,In_2275);
xnor U629 (N_629,In_1230,In_1154);
nand U630 (N_630,In_2812,In_1216);
xnor U631 (N_631,In_1337,In_2165);
nand U632 (N_632,In_1690,In_2870);
or U633 (N_633,In_2237,In_2440);
or U634 (N_634,In_386,In_2335);
xnor U635 (N_635,In_522,In_2272);
nor U636 (N_636,In_909,In_1023);
nor U637 (N_637,In_2303,In_188);
or U638 (N_638,In_726,In_1265);
nand U639 (N_639,In_2888,In_1752);
and U640 (N_640,In_246,In_2882);
or U641 (N_641,In_2159,In_1676);
nand U642 (N_642,In_2770,In_1316);
nand U643 (N_643,In_1022,In_2555);
and U644 (N_644,In_203,In_1995);
and U645 (N_645,In_929,In_2462);
or U646 (N_646,In_2013,In_2724);
or U647 (N_647,In_2194,In_2248);
nor U648 (N_648,In_2679,In_1044);
nand U649 (N_649,In_2487,In_250);
or U650 (N_650,In_2564,In_1197);
and U651 (N_651,In_1919,In_1903);
or U652 (N_652,In_771,In_712);
or U653 (N_653,In_2287,In_1913);
and U654 (N_654,In_1917,In_655);
nor U655 (N_655,In_556,In_1442);
or U656 (N_656,In_1784,In_1097);
nand U657 (N_657,In_992,In_416);
or U658 (N_658,In_2993,In_2975);
or U659 (N_659,In_2292,In_272);
and U660 (N_660,In_2363,In_2835);
and U661 (N_661,In_397,In_1443);
or U662 (N_662,In_317,In_1817);
or U663 (N_663,In_1687,In_2003);
xnor U664 (N_664,In_2658,In_1623);
xnor U665 (N_665,In_919,In_2507);
xnor U666 (N_666,In_71,In_1694);
or U667 (N_667,In_1745,In_2719);
nor U668 (N_668,In_1759,In_1866);
nand U669 (N_669,In_782,In_979);
nand U670 (N_670,In_621,In_2309);
or U671 (N_671,In_2168,In_211);
and U672 (N_672,In_707,In_1765);
and U673 (N_673,In_232,In_646);
or U674 (N_674,In_996,In_1122);
and U675 (N_675,In_1629,In_2064);
and U676 (N_676,In_2490,In_2249);
nor U677 (N_677,In_908,In_204);
and U678 (N_678,In_2718,In_482);
and U679 (N_679,In_705,In_1869);
or U680 (N_680,In_2222,In_1034);
and U681 (N_681,In_626,In_980);
xnor U682 (N_682,In_26,In_2568);
nor U683 (N_683,In_1648,In_199);
xor U684 (N_684,In_792,In_2645);
nor U685 (N_685,In_1234,In_1279);
nand U686 (N_686,In_1141,In_2768);
xnor U687 (N_687,In_2240,In_377);
or U688 (N_688,In_1448,In_1815);
or U689 (N_689,In_683,In_171);
or U690 (N_690,In_2977,In_634);
nor U691 (N_691,In_1960,In_2816);
and U692 (N_692,In_1521,In_462);
nor U693 (N_693,In_1464,In_412);
xnor U694 (N_694,In_2405,In_162);
nor U695 (N_695,In_319,In_2877);
xnor U696 (N_696,In_2057,In_2771);
and U697 (N_697,In_2684,In_1660);
xnor U698 (N_698,In_2741,In_159);
nand U699 (N_699,In_1997,In_1563);
nand U700 (N_700,In_2143,In_585);
nor U701 (N_701,In_2418,In_2644);
nand U702 (N_702,In_648,In_2435);
nand U703 (N_703,In_701,In_332);
xnor U704 (N_704,In_2043,In_2545);
nand U705 (N_705,In_692,In_328);
nor U706 (N_706,In_2605,In_2583);
nand U707 (N_707,In_1053,In_2530);
and U708 (N_708,In_2311,In_1378);
or U709 (N_709,In_2596,In_1150);
and U710 (N_710,In_1166,In_2826);
nor U711 (N_711,In_2273,In_155);
xor U712 (N_712,In_936,In_1308);
and U713 (N_713,In_24,In_549);
or U714 (N_714,In_1190,In_735);
xor U715 (N_715,In_1399,In_593);
nor U716 (N_716,In_1236,In_813);
nand U717 (N_717,In_50,In_1887);
or U718 (N_718,In_1762,In_1208);
or U719 (N_719,In_2185,In_2105);
xor U720 (N_720,In_2773,In_1845);
nor U721 (N_721,In_367,In_896);
xor U722 (N_722,In_1918,In_612);
or U723 (N_723,In_2153,In_2321);
nand U724 (N_724,In_1106,In_4);
nand U725 (N_725,In_1401,In_134);
and U726 (N_726,In_355,In_345);
xnor U727 (N_727,In_80,In_2799);
or U728 (N_728,In_995,In_1972);
nand U729 (N_729,In_610,In_236);
and U730 (N_730,In_748,In_545);
xor U731 (N_731,In_682,In_485);
xor U732 (N_732,In_2350,In_340);
or U733 (N_733,In_2905,In_2938);
nand U734 (N_734,In_1167,In_519);
nand U735 (N_735,In_2052,In_1935);
and U736 (N_736,In_862,In_660);
or U737 (N_737,In_501,In_2686);
nand U738 (N_738,In_469,In_175);
nor U739 (N_739,In_194,In_59);
nor U740 (N_740,In_2107,In_2878);
and U741 (N_741,In_2803,In_1930);
nand U742 (N_742,In_494,In_1487);
nand U743 (N_743,In_1980,In_2548);
xor U744 (N_744,In_1272,In_73);
nand U745 (N_745,In_2025,In_191);
and U746 (N_746,In_1137,In_2969);
nand U747 (N_747,In_953,In_1152);
nor U748 (N_748,In_437,In_1539);
xor U749 (N_749,In_540,In_2094);
and U750 (N_750,In_2473,In_1726);
and U751 (N_751,In_603,In_510);
and U752 (N_752,In_1685,In_334);
xnor U753 (N_753,In_2367,In_2109);
and U754 (N_754,In_109,In_1418);
xnor U755 (N_755,In_407,In_1667);
nor U756 (N_756,In_2104,In_1663);
nor U757 (N_757,In_1856,In_736);
nor U758 (N_758,In_1692,In_2478);
and U759 (N_759,In_233,In_2845);
nand U760 (N_760,In_516,In_106);
and U761 (N_761,In_1242,In_2769);
nand U762 (N_762,In_2291,In_2566);
nor U763 (N_763,In_1790,In_1585);
nor U764 (N_764,In_2573,In_2593);
nor U765 (N_765,In_2524,In_2201);
nand U766 (N_766,In_2456,In_583);
and U767 (N_767,In_350,In_1704);
xnor U768 (N_768,In_447,In_1502);
and U769 (N_769,In_2680,In_950);
nand U770 (N_770,In_1430,In_1388);
xor U771 (N_771,In_2073,In_1955);
nor U772 (N_772,In_1802,In_1321);
xnor U773 (N_773,In_2277,In_57);
or U774 (N_774,In_1419,In_2453);
or U775 (N_775,In_1136,In_1156);
or U776 (N_776,In_2553,In_1620);
nand U777 (N_777,In_2649,In_2537);
xnor U778 (N_778,In_767,In_578);
or U779 (N_779,In_122,In_2790);
nand U780 (N_780,In_182,In_5);
or U781 (N_781,In_711,In_2445);
nor U782 (N_782,In_2777,In_818);
or U783 (N_783,In_2496,In_2876);
xnor U784 (N_784,In_244,In_227);
or U785 (N_785,In_499,In_104);
nand U786 (N_786,In_717,In_1454);
or U787 (N_787,In_1214,In_2931);
xnor U788 (N_788,In_2160,In_1070);
nand U789 (N_789,In_439,In_1882);
and U790 (N_790,In_733,In_698);
nand U791 (N_791,In_849,In_2832);
and U792 (N_792,In_2060,In_1436);
and U793 (N_793,In_2785,In_562);
xor U794 (N_794,In_2245,In_458);
nor U795 (N_795,In_2006,In_1559);
nor U796 (N_796,In_2155,In_885);
xnor U797 (N_797,In_1680,In_2778);
and U798 (N_798,In_1848,In_1441);
xor U799 (N_799,In_805,In_1196);
and U800 (N_800,In_451,In_1833);
and U801 (N_801,In_220,In_537);
xnor U802 (N_802,In_2534,In_2032);
xor U803 (N_803,In_1050,In_2409);
or U804 (N_804,In_213,In_2632);
or U805 (N_805,In_299,In_647);
xor U806 (N_806,In_1055,In_1508);
nand U807 (N_807,In_525,In_957);
and U808 (N_808,In_2543,In_965);
xor U809 (N_809,In_2527,In_1957);
or U810 (N_810,In_2615,In_2252);
and U811 (N_811,In_2129,In_880);
or U812 (N_812,In_330,In_986);
or U813 (N_813,In_1598,In_722);
or U814 (N_814,In_360,In_951);
nand U815 (N_815,In_2175,In_1398);
or U816 (N_816,In_2514,In_413);
xor U817 (N_817,In_2379,In_2217);
xnor U818 (N_818,In_1421,In_1447);
or U819 (N_819,In_1688,In_25);
nor U820 (N_820,In_2455,In_637);
and U821 (N_821,In_2687,In_1274);
and U822 (N_822,In_2134,In_1235);
xor U823 (N_823,In_1835,In_1732);
and U824 (N_824,In_663,In_60);
and U825 (N_825,In_2901,In_2098);
nor U826 (N_826,In_2074,In_558);
or U827 (N_827,In_2791,In_2208);
nor U828 (N_828,In_2276,In_2660);
and U829 (N_829,In_650,In_954);
or U830 (N_830,In_2887,In_2029);
nor U831 (N_831,In_1703,In_2846);
xor U832 (N_832,In_445,In_1457);
xnor U833 (N_833,In_2752,In_847);
and U834 (N_834,In_1884,In_388);
or U835 (N_835,In_2962,In_1782);
nor U836 (N_836,In_1785,In_1636);
nand U837 (N_837,In_2963,In_1048);
or U838 (N_838,In_247,In_442);
or U839 (N_839,In_477,In_533);
and U840 (N_840,In_624,In_2412);
xnor U841 (N_841,In_1803,In_2196);
and U842 (N_842,In_1883,In_557);
and U843 (N_843,In_1718,In_2839);
xnor U844 (N_844,In_387,In_2841);
nor U845 (N_845,In_922,In_375);
nand U846 (N_846,In_69,In_1924);
nand U847 (N_847,In_1270,In_2442);
and U848 (N_848,In_2935,In_2668);
or U849 (N_849,In_797,In_1381);
or U850 (N_850,In_1894,In_1315);
nand U851 (N_851,In_2426,In_2065);
xnor U852 (N_852,In_1907,In_2419);
nand U853 (N_853,In_1471,In_809);
nand U854 (N_854,In_1331,In_2671);
nor U855 (N_855,In_871,In_2390);
nand U856 (N_856,In_2979,In_2699);
and U857 (N_857,In_1251,In_255);
nor U858 (N_858,In_1876,In_2039);
and U859 (N_859,In_2339,In_2007);
and U860 (N_860,In_2449,In_2731);
or U861 (N_861,In_2674,In_2071);
xor U862 (N_862,In_325,In_133);
and U863 (N_863,In_2156,In_881);
nand U864 (N_864,In_1294,In_904);
nor U865 (N_865,In_1506,In_2784);
nor U866 (N_866,In_1800,In_2061);
xor U867 (N_867,In_2079,In_101);
nor U868 (N_868,In_1090,In_353);
or U869 (N_869,In_8,In_2476);
xor U870 (N_870,In_1872,In_2561);
or U871 (N_871,In_1709,In_30);
or U872 (N_872,In_677,In_2464);
and U873 (N_873,In_1266,In_132);
and U874 (N_874,In_2508,In_2167);
and U875 (N_875,In_2137,In_1012);
nand U876 (N_876,In_1082,In_636);
xnor U877 (N_877,In_1786,In_1600);
nor U878 (N_878,In_1896,In_2869);
xnor U879 (N_879,In_342,In_2860);
nand U880 (N_880,In_875,In_1434);
nor U881 (N_881,In_716,In_2863);
nand U882 (N_882,In_2447,In_214);
or U883 (N_883,In_577,In_1601);
or U884 (N_884,In_42,In_1153);
or U885 (N_885,In_2828,In_961);
nor U886 (N_886,In_119,In_1091);
nand U887 (N_887,In_1131,In_2884);
and U888 (N_888,In_1123,In_1702);
and U889 (N_889,In_70,In_1959);
nand U890 (N_890,In_1348,In_828);
nand U891 (N_891,In_2215,In_2008);
nor U892 (N_892,In_1188,In_2898);
or U893 (N_893,In_240,In_1445);
xnor U894 (N_894,In_1177,In_2643);
or U895 (N_895,In_2982,In_2136);
and U896 (N_896,In_1908,In_392);
nor U897 (N_897,In_2638,In_2959);
nor U898 (N_898,In_2957,In_1747);
xor U899 (N_899,In_2544,In_2970);
xor U900 (N_900,In_148,In_1417);
nand U901 (N_901,In_2973,In_1767);
nand U902 (N_902,In_304,In_98);
or U903 (N_903,In_1810,In_339);
nor U904 (N_904,In_1857,In_2243);
nor U905 (N_905,In_1937,In_2804);
or U906 (N_906,In_1110,In_2786);
nor U907 (N_907,In_2009,In_2673);
nand U908 (N_908,In_84,In_1203);
and U909 (N_909,In_2213,In_1812);
nor U910 (N_910,In_2756,In_1596);
nor U911 (N_911,In_2285,In_1223);
or U912 (N_912,In_459,In_2023);
nand U913 (N_913,In_135,In_695);
nand U914 (N_914,In_1184,In_289);
and U915 (N_915,In_1591,In_1412);
nor U916 (N_916,In_1664,In_1404);
nand U917 (N_917,In_1148,In_1340);
nor U918 (N_918,In_385,In_1409);
nor U919 (N_919,In_2862,In_260);
or U920 (N_920,In_2766,In_690);
nand U921 (N_921,In_2002,In_1556);
and U922 (N_922,In_2939,In_1729);
nand U923 (N_923,In_33,In_1737);
xor U924 (N_924,In_1047,In_1939);
xor U925 (N_925,In_2112,In_2748);
and U926 (N_926,In_1564,In_879);
nand U927 (N_927,In_2438,In_1828);
nand U928 (N_928,In_2754,In_1743);
nand U929 (N_929,In_2355,In_2261);
nand U930 (N_930,In_197,In_2852);
nand U931 (N_931,In_1093,In_684);
and U932 (N_932,In_2209,In_464);
xor U933 (N_933,In_644,In_2782);
and U934 (N_934,In_1394,In_1354);
nand U935 (N_935,In_2099,In_2991);
xor U936 (N_936,In_799,In_1548);
or U937 (N_937,In_2488,In_2663);
xnor U938 (N_938,In_234,In_12);
and U939 (N_939,In_752,In_424);
and U940 (N_940,In_2609,In_1001);
nand U941 (N_941,In_2289,In_1218);
and U942 (N_942,In_2054,In_539);
nor U943 (N_943,In_1722,In_2242);
or U944 (N_944,In_1320,In_895);
or U945 (N_945,In_1546,In_2946);
and U946 (N_946,In_974,In_335);
nand U947 (N_947,In_1198,In_102);
and U948 (N_948,In_2518,In_1978);
or U949 (N_949,In_1377,In_294);
xor U950 (N_950,In_2212,In_699);
nand U951 (N_951,In_2691,In_357);
xor U952 (N_952,In_1387,In_1948);
nand U953 (N_953,In_1032,In_2480);
and U954 (N_954,In_1713,In_376);
nand U955 (N_955,In_1370,In_373);
nand U956 (N_956,In_1494,In_1628);
and U957 (N_957,In_1542,In_2712);
nand U958 (N_958,In_409,In_659);
nand U959 (N_959,In_685,In_1744);
or U960 (N_960,In_320,In_1565);
or U961 (N_961,In_1174,In_2662);
and U962 (N_962,In_584,In_2813);
nor U963 (N_963,In_2936,In_278);
nand U964 (N_964,In_51,In_1738);
and U965 (N_965,In_1906,In_1041);
xnor U966 (N_966,In_827,In_2986);
or U967 (N_967,In_1842,In_166);
or U968 (N_968,In_189,In_2279);
xnor U969 (N_969,In_2903,In_1853);
xnor U970 (N_970,In_341,In_1668);
nand U971 (N_971,In_1635,In_638);
nor U972 (N_972,In_474,In_1689);
and U973 (N_973,In_2955,In_914);
nand U974 (N_974,In_2914,In_2625);
xor U975 (N_975,In_438,In_2795);
nor U976 (N_976,In_144,In_756);
and U977 (N_977,In_2614,In_2199);
nand U978 (N_978,In_2376,In_1440);
and U979 (N_979,In_2031,In_1303);
xor U980 (N_980,In_351,In_2427);
nand U981 (N_981,In_2510,In_738);
nor U982 (N_982,In_2672,In_1515);
and U983 (N_983,In_1081,In_807);
or U984 (N_984,In_2700,In_689);
nor U985 (N_985,In_1353,In_2132);
and U986 (N_986,In_1293,In_1193);
nor U987 (N_987,In_72,In_1999);
or U988 (N_988,In_1811,In_764);
nor U989 (N_989,In_1533,In_2967);
and U990 (N_990,In_1941,In_933);
or U991 (N_991,In_2010,In_2214);
xor U992 (N_992,In_1974,In_775);
nand U993 (N_993,In_201,In_1851);
xnor U994 (N_994,In_694,In_1746);
nor U995 (N_995,In_1892,In_2811);
or U996 (N_996,In_804,In_2232);
xor U997 (N_997,In_196,In_1376);
nor U998 (N_998,In_1517,In_79);
or U999 (N_999,In_2169,In_2683);
or U1000 (N_1000,In_758,In_2227);
nor U1001 (N_1001,In_1169,In_639);
nand U1002 (N_1002,In_450,In_2831);
nand U1003 (N_1003,In_2468,In_256);
xor U1004 (N_1004,In_2413,In_366);
nand U1005 (N_1005,In_998,In_2198);
or U1006 (N_1006,In_1254,In_2779);
xnor U1007 (N_1007,In_536,In_2184);
xnor U1008 (N_1008,In_1805,In_882);
or U1009 (N_1009,In_1748,In_1932);
xnor U1010 (N_1010,In_1622,In_2088);
nor U1011 (N_1011,In_266,In_1575);
and U1012 (N_1012,In_2722,In_120);
xnor U1013 (N_1013,In_327,In_2504);
and U1014 (N_1014,In_2735,In_947);
xnor U1015 (N_1015,In_282,In_729);
and U1016 (N_1016,In_2354,In_1679);
nand U1017 (N_1017,In_2592,In_1615);
and U1018 (N_1018,In_2408,In_816);
nand U1019 (N_1019,In_508,In_1799);
and U1020 (N_1020,In_534,In_1492);
or U1021 (N_1021,In_1006,In_2549);
xnor U1022 (N_1022,In_680,In_1073);
and U1023 (N_1023,In_1953,In_1772);
xor U1024 (N_1024,In_2947,In_2325);
or U1025 (N_1025,In_314,In_205);
nor U1026 (N_1026,In_45,In_1176);
and U1027 (N_1027,In_1356,In_559);
nor U1028 (N_1028,In_2040,In_1474);
nor U1029 (N_1029,In_10,In_668);
or U1030 (N_1030,In_2246,In_1849);
nor U1031 (N_1031,In_594,In_2360);
nand U1032 (N_1032,In_1695,In_674);
nand U1033 (N_1033,In_1673,In_732);
nor U1034 (N_1034,In_1479,In_1126);
and U1035 (N_1035,In_2506,In_2158);
nand U1036 (N_1036,In_506,In_1674);
xor U1037 (N_1037,In_2113,In_1586);
and U1038 (N_1038,In_2262,In_1329);
or U1039 (N_1039,In_1684,In_1211);
and U1040 (N_1040,In_912,In_1095);
and U1041 (N_1041,In_872,In_55);
nand U1042 (N_1042,In_569,In_93);
nand U1043 (N_1043,In_1981,In_2499);
nor U1044 (N_1044,In_1574,In_2624);
xor U1045 (N_1045,In_1639,In_2711);
or U1046 (N_1046,In_432,In_1781);
and U1047 (N_1047,In_2188,In_311);
nand U1048 (N_1048,In_527,In_1347);
and U1049 (N_1049,In_1899,In_1742);
xor U1050 (N_1050,In_2763,In_2917);
nor U1051 (N_1051,In_967,In_1173);
and U1052 (N_1052,In_1510,In_1940);
nand U1053 (N_1053,In_719,In_2796);
nand U1054 (N_1054,In_1949,In_298);
or U1055 (N_1055,In_2264,In_831);
nand U1056 (N_1056,In_2172,In_1996);
nor U1057 (N_1057,In_1035,In_105);
xnor U1058 (N_1058,In_2627,In_1424);
nand U1059 (N_1059,In_2858,In_1275);
xnor U1060 (N_1060,In_2434,In_2475);
nor U1061 (N_1061,In_2511,In_2182);
nor U1062 (N_1062,In_1420,In_1252);
or U1063 (N_1063,In_1808,In_2562);
nand U1064 (N_1064,In_150,In_2463);
xor U1065 (N_1065,In_2764,In_1519);
or U1066 (N_1066,In_1455,In_1985);
xnor U1067 (N_1067,In_960,In_408);
and U1068 (N_1068,In_2085,In_2189);
nor U1069 (N_1069,In_2026,In_1555);
nand U1070 (N_1070,In_483,In_2570);
xnor U1071 (N_1071,In_124,In_2809);
or U1072 (N_1072,In_2020,In_1529);
or U1073 (N_1073,In_2667,In_2983);
xor U1074 (N_1074,In_2909,In_1118);
nand U1075 (N_1075,In_1988,In_780);
xor U1076 (N_1076,In_1998,In_1260);
nor U1077 (N_1077,In_1641,In_2056);
nand U1078 (N_1078,In_285,In_2753);
nor U1079 (N_1079,In_1225,In_1313);
xor U1080 (N_1080,In_2146,In_643);
nand U1081 (N_1081,In_1054,In_1771);
nand U1082 (N_1082,In_1654,In_2388);
xnor U1083 (N_1083,In_2981,In_1379);
xor U1084 (N_1084,In_173,In_887);
and U1085 (N_1085,In_1046,In_1268);
and U1086 (N_1086,In_1365,In_970);
nor U1087 (N_1087,In_1452,In_430);
xor U1088 (N_1088,In_1488,In_920);
nor U1089 (N_1089,In_2580,In_870);
nand U1090 (N_1090,In_662,In_2808);
xor U1091 (N_1091,In_2535,In_2);
xnor U1092 (N_1092,In_645,In_2704);
or U1093 (N_1093,In_1138,In_2919);
nand U1094 (N_1094,In_2051,In_903);
xor U1095 (N_1095,In_2997,In_2723);
or U1096 (N_1096,In_1289,In_1175);
or U1097 (N_1097,In_306,In_1619);
nand U1098 (N_1098,In_190,In_1719);
xor U1099 (N_1099,In_2116,In_470);
nor U1100 (N_1100,In_263,In_448);
and U1101 (N_1101,In_2495,In_2597);
and U1102 (N_1102,In_1033,In_1416);
xnor U1103 (N_1103,In_1766,In_1408);
nor U1104 (N_1104,In_550,In_262);
or U1105 (N_1105,In_1952,In_1950);
and U1106 (N_1106,In_147,In_2864);
xor U1107 (N_1107,In_2067,In_2399);
and U1108 (N_1108,In_2576,In_2226);
or U1109 (N_1109,In_971,In_2952);
and U1110 (N_1110,In_511,In_543);
nor U1111 (N_1111,In_487,In_1993);
xor U1112 (N_1112,In_177,In_791);
or U1113 (N_1113,In_1020,In_715);
and U1114 (N_1114,In_1358,In_2386);
nand U1115 (N_1115,In_1201,In_2221);
nor U1116 (N_1116,In_1068,In_2121);
nand U1117 (N_1117,In_1874,In_567);
and U1118 (N_1118,In_146,In_425);
nor U1119 (N_1119,In_179,In_1267);
nand U1120 (N_1120,In_898,In_768);
xnor U1121 (N_1121,In_1513,In_2081);
nor U1122 (N_1122,In_7,In_1036);
and U1123 (N_1123,In_2195,In_1708);
nor U1124 (N_1124,In_1656,In_1187);
xor U1125 (N_1125,In_2318,In_1902);
xor U1126 (N_1126,In_1962,In_1302);
xnor U1127 (N_1127,In_2725,In_1928);
and U1128 (N_1128,In_2623,In_468);
xnor U1129 (N_1129,In_2131,In_2681);
xnor U1130 (N_1130,In_77,In_2186);
nand U1131 (N_1131,In_1984,In_1927);
nand U1132 (N_1132,In_1056,In_2077);
nor U1133 (N_1133,In_1410,In_2312);
and U1134 (N_1134,In_2847,In_560);
xor U1135 (N_1135,In_641,In_2322);
and U1136 (N_1136,In_990,In_207);
xor U1137 (N_1137,In_2063,In_454);
or U1138 (N_1138,In_1841,In_671);
xnor U1139 (N_1139,In_1461,In_502);
nor U1140 (N_1140,In_91,In_2928);
nor U1141 (N_1141,In_2666,In_942);
xor U1142 (N_1142,In_1481,In_2709);
and U1143 (N_1143,In_546,In_994);
and U1144 (N_1144,In_406,In_1595);
or U1145 (N_1145,In_640,In_2833);
nand U1146 (N_1146,In_495,In_2357);
and U1147 (N_1147,In_579,In_258);
and U1148 (N_1148,In_1199,In_2458);
nand U1149 (N_1149,In_2883,In_2972);
nor U1150 (N_1150,In_789,In_1877);
nor U1151 (N_1151,In_2600,In_1018);
and U1152 (N_1152,In_2749,In_2218);
xor U1153 (N_1153,In_1875,In_321);
nand U1154 (N_1154,In_2546,In_1483);
xnor U1155 (N_1155,In_17,In_1121);
nor U1156 (N_1156,In_178,In_2382);
or U1157 (N_1157,In_2988,In_1005);
xor U1158 (N_1158,In_2424,In_675);
nand U1159 (N_1159,In_1397,In_837);
nand U1160 (N_1160,In_1543,In_565);
xor U1161 (N_1161,In_931,In_811);
and U1162 (N_1162,In_1243,In_2157);
and U1163 (N_1163,In_1215,In_414);
xor U1164 (N_1164,In_728,In_1077);
or U1165 (N_1165,In_2324,In_1607);
and U1166 (N_1166,In_192,In_2820);
nor U1167 (N_1167,In_1516,In_605);
xor U1168 (N_1168,In_267,In_2902);
nor U1169 (N_1169,In_604,In_198);
and U1170 (N_1170,In_1753,In_2824);
xnor U1171 (N_1171,In_2124,In_2998);
or U1172 (N_1172,In_472,In_955);
and U1173 (N_1173,In_2892,In_1373);
nand U1174 (N_1174,In_2560,In_1031);
or U1175 (N_1175,In_555,In_1300);
xor U1176 (N_1176,In_1017,In_2391);
xnor U1177 (N_1177,In_2078,In_65);
nand U1178 (N_1178,In_1528,In_582);
and U1179 (N_1179,In_2268,In_1847);
and U1180 (N_1180,In_665,In_2441);
or U1181 (N_1181,In_2676,In_1227);
xor U1182 (N_1182,In_435,In_547);
or U1183 (N_1183,In_443,In_907);
nand U1184 (N_1184,In_1295,In_1071);
and U1185 (N_1185,In_2164,In_2389);
or U1186 (N_1186,In_2448,In_623);
xor U1187 (N_1187,In_2904,In_1206);
nor U1188 (N_1188,In_123,In_1311);
or U1189 (N_1189,In_2110,In_620);
xnor U1190 (N_1190,In_1640,In_2481);
nor U1191 (N_1191,In_590,In_1345);
and U1192 (N_1192,In_1114,In_528);
nor U1193 (N_1193,In_2726,In_1645);
and U1194 (N_1194,In_2798,In_1324);
nand U1195 (N_1195,In_2482,In_2494);
xnor U1196 (N_1196,In_1584,In_1273);
nor U1197 (N_1197,In_1778,In_1075);
and U1198 (N_1198,In_1733,In_1058);
and U1199 (N_1199,In_978,In_302);
or U1200 (N_1200,In_1258,In_2117);
and U1201 (N_1201,In_574,In_2365);
and U1202 (N_1202,In_2999,In_2118);
nor U1203 (N_1203,In_433,In_653);
nor U1204 (N_1204,In_2873,In_1934);
and U1205 (N_1205,In_1383,In_2301);
nand U1206 (N_1206,In_2358,In_478);
and U1207 (N_1207,In_1971,In_2016);
and U1208 (N_1208,In_372,In_1966);
xnor U1209 (N_1209,In_2474,In_218);
or U1210 (N_1210,In_2814,In_2371);
and U1211 (N_1211,In_329,In_2392);
and U1212 (N_1212,In_720,In_176);
xor U1213 (N_1213,In_1831,In_1758);
or U1214 (N_1214,In_2520,In_1446);
xor U1215 (N_1215,In_2140,In_1592);
nor U1216 (N_1216,In_1739,In_554);
xnor U1217 (N_1217,In_852,In_1540);
and U1218 (N_1218,In_854,In_2669);
nor U1219 (N_1219,In_563,In_46);
nor U1220 (N_1220,In_27,In_2547);
and U1221 (N_1221,In_418,In_1897);
xnor U1222 (N_1222,In_2122,In_2050);
nand U1223 (N_1223,In_1181,In_2551);
and U1224 (N_1224,In_796,In_2974);
or U1225 (N_1225,In_890,In_2151);
xnor U1226 (N_1226,In_1438,In_869);
or U1227 (N_1227,In_2103,In_2907);
nor U1228 (N_1228,In_2037,In_2274);
or U1229 (N_1229,In_1332,In_1518);
and U1230 (N_1230,In_2220,In_1666);
or U1231 (N_1231,In_2834,In_2469);
nor U1232 (N_1232,In_1578,In_2948);
and U1233 (N_1233,In_1351,In_1282);
nand U1234 (N_1234,In_434,In_1449);
and U1235 (N_1235,In_505,In_2589);
nor U1236 (N_1236,In_2461,In_1819);
and U1237 (N_1237,In_2885,In_1210);
nand U1238 (N_1238,In_2423,In_136);
nand U1239 (N_1239,In_497,In_2470);
nor U1240 (N_1240,In_1886,In_1675);
or U1241 (N_1241,In_405,In_1638);
and U1242 (N_1242,In_1080,In_2417);
and U1243 (N_1243,In_1292,In_2432);
or U1244 (N_1244,In_2789,In_1890);
or U1245 (N_1245,In_2759,In_835);
nand U1246 (N_1246,In_1893,In_924);
or U1247 (N_1247,In_2224,In_2921);
nor U1248 (N_1248,In_2406,In_2890);
nand U1249 (N_1249,In_2253,In_184);
xnor U1250 (N_1250,In_2086,In_581);
or U1251 (N_1251,In_479,In_1929);
nor U1252 (N_1252,In_1714,In_1627);
nor U1253 (N_1253,In_2439,In_1933);
and U1254 (N_1254,In_1189,In_2139);
xnor U1255 (N_1255,In_2503,In_2072);
and U1256 (N_1256,In_2320,In_2690);
or U1257 (N_1257,In_1524,In_1721);
and U1258 (N_1258,In_2815,In_2048);
or U1259 (N_1259,In_1016,In_1823);
nand U1260 (N_1260,In_1969,In_1562);
nor U1261 (N_1261,In_1570,In_2523);
or U1262 (N_1262,In_2776,In_1860);
nor U1263 (N_1263,In_608,In_1843);
or U1264 (N_1264,In_714,In_2446);
and U1265 (N_1265,In_186,In_1476);
nand U1266 (N_1266,In_1975,In_1760);
nand U1267 (N_1267,In_2954,In_774);
nand U1268 (N_1268,In_750,In_2340);
nor U1269 (N_1269,In_301,In_410);
nand U1270 (N_1270,In_1283,In_36);
or U1271 (N_1271,In_2738,In_1414);
or U1272 (N_1272,In_1489,In_2817);
nand U1273 (N_1273,In_1631,In_2361);
nand U1274 (N_1274,In_1369,In_48);
nand U1275 (N_1275,In_153,In_403);
and U1276 (N_1276,In_1284,In_874);
and U1277 (N_1277,In_68,In_331);
or U1278 (N_1278,In_2515,In_1087);
and U1279 (N_1279,In_426,In_1898);
xor U1280 (N_1280,In_834,In_1346);
nand U1281 (N_1281,In_28,In_798);
nand U1282 (N_1282,In_1696,In_2011);
nand U1283 (N_1283,In_1015,In_1670);
and U1284 (N_1284,In_43,In_609);
or U1285 (N_1285,In_2178,In_2255);
nand U1286 (N_1286,In_156,In_1219);
xnor U1287 (N_1287,In_2457,In_187);
nor U1288 (N_1288,In_476,In_2316);
and U1289 (N_1289,In_446,In_112);
nor U1290 (N_1290,In_110,In_444);
nand U1291 (N_1291,In_1079,In_223);
and U1292 (N_1292,In_384,In_251);
nor U1293 (N_1293,In_855,In_1777);
xor U1294 (N_1294,In_142,In_1754);
xor U1295 (N_1295,In_1633,In_761);
nor U1296 (N_1296,In_607,In_910);
nand U1297 (N_1297,In_2012,In_362);
or U1298 (N_1298,In_888,In_2211);
nor U1299 (N_1299,In_305,In_2163);
xnor U1300 (N_1300,In_1428,In_1535);
or U1301 (N_1301,In_2635,In_2654);
nand U1302 (N_1302,In_2402,In_1871);
nand U1303 (N_1303,In_1393,In_836);
nor U1304 (N_1304,In_2867,In_1229);
nor U1305 (N_1305,In_788,In_2968);
xor U1306 (N_1306,In_1657,In_2650);
or U1307 (N_1307,In_2394,In_1343);
nand U1308 (N_1308,In_820,In_2571);
and U1309 (N_1309,In_2326,In_1158);
nand U1310 (N_1310,In_1278,In_1147);
nor U1311 (N_1311,In_457,In_195);
nor U1312 (N_1312,In_2497,In_1309);
xnor U1313 (N_1313,In_1915,In_1112);
nor U1314 (N_1314,In_1512,In_2830);
nand U1315 (N_1315,In_2028,In_1779);
and U1316 (N_1316,In_2415,In_1098);
or U1317 (N_1317,In_1662,In_2601);
or U1318 (N_1318,In_686,In_1554);
nand U1319 (N_1319,In_591,In_2231);
nor U1320 (N_1320,In_783,In_2664);
nor U1321 (N_1321,In_1280,In_1244);
xor U1322 (N_1322,In_952,In_1120);
and U1323 (N_1323,In_2230,In_449);
or U1324 (N_1324,In_40,In_2062);
xor U1325 (N_1325,In_2772,In_1149);
nand U1326 (N_1326,In_2805,In_669);
nand U1327 (N_1327,In_857,In_303);
xnor U1328 (N_1328,In_1593,In_2744);
or U1329 (N_1329,In_1867,In_2254);
nor U1330 (N_1330,In_1683,In_62);
and U1331 (N_1331,In_600,In_902);
nand U1332 (N_1332,In_1979,In_400);
nor U1333 (N_1333,In_2100,In_461);
and U1334 (N_1334,In_2542,In_1062);
nand U1335 (N_1335,In_463,In_2539);
nand U1336 (N_1336,In_1480,In_514);
nor U1337 (N_1337,In_2170,In_404);
xor U1338 (N_1338,In_2540,In_1228);
and U1339 (N_1339,In_1821,In_359);
xnor U1340 (N_1340,In_889,In_934);
nand U1341 (N_1341,In_1793,In_2410);
or U1342 (N_1342,In_749,In_982);
or U1343 (N_1343,In_757,In_2880);
nand U1344 (N_1344,In_1837,In_2861);
or U1345 (N_1345,In_2767,In_1135);
xor U1346 (N_1346,In_2807,In_940);
xnor U1347 (N_1347,In_1579,In_2091);
and U1348 (N_1348,In_1612,In_1074);
and U1349 (N_1349,In_2745,In_421);
xnor U1350 (N_1350,In_1911,In_1286);
and U1351 (N_1351,In_1029,In_1769);
nand U1352 (N_1352,In_1444,In_814);
or U1353 (N_1353,In_287,In_755);
nor U1354 (N_1354,In_2397,In_1813);
and U1355 (N_1355,In_1523,In_1262);
and U1356 (N_1356,In_657,In_415);
nor U1357 (N_1357,In_2479,In_1642);
xnor U1358 (N_1358,In_2647,In_352);
nand U1359 (N_1359,In_1868,In_734);
nor U1360 (N_1360,In_318,In_2874);
or U1361 (N_1361,In_2637,In_1912);
xor U1362 (N_1362,In_2823,In_1086);
nand U1363 (N_1363,In_635,In_1185);
nor U1364 (N_1364,In_2115,In_2616);
or U1365 (N_1365,In_492,In_666);
nor U1366 (N_1366,In_2362,In_1525);
and U1367 (N_1367,In_1063,In_2965);
and U1368 (N_1368,In_2526,In_2512);
or U1369 (N_1369,In_1816,In_1361);
or U1370 (N_1370,In_1213,In_589);
and U1371 (N_1371,In_570,In_642);
nor U1372 (N_1372,In_2927,In_390);
nand U1373 (N_1373,In_1076,In_498);
xor U1374 (N_1374,In_2758,In_597);
nand U1375 (N_1375,In_206,In_2692);
xor U1376 (N_1376,In_1829,In_1429);
or U1377 (N_1377,In_291,In_1143);
xor U1378 (N_1378,In_269,In_160);
nor U1379 (N_1379,In_1832,In_2329);
nor U1380 (N_1380,In_571,In_1827);
and U1381 (N_1381,In_165,In_706);
and U1382 (N_1382,In_897,In_1349);
or U1383 (N_1383,In_542,In_2941);
or U1384 (N_1384,In_1498,In_1241);
nand U1385 (N_1385,In_1501,In_2802);
xnor U1386 (N_1386,In_832,In_561);
or U1387 (N_1387,In_1217,In_1269);
nor U1388 (N_1388,In_762,In_2513);
nand U1389 (N_1389,In_1818,In_702);
nand U1390 (N_1390,In_2572,In_844);
or U1391 (N_1391,In_431,In_1731);
xor U1392 (N_1392,In_1287,In_2910);
xor U1393 (N_1393,In_1231,In_1256);
nand U1394 (N_1394,In_44,In_92);
and U1395 (N_1395,In_524,In_277);
nor U1396 (N_1396,In_82,In_1342);
xnor U1397 (N_1397,In_1573,In_2879);
and U1398 (N_1398,In_803,In_2577);
xor U1399 (N_1399,In_1168,In_915);
and U1400 (N_1400,In_2022,In_1249);
nand U1401 (N_1401,In_1460,In_2501);
nand U1402 (N_1402,In_32,In_1807);
nor U1403 (N_1403,In_1650,In_523);
and U1404 (N_1404,In_1146,In_658);
nand U1405 (N_1405,In_1021,In_369);
nor U1406 (N_1406,In_2148,In_1132);
nand U1407 (N_1407,In_2945,In_900);
xor U1408 (N_1408,In_1532,In_2351);
and U1409 (N_1409,In_1840,In_956);
nor U1410 (N_1410,In_2018,In_2612);
and U1411 (N_1411,In_114,In_2114);
nand U1412 (N_1412,In_2489,In_1522);
nand U1413 (N_1413,In_1380,In_751);
nor U1414 (N_1414,In_925,In_1870);
or U1415 (N_1415,In_911,In_336);
xnor U1416 (N_1416,In_943,In_354);
xor U1417 (N_1417,In_861,In_1712);
xor U1418 (N_1418,In_2257,In_1456);
and U1419 (N_1419,In_2428,In_300);
nand U1420 (N_1420,In_1496,In_475);
nand U1421 (N_1421,In_1568,In_13);
or U1422 (N_1422,In_1963,In_941);
and U1423 (N_1423,In_564,In_2591);
nand U1424 (N_1424,In_718,In_2414);
and U1425 (N_1425,In_2256,In_864);
and U1426 (N_1426,In_848,In_2138);
xnor U1427 (N_1427,In_963,In_2702);
xor U1428 (N_1428,In_1172,In_840);
and U1429 (N_1429,In_1101,In_696);
nand U1430 (N_1430,In_1621,In_2295);
nor U1431 (N_1431,In_1328,In_1824);
nor U1432 (N_1432,In_138,In_2087);
nor U1433 (N_1433,In_66,In_531);
nor U1434 (N_1434,In_2027,In_2135);
nand U1435 (N_1435,In_1756,In_945);
nor U1436 (N_1436,In_41,In_1925);
xor U1437 (N_1437,In_1233,In_1861);
nor U1438 (N_1438,In_2377,In_2359);
nor U1439 (N_1439,In_1938,In_2659);
and U1440 (N_1440,In_2689,In_697);
nor U1441 (N_1441,In_6,In_2004);
xor U1442 (N_1442,In_2437,In_343);
and U1443 (N_1443,In_2827,In_2401);
xnor U1444 (N_1444,In_1637,In_987);
or U1445 (N_1445,In_1789,In_1051);
or U1446 (N_1446,In_2854,In_572);
nand U1447 (N_1447,In_2396,In_2710);
xnor U1448 (N_1448,In_394,In_323);
nand U1449 (N_1449,In_1407,In_727);
nor U1450 (N_1450,In_2047,In_2206);
nor U1451 (N_1451,In_2728,In_1557);
nor U1452 (N_1452,In_97,In_1334);
xor U1453 (N_1453,In_917,In_2840);
and U1454 (N_1454,In_137,In_754);
nor U1455 (N_1455,In_2915,In_2920);
nand U1456 (N_1456,In_163,In_1333);
and U1457 (N_1457,In_452,In_1359);
or U1458 (N_1458,In_810,In_1520);
nor U1459 (N_1459,In_1646,In_1626);
xnor U1460 (N_1460,In_2393,In_396);
nor U1461 (N_1461,In_2651,In_1008);
nand U1462 (N_1462,In_985,In_2125);
nand U1463 (N_1463,In_2177,In_76);
or U1464 (N_1464,In_242,In_1632);
nand U1465 (N_1465,In_2522,In_2822);
xor U1466 (N_1466,In_1155,In_2425);
and U1467 (N_1467,In_2942,In_2958);
and U1468 (N_1468,In_2793,In_1916);
xnor U1469 (N_1469,In_1140,In_1943);
xnor U1470 (N_1470,In_2471,In_1830);
and U1471 (N_1471,In_2713,In_2721);
or U1472 (N_1472,In_2630,In_230);
or U1473 (N_1473,In_210,In_886);
nor U1474 (N_1474,In_2618,In_94);
or U1475 (N_1475,In_759,In_1500);
nor U1476 (N_1476,In_785,In_1858);
and U1477 (N_1477,In_2130,In_1085);
nor U1478 (N_1478,In_14,In_1478);
nor U1479 (N_1479,In_1576,In_1341);
xor U1480 (N_1480,In_292,In_1002);
nor U1481 (N_1481,In_977,In_2557);
or U1482 (N_1482,In_1312,In_1468);
or U1483 (N_1483,In_1503,In_1127);
nor U1484 (N_1484,In_2123,In_1010);
nand U1485 (N_1485,In_2762,In_1798);
nor U1486 (N_1486,In_1603,In_833);
or U1487 (N_1487,In_1003,In_2550);
xor U1488 (N_1488,In_1092,In_801);
nor U1489 (N_1489,In_1774,In_337);
and U1490 (N_1490,In_368,In_851);
or U1491 (N_1491,In_217,In_231);
nand U1492 (N_1492,In_308,In_1119);
nand U1493 (N_1493,In_2868,In_1968);
or U1494 (N_1494,In_1125,In_145);
and U1495 (N_1495,In_2336,In_2477);
and U1496 (N_1496,In_741,In_573);
xnor U1497 (N_1497,In_989,In_843);
and U1498 (N_1498,In_1257,In_2747);
or U1499 (N_1499,In_1291,In_1375);
and U1500 (N_1500,In_1201,In_682);
xnor U1501 (N_1501,In_2402,In_2365);
nand U1502 (N_1502,In_428,In_1026);
and U1503 (N_1503,In_1832,In_1434);
and U1504 (N_1504,In_310,In_651);
and U1505 (N_1505,In_873,In_977);
xnor U1506 (N_1506,In_1139,In_223);
xnor U1507 (N_1507,In_1944,In_1910);
nand U1508 (N_1508,In_1133,In_643);
nand U1509 (N_1509,In_1391,In_1591);
nor U1510 (N_1510,In_2224,In_239);
and U1511 (N_1511,In_169,In_1993);
and U1512 (N_1512,In_2183,In_2854);
nor U1513 (N_1513,In_728,In_2115);
xor U1514 (N_1514,In_2888,In_1023);
nor U1515 (N_1515,In_446,In_2724);
nor U1516 (N_1516,In_1252,In_728);
xor U1517 (N_1517,In_413,In_2876);
xor U1518 (N_1518,In_2184,In_838);
xor U1519 (N_1519,In_2013,In_579);
or U1520 (N_1520,In_1380,In_2512);
or U1521 (N_1521,In_1757,In_2958);
nand U1522 (N_1522,In_212,In_750);
or U1523 (N_1523,In_2026,In_2727);
nand U1524 (N_1524,In_2705,In_1184);
nand U1525 (N_1525,In_220,In_1620);
nor U1526 (N_1526,In_2260,In_784);
xnor U1527 (N_1527,In_801,In_892);
nand U1528 (N_1528,In_545,In_38);
nor U1529 (N_1529,In_254,In_1254);
xnor U1530 (N_1530,In_917,In_2204);
or U1531 (N_1531,In_2647,In_2085);
nand U1532 (N_1532,In_223,In_949);
or U1533 (N_1533,In_1099,In_599);
or U1534 (N_1534,In_2327,In_2906);
xor U1535 (N_1535,In_1153,In_1736);
xnor U1536 (N_1536,In_2505,In_91);
nand U1537 (N_1537,In_1917,In_1916);
or U1538 (N_1538,In_882,In_424);
nor U1539 (N_1539,In_565,In_1765);
xor U1540 (N_1540,In_405,In_2066);
nand U1541 (N_1541,In_456,In_14);
or U1542 (N_1542,In_1931,In_1181);
xor U1543 (N_1543,In_209,In_1644);
or U1544 (N_1544,In_1512,In_1087);
and U1545 (N_1545,In_1778,In_2110);
nor U1546 (N_1546,In_1547,In_2155);
nor U1547 (N_1547,In_470,In_427);
or U1548 (N_1548,In_1434,In_1516);
and U1549 (N_1549,In_273,In_360);
and U1550 (N_1550,In_1954,In_2566);
xor U1551 (N_1551,In_1669,In_389);
nor U1552 (N_1552,In_1869,In_52);
and U1553 (N_1553,In_2418,In_524);
nand U1554 (N_1554,In_18,In_1753);
nand U1555 (N_1555,In_2995,In_1527);
or U1556 (N_1556,In_287,In_2967);
or U1557 (N_1557,In_1874,In_470);
or U1558 (N_1558,In_406,In_1235);
or U1559 (N_1559,In_2435,In_2411);
and U1560 (N_1560,In_907,In_2813);
nand U1561 (N_1561,In_2837,In_960);
and U1562 (N_1562,In_1192,In_727);
nand U1563 (N_1563,In_2346,In_2397);
nor U1564 (N_1564,In_2275,In_2934);
or U1565 (N_1565,In_1302,In_112);
xnor U1566 (N_1566,In_259,In_2346);
nor U1567 (N_1567,In_414,In_2945);
xnor U1568 (N_1568,In_2764,In_2661);
xor U1569 (N_1569,In_2940,In_1640);
nand U1570 (N_1570,In_887,In_2714);
nand U1571 (N_1571,In_1803,In_2277);
and U1572 (N_1572,In_126,In_750);
xnor U1573 (N_1573,In_2953,In_337);
xor U1574 (N_1574,In_1314,In_1270);
nand U1575 (N_1575,In_249,In_901);
or U1576 (N_1576,In_1626,In_1245);
or U1577 (N_1577,In_925,In_368);
xnor U1578 (N_1578,In_1655,In_374);
and U1579 (N_1579,In_2381,In_1759);
and U1580 (N_1580,In_1917,In_1940);
or U1581 (N_1581,In_1701,In_1140);
nor U1582 (N_1582,In_1835,In_595);
xor U1583 (N_1583,In_1766,In_163);
nor U1584 (N_1584,In_143,In_1054);
nor U1585 (N_1585,In_2441,In_1505);
xnor U1586 (N_1586,In_2868,In_1112);
nand U1587 (N_1587,In_1900,In_2003);
nand U1588 (N_1588,In_1775,In_2881);
and U1589 (N_1589,In_2206,In_1070);
nor U1590 (N_1590,In_2203,In_1505);
or U1591 (N_1591,In_2384,In_714);
nor U1592 (N_1592,In_1075,In_1090);
nand U1593 (N_1593,In_249,In_594);
xnor U1594 (N_1594,In_2262,In_2945);
xor U1595 (N_1595,In_1382,In_2142);
and U1596 (N_1596,In_428,In_1244);
or U1597 (N_1597,In_1983,In_348);
and U1598 (N_1598,In_2387,In_409);
or U1599 (N_1599,In_487,In_651);
nand U1600 (N_1600,In_467,In_267);
or U1601 (N_1601,In_1063,In_2562);
xnor U1602 (N_1602,In_1777,In_1381);
and U1603 (N_1603,In_1790,In_2912);
or U1604 (N_1604,In_2143,In_2947);
xnor U1605 (N_1605,In_1823,In_314);
nand U1606 (N_1606,In_1989,In_69);
xor U1607 (N_1607,In_533,In_1702);
and U1608 (N_1608,In_613,In_2664);
or U1609 (N_1609,In_1729,In_2981);
xor U1610 (N_1610,In_1126,In_871);
and U1611 (N_1611,In_1881,In_117);
xor U1612 (N_1612,In_1591,In_1404);
nand U1613 (N_1613,In_1987,In_2726);
xor U1614 (N_1614,In_395,In_2425);
nand U1615 (N_1615,In_1151,In_2916);
nor U1616 (N_1616,In_294,In_1705);
and U1617 (N_1617,In_182,In_2987);
or U1618 (N_1618,In_721,In_1177);
nand U1619 (N_1619,In_222,In_572);
nand U1620 (N_1620,In_1269,In_2462);
or U1621 (N_1621,In_87,In_1259);
or U1622 (N_1622,In_2057,In_1090);
or U1623 (N_1623,In_436,In_590);
nor U1624 (N_1624,In_2476,In_628);
xnor U1625 (N_1625,In_1725,In_135);
nor U1626 (N_1626,In_2687,In_295);
nand U1627 (N_1627,In_1621,In_2796);
nor U1628 (N_1628,In_770,In_2469);
nand U1629 (N_1629,In_461,In_1071);
and U1630 (N_1630,In_1809,In_2466);
nand U1631 (N_1631,In_542,In_506);
xnor U1632 (N_1632,In_135,In_576);
xor U1633 (N_1633,In_898,In_1999);
and U1634 (N_1634,In_2877,In_498);
or U1635 (N_1635,In_1093,In_1687);
nor U1636 (N_1636,In_2537,In_229);
and U1637 (N_1637,In_2662,In_2590);
xnor U1638 (N_1638,In_826,In_2463);
and U1639 (N_1639,In_2523,In_947);
or U1640 (N_1640,In_2517,In_2980);
nand U1641 (N_1641,In_180,In_2688);
nor U1642 (N_1642,In_227,In_2501);
or U1643 (N_1643,In_2902,In_2818);
nand U1644 (N_1644,In_679,In_1951);
nand U1645 (N_1645,In_2635,In_2904);
xor U1646 (N_1646,In_409,In_1699);
and U1647 (N_1647,In_704,In_2556);
xnor U1648 (N_1648,In_2370,In_1329);
xor U1649 (N_1649,In_254,In_1982);
xnor U1650 (N_1650,In_1898,In_2238);
and U1651 (N_1651,In_115,In_177);
xor U1652 (N_1652,In_1932,In_2190);
xor U1653 (N_1653,In_1294,In_38);
nor U1654 (N_1654,In_2103,In_2270);
nor U1655 (N_1655,In_178,In_2589);
xor U1656 (N_1656,In_617,In_581);
xnor U1657 (N_1657,In_554,In_429);
and U1658 (N_1658,In_523,In_1598);
nand U1659 (N_1659,In_1064,In_644);
xor U1660 (N_1660,In_1141,In_2121);
and U1661 (N_1661,In_1908,In_2871);
nor U1662 (N_1662,In_1367,In_677);
or U1663 (N_1663,In_593,In_595);
nand U1664 (N_1664,In_2458,In_1876);
xor U1665 (N_1665,In_2302,In_880);
or U1666 (N_1666,In_1501,In_1836);
nor U1667 (N_1667,In_882,In_937);
xnor U1668 (N_1668,In_2791,In_895);
nand U1669 (N_1669,In_1265,In_2465);
or U1670 (N_1670,In_592,In_2207);
or U1671 (N_1671,In_804,In_882);
and U1672 (N_1672,In_1197,In_1232);
or U1673 (N_1673,In_482,In_2297);
nor U1674 (N_1674,In_1809,In_151);
or U1675 (N_1675,In_1058,In_1991);
or U1676 (N_1676,In_2371,In_1629);
nand U1677 (N_1677,In_1702,In_1409);
and U1678 (N_1678,In_92,In_485);
or U1679 (N_1679,In_1347,In_2373);
and U1680 (N_1680,In_483,In_2907);
or U1681 (N_1681,In_528,In_2968);
nand U1682 (N_1682,In_92,In_1461);
xnor U1683 (N_1683,In_1095,In_2816);
nand U1684 (N_1684,In_448,In_906);
and U1685 (N_1685,In_2191,In_1438);
or U1686 (N_1686,In_2405,In_321);
or U1687 (N_1687,In_487,In_1172);
or U1688 (N_1688,In_2887,In_1408);
nand U1689 (N_1689,In_1369,In_987);
xor U1690 (N_1690,In_2437,In_1114);
xor U1691 (N_1691,In_2653,In_871);
or U1692 (N_1692,In_1255,In_2346);
xor U1693 (N_1693,In_2516,In_1775);
xor U1694 (N_1694,In_123,In_337);
xor U1695 (N_1695,In_221,In_2459);
and U1696 (N_1696,In_15,In_536);
nor U1697 (N_1697,In_1536,In_1270);
nor U1698 (N_1698,In_909,In_1385);
or U1699 (N_1699,In_676,In_589);
or U1700 (N_1700,In_258,In_1758);
and U1701 (N_1701,In_1940,In_1657);
xnor U1702 (N_1702,In_2830,In_2574);
nor U1703 (N_1703,In_2016,In_1730);
nor U1704 (N_1704,In_1210,In_2391);
or U1705 (N_1705,In_1472,In_125);
or U1706 (N_1706,In_204,In_1694);
nand U1707 (N_1707,In_435,In_1607);
and U1708 (N_1708,In_2489,In_509);
or U1709 (N_1709,In_2891,In_415);
nor U1710 (N_1710,In_1126,In_2144);
nor U1711 (N_1711,In_1104,In_1772);
and U1712 (N_1712,In_764,In_1780);
nor U1713 (N_1713,In_2278,In_554);
nor U1714 (N_1714,In_530,In_1091);
xnor U1715 (N_1715,In_2987,In_1935);
nand U1716 (N_1716,In_1951,In_1026);
xor U1717 (N_1717,In_932,In_929);
xor U1718 (N_1718,In_1532,In_2300);
xor U1719 (N_1719,In_1218,In_2731);
xor U1720 (N_1720,In_2403,In_2269);
xnor U1721 (N_1721,In_1535,In_1925);
and U1722 (N_1722,In_990,In_2171);
xnor U1723 (N_1723,In_338,In_895);
xnor U1724 (N_1724,In_680,In_1845);
xor U1725 (N_1725,In_2799,In_2965);
xnor U1726 (N_1726,In_2638,In_2603);
nand U1727 (N_1727,In_856,In_2904);
nand U1728 (N_1728,In_401,In_2278);
and U1729 (N_1729,In_107,In_67);
and U1730 (N_1730,In_2622,In_2721);
nor U1731 (N_1731,In_1244,In_717);
nand U1732 (N_1732,In_1114,In_2041);
xor U1733 (N_1733,In_888,In_2227);
and U1734 (N_1734,In_926,In_2463);
xor U1735 (N_1735,In_733,In_1018);
or U1736 (N_1736,In_2659,In_1114);
and U1737 (N_1737,In_2456,In_1472);
nor U1738 (N_1738,In_961,In_2619);
nand U1739 (N_1739,In_1948,In_1825);
or U1740 (N_1740,In_90,In_2730);
or U1741 (N_1741,In_2464,In_293);
xnor U1742 (N_1742,In_2294,In_1210);
or U1743 (N_1743,In_1681,In_1981);
and U1744 (N_1744,In_966,In_1221);
nand U1745 (N_1745,In_2900,In_930);
nand U1746 (N_1746,In_1373,In_1492);
and U1747 (N_1747,In_539,In_1749);
or U1748 (N_1748,In_2387,In_1816);
and U1749 (N_1749,In_964,In_1136);
nor U1750 (N_1750,In_1665,In_76);
and U1751 (N_1751,In_1634,In_1622);
or U1752 (N_1752,In_1428,In_1898);
or U1753 (N_1753,In_2206,In_1610);
nor U1754 (N_1754,In_2929,In_190);
nor U1755 (N_1755,In_963,In_1607);
or U1756 (N_1756,In_2046,In_958);
nand U1757 (N_1757,In_367,In_1226);
nor U1758 (N_1758,In_852,In_37);
and U1759 (N_1759,In_1284,In_2259);
nand U1760 (N_1760,In_2269,In_2721);
nor U1761 (N_1761,In_2035,In_2765);
nor U1762 (N_1762,In_1966,In_2677);
xor U1763 (N_1763,In_1262,In_1473);
nor U1764 (N_1764,In_2405,In_1780);
xnor U1765 (N_1765,In_2609,In_2505);
or U1766 (N_1766,In_2980,In_1125);
xnor U1767 (N_1767,In_2747,In_335);
nand U1768 (N_1768,In_1548,In_62);
and U1769 (N_1769,In_100,In_2575);
or U1770 (N_1770,In_1755,In_496);
and U1771 (N_1771,In_2853,In_1734);
and U1772 (N_1772,In_310,In_1787);
xnor U1773 (N_1773,In_883,In_2321);
and U1774 (N_1774,In_590,In_2656);
xnor U1775 (N_1775,In_1826,In_1436);
nand U1776 (N_1776,In_2647,In_958);
and U1777 (N_1777,In_2379,In_6);
nand U1778 (N_1778,In_438,In_655);
nor U1779 (N_1779,In_1048,In_2956);
xnor U1780 (N_1780,In_1693,In_1101);
nor U1781 (N_1781,In_1748,In_595);
xnor U1782 (N_1782,In_30,In_1521);
nand U1783 (N_1783,In_2850,In_1253);
or U1784 (N_1784,In_2841,In_375);
nor U1785 (N_1785,In_2647,In_2861);
nor U1786 (N_1786,In_2966,In_988);
xor U1787 (N_1787,In_1846,In_829);
or U1788 (N_1788,In_1060,In_2970);
and U1789 (N_1789,In_1454,In_666);
nand U1790 (N_1790,In_1191,In_966);
nand U1791 (N_1791,In_1928,In_685);
and U1792 (N_1792,In_1653,In_2812);
and U1793 (N_1793,In_2195,In_1973);
or U1794 (N_1794,In_2145,In_2309);
nand U1795 (N_1795,In_2673,In_1912);
and U1796 (N_1796,In_2795,In_1046);
or U1797 (N_1797,In_2929,In_2711);
or U1798 (N_1798,In_2675,In_2305);
xor U1799 (N_1799,In_1587,In_973);
nor U1800 (N_1800,In_1839,In_1072);
and U1801 (N_1801,In_2516,In_1627);
and U1802 (N_1802,In_1000,In_2166);
or U1803 (N_1803,In_693,In_431);
nor U1804 (N_1804,In_1732,In_2417);
xnor U1805 (N_1805,In_134,In_2196);
nor U1806 (N_1806,In_163,In_679);
xor U1807 (N_1807,In_533,In_1371);
nor U1808 (N_1808,In_1278,In_1396);
or U1809 (N_1809,In_2218,In_77);
nand U1810 (N_1810,In_1790,In_2951);
xnor U1811 (N_1811,In_1374,In_814);
nor U1812 (N_1812,In_1085,In_2805);
or U1813 (N_1813,In_2316,In_2157);
or U1814 (N_1814,In_2439,In_38);
or U1815 (N_1815,In_182,In_638);
xnor U1816 (N_1816,In_538,In_2834);
nand U1817 (N_1817,In_1686,In_2118);
nand U1818 (N_1818,In_2737,In_1787);
or U1819 (N_1819,In_2104,In_218);
nand U1820 (N_1820,In_180,In_1306);
xnor U1821 (N_1821,In_2984,In_2730);
and U1822 (N_1822,In_1873,In_2965);
xor U1823 (N_1823,In_1090,In_2213);
or U1824 (N_1824,In_2942,In_1432);
xor U1825 (N_1825,In_2240,In_2833);
and U1826 (N_1826,In_233,In_86);
nand U1827 (N_1827,In_2251,In_2721);
nand U1828 (N_1828,In_20,In_1035);
or U1829 (N_1829,In_2135,In_1200);
xnor U1830 (N_1830,In_1117,In_2024);
and U1831 (N_1831,In_1275,In_1691);
nor U1832 (N_1832,In_788,In_804);
nor U1833 (N_1833,In_2123,In_2708);
and U1834 (N_1834,In_1904,In_2880);
nor U1835 (N_1835,In_104,In_639);
nor U1836 (N_1836,In_607,In_2719);
xor U1837 (N_1837,In_767,In_2526);
nor U1838 (N_1838,In_1057,In_1417);
xnor U1839 (N_1839,In_935,In_121);
and U1840 (N_1840,In_1482,In_2080);
and U1841 (N_1841,In_1262,In_2560);
xor U1842 (N_1842,In_1855,In_1039);
xor U1843 (N_1843,In_660,In_1044);
nand U1844 (N_1844,In_1906,In_871);
xnor U1845 (N_1845,In_2722,In_1503);
and U1846 (N_1846,In_638,In_497);
xor U1847 (N_1847,In_1158,In_137);
and U1848 (N_1848,In_1273,In_526);
xnor U1849 (N_1849,In_137,In_2302);
xnor U1850 (N_1850,In_2905,In_2168);
or U1851 (N_1851,In_1773,In_406);
and U1852 (N_1852,In_1813,In_1226);
xnor U1853 (N_1853,In_2460,In_2243);
xor U1854 (N_1854,In_2734,In_314);
xor U1855 (N_1855,In_2019,In_1747);
xor U1856 (N_1856,In_1541,In_1184);
or U1857 (N_1857,In_549,In_1749);
nand U1858 (N_1858,In_1442,In_1441);
xor U1859 (N_1859,In_948,In_525);
nand U1860 (N_1860,In_429,In_334);
or U1861 (N_1861,In_1188,In_2956);
and U1862 (N_1862,In_2072,In_2693);
nand U1863 (N_1863,In_372,In_2121);
or U1864 (N_1864,In_2591,In_772);
nor U1865 (N_1865,In_2302,In_1372);
or U1866 (N_1866,In_2497,In_1115);
nor U1867 (N_1867,In_271,In_1374);
and U1868 (N_1868,In_1436,In_2074);
nand U1869 (N_1869,In_315,In_2688);
and U1870 (N_1870,In_2785,In_1712);
nand U1871 (N_1871,In_454,In_1708);
nor U1872 (N_1872,In_955,In_412);
or U1873 (N_1873,In_1829,In_540);
nand U1874 (N_1874,In_1938,In_2997);
xor U1875 (N_1875,In_1553,In_1006);
nor U1876 (N_1876,In_51,In_1540);
or U1877 (N_1877,In_2822,In_307);
and U1878 (N_1878,In_2526,In_1626);
xnor U1879 (N_1879,In_1243,In_1793);
xor U1880 (N_1880,In_1049,In_2423);
and U1881 (N_1881,In_459,In_1266);
nand U1882 (N_1882,In_2872,In_2808);
or U1883 (N_1883,In_1007,In_2489);
nand U1884 (N_1884,In_2652,In_1093);
xor U1885 (N_1885,In_1687,In_2197);
and U1886 (N_1886,In_138,In_363);
or U1887 (N_1887,In_2227,In_2295);
and U1888 (N_1888,In_1972,In_1525);
xnor U1889 (N_1889,In_259,In_562);
nand U1890 (N_1890,In_1755,In_2670);
nor U1891 (N_1891,In_954,In_554);
xnor U1892 (N_1892,In_1416,In_561);
or U1893 (N_1893,In_1253,In_2493);
nor U1894 (N_1894,In_2475,In_1481);
nor U1895 (N_1895,In_1958,In_438);
nand U1896 (N_1896,In_598,In_810);
nand U1897 (N_1897,In_2713,In_1197);
or U1898 (N_1898,In_2406,In_574);
or U1899 (N_1899,In_1007,In_67);
xnor U1900 (N_1900,In_758,In_1533);
nand U1901 (N_1901,In_1338,In_2454);
xnor U1902 (N_1902,In_2502,In_2984);
nand U1903 (N_1903,In_146,In_1920);
and U1904 (N_1904,In_2670,In_2984);
or U1905 (N_1905,In_2525,In_999);
nand U1906 (N_1906,In_453,In_2302);
and U1907 (N_1907,In_222,In_1268);
or U1908 (N_1908,In_2933,In_90);
nand U1909 (N_1909,In_303,In_1483);
nor U1910 (N_1910,In_951,In_2773);
and U1911 (N_1911,In_1136,In_707);
and U1912 (N_1912,In_2235,In_2076);
nand U1913 (N_1913,In_2104,In_2950);
or U1914 (N_1914,In_2497,In_303);
nand U1915 (N_1915,In_1535,In_829);
and U1916 (N_1916,In_1589,In_278);
or U1917 (N_1917,In_1688,In_1777);
or U1918 (N_1918,In_114,In_1209);
nor U1919 (N_1919,In_1560,In_2098);
xnor U1920 (N_1920,In_1844,In_964);
nand U1921 (N_1921,In_2071,In_2143);
nor U1922 (N_1922,In_1625,In_893);
xor U1923 (N_1923,In_2645,In_867);
xor U1924 (N_1924,In_1643,In_1000);
or U1925 (N_1925,In_1565,In_1429);
nand U1926 (N_1926,In_2092,In_88);
nand U1927 (N_1927,In_2339,In_2624);
nor U1928 (N_1928,In_350,In_809);
and U1929 (N_1929,In_469,In_1427);
xnor U1930 (N_1930,In_904,In_1213);
nor U1931 (N_1931,In_817,In_1941);
nor U1932 (N_1932,In_2008,In_1120);
xor U1933 (N_1933,In_2158,In_2295);
nand U1934 (N_1934,In_2513,In_2090);
nor U1935 (N_1935,In_2194,In_9);
nand U1936 (N_1936,In_1942,In_1060);
nor U1937 (N_1937,In_2072,In_2190);
and U1938 (N_1938,In_2481,In_2613);
and U1939 (N_1939,In_645,In_1643);
nor U1940 (N_1940,In_1667,In_2529);
nand U1941 (N_1941,In_301,In_1495);
or U1942 (N_1942,In_884,In_416);
or U1943 (N_1943,In_900,In_290);
nand U1944 (N_1944,In_1888,In_2050);
xnor U1945 (N_1945,In_1672,In_1977);
xnor U1946 (N_1946,In_2210,In_2930);
nand U1947 (N_1947,In_506,In_2508);
nand U1948 (N_1948,In_8,In_481);
xor U1949 (N_1949,In_1094,In_1677);
nor U1950 (N_1950,In_2030,In_2768);
xor U1951 (N_1951,In_2423,In_2750);
or U1952 (N_1952,In_2138,In_1442);
and U1953 (N_1953,In_2289,In_1227);
nand U1954 (N_1954,In_1019,In_1343);
nor U1955 (N_1955,In_2944,In_2331);
nor U1956 (N_1956,In_155,In_798);
and U1957 (N_1957,In_1108,In_2010);
or U1958 (N_1958,In_1809,In_1602);
nor U1959 (N_1959,In_2139,In_647);
or U1960 (N_1960,In_2887,In_276);
and U1961 (N_1961,In_1672,In_2775);
nor U1962 (N_1962,In_2902,In_2132);
and U1963 (N_1963,In_2498,In_1069);
nor U1964 (N_1964,In_460,In_2046);
xnor U1965 (N_1965,In_2955,In_840);
xnor U1966 (N_1966,In_2600,In_4);
nand U1967 (N_1967,In_37,In_1675);
or U1968 (N_1968,In_2332,In_2121);
and U1969 (N_1969,In_444,In_1213);
nor U1970 (N_1970,In_2008,In_811);
xor U1971 (N_1971,In_1487,In_1763);
or U1972 (N_1972,In_476,In_2922);
or U1973 (N_1973,In_50,In_1489);
and U1974 (N_1974,In_2174,In_2494);
nor U1975 (N_1975,In_266,In_2023);
or U1976 (N_1976,In_1476,In_1434);
xnor U1977 (N_1977,In_2998,In_1465);
nor U1978 (N_1978,In_2558,In_808);
xor U1979 (N_1979,In_1335,In_740);
xor U1980 (N_1980,In_619,In_751);
and U1981 (N_1981,In_1403,In_598);
or U1982 (N_1982,In_660,In_1060);
xor U1983 (N_1983,In_2956,In_2541);
nor U1984 (N_1984,In_2602,In_963);
xnor U1985 (N_1985,In_869,In_1967);
nand U1986 (N_1986,In_828,In_75);
nor U1987 (N_1987,In_1462,In_221);
nand U1988 (N_1988,In_1511,In_636);
xnor U1989 (N_1989,In_665,In_47);
or U1990 (N_1990,In_2737,In_1298);
or U1991 (N_1991,In_1292,In_631);
xnor U1992 (N_1992,In_631,In_751);
nor U1993 (N_1993,In_1975,In_2545);
and U1994 (N_1994,In_435,In_2273);
and U1995 (N_1995,In_879,In_2859);
xnor U1996 (N_1996,In_1979,In_1481);
nand U1997 (N_1997,In_649,In_973);
xnor U1998 (N_1998,In_500,In_176);
or U1999 (N_1999,In_2941,In_801);
nor U2000 (N_2000,In_2140,In_1186);
nor U2001 (N_2001,In_429,In_2961);
or U2002 (N_2002,In_2240,In_1723);
nand U2003 (N_2003,In_1959,In_2380);
nand U2004 (N_2004,In_557,In_1531);
xor U2005 (N_2005,In_255,In_2124);
or U2006 (N_2006,In_2459,In_224);
or U2007 (N_2007,In_1983,In_1096);
nand U2008 (N_2008,In_1292,In_1752);
or U2009 (N_2009,In_1604,In_704);
nor U2010 (N_2010,In_2281,In_1913);
xnor U2011 (N_2011,In_1014,In_1402);
nor U2012 (N_2012,In_1889,In_1980);
nand U2013 (N_2013,In_1441,In_2071);
xor U2014 (N_2014,In_2979,In_1998);
nand U2015 (N_2015,In_485,In_1256);
nor U2016 (N_2016,In_2158,In_565);
and U2017 (N_2017,In_1656,In_1016);
nor U2018 (N_2018,In_1143,In_2453);
or U2019 (N_2019,In_2425,In_1446);
nor U2020 (N_2020,In_2874,In_2164);
and U2021 (N_2021,In_2095,In_640);
and U2022 (N_2022,In_2076,In_2179);
and U2023 (N_2023,In_2138,In_2694);
or U2024 (N_2024,In_878,In_163);
and U2025 (N_2025,In_1750,In_2183);
nor U2026 (N_2026,In_920,In_545);
and U2027 (N_2027,In_1367,In_2112);
or U2028 (N_2028,In_1019,In_416);
or U2029 (N_2029,In_2422,In_1272);
and U2030 (N_2030,In_1206,In_2649);
and U2031 (N_2031,In_2317,In_2712);
xor U2032 (N_2032,In_2042,In_2100);
and U2033 (N_2033,In_732,In_933);
and U2034 (N_2034,In_847,In_1078);
nand U2035 (N_2035,In_490,In_1055);
nor U2036 (N_2036,In_2819,In_441);
nand U2037 (N_2037,In_2304,In_457);
and U2038 (N_2038,In_3,In_1811);
and U2039 (N_2039,In_2168,In_45);
nand U2040 (N_2040,In_1061,In_2182);
and U2041 (N_2041,In_1809,In_2616);
nor U2042 (N_2042,In_697,In_1794);
and U2043 (N_2043,In_1467,In_2371);
nor U2044 (N_2044,In_179,In_348);
xor U2045 (N_2045,In_1298,In_5);
nor U2046 (N_2046,In_2386,In_1473);
and U2047 (N_2047,In_1440,In_1307);
nor U2048 (N_2048,In_758,In_2740);
nand U2049 (N_2049,In_2391,In_2038);
or U2050 (N_2050,In_865,In_2992);
nor U2051 (N_2051,In_2373,In_2385);
or U2052 (N_2052,In_74,In_2665);
xnor U2053 (N_2053,In_1272,In_2124);
xor U2054 (N_2054,In_199,In_1461);
or U2055 (N_2055,In_1794,In_1732);
or U2056 (N_2056,In_1689,In_2156);
xnor U2057 (N_2057,In_2810,In_2764);
or U2058 (N_2058,In_300,In_2993);
and U2059 (N_2059,In_2261,In_240);
or U2060 (N_2060,In_1810,In_891);
and U2061 (N_2061,In_1413,In_1096);
nor U2062 (N_2062,In_77,In_2814);
nor U2063 (N_2063,In_1044,In_2257);
nor U2064 (N_2064,In_1056,In_2521);
nand U2065 (N_2065,In_1830,In_1311);
nor U2066 (N_2066,In_2797,In_1718);
and U2067 (N_2067,In_81,In_1593);
or U2068 (N_2068,In_2949,In_2271);
xor U2069 (N_2069,In_1297,In_2870);
or U2070 (N_2070,In_243,In_574);
xnor U2071 (N_2071,In_1695,In_2602);
xor U2072 (N_2072,In_167,In_113);
and U2073 (N_2073,In_1280,In_1666);
and U2074 (N_2074,In_1567,In_1795);
nand U2075 (N_2075,In_2290,In_1423);
xor U2076 (N_2076,In_2143,In_1490);
xor U2077 (N_2077,In_321,In_1836);
nor U2078 (N_2078,In_1009,In_784);
xnor U2079 (N_2079,In_2767,In_2584);
nand U2080 (N_2080,In_2894,In_2491);
and U2081 (N_2081,In_1192,In_196);
or U2082 (N_2082,In_2150,In_627);
nor U2083 (N_2083,In_1364,In_2104);
or U2084 (N_2084,In_399,In_2324);
or U2085 (N_2085,In_2527,In_907);
nand U2086 (N_2086,In_642,In_1010);
nand U2087 (N_2087,In_1806,In_84);
nor U2088 (N_2088,In_2959,In_528);
nor U2089 (N_2089,In_1912,In_1625);
and U2090 (N_2090,In_1729,In_1987);
nand U2091 (N_2091,In_1671,In_2097);
nand U2092 (N_2092,In_1447,In_2945);
or U2093 (N_2093,In_2500,In_1711);
and U2094 (N_2094,In_2017,In_2132);
nand U2095 (N_2095,In_100,In_242);
xor U2096 (N_2096,In_2720,In_978);
or U2097 (N_2097,In_1046,In_1160);
nor U2098 (N_2098,In_525,In_2057);
or U2099 (N_2099,In_1756,In_542);
nand U2100 (N_2100,In_636,In_322);
or U2101 (N_2101,In_763,In_2403);
or U2102 (N_2102,In_558,In_248);
or U2103 (N_2103,In_869,In_807);
and U2104 (N_2104,In_2760,In_2716);
nor U2105 (N_2105,In_2386,In_2470);
or U2106 (N_2106,In_2976,In_2212);
xor U2107 (N_2107,In_2943,In_2937);
nor U2108 (N_2108,In_2653,In_1657);
and U2109 (N_2109,In_2793,In_702);
nor U2110 (N_2110,In_157,In_1320);
and U2111 (N_2111,In_1743,In_1598);
and U2112 (N_2112,In_1735,In_1527);
or U2113 (N_2113,In_1110,In_69);
and U2114 (N_2114,In_813,In_2082);
or U2115 (N_2115,In_403,In_2385);
and U2116 (N_2116,In_1626,In_156);
nand U2117 (N_2117,In_930,In_1102);
and U2118 (N_2118,In_2694,In_1063);
xnor U2119 (N_2119,In_2484,In_2812);
nor U2120 (N_2120,In_2087,In_2935);
and U2121 (N_2121,In_2969,In_2731);
xor U2122 (N_2122,In_2030,In_910);
nand U2123 (N_2123,In_620,In_2388);
xor U2124 (N_2124,In_745,In_1484);
xnor U2125 (N_2125,In_595,In_482);
or U2126 (N_2126,In_995,In_2303);
xor U2127 (N_2127,In_511,In_137);
and U2128 (N_2128,In_72,In_933);
xnor U2129 (N_2129,In_2652,In_2302);
xnor U2130 (N_2130,In_2086,In_1415);
xor U2131 (N_2131,In_315,In_854);
or U2132 (N_2132,In_2970,In_2163);
xor U2133 (N_2133,In_20,In_962);
nor U2134 (N_2134,In_1618,In_292);
and U2135 (N_2135,In_256,In_1521);
nor U2136 (N_2136,In_2229,In_1035);
nor U2137 (N_2137,In_751,In_2789);
or U2138 (N_2138,In_615,In_579);
or U2139 (N_2139,In_929,In_2208);
xnor U2140 (N_2140,In_1076,In_2860);
or U2141 (N_2141,In_659,In_1623);
nor U2142 (N_2142,In_69,In_725);
and U2143 (N_2143,In_172,In_569);
or U2144 (N_2144,In_1015,In_1689);
or U2145 (N_2145,In_2817,In_793);
nor U2146 (N_2146,In_2732,In_2589);
xnor U2147 (N_2147,In_799,In_1220);
and U2148 (N_2148,In_839,In_391);
or U2149 (N_2149,In_2756,In_2228);
nand U2150 (N_2150,In_1225,In_1956);
nor U2151 (N_2151,In_506,In_628);
xor U2152 (N_2152,In_2192,In_1657);
xor U2153 (N_2153,In_2854,In_2436);
and U2154 (N_2154,In_1727,In_960);
xor U2155 (N_2155,In_641,In_2305);
nor U2156 (N_2156,In_2957,In_406);
nor U2157 (N_2157,In_298,In_1160);
nor U2158 (N_2158,In_2481,In_482);
or U2159 (N_2159,In_1975,In_2886);
nand U2160 (N_2160,In_1492,In_2153);
nand U2161 (N_2161,In_665,In_767);
nand U2162 (N_2162,In_843,In_2729);
xor U2163 (N_2163,In_1580,In_1505);
or U2164 (N_2164,In_1382,In_1670);
and U2165 (N_2165,In_186,In_2658);
and U2166 (N_2166,In_2107,In_2044);
or U2167 (N_2167,In_762,In_2080);
nand U2168 (N_2168,In_1009,In_1367);
nand U2169 (N_2169,In_1318,In_2111);
and U2170 (N_2170,In_1831,In_1328);
nand U2171 (N_2171,In_22,In_2104);
and U2172 (N_2172,In_1938,In_2513);
xnor U2173 (N_2173,In_484,In_2937);
nor U2174 (N_2174,In_2331,In_2138);
and U2175 (N_2175,In_1863,In_571);
and U2176 (N_2176,In_1103,In_2643);
nand U2177 (N_2177,In_2925,In_742);
nor U2178 (N_2178,In_2751,In_534);
or U2179 (N_2179,In_1289,In_2933);
nor U2180 (N_2180,In_668,In_2503);
nand U2181 (N_2181,In_539,In_1866);
nand U2182 (N_2182,In_2565,In_2382);
or U2183 (N_2183,In_2569,In_1163);
xor U2184 (N_2184,In_244,In_687);
xnor U2185 (N_2185,In_189,In_203);
nand U2186 (N_2186,In_1473,In_2020);
nor U2187 (N_2187,In_1741,In_1111);
nand U2188 (N_2188,In_551,In_1621);
nor U2189 (N_2189,In_2387,In_1657);
nand U2190 (N_2190,In_1799,In_408);
nor U2191 (N_2191,In_2904,In_403);
or U2192 (N_2192,In_1634,In_1256);
nor U2193 (N_2193,In_1776,In_196);
and U2194 (N_2194,In_828,In_2458);
and U2195 (N_2195,In_1563,In_1567);
and U2196 (N_2196,In_1973,In_449);
nand U2197 (N_2197,In_2368,In_1367);
nand U2198 (N_2198,In_114,In_943);
or U2199 (N_2199,In_1253,In_2475);
or U2200 (N_2200,In_1266,In_244);
or U2201 (N_2201,In_1958,In_2414);
nand U2202 (N_2202,In_2788,In_2327);
and U2203 (N_2203,In_2695,In_2336);
and U2204 (N_2204,In_270,In_166);
xor U2205 (N_2205,In_79,In_507);
and U2206 (N_2206,In_224,In_2981);
nand U2207 (N_2207,In_2295,In_2528);
and U2208 (N_2208,In_1450,In_1227);
nand U2209 (N_2209,In_2617,In_2833);
or U2210 (N_2210,In_556,In_2804);
nand U2211 (N_2211,In_58,In_2211);
or U2212 (N_2212,In_1683,In_2194);
nor U2213 (N_2213,In_749,In_77);
nand U2214 (N_2214,In_942,In_2901);
or U2215 (N_2215,In_2602,In_2877);
nor U2216 (N_2216,In_1604,In_1431);
nand U2217 (N_2217,In_949,In_568);
nor U2218 (N_2218,In_252,In_437);
and U2219 (N_2219,In_2416,In_571);
and U2220 (N_2220,In_330,In_705);
nand U2221 (N_2221,In_596,In_1821);
or U2222 (N_2222,In_793,In_1011);
xnor U2223 (N_2223,In_965,In_450);
nor U2224 (N_2224,In_624,In_40);
nand U2225 (N_2225,In_189,In_790);
or U2226 (N_2226,In_2984,In_2976);
nor U2227 (N_2227,In_1817,In_976);
nand U2228 (N_2228,In_295,In_1354);
nand U2229 (N_2229,In_1966,In_2965);
nand U2230 (N_2230,In_595,In_1945);
and U2231 (N_2231,In_232,In_154);
and U2232 (N_2232,In_113,In_2688);
and U2233 (N_2233,In_1784,In_2414);
nor U2234 (N_2234,In_777,In_900);
and U2235 (N_2235,In_1027,In_1137);
and U2236 (N_2236,In_2281,In_2861);
nor U2237 (N_2237,In_2687,In_1642);
nor U2238 (N_2238,In_2709,In_926);
and U2239 (N_2239,In_389,In_1475);
or U2240 (N_2240,In_321,In_2544);
and U2241 (N_2241,In_2513,In_2651);
nor U2242 (N_2242,In_397,In_653);
nor U2243 (N_2243,In_1369,In_2821);
nand U2244 (N_2244,In_2455,In_1554);
nand U2245 (N_2245,In_340,In_2298);
or U2246 (N_2246,In_1109,In_779);
and U2247 (N_2247,In_335,In_2697);
nor U2248 (N_2248,In_657,In_2767);
and U2249 (N_2249,In_1272,In_352);
and U2250 (N_2250,In_1113,In_1799);
nor U2251 (N_2251,In_982,In_586);
nor U2252 (N_2252,In_854,In_2499);
xnor U2253 (N_2253,In_2970,In_1518);
nor U2254 (N_2254,In_1021,In_1786);
xnor U2255 (N_2255,In_1590,In_1076);
xor U2256 (N_2256,In_1175,In_804);
xnor U2257 (N_2257,In_1549,In_829);
nand U2258 (N_2258,In_2543,In_707);
xnor U2259 (N_2259,In_2119,In_2820);
nand U2260 (N_2260,In_1752,In_1596);
and U2261 (N_2261,In_35,In_932);
or U2262 (N_2262,In_2159,In_2294);
xnor U2263 (N_2263,In_1091,In_819);
or U2264 (N_2264,In_2396,In_1135);
nand U2265 (N_2265,In_68,In_1067);
and U2266 (N_2266,In_643,In_219);
nand U2267 (N_2267,In_1292,In_2813);
xnor U2268 (N_2268,In_1044,In_1485);
nor U2269 (N_2269,In_2212,In_1364);
nor U2270 (N_2270,In_1432,In_796);
xor U2271 (N_2271,In_1621,In_553);
nor U2272 (N_2272,In_2412,In_145);
xnor U2273 (N_2273,In_2795,In_1343);
nor U2274 (N_2274,In_2558,In_1182);
nand U2275 (N_2275,In_2863,In_2363);
nand U2276 (N_2276,In_1579,In_1265);
and U2277 (N_2277,In_1098,In_2444);
nand U2278 (N_2278,In_1060,In_956);
or U2279 (N_2279,In_461,In_800);
and U2280 (N_2280,In_844,In_819);
nor U2281 (N_2281,In_1639,In_1864);
xor U2282 (N_2282,In_1372,In_1671);
and U2283 (N_2283,In_660,In_1921);
nor U2284 (N_2284,In_826,In_454);
and U2285 (N_2285,In_1230,In_873);
and U2286 (N_2286,In_1628,In_2209);
xnor U2287 (N_2287,In_2325,In_265);
and U2288 (N_2288,In_2715,In_2070);
xnor U2289 (N_2289,In_2595,In_1749);
xnor U2290 (N_2290,In_2674,In_2568);
xor U2291 (N_2291,In_1038,In_1911);
nor U2292 (N_2292,In_2031,In_1404);
nor U2293 (N_2293,In_2596,In_92);
nor U2294 (N_2294,In_991,In_2014);
or U2295 (N_2295,In_331,In_2384);
or U2296 (N_2296,In_943,In_456);
nor U2297 (N_2297,In_292,In_460);
and U2298 (N_2298,In_926,In_951);
nand U2299 (N_2299,In_2381,In_237);
and U2300 (N_2300,In_2349,In_2487);
or U2301 (N_2301,In_1823,In_2384);
or U2302 (N_2302,In_879,In_869);
xnor U2303 (N_2303,In_2756,In_2314);
and U2304 (N_2304,In_212,In_2743);
nand U2305 (N_2305,In_2761,In_1385);
nor U2306 (N_2306,In_2986,In_749);
nor U2307 (N_2307,In_2304,In_488);
and U2308 (N_2308,In_1045,In_81);
nand U2309 (N_2309,In_2933,In_1698);
nor U2310 (N_2310,In_1716,In_651);
and U2311 (N_2311,In_1073,In_2308);
and U2312 (N_2312,In_1857,In_2070);
nor U2313 (N_2313,In_672,In_2977);
nand U2314 (N_2314,In_1040,In_1574);
or U2315 (N_2315,In_1533,In_334);
xnor U2316 (N_2316,In_1437,In_2803);
nand U2317 (N_2317,In_2390,In_2472);
and U2318 (N_2318,In_960,In_1348);
nand U2319 (N_2319,In_440,In_2334);
nor U2320 (N_2320,In_1683,In_548);
or U2321 (N_2321,In_614,In_2738);
nand U2322 (N_2322,In_1675,In_1477);
xor U2323 (N_2323,In_133,In_1158);
xor U2324 (N_2324,In_2944,In_701);
and U2325 (N_2325,In_2585,In_2820);
nand U2326 (N_2326,In_2858,In_2022);
xor U2327 (N_2327,In_2554,In_1363);
xor U2328 (N_2328,In_1954,In_176);
or U2329 (N_2329,In_2450,In_2885);
or U2330 (N_2330,In_2920,In_1794);
and U2331 (N_2331,In_1909,In_1872);
nand U2332 (N_2332,In_2194,In_1164);
nor U2333 (N_2333,In_2267,In_1481);
or U2334 (N_2334,In_1141,In_2145);
and U2335 (N_2335,In_2050,In_2065);
xnor U2336 (N_2336,In_160,In_2129);
xnor U2337 (N_2337,In_256,In_2502);
nand U2338 (N_2338,In_2037,In_1112);
or U2339 (N_2339,In_181,In_1449);
nor U2340 (N_2340,In_736,In_560);
and U2341 (N_2341,In_2786,In_435);
or U2342 (N_2342,In_408,In_2642);
nor U2343 (N_2343,In_249,In_2446);
nand U2344 (N_2344,In_1023,In_1501);
and U2345 (N_2345,In_2889,In_1586);
or U2346 (N_2346,In_2370,In_2068);
nor U2347 (N_2347,In_303,In_726);
and U2348 (N_2348,In_1156,In_1682);
or U2349 (N_2349,In_1663,In_815);
nor U2350 (N_2350,In_2188,In_322);
or U2351 (N_2351,In_1588,In_2519);
or U2352 (N_2352,In_1776,In_1421);
nor U2353 (N_2353,In_2379,In_1266);
nor U2354 (N_2354,In_2349,In_2055);
and U2355 (N_2355,In_2075,In_801);
and U2356 (N_2356,In_1833,In_2836);
nor U2357 (N_2357,In_464,In_73);
nand U2358 (N_2358,In_2689,In_906);
nor U2359 (N_2359,In_2414,In_2573);
xor U2360 (N_2360,In_2806,In_1541);
xor U2361 (N_2361,In_1086,In_1675);
or U2362 (N_2362,In_1601,In_1110);
nor U2363 (N_2363,In_268,In_184);
xnor U2364 (N_2364,In_700,In_36);
nor U2365 (N_2365,In_656,In_947);
xor U2366 (N_2366,In_646,In_2986);
xor U2367 (N_2367,In_1307,In_1837);
nor U2368 (N_2368,In_608,In_474);
and U2369 (N_2369,In_2480,In_1146);
or U2370 (N_2370,In_1035,In_576);
nor U2371 (N_2371,In_1857,In_1485);
and U2372 (N_2372,In_1375,In_1155);
nand U2373 (N_2373,In_2186,In_299);
or U2374 (N_2374,In_2867,In_2484);
nor U2375 (N_2375,In_976,In_2082);
xnor U2376 (N_2376,In_901,In_2576);
or U2377 (N_2377,In_766,In_1698);
xnor U2378 (N_2378,In_1974,In_2816);
xor U2379 (N_2379,In_2040,In_1646);
xnor U2380 (N_2380,In_2463,In_2694);
or U2381 (N_2381,In_67,In_2488);
nand U2382 (N_2382,In_1271,In_1276);
xnor U2383 (N_2383,In_1786,In_1498);
xor U2384 (N_2384,In_2937,In_2183);
or U2385 (N_2385,In_2464,In_2918);
and U2386 (N_2386,In_975,In_1256);
nand U2387 (N_2387,In_1447,In_641);
nor U2388 (N_2388,In_420,In_2808);
xnor U2389 (N_2389,In_2824,In_1412);
and U2390 (N_2390,In_2089,In_2919);
nor U2391 (N_2391,In_863,In_1823);
and U2392 (N_2392,In_350,In_2578);
xor U2393 (N_2393,In_1685,In_1635);
or U2394 (N_2394,In_1139,In_2639);
nor U2395 (N_2395,In_1962,In_900);
or U2396 (N_2396,In_1856,In_662);
nand U2397 (N_2397,In_1830,In_2872);
and U2398 (N_2398,In_929,In_115);
or U2399 (N_2399,In_1350,In_2277);
nor U2400 (N_2400,In_2261,In_2620);
nor U2401 (N_2401,In_2341,In_1672);
nor U2402 (N_2402,In_2650,In_1438);
xor U2403 (N_2403,In_715,In_2372);
nor U2404 (N_2404,In_326,In_822);
nor U2405 (N_2405,In_290,In_2702);
xor U2406 (N_2406,In_1168,In_2905);
or U2407 (N_2407,In_1743,In_1003);
or U2408 (N_2408,In_1255,In_712);
nand U2409 (N_2409,In_469,In_1175);
nand U2410 (N_2410,In_2435,In_1731);
xnor U2411 (N_2411,In_1823,In_625);
nor U2412 (N_2412,In_2898,In_2239);
xor U2413 (N_2413,In_1890,In_870);
and U2414 (N_2414,In_740,In_1083);
and U2415 (N_2415,In_2672,In_1687);
nand U2416 (N_2416,In_2528,In_103);
and U2417 (N_2417,In_786,In_2762);
or U2418 (N_2418,In_854,In_2253);
and U2419 (N_2419,In_977,In_2839);
or U2420 (N_2420,In_2815,In_859);
nand U2421 (N_2421,In_1107,In_477);
nand U2422 (N_2422,In_1569,In_521);
xor U2423 (N_2423,In_1938,In_840);
and U2424 (N_2424,In_1639,In_2333);
xnor U2425 (N_2425,In_1263,In_1941);
and U2426 (N_2426,In_1567,In_599);
nor U2427 (N_2427,In_34,In_1363);
and U2428 (N_2428,In_102,In_1184);
nor U2429 (N_2429,In_1747,In_2368);
or U2430 (N_2430,In_1130,In_2865);
xnor U2431 (N_2431,In_96,In_1865);
and U2432 (N_2432,In_2943,In_1381);
and U2433 (N_2433,In_1774,In_913);
nand U2434 (N_2434,In_1359,In_1279);
and U2435 (N_2435,In_2989,In_1389);
xor U2436 (N_2436,In_479,In_1717);
nand U2437 (N_2437,In_1233,In_1812);
nor U2438 (N_2438,In_1025,In_236);
nor U2439 (N_2439,In_726,In_1062);
xor U2440 (N_2440,In_748,In_1169);
or U2441 (N_2441,In_83,In_1802);
and U2442 (N_2442,In_2584,In_2404);
and U2443 (N_2443,In_2428,In_1145);
nand U2444 (N_2444,In_2211,In_215);
xor U2445 (N_2445,In_1982,In_1650);
nor U2446 (N_2446,In_1641,In_354);
xor U2447 (N_2447,In_491,In_597);
nand U2448 (N_2448,In_1360,In_879);
or U2449 (N_2449,In_779,In_417);
nor U2450 (N_2450,In_518,In_2447);
xor U2451 (N_2451,In_136,In_1310);
nand U2452 (N_2452,In_1426,In_1323);
and U2453 (N_2453,In_1828,In_279);
or U2454 (N_2454,In_2690,In_2856);
xnor U2455 (N_2455,In_1247,In_2731);
xor U2456 (N_2456,In_1885,In_324);
and U2457 (N_2457,In_246,In_1452);
nor U2458 (N_2458,In_1259,In_510);
or U2459 (N_2459,In_2961,In_1388);
xnor U2460 (N_2460,In_1042,In_730);
and U2461 (N_2461,In_706,In_160);
xnor U2462 (N_2462,In_2530,In_1162);
nor U2463 (N_2463,In_1850,In_1463);
or U2464 (N_2464,In_232,In_2296);
and U2465 (N_2465,In_675,In_2486);
nand U2466 (N_2466,In_1354,In_578);
or U2467 (N_2467,In_311,In_1265);
xnor U2468 (N_2468,In_2519,In_2246);
nor U2469 (N_2469,In_29,In_1309);
or U2470 (N_2470,In_969,In_342);
nand U2471 (N_2471,In_1801,In_1860);
nand U2472 (N_2472,In_2087,In_733);
and U2473 (N_2473,In_2188,In_105);
nand U2474 (N_2474,In_1731,In_2421);
and U2475 (N_2475,In_1432,In_2071);
and U2476 (N_2476,In_1564,In_478);
nor U2477 (N_2477,In_680,In_2606);
or U2478 (N_2478,In_1182,In_171);
and U2479 (N_2479,In_667,In_1745);
nor U2480 (N_2480,In_1345,In_2742);
xnor U2481 (N_2481,In_2461,In_1635);
nand U2482 (N_2482,In_390,In_407);
and U2483 (N_2483,In_784,In_816);
nor U2484 (N_2484,In_270,In_176);
nand U2485 (N_2485,In_2809,In_701);
xor U2486 (N_2486,In_2191,In_498);
nor U2487 (N_2487,In_2606,In_583);
and U2488 (N_2488,In_2836,In_1116);
or U2489 (N_2489,In_231,In_1426);
and U2490 (N_2490,In_1357,In_379);
nand U2491 (N_2491,In_543,In_1189);
nand U2492 (N_2492,In_1837,In_1862);
xnor U2493 (N_2493,In_2937,In_1669);
and U2494 (N_2494,In_640,In_1359);
or U2495 (N_2495,In_1044,In_1046);
and U2496 (N_2496,In_524,In_2883);
and U2497 (N_2497,In_988,In_2473);
or U2498 (N_2498,In_725,In_2995);
nand U2499 (N_2499,In_613,In_1792);
and U2500 (N_2500,In_2018,In_1512);
and U2501 (N_2501,In_1975,In_1252);
and U2502 (N_2502,In_2035,In_2271);
nand U2503 (N_2503,In_2021,In_203);
or U2504 (N_2504,In_2058,In_1185);
xnor U2505 (N_2505,In_2217,In_2366);
nor U2506 (N_2506,In_2506,In_1032);
nor U2507 (N_2507,In_2945,In_1661);
xor U2508 (N_2508,In_818,In_671);
xor U2509 (N_2509,In_2025,In_37);
and U2510 (N_2510,In_2933,In_15);
or U2511 (N_2511,In_1764,In_2811);
and U2512 (N_2512,In_163,In_46);
and U2513 (N_2513,In_1445,In_2012);
and U2514 (N_2514,In_292,In_1945);
xor U2515 (N_2515,In_1490,In_2426);
and U2516 (N_2516,In_2121,In_1993);
xor U2517 (N_2517,In_1469,In_2632);
or U2518 (N_2518,In_2269,In_2456);
or U2519 (N_2519,In_1917,In_1759);
and U2520 (N_2520,In_1524,In_1066);
nand U2521 (N_2521,In_39,In_2140);
or U2522 (N_2522,In_259,In_855);
or U2523 (N_2523,In_90,In_1362);
or U2524 (N_2524,In_1073,In_2110);
and U2525 (N_2525,In_1523,In_2006);
and U2526 (N_2526,In_65,In_168);
or U2527 (N_2527,In_1530,In_323);
and U2528 (N_2528,In_1447,In_1924);
nor U2529 (N_2529,In_2898,In_814);
or U2530 (N_2530,In_809,In_2351);
or U2531 (N_2531,In_2848,In_614);
and U2532 (N_2532,In_1848,In_1089);
xor U2533 (N_2533,In_2928,In_1188);
nand U2534 (N_2534,In_1698,In_2303);
and U2535 (N_2535,In_747,In_377);
xnor U2536 (N_2536,In_581,In_544);
and U2537 (N_2537,In_1238,In_1342);
xnor U2538 (N_2538,In_877,In_852);
and U2539 (N_2539,In_35,In_2198);
and U2540 (N_2540,In_628,In_287);
nor U2541 (N_2541,In_1303,In_2978);
or U2542 (N_2542,In_1352,In_1079);
nand U2543 (N_2543,In_1523,In_1953);
nor U2544 (N_2544,In_2304,In_1030);
or U2545 (N_2545,In_2553,In_599);
and U2546 (N_2546,In_1274,In_2133);
xnor U2547 (N_2547,In_1469,In_2008);
nor U2548 (N_2548,In_242,In_346);
or U2549 (N_2549,In_2404,In_1724);
nand U2550 (N_2550,In_1982,In_1634);
or U2551 (N_2551,In_1742,In_1297);
nor U2552 (N_2552,In_2226,In_1648);
nor U2553 (N_2553,In_2025,In_2463);
nor U2554 (N_2554,In_55,In_984);
and U2555 (N_2555,In_2145,In_1351);
nand U2556 (N_2556,In_399,In_1976);
nand U2557 (N_2557,In_1221,In_1953);
or U2558 (N_2558,In_267,In_2549);
and U2559 (N_2559,In_2215,In_1451);
and U2560 (N_2560,In_2123,In_1129);
xnor U2561 (N_2561,In_1434,In_1548);
xor U2562 (N_2562,In_2339,In_2457);
and U2563 (N_2563,In_603,In_2197);
nand U2564 (N_2564,In_2254,In_385);
nand U2565 (N_2565,In_2400,In_1473);
nor U2566 (N_2566,In_1151,In_1829);
and U2567 (N_2567,In_1525,In_556);
or U2568 (N_2568,In_2552,In_1713);
xor U2569 (N_2569,In_1323,In_916);
or U2570 (N_2570,In_1982,In_2872);
and U2571 (N_2571,In_355,In_2253);
nor U2572 (N_2572,In_1557,In_1801);
xor U2573 (N_2573,In_2252,In_1880);
nor U2574 (N_2574,In_1798,In_124);
nor U2575 (N_2575,In_1624,In_2963);
nand U2576 (N_2576,In_2913,In_2136);
nand U2577 (N_2577,In_1795,In_1860);
nand U2578 (N_2578,In_685,In_472);
nor U2579 (N_2579,In_1603,In_2337);
xor U2580 (N_2580,In_2812,In_790);
xor U2581 (N_2581,In_2445,In_1482);
xnor U2582 (N_2582,In_722,In_2988);
and U2583 (N_2583,In_492,In_1287);
and U2584 (N_2584,In_1538,In_2682);
xnor U2585 (N_2585,In_1975,In_1634);
and U2586 (N_2586,In_77,In_1321);
and U2587 (N_2587,In_1243,In_492);
nor U2588 (N_2588,In_2056,In_1612);
xor U2589 (N_2589,In_884,In_2573);
nand U2590 (N_2590,In_294,In_319);
and U2591 (N_2591,In_15,In_2142);
xor U2592 (N_2592,In_1156,In_2135);
and U2593 (N_2593,In_85,In_866);
or U2594 (N_2594,In_121,In_1858);
nand U2595 (N_2595,In_1262,In_347);
nand U2596 (N_2596,In_2693,In_890);
nor U2597 (N_2597,In_1593,In_2593);
and U2598 (N_2598,In_24,In_486);
xor U2599 (N_2599,In_1769,In_2188);
xnor U2600 (N_2600,In_2163,In_1467);
or U2601 (N_2601,In_1397,In_72);
nor U2602 (N_2602,In_311,In_2035);
xor U2603 (N_2603,In_2614,In_2695);
xnor U2604 (N_2604,In_1081,In_713);
nor U2605 (N_2605,In_1226,In_831);
and U2606 (N_2606,In_376,In_1991);
or U2607 (N_2607,In_2023,In_2525);
xor U2608 (N_2608,In_486,In_2019);
or U2609 (N_2609,In_415,In_2546);
or U2610 (N_2610,In_897,In_401);
nor U2611 (N_2611,In_2267,In_1151);
or U2612 (N_2612,In_2285,In_2079);
nand U2613 (N_2613,In_404,In_949);
nor U2614 (N_2614,In_1583,In_669);
nor U2615 (N_2615,In_993,In_896);
xor U2616 (N_2616,In_403,In_1319);
nor U2617 (N_2617,In_1019,In_2789);
nor U2618 (N_2618,In_1038,In_76);
or U2619 (N_2619,In_1762,In_2003);
xor U2620 (N_2620,In_2776,In_797);
nor U2621 (N_2621,In_1488,In_2296);
and U2622 (N_2622,In_289,In_583);
or U2623 (N_2623,In_2228,In_1458);
nand U2624 (N_2624,In_1727,In_2256);
or U2625 (N_2625,In_2301,In_707);
nand U2626 (N_2626,In_1482,In_1969);
or U2627 (N_2627,In_1190,In_904);
nor U2628 (N_2628,In_1474,In_1339);
or U2629 (N_2629,In_329,In_1843);
and U2630 (N_2630,In_1452,In_1381);
xor U2631 (N_2631,In_2239,In_1245);
and U2632 (N_2632,In_489,In_1557);
nand U2633 (N_2633,In_332,In_1536);
nand U2634 (N_2634,In_2817,In_2083);
and U2635 (N_2635,In_2305,In_45);
nand U2636 (N_2636,In_1023,In_2896);
nor U2637 (N_2637,In_1059,In_1883);
xnor U2638 (N_2638,In_782,In_1021);
or U2639 (N_2639,In_581,In_942);
or U2640 (N_2640,In_1783,In_407);
nand U2641 (N_2641,In_1245,In_309);
xnor U2642 (N_2642,In_340,In_1345);
xnor U2643 (N_2643,In_2695,In_159);
nor U2644 (N_2644,In_2290,In_831);
nor U2645 (N_2645,In_2102,In_1997);
and U2646 (N_2646,In_730,In_2940);
and U2647 (N_2647,In_1416,In_1512);
nor U2648 (N_2648,In_1350,In_372);
or U2649 (N_2649,In_588,In_1025);
nand U2650 (N_2650,In_2123,In_2603);
nand U2651 (N_2651,In_1222,In_99);
and U2652 (N_2652,In_338,In_765);
nand U2653 (N_2653,In_2644,In_469);
xnor U2654 (N_2654,In_1513,In_1622);
xor U2655 (N_2655,In_2814,In_2806);
xnor U2656 (N_2656,In_230,In_2752);
or U2657 (N_2657,In_258,In_2876);
nor U2658 (N_2658,In_2441,In_2209);
and U2659 (N_2659,In_1254,In_326);
and U2660 (N_2660,In_1816,In_1434);
nor U2661 (N_2661,In_1895,In_1321);
xnor U2662 (N_2662,In_2545,In_2767);
and U2663 (N_2663,In_1750,In_2643);
or U2664 (N_2664,In_571,In_2523);
xnor U2665 (N_2665,In_1674,In_2410);
and U2666 (N_2666,In_2435,In_1501);
and U2667 (N_2667,In_1364,In_2022);
and U2668 (N_2668,In_982,In_1377);
xnor U2669 (N_2669,In_695,In_2412);
nand U2670 (N_2670,In_1129,In_2853);
and U2671 (N_2671,In_2039,In_2495);
and U2672 (N_2672,In_310,In_2553);
xnor U2673 (N_2673,In_2176,In_550);
nand U2674 (N_2674,In_2544,In_575);
and U2675 (N_2675,In_2815,In_2401);
xnor U2676 (N_2676,In_325,In_308);
or U2677 (N_2677,In_2748,In_1023);
nand U2678 (N_2678,In_2495,In_1914);
nand U2679 (N_2679,In_542,In_2319);
and U2680 (N_2680,In_412,In_190);
nand U2681 (N_2681,In_607,In_2798);
xor U2682 (N_2682,In_661,In_1771);
nor U2683 (N_2683,In_2507,In_2406);
xor U2684 (N_2684,In_1833,In_154);
nand U2685 (N_2685,In_2773,In_265);
nor U2686 (N_2686,In_2395,In_979);
and U2687 (N_2687,In_1059,In_2924);
nor U2688 (N_2688,In_576,In_1861);
xnor U2689 (N_2689,In_2320,In_2479);
xnor U2690 (N_2690,In_2408,In_2591);
nor U2691 (N_2691,In_800,In_776);
xor U2692 (N_2692,In_992,In_2706);
nor U2693 (N_2693,In_2082,In_1601);
nand U2694 (N_2694,In_1867,In_1540);
xor U2695 (N_2695,In_2861,In_1810);
xor U2696 (N_2696,In_426,In_1737);
xor U2697 (N_2697,In_1724,In_1914);
nor U2698 (N_2698,In_963,In_2454);
and U2699 (N_2699,In_2184,In_850);
nor U2700 (N_2700,In_1073,In_428);
nor U2701 (N_2701,In_2542,In_2773);
or U2702 (N_2702,In_1791,In_1417);
or U2703 (N_2703,In_535,In_471);
and U2704 (N_2704,In_2392,In_321);
xor U2705 (N_2705,In_2045,In_871);
and U2706 (N_2706,In_613,In_1632);
xnor U2707 (N_2707,In_2026,In_2125);
nor U2708 (N_2708,In_641,In_347);
nor U2709 (N_2709,In_1105,In_314);
and U2710 (N_2710,In_1922,In_2633);
nand U2711 (N_2711,In_2079,In_1934);
nor U2712 (N_2712,In_2855,In_2034);
xor U2713 (N_2713,In_1601,In_297);
xnor U2714 (N_2714,In_2626,In_835);
xor U2715 (N_2715,In_618,In_2281);
and U2716 (N_2716,In_1134,In_796);
or U2717 (N_2717,In_1632,In_843);
nand U2718 (N_2718,In_54,In_1318);
nor U2719 (N_2719,In_2971,In_1863);
nand U2720 (N_2720,In_510,In_1922);
and U2721 (N_2721,In_873,In_393);
nor U2722 (N_2722,In_2845,In_542);
nand U2723 (N_2723,In_741,In_2038);
or U2724 (N_2724,In_2996,In_992);
or U2725 (N_2725,In_152,In_180);
and U2726 (N_2726,In_1057,In_236);
xor U2727 (N_2727,In_1056,In_2703);
and U2728 (N_2728,In_2353,In_2364);
xnor U2729 (N_2729,In_1494,In_259);
and U2730 (N_2730,In_215,In_1364);
xnor U2731 (N_2731,In_2172,In_1543);
nand U2732 (N_2732,In_1644,In_2292);
and U2733 (N_2733,In_2839,In_2099);
nor U2734 (N_2734,In_1127,In_2202);
nor U2735 (N_2735,In_2045,In_847);
xor U2736 (N_2736,In_2996,In_2912);
nand U2737 (N_2737,In_622,In_2341);
or U2738 (N_2738,In_2045,In_22);
or U2739 (N_2739,In_657,In_2129);
or U2740 (N_2740,In_1353,In_2982);
and U2741 (N_2741,In_588,In_23);
xor U2742 (N_2742,In_2775,In_1919);
or U2743 (N_2743,In_792,In_1044);
nor U2744 (N_2744,In_983,In_2384);
nor U2745 (N_2745,In_1772,In_2566);
xor U2746 (N_2746,In_284,In_303);
or U2747 (N_2747,In_296,In_1304);
xor U2748 (N_2748,In_1739,In_1114);
nand U2749 (N_2749,In_2901,In_1321);
and U2750 (N_2750,In_77,In_287);
and U2751 (N_2751,In_1968,In_1982);
xnor U2752 (N_2752,In_1199,In_2675);
xor U2753 (N_2753,In_20,In_1884);
nor U2754 (N_2754,In_742,In_780);
and U2755 (N_2755,In_2023,In_1307);
or U2756 (N_2756,In_250,In_434);
and U2757 (N_2757,In_981,In_1826);
or U2758 (N_2758,In_2733,In_146);
xor U2759 (N_2759,In_969,In_2010);
and U2760 (N_2760,In_1468,In_1525);
and U2761 (N_2761,In_132,In_1546);
and U2762 (N_2762,In_957,In_2054);
xor U2763 (N_2763,In_1402,In_612);
or U2764 (N_2764,In_2235,In_895);
and U2765 (N_2765,In_1943,In_2260);
and U2766 (N_2766,In_2976,In_1542);
xor U2767 (N_2767,In_1387,In_1443);
nor U2768 (N_2768,In_1194,In_1858);
and U2769 (N_2769,In_1177,In_504);
and U2770 (N_2770,In_1932,In_2513);
and U2771 (N_2771,In_2663,In_2005);
nand U2772 (N_2772,In_1634,In_1360);
or U2773 (N_2773,In_1658,In_735);
xnor U2774 (N_2774,In_1935,In_923);
nand U2775 (N_2775,In_2676,In_2019);
nand U2776 (N_2776,In_2658,In_2246);
nor U2777 (N_2777,In_2783,In_957);
xnor U2778 (N_2778,In_362,In_1338);
or U2779 (N_2779,In_1907,In_1144);
nand U2780 (N_2780,In_1688,In_2584);
nor U2781 (N_2781,In_2244,In_383);
nand U2782 (N_2782,In_1093,In_395);
nand U2783 (N_2783,In_752,In_1548);
xnor U2784 (N_2784,In_1421,In_236);
nor U2785 (N_2785,In_2599,In_2804);
xnor U2786 (N_2786,In_981,In_1737);
xnor U2787 (N_2787,In_2321,In_308);
and U2788 (N_2788,In_41,In_698);
nor U2789 (N_2789,In_2382,In_2299);
xor U2790 (N_2790,In_1882,In_2349);
and U2791 (N_2791,In_1419,In_73);
and U2792 (N_2792,In_2567,In_1474);
xor U2793 (N_2793,In_2533,In_2268);
nand U2794 (N_2794,In_796,In_2103);
and U2795 (N_2795,In_950,In_2801);
nor U2796 (N_2796,In_2660,In_1068);
xnor U2797 (N_2797,In_288,In_1726);
and U2798 (N_2798,In_2203,In_1529);
and U2799 (N_2799,In_2818,In_2489);
nand U2800 (N_2800,In_1729,In_2582);
xor U2801 (N_2801,In_483,In_2322);
nand U2802 (N_2802,In_2099,In_487);
and U2803 (N_2803,In_1360,In_382);
and U2804 (N_2804,In_372,In_1055);
xor U2805 (N_2805,In_1357,In_631);
nor U2806 (N_2806,In_2728,In_580);
or U2807 (N_2807,In_2877,In_1007);
xnor U2808 (N_2808,In_2709,In_1952);
and U2809 (N_2809,In_895,In_2191);
and U2810 (N_2810,In_2939,In_294);
or U2811 (N_2811,In_45,In_66);
and U2812 (N_2812,In_781,In_2379);
nor U2813 (N_2813,In_667,In_2466);
or U2814 (N_2814,In_444,In_966);
or U2815 (N_2815,In_2556,In_2734);
nand U2816 (N_2816,In_1539,In_2237);
nand U2817 (N_2817,In_1221,In_540);
and U2818 (N_2818,In_79,In_2693);
nor U2819 (N_2819,In_2022,In_1514);
nand U2820 (N_2820,In_758,In_2665);
nand U2821 (N_2821,In_438,In_2377);
or U2822 (N_2822,In_2005,In_1786);
nand U2823 (N_2823,In_2219,In_1599);
xnor U2824 (N_2824,In_668,In_1331);
and U2825 (N_2825,In_1992,In_191);
nand U2826 (N_2826,In_1942,In_20);
and U2827 (N_2827,In_896,In_1524);
or U2828 (N_2828,In_2306,In_3);
nand U2829 (N_2829,In_1168,In_1955);
nor U2830 (N_2830,In_395,In_620);
or U2831 (N_2831,In_2466,In_1460);
xor U2832 (N_2832,In_755,In_893);
and U2833 (N_2833,In_647,In_2589);
nand U2834 (N_2834,In_805,In_1645);
nand U2835 (N_2835,In_1783,In_2108);
nor U2836 (N_2836,In_2467,In_1264);
nand U2837 (N_2837,In_1001,In_1919);
and U2838 (N_2838,In_1802,In_1142);
and U2839 (N_2839,In_1197,In_1738);
and U2840 (N_2840,In_2323,In_1774);
or U2841 (N_2841,In_2314,In_447);
and U2842 (N_2842,In_2819,In_881);
nor U2843 (N_2843,In_2397,In_2968);
or U2844 (N_2844,In_1851,In_1606);
xor U2845 (N_2845,In_1666,In_736);
nor U2846 (N_2846,In_2990,In_1551);
nor U2847 (N_2847,In_1554,In_740);
nor U2848 (N_2848,In_2046,In_2831);
nor U2849 (N_2849,In_1309,In_209);
and U2850 (N_2850,In_2395,In_2898);
and U2851 (N_2851,In_609,In_2561);
and U2852 (N_2852,In_2035,In_1299);
nand U2853 (N_2853,In_1817,In_659);
nand U2854 (N_2854,In_2317,In_1492);
nand U2855 (N_2855,In_2645,In_941);
and U2856 (N_2856,In_838,In_701);
nand U2857 (N_2857,In_84,In_2795);
or U2858 (N_2858,In_1999,In_1470);
xnor U2859 (N_2859,In_519,In_443);
nor U2860 (N_2860,In_2183,In_1191);
and U2861 (N_2861,In_2989,In_1018);
nand U2862 (N_2862,In_800,In_2914);
and U2863 (N_2863,In_1836,In_922);
or U2864 (N_2864,In_2818,In_1959);
xnor U2865 (N_2865,In_2655,In_539);
or U2866 (N_2866,In_1270,In_2604);
and U2867 (N_2867,In_2526,In_145);
nand U2868 (N_2868,In_2790,In_248);
or U2869 (N_2869,In_1001,In_1285);
and U2870 (N_2870,In_2156,In_1084);
xnor U2871 (N_2871,In_1759,In_2040);
or U2872 (N_2872,In_634,In_402);
nor U2873 (N_2873,In_2691,In_1811);
nor U2874 (N_2874,In_1654,In_866);
xnor U2875 (N_2875,In_2750,In_1456);
xnor U2876 (N_2876,In_2698,In_2020);
nand U2877 (N_2877,In_2810,In_979);
xor U2878 (N_2878,In_2613,In_330);
nand U2879 (N_2879,In_2488,In_1127);
nand U2880 (N_2880,In_699,In_1821);
xor U2881 (N_2881,In_2783,In_1109);
nor U2882 (N_2882,In_1949,In_1816);
and U2883 (N_2883,In_536,In_300);
xnor U2884 (N_2884,In_2553,In_1163);
xnor U2885 (N_2885,In_2822,In_2476);
xnor U2886 (N_2886,In_2954,In_105);
and U2887 (N_2887,In_2142,In_1538);
xnor U2888 (N_2888,In_1817,In_606);
nor U2889 (N_2889,In_816,In_719);
nor U2890 (N_2890,In_177,In_2060);
nand U2891 (N_2891,In_2767,In_400);
xor U2892 (N_2892,In_1478,In_818);
nand U2893 (N_2893,In_2674,In_352);
or U2894 (N_2894,In_2143,In_713);
nand U2895 (N_2895,In_547,In_1092);
nor U2896 (N_2896,In_1727,In_2660);
and U2897 (N_2897,In_1491,In_2762);
nand U2898 (N_2898,In_1946,In_626);
or U2899 (N_2899,In_585,In_902);
and U2900 (N_2900,In_1053,In_1503);
or U2901 (N_2901,In_532,In_1657);
xor U2902 (N_2902,In_1735,In_231);
nor U2903 (N_2903,In_2241,In_2488);
or U2904 (N_2904,In_2127,In_2116);
and U2905 (N_2905,In_2888,In_783);
and U2906 (N_2906,In_134,In_30);
nand U2907 (N_2907,In_638,In_2735);
nor U2908 (N_2908,In_342,In_2233);
nor U2909 (N_2909,In_1028,In_1059);
and U2910 (N_2910,In_1623,In_1885);
and U2911 (N_2911,In_1865,In_2721);
nand U2912 (N_2912,In_2927,In_2548);
and U2913 (N_2913,In_826,In_731);
and U2914 (N_2914,In_2696,In_1844);
or U2915 (N_2915,In_170,In_195);
nor U2916 (N_2916,In_1925,In_1433);
nand U2917 (N_2917,In_2023,In_862);
xor U2918 (N_2918,In_1139,In_89);
and U2919 (N_2919,In_66,In_847);
nor U2920 (N_2920,In_106,In_1906);
nor U2921 (N_2921,In_548,In_1632);
nand U2922 (N_2922,In_2166,In_1135);
xor U2923 (N_2923,In_1285,In_2251);
or U2924 (N_2924,In_186,In_1466);
and U2925 (N_2925,In_51,In_102);
and U2926 (N_2926,In_1529,In_1901);
and U2927 (N_2927,In_1105,In_1198);
xor U2928 (N_2928,In_688,In_2647);
nor U2929 (N_2929,In_505,In_313);
and U2930 (N_2930,In_1736,In_2338);
or U2931 (N_2931,In_463,In_1289);
or U2932 (N_2932,In_287,In_2528);
nor U2933 (N_2933,In_2922,In_16);
and U2934 (N_2934,In_1373,In_381);
nor U2935 (N_2935,In_1963,In_352);
nor U2936 (N_2936,In_2717,In_1104);
nand U2937 (N_2937,In_2596,In_877);
and U2938 (N_2938,In_691,In_1112);
or U2939 (N_2939,In_1055,In_2843);
nor U2940 (N_2940,In_1369,In_550);
xnor U2941 (N_2941,In_2704,In_2302);
nor U2942 (N_2942,In_2346,In_580);
nor U2943 (N_2943,In_1218,In_1651);
or U2944 (N_2944,In_1789,In_1616);
nand U2945 (N_2945,In_2586,In_1161);
nand U2946 (N_2946,In_2465,In_2708);
and U2947 (N_2947,In_1359,In_893);
xnor U2948 (N_2948,In_616,In_760);
xnor U2949 (N_2949,In_337,In_512);
nor U2950 (N_2950,In_2965,In_1720);
nand U2951 (N_2951,In_1939,In_1123);
or U2952 (N_2952,In_1873,In_2740);
and U2953 (N_2953,In_691,In_2571);
or U2954 (N_2954,In_962,In_691);
nor U2955 (N_2955,In_924,In_1564);
nand U2956 (N_2956,In_1490,In_1627);
nor U2957 (N_2957,In_2718,In_2204);
or U2958 (N_2958,In_648,In_1781);
or U2959 (N_2959,In_63,In_31);
xor U2960 (N_2960,In_1245,In_604);
xnor U2961 (N_2961,In_547,In_2787);
and U2962 (N_2962,In_2699,In_2993);
xor U2963 (N_2963,In_2033,In_1669);
or U2964 (N_2964,In_2354,In_1325);
nand U2965 (N_2965,In_656,In_2509);
nor U2966 (N_2966,In_860,In_1040);
nand U2967 (N_2967,In_224,In_1601);
nor U2968 (N_2968,In_1611,In_1958);
nand U2969 (N_2969,In_1699,In_2287);
or U2970 (N_2970,In_2738,In_2449);
nand U2971 (N_2971,In_1603,In_1552);
or U2972 (N_2972,In_25,In_2939);
nor U2973 (N_2973,In_898,In_2160);
or U2974 (N_2974,In_1867,In_1840);
or U2975 (N_2975,In_956,In_443);
nor U2976 (N_2976,In_1405,In_196);
xnor U2977 (N_2977,In_2525,In_2707);
nor U2978 (N_2978,In_307,In_2802);
and U2979 (N_2979,In_2637,In_1733);
or U2980 (N_2980,In_2043,In_2442);
nand U2981 (N_2981,In_2835,In_1609);
nor U2982 (N_2982,In_2558,In_270);
xor U2983 (N_2983,In_1522,In_2017);
nor U2984 (N_2984,In_2194,In_827);
nor U2985 (N_2985,In_2231,In_1687);
or U2986 (N_2986,In_866,In_2606);
nand U2987 (N_2987,In_2827,In_1657);
or U2988 (N_2988,In_1528,In_2606);
and U2989 (N_2989,In_2720,In_2979);
or U2990 (N_2990,In_1090,In_200);
nor U2991 (N_2991,In_2126,In_606);
or U2992 (N_2992,In_210,In_1265);
or U2993 (N_2993,In_2846,In_1320);
xnor U2994 (N_2994,In_2657,In_2240);
and U2995 (N_2995,In_2997,In_1128);
and U2996 (N_2996,In_2504,In_286);
xor U2997 (N_2997,In_2555,In_879);
or U2998 (N_2998,In_2360,In_1265);
nand U2999 (N_2999,In_591,In_563);
nand U3000 (N_3000,In_1760,In_718);
nand U3001 (N_3001,In_1934,In_571);
and U3002 (N_3002,In_2986,In_1689);
or U3003 (N_3003,In_1336,In_1739);
nand U3004 (N_3004,In_408,In_2532);
nor U3005 (N_3005,In_2083,In_2531);
and U3006 (N_3006,In_549,In_1731);
or U3007 (N_3007,In_439,In_59);
xor U3008 (N_3008,In_2745,In_1977);
xor U3009 (N_3009,In_2318,In_1118);
nor U3010 (N_3010,In_2221,In_320);
and U3011 (N_3011,In_2424,In_1722);
nand U3012 (N_3012,In_1324,In_1280);
and U3013 (N_3013,In_2359,In_1225);
nor U3014 (N_3014,In_1402,In_2962);
nor U3015 (N_3015,In_1504,In_2567);
and U3016 (N_3016,In_2251,In_830);
nand U3017 (N_3017,In_2026,In_1631);
xor U3018 (N_3018,In_1513,In_1501);
and U3019 (N_3019,In_450,In_676);
nor U3020 (N_3020,In_1611,In_654);
or U3021 (N_3021,In_463,In_1869);
or U3022 (N_3022,In_939,In_589);
nor U3023 (N_3023,In_1293,In_713);
and U3024 (N_3024,In_2870,In_1572);
and U3025 (N_3025,In_2424,In_361);
xor U3026 (N_3026,In_563,In_1540);
and U3027 (N_3027,In_2933,In_2687);
nand U3028 (N_3028,In_2303,In_2148);
xnor U3029 (N_3029,In_1620,In_61);
and U3030 (N_3030,In_1045,In_1909);
nor U3031 (N_3031,In_1355,In_2583);
nand U3032 (N_3032,In_1870,In_2265);
nand U3033 (N_3033,In_1712,In_631);
xor U3034 (N_3034,In_43,In_1935);
nor U3035 (N_3035,In_808,In_1329);
and U3036 (N_3036,In_732,In_376);
nand U3037 (N_3037,In_820,In_1741);
or U3038 (N_3038,In_2035,In_494);
xor U3039 (N_3039,In_441,In_789);
or U3040 (N_3040,In_2513,In_959);
nor U3041 (N_3041,In_1262,In_182);
nand U3042 (N_3042,In_255,In_2035);
or U3043 (N_3043,In_1822,In_2900);
nand U3044 (N_3044,In_2788,In_367);
and U3045 (N_3045,In_2679,In_1744);
nor U3046 (N_3046,In_518,In_2612);
nand U3047 (N_3047,In_2858,In_1126);
or U3048 (N_3048,In_2963,In_304);
or U3049 (N_3049,In_1864,In_1786);
nand U3050 (N_3050,In_1409,In_2762);
nor U3051 (N_3051,In_1063,In_257);
nor U3052 (N_3052,In_641,In_1396);
or U3053 (N_3053,In_2316,In_1164);
or U3054 (N_3054,In_2518,In_1795);
xor U3055 (N_3055,In_1244,In_1524);
and U3056 (N_3056,In_2381,In_168);
or U3057 (N_3057,In_1993,In_1212);
nor U3058 (N_3058,In_2576,In_1783);
nor U3059 (N_3059,In_630,In_2754);
xnor U3060 (N_3060,In_2877,In_1400);
nand U3061 (N_3061,In_2622,In_1118);
nor U3062 (N_3062,In_2405,In_2726);
xnor U3063 (N_3063,In_1260,In_2275);
and U3064 (N_3064,In_2817,In_403);
nand U3065 (N_3065,In_2784,In_2838);
or U3066 (N_3066,In_425,In_1063);
and U3067 (N_3067,In_2255,In_545);
nor U3068 (N_3068,In_2665,In_851);
and U3069 (N_3069,In_27,In_1512);
nor U3070 (N_3070,In_1557,In_2622);
nand U3071 (N_3071,In_2197,In_1300);
nor U3072 (N_3072,In_2514,In_2938);
xnor U3073 (N_3073,In_630,In_926);
nand U3074 (N_3074,In_1812,In_1582);
and U3075 (N_3075,In_2874,In_1912);
and U3076 (N_3076,In_2009,In_2357);
and U3077 (N_3077,In_1630,In_2788);
nand U3078 (N_3078,In_432,In_2401);
xor U3079 (N_3079,In_858,In_1410);
nor U3080 (N_3080,In_1392,In_1927);
nor U3081 (N_3081,In_313,In_1548);
and U3082 (N_3082,In_6,In_1948);
xor U3083 (N_3083,In_2993,In_977);
nor U3084 (N_3084,In_1143,In_2016);
or U3085 (N_3085,In_335,In_658);
nand U3086 (N_3086,In_2576,In_2558);
xor U3087 (N_3087,In_588,In_267);
nand U3088 (N_3088,In_1645,In_573);
or U3089 (N_3089,In_1508,In_1533);
and U3090 (N_3090,In_404,In_2067);
nor U3091 (N_3091,In_2013,In_1783);
nor U3092 (N_3092,In_427,In_802);
xor U3093 (N_3093,In_52,In_2272);
xor U3094 (N_3094,In_5,In_426);
and U3095 (N_3095,In_1000,In_2508);
xnor U3096 (N_3096,In_116,In_402);
and U3097 (N_3097,In_280,In_2007);
xor U3098 (N_3098,In_27,In_787);
nor U3099 (N_3099,In_2451,In_1965);
and U3100 (N_3100,In_2573,In_831);
nand U3101 (N_3101,In_1837,In_765);
nor U3102 (N_3102,In_389,In_2054);
xor U3103 (N_3103,In_2319,In_351);
and U3104 (N_3104,In_229,In_902);
xnor U3105 (N_3105,In_1961,In_19);
nand U3106 (N_3106,In_2862,In_1422);
and U3107 (N_3107,In_2577,In_2638);
or U3108 (N_3108,In_735,In_1252);
or U3109 (N_3109,In_1973,In_122);
and U3110 (N_3110,In_109,In_2011);
xnor U3111 (N_3111,In_85,In_2247);
nand U3112 (N_3112,In_1438,In_2505);
nand U3113 (N_3113,In_1716,In_2824);
and U3114 (N_3114,In_2362,In_105);
nand U3115 (N_3115,In_1050,In_2335);
xnor U3116 (N_3116,In_1544,In_376);
nor U3117 (N_3117,In_443,In_270);
nor U3118 (N_3118,In_2067,In_1068);
nor U3119 (N_3119,In_2875,In_187);
xor U3120 (N_3120,In_2456,In_2975);
xnor U3121 (N_3121,In_551,In_832);
nand U3122 (N_3122,In_2067,In_1418);
nor U3123 (N_3123,In_2109,In_1503);
nor U3124 (N_3124,In_1915,In_7);
nor U3125 (N_3125,In_2962,In_1837);
nand U3126 (N_3126,In_682,In_1119);
nand U3127 (N_3127,In_2829,In_1881);
and U3128 (N_3128,In_2236,In_2579);
nand U3129 (N_3129,In_490,In_2904);
nand U3130 (N_3130,In_2743,In_1163);
or U3131 (N_3131,In_316,In_2851);
nor U3132 (N_3132,In_2178,In_552);
xnor U3133 (N_3133,In_161,In_23);
xnor U3134 (N_3134,In_2286,In_1127);
or U3135 (N_3135,In_2286,In_2436);
nand U3136 (N_3136,In_1281,In_1322);
nor U3137 (N_3137,In_568,In_74);
or U3138 (N_3138,In_2893,In_1327);
and U3139 (N_3139,In_867,In_452);
or U3140 (N_3140,In_2496,In_316);
nand U3141 (N_3141,In_1215,In_1436);
nand U3142 (N_3142,In_2037,In_160);
xnor U3143 (N_3143,In_2387,In_1260);
nor U3144 (N_3144,In_2538,In_1374);
xor U3145 (N_3145,In_2507,In_619);
and U3146 (N_3146,In_451,In_2070);
nand U3147 (N_3147,In_1471,In_1242);
or U3148 (N_3148,In_1852,In_1346);
nor U3149 (N_3149,In_2836,In_979);
or U3150 (N_3150,In_2429,In_2012);
or U3151 (N_3151,In_126,In_122);
xor U3152 (N_3152,In_151,In_1839);
xnor U3153 (N_3153,In_1623,In_2511);
nor U3154 (N_3154,In_538,In_1978);
nor U3155 (N_3155,In_1394,In_1087);
nand U3156 (N_3156,In_1194,In_492);
or U3157 (N_3157,In_2496,In_452);
nor U3158 (N_3158,In_2308,In_720);
xnor U3159 (N_3159,In_518,In_879);
xnor U3160 (N_3160,In_271,In_1443);
xnor U3161 (N_3161,In_2798,In_1813);
and U3162 (N_3162,In_1912,In_1708);
or U3163 (N_3163,In_868,In_2204);
and U3164 (N_3164,In_1714,In_494);
xor U3165 (N_3165,In_1828,In_644);
nand U3166 (N_3166,In_1960,In_1659);
or U3167 (N_3167,In_681,In_787);
nor U3168 (N_3168,In_368,In_753);
xor U3169 (N_3169,In_2961,In_2709);
or U3170 (N_3170,In_2643,In_1989);
xor U3171 (N_3171,In_2593,In_1702);
and U3172 (N_3172,In_2027,In_1556);
and U3173 (N_3173,In_2238,In_1271);
xor U3174 (N_3174,In_725,In_1382);
nand U3175 (N_3175,In_199,In_349);
or U3176 (N_3176,In_818,In_2270);
or U3177 (N_3177,In_761,In_2538);
and U3178 (N_3178,In_865,In_202);
and U3179 (N_3179,In_1752,In_2870);
nor U3180 (N_3180,In_2786,In_202);
or U3181 (N_3181,In_727,In_2826);
nor U3182 (N_3182,In_924,In_1340);
xnor U3183 (N_3183,In_1851,In_2063);
nand U3184 (N_3184,In_1827,In_1668);
nand U3185 (N_3185,In_1213,In_376);
or U3186 (N_3186,In_1780,In_176);
xnor U3187 (N_3187,In_732,In_1638);
nand U3188 (N_3188,In_1374,In_695);
and U3189 (N_3189,In_989,In_2313);
nor U3190 (N_3190,In_2049,In_2151);
or U3191 (N_3191,In_1311,In_850);
or U3192 (N_3192,In_1327,In_346);
and U3193 (N_3193,In_104,In_790);
nor U3194 (N_3194,In_629,In_1263);
xnor U3195 (N_3195,In_2621,In_2053);
xnor U3196 (N_3196,In_1668,In_355);
nor U3197 (N_3197,In_1578,In_2873);
nand U3198 (N_3198,In_657,In_2562);
and U3199 (N_3199,In_2520,In_564);
xnor U3200 (N_3200,In_418,In_212);
or U3201 (N_3201,In_127,In_1891);
xor U3202 (N_3202,In_198,In_1134);
nand U3203 (N_3203,In_871,In_597);
and U3204 (N_3204,In_1821,In_406);
nand U3205 (N_3205,In_1597,In_1284);
or U3206 (N_3206,In_2290,In_634);
or U3207 (N_3207,In_2553,In_1566);
or U3208 (N_3208,In_2278,In_900);
nand U3209 (N_3209,In_2540,In_2356);
or U3210 (N_3210,In_1056,In_1809);
nor U3211 (N_3211,In_1092,In_192);
nand U3212 (N_3212,In_1579,In_1056);
xor U3213 (N_3213,In_2138,In_119);
xnor U3214 (N_3214,In_307,In_2963);
xnor U3215 (N_3215,In_2975,In_1433);
and U3216 (N_3216,In_1836,In_2000);
xor U3217 (N_3217,In_1209,In_2042);
xnor U3218 (N_3218,In_2164,In_133);
nand U3219 (N_3219,In_195,In_635);
and U3220 (N_3220,In_2534,In_1965);
xor U3221 (N_3221,In_40,In_1145);
nor U3222 (N_3222,In_2156,In_1982);
xor U3223 (N_3223,In_1905,In_2670);
or U3224 (N_3224,In_924,In_1357);
or U3225 (N_3225,In_736,In_110);
or U3226 (N_3226,In_2281,In_1611);
and U3227 (N_3227,In_1036,In_2700);
nand U3228 (N_3228,In_2540,In_770);
nor U3229 (N_3229,In_576,In_1455);
and U3230 (N_3230,In_2676,In_485);
or U3231 (N_3231,In_836,In_2843);
nand U3232 (N_3232,In_628,In_633);
nand U3233 (N_3233,In_2523,In_786);
nand U3234 (N_3234,In_296,In_2193);
or U3235 (N_3235,In_2654,In_1787);
or U3236 (N_3236,In_1753,In_2287);
or U3237 (N_3237,In_681,In_1273);
and U3238 (N_3238,In_1517,In_1836);
nand U3239 (N_3239,In_1948,In_2538);
or U3240 (N_3240,In_1900,In_2057);
nand U3241 (N_3241,In_73,In_1524);
and U3242 (N_3242,In_1693,In_751);
and U3243 (N_3243,In_2246,In_97);
or U3244 (N_3244,In_561,In_759);
nand U3245 (N_3245,In_1204,In_2106);
and U3246 (N_3246,In_579,In_1650);
or U3247 (N_3247,In_1947,In_1071);
xor U3248 (N_3248,In_70,In_1786);
nand U3249 (N_3249,In_957,In_323);
nor U3250 (N_3250,In_1236,In_2267);
nor U3251 (N_3251,In_294,In_1719);
nand U3252 (N_3252,In_1794,In_1676);
xor U3253 (N_3253,In_2130,In_1419);
and U3254 (N_3254,In_246,In_348);
and U3255 (N_3255,In_2699,In_1050);
xor U3256 (N_3256,In_554,In_1866);
and U3257 (N_3257,In_1113,In_2431);
nor U3258 (N_3258,In_1271,In_2679);
and U3259 (N_3259,In_826,In_1854);
xnor U3260 (N_3260,In_1180,In_346);
or U3261 (N_3261,In_1565,In_12);
xor U3262 (N_3262,In_127,In_2930);
and U3263 (N_3263,In_1767,In_1505);
xor U3264 (N_3264,In_1501,In_869);
nand U3265 (N_3265,In_1663,In_2866);
or U3266 (N_3266,In_1180,In_2515);
or U3267 (N_3267,In_1343,In_2135);
xor U3268 (N_3268,In_2644,In_392);
or U3269 (N_3269,In_347,In_2050);
or U3270 (N_3270,In_882,In_177);
nand U3271 (N_3271,In_2428,In_2076);
xor U3272 (N_3272,In_2124,In_995);
and U3273 (N_3273,In_585,In_1841);
and U3274 (N_3274,In_940,In_1687);
or U3275 (N_3275,In_2656,In_518);
nand U3276 (N_3276,In_372,In_130);
and U3277 (N_3277,In_2508,In_726);
xor U3278 (N_3278,In_911,In_28);
xor U3279 (N_3279,In_1795,In_1568);
xnor U3280 (N_3280,In_2359,In_1105);
xnor U3281 (N_3281,In_225,In_2635);
and U3282 (N_3282,In_245,In_174);
nand U3283 (N_3283,In_901,In_1649);
or U3284 (N_3284,In_2529,In_170);
xor U3285 (N_3285,In_1360,In_1679);
and U3286 (N_3286,In_1958,In_578);
nand U3287 (N_3287,In_2681,In_2004);
or U3288 (N_3288,In_48,In_1969);
or U3289 (N_3289,In_1836,In_2384);
nor U3290 (N_3290,In_657,In_166);
nand U3291 (N_3291,In_1508,In_2014);
and U3292 (N_3292,In_697,In_1359);
or U3293 (N_3293,In_857,In_637);
or U3294 (N_3294,In_2568,In_2120);
xor U3295 (N_3295,In_572,In_1347);
and U3296 (N_3296,In_2543,In_2301);
or U3297 (N_3297,In_1590,In_2957);
nor U3298 (N_3298,In_2680,In_1638);
and U3299 (N_3299,In_2028,In_78);
or U3300 (N_3300,In_1750,In_894);
nand U3301 (N_3301,In_167,In_944);
xnor U3302 (N_3302,In_2963,In_2147);
xnor U3303 (N_3303,In_815,In_96);
or U3304 (N_3304,In_1882,In_2830);
nor U3305 (N_3305,In_959,In_323);
xor U3306 (N_3306,In_364,In_321);
and U3307 (N_3307,In_26,In_1201);
and U3308 (N_3308,In_2156,In_1871);
nor U3309 (N_3309,In_117,In_2019);
nand U3310 (N_3310,In_1986,In_709);
nor U3311 (N_3311,In_1413,In_2347);
nor U3312 (N_3312,In_232,In_1151);
nor U3313 (N_3313,In_1366,In_1961);
nand U3314 (N_3314,In_1758,In_2965);
xnor U3315 (N_3315,In_1458,In_2916);
nor U3316 (N_3316,In_2935,In_29);
and U3317 (N_3317,In_2769,In_263);
or U3318 (N_3318,In_562,In_1125);
or U3319 (N_3319,In_414,In_2662);
and U3320 (N_3320,In_301,In_1815);
nand U3321 (N_3321,In_2191,In_1971);
or U3322 (N_3322,In_483,In_2574);
nor U3323 (N_3323,In_1610,In_2925);
nor U3324 (N_3324,In_2260,In_2857);
nor U3325 (N_3325,In_190,In_990);
xnor U3326 (N_3326,In_1000,In_1008);
nand U3327 (N_3327,In_1754,In_193);
nor U3328 (N_3328,In_418,In_1043);
nor U3329 (N_3329,In_724,In_798);
xor U3330 (N_3330,In_2062,In_533);
xnor U3331 (N_3331,In_727,In_1531);
nand U3332 (N_3332,In_1686,In_804);
or U3333 (N_3333,In_28,In_531);
nor U3334 (N_3334,In_2219,In_2045);
xor U3335 (N_3335,In_80,In_1785);
nand U3336 (N_3336,In_465,In_2537);
and U3337 (N_3337,In_2082,In_132);
or U3338 (N_3338,In_2658,In_1064);
nor U3339 (N_3339,In_2012,In_754);
nand U3340 (N_3340,In_2259,In_1995);
xor U3341 (N_3341,In_924,In_739);
nor U3342 (N_3342,In_1654,In_2016);
nor U3343 (N_3343,In_1982,In_2836);
and U3344 (N_3344,In_86,In_1522);
nand U3345 (N_3345,In_1385,In_2013);
or U3346 (N_3346,In_745,In_1724);
and U3347 (N_3347,In_1299,In_618);
xor U3348 (N_3348,In_2613,In_2863);
or U3349 (N_3349,In_680,In_84);
xnor U3350 (N_3350,In_2526,In_611);
xnor U3351 (N_3351,In_1295,In_2152);
xnor U3352 (N_3352,In_2700,In_714);
nor U3353 (N_3353,In_1178,In_43);
nand U3354 (N_3354,In_686,In_1343);
nor U3355 (N_3355,In_1601,In_1996);
and U3356 (N_3356,In_974,In_1005);
nand U3357 (N_3357,In_1154,In_2812);
and U3358 (N_3358,In_1064,In_824);
xnor U3359 (N_3359,In_407,In_1579);
and U3360 (N_3360,In_1701,In_431);
and U3361 (N_3361,In_2559,In_558);
nor U3362 (N_3362,In_2438,In_959);
and U3363 (N_3363,In_1166,In_728);
xnor U3364 (N_3364,In_1743,In_2896);
or U3365 (N_3365,In_345,In_558);
or U3366 (N_3366,In_1790,In_472);
nand U3367 (N_3367,In_347,In_196);
xor U3368 (N_3368,In_373,In_1642);
and U3369 (N_3369,In_2076,In_1239);
nor U3370 (N_3370,In_356,In_1960);
nand U3371 (N_3371,In_2041,In_2157);
nor U3372 (N_3372,In_1410,In_1078);
or U3373 (N_3373,In_1315,In_1839);
xor U3374 (N_3374,In_637,In_2830);
nor U3375 (N_3375,In_2105,In_376);
xnor U3376 (N_3376,In_2432,In_1119);
or U3377 (N_3377,In_825,In_2314);
xor U3378 (N_3378,In_678,In_2092);
xor U3379 (N_3379,In_2,In_599);
nor U3380 (N_3380,In_79,In_1946);
xnor U3381 (N_3381,In_1524,In_2359);
or U3382 (N_3382,In_156,In_2769);
and U3383 (N_3383,In_959,In_577);
and U3384 (N_3384,In_2124,In_2182);
nand U3385 (N_3385,In_2024,In_2911);
nand U3386 (N_3386,In_1415,In_811);
or U3387 (N_3387,In_967,In_1795);
or U3388 (N_3388,In_1782,In_1901);
xnor U3389 (N_3389,In_2802,In_2235);
and U3390 (N_3390,In_1820,In_827);
and U3391 (N_3391,In_770,In_1829);
and U3392 (N_3392,In_43,In_2603);
and U3393 (N_3393,In_2541,In_158);
nor U3394 (N_3394,In_2018,In_1790);
xnor U3395 (N_3395,In_75,In_2615);
or U3396 (N_3396,In_1869,In_2551);
nand U3397 (N_3397,In_2905,In_2102);
nor U3398 (N_3398,In_2687,In_1191);
xnor U3399 (N_3399,In_569,In_2425);
and U3400 (N_3400,In_2078,In_1140);
nor U3401 (N_3401,In_357,In_2858);
nand U3402 (N_3402,In_138,In_86);
nand U3403 (N_3403,In_1654,In_214);
nor U3404 (N_3404,In_1336,In_2204);
nor U3405 (N_3405,In_552,In_987);
or U3406 (N_3406,In_17,In_2563);
nand U3407 (N_3407,In_2652,In_1155);
nand U3408 (N_3408,In_1181,In_2918);
nand U3409 (N_3409,In_2837,In_1986);
and U3410 (N_3410,In_174,In_2324);
nand U3411 (N_3411,In_109,In_263);
or U3412 (N_3412,In_1867,In_2523);
and U3413 (N_3413,In_1570,In_1528);
or U3414 (N_3414,In_2415,In_180);
and U3415 (N_3415,In_1564,In_1698);
or U3416 (N_3416,In_918,In_1515);
nor U3417 (N_3417,In_2802,In_1904);
xor U3418 (N_3418,In_2382,In_531);
nor U3419 (N_3419,In_1872,In_2059);
xor U3420 (N_3420,In_2576,In_116);
xor U3421 (N_3421,In_2688,In_407);
nor U3422 (N_3422,In_2838,In_262);
xnor U3423 (N_3423,In_2806,In_2986);
nand U3424 (N_3424,In_1813,In_1642);
or U3425 (N_3425,In_1752,In_2453);
nor U3426 (N_3426,In_1391,In_2992);
nand U3427 (N_3427,In_2889,In_1832);
and U3428 (N_3428,In_1094,In_2173);
nand U3429 (N_3429,In_1715,In_551);
and U3430 (N_3430,In_990,In_266);
nor U3431 (N_3431,In_2341,In_1724);
or U3432 (N_3432,In_1903,In_1521);
and U3433 (N_3433,In_2482,In_1506);
or U3434 (N_3434,In_2004,In_2970);
or U3435 (N_3435,In_999,In_233);
nor U3436 (N_3436,In_1503,In_2587);
and U3437 (N_3437,In_1856,In_702);
and U3438 (N_3438,In_2205,In_471);
xnor U3439 (N_3439,In_1583,In_1972);
xor U3440 (N_3440,In_567,In_191);
nand U3441 (N_3441,In_832,In_2239);
xnor U3442 (N_3442,In_478,In_1534);
or U3443 (N_3443,In_1494,In_2326);
nand U3444 (N_3444,In_369,In_815);
and U3445 (N_3445,In_1838,In_1207);
nor U3446 (N_3446,In_326,In_2895);
nor U3447 (N_3447,In_1704,In_1099);
nor U3448 (N_3448,In_2333,In_1199);
and U3449 (N_3449,In_2779,In_2495);
nand U3450 (N_3450,In_826,In_912);
xor U3451 (N_3451,In_2229,In_2315);
or U3452 (N_3452,In_2548,In_2317);
nor U3453 (N_3453,In_422,In_543);
nor U3454 (N_3454,In_2135,In_620);
or U3455 (N_3455,In_798,In_1981);
nand U3456 (N_3456,In_1130,In_2522);
and U3457 (N_3457,In_232,In_2341);
or U3458 (N_3458,In_2888,In_750);
xnor U3459 (N_3459,In_1620,In_2734);
xor U3460 (N_3460,In_1635,In_1203);
nor U3461 (N_3461,In_2120,In_786);
nand U3462 (N_3462,In_857,In_1173);
nand U3463 (N_3463,In_2046,In_1074);
nand U3464 (N_3464,In_2555,In_105);
xor U3465 (N_3465,In_397,In_2957);
nand U3466 (N_3466,In_2718,In_1804);
xnor U3467 (N_3467,In_1737,In_902);
or U3468 (N_3468,In_971,In_789);
nor U3469 (N_3469,In_107,In_1318);
nor U3470 (N_3470,In_1853,In_33);
nor U3471 (N_3471,In_2295,In_171);
xnor U3472 (N_3472,In_2933,In_3);
xnor U3473 (N_3473,In_1284,In_1356);
nor U3474 (N_3474,In_1314,In_2343);
and U3475 (N_3475,In_1451,In_2891);
xnor U3476 (N_3476,In_2167,In_1431);
or U3477 (N_3477,In_1173,In_1784);
or U3478 (N_3478,In_2942,In_2937);
nor U3479 (N_3479,In_1070,In_1763);
xnor U3480 (N_3480,In_2057,In_1380);
nand U3481 (N_3481,In_1467,In_2302);
xor U3482 (N_3482,In_2602,In_2142);
and U3483 (N_3483,In_74,In_2476);
nor U3484 (N_3484,In_1121,In_1323);
nand U3485 (N_3485,In_1768,In_2715);
and U3486 (N_3486,In_2499,In_1417);
nor U3487 (N_3487,In_399,In_1387);
and U3488 (N_3488,In_301,In_1801);
nand U3489 (N_3489,In_996,In_1489);
nor U3490 (N_3490,In_1396,In_1021);
nand U3491 (N_3491,In_2479,In_598);
nand U3492 (N_3492,In_496,In_1116);
xor U3493 (N_3493,In_1200,In_2370);
or U3494 (N_3494,In_2552,In_1213);
xor U3495 (N_3495,In_1244,In_2069);
xnor U3496 (N_3496,In_300,In_28);
xor U3497 (N_3497,In_1582,In_1999);
and U3498 (N_3498,In_1329,In_1381);
xnor U3499 (N_3499,In_894,In_840);
nor U3500 (N_3500,In_2429,In_1351);
nand U3501 (N_3501,In_1864,In_650);
nor U3502 (N_3502,In_2140,In_1691);
nor U3503 (N_3503,In_2592,In_1936);
or U3504 (N_3504,In_1601,In_2765);
xor U3505 (N_3505,In_1774,In_1089);
or U3506 (N_3506,In_1654,In_2124);
and U3507 (N_3507,In_1845,In_2827);
xnor U3508 (N_3508,In_555,In_1232);
xor U3509 (N_3509,In_1644,In_1888);
nand U3510 (N_3510,In_322,In_2450);
nand U3511 (N_3511,In_364,In_149);
xor U3512 (N_3512,In_671,In_230);
nor U3513 (N_3513,In_971,In_1053);
nand U3514 (N_3514,In_2871,In_2947);
nand U3515 (N_3515,In_520,In_2743);
nor U3516 (N_3516,In_1304,In_2835);
or U3517 (N_3517,In_910,In_663);
nor U3518 (N_3518,In_123,In_2372);
xor U3519 (N_3519,In_1966,In_2088);
nand U3520 (N_3520,In_45,In_1899);
and U3521 (N_3521,In_1742,In_2360);
xor U3522 (N_3522,In_324,In_446);
nand U3523 (N_3523,In_709,In_2137);
or U3524 (N_3524,In_364,In_1043);
nor U3525 (N_3525,In_1811,In_2015);
xnor U3526 (N_3526,In_1977,In_2759);
xnor U3527 (N_3527,In_1369,In_1124);
and U3528 (N_3528,In_61,In_882);
nor U3529 (N_3529,In_1990,In_1239);
nor U3530 (N_3530,In_1909,In_992);
nand U3531 (N_3531,In_1758,In_984);
nand U3532 (N_3532,In_2869,In_2169);
or U3533 (N_3533,In_2484,In_2639);
or U3534 (N_3534,In_1878,In_1463);
xor U3535 (N_3535,In_1212,In_2809);
and U3536 (N_3536,In_1937,In_1322);
and U3537 (N_3537,In_1084,In_2798);
nand U3538 (N_3538,In_680,In_2664);
nor U3539 (N_3539,In_2906,In_2007);
nand U3540 (N_3540,In_33,In_956);
or U3541 (N_3541,In_883,In_834);
nand U3542 (N_3542,In_1337,In_2600);
or U3543 (N_3543,In_1013,In_500);
nor U3544 (N_3544,In_2706,In_385);
xor U3545 (N_3545,In_1052,In_2059);
and U3546 (N_3546,In_2996,In_1908);
and U3547 (N_3547,In_1071,In_2307);
nor U3548 (N_3548,In_138,In_1405);
nor U3549 (N_3549,In_285,In_2375);
or U3550 (N_3550,In_1401,In_1653);
xor U3551 (N_3551,In_878,In_870);
and U3552 (N_3552,In_1000,In_2550);
and U3553 (N_3553,In_1123,In_1487);
nand U3554 (N_3554,In_652,In_2695);
nand U3555 (N_3555,In_1257,In_1866);
or U3556 (N_3556,In_1944,In_2161);
and U3557 (N_3557,In_260,In_1351);
nor U3558 (N_3558,In_1385,In_698);
nor U3559 (N_3559,In_209,In_2958);
or U3560 (N_3560,In_2117,In_962);
nor U3561 (N_3561,In_2852,In_740);
nand U3562 (N_3562,In_1780,In_2239);
nor U3563 (N_3563,In_2748,In_1974);
xor U3564 (N_3564,In_145,In_2181);
or U3565 (N_3565,In_2809,In_2053);
nand U3566 (N_3566,In_2654,In_2945);
xnor U3567 (N_3567,In_1587,In_2858);
or U3568 (N_3568,In_2472,In_1396);
and U3569 (N_3569,In_1236,In_615);
and U3570 (N_3570,In_791,In_2049);
nand U3571 (N_3571,In_309,In_1045);
xor U3572 (N_3572,In_2865,In_2269);
xnor U3573 (N_3573,In_1917,In_118);
nand U3574 (N_3574,In_1174,In_865);
and U3575 (N_3575,In_225,In_956);
nor U3576 (N_3576,In_1868,In_2501);
nor U3577 (N_3577,In_1819,In_2026);
or U3578 (N_3578,In_1893,In_2272);
and U3579 (N_3579,In_236,In_2422);
and U3580 (N_3580,In_2519,In_986);
xnor U3581 (N_3581,In_2295,In_436);
xnor U3582 (N_3582,In_461,In_2889);
nor U3583 (N_3583,In_1087,In_2488);
or U3584 (N_3584,In_741,In_1444);
and U3585 (N_3585,In_1641,In_780);
nor U3586 (N_3586,In_711,In_319);
xor U3587 (N_3587,In_1509,In_2257);
nor U3588 (N_3588,In_1542,In_2975);
or U3589 (N_3589,In_211,In_2646);
nand U3590 (N_3590,In_2910,In_2953);
or U3591 (N_3591,In_2886,In_2394);
xnor U3592 (N_3592,In_700,In_1202);
and U3593 (N_3593,In_2398,In_2873);
nand U3594 (N_3594,In_1667,In_729);
and U3595 (N_3595,In_1,In_1169);
xnor U3596 (N_3596,In_2957,In_2530);
and U3597 (N_3597,In_1830,In_1081);
or U3598 (N_3598,In_2276,In_2708);
and U3599 (N_3599,In_907,In_645);
nor U3600 (N_3600,In_645,In_1971);
xnor U3601 (N_3601,In_1563,In_665);
nand U3602 (N_3602,In_1225,In_1250);
xnor U3603 (N_3603,In_1675,In_1622);
xnor U3604 (N_3604,In_279,In_1103);
nand U3605 (N_3605,In_1582,In_2704);
or U3606 (N_3606,In_224,In_597);
nor U3607 (N_3607,In_1640,In_1398);
nand U3608 (N_3608,In_2536,In_1837);
xor U3609 (N_3609,In_422,In_2035);
or U3610 (N_3610,In_655,In_1448);
or U3611 (N_3611,In_919,In_2201);
nand U3612 (N_3612,In_1554,In_281);
and U3613 (N_3613,In_418,In_40);
xor U3614 (N_3614,In_2463,In_2348);
xnor U3615 (N_3615,In_2454,In_1589);
nor U3616 (N_3616,In_732,In_1770);
xnor U3617 (N_3617,In_1564,In_2250);
nor U3618 (N_3618,In_1489,In_2351);
nor U3619 (N_3619,In_1837,In_1378);
and U3620 (N_3620,In_1154,In_2520);
and U3621 (N_3621,In_576,In_549);
nor U3622 (N_3622,In_1548,In_1079);
or U3623 (N_3623,In_438,In_2890);
nor U3624 (N_3624,In_1812,In_710);
nor U3625 (N_3625,In_2617,In_1257);
and U3626 (N_3626,In_395,In_1281);
xnor U3627 (N_3627,In_637,In_2944);
or U3628 (N_3628,In_2091,In_1131);
and U3629 (N_3629,In_2812,In_641);
and U3630 (N_3630,In_2282,In_724);
and U3631 (N_3631,In_158,In_1676);
nor U3632 (N_3632,In_2859,In_1347);
or U3633 (N_3633,In_2938,In_1536);
nor U3634 (N_3634,In_2209,In_632);
and U3635 (N_3635,In_1820,In_1616);
nor U3636 (N_3636,In_11,In_295);
and U3637 (N_3637,In_195,In_1079);
nor U3638 (N_3638,In_723,In_2281);
nand U3639 (N_3639,In_288,In_1625);
or U3640 (N_3640,In_2422,In_2535);
or U3641 (N_3641,In_357,In_1515);
xor U3642 (N_3642,In_108,In_1366);
or U3643 (N_3643,In_193,In_608);
or U3644 (N_3644,In_1115,In_176);
or U3645 (N_3645,In_1008,In_1818);
nand U3646 (N_3646,In_58,In_1427);
or U3647 (N_3647,In_2791,In_2576);
nor U3648 (N_3648,In_2302,In_1572);
or U3649 (N_3649,In_1439,In_1097);
xnor U3650 (N_3650,In_1164,In_928);
nor U3651 (N_3651,In_1228,In_654);
and U3652 (N_3652,In_2479,In_2773);
nand U3653 (N_3653,In_696,In_1170);
xor U3654 (N_3654,In_1546,In_1629);
and U3655 (N_3655,In_1154,In_987);
or U3656 (N_3656,In_1535,In_2525);
xnor U3657 (N_3657,In_110,In_148);
and U3658 (N_3658,In_1986,In_1277);
nand U3659 (N_3659,In_1880,In_339);
xnor U3660 (N_3660,In_1752,In_1705);
or U3661 (N_3661,In_1301,In_693);
nor U3662 (N_3662,In_458,In_1137);
nand U3663 (N_3663,In_1265,In_594);
or U3664 (N_3664,In_2144,In_312);
nand U3665 (N_3665,In_306,In_1313);
nor U3666 (N_3666,In_2295,In_1672);
xnor U3667 (N_3667,In_1061,In_265);
and U3668 (N_3668,In_816,In_2059);
nor U3669 (N_3669,In_2532,In_197);
xor U3670 (N_3670,In_2138,In_2242);
xor U3671 (N_3671,In_460,In_1104);
nor U3672 (N_3672,In_2200,In_361);
or U3673 (N_3673,In_2598,In_954);
and U3674 (N_3674,In_2027,In_2264);
or U3675 (N_3675,In_1603,In_1504);
xnor U3676 (N_3676,In_1365,In_2417);
and U3677 (N_3677,In_2466,In_551);
nand U3678 (N_3678,In_2154,In_2258);
or U3679 (N_3679,In_2919,In_738);
and U3680 (N_3680,In_2519,In_1075);
nand U3681 (N_3681,In_1594,In_456);
nand U3682 (N_3682,In_18,In_2031);
nor U3683 (N_3683,In_1168,In_1274);
nand U3684 (N_3684,In_103,In_2174);
nand U3685 (N_3685,In_2230,In_2433);
xor U3686 (N_3686,In_1844,In_870);
nand U3687 (N_3687,In_1778,In_1319);
or U3688 (N_3688,In_1276,In_1535);
or U3689 (N_3689,In_546,In_1598);
or U3690 (N_3690,In_2884,In_1520);
xor U3691 (N_3691,In_2415,In_53);
xor U3692 (N_3692,In_568,In_2267);
xnor U3693 (N_3693,In_2329,In_2401);
or U3694 (N_3694,In_2910,In_1939);
nand U3695 (N_3695,In_2813,In_2570);
nand U3696 (N_3696,In_1602,In_2068);
nor U3697 (N_3697,In_2755,In_2870);
and U3698 (N_3698,In_1937,In_521);
nor U3699 (N_3699,In_1173,In_2769);
nor U3700 (N_3700,In_1406,In_2699);
nand U3701 (N_3701,In_281,In_2882);
xnor U3702 (N_3702,In_1335,In_2378);
xnor U3703 (N_3703,In_2066,In_1789);
nand U3704 (N_3704,In_375,In_1918);
or U3705 (N_3705,In_2814,In_1027);
xor U3706 (N_3706,In_580,In_2683);
nor U3707 (N_3707,In_1623,In_1351);
and U3708 (N_3708,In_1909,In_451);
xor U3709 (N_3709,In_1335,In_1150);
nor U3710 (N_3710,In_1684,In_308);
or U3711 (N_3711,In_885,In_1241);
xnor U3712 (N_3712,In_695,In_2489);
nor U3713 (N_3713,In_2455,In_93);
and U3714 (N_3714,In_1722,In_320);
or U3715 (N_3715,In_123,In_1566);
nor U3716 (N_3716,In_1918,In_392);
and U3717 (N_3717,In_2459,In_1678);
or U3718 (N_3718,In_1855,In_2426);
xnor U3719 (N_3719,In_1114,In_544);
xor U3720 (N_3720,In_1890,In_413);
nand U3721 (N_3721,In_2045,In_425);
and U3722 (N_3722,In_461,In_1456);
nand U3723 (N_3723,In_2085,In_2148);
or U3724 (N_3724,In_1144,In_258);
and U3725 (N_3725,In_1886,In_2828);
and U3726 (N_3726,In_1475,In_530);
nand U3727 (N_3727,In_628,In_2239);
xor U3728 (N_3728,In_1358,In_314);
nor U3729 (N_3729,In_141,In_345);
and U3730 (N_3730,In_1367,In_2533);
and U3731 (N_3731,In_2881,In_2965);
and U3732 (N_3732,In_2334,In_305);
xnor U3733 (N_3733,In_200,In_2262);
nand U3734 (N_3734,In_588,In_2744);
nor U3735 (N_3735,In_1509,In_2878);
and U3736 (N_3736,In_2860,In_2711);
and U3737 (N_3737,In_1973,In_265);
nand U3738 (N_3738,In_1848,In_1035);
nand U3739 (N_3739,In_294,In_2416);
or U3740 (N_3740,In_1919,In_2884);
xor U3741 (N_3741,In_810,In_1252);
xnor U3742 (N_3742,In_1480,In_2269);
xor U3743 (N_3743,In_1213,In_2193);
and U3744 (N_3744,In_89,In_153);
xor U3745 (N_3745,In_98,In_2424);
xor U3746 (N_3746,In_2257,In_2332);
xor U3747 (N_3747,In_2327,In_2235);
nand U3748 (N_3748,In_1550,In_2227);
or U3749 (N_3749,In_83,In_2104);
nor U3750 (N_3750,In_2223,In_1036);
nor U3751 (N_3751,In_618,In_168);
or U3752 (N_3752,In_1441,In_605);
xnor U3753 (N_3753,In_30,In_2135);
or U3754 (N_3754,In_2821,In_1985);
xor U3755 (N_3755,In_213,In_1646);
or U3756 (N_3756,In_2331,In_822);
xnor U3757 (N_3757,In_2128,In_720);
xnor U3758 (N_3758,In_1971,In_2978);
nand U3759 (N_3759,In_688,In_1426);
nand U3760 (N_3760,In_828,In_1000);
nor U3761 (N_3761,In_1755,In_1218);
or U3762 (N_3762,In_2777,In_1394);
or U3763 (N_3763,In_567,In_2700);
nand U3764 (N_3764,In_2252,In_1514);
and U3765 (N_3765,In_168,In_2343);
xor U3766 (N_3766,In_196,In_2697);
nand U3767 (N_3767,In_2656,In_2850);
nor U3768 (N_3768,In_410,In_115);
xnor U3769 (N_3769,In_807,In_2751);
nand U3770 (N_3770,In_854,In_703);
or U3771 (N_3771,In_2691,In_1254);
xnor U3772 (N_3772,In_1201,In_1189);
xnor U3773 (N_3773,In_2442,In_1585);
and U3774 (N_3774,In_1407,In_1515);
nand U3775 (N_3775,In_1602,In_2921);
or U3776 (N_3776,In_946,In_261);
nand U3777 (N_3777,In_2285,In_1194);
or U3778 (N_3778,In_30,In_1093);
and U3779 (N_3779,In_1081,In_2108);
nand U3780 (N_3780,In_2332,In_2295);
nand U3781 (N_3781,In_2299,In_109);
nor U3782 (N_3782,In_2569,In_140);
nor U3783 (N_3783,In_1700,In_1571);
xor U3784 (N_3784,In_2760,In_1128);
and U3785 (N_3785,In_1671,In_1295);
and U3786 (N_3786,In_2449,In_755);
and U3787 (N_3787,In_683,In_1940);
and U3788 (N_3788,In_1611,In_1596);
and U3789 (N_3789,In_2988,In_1286);
nor U3790 (N_3790,In_1321,In_933);
or U3791 (N_3791,In_776,In_965);
and U3792 (N_3792,In_1315,In_1336);
or U3793 (N_3793,In_20,In_1918);
nor U3794 (N_3794,In_154,In_1297);
nor U3795 (N_3795,In_1745,In_1100);
nor U3796 (N_3796,In_1307,In_1251);
xnor U3797 (N_3797,In_1118,In_2924);
nor U3798 (N_3798,In_2135,In_2081);
nor U3799 (N_3799,In_2062,In_363);
nor U3800 (N_3800,In_2200,In_2728);
nor U3801 (N_3801,In_1163,In_850);
nor U3802 (N_3802,In_1369,In_2845);
nand U3803 (N_3803,In_2295,In_2792);
xor U3804 (N_3804,In_2104,In_1954);
nor U3805 (N_3805,In_1622,In_1101);
nor U3806 (N_3806,In_1395,In_151);
or U3807 (N_3807,In_2285,In_2866);
or U3808 (N_3808,In_1980,In_2944);
xnor U3809 (N_3809,In_2026,In_266);
nand U3810 (N_3810,In_105,In_185);
nor U3811 (N_3811,In_1570,In_2212);
and U3812 (N_3812,In_2244,In_505);
nor U3813 (N_3813,In_2193,In_479);
and U3814 (N_3814,In_1790,In_307);
or U3815 (N_3815,In_805,In_872);
nand U3816 (N_3816,In_344,In_433);
or U3817 (N_3817,In_2318,In_357);
nor U3818 (N_3818,In_1858,In_2170);
nand U3819 (N_3819,In_1948,In_1841);
or U3820 (N_3820,In_2260,In_1826);
nor U3821 (N_3821,In_62,In_923);
or U3822 (N_3822,In_295,In_2780);
and U3823 (N_3823,In_102,In_2445);
and U3824 (N_3824,In_93,In_2247);
or U3825 (N_3825,In_1274,In_507);
or U3826 (N_3826,In_2761,In_2098);
xnor U3827 (N_3827,In_2399,In_2571);
and U3828 (N_3828,In_1006,In_2507);
and U3829 (N_3829,In_218,In_411);
and U3830 (N_3830,In_1175,In_21);
and U3831 (N_3831,In_1262,In_2320);
nand U3832 (N_3832,In_780,In_167);
xor U3833 (N_3833,In_857,In_101);
nor U3834 (N_3834,In_8,In_2090);
xor U3835 (N_3835,In_92,In_2768);
and U3836 (N_3836,In_2443,In_1785);
nand U3837 (N_3837,In_1835,In_2999);
or U3838 (N_3838,In_1824,In_1413);
xor U3839 (N_3839,In_1780,In_1494);
nor U3840 (N_3840,In_1338,In_1991);
and U3841 (N_3841,In_200,In_943);
and U3842 (N_3842,In_872,In_30);
nor U3843 (N_3843,In_85,In_2453);
and U3844 (N_3844,In_2917,In_92);
nor U3845 (N_3845,In_5,In_1121);
xor U3846 (N_3846,In_790,In_1630);
nand U3847 (N_3847,In_984,In_2948);
xnor U3848 (N_3848,In_1514,In_1135);
nand U3849 (N_3849,In_908,In_1367);
nor U3850 (N_3850,In_1563,In_1455);
nand U3851 (N_3851,In_1932,In_1327);
xnor U3852 (N_3852,In_1276,In_618);
nor U3853 (N_3853,In_275,In_2920);
nand U3854 (N_3854,In_880,In_271);
or U3855 (N_3855,In_1178,In_1890);
and U3856 (N_3856,In_771,In_481);
or U3857 (N_3857,In_2977,In_2350);
nand U3858 (N_3858,In_350,In_152);
and U3859 (N_3859,In_1501,In_1825);
or U3860 (N_3860,In_2591,In_1642);
xor U3861 (N_3861,In_895,In_258);
xor U3862 (N_3862,In_905,In_1805);
nand U3863 (N_3863,In_2526,In_327);
and U3864 (N_3864,In_1867,In_2816);
xnor U3865 (N_3865,In_2550,In_1598);
nor U3866 (N_3866,In_645,In_2832);
nand U3867 (N_3867,In_1444,In_1787);
or U3868 (N_3868,In_2089,In_420);
or U3869 (N_3869,In_1908,In_1500);
nor U3870 (N_3870,In_337,In_917);
or U3871 (N_3871,In_1377,In_2557);
xnor U3872 (N_3872,In_619,In_924);
nor U3873 (N_3873,In_259,In_2922);
nor U3874 (N_3874,In_285,In_2456);
or U3875 (N_3875,In_627,In_1465);
or U3876 (N_3876,In_2736,In_254);
nand U3877 (N_3877,In_2008,In_2186);
or U3878 (N_3878,In_450,In_2589);
or U3879 (N_3879,In_1745,In_2221);
or U3880 (N_3880,In_2264,In_932);
nor U3881 (N_3881,In_937,In_2174);
or U3882 (N_3882,In_1854,In_2698);
nor U3883 (N_3883,In_1551,In_260);
nor U3884 (N_3884,In_2058,In_2723);
nor U3885 (N_3885,In_951,In_166);
nor U3886 (N_3886,In_1474,In_1681);
xor U3887 (N_3887,In_2174,In_2518);
or U3888 (N_3888,In_870,In_1593);
xor U3889 (N_3889,In_2863,In_2684);
xor U3890 (N_3890,In_2821,In_2978);
xor U3891 (N_3891,In_2830,In_2994);
nand U3892 (N_3892,In_2189,In_87);
nand U3893 (N_3893,In_2919,In_2653);
xor U3894 (N_3894,In_2118,In_2247);
xor U3895 (N_3895,In_336,In_1402);
xor U3896 (N_3896,In_2288,In_520);
nor U3897 (N_3897,In_2712,In_209);
nand U3898 (N_3898,In_1598,In_1902);
nor U3899 (N_3899,In_1250,In_2298);
and U3900 (N_3900,In_915,In_2195);
and U3901 (N_3901,In_1232,In_2806);
nor U3902 (N_3902,In_1087,In_1250);
nor U3903 (N_3903,In_2475,In_2608);
or U3904 (N_3904,In_2551,In_2803);
nand U3905 (N_3905,In_360,In_2075);
or U3906 (N_3906,In_2024,In_2984);
nand U3907 (N_3907,In_1372,In_2099);
xor U3908 (N_3908,In_1090,In_1847);
xor U3909 (N_3909,In_2463,In_1378);
and U3910 (N_3910,In_1958,In_896);
or U3911 (N_3911,In_2737,In_931);
nor U3912 (N_3912,In_435,In_1835);
or U3913 (N_3913,In_1738,In_466);
nand U3914 (N_3914,In_2694,In_1359);
nor U3915 (N_3915,In_1169,In_1517);
xnor U3916 (N_3916,In_266,In_1452);
and U3917 (N_3917,In_32,In_2482);
nand U3918 (N_3918,In_568,In_639);
and U3919 (N_3919,In_302,In_86);
or U3920 (N_3920,In_2845,In_1038);
xnor U3921 (N_3921,In_2288,In_2592);
nor U3922 (N_3922,In_2189,In_800);
xor U3923 (N_3923,In_1691,In_501);
or U3924 (N_3924,In_891,In_1655);
xor U3925 (N_3925,In_116,In_2976);
and U3926 (N_3926,In_554,In_971);
nor U3927 (N_3927,In_528,In_1260);
xnor U3928 (N_3928,In_2716,In_1009);
or U3929 (N_3929,In_1935,In_586);
and U3930 (N_3930,In_2027,In_1270);
nand U3931 (N_3931,In_2880,In_1679);
nand U3932 (N_3932,In_768,In_1302);
or U3933 (N_3933,In_356,In_416);
nand U3934 (N_3934,In_324,In_2051);
nor U3935 (N_3935,In_256,In_1022);
nand U3936 (N_3936,In_2787,In_482);
and U3937 (N_3937,In_2654,In_859);
nor U3938 (N_3938,In_362,In_137);
nor U3939 (N_3939,In_2076,In_2095);
nor U3940 (N_3940,In_1723,In_2529);
or U3941 (N_3941,In_2081,In_756);
nor U3942 (N_3942,In_767,In_1863);
or U3943 (N_3943,In_649,In_1192);
xor U3944 (N_3944,In_1383,In_1540);
nor U3945 (N_3945,In_196,In_1284);
or U3946 (N_3946,In_1178,In_1487);
nand U3947 (N_3947,In_2828,In_1444);
and U3948 (N_3948,In_2281,In_2972);
nor U3949 (N_3949,In_260,In_498);
or U3950 (N_3950,In_1143,In_55);
or U3951 (N_3951,In_2190,In_934);
or U3952 (N_3952,In_1293,In_2828);
or U3953 (N_3953,In_1511,In_2572);
nand U3954 (N_3954,In_266,In_1632);
or U3955 (N_3955,In_954,In_1379);
nand U3956 (N_3956,In_1884,In_145);
or U3957 (N_3957,In_2694,In_1983);
xnor U3958 (N_3958,In_682,In_1601);
xor U3959 (N_3959,In_2359,In_825);
nor U3960 (N_3960,In_2712,In_1299);
nand U3961 (N_3961,In_39,In_1493);
and U3962 (N_3962,In_1391,In_1220);
nor U3963 (N_3963,In_1912,In_2644);
or U3964 (N_3964,In_1707,In_1875);
nand U3965 (N_3965,In_225,In_1697);
nand U3966 (N_3966,In_1473,In_788);
xor U3967 (N_3967,In_1749,In_996);
xor U3968 (N_3968,In_2851,In_1351);
nor U3969 (N_3969,In_1087,In_2292);
nor U3970 (N_3970,In_645,In_358);
xnor U3971 (N_3971,In_2136,In_931);
xnor U3972 (N_3972,In_2618,In_358);
and U3973 (N_3973,In_1088,In_2342);
and U3974 (N_3974,In_1191,In_752);
xnor U3975 (N_3975,In_504,In_2751);
nand U3976 (N_3976,In_2679,In_2963);
nor U3977 (N_3977,In_2611,In_1622);
and U3978 (N_3978,In_399,In_720);
and U3979 (N_3979,In_1158,In_170);
or U3980 (N_3980,In_1474,In_2914);
or U3981 (N_3981,In_87,In_2231);
and U3982 (N_3982,In_2732,In_1475);
nor U3983 (N_3983,In_2956,In_2546);
and U3984 (N_3984,In_2546,In_579);
xor U3985 (N_3985,In_2430,In_2240);
nand U3986 (N_3986,In_2112,In_967);
and U3987 (N_3987,In_231,In_1064);
nor U3988 (N_3988,In_533,In_744);
nor U3989 (N_3989,In_2230,In_570);
or U3990 (N_3990,In_1118,In_2094);
xor U3991 (N_3991,In_814,In_2511);
and U3992 (N_3992,In_42,In_147);
nor U3993 (N_3993,In_1825,In_2790);
nor U3994 (N_3994,In_933,In_1175);
and U3995 (N_3995,In_1843,In_2645);
nand U3996 (N_3996,In_2305,In_2527);
nor U3997 (N_3997,In_336,In_738);
or U3998 (N_3998,In_2539,In_2567);
and U3999 (N_3999,In_1351,In_2817);
nor U4000 (N_4000,In_1032,In_2754);
and U4001 (N_4001,In_1015,In_2413);
and U4002 (N_4002,In_2817,In_1148);
and U4003 (N_4003,In_1991,In_1697);
and U4004 (N_4004,In_2023,In_2881);
and U4005 (N_4005,In_1494,In_1104);
nand U4006 (N_4006,In_576,In_271);
and U4007 (N_4007,In_2741,In_2798);
xor U4008 (N_4008,In_320,In_2809);
or U4009 (N_4009,In_2451,In_1814);
xnor U4010 (N_4010,In_442,In_496);
xnor U4011 (N_4011,In_1958,In_593);
and U4012 (N_4012,In_319,In_2690);
nand U4013 (N_4013,In_2223,In_310);
and U4014 (N_4014,In_288,In_2156);
xor U4015 (N_4015,In_1528,In_2220);
nand U4016 (N_4016,In_2320,In_1846);
or U4017 (N_4017,In_1907,In_1720);
nand U4018 (N_4018,In_1061,In_2869);
xnor U4019 (N_4019,In_798,In_1841);
nand U4020 (N_4020,In_2172,In_2061);
nand U4021 (N_4021,In_2888,In_1902);
nand U4022 (N_4022,In_1682,In_1691);
xnor U4023 (N_4023,In_1249,In_677);
or U4024 (N_4024,In_1098,In_688);
nand U4025 (N_4025,In_1641,In_708);
xor U4026 (N_4026,In_2240,In_1699);
nor U4027 (N_4027,In_900,In_674);
and U4028 (N_4028,In_2674,In_2690);
or U4029 (N_4029,In_1938,In_2106);
and U4030 (N_4030,In_2883,In_1797);
and U4031 (N_4031,In_2845,In_2449);
nor U4032 (N_4032,In_2574,In_1693);
or U4033 (N_4033,In_1852,In_1776);
or U4034 (N_4034,In_402,In_1133);
or U4035 (N_4035,In_1732,In_483);
nor U4036 (N_4036,In_1262,In_504);
or U4037 (N_4037,In_2311,In_1105);
nand U4038 (N_4038,In_218,In_475);
nand U4039 (N_4039,In_2533,In_2850);
xnor U4040 (N_4040,In_437,In_417);
nand U4041 (N_4041,In_640,In_637);
or U4042 (N_4042,In_1068,In_1277);
nand U4043 (N_4043,In_287,In_1255);
xnor U4044 (N_4044,In_2373,In_945);
or U4045 (N_4045,In_1362,In_2125);
or U4046 (N_4046,In_449,In_318);
nor U4047 (N_4047,In_2824,In_2944);
xor U4048 (N_4048,In_1759,In_2477);
and U4049 (N_4049,In_1793,In_1730);
xor U4050 (N_4050,In_1066,In_2757);
nand U4051 (N_4051,In_217,In_779);
or U4052 (N_4052,In_1946,In_1421);
nor U4053 (N_4053,In_2543,In_1652);
nand U4054 (N_4054,In_2581,In_860);
xor U4055 (N_4055,In_1063,In_917);
and U4056 (N_4056,In_779,In_2794);
or U4057 (N_4057,In_624,In_1756);
xor U4058 (N_4058,In_1820,In_480);
and U4059 (N_4059,In_2019,In_2305);
nand U4060 (N_4060,In_1357,In_76);
nand U4061 (N_4061,In_2746,In_270);
nand U4062 (N_4062,In_2051,In_1329);
xor U4063 (N_4063,In_317,In_36);
and U4064 (N_4064,In_2176,In_1125);
nand U4065 (N_4065,In_661,In_1419);
nand U4066 (N_4066,In_145,In_2410);
nand U4067 (N_4067,In_1475,In_2137);
and U4068 (N_4068,In_483,In_479);
and U4069 (N_4069,In_931,In_1665);
and U4070 (N_4070,In_2879,In_1524);
xor U4071 (N_4071,In_201,In_44);
xor U4072 (N_4072,In_1785,In_1161);
nor U4073 (N_4073,In_2253,In_1748);
xnor U4074 (N_4074,In_2484,In_2739);
nand U4075 (N_4075,In_349,In_930);
or U4076 (N_4076,In_510,In_1445);
xnor U4077 (N_4077,In_2468,In_1546);
or U4078 (N_4078,In_592,In_1257);
xnor U4079 (N_4079,In_1003,In_714);
xor U4080 (N_4080,In_2696,In_2974);
nor U4081 (N_4081,In_1415,In_806);
nor U4082 (N_4082,In_2136,In_673);
nor U4083 (N_4083,In_1742,In_1668);
nand U4084 (N_4084,In_1781,In_2698);
and U4085 (N_4085,In_1901,In_1626);
xnor U4086 (N_4086,In_450,In_420);
nand U4087 (N_4087,In_512,In_1977);
xor U4088 (N_4088,In_946,In_684);
nand U4089 (N_4089,In_2434,In_1107);
or U4090 (N_4090,In_483,In_456);
xnor U4091 (N_4091,In_2105,In_129);
nor U4092 (N_4092,In_2002,In_2212);
or U4093 (N_4093,In_2271,In_2325);
nor U4094 (N_4094,In_908,In_1892);
and U4095 (N_4095,In_872,In_1056);
nor U4096 (N_4096,In_937,In_1939);
xnor U4097 (N_4097,In_241,In_497);
or U4098 (N_4098,In_1716,In_2616);
xor U4099 (N_4099,In_2857,In_1136);
nand U4100 (N_4100,In_431,In_1415);
or U4101 (N_4101,In_107,In_147);
nor U4102 (N_4102,In_473,In_856);
and U4103 (N_4103,In_92,In_275);
nor U4104 (N_4104,In_236,In_830);
or U4105 (N_4105,In_950,In_2337);
and U4106 (N_4106,In_849,In_1322);
or U4107 (N_4107,In_2379,In_305);
nor U4108 (N_4108,In_2663,In_2263);
nor U4109 (N_4109,In_772,In_753);
nand U4110 (N_4110,In_2971,In_2979);
nand U4111 (N_4111,In_838,In_2963);
xor U4112 (N_4112,In_2245,In_2960);
nand U4113 (N_4113,In_1403,In_1413);
and U4114 (N_4114,In_2120,In_50);
xnor U4115 (N_4115,In_1089,In_1444);
xnor U4116 (N_4116,In_659,In_609);
and U4117 (N_4117,In_526,In_1487);
or U4118 (N_4118,In_153,In_91);
or U4119 (N_4119,In_927,In_2735);
nor U4120 (N_4120,In_627,In_939);
xor U4121 (N_4121,In_2751,In_997);
nand U4122 (N_4122,In_1654,In_456);
nor U4123 (N_4123,In_2383,In_693);
or U4124 (N_4124,In_820,In_279);
xor U4125 (N_4125,In_2663,In_2610);
xor U4126 (N_4126,In_1337,In_404);
xor U4127 (N_4127,In_1616,In_2901);
nor U4128 (N_4128,In_2141,In_815);
xor U4129 (N_4129,In_1385,In_2737);
nor U4130 (N_4130,In_119,In_1507);
or U4131 (N_4131,In_755,In_320);
xnor U4132 (N_4132,In_594,In_1109);
xnor U4133 (N_4133,In_2806,In_2199);
xnor U4134 (N_4134,In_1282,In_2033);
and U4135 (N_4135,In_1471,In_1285);
or U4136 (N_4136,In_189,In_2310);
nor U4137 (N_4137,In_2623,In_640);
and U4138 (N_4138,In_841,In_756);
nand U4139 (N_4139,In_1566,In_2067);
and U4140 (N_4140,In_2426,In_445);
xor U4141 (N_4141,In_2022,In_2984);
nor U4142 (N_4142,In_516,In_1458);
and U4143 (N_4143,In_310,In_2518);
xnor U4144 (N_4144,In_2244,In_1457);
nand U4145 (N_4145,In_280,In_2494);
and U4146 (N_4146,In_1910,In_2080);
and U4147 (N_4147,In_279,In_790);
and U4148 (N_4148,In_2615,In_2649);
nor U4149 (N_4149,In_1984,In_242);
and U4150 (N_4150,In_2879,In_2610);
xnor U4151 (N_4151,In_809,In_551);
or U4152 (N_4152,In_1783,In_412);
or U4153 (N_4153,In_2886,In_1262);
or U4154 (N_4154,In_267,In_912);
nand U4155 (N_4155,In_658,In_1462);
nor U4156 (N_4156,In_1029,In_895);
xor U4157 (N_4157,In_2214,In_988);
and U4158 (N_4158,In_1051,In_200);
and U4159 (N_4159,In_1286,In_2311);
nand U4160 (N_4160,In_1201,In_1954);
nor U4161 (N_4161,In_2961,In_1905);
and U4162 (N_4162,In_542,In_241);
and U4163 (N_4163,In_1741,In_2432);
nor U4164 (N_4164,In_1910,In_2769);
xor U4165 (N_4165,In_1064,In_1608);
and U4166 (N_4166,In_2812,In_2113);
nand U4167 (N_4167,In_945,In_1225);
and U4168 (N_4168,In_294,In_2871);
nand U4169 (N_4169,In_1427,In_358);
and U4170 (N_4170,In_2388,In_574);
xnor U4171 (N_4171,In_101,In_1737);
nor U4172 (N_4172,In_70,In_2454);
xor U4173 (N_4173,In_2290,In_1272);
and U4174 (N_4174,In_1677,In_817);
nor U4175 (N_4175,In_915,In_2747);
nand U4176 (N_4176,In_839,In_2512);
nand U4177 (N_4177,In_219,In_1302);
nor U4178 (N_4178,In_1787,In_1799);
or U4179 (N_4179,In_2437,In_1262);
nand U4180 (N_4180,In_24,In_2439);
nor U4181 (N_4181,In_85,In_633);
xnor U4182 (N_4182,In_1052,In_2987);
and U4183 (N_4183,In_1698,In_65);
and U4184 (N_4184,In_2855,In_314);
and U4185 (N_4185,In_2505,In_1124);
nor U4186 (N_4186,In_1771,In_1665);
xor U4187 (N_4187,In_2229,In_322);
nand U4188 (N_4188,In_273,In_356);
or U4189 (N_4189,In_2482,In_2337);
and U4190 (N_4190,In_322,In_1974);
nor U4191 (N_4191,In_1129,In_2255);
nand U4192 (N_4192,In_1650,In_911);
nand U4193 (N_4193,In_57,In_2894);
and U4194 (N_4194,In_2323,In_1554);
nand U4195 (N_4195,In_219,In_2386);
xnor U4196 (N_4196,In_2554,In_2440);
xor U4197 (N_4197,In_531,In_1745);
xnor U4198 (N_4198,In_560,In_644);
nand U4199 (N_4199,In_1916,In_1111);
xnor U4200 (N_4200,In_2537,In_2856);
xnor U4201 (N_4201,In_2125,In_2299);
xnor U4202 (N_4202,In_2686,In_2753);
nand U4203 (N_4203,In_1978,In_1944);
and U4204 (N_4204,In_919,In_1347);
nand U4205 (N_4205,In_1365,In_1391);
xor U4206 (N_4206,In_2055,In_2761);
nor U4207 (N_4207,In_2525,In_2034);
and U4208 (N_4208,In_2538,In_1763);
or U4209 (N_4209,In_1649,In_312);
nand U4210 (N_4210,In_1624,In_274);
xor U4211 (N_4211,In_1498,In_1953);
nand U4212 (N_4212,In_2285,In_2877);
and U4213 (N_4213,In_1362,In_1116);
nand U4214 (N_4214,In_2096,In_105);
or U4215 (N_4215,In_403,In_2097);
nor U4216 (N_4216,In_632,In_1110);
xnor U4217 (N_4217,In_1738,In_747);
xor U4218 (N_4218,In_2742,In_1001);
xor U4219 (N_4219,In_2082,In_842);
nand U4220 (N_4220,In_2836,In_2066);
or U4221 (N_4221,In_2120,In_2677);
nand U4222 (N_4222,In_634,In_2805);
xnor U4223 (N_4223,In_2442,In_1386);
xor U4224 (N_4224,In_2606,In_464);
or U4225 (N_4225,In_2966,In_1741);
or U4226 (N_4226,In_1652,In_1076);
or U4227 (N_4227,In_2300,In_2324);
nor U4228 (N_4228,In_2524,In_2177);
nand U4229 (N_4229,In_2809,In_2833);
and U4230 (N_4230,In_1836,In_610);
nand U4231 (N_4231,In_1577,In_694);
nand U4232 (N_4232,In_2379,In_2953);
nor U4233 (N_4233,In_1138,In_2250);
nor U4234 (N_4234,In_341,In_2008);
nor U4235 (N_4235,In_1763,In_2055);
nor U4236 (N_4236,In_849,In_2892);
or U4237 (N_4237,In_587,In_1816);
xor U4238 (N_4238,In_1708,In_675);
nor U4239 (N_4239,In_462,In_1681);
nand U4240 (N_4240,In_441,In_2814);
or U4241 (N_4241,In_1356,In_818);
nor U4242 (N_4242,In_581,In_799);
nand U4243 (N_4243,In_2883,In_1472);
xor U4244 (N_4244,In_914,In_1893);
or U4245 (N_4245,In_2452,In_994);
or U4246 (N_4246,In_785,In_234);
and U4247 (N_4247,In_2967,In_899);
nand U4248 (N_4248,In_1424,In_2539);
xor U4249 (N_4249,In_833,In_674);
nor U4250 (N_4250,In_2966,In_2340);
or U4251 (N_4251,In_384,In_1206);
and U4252 (N_4252,In_692,In_2478);
nand U4253 (N_4253,In_2048,In_2558);
nand U4254 (N_4254,In_2891,In_1822);
nor U4255 (N_4255,In_1698,In_469);
xnor U4256 (N_4256,In_392,In_1586);
or U4257 (N_4257,In_2795,In_1369);
nor U4258 (N_4258,In_2196,In_2189);
nand U4259 (N_4259,In_2472,In_266);
or U4260 (N_4260,In_2159,In_2949);
nand U4261 (N_4261,In_1340,In_1960);
nor U4262 (N_4262,In_2610,In_722);
or U4263 (N_4263,In_250,In_2338);
and U4264 (N_4264,In_1606,In_1488);
or U4265 (N_4265,In_2495,In_2649);
nand U4266 (N_4266,In_2935,In_432);
or U4267 (N_4267,In_923,In_816);
nor U4268 (N_4268,In_2380,In_482);
xnor U4269 (N_4269,In_71,In_667);
nand U4270 (N_4270,In_2056,In_2638);
nor U4271 (N_4271,In_1405,In_2735);
nor U4272 (N_4272,In_2924,In_2431);
xor U4273 (N_4273,In_1799,In_2901);
nor U4274 (N_4274,In_330,In_344);
nor U4275 (N_4275,In_1904,In_2529);
and U4276 (N_4276,In_187,In_1862);
and U4277 (N_4277,In_1414,In_2633);
nand U4278 (N_4278,In_2374,In_1589);
xnor U4279 (N_4279,In_1322,In_502);
or U4280 (N_4280,In_1045,In_2043);
nor U4281 (N_4281,In_1132,In_2029);
or U4282 (N_4282,In_2957,In_2535);
or U4283 (N_4283,In_651,In_345);
nor U4284 (N_4284,In_2041,In_1224);
or U4285 (N_4285,In_670,In_2224);
or U4286 (N_4286,In_1909,In_253);
xnor U4287 (N_4287,In_948,In_2139);
and U4288 (N_4288,In_270,In_672);
nor U4289 (N_4289,In_623,In_1826);
nand U4290 (N_4290,In_616,In_2024);
and U4291 (N_4291,In_416,In_988);
nor U4292 (N_4292,In_2586,In_618);
xor U4293 (N_4293,In_2559,In_2437);
nor U4294 (N_4294,In_2352,In_1379);
xor U4295 (N_4295,In_1113,In_216);
nor U4296 (N_4296,In_1040,In_1351);
and U4297 (N_4297,In_1466,In_2633);
or U4298 (N_4298,In_2852,In_2846);
nor U4299 (N_4299,In_2292,In_93);
and U4300 (N_4300,In_1726,In_1282);
and U4301 (N_4301,In_2184,In_662);
or U4302 (N_4302,In_1736,In_2578);
and U4303 (N_4303,In_394,In_1830);
xor U4304 (N_4304,In_684,In_2453);
or U4305 (N_4305,In_809,In_1112);
nand U4306 (N_4306,In_1609,In_2397);
nand U4307 (N_4307,In_619,In_2567);
and U4308 (N_4308,In_1931,In_2286);
nor U4309 (N_4309,In_1467,In_1743);
nor U4310 (N_4310,In_113,In_900);
nand U4311 (N_4311,In_775,In_2747);
or U4312 (N_4312,In_355,In_318);
nand U4313 (N_4313,In_1003,In_1605);
and U4314 (N_4314,In_2996,In_267);
nor U4315 (N_4315,In_527,In_2032);
or U4316 (N_4316,In_987,In_1672);
and U4317 (N_4317,In_1606,In_2472);
or U4318 (N_4318,In_2734,In_266);
nor U4319 (N_4319,In_189,In_666);
nor U4320 (N_4320,In_781,In_1251);
or U4321 (N_4321,In_941,In_898);
nand U4322 (N_4322,In_2185,In_1678);
and U4323 (N_4323,In_2300,In_1755);
nand U4324 (N_4324,In_284,In_2962);
or U4325 (N_4325,In_1118,In_1778);
and U4326 (N_4326,In_2213,In_1242);
xnor U4327 (N_4327,In_291,In_2826);
or U4328 (N_4328,In_521,In_2893);
xnor U4329 (N_4329,In_1550,In_951);
xnor U4330 (N_4330,In_2093,In_265);
nor U4331 (N_4331,In_1833,In_491);
nor U4332 (N_4332,In_1790,In_1128);
nor U4333 (N_4333,In_2569,In_562);
nand U4334 (N_4334,In_1329,In_1510);
or U4335 (N_4335,In_1530,In_1957);
or U4336 (N_4336,In_1564,In_2509);
or U4337 (N_4337,In_921,In_668);
nor U4338 (N_4338,In_82,In_904);
or U4339 (N_4339,In_695,In_2638);
or U4340 (N_4340,In_1621,In_693);
nor U4341 (N_4341,In_326,In_2268);
nor U4342 (N_4342,In_272,In_2049);
nand U4343 (N_4343,In_1626,In_1121);
nand U4344 (N_4344,In_573,In_1741);
nand U4345 (N_4345,In_1550,In_2812);
and U4346 (N_4346,In_1799,In_1247);
xnor U4347 (N_4347,In_1376,In_77);
nand U4348 (N_4348,In_2086,In_1651);
xnor U4349 (N_4349,In_1920,In_1252);
and U4350 (N_4350,In_1906,In_1175);
or U4351 (N_4351,In_1561,In_219);
nor U4352 (N_4352,In_25,In_2399);
nor U4353 (N_4353,In_373,In_140);
nor U4354 (N_4354,In_2100,In_467);
nand U4355 (N_4355,In_2652,In_1800);
xor U4356 (N_4356,In_1816,In_211);
nand U4357 (N_4357,In_2785,In_1151);
nor U4358 (N_4358,In_2876,In_1245);
nor U4359 (N_4359,In_1477,In_2725);
or U4360 (N_4360,In_2107,In_1614);
xnor U4361 (N_4361,In_998,In_1921);
nand U4362 (N_4362,In_129,In_1486);
nor U4363 (N_4363,In_184,In_732);
and U4364 (N_4364,In_1886,In_2709);
nor U4365 (N_4365,In_2557,In_1154);
nor U4366 (N_4366,In_923,In_2510);
xnor U4367 (N_4367,In_1488,In_1162);
nor U4368 (N_4368,In_910,In_250);
nor U4369 (N_4369,In_51,In_1761);
nor U4370 (N_4370,In_1422,In_1793);
xnor U4371 (N_4371,In_885,In_712);
nand U4372 (N_4372,In_837,In_2728);
nand U4373 (N_4373,In_653,In_768);
nor U4374 (N_4374,In_2295,In_2320);
or U4375 (N_4375,In_2838,In_2618);
xor U4376 (N_4376,In_835,In_49);
xor U4377 (N_4377,In_1029,In_298);
nand U4378 (N_4378,In_2330,In_1469);
nor U4379 (N_4379,In_1241,In_1755);
nor U4380 (N_4380,In_1159,In_1933);
nor U4381 (N_4381,In_1565,In_2396);
nand U4382 (N_4382,In_612,In_1072);
and U4383 (N_4383,In_513,In_1276);
xor U4384 (N_4384,In_69,In_2718);
xor U4385 (N_4385,In_1382,In_1526);
or U4386 (N_4386,In_2143,In_863);
xor U4387 (N_4387,In_2344,In_1262);
and U4388 (N_4388,In_617,In_545);
nand U4389 (N_4389,In_1969,In_182);
or U4390 (N_4390,In_2288,In_2193);
and U4391 (N_4391,In_1455,In_1971);
and U4392 (N_4392,In_2884,In_2507);
or U4393 (N_4393,In_702,In_2029);
and U4394 (N_4394,In_2427,In_2713);
and U4395 (N_4395,In_1967,In_1673);
xor U4396 (N_4396,In_268,In_2825);
nor U4397 (N_4397,In_271,In_396);
xor U4398 (N_4398,In_1010,In_92);
xnor U4399 (N_4399,In_1022,In_895);
nor U4400 (N_4400,In_1928,In_1548);
nand U4401 (N_4401,In_353,In_2439);
or U4402 (N_4402,In_1504,In_312);
nor U4403 (N_4403,In_785,In_755);
nand U4404 (N_4404,In_334,In_2189);
and U4405 (N_4405,In_171,In_381);
nor U4406 (N_4406,In_1848,In_2608);
nor U4407 (N_4407,In_1402,In_1331);
nand U4408 (N_4408,In_2037,In_1884);
and U4409 (N_4409,In_492,In_2159);
xor U4410 (N_4410,In_1965,In_657);
nor U4411 (N_4411,In_2463,In_1252);
xor U4412 (N_4412,In_2959,In_2212);
nand U4413 (N_4413,In_2732,In_1602);
or U4414 (N_4414,In_230,In_285);
and U4415 (N_4415,In_1076,In_472);
or U4416 (N_4416,In_1158,In_2430);
nor U4417 (N_4417,In_2426,In_1306);
and U4418 (N_4418,In_2058,In_1671);
or U4419 (N_4419,In_1986,In_1006);
or U4420 (N_4420,In_419,In_1886);
and U4421 (N_4421,In_1054,In_1278);
xor U4422 (N_4422,In_94,In_1049);
and U4423 (N_4423,In_2693,In_343);
xnor U4424 (N_4424,In_916,In_1885);
xor U4425 (N_4425,In_352,In_2951);
nand U4426 (N_4426,In_1479,In_1439);
nor U4427 (N_4427,In_2372,In_2115);
nand U4428 (N_4428,In_1735,In_2718);
nand U4429 (N_4429,In_479,In_1689);
nand U4430 (N_4430,In_2377,In_1045);
or U4431 (N_4431,In_130,In_1974);
nand U4432 (N_4432,In_60,In_1349);
nand U4433 (N_4433,In_2241,In_31);
and U4434 (N_4434,In_817,In_2199);
xnor U4435 (N_4435,In_2146,In_1718);
and U4436 (N_4436,In_1664,In_675);
xnor U4437 (N_4437,In_1758,In_2041);
xnor U4438 (N_4438,In_1592,In_1393);
and U4439 (N_4439,In_1426,In_1589);
nand U4440 (N_4440,In_2228,In_1067);
and U4441 (N_4441,In_2391,In_1966);
nor U4442 (N_4442,In_1329,In_264);
nor U4443 (N_4443,In_801,In_2970);
or U4444 (N_4444,In_2001,In_624);
or U4445 (N_4445,In_2,In_996);
and U4446 (N_4446,In_1749,In_1249);
nor U4447 (N_4447,In_1223,In_1103);
and U4448 (N_4448,In_995,In_990);
xnor U4449 (N_4449,In_562,In_907);
nor U4450 (N_4450,In_2488,In_2097);
nor U4451 (N_4451,In_1286,In_2604);
or U4452 (N_4452,In_1678,In_2542);
and U4453 (N_4453,In_1428,In_202);
and U4454 (N_4454,In_1937,In_566);
or U4455 (N_4455,In_1243,In_452);
nor U4456 (N_4456,In_1919,In_2749);
and U4457 (N_4457,In_2785,In_72);
nand U4458 (N_4458,In_984,In_737);
or U4459 (N_4459,In_195,In_230);
nand U4460 (N_4460,In_1061,In_2813);
nor U4461 (N_4461,In_1006,In_488);
and U4462 (N_4462,In_719,In_1534);
nand U4463 (N_4463,In_1544,In_1701);
nor U4464 (N_4464,In_2593,In_272);
xnor U4465 (N_4465,In_2172,In_1206);
xnor U4466 (N_4466,In_189,In_2515);
nand U4467 (N_4467,In_113,In_2802);
xnor U4468 (N_4468,In_363,In_1327);
nand U4469 (N_4469,In_19,In_1169);
nand U4470 (N_4470,In_1510,In_2069);
and U4471 (N_4471,In_1375,In_1184);
and U4472 (N_4472,In_1413,In_630);
or U4473 (N_4473,In_62,In_415);
nand U4474 (N_4474,In_2863,In_2642);
or U4475 (N_4475,In_1478,In_2759);
and U4476 (N_4476,In_1228,In_2101);
nand U4477 (N_4477,In_2971,In_2640);
and U4478 (N_4478,In_2135,In_257);
nand U4479 (N_4479,In_982,In_910);
and U4480 (N_4480,In_1554,In_2746);
nand U4481 (N_4481,In_1008,In_2515);
xnor U4482 (N_4482,In_2296,In_1487);
and U4483 (N_4483,In_1874,In_1253);
nor U4484 (N_4484,In_2119,In_2614);
nor U4485 (N_4485,In_1039,In_1368);
nor U4486 (N_4486,In_256,In_1005);
nor U4487 (N_4487,In_1210,In_2275);
xnor U4488 (N_4488,In_2232,In_1071);
and U4489 (N_4489,In_58,In_2405);
or U4490 (N_4490,In_2135,In_1090);
and U4491 (N_4491,In_2810,In_267);
and U4492 (N_4492,In_2902,In_93);
xnor U4493 (N_4493,In_934,In_1558);
nor U4494 (N_4494,In_51,In_358);
or U4495 (N_4495,In_1597,In_2910);
or U4496 (N_4496,In_2627,In_1);
or U4497 (N_4497,In_1537,In_461);
nor U4498 (N_4498,In_695,In_554);
nand U4499 (N_4499,In_2342,In_2257);
or U4500 (N_4500,In_2917,In_1557);
xor U4501 (N_4501,In_627,In_2824);
or U4502 (N_4502,In_2392,In_2879);
nor U4503 (N_4503,In_1015,In_705);
or U4504 (N_4504,In_1899,In_2513);
xor U4505 (N_4505,In_1720,In_243);
nand U4506 (N_4506,In_1946,In_1119);
or U4507 (N_4507,In_1009,In_582);
and U4508 (N_4508,In_365,In_302);
nand U4509 (N_4509,In_1526,In_920);
nor U4510 (N_4510,In_528,In_1379);
or U4511 (N_4511,In_2676,In_1345);
or U4512 (N_4512,In_2031,In_1455);
and U4513 (N_4513,In_1047,In_2509);
xor U4514 (N_4514,In_1623,In_2646);
or U4515 (N_4515,In_2473,In_2635);
and U4516 (N_4516,In_1537,In_2388);
xor U4517 (N_4517,In_2907,In_124);
or U4518 (N_4518,In_890,In_499);
and U4519 (N_4519,In_1788,In_1981);
nand U4520 (N_4520,In_1719,In_253);
or U4521 (N_4521,In_1580,In_1937);
and U4522 (N_4522,In_1787,In_1296);
nor U4523 (N_4523,In_875,In_1056);
nand U4524 (N_4524,In_2878,In_1534);
xnor U4525 (N_4525,In_2635,In_755);
nor U4526 (N_4526,In_510,In_1063);
xnor U4527 (N_4527,In_1880,In_512);
xnor U4528 (N_4528,In_2234,In_397);
and U4529 (N_4529,In_712,In_1682);
or U4530 (N_4530,In_1962,In_2767);
and U4531 (N_4531,In_2167,In_1998);
and U4532 (N_4532,In_1702,In_2520);
nor U4533 (N_4533,In_1447,In_912);
xnor U4534 (N_4534,In_118,In_627);
or U4535 (N_4535,In_1415,In_1547);
or U4536 (N_4536,In_1576,In_1572);
nor U4537 (N_4537,In_1751,In_2635);
xor U4538 (N_4538,In_1654,In_274);
xnor U4539 (N_4539,In_17,In_2082);
and U4540 (N_4540,In_915,In_1613);
or U4541 (N_4541,In_263,In_1994);
xor U4542 (N_4542,In_2904,In_1812);
xnor U4543 (N_4543,In_2136,In_310);
and U4544 (N_4544,In_2941,In_2748);
and U4545 (N_4545,In_468,In_1747);
or U4546 (N_4546,In_672,In_1035);
or U4547 (N_4547,In_1312,In_579);
nor U4548 (N_4548,In_1113,In_2421);
xnor U4549 (N_4549,In_2311,In_2520);
nor U4550 (N_4550,In_1270,In_751);
nand U4551 (N_4551,In_1555,In_2591);
nor U4552 (N_4552,In_978,In_351);
nand U4553 (N_4553,In_2885,In_911);
xnor U4554 (N_4554,In_773,In_1165);
nand U4555 (N_4555,In_1708,In_2424);
xnor U4556 (N_4556,In_2001,In_1874);
or U4557 (N_4557,In_984,In_1042);
and U4558 (N_4558,In_661,In_2626);
nand U4559 (N_4559,In_1217,In_1382);
and U4560 (N_4560,In_2214,In_1392);
nand U4561 (N_4561,In_265,In_1025);
xor U4562 (N_4562,In_1317,In_1610);
or U4563 (N_4563,In_1448,In_461);
nor U4564 (N_4564,In_1623,In_2211);
xnor U4565 (N_4565,In_720,In_2823);
or U4566 (N_4566,In_539,In_2706);
or U4567 (N_4567,In_996,In_1295);
nand U4568 (N_4568,In_2938,In_284);
xnor U4569 (N_4569,In_1764,In_2230);
nor U4570 (N_4570,In_2565,In_2855);
nor U4571 (N_4571,In_2722,In_219);
xor U4572 (N_4572,In_366,In_2342);
and U4573 (N_4573,In_2300,In_2205);
or U4574 (N_4574,In_1385,In_131);
and U4575 (N_4575,In_1504,In_387);
or U4576 (N_4576,In_680,In_132);
or U4577 (N_4577,In_2199,In_394);
or U4578 (N_4578,In_1476,In_1976);
or U4579 (N_4579,In_1596,In_667);
or U4580 (N_4580,In_2628,In_2537);
nand U4581 (N_4581,In_1627,In_2280);
nand U4582 (N_4582,In_330,In_2505);
or U4583 (N_4583,In_1723,In_737);
nand U4584 (N_4584,In_2396,In_2100);
nand U4585 (N_4585,In_1726,In_1732);
and U4586 (N_4586,In_2263,In_2559);
nor U4587 (N_4587,In_58,In_1615);
nor U4588 (N_4588,In_1942,In_41);
xnor U4589 (N_4589,In_1032,In_2430);
xnor U4590 (N_4590,In_1886,In_261);
nand U4591 (N_4591,In_415,In_223);
nor U4592 (N_4592,In_941,In_146);
nand U4593 (N_4593,In_1234,In_2836);
or U4594 (N_4594,In_1080,In_1674);
nand U4595 (N_4595,In_1351,In_685);
xnor U4596 (N_4596,In_2344,In_1044);
nand U4597 (N_4597,In_2737,In_2929);
xor U4598 (N_4598,In_233,In_2269);
or U4599 (N_4599,In_1015,In_866);
nor U4600 (N_4600,In_827,In_58);
nor U4601 (N_4601,In_203,In_1769);
nand U4602 (N_4602,In_1306,In_2930);
nand U4603 (N_4603,In_1483,In_2282);
or U4604 (N_4604,In_180,In_2144);
and U4605 (N_4605,In_1463,In_416);
nand U4606 (N_4606,In_1080,In_1935);
xor U4607 (N_4607,In_842,In_2198);
and U4608 (N_4608,In_234,In_2211);
xor U4609 (N_4609,In_1619,In_2113);
nand U4610 (N_4610,In_793,In_474);
or U4611 (N_4611,In_697,In_2519);
or U4612 (N_4612,In_501,In_2047);
and U4613 (N_4613,In_2402,In_2706);
nand U4614 (N_4614,In_1833,In_617);
or U4615 (N_4615,In_2775,In_911);
nor U4616 (N_4616,In_977,In_673);
nor U4617 (N_4617,In_171,In_1227);
xnor U4618 (N_4618,In_2056,In_2716);
and U4619 (N_4619,In_1010,In_1657);
xnor U4620 (N_4620,In_2276,In_1539);
nand U4621 (N_4621,In_2996,In_1027);
or U4622 (N_4622,In_977,In_1309);
nand U4623 (N_4623,In_2517,In_1081);
or U4624 (N_4624,In_5,In_573);
and U4625 (N_4625,In_2768,In_2884);
nor U4626 (N_4626,In_2804,In_1870);
nor U4627 (N_4627,In_2342,In_1071);
or U4628 (N_4628,In_1710,In_1071);
and U4629 (N_4629,In_2794,In_449);
xor U4630 (N_4630,In_1931,In_1132);
xnor U4631 (N_4631,In_244,In_1287);
and U4632 (N_4632,In_2735,In_2032);
xor U4633 (N_4633,In_2302,In_631);
xnor U4634 (N_4634,In_631,In_326);
or U4635 (N_4635,In_608,In_2145);
or U4636 (N_4636,In_1091,In_917);
nor U4637 (N_4637,In_1501,In_502);
xnor U4638 (N_4638,In_2334,In_1890);
and U4639 (N_4639,In_2278,In_2727);
xor U4640 (N_4640,In_1012,In_2071);
xnor U4641 (N_4641,In_2067,In_5);
nand U4642 (N_4642,In_2309,In_1743);
or U4643 (N_4643,In_542,In_408);
and U4644 (N_4644,In_1144,In_77);
xor U4645 (N_4645,In_39,In_971);
or U4646 (N_4646,In_1521,In_1229);
nor U4647 (N_4647,In_2394,In_2371);
nand U4648 (N_4648,In_2279,In_2330);
nand U4649 (N_4649,In_1926,In_2848);
nor U4650 (N_4650,In_733,In_1758);
nand U4651 (N_4651,In_922,In_87);
nand U4652 (N_4652,In_2647,In_747);
and U4653 (N_4653,In_1857,In_96);
nor U4654 (N_4654,In_2750,In_115);
xor U4655 (N_4655,In_2389,In_2724);
nand U4656 (N_4656,In_187,In_1478);
and U4657 (N_4657,In_822,In_1267);
and U4658 (N_4658,In_941,In_2086);
xor U4659 (N_4659,In_769,In_2272);
nor U4660 (N_4660,In_2787,In_368);
xnor U4661 (N_4661,In_324,In_315);
or U4662 (N_4662,In_1753,In_1005);
nor U4663 (N_4663,In_900,In_1598);
and U4664 (N_4664,In_217,In_2735);
nor U4665 (N_4665,In_774,In_2657);
nor U4666 (N_4666,In_1920,In_405);
nand U4667 (N_4667,In_1873,In_840);
and U4668 (N_4668,In_967,In_1357);
xor U4669 (N_4669,In_2882,In_2301);
or U4670 (N_4670,In_1895,In_1318);
nor U4671 (N_4671,In_1224,In_1795);
nand U4672 (N_4672,In_1970,In_2515);
nand U4673 (N_4673,In_2903,In_506);
nor U4674 (N_4674,In_1361,In_2944);
or U4675 (N_4675,In_2052,In_759);
xor U4676 (N_4676,In_1208,In_2189);
nand U4677 (N_4677,In_2024,In_1834);
and U4678 (N_4678,In_1905,In_197);
nor U4679 (N_4679,In_1131,In_1962);
or U4680 (N_4680,In_437,In_706);
xnor U4681 (N_4681,In_252,In_1967);
nand U4682 (N_4682,In_2834,In_75);
xnor U4683 (N_4683,In_583,In_2742);
nor U4684 (N_4684,In_428,In_941);
xor U4685 (N_4685,In_192,In_828);
or U4686 (N_4686,In_1036,In_598);
nor U4687 (N_4687,In_1454,In_434);
nor U4688 (N_4688,In_1165,In_2874);
or U4689 (N_4689,In_1490,In_2680);
nand U4690 (N_4690,In_2790,In_793);
xnor U4691 (N_4691,In_1167,In_1243);
nand U4692 (N_4692,In_2814,In_2491);
and U4693 (N_4693,In_746,In_1790);
and U4694 (N_4694,In_2157,In_1985);
nor U4695 (N_4695,In_2531,In_2972);
and U4696 (N_4696,In_876,In_1994);
nand U4697 (N_4697,In_1913,In_2684);
xor U4698 (N_4698,In_250,In_2928);
nand U4699 (N_4699,In_1973,In_696);
xnor U4700 (N_4700,In_1499,In_2704);
xor U4701 (N_4701,In_2625,In_1964);
nor U4702 (N_4702,In_1334,In_2119);
and U4703 (N_4703,In_2946,In_1775);
nand U4704 (N_4704,In_2681,In_2771);
and U4705 (N_4705,In_1815,In_937);
nor U4706 (N_4706,In_269,In_406);
or U4707 (N_4707,In_1318,In_2117);
nand U4708 (N_4708,In_2241,In_84);
or U4709 (N_4709,In_1486,In_282);
nand U4710 (N_4710,In_2697,In_829);
or U4711 (N_4711,In_670,In_2495);
nor U4712 (N_4712,In_2276,In_2752);
and U4713 (N_4713,In_887,In_1033);
and U4714 (N_4714,In_2403,In_635);
nand U4715 (N_4715,In_513,In_2369);
nor U4716 (N_4716,In_657,In_1739);
nor U4717 (N_4717,In_782,In_668);
and U4718 (N_4718,In_2879,In_1510);
or U4719 (N_4719,In_1581,In_81);
xor U4720 (N_4720,In_1822,In_1290);
nor U4721 (N_4721,In_2864,In_2057);
or U4722 (N_4722,In_635,In_81);
or U4723 (N_4723,In_2434,In_2775);
nand U4724 (N_4724,In_1485,In_1673);
xnor U4725 (N_4725,In_469,In_203);
and U4726 (N_4726,In_1184,In_2126);
nor U4727 (N_4727,In_2350,In_2393);
or U4728 (N_4728,In_2215,In_171);
and U4729 (N_4729,In_2854,In_1957);
nand U4730 (N_4730,In_224,In_2505);
or U4731 (N_4731,In_1758,In_792);
or U4732 (N_4732,In_2534,In_1191);
nand U4733 (N_4733,In_2149,In_2015);
nand U4734 (N_4734,In_2052,In_2278);
xor U4735 (N_4735,In_544,In_2184);
nor U4736 (N_4736,In_2302,In_1534);
xor U4737 (N_4737,In_2773,In_2386);
or U4738 (N_4738,In_215,In_885);
or U4739 (N_4739,In_1668,In_2589);
nor U4740 (N_4740,In_194,In_840);
nor U4741 (N_4741,In_2194,In_1876);
or U4742 (N_4742,In_2396,In_1514);
nand U4743 (N_4743,In_935,In_259);
or U4744 (N_4744,In_1244,In_982);
and U4745 (N_4745,In_2679,In_529);
and U4746 (N_4746,In_443,In_577);
or U4747 (N_4747,In_1736,In_208);
nand U4748 (N_4748,In_1652,In_351);
nand U4749 (N_4749,In_2546,In_1561);
or U4750 (N_4750,In_1817,In_8);
and U4751 (N_4751,In_1481,In_718);
nor U4752 (N_4752,In_2289,In_1613);
nand U4753 (N_4753,In_2495,In_1582);
nor U4754 (N_4754,In_1728,In_239);
nand U4755 (N_4755,In_166,In_1640);
and U4756 (N_4756,In_1273,In_2935);
xor U4757 (N_4757,In_1546,In_1152);
xor U4758 (N_4758,In_1265,In_1650);
xnor U4759 (N_4759,In_2579,In_2790);
and U4760 (N_4760,In_1053,In_1583);
or U4761 (N_4761,In_2753,In_769);
nor U4762 (N_4762,In_570,In_732);
and U4763 (N_4763,In_1068,In_2285);
nand U4764 (N_4764,In_2514,In_2961);
nand U4765 (N_4765,In_877,In_1814);
or U4766 (N_4766,In_1897,In_2542);
xor U4767 (N_4767,In_430,In_2265);
and U4768 (N_4768,In_1859,In_2555);
nand U4769 (N_4769,In_2780,In_304);
xor U4770 (N_4770,In_1309,In_1781);
and U4771 (N_4771,In_2388,In_1597);
or U4772 (N_4772,In_1200,In_586);
nor U4773 (N_4773,In_2400,In_114);
and U4774 (N_4774,In_2119,In_756);
nor U4775 (N_4775,In_2992,In_288);
nor U4776 (N_4776,In_2916,In_1675);
nand U4777 (N_4777,In_865,In_491);
nand U4778 (N_4778,In_192,In_2148);
xor U4779 (N_4779,In_1631,In_335);
nand U4780 (N_4780,In_2944,In_400);
nand U4781 (N_4781,In_1577,In_1922);
and U4782 (N_4782,In_907,In_385);
xnor U4783 (N_4783,In_2615,In_2260);
nand U4784 (N_4784,In_784,In_1000);
xnor U4785 (N_4785,In_2522,In_927);
xnor U4786 (N_4786,In_1681,In_973);
or U4787 (N_4787,In_35,In_636);
xor U4788 (N_4788,In_2311,In_1677);
nor U4789 (N_4789,In_2633,In_764);
nand U4790 (N_4790,In_1216,In_2128);
nand U4791 (N_4791,In_1671,In_2914);
nand U4792 (N_4792,In_2864,In_200);
and U4793 (N_4793,In_1598,In_461);
nor U4794 (N_4794,In_268,In_1695);
xor U4795 (N_4795,In_572,In_1747);
xnor U4796 (N_4796,In_321,In_1939);
nor U4797 (N_4797,In_1562,In_33);
and U4798 (N_4798,In_549,In_2581);
nor U4799 (N_4799,In_927,In_1401);
nand U4800 (N_4800,In_145,In_1477);
xnor U4801 (N_4801,In_2116,In_345);
xor U4802 (N_4802,In_600,In_1847);
nand U4803 (N_4803,In_1505,In_1430);
xor U4804 (N_4804,In_321,In_1351);
nor U4805 (N_4805,In_1779,In_1045);
or U4806 (N_4806,In_2210,In_554);
or U4807 (N_4807,In_580,In_2797);
and U4808 (N_4808,In_1090,In_659);
or U4809 (N_4809,In_938,In_1190);
and U4810 (N_4810,In_1809,In_103);
xnor U4811 (N_4811,In_699,In_449);
xor U4812 (N_4812,In_2362,In_2891);
or U4813 (N_4813,In_1132,In_456);
or U4814 (N_4814,In_576,In_1130);
and U4815 (N_4815,In_2542,In_1528);
xnor U4816 (N_4816,In_2161,In_1445);
nor U4817 (N_4817,In_421,In_2729);
nor U4818 (N_4818,In_773,In_305);
and U4819 (N_4819,In_2026,In_820);
xnor U4820 (N_4820,In_654,In_2934);
nor U4821 (N_4821,In_2131,In_1779);
nor U4822 (N_4822,In_2497,In_222);
or U4823 (N_4823,In_393,In_658);
nand U4824 (N_4824,In_1270,In_2989);
nor U4825 (N_4825,In_2593,In_91);
or U4826 (N_4826,In_1498,In_568);
nor U4827 (N_4827,In_1523,In_383);
and U4828 (N_4828,In_54,In_447);
or U4829 (N_4829,In_1928,In_1066);
xor U4830 (N_4830,In_902,In_2457);
nor U4831 (N_4831,In_2871,In_2075);
nand U4832 (N_4832,In_367,In_1906);
or U4833 (N_4833,In_1013,In_1152);
nor U4834 (N_4834,In_2701,In_1554);
nand U4835 (N_4835,In_2082,In_2267);
or U4836 (N_4836,In_2825,In_642);
nor U4837 (N_4837,In_154,In_1608);
nand U4838 (N_4838,In_161,In_109);
xor U4839 (N_4839,In_760,In_738);
xor U4840 (N_4840,In_423,In_503);
nand U4841 (N_4841,In_1311,In_2908);
and U4842 (N_4842,In_1502,In_2405);
nor U4843 (N_4843,In_1951,In_2807);
nand U4844 (N_4844,In_2203,In_258);
nand U4845 (N_4845,In_890,In_1872);
nor U4846 (N_4846,In_1455,In_1189);
nand U4847 (N_4847,In_733,In_2331);
nor U4848 (N_4848,In_1371,In_2641);
nand U4849 (N_4849,In_131,In_1754);
nand U4850 (N_4850,In_1639,In_1550);
nand U4851 (N_4851,In_2911,In_47);
xnor U4852 (N_4852,In_2675,In_1002);
nor U4853 (N_4853,In_1789,In_1808);
nand U4854 (N_4854,In_1889,In_1787);
nor U4855 (N_4855,In_2019,In_2120);
nand U4856 (N_4856,In_1543,In_1574);
nor U4857 (N_4857,In_2850,In_2160);
and U4858 (N_4858,In_546,In_2012);
xor U4859 (N_4859,In_1981,In_1717);
nor U4860 (N_4860,In_2441,In_2980);
nand U4861 (N_4861,In_1656,In_2791);
and U4862 (N_4862,In_1195,In_112);
or U4863 (N_4863,In_271,In_113);
or U4864 (N_4864,In_33,In_1892);
nor U4865 (N_4865,In_1795,In_2029);
xor U4866 (N_4866,In_169,In_486);
or U4867 (N_4867,In_1870,In_2698);
or U4868 (N_4868,In_1741,In_1163);
and U4869 (N_4869,In_656,In_1481);
or U4870 (N_4870,In_1349,In_2633);
nand U4871 (N_4871,In_1519,In_2261);
nor U4872 (N_4872,In_2693,In_1111);
nand U4873 (N_4873,In_1468,In_733);
or U4874 (N_4874,In_1763,In_1505);
nor U4875 (N_4875,In_2640,In_2059);
nand U4876 (N_4876,In_384,In_142);
and U4877 (N_4877,In_1623,In_1410);
xor U4878 (N_4878,In_879,In_1593);
or U4879 (N_4879,In_1765,In_362);
nor U4880 (N_4880,In_2030,In_2965);
or U4881 (N_4881,In_1501,In_210);
nand U4882 (N_4882,In_750,In_1133);
xor U4883 (N_4883,In_2864,In_1449);
nor U4884 (N_4884,In_350,In_2206);
or U4885 (N_4885,In_2604,In_1493);
xnor U4886 (N_4886,In_2650,In_672);
xor U4887 (N_4887,In_1182,In_470);
and U4888 (N_4888,In_1722,In_1858);
and U4889 (N_4889,In_1695,In_200);
nor U4890 (N_4890,In_2012,In_1212);
or U4891 (N_4891,In_2640,In_1553);
nand U4892 (N_4892,In_430,In_2635);
xor U4893 (N_4893,In_947,In_1742);
or U4894 (N_4894,In_2570,In_1202);
nand U4895 (N_4895,In_960,In_1481);
xor U4896 (N_4896,In_336,In_1978);
xor U4897 (N_4897,In_1909,In_1012);
and U4898 (N_4898,In_2841,In_930);
nand U4899 (N_4899,In_1044,In_2226);
and U4900 (N_4900,In_986,In_1459);
and U4901 (N_4901,In_2711,In_2654);
and U4902 (N_4902,In_2481,In_1739);
or U4903 (N_4903,In_2124,In_1823);
nand U4904 (N_4904,In_2478,In_1831);
xnor U4905 (N_4905,In_42,In_1446);
nor U4906 (N_4906,In_1789,In_1864);
xor U4907 (N_4907,In_1582,In_2124);
xor U4908 (N_4908,In_2826,In_1006);
nand U4909 (N_4909,In_2892,In_2963);
nor U4910 (N_4910,In_360,In_1485);
nor U4911 (N_4911,In_2122,In_2988);
and U4912 (N_4912,In_1727,In_113);
and U4913 (N_4913,In_543,In_470);
nor U4914 (N_4914,In_1209,In_1346);
xor U4915 (N_4915,In_2003,In_2933);
and U4916 (N_4916,In_1826,In_860);
nand U4917 (N_4917,In_2934,In_2728);
nand U4918 (N_4918,In_942,In_1160);
or U4919 (N_4919,In_1487,In_2111);
and U4920 (N_4920,In_2652,In_1204);
or U4921 (N_4921,In_1300,In_1892);
and U4922 (N_4922,In_2320,In_1676);
xnor U4923 (N_4923,In_895,In_1897);
xnor U4924 (N_4924,In_2597,In_2851);
and U4925 (N_4925,In_2144,In_937);
nand U4926 (N_4926,In_2049,In_2538);
nand U4927 (N_4927,In_1794,In_2440);
nor U4928 (N_4928,In_2351,In_392);
or U4929 (N_4929,In_1329,In_1585);
or U4930 (N_4930,In_533,In_2237);
nor U4931 (N_4931,In_369,In_640);
nor U4932 (N_4932,In_205,In_2246);
or U4933 (N_4933,In_1007,In_816);
xnor U4934 (N_4934,In_1298,In_2322);
nor U4935 (N_4935,In_1094,In_1902);
xnor U4936 (N_4936,In_2916,In_2273);
or U4937 (N_4937,In_404,In_1950);
nand U4938 (N_4938,In_2524,In_919);
nor U4939 (N_4939,In_343,In_2114);
nor U4940 (N_4940,In_19,In_1411);
xor U4941 (N_4941,In_1089,In_1389);
xor U4942 (N_4942,In_2702,In_233);
nor U4943 (N_4943,In_2807,In_2542);
xnor U4944 (N_4944,In_2735,In_1163);
nor U4945 (N_4945,In_2396,In_2155);
or U4946 (N_4946,In_919,In_42);
and U4947 (N_4947,In_1801,In_2848);
nand U4948 (N_4948,In_1278,In_1088);
nor U4949 (N_4949,In_622,In_1972);
nand U4950 (N_4950,In_602,In_255);
and U4951 (N_4951,In_2074,In_437);
and U4952 (N_4952,In_1017,In_1299);
and U4953 (N_4953,In_947,In_1358);
and U4954 (N_4954,In_959,In_714);
or U4955 (N_4955,In_2024,In_683);
nand U4956 (N_4956,In_2799,In_2067);
nor U4957 (N_4957,In_1330,In_100);
xor U4958 (N_4958,In_2681,In_402);
nor U4959 (N_4959,In_2465,In_2601);
and U4960 (N_4960,In_1656,In_757);
xnor U4961 (N_4961,In_2004,In_733);
nand U4962 (N_4962,In_1299,In_2315);
xnor U4963 (N_4963,In_1844,In_202);
and U4964 (N_4964,In_2540,In_1334);
nand U4965 (N_4965,In_2747,In_2946);
nor U4966 (N_4966,In_799,In_2359);
xor U4967 (N_4967,In_2633,In_1502);
nor U4968 (N_4968,In_1520,In_1786);
or U4969 (N_4969,In_167,In_731);
nor U4970 (N_4970,In_990,In_2443);
or U4971 (N_4971,In_593,In_1080);
and U4972 (N_4972,In_2480,In_1922);
and U4973 (N_4973,In_2783,In_174);
nand U4974 (N_4974,In_97,In_925);
and U4975 (N_4975,In_2690,In_2865);
nor U4976 (N_4976,In_1549,In_2808);
or U4977 (N_4977,In_2703,In_2518);
and U4978 (N_4978,In_67,In_657);
nand U4979 (N_4979,In_1593,In_1508);
nor U4980 (N_4980,In_1581,In_300);
nand U4981 (N_4981,In_1308,In_821);
xor U4982 (N_4982,In_1245,In_644);
and U4983 (N_4983,In_372,In_1955);
and U4984 (N_4984,In_534,In_2530);
or U4985 (N_4985,In_1154,In_460);
nor U4986 (N_4986,In_988,In_1284);
and U4987 (N_4987,In_596,In_1296);
nand U4988 (N_4988,In_1851,In_119);
xor U4989 (N_4989,In_1251,In_500);
nor U4990 (N_4990,In_37,In_295);
or U4991 (N_4991,In_1278,In_390);
nand U4992 (N_4992,In_96,In_513);
or U4993 (N_4993,In_2735,In_2543);
xor U4994 (N_4994,In_510,In_1681);
xor U4995 (N_4995,In_948,In_1552);
and U4996 (N_4996,In_2529,In_1437);
xor U4997 (N_4997,In_2871,In_2858);
xor U4998 (N_4998,In_2593,In_2337);
nor U4999 (N_4999,In_1949,In_2439);
nor U5000 (N_5000,In_2789,In_2321);
and U5001 (N_5001,In_2753,In_2945);
or U5002 (N_5002,In_1465,In_47);
xnor U5003 (N_5003,In_1344,In_1564);
and U5004 (N_5004,In_1882,In_1160);
xnor U5005 (N_5005,In_1889,In_1628);
or U5006 (N_5006,In_2513,In_908);
nand U5007 (N_5007,In_2776,In_1025);
or U5008 (N_5008,In_447,In_2830);
nand U5009 (N_5009,In_2480,In_440);
nor U5010 (N_5010,In_2839,In_2396);
xor U5011 (N_5011,In_1604,In_808);
or U5012 (N_5012,In_1510,In_922);
or U5013 (N_5013,In_2453,In_1856);
or U5014 (N_5014,In_411,In_1154);
nand U5015 (N_5015,In_433,In_1809);
and U5016 (N_5016,In_1952,In_714);
xor U5017 (N_5017,In_593,In_986);
nand U5018 (N_5018,In_1882,In_954);
and U5019 (N_5019,In_1947,In_2940);
or U5020 (N_5020,In_264,In_1065);
or U5021 (N_5021,In_128,In_1934);
or U5022 (N_5022,In_794,In_695);
nor U5023 (N_5023,In_719,In_1313);
and U5024 (N_5024,In_2819,In_228);
and U5025 (N_5025,In_2005,In_1323);
nand U5026 (N_5026,In_2389,In_1496);
nand U5027 (N_5027,In_950,In_249);
or U5028 (N_5028,In_1084,In_1184);
nand U5029 (N_5029,In_2346,In_2515);
nand U5030 (N_5030,In_1295,In_875);
nand U5031 (N_5031,In_1211,In_2193);
nor U5032 (N_5032,In_352,In_249);
xor U5033 (N_5033,In_948,In_668);
nor U5034 (N_5034,In_2319,In_2219);
xor U5035 (N_5035,In_1841,In_601);
or U5036 (N_5036,In_191,In_1486);
nand U5037 (N_5037,In_506,In_1482);
and U5038 (N_5038,In_455,In_1267);
or U5039 (N_5039,In_1781,In_2417);
and U5040 (N_5040,In_459,In_1000);
xor U5041 (N_5041,In_103,In_1018);
nor U5042 (N_5042,In_1327,In_1571);
nor U5043 (N_5043,In_2767,In_1990);
or U5044 (N_5044,In_87,In_1273);
or U5045 (N_5045,In_2195,In_1753);
and U5046 (N_5046,In_633,In_617);
or U5047 (N_5047,In_2787,In_2692);
xor U5048 (N_5048,In_2326,In_1814);
xor U5049 (N_5049,In_633,In_469);
or U5050 (N_5050,In_1996,In_410);
nor U5051 (N_5051,In_1271,In_2042);
nand U5052 (N_5052,In_1112,In_1670);
and U5053 (N_5053,In_2066,In_1445);
nor U5054 (N_5054,In_1613,In_2681);
nor U5055 (N_5055,In_699,In_1967);
and U5056 (N_5056,In_2283,In_1039);
nor U5057 (N_5057,In_326,In_2027);
or U5058 (N_5058,In_1345,In_1784);
nor U5059 (N_5059,In_471,In_1555);
nand U5060 (N_5060,In_2746,In_1185);
nor U5061 (N_5061,In_1486,In_240);
and U5062 (N_5062,In_2839,In_2913);
or U5063 (N_5063,In_2788,In_2201);
nand U5064 (N_5064,In_1087,In_2582);
nand U5065 (N_5065,In_2735,In_683);
nor U5066 (N_5066,In_707,In_2994);
nand U5067 (N_5067,In_1326,In_361);
nand U5068 (N_5068,In_2119,In_1075);
or U5069 (N_5069,In_2382,In_1916);
nand U5070 (N_5070,In_1273,In_2118);
or U5071 (N_5071,In_1045,In_1067);
nor U5072 (N_5072,In_2362,In_843);
or U5073 (N_5073,In_807,In_1470);
nand U5074 (N_5074,In_1058,In_1730);
nand U5075 (N_5075,In_816,In_2464);
and U5076 (N_5076,In_429,In_275);
and U5077 (N_5077,In_2539,In_2893);
and U5078 (N_5078,In_2363,In_64);
nor U5079 (N_5079,In_1679,In_2335);
xor U5080 (N_5080,In_2556,In_1513);
xor U5081 (N_5081,In_339,In_218);
or U5082 (N_5082,In_1919,In_628);
xor U5083 (N_5083,In_2020,In_1987);
nand U5084 (N_5084,In_1415,In_1985);
or U5085 (N_5085,In_2897,In_565);
and U5086 (N_5086,In_1965,In_1353);
and U5087 (N_5087,In_157,In_621);
and U5088 (N_5088,In_2046,In_2877);
or U5089 (N_5089,In_1866,In_2596);
or U5090 (N_5090,In_812,In_2370);
or U5091 (N_5091,In_526,In_620);
and U5092 (N_5092,In_2101,In_1583);
or U5093 (N_5093,In_360,In_2588);
xnor U5094 (N_5094,In_2402,In_1076);
nor U5095 (N_5095,In_2552,In_1492);
and U5096 (N_5096,In_364,In_221);
and U5097 (N_5097,In_602,In_2677);
nor U5098 (N_5098,In_962,In_703);
nor U5099 (N_5099,In_1002,In_706);
and U5100 (N_5100,In_838,In_2575);
nor U5101 (N_5101,In_1797,In_2477);
or U5102 (N_5102,In_52,In_1223);
nor U5103 (N_5103,In_1430,In_900);
or U5104 (N_5104,In_397,In_2388);
nand U5105 (N_5105,In_965,In_654);
nand U5106 (N_5106,In_1200,In_1527);
or U5107 (N_5107,In_2030,In_2990);
nand U5108 (N_5108,In_822,In_2842);
nand U5109 (N_5109,In_295,In_1934);
or U5110 (N_5110,In_2177,In_1173);
xor U5111 (N_5111,In_2596,In_2316);
or U5112 (N_5112,In_300,In_2979);
or U5113 (N_5113,In_2348,In_2133);
and U5114 (N_5114,In_478,In_1264);
nand U5115 (N_5115,In_2817,In_2945);
nand U5116 (N_5116,In_1701,In_2664);
nor U5117 (N_5117,In_1444,In_564);
and U5118 (N_5118,In_641,In_2296);
nand U5119 (N_5119,In_857,In_1867);
and U5120 (N_5120,In_2200,In_1644);
xnor U5121 (N_5121,In_2478,In_2280);
xor U5122 (N_5122,In_2900,In_438);
or U5123 (N_5123,In_1643,In_474);
or U5124 (N_5124,In_916,In_1820);
nand U5125 (N_5125,In_2750,In_762);
nor U5126 (N_5126,In_801,In_1893);
or U5127 (N_5127,In_2262,In_1814);
xnor U5128 (N_5128,In_2566,In_2356);
xnor U5129 (N_5129,In_2985,In_263);
nand U5130 (N_5130,In_907,In_626);
nand U5131 (N_5131,In_2724,In_1794);
xor U5132 (N_5132,In_2149,In_2734);
nor U5133 (N_5133,In_635,In_1323);
nand U5134 (N_5134,In_964,In_2319);
xnor U5135 (N_5135,In_1336,In_2667);
nand U5136 (N_5136,In_550,In_94);
xnor U5137 (N_5137,In_1991,In_1896);
or U5138 (N_5138,In_2672,In_222);
or U5139 (N_5139,In_2997,In_2662);
nor U5140 (N_5140,In_1563,In_2212);
and U5141 (N_5141,In_1752,In_689);
or U5142 (N_5142,In_1177,In_1161);
nor U5143 (N_5143,In_2639,In_2480);
xnor U5144 (N_5144,In_2002,In_657);
or U5145 (N_5145,In_2599,In_2255);
or U5146 (N_5146,In_1528,In_921);
or U5147 (N_5147,In_876,In_628);
or U5148 (N_5148,In_2677,In_645);
and U5149 (N_5149,In_1620,In_254);
xor U5150 (N_5150,In_954,In_2943);
or U5151 (N_5151,In_353,In_1583);
nor U5152 (N_5152,In_1346,In_990);
and U5153 (N_5153,In_1373,In_161);
and U5154 (N_5154,In_2387,In_2748);
xnor U5155 (N_5155,In_2385,In_853);
nor U5156 (N_5156,In_2684,In_1714);
xnor U5157 (N_5157,In_2792,In_512);
and U5158 (N_5158,In_1497,In_2899);
nand U5159 (N_5159,In_1964,In_1053);
xor U5160 (N_5160,In_837,In_414);
nand U5161 (N_5161,In_347,In_449);
xor U5162 (N_5162,In_1668,In_2452);
and U5163 (N_5163,In_430,In_1663);
or U5164 (N_5164,In_1195,In_2864);
or U5165 (N_5165,In_316,In_1719);
nor U5166 (N_5166,In_1893,In_2022);
or U5167 (N_5167,In_1039,In_1009);
xnor U5168 (N_5168,In_2122,In_1136);
nand U5169 (N_5169,In_2357,In_172);
and U5170 (N_5170,In_1416,In_2003);
xor U5171 (N_5171,In_2243,In_2300);
or U5172 (N_5172,In_383,In_2247);
nand U5173 (N_5173,In_1738,In_12);
nor U5174 (N_5174,In_759,In_2358);
xnor U5175 (N_5175,In_2621,In_307);
xor U5176 (N_5176,In_2170,In_2769);
xnor U5177 (N_5177,In_1986,In_766);
xnor U5178 (N_5178,In_838,In_609);
and U5179 (N_5179,In_708,In_369);
nor U5180 (N_5180,In_1943,In_1767);
nand U5181 (N_5181,In_1353,In_2105);
nand U5182 (N_5182,In_1750,In_868);
xor U5183 (N_5183,In_2149,In_702);
or U5184 (N_5184,In_859,In_2668);
and U5185 (N_5185,In_509,In_443);
or U5186 (N_5186,In_1893,In_13);
or U5187 (N_5187,In_1066,In_958);
and U5188 (N_5188,In_1294,In_651);
nand U5189 (N_5189,In_1150,In_2278);
or U5190 (N_5190,In_2967,In_594);
nor U5191 (N_5191,In_1423,In_589);
and U5192 (N_5192,In_935,In_149);
and U5193 (N_5193,In_1722,In_2953);
nand U5194 (N_5194,In_2377,In_267);
or U5195 (N_5195,In_2661,In_1212);
xor U5196 (N_5196,In_349,In_2238);
and U5197 (N_5197,In_1890,In_411);
nor U5198 (N_5198,In_282,In_507);
or U5199 (N_5199,In_1234,In_331);
nor U5200 (N_5200,In_2210,In_1305);
nor U5201 (N_5201,In_1683,In_1853);
nand U5202 (N_5202,In_2408,In_1040);
or U5203 (N_5203,In_1569,In_769);
nand U5204 (N_5204,In_140,In_1563);
nor U5205 (N_5205,In_2710,In_2863);
or U5206 (N_5206,In_2261,In_1713);
or U5207 (N_5207,In_679,In_2044);
and U5208 (N_5208,In_309,In_1360);
nand U5209 (N_5209,In_814,In_1450);
nor U5210 (N_5210,In_1216,In_2207);
xnor U5211 (N_5211,In_1605,In_1852);
and U5212 (N_5212,In_159,In_1891);
and U5213 (N_5213,In_1847,In_1962);
nand U5214 (N_5214,In_1860,In_6);
nor U5215 (N_5215,In_1806,In_2654);
nand U5216 (N_5216,In_1640,In_1413);
nand U5217 (N_5217,In_2043,In_2926);
nor U5218 (N_5218,In_2278,In_1254);
xor U5219 (N_5219,In_1146,In_2961);
nor U5220 (N_5220,In_2634,In_1216);
and U5221 (N_5221,In_2616,In_2318);
and U5222 (N_5222,In_505,In_2017);
nand U5223 (N_5223,In_529,In_1698);
or U5224 (N_5224,In_1505,In_712);
nor U5225 (N_5225,In_86,In_2635);
nand U5226 (N_5226,In_2548,In_2001);
nor U5227 (N_5227,In_622,In_416);
nand U5228 (N_5228,In_1110,In_1049);
or U5229 (N_5229,In_1799,In_1114);
nand U5230 (N_5230,In_2535,In_396);
xnor U5231 (N_5231,In_1484,In_200);
and U5232 (N_5232,In_1715,In_608);
or U5233 (N_5233,In_1355,In_473);
nor U5234 (N_5234,In_1159,In_2717);
or U5235 (N_5235,In_1852,In_205);
or U5236 (N_5236,In_2701,In_1694);
nor U5237 (N_5237,In_160,In_2617);
and U5238 (N_5238,In_2679,In_2861);
and U5239 (N_5239,In_1184,In_2148);
xnor U5240 (N_5240,In_1580,In_820);
xor U5241 (N_5241,In_2292,In_2726);
nand U5242 (N_5242,In_2193,In_656);
nand U5243 (N_5243,In_310,In_1851);
nand U5244 (N_5244,In_2187,In_960);
xor U5245 (N_5245,In_1865,In_100);
or U5246 (N_5246,In_2515,In_2775);
and U5247 (N_5247,In_1583,In_1902);
nor U5248 (N_5248,In_1076,In_2092);
and U5249 (N_5249,In_391,In_958);
xor U5250 (N_5250,In_2552,In_2778);
nor U5251 (N_5251,In_763,In_1678);
nand U5252 (N_5252,In_2445,In_2332);
xor U5253 (N_5253,In_1921,In_1192);
or U5254 (N_5254,In_1999,In_321);
nand U5255 (N_5255,In_1784,In_720);
or U5256 (N_5256,In_2981,In_1644);
nand U5257 (N_5257,In_1467,In_1016);
xnor U5258 (N_5258,In_1322,In_588);
xnor U5259 (N_5259,In_229,In_2215);
nand U5260 (N_5260,In_1736,In_2515);
nor U5261 (N_5261,In_1408,In_2889);
xnor U5262 (N_5262,In_1101,In_470);
nand U5263 (N_5263,In_2555,In_245);
and U5264 (N_5264,In_202,In_462);
or U5265 (N_5265,In_694,In_1170);
or U5266 (N_5266,In_2804,In_913);
or U5267 (N_5267,In_2887,In_983);
xor U5268 (N_5268,In_825,In_2806);
xor U5269 (N_5269,In_1062,In_722);
and U5270 (N_5270,In_1533,In_2649);
and U5271 (N_5271,In_2254,In_2547);
xnor U5272 (N_5272,In_751,In_1976);
and U5273 (N_5273,In_1570,In_1157);
and U5274 (N_5274,In_2479,In_2807);
or U5275 (N_5275,In_515,In_2197);
and U5276 (N_5276,In_1720,In_714);
and U5277 (N_5277,In_1092,In_580);
and U5278 (N_5278,In_36,In_638);
or U5279 (N_5279,In_1316,In_408);
and U5280 (N_5280,In_927,In_424);
nand U5281 (N_5281,In_2429,In_694);
nor U5282 (N_5282,In_1239,In_561);
nor U5283 (N_5283,In_1904,In_913);
and U5284 (N_5284,In_1208,In_238);
or U5285 (N_5285,In_603,In_959);
or U5286 (N_5286,In_1670,In_420);
or U5287 (N_5287,In_2129,In_353);
nor U5288 (N_5288,In_1905,In_557);
xor U5289 (N_5289,In_2627,In_1636);
or U5290 (N_5290,In_1264,In_1388);
nand U5291 (N_5291,In_825,In_86);
nand U5292 (N_5292,In_1405,In_920);
nor U5293 (N_5293,In_2372,In_356);
xnor U5294 (N_5294,In_593,In_789);
and U5295 (N_5295,In_1581,In_685);
and U5296 (N_5296,In_1826,In_2849);
and U5297 (N_5297,In_272,In_2579);
xor U5298 (N_5298,In_355,In_2797);
or U5299 (N_5299,In_2399,In_2844);
nor U5300 (N_5300,In_463,In_420);
or U5301 (N_5301,In_801,In_660);
nor U5302 (N_5302,In_1360,In_572);
xnor U5303 (N_5303,In_1683,In_1478);
nor U5304 (N_5304,In_2116,In_2827);
or U5305 (N_5305,In_2162,In_2516);
xnor U5306 (N_5306,In_109,In_2686);
xor U5307 (N_5307,In_2171,In_161);
xor U5308 (N_5308,In_1559,In_265);
and U5309 (N_5309,In_567,In_1009);
xnor U5310 (N_5310,In_1505,In_120);
or U5311 (N_5311,In_1245,In_1375);
xor U5312 (N_5312,In_1387,In_815);
nor U5313 (N_5313,In_2521,In_2567);
xor U5314 (N_5314,In_2452,In_860);
nor U5315 (N_5315,In_2628,In_103);
or U5316 (N_5316,In_109,In_2029);
or U5317 (N_5317,In_157,In_2952);
nand U5318 (N_5318,In_692,In_2811);
or U5319 (N_5319,In_942,In_546);
xor U5320 (N_5320,In_1973,In_1499);
xnor U5321 (N_5321,In_245,In_2535);
xor U5322 (N_5322,In_1801,In_2102);
and U5323 (N_5323,In_2126,In_1861);
xnor U5324 (N_5324,In_328,In_1264);
nand U5325 (N_5325,In_2045,In_1537);
or U5326 (N_5326,In_1898,In_1727);
nand U5327 (N_5327,In_1112,In_1410);
nor U5328 (N_5328,In_2585,In_2604);
or U5329 (N_5329,In_541,In_1322);
nand U5330 (N_5330,In_142,In_297);
and U5331 (N_5331,In_2603,In_1628);
nand U5332 (N_5332,In_215,In_1784);
nor U5333 (N_5333,In_252,In_1172);
and U5334 (N_5334,In_1472,In_2281);
or U5335 (N_5335,In_1146,In_2933);
xnor U5336 (N_5336,In_1208,In_502);
nand U5337 (N_5337,In_2458,In_1190);
nor U5338 (N_5338,In_527,In_2461);
xor U5339 (N_5339,In_196,In_2511);
nor U5340 (N_5340,In_2646,In_242);
nor U5341 (N_5341,In_1770,In_1372);
nand U5342 (N_5342,In_1850,In_634);
and U5343 (N_5343,In_2352,In_934);
nand U5344 (N_5344,In_109,In_2814);
xor U5345 (N_5345,In_2534,In_52);
nand U5346 (N_5346,In_832,In_286);
nand U5347 (N_5347,In_2529,In_2606);
xnor U5348 (N_5348,In_1097,In_1150);
xor U5349 (N_5349,In_2377,In_2793);
nand U5350 (N_5350,In_974,In_1734);
nor U5351 (N_5351,In_2300,In_1265);
xor U5352 (N_5352,In_2710,In_420);
or U5353 (N_5353,In_2187,In_1982);
or U5354 (N_5354,In_201,In_1701);
and U5355 (N_5355,In_1629,In_1114);
nand U5356 (N_5356,In_1039,In_2216);
xnor U5357 (N_5357,In_2971,In_1717);
xnor U5358 (N_5358,In_2926,In_363);
or U5359 (N_5359,In_1522,In_352);
and U5360 (N_5360,In_986,In_384);
nor U5361 (N_5361,In_463,In_181);
or U5362 (N_5362,In_1217,In_2584);
nand U5363 (N_5363,In_1032,In_2587);
and U5364 (N_5364,In_1088,In_1561);
xnor U5365 (N_5365,In_1528,In_843);
and U5366 (N_5366,In_1206,In_1480);
nor U5367 (N_5367,In_1579,In_1121);
xnor U5368 (N_5368,In_2610,In_2476);
and U5369 (N_5369,In_329,In_723);
xnor U5370 (N_5370,In_2233,In_1720);
or U5371 (N_5371,In_784,In_1742);
or U5372 (N_5372,In_1583,In_151);
xnor U5373 (N_5373,In_1270,In_1830);
xnor U5374 (N_5374,In_1624,In_1768);
nor U5375 (N_5375,In_2517,In_2953);
and U5376 (N_5376,In_517,In_1141);
nand U5377 (N_5377,In_2539,In_790);
xnor U5378 (N_5378,In_2704,In_2277);
or U5379 (N_5379,In_227,In_1577);
xnor U5380 (N_5380,In_596,In_1929);
and U5381 (N_5381,In_624,In_529);
or U5382 (N_5382,In_1213,In_1683);
nand U5383 (N_5383,In_297,In_190);
nand U5384 (N_5384,In_1772,In_1696);
or U5385 (N_5385,In_919,In_565);
nand U5386 (N_5386,In_1192,In_19);
nor U5387 (N_5387,In_976,In_1609);
and U5388 (N_5388,In_958,In_1985);
or U5389 (N_5389,In_2233,In_1382);
nand U5390 (N_5390,In_87,In_2356);
xor U5391 (N_5391,In_932,In_2920);
or U5392 (N_5392,In_2501,In_665);
xor U5393 (N_5393,In_1648,In_647);
nand U5394 (N_5394,In_2155,In_343);
or U5395 (N_5395,In_850,In_2362);
xor U5396 (N_5396,In_2342,In_429);
or U5397 (N_5397,In_1346,In_895);
xnor U5398 (N_5398,In_28,In_2166);
and U5399 (N_5399,In_1797,In_857);
xor U5400 (N_5400,In_2028,In_1616);
nor U5401 (N_5401,In_1325,In_984);
nor U5402 (N_5402,In_1165,In_2016);
nand U5403 (N_5403,In_1430,In_2456);
or U5404 (N_5404,In_1921,In_1733);
or U5405 (N_5405,In_239,In_2099);
nand U5406 (N_5406,In_561,In_762);
or U5407 (N_5407,In_2923,In_9);
nand U5408 (N_5408,In_2628,In_2992);
or U5409 (N_5409,In_2689,In_1259);
nor U5410 (N_5410,In_1902,In_2460);
nand U5411 (N_5411,In_2767,In_494);
and U5412 (N_5412,In_1711,In_726);
and U5413 (N_5413,In_380,In_1088);
xor U5414 (N_5414,In_2032,In_626);
xnor U5415 (N_5415,In_1359,In_2664);
nor U5416 (N_5416,In_223,In_924);
and U5417 (N_5417,In_1060,In_1169);
or U5418 (N_5418,In_2990,In_2557);
xnor U5419 (N_5419,In_2919,In_2237);
nand U5420 (N_5420,In_1791,In_139);
or U5421 (N_5421,In_1960,In_237);
or U5422 (N_5422,In_697,In_504);
nand U5423 (N_5423,In_2149,In_1070);
and U5424 (N_5424,In_1151,In_2953);
nor U5425 (N_5425,In_2526,In_122);
or U5426 (N_5426,In_2176,In_2512);
or U5427 (N_5427,In_790,In_1292);
nor U5428 (N_5428,In_2919,In_814);
or U5429 (N_5429,In_585,In_1354);
xor U5430 (N_5430,In_1084,In_407);
nor U5431 (N_5431,In_2679,In_1176);
nor U5432 (N_5432,In_1059,In_1556);
nand U5433 (N_5433,In_2152,In_756);
and U5434 (N_5434,In_1983,In_899);
and U5435 (N_5435,In_392,In_570);
and U5436 (N_5436,In_2583,In_2874);
or U5437 (N_5437,In_270,In_266);
and U5438 (N_5438,In_1878,In_2833);
or U5439 (N_5439,In_88,In_656);
nor U5440 (N_5440,In_1941,In_2131);
nor U5441 (N_5441,In_2324,In_2388);
and U5442 (N_5442,In_1121,In_2737);
nand U5443 (N_5443,In_2750,In_1441);
nand U5444 (N_5444,In_1437,In_664);
nand U5445 (N_5445,In_2415,In_2056);
or U5446 (N_5446,In_277,In_1678);
and U5447 (N_5447,In_1698,In_1683);
and U5448 (N_5448,In_837,In_2209);
nand U5449 (N_5449,In_1833,In_690);
and U5450 (N_5450,In_564,In_2461);
xnor U5451 (N_5451,In_2923,In_2233);
and U5452 (N_5452,In_568,In_586);
and U5453 (N_5453,In_2228,In_2050);
nand U5454 (N_5454,In_2830,In_1804);
and U5455 (N_5455,In_2323,In_525);
nor U5456 (N_5456,In_1040,In_100);
or U5457 (N_5457,In_717,In_1249);
xor U5458 (N_5458,In_886,In_2414);
nand U5459 (N_5459,In_920,In_2083);
nand U5460 (N_5460,In_1628,In_1599);
and U5461 (N_5461,In_611,In_1617);
xnor U5462 (N_5462,In_28,In_1476);
nor U5463 (N_5463,In_951,In_1924);
nand U5464 (N_5464,In_2469,In_486);
nand U5465 (N_5465,In_2489,In_790);
xnor U5466 (N_5466,In_2572,In_2217);
or U5467 (N_5467,In_2051,In_208);
and U5468 (N_5468,In_2035,In_19);
nor U5469 (N_5469,In_2917,In_1880);
nand U5470 (N_5470,In_1042,In_1688);
nor U5471 (N_5471,In_1382,In_1062);
nor U5472 (N_5472,In_2256,In_1606);
or U5473 (N_5473,In_480,In_1815);
xnor U5474 (N_5474,In_2676,In_1658);
nor U5475 (N_5475,In_161,In_1908);
and U5476 (N_5476,In_806,In_2362);
and U5477 (N_5477,In_1059,In_2756);
nand U5478 (N_5478,In_2086,In_2933);
nand U5479 (N_5479,In_2658,In_2149);
nand U5480 (N_5480,In_2013,In_1643);
and U5481 (N_5481,In_2649,In_1809);
and U5482 (N_5482,In_1640,In_272);
nand U5483 (N_5483,In_1025,In_2730);
and U5484 (N_5484,In_2672,In_1263);
or U5485 (N_5485,In_1446,In_1958);
nor U5486 (N_5486,In_1243,In_2826);
nor U5487 (N_5487,In_1741,In_1573);
and U5488 (N_5488,In_1551,In_184);
nor U5489 (N_5489,In_2782,In_2507);
and U5490 (N_5490,In_1040,In_783);
xnor U5491 (N_5491,In_387,In_687);
and U5492 (N_5492,In_2146,In_1164);
nand U5493 (N_5493,In_1439,In_1746);
or U5494 (N_5494,In_474,In_2661);
nand U5495 (N_5495,In_1090,In_611);
nand U5496 (N_5496,In_2383,In_714);
or U5497 (N_5497,In_2767,In_2250);
and U5498 (N_5498,In_2192,In_675);
xnor U5499 (N_5499,In_265,In_2351);
and U5500 (N_5500,In_2132,In_2995);
nand U5501 (N_5501,In_18,In_1692);
nand U5502 (N_5502,In_2293,In_2572);
nand U5503 (N_5503,In_2856,In_846);
or U5504 (N_5504,In_2595,In_2159);
nor U5505 (N_5505,In_816,In_709);
and U5506 (N_5506,In_946,In_1093);
nor U5507 (N_5507,In_851,In_1410);
nand U5508 (N_5508,In_439,In_1946);
and U5509 (N_5509,In_623,In_743);
or U5510 (N_5510,In_216,In_2980);
xnor U5511 (N_5511,In_798,In_686);
and U5512 (N_5512,In_586,In_2008);
or U5513 (N_5513,In_2212,In_273);
and U5514 (N_5514,In_2594,In_149);
or U5515 (N_5515,In_2610,In_806);
xnor U5516 (N_5516,In_2627,In_2223);
nor U5517 (N_5517,In_2409,In_1027);
and U5518 (N_5518,In_1782,In_2067);
xnor U5519 (N_5519,In_1500,In_2546);
or U5520 (N_5520,In_2312,In_1501);
and U5521 (N_5521,In_8,In_1264);
nor U5522 (N_5522,In_421,In_1171);
nand U5523 (N_5523,In_2746,In_1071);
xnor U5524 (N_5524,In_1643,In_2569);
xor U5525 (N_5525,In_506,In_370);
and U5526 (N_5526,In_1029,In_1844);
and U5527 (N_5527,In_169,In_1004);
nand U5528 (N_5528,In_1458,In_2123);
nor U5529 (N_5529,In_367,In_582);
nand U5530 (N_5530,In_1131,In_906);
xnor U5531 (N_5531,In_1883,In_657);
or U5532 (N_5532,In_1890,In_1752);
xor U5533 (N_5533,In_496,In_1512);
and U5534 (N_5534,In_2957,In_2805);
nand U5535 (N_5535,In_1953,In_2448);
or U5536 (N_5536,In_1537,In_1349);
or U5537 (N_5537,In_2755,In_1059);
or U5538 (N_5538,In_839,In_2828);
nand U5539 (N_5539,In_105,In_2107);
nand U5540 (N_5540,In_1996,In_2009);
and U5541 (N_5541,In_1017,In_68);
and U5542 (N_5542,In_675,In_1926);
nor U5543 (N_5543,In_2864,In_555);
nand U5544 (N_5544,In_601,In_2842);
nor U5545 (N_5545,In_2526,In_940);
nand U5546 (N_5546,In_2337,In_682);
or U5547 (N_5547,In_1439,In_1330);
nand U5548 (N_5548,In_2103,In_1207);
nor U5549 (N_5549,In_1679,In_1811);
xnor U5550 (N_5550,In_716,In_2685);
or U5551 (N_5551,In_463,In_153);
nor U5552 (N_5552,In_1798,In_333);
xnor U5553 (N_5553,In_1066,In_762);
or U5554 (N_5554,In_2304,In_1995);
and U5555 (N_5555,In_2920,In_880);
or U5556 (N_5556,In_1280,In_2095);
nor U5557 (N_5557,In_1787,In_1450);
xor U5558 (N_5558,In_2769,In_1348);
nor U5559 (N_5559,In_2500,In_335);
nor U5560 (N_5560,In_1901,In_964);
nand U5561 (N_5561,In_1841,In_312);
nor U5562 (N_5562,In_2820,In_957);
nand U5563 (N_5563,In_492,In_1503);
nand U5564 (N_5564,In_1802,In_683);
and U5565 (N_5565,In_1262,In_743);
nand U5566 (N_5566,In_1339,In_1778);
or U5567 (N_5567,In_1816,In_1680);
xor U5568 (N_5568,In_2851,In_902);
or U5569 (N_5569,In_426,In_756);
xnor U5570 (N_5570,In_594,In_2451);
or U5571 (N_5571,In_234,In_2772);
nor U5572 (N_5572,In_2902,In_1816);
or U5573 (N_5573,In_1389,In_271);
xnor U5574 (N_5574,In_306,In_456);
nor U5575 (N_5575,In_2362,In_2068);
nand U5576 (N_5576,In_323,In_218);
or U5577 (N_5577,In_1320,In_1641);
or U5578 (N_5578,In_1635,In_1202);
nand U5579 (N_5579,In_2813,In_2410);
xnor U5580 (N_5580,In_2990,In_1189);
nor U5581 (N_5581,In_664,In_1178);
nand U5582 (N_5582,In_2244,In_2434);
nand U5583 (N_5583,In_813,In_862);
nor U5584 (N_5584,In_388,In_841);
and U5585 (N_5585,In_1349,In_968);
and U5586 (N_5586,In_793,In_2865);
or U5587 (N_5587,In_2579,In_823);
and U5588 (N_5588,In_46,In_2307);
or U5589 (N_5589,In_1121,In_1584);
or U5590 (N_5590,In_1647,In_2815);
and U5591 (N_5591,In_2758,In_1176);
nand U5592 (N_5592,In_1185,In_641);
or U5593 (N_5593,In_1722,In_2130);
xor U5594 (N_5594,In_1957,In_1964);
and U5595 (N_5595,In_1841,In_2427);
or U5596 (N_5596,In_396,In_2288);
xnor U5597 (N_5597,In_1563,In_294);
nor U5598 (N_5598,In_2355,In_1282);
nor U5599 (N_5599,In_939,In_602);
nor U5600 (N_5600,In_2083,In_283);
nand U5601 (N_5601,In_2270,In_1076);
nand U5602 (N_5602,In_771,In_2818);
or U5603 (N_5603,In_1559,In_2915);
xor U5604 (N_5604,In_1888,In_2559);
nor U5605 (N_5605,In_522,In_1888);
nor U5606 (N_5606,In_917,In_2542);
xor U5607 (N_5607,In_1142,In_1691);
or U5608 (N_5608,In_407,In_16);
nor U5609 (N_5609,In_1482,In_1820);
xnor U5610 (N_5610,In_579,In_2450);
and U5611 (N_5611,In_2568,In_2484);
nand U5612 (N_5612,In_1695,In_571);
or U5613 (N_5613,In_1436,In_264);
or U5614 (N_5614,In_2330,In_1660);
nand U5615 (N_5615,In_2360,In_1286);
or U5616 (N_5616,In_1249,In_645);
and U5617 (N_5617,In_1054,In_1618);
and U5618 (N_5618,In_1779,In_2928);
nor U5619 (N_5619,In_1867,In_2338);
nor U5620 (N_5620,In_1602,In_557);
xor U5621 (N_5621,In_2789,In_644);
and U5622 (N_5622,In_1178,In_26);
xor U5623 (N_5623,In_44,In_467);
and U5624 (N_5624,In_2110,In_2192);
nor U5625 (N_5625,In_2856,In_1931);
or U5626 (N_5626,In_2412,In_226);
nor U5627 (N_5627,In_1004,In_1392);
and U5628 (N_5628,In_1830,In_2122);
and U5629 (N_5629,In_1282,In_2725);
nor U5630 (N_5630,In_2670,In_1047);
or U5631 (N_5631,In_330,In_893);
nor U5632 (N_5632,In_1759,In_1603);
nor U5633 (N_5633,In_447,In_775);
nand U5634 (N_5634,In_179,In_27);
and U5635 (N_5635,In_127,In_2028);
nor U5636 (N_5636,In_2607,In_1933);
and U5637 (N_5637,In_1427,In_1278);
nand U5638 (N_5638,In_2038,In_2726);
nor U5639 (N_5639,In_2777,In_376);
nor U5640 (N_5640,In_2757,In_811);
and U5641 (N_5641,In_1207,In_258);
nand U5642 (N_5642,In_1186,In_311);
xnor U5643 (N_5643,In_2434,In_2873);
or U5644 (N_5644,In_2078,In_2532);
nor U5645 (N_5645,In_1465,In_1500);
nor U5646 (N_5646,In_1615,In_2039);
nand U5647 (N_5647,In_823,In_1060);
or U5648 (N_5648,In_162,In_341);
xnor U5649 (N_5649,In_2937,In_1242);
nand U5650 (N_5650,In_2730,In_2773);
and U5651 (N_5651,In_2636,In_254);
or U5652 (N_5652,In_462,In_1546);
nor U5653 (N_5653,In_2952,In_1016);
nand U5654 (N_5654,In_1085,In_2954);
xnor U5655 (N_5655,In_2059,In_2895);
nor U5656 (N_5656,In_1472,In_1688);
and U5657 (N_5657,In_722,In_204);
nor U5658 (N_5658,In_1575,In_1390);
and U5659 (N_5659,In_2870,In_441);
nand U5660 (N_5660,In_2531,In_2517);
and U5661 (N_5661,In_530,In_2217);
and U5662 (N_5662,In_642,In_214);
nand U5663 (N_5663,In_2443,In_2869);
and U5664 (N_5664,In_659,In_2601);
or U5665 (N_5665,In_1117,In_2276);
xnor U5666 (N_5666,In_434,In_2445);
nor U5667 (N_5667,In_721,In_587);
nor U5668 (N_5668,In_1072,In_1999);
nor U5669 (N_5669,In_2510,In_1471);
nor U5670 (N_5670,In_49,In_1025);
nand U5671 (N_5671,In_2330,In_732);
and U5672 (N_5672,In_1388,In_273);
or U5673 (N_5673,In_336,In_1996);
xnor U5674 (N_5674,In_435,In_937);
and U5675 (N_5675,In_2495,In_933);
nor U5676 (N_5676,In_843,In_1428);
nor U5677 (N_5677,In_1251,In_2445);
and U5678 (N_5678,In_1584,In_2859);
nor U5679 (N_5679,In_1117,In_2113);
nor U5680 (N_5680,In_490,In_1220);
or U5681 (N_5681,In_1684,In_67);
xor U5682 (N_5682,In_2956,In_720);
nand U5683 (N_5683,In_2921,In_2826);
and U5684 (N_5684,In_2796,In_408);
nand U5685 (N_5685,In_1693,In_2611);
or U5686 (N_5686,In_1503,In_283);
xnor U5687 (N_5687,In_846,In_2829);
xor U5688 (N_5688,In_1505,In_1548);
nand U5689 (N_5689,In_2793,In_2897);
nor U5690 (N_5690,In_713,In_2210);
or U5691 (N_5691,In_847,In_1449);
nor U5692 (N_5692,In_1297,In_1462);
nand U5693 (N_5693,In_2564,In_1748);
nor U5694 (N_5694,In_669,In_1320);
nor U5695 (N_5695,In_2218,In_988);
and U5696 (N_5696,In_2231,In_1768);
xnor U5697 (N_5697,In_2697,In_513);
nand U5698 (N_5698,In_2670,In_204);
and U5699 (N_5699,In_462,In_2194);
nand U5700 (N_5700,In_1603,In_943);
nand U5701 (N_5701,In_2472,In_2770);
and U5702 (N_5702,In_47,In_1094);
xnor U5703 (N_5703,In_2126,In_2808);
nor U5704 (N_5704,In_350,In_2746);
or U5705 (N_5705,In_2704,In_2407);
and U5706 (N_5706,In_928,In_1254);
and U5707 (N_5707,In_1510,In_2563);
nor U5708 (N_5708,In_2234,In_2077);
xor U5709 (N_5709,In_115,In_1057);
xor U5710 (N_5710,In_2488,In_283);
xor U5711 (N_5711,In_2367,In_95);
nand U5712 (N_5712,In_1557,In_541);
nor U5713 (N_5713,In_589,In_706);
nor U5714 (N_5714,In_1177,In_1061);
nand U5715 (N_5715,In_1826,In_2261);
nor U5716 (N_5716,In_2144,In_1833);
and U5717 (N_5717,In_1155,In_265);
and U5718 (N_5718,In_157,In_2772);
nand U5719 (N_5719,In_2324,In_2532);
nand U5720 (N_5720,In_2206,In_1576);
nand U5721 (N_5721,In_2731,In_1585);
nor U5722 (N_5722,In_516,In_1468);
nor U5723 (N_5723,In_2798,In_1120);
or U5724 (N_5724,In_599,In_2644);
xnor U5725 (N_5725,In_671,In_307);
or U5726 (N_5726,In_2061,In_1508);
or U5727 (N_5727,In_456,In_1195);
and U5728 (N_5728,In_2925,In_914);
xnor U5729 (N_5729,In_2077,In_2539);
nand U5730 (N_5730,In_2966,In_1919);
or U5731 (N_5731,In_2165,In_2775);
nand U5732 (N_5732,In_649,In_1927);
nor U5733 (N_5733,In_1242,In_1753);
or U5734 (N_5734,In_1228,In_2314);
and U5735 (N_5735,In_269,In_1024);
and U5736 (N_5736,In_343,In_2140);
xor U5737 (N_5737,In_970,In_2644);
and U5738 (N_5738,In_2539,In_1798);
and U5739 (N_5739,In_1567,In_2653);
xnor U5740 (N_5740,In_397,In_99);
xnor U5741 (N_5741,In_144,In_1482);
nand U5742 (N_5742,In_2615,In_881);
xnor U5743 (N_5743,In_2007,In_1610);
and U5744 (N_5744,In_1118,In_135);
or U5745 (N_5745,In_1309,In_1722);
or U5746 (N_5746,In_2199,In_976);
and U5747 (N_5747,In_2676,In_2609);
nor U5748 (N_5748,In_796,In_2890);
xnor U5749 (N_5749,In_2045,In_2309);
and U5750 (N_5750,In_997,In_210);
and U5751 (N_5751,In_2777,In_668);
xor U5752 (N_5752,In_1810,In_2498);
and U5753 (N_5753,In_2470,In_300);
nand U5754 (N_5754,In_2398,In_2341);
or U5755 (N_5755,In_1944,In_943);
and U5756 (N_5756,In_1800,In_553);
and U5757 (N_5757,In_2333,In_437);
or U5758 (N_5758,In_76,In_245);
or U5759 (N_5759,In_1831,In_2090);
and U5760 (N_5760,In_997,In_2860);
and U5761 (N_5761,In_999,In_2687);
xor U5762 (N_5762,In_1375,In_527);
nand U5763 (N_5763,In_2832,In_1542);
nor U5764 (N_5764,In_2598,In_2724);
nor U5765 (N_5765,In_2089,In_886);
nor U5766 (N_5766,In_517,In_359);
and U5767 (N_5767,In_2365,In_1417);
nor U5768 (N_5768,In_1575,In_2736);
nand U5769 (N_5769,In_2639,In_2850);
nand U5770 (N_5770,In_1568,In_2309);
and U5771 (N_5771,In_2095,In_1838);
nand U5772 (N_5772,In_2655,In_1654);
nor U5773 (N_5773,In_2858,In_1860);
or U5774 (N_5774,In_762,In_1419);
and U5775 (N_5775,In_822,In_76);
nor U5776 (N_5776,In_826,In_234);
xnor U5777 (N_5777,In_2161,In_283);
and U5778 (N_5778,In_1460,In_2908);
xnor U5779 (N_5779,In_1272,In_2827);
nand U5780 (N_5780,In_471,In_1004);
xnor U5781 (N_5781,In_184,In_1495);
or U5782 (N_5782,In_2632,In_49);
xor U5783 (N_5783,In_555,In_1383);
nor U5784 (N_5784,In_1933,In_1036);
xnor U5785 (N_5785,In_812,In_1066);
nand U5786 (N_5786,In_2967,In_876);
and U5787 (N_5787,In_930,In_2660);
nand U5788 (N_5788,In_732,In_436);
xnor U5789 (N_5789,In_874,In_447);
nand U5790 (N_5790,In_1957,In_1328);
or U5791 (N_5791,In_2173,In_1554);
and U5792 (N_5792,In_1092,In_183);
or U5793 (N_5793,In_757,In_1350);
xnor U5794 (N_5794,In_205,In_2);
nor U5795 (N_5795,In_1928,In_2930);
and U5796 (N_5796,In_2940,In_784);
nand U5797 (N_5797,In_449,In_2426);
nor U5798 (N_5798,In_1529,In_1736);
nand U5799 (N_5799,In_2647,In_2335);
or U5800 (N_5800,In_2580,In_1472);
or U5801 (N_5801,In_327,In_1979);
and U5802 (N_5802,In_1323,In_489);
xor U5803 (N_5803,In_2976,In_2885);
nor U5804 (N_5804,In_2290,In_381);
or U5805 (N_5805,In_1698,In_2357);
nand U5806 (N_5806,In_1716,In_1714);
xnor U5807 (N_5807,In_1510,In_1006);
nor U5808 (N_5808,In_2796,In_2204);
xor U5809 (N_5809,In_2852,In_1029);
and U5810 (N_5810,In_2127,In_2311);
nor U5811 (N_5811,In_2109,In_580);
nor U5812 (N_5812,In_2103,In_2143);
nand U5813 (N_5813,In_769,In_2045);
nand U5814 (N_5814,In_2899,In_345);
xnor U5815 (N_5815,In_734,In_1799);
or U5816 (N_5816,In_2506,In_1491);
nor U5817 (N_5817,In_2119,In_2074);
nand U5818 (N_5818,In_538,In_381);
nor U5819 (N_5819,In_113,In_1173);
xnor U5820 (N_5820,In_937,In_283);
nand U5821 (N_5821,In_398,In_733);
and U5822 (N_5822,In_565,In_75);
and U5823 (N_5823,In_1828,In_134);
xnor U5824 (N_5824,In_1417,In_2528);
xnor U5825 (N_5825,In_591,In_675);
or U5826 (N_5826,In_890,In_1812);
xnor U5827 (N_5827,In_2486,In_1389);
nor U5828 (N_5828,In_2475,In_2933);
nor U5829 (N_5829,In_2297,In_1984);
nand U5830 (N_5830,In_2121,In_465);
and U5831 (N_5831,In_6,In_2723);
nand U5832 (N_5832,In_1805,In_2570);
xnor U5833 (N_5833,In_1326,In_2634);
xnor U5834 (N_5834,In_1133,In_2009);
and U5835 (N_5835,In_2749,In_528);
xnor U5836 (N_5836,In_2334,In_876);
and U5837 (N_5837,In_739,In_1992);
or U5838 (N_5838,In_1335,In_2357);
and U5839 (N_5839,In_292,In_2784);
or U5840 (N_5840,In_1101,In_909);
nor U5841 (N_5841,In_1253,In_1662);
nand U5842 (N_5842,In_109,In_1167);
and U5843 (N_5843,In_2967,In_2588);
and U5844 (N_5844,In_612,In_541);
or U5845 (N_5845,In_1091,In_2699);
and U5846 (N_5846,In_2839,In_396);
and U5847 (N_5847,In_2013,In_920);
xnor U5848 (N_5848,In_1622,In_2216);
or U5849 (N_5849,In_2595,In_1021);
xor U5850 (N_5850,In_1032,In_584);
nand U5851 (N_5851,In_2229,In_2659);
or U5852 (N_5852,In_1516,In_1027);
and U5853 (N_5853,In_1258,In_306);
nand U5854 (N_5854,In_2892,In_2935);
and U5855 (N_5855,In_2858,In_2067);
or U5856 (N_5856,In_952,In_10);
or U5857 (N_5857,In_1523,In_2905);
xor U5858 (N_5858,In_98,In_2358);
nand U5859 (N_5859,In_142,In_177);
xnor U5860 (N_5860,In_2724,In_785);
or U5861 (N_5861,In_1798,In_518);
and U5862 (N_5862,In_1373,In_2466);
and U5863 (N_5863,In_1670,In_310);
or U5864 (N_5864,In_1051,In_1200);
nor U5865 (N_5865,In_2119,In_177);
and U5866 (N_5866,In_824,In_625);
or U5867 (N_5867,In_266,In_515);
and U5868 (N_5868,In_2627,In_1419);
nor U5869 (N_5869,In_882,In_2015);
xor U5870 (N_5870,In_354,In_567);
nand U5871 (N_5871,In_1925,In_43);
and U5872 (N_5872,In_2989,In_2503);
or U5873 (N_5873,In_1337,In_1222);
or U5874 (N_5874,In_2119,In_2979);
and U5875 (N_5875,In_2586,In_628);
xnor U5876 (N_5876,In_609,In_1448);
nand U5877 (N_5877,In_2346,In_1460);
nor U5878 (N_5878,In_35,In_1945);
and U5879 (N_5879,In_2547,In_623);
xor U5880 (N_5880,In_1687,In_2304);
or U5881 (N_5881,In_467,In_2671);
nand U5882 (N_5882,In_1020,In_2931);
or U5883 (N_5883,In_574,In_994);
nand U5884 (N_5884,In_548,In_890);
or U5885 (N_5885,In_2805,In_2157);
xnor U5886 (N_5886,In_246,In_2001);
xnor U5887 (N_5887,In_1318,In_1260);
nand U5888 (N_5888,In_8,In_1916);
xor U5889 (N_5889,In_46,In_1861);
and U5890 (N_5890,In_2226,In_1429);
nand U5891 (N_5891,In_1815,In_1710);
xor U5892 (N_5892,In_1286,In_2451);
nand U5893 (N_5893,In_299,In_2937);
nand U5894 (N_5894,In_2606,In_138);
and U5895 (N_5895,In_259,In_2912);
nor U5896 (N_5896,In_1780,In_618);
or U5897 (N_5897,In_2802,In_2636);
nor U5898 (N_5898,In_967,In_509);
and U5899 (N_5899,In_2126,In_2511);
nand U5900 (N_5900,In_1585,In_1198);
or U5901 (N_5901,In_903,In_2932);
and U5902 (N_5902,In_2825,In_1691);
nand U5903 (N_5903,In_966,In_1844);
nor U5904 (N_5904,In_596,In_2355);
nor U5905 (N_5905,In_1120,In_2718);
nand U5906 (N_5906,In_1449,In_2792);
xnor U5907 (N_5907,In_1700,In_2420);
or U5908 (N_5908,In_1479,In_2460);
nand U5909 (N_5909,In_368,In_1907);
nand U5910 (N_5910,In_1446,In_2358);
xor U5911 (N_5911,In_2183,In_1609);
nand U5912 (N_5912,In_374,In_950);
or U5913 (N_5913,In_2931,In_2703);
nor U5914 (N_5914,In_2687,In_2857);
and U5915 (N_5915,In_2585,In_2213);
or U5916 (N_5916,In_2286,In_2049);
and U5917 (N_5917,In_2017,In_2804);
xnor U5918 (N_5918,In_2010,In_2677);
xnor U5919 (N_5919,In_1092,In_62);
or U5920 (N_5920,In_581,In_946);
nor U5921 (N_5921,In_616,In_2508);
nand U5922 (N_5922,In_2976,In_364);
nand U5923 (N_5923,In_914,In_799);
or U5924 (N_5924,In_2339,In_1395);
and U5925 (N_5925,In_1854,In_286);
nand U5926 (N_5926,In_293,In_249);
or U5927 (N_5927,In_1324,In_98);
nor U5928 (N_5928,In_2398,In_2106);
and U5929 (N_5929,In_1903,In_1868);
nand U5930 (N_5930,In_1320,In_1906);
or U5931 (N_5931,In_2739,In_2035);
nand U5932 (N_5932,In_2597,In_2814);
xnor U5933 (N_5933,In_2944,In_2829);
nor U5934 (N_5934,In_1110,In_2038);
nand U5935 (N_5935,In_885,In_1082);
or U5936 (N_5936,In_2013,In_2003);
xnor U5937 (N_5937,In_1189,In_487);
and U5938 (N_5938,In_2985,In_217);
nand U5939 (N_5939,In_801,In_1740);
xnor U5940 (N_5940,In_40,In_2262);
xnor U5941 (N_5941,In_476,In_2533);
xnor U5942 (N_5942,In_1230,In_2685);
and U5943 (N_5943,In_715,In_1207);
and U5944 (N_5944,In_1938,In_2506);
xor U5945 (N_5945,In_1080,In_1983);
nand U5946 (N_5946,In_2226,In_108);
xnor U5947 (N_5947,In_2096,In_1229);
nor U5948 (N_5948,In_1303,In_1588);
nor U5949 (N_5949,In_2850,In_96);
nor U5950 (N_5950,In_2045,In_2934);
nand U5951 (N_5951,In_987,In_1255);
nand U5952 (N_5952,In_920,In_396);
nand U5953 (N_5953,In_1521,In_1320);
and U5954 (N_5954,In_2507,In_2812);
nand U5955 (N_5955,In_1760,In_1492);
nand U5956 (N_5956,In_2432,In_601);
nand U5957 (N_5957,In_537,In_1525);
nor U5958 (N_5958,In_722,In_1658);
nor U5959 (N_5959,In_1764,In_2101);
xor U5960 (N_5960,In_2758,In_218);
nand U5961 (N_5961,In_2828,In_289);
nand U5962 (N_5962,In_1080,In_456);
xnor U5963 (N_5963,In_2186,In_1176);
nand U5964 (N_5964,In_2960,In_832);
xor U5965 (N_5965,In_1764,In_1002);
nand U5966 (N_5966,In_650,In_579);
or U5967 (N_5967,In_256,In_2490);
xor U5968 (N_5968,In_2218,In_1573);
or U5969 (N_5969,In_335,In_1653);
and U5970 (N_5970,In_50,In_2430);
nand U5971 (N_5971,In_2999,In_1029);
and U5972 (N_5972,In_1360,In_1677);
or U5973 (N_5973,In_359,In_1227);
nand U5974 (N_5974,In_32,In_1290);
nand U5975 (N_5975,In_412,In_818);
nor U5976 (N_5976,In_1379,In_985);
nand U5977 (N_5977,In_179,In_2398);
nor U5978 (N_5978,In_1832,In_1160);
or U5979 (N_5979,In_2940,In_1895);
xor U5980 (N_5980,In_1341,In_1787);
or U5981 (N_5981,In_1239,In_2017);
or U5982 (N_5982,In_1967,In_682);
or U5983 (N_5983,In_1017,In_2368);
nand U5984 (N_5984,In_1394,In_1476);
nor U5985 (N_5985,In_1212,In_1645);
nand U5986 (N_5986,In_360,In_1041);
and U5987 (N_5987,In_2878,In_266);
nand U5988 (N_5988,In_2613,In_1096);
and U5989 (N_5989,In_411,In_2515);
nand U5990 (N_5990,In_2813,In_1904);
xnor U5991 (N_5991,In_2358,In_1245);
xnor U5992 (N_5992,In_1623,In_716);
or U5993 (N_5993,In_378,In_1053);
nor U5994 (N_5994,In_2479,In_9);
nand U5995 (N_5995,In_886,In_2486);
or U5996 (N_5996,In_946,In_1049);
nand U5997 (N_5997,In_1240,In_368);
and U5998 (N_5998,In_1755,In_1518);
xnor U5999 (N_5999,In_2604,In_295);
and U6000 (N_6000,N_4230,N_274);
xnor U6001 (N_6001,N_4107,N_2543);
nand U6002 (N_6002,N_5413,N_89);
nor U6003 (N_6003,N_1420,N_4478);
xnor U6004 (N_6004,N_4277,N_2667);
xor U6005 (N_6005,N_5773,N_4196);
xnor U6006 (N_6006,N_556,N_768);
nand U6007 (N_6007,N_3867,N_2856);
and U6008 (N_6008,N_3395,N_2273);
and U6009 (N_6009,N_3797,N_4202);
nor U6010 (N_6010,N_4706,N_4036);
and U6011 (N_6011,N_3682,N_1450);
or U6012 (N_6012,N_1237,N_1762);
or U6013 (N_6013,N_5264,N_1020);
and U6014 (N_6014,N_1586,N_2737);
xnor U6015 (N_6015,N_2008,N_5458);
nand U6016 (N_6016,N_3231,N_4805);
nor U6017 (N_6017,N_4042,N_2266);
xor U6018 (N_6018,N_4345,N_5422);
nand U6019 (N_6019,N_5908,N_1238);
and U6020 (N_6020,N_3576,N_5401);
nor U6021 (N_6021,N_93,N_3195);
xnor U6022 (N_6022,N_3675,N_4873);
nand U6023 (N_6023,N_3507,N_4405);
and U6024 (N_6024,N_2231,N_3178);
nor U6025 (N_6025,N_3976,N_791);
nor U6026 (N_6026,N_5251,N_1997);
and U6027 (N_6027,N_4882,N_924);
nand U6028 (N_6028,N_5728,N_2686);
nand U6029 (N_6029,N_2953,N_216);
and U6030 (N_6030,N_2896,N_3424);
nand U6031 (N_6031,N_573,N_3447);
xor U6032 (N_6032,N_1977,N_98);
or U6033 (N_6033,N_1448,N_1918);
nand U6034 (N_6034,N_4408,N_4261);
or U6035 (N_6035,N_5989,N_1011);
nor U6036 (N_6036,N_4470,N_1151);
nand U6037 (N_6037,N_2436,N_235);
nor U6038 (N_6038,N_905,N_3311);
xor U6039 (N_6039,N_3679,N_2264);
and U6040 (N_6040,N_56,N_4916);
or U6041 (N_6041,N_4495,N_5022);
nand U6042 (N_6042,N_3446,N_1489);
and U6043 (N_6043,N_606,N_2111);
nor U6044 (N_6044,N_1023,N_557);
nor U6045 (N_6045,N_5994,N_1098);
nand U6046 (N_6046,N_2731,N_5973);
or U6047 (N_6047,N_343,N_3508);
nand U6048 (N_6048,N_1700,N_5996);
nor U6049 (N_6049,N_2645,N_5131);
or U6050 (N_6050,N_5577,N_4200);
and U6051 (N_6051,N_2559,N_3946);
xnor U6052 (N_6052,N_5800,N_2872);
xnor U6053 (N_6053,N_3815,N_5572);
or U6054 (N_6054,N_5755,N_5202);
and U6055 (N_6055,N_3406,N_3152);
nor U6056 (N_6056,N_2729,N_5034);
and U6057 (N_6057,N_3936,N_5813);
xor U6058 (N_6058,N_3294,N_192);
and U6059 (N_6059,N_3990,N_5938);
or U6060 (N_6060,N_4371,N_4289);
and U6061 (N_6061,N_4360,N_1785);
xor U6062 (N_6062,N_5114,N_2713);
or U6063 (N_6063,N_5753,N_1393);
nor U6064 (N_6064,N_4709,N_159);
nand U6065 (N_6065,N_4006,N_1046);
nor U6066 (N_6066,N_1640,N_603);
and U6067 (N_6067,N_5497,N_3389);
nand U6068 (N_6068,N_4960,N_4410);
and U6069 (N_6069,N_4430,N_2244);
xnor U6070 (N_6070,N_1371,N_1192);
or U6071 (N_6071,N_3578,N_4819);
or U6072 (N_6072,N_5157,N_80);
and U6073 (N_6073,N_2692,N_2029);
or U6074 (N_6074,N_5913,N_2711);
or U6075 (N_6075,N_1765,N_518);
nand U6076 (N_6076,N_3428,N_5979);
or U6077 (N_6077,N_4714,N_5730);
nor U6078 (N_6078,N_5410,N_4283);
nand U6079 (N_6079,N_1874,N_4178);
nand U6080 (N_6080,N_1477,N_4119);
and U6081 (N_6081,N_4118,N_5560);
xor U6082 (N_6082,N_5660,N_5392);
or U6083 (N_6083,N_1920,N_1738);
nand U6084 (N_6084,N_3809,N_1457);
and U6085 (N_6085,N_1168,N_3676);
xor U6086 (N_6086,N_4038,N_303);
nand U6087 (N_6087,N_493,N_478);
nand U6088 (N_6088,N_2699,N_638);
and U6089 (N_6089,N_4518,N_1875);
nand U6090 (N_6090,N_5126,N_5568);
nand U6091 (N_6091,N_2039,N_5543);
xnor U6092 (N_6092,N_5437,N_2168);
and U6093 (N_6093,N_2417,N_316);
and U6094 (N_6094,N_3498,N_2595);
nand U6095 (N_6095,N_5872,N_2516);
and U6096 (N_6096,N_4638,N_3314);
and U6097 (N_6097,N_4759,N_3648);
or U6098 (N_6098,N_3257,N_3645);
nand U6099 (N_6099,N_1719,N_5983);
and U6100 (N_6100,N_4886,N_1344);
or U6101 (N_6101,N_4151,N_2779);
nor U6102 (N_6102,N_2331,N_2083);
xor U6103 (N_6103,N_4016,N_30);
and U6104 (N_6104,N_3620,N_591);
xnor U6105 (N_6105,N_361,N_2893);
xnor U6106 (N_6106,N_2243,N_5395);
and U6107 (N_6107,N_4077,N_262);
and U6108 (N_6108,N_1650,N_5304);
nand U6109 (N_6109,N_2439,N_3667);
and U6110 (N_6110,N_996,N_3065);
xor U6111 (N_6111,N_1321,N_3969);
xor U6112 (N_6112,N_2472,N_685);
nor U6113 (N_6113,N_2362,N_521);
nand U6114 (N_6114,N_1065,N_2075);
nor U6115 (N_6115,N_3156,N_4362);
or U6116 (N_6116,N_19,N_2619);
and U6117 (N_6117,N_1367,N_2821);
or U6118 (N_6118,N_1733,N_3222);
nor U6119 (N_6119,N_4885,N_426);
nand U6120 (N_6120,N_597,N_4254);
nor U6121 (N_6121,N_1194,N_4183);
xnor U6122 (N_6122,N_5279,N_2640);
nor U6123 (N_6123,N_3217,N_3573);
and U6124 (N_6124,N_3471,N_2064);
xor U6125 (N_6125,N_3847,N_272);
xor U6126 (N_6126,N_3036,N_3562);
and U6127 (N_6127,N_4433,N_2652);
or U6128 (N_6128,N_4705,N_5659);
and U6129 (N_6129,N_3674,N_541);
nand U6130 (N_6130,N_1561,N_85);
nor U6131 (N_6131,N_2909,N_5622);
nand U6132 (N_6132,N_4521,N_484);
nand U6133 (N_6133,N_2385,N_5581);
or U6134 (N_6134,N_3417,N_5085);
and U6135 (N_6135,N_3841,N_3372);
and U6136 (N_6136,N_5370,N_4003);
or U6137 (N_6137,N_2991,N_4295);
xor U6138 (N_6138,N_4041,N_3541);
or U6139 (N_6139,N_830,N_5842);
nand U6140 (N_6140,N_1860,N_817);
and U6141 (N_6141,N_699,N_1258);
nor U6142 (N_6142,N_4949,N_488);
and U6143 (N_6143,N_1871,N_4064);
xnor U6144 (N_6144,N_553,N_3080);
xnor U6145 (N_6145,N_5701,N_1166);
or U6146 (N_6146,N_5718,N_3866);
and U6147 (N_6147,N_198,N_3731);
xnor U6148 (N_6148,N_302,N_4866);
nand U6149 (N_6149,N_2453,N_3862);
nor U6150 (N_6150,N_1759,N_3386);
and U6151 (N_6151,N_724,N_1642);
and U6152 (N_6152,N_566,N_4161);
or U6153 (N_6153,N_4531,N_2934);
nand U6154 (N_6154,N_1625,N_3017);
xnor U6155 (N_6155,N_542,N_2060);
xnor U6156 (N_6156,N_4600,N_237);
nor U6157 (N_6157,N_3117,N_1979);
nand U6158 (N_6158,N_3773,N_2968);
or U6159 (N_6159,N_4192,N_415);
xnor U6160 (N_6160,N_1278,N_3202);
or U6161 (N_6161,N_3999,N_1357);
xor U6162 (N_6162,N_2093,N_3884);
xnor U6163 (N_6163,N_5048,N_1731);
nand U6164 (N_6164,N_5104,N_3187);
xor U6165 (N_6165,N_633,N_2873);
xnor U6166 (N_6166,N_3244,N_4089);
nor U6167 (N_6167,N_374,N_5781);
nor U6168 (N_6168,N_1697,N_2465);
xnor U6169 (N_6169,N_2343,N_171);
and U6170 (N_6170,N_4498,N_5561);
or U6171 (N_6171,N_5613,N_5633);
or U6172 (N_6172,N_345,N_1974);
xnor U6173 (N_6173,N_1200,N_2723);
and U6174 (N_6174,N_341,N_3338);
nor U6175 (N_6175,N_2862,N_2188);
or U6176 (N_6176,N_4215,N_423);
or U6177 (N_6177,N_2982,N_4144);
nand U6178 (N_6178,N_2267,N_5564);
or U6179 (N_6179,N_5513,N_4884);
or U6180 (N_6180,N_5953,N_4488);
and U6181 (N_6181,N_4617,N_448);
nor U6182 (N_6182,N_2749,N_1245);
or U6183 (N_6183,N_4483,N_5741);
and U6184 (N_6184,N_4844,N_1828);
or U6185 (N_6185,N_964,N_2664);
or U6186 (N_6186,N_1821,N_2178);
nand U6187 (N_6187,N_3913,N_2329);
nand U6188 (N_6188,N_2901,N_4102);
nand U6189 (N_6189,N_5470,N_4861);
or U6190 (N_6190,N_4995,N_3167);
xor U6191 (N_6191,N_3844,N_1063);
nor U6192 (N_6192,N_3531,N_104);
or U6193 (N_6193,N_5522,N_885);
nand U6194 (N_6194,N_2360,N_2120);
nand U6195 (N_6195,N_2826,N_5307);
and U6196 (N_6196,N_1732,N_4288);
and U6197 (N_6197,N_4734,N_5376);
nor U6198 (N_6198,N_326,N_3747);
and U6199 (N_6199,N_3941,N_3004);
or U6200 (N_6200,N_136,N_5076);
xor U6201 (N_6201,N_1350,N_926);
nand U6202 (N_6202,N_2671,N_982);
nor U6203 (N_6203,N_2592,N_1752);
or U6204 (N_6204,N_2969,N_3255);
or U6205 (N_6205,N_5312,N_3213);
nand U6206 (N_6206,N_3169,N_2883);
and U6207 (N_6207,N_460,N_180);
nor U6208 (N_6208,N_1867,N_255);
xor U6209 (N_6209,N_3712,N_2615);
nor U6210 (N_6210,N_3356,N_5285);
or U6211 (N_6211,N_5274,N_2677);
nor U6212 (N_6212,N_2209,N_2925);
and U6213 (N_6213,N_2604,N_3344);
or U6214 (N_6214,N_4052,N_2444);
or U6215 (N_6215,N_3971,N_4865);
and U6216 (N_6216,N_910,N_679);
nor U6217 (N_6217,N_5957,N_2073);
xnor U6218 (N_6218,N_299,N_4991);
and U6219 (N_6219,N_2744,N_1521);
or U6220 (N_6220,N_3566,N_2603);
nand U6221 (N_6221,N_2815,N_5221);
and U6222 (N_6222,N_1348,N_1188);
nand U6223 (N_6223,N_2136,N_2644);
and U6224 (N_6224,N_2222,N_4738);
and U6225 (N_6225,N_3245,N_2551);
xnor U6226 (N_6226,N_4900,N_5419);
xnor U6227 (N_6227,N_5381,N_1147);
nand U6228 (N_6228,N_4787,N_2684);
nand U6229 (N_6229,N_947,N_3120);
xor U6230 (N_6230,N_5489,N_186);
nor U6231 (N_6231,N_5242,N_5071);
nand U6232 (N_6232,N_3820,N_794);
or U6233 (N_6233,N_5615,N_3405);
xnor U6234 (N_6234,N_5394,N_4735);
xor U6235 (N_6235,N_5514,N_4060);
and U6236 (N_6236,N_1659,N_2789);
nor U6237 (N_6237,N_1366,N_1500);
nor U6238 (N_6238,N_766,N_803);
nand U6239 (N_6239,N_2214,N_5565);
nor U6240 (N_6240,N_2771,N_1773);
xnor U6241 (N_6241,N_126,N_111);
nand U6242 (N_6242,N_2981,N_5754);
xor U6243 (N_6243,N_16,N_5592);
and U6244 (N_6244,N_787,N_5123);
and U6245 (N_6245,N_4857,N_1180);
nor U6246 (N_6246,N_4383,N_4814);
or U6247 (N_6247,N_2312,N_2260);
xor U6248 (N_6248,N_3864,N_2910);
and U6249 (N_6249,N_2786,N_3072);
xor U6250 (N_6250,N_4975,N_949);
or U6251 (N_6251,N_381,N_2858);
xor U6252 (N_6252,N_4835,N_3336);
xnor U6253 (N_6253,N_661,N_5607);
or U6254 (N_6254,N_5848,N_4236);
and U6255 (N_6255,N_1895,N_2030);
nor U6256 (N_6256,N_1134,N_4629);
nand U6257 (N_6257,N_2569,N_42);
xor U6258 (N_6258,N_3713,N_833);
nor U6259 (N_6259,N_2919,N_4141);
and U6260 (N_6260,N_1402,N_5125);
nor U6261 (N_6261,N_5344,N_2582);
and U6262 (N_6262,N_2889,N_3759);
and U6263 (N_6263,N_4112,N_3590);
xor U6264 (N_6264,N_3019,N_950);
or U6265 (N_6265,N_1469,N_1717);
xor U6266 (N_6266,N_2258,N_4506);
and U6267 (N_6267,N_5435,N_2738);
xnor U6268 (N_6268,N_1162,N_3381);
nor U6269 (N_6269,N_5492,N_1191);
nor U6270 (N_6270,N_4287,N_2277);
xnor U6271 (N_6271,N_3579,N_655);
and U6272 (N_6272,N_5997,N_2367);
and U6273 (N_6273,N_711,N_3736);
or U6274 (N_6274,N_1049,N_3932);
and U6275 (N_6275,N_2511,N_2053);
nand U6276 (N_6276,N_2674,N_2124);
nand U6277 (N_6277,N_4413,N_1849);
and U6278 (N_6278,N_5473,N_4179);
xor U6279 (N_6279,N_900,N_3730);
or U6280 (N_6280,N_5468,N_5998);
xnor U6281 (N_6281,N_3545,N_2042);
nand U6282 (N_6282,N_2303,N_1337);
nor U6283 (N_6283,N_761,N_1781);
or U6284 (N_6284,N_2947,N_1171);
xor U6285 (N_6285,N_3241,N_2418);
and U6286 (N_6286,N_5706,N_5383);
nand U6287 (N_6287,N_3934,N_4216);
or U6288 (N_6288,N_5610,N_684);
or U6289 (N_6289,N_5057,N_5469);
xor U6290 (N_6290,N_3432,N_580);
nor U6291 (N_6291,N_4123,N_296);
nand U6292 (N_6292,N_2221,N_721);
and U6293 (N_6293,N_2570,N_666);
or U6294 (N_6294,N_1506,N_2212);
nor U6295 (N_6295,N_1532,N_4504);
nand U6296 (N_6296,N_5725,N_1464);
or U6297 (N_6297,N_450,N_3938);
xnor U6298 (N_6298,N_3491,N_267);
or U6299 (N_6299,N_4124,N_598);
and U6300 (N_6300,N_4347,N_1846);
nor U6301 (N_6301,N_5723,N_4019);
xnor U6302 (N_6302,N_4562,N_2700);
nor U6303 (N_6303,N_1019,N_1296);
and U6304 (N_6304,N_1293,N_4166);
or U6305 (N_6305,N_1160,N_147);
xnor U6306 (N_6306,N_4690,N_2491);
nand U6307 (N_6307,N_1185,N_5191);
xor U6308 (N_6308,N_3168,N_1285);
nand U6309 (N_6309,N_3678,N_2422);
and U6310 (N_6310,N_5029,N_4175);
xor U6311 (N_6311,N_120,N_2131);
xor U6312 (N_6312,N_50,N_3523);
nand U6313 (N_6313,N_5775,N_1587);
nor U6314 (N_6314,N_4464,N_3394);
nand U6315 (N_6315,N_1713,N_1341);
nand U6316 (N_6316,N_3619,N_2648);
nand U6317 (N_6317,N_2263,N_801);
xnor U6318 (N_6318,N_3046,N_3570);
nand U6319 (N_6319,N_4936,N_5883);
or U6320 (N_6320,N_97,N_1545);
nor U6321 (N_6321,N_1050,N_5211);
nand U6322 (N_6322,N_625,N_393);
or U6323 (N_6323,N_4270,N_39);
and U6324 (N_6324,N_128,N_1239);
xor U6325 (N_6325,N_5447,N_2252);
xnor U6326 (N_6326,N_3827,N_199);
and U6327 (N_6327,N_1924,N_413);
nor U6328 (N_6328,N_4044,N_5145);
nand U6329 (N_6329,N_5559,N_3391);
and U6330 (N_6330,N_5173,N_148);
nor U6331 (N_6331,N_1220,N_4070);
nand U6332 (N_6332,N_4806,N_4377);
nor U6333 (N_6333,N_3559,N_5758);
or U6334 (N_6334,N_3124,N_2176);
xnor U6335 (N_6335,N_1289,N_1809);
or U6336 (N_6336,N_1503,N_650);
nand U6337 (N_6337,N_607,N_3542);
and U6338 (N_6338,N_1987,N_2330);
xor U6339 (N_6339,N_3829,N_4711);
or U6340 (N_6340,N_2623,N_1858);
nand U6341 (N_6341,N_5964,N_944);
xor U6342 (N_6342,N_1743,N_1433);
and U6343 (N_6343,N_1437,N_3280);
nor U6344 (N_6344,N_3249,N_1042);
and U6345 (N_6345,N_3571,N_116);
and U6346 (N_6346,N_1325,N_4914);
nand U6347 (N_6347,N_912,N_1317);
xnor U6348 (N_6348,N_3096,N_5027);
and U6349 (N_6349,N_3115,N_1658);
and U6350 (N_6350,N_1859,N_3514);
nor U6351 (N_6351,N_1919,N_2798);
nor U6352 (N_6352,N_4284,N_2204);
nand U6353 (N_6353,N_5268,N_360);
and U6354 (N_6354,N_1222,N_4956);
nand U6355 (N_6355,N_4969,N_1323);
nand U6356 (N_6356,N_2276,N_927);
and U6357 (N_6357,N_1078,N_5007);
nand U6358 (N_6358,N_4248,N_4406);
nor U6359 (N_6359,N_5790,N_3282);
nand U6360 (N_6360,N_5729,N_1345);
nand U6361 (N_6361,N_1079,N_2793);
and U6362 (N_6362,N_5089,N_4320);
or U6363 (N_6363,N_1985,N_616);
and U6364 (N_6364,N_3569,N_3808);
or U6365 (N_6365,N_1304,N_1630);
and U6366 (N_6366,N_403,N_742);
nor U6367 (N_6367,N_520,N_3807);
nand U6368 (N_6368,N_2341,N_1699);
or U6369 (N_6369,N_4670,N_4104);
and U6370 (N_6370,N_2555,N_4133);
and U6371 (N_6371,N_3182,N_273);
xor U6372 (N_6372,N_5314,N_4809);
nor U6373 (N_6373,N_5768,N_3921);
xnor U6374 (N_6374,N_443,N_3874);
xor U6375 (N_6375,N_2442,N_2139);
xnor U6376 (N_6376,N_1182,N_5537);
nor U6377 (N_6377,N_4515,N_3146);
or U6378 (N_6378,N_5590,N_5510);
xnor U6379 (N_6379,N_3277,N_3706);
nand U6380 (N_6380,N_3327,N_965);
and U6381 (N_6381,N_5079,N_560);
xnor U6382 (N_6382,N_5937,N_1379);
xnor U6383 (N_6383,N_1568,N_5445);
xor U6384 (N_6384,N_3822,N_3882);
nor U6385 (N_6385,N_4658,N_422);
xor U6386 (N_6386,N_1960,N_1651);
nand U6387 (N_6387,N_758,N_3153);
and U6388 (N_6388,N_3362,N_2262);
nand U6389 (N_6389,N_4240,N_1218);
nor U6390 (N_6390,N_954,N_4692);
xor U6391 (N_6391,N_3918,N_4838);
nand U6392 (N_6392,N_4376,N_2608);
nand U6393 (N_6393,N_5747,N_2661);
nand U6394 (N_6394,N_4720,N_2666);
nor U6395 (N_6395,N_936,N_883);
or U6396 (N_6396,N_3042,N_5733);
nor U6397 (N_6397,N_5069,N_3521);
or U6398 (N_6398,N_4683,N_2187);
nand U6399 (N_6399,N_1173,N_4781);
or U6400 (N_6400,N_1407,N_4204);
xnor U6401 (N_6401,N_290,N_1170);
nor U6402 (N_6402,N_3517,N_5627);
and U6403 (N_6403,N_3640,N_969);
nor U6404 (N_6404,N_1887,N_4108);
xnor U6405 (N_6405,N_442,N_3816);
and U6406 (N_6406,N_4669,N_4940);
nor U6407 (N_6407,N_5358,N_2609);
and U6408 (N_6408,N_2933,N_5283);
nor U6409 (N_6409,N_2346,N_69);
xnor U6410 (N_6410,N_2234,N_4780);
nand U6411 (N_6411,N_4789,N_4996);
nor U6412 (N_6412,N_645,N_1483);
or U6413 (N_6413,N_895,N_1066);
nand U6414 (N_6414,N_1562,N_1963);
xor U6415 (N_6415,N_5111,N_4534);
xnor U6416 (N_6416,N_1312,N_166);
or U6417 (N_6417,N_2750,N_24);
xor U6418 (N_6418,N_4252,N_4769);
nor U6419 (N_6419,N_5263,N_3301);
nand U6420 (N_6420,N_2647,N_5796);
nand U6421 (N_6421,N_3269,N_2502);
nand U6422 (N_6422,N_4313,N_5618);
nand U6423 (N_6423,N_2599,N_2790);
or U6424 (N_6424,N_1115,N_3777);
nand U6425 (N_6425,N_3661,N_3454);
xor U6426 (N_6426,N_3263,N_612);
nor U6427 (N_6427,N_2328,N_2045);
nor U6428 (N_6428,N_5012,N_2732);
nor U6429 (N_6429,N_2780,N_2350);
nor U6430 (N_6430,N_2335,N_2528);
and U6431 (N_6431,N_4667,N_3937);
nand U6432 (N_6432,N_4138,N_5902);
and U6433 (N_6433,N_5856,N_4796);
xor U6434 (N_6434,N_4530,N_4032);
nor U6435 (N_6435,N_1067,N_3433);
or U6436 (N_6436,N_1369,N_4424);
or U6437 (N_6437,N_934,N_5570);
or U6438 (N_6438,N_3016,N_1533);
xnor U6439 (N_6439,N_5525,N_2372);
nor U6440 (N_6440,N_1320,N_3942);
nor U6441 (N_6441,N_5323,N_1363);
and U6442 (N_6442,N_3906,N_5806);
xor U6443 (N_6443,N_5219,N_1252);
xnor U6444 (N_6444,N_710,N_2458);
and U6445 (N_6445,N_3550,N_1275);
and U6446 (N_6446,N_1780,N_2719);
xor U6447 (N_6447,N_894,N_1988);
nor U6448 (N_6448,N_142,N_4625);
nor U6449 (N_6449,N_5788,N_5520);
nor U6450 (N_6450,N_2344,N_205);
and U6451 (N_6451,N_3767,N_977);
nor U6452 (N_6452,N_4004,N_3895);
and U6453 (N_6453,N_1299,N_2411);
or U6454 (N_6454,N_1579,N_867);
nor U6455 (N_6455,N_2205,N_5464);
nand U6456 (N_6456,N_583,N_4674);
nand U6457 (N_6457,N_2043,N_4499);
nor U6458 (N_6458,N_3537,N_3463);
or U6459 (N_6459,N_2690,N_538);
and U6460 (N_6460,N_2435,N_408);
or U6461 (N_6461,N_1029,N_2446);
nand U6462 (N_6462,N_4385,N_138);
xor U6463 (N_6463,N_1032,N_1788);
and U6464 (N_6464,N_5962,N_5932);
or U6465 (N_6465,N_4197,N_2529);
xnor U6466 (N_6466,N_1791,N_1638);
xor U6467 (N_6467,N_3544,N_5137);
and U6468 (N_6468,N_309,N_3141);
nand U6469 (N_6469,N_197,N_4427);
or U6470 (N_6470,N_4905,N_4435);
nor U6471 (N_6471,N_3642,N_2006);
nand U6472 (N_6472,N_5398,N_1853);
nand U6473 (N_6473,N_2832,N_1132);
xor U6474 (N_6474,N_4718,N_2942);
or U6475 (N_6475,N_1766,N_3750);
xnor U6476 (N_6476,N_702,N_2080);
nor U6477 (N_6477,N_2369,N_253);
nand U6478 (N_6478,N_2416,N_3870);
xor U6479 (N_6479,N_1556,N_5443);
or U6480 (N_6480,N_4260,N_5614);
or U6481 (N_6481,N_1081,N_1460);
xor U6482 (N_6482,N_1070,N_4130);
or U6483 (N_6483,N_3125,N_1288);
or U6484 (N_6484,N_3853,N_1361);
and U6485 (N_6485,N_1471,N_975);
or U6486 (N_6486,N_4058,N_3910);
xor U6487 (N_6487,N_4876,N_2876);
xnor U6488 (N_6488,N_5714,N_5337);
nand U6489 (N_6489,N_5326,N_4887);
and U6490 (N_6490,N_3819,N_349);
and U6491 (N_6491,N_2958,N_1549);
or U6492 (N_6492,N_5616,N_3320);
or U6493 (N_6493,N_2642,N_4557);
and U6494 (N_6494,N_1864,N_2479);
nor U6495 (N_6495,N_5282,N_4980);
nor U6496 (N_6496,N_5782,N_848);
xor U6497 (N_6497,N_1260,N_4543);
xor U6498 (N_6498,N_4522,N_2069);
and U6499 (N_6499,N_2879,N_4246);
nand U6500 (N_6500,N_5321,N_3764);
nor U6501 (N_6501,N_3868,N_5192);
or U6502 (N_6502,N_5190,N_4474);
nor U6503 (N_6503,N_763,N_5350);
and U6504 (N_6504,N_1426,N_579);
nor U6505 (N_6505,N_1739,N_3349);
nand U6506 (N_6506,N_1654,N_3281);
and U6507 (N_6507,N_1075,N_3806);
xor U6508 (N_6508,N_5692,N_1940);
nor U6509 (N_6509,N_1877,N_4221);
nor U6510 (N_6510,N_2361,N_5707);
or U6511 (N_6511,N_406,N_5904);
nor U6512 (N_6512,N_5992,N_2097);
xnor U6513 (N_6513,N_1879,N_5456);
or U6514 (N_6514,N_2211,N_1611);
xor U6515 (N_6515,N_5042,N_1085);
nor U6516 (N_6516,N_1905,N_2059);
and U6517 (N_6517,N_2112,N_5648);
nand U6518 (N_6518,N_5955,N_124);
and U6519 (N_6519,N_1836,N_5484);
and U6520 (N_6520,N_333,N_4850);
nor U6521 (N_6521,N_1465,N_4672);
nand U6522 (N_6522,N_2192,N_2795);
xor U6523 (N_6523,N_132,N_515);
and U6524 (N_6524,N_5512,N_3778);
and U6525 (N_6525,N_1164,N_4962);
and U6526 (N_6526,N_1211,N_4400);
or U6527 (N_6527,N_311,N_384);
and U6528 (N_6528,N_5669,N_4457);
and U6529 (N_6529,N_3266,N_2627);
or U6530 (N_6530,N_5231,N_5207);
and U6531 (N_6531,N_4702,N_5906);
or U6532 (N_6532,N_3917,N_701);
nand U6533 (N_6533,N_5884,N_3483);
nand U6534 (N_6534,N_5642,N_2158);
xor U6535 (N_6535,N_5837,N_1909);
and U6536 (N_6536,N_4055,N_2373);
xnor U6537 (N_6537,N_3307,N_807);
or U6538 (N_6538,N_2468,N_800);
nand U6539 (N_6539,N_4957,N_5911);
nor U6540 (N_6540,N_629,N_2743);
or U6541 (N_6541,N_3539,N_3516);
nand U6542 (N_6542,N_4793,N_3961);
nand U6543 (N_6543,N_1394,N_2767);
xor U6544 (N_6544,N_3846,N_2134);
nand U6545 (N_6545,N_2532,N_2945);
nor U6546 (N_6546,N_2510,N_1055);
nand U6547 (N_6547,N_562,N_2712);
or U6548 (N_6548,N_5786,N_388);
nand U6549 (N_6549,N_568,N_1832);
nor U6550 (N_6550,N_2656,N_1362);
or U6551 (N_6551,N_3393,N_5288);
and U6552 (N_6552,N_698,N_3385);
or U6553 (N_6553,N_3987,N_3071);
nor U6554 (N_6554,N_2433,N_5176);
nand U6555 (N_6555,N_4613,N_3518);
and U6556 (N_6556,N_2497,N_1443);
and U6557 (N_6557,N_2586,N_559);
nor U6558 (N_6558,N_1777,N_4921);
nand U6559 (N_6559,N_5115,N_1311);
and U6560 (N_6560,N_458,N_1476);
and U6561 (N_6561,N_4988,N_2784);
and U6562 (N_6562,N_4574,N_3779);
xor U6563 (N_6563,N_4675,N_810);
or U6564 (N_6564,N_2393,N_2906);
xor U6565 (N_6565,N_2023,N_3103);
or U6566 (N_6566,N_3190,N_4441);
or U6567 (N_6567,N_5154,N_3532);
and U6568 (N_6568,N_3059,N_5982);
or U6569 (N_6569,N_169,N_5859);
or U6570 (N_6570,N_5055,N_3479);
xor U6571 (N_6571,N_3948,N_5757);
or U6572 (N_6572,N_4685,N_2695);
nand U6573 (N_6573,N_1324,N_3375);
or U6574 (N_6574,N_5475,N_2368);
or U6575 (N_6575,N_2462,N_2875);
xnor U6576 (N_6576,N_2733,N_3632);
nand U6577 (N_6577,N_4253,N_1490);
xor U6578 (N_6578,N_4460,N_1825);
or U6579 (N_6579,N_4222,N_1400);
and U6580 (N_6580,N_3848,N_3510);
nor U6581 (N_6581,N_2506,N_1048);
or U6582 (N_6582,N_1144,N_5910);
or U6583 (N_6583,N_860,N_5776);
or U6584 (N_6584,N_2899,N_3326);
xnor U6585 (N_6585,N_2633,N_2636);
xor U6586 (N_6586,N_755,N_3488);
nor U6587 (N_6587,N_55,N_4365);
or U6588 (N_6588,N_5159,N_2283);
or U6589 (N_6589,N_3123,N_2709);
and U6590 (N_6590,N_2998,N_1626);
and U6591 (N_6591,N_307,N_1157);
xor U6592 (N_6592,N_2672,N_4001);
or U6593 (N_6593,N_68,N_4007);
xnor U6594 (N_6594,N_3370,N_4306);
xnor U6595 (N_6595,N_3094,N_4205);
nor U6596 (N_6596,N_3401,N_2707);
or U6597 (N_6597,N_5014,N_764);
nor U6598 (N_6598,N_4176,N_4568);
and U6599 (N_6599,N_4338,N_4641);
nand U6600 (N_6600,N_4966,N_176);
and U6601 (N_6601,N_3199,N_2602);
and U6602 (N_6602,N_4618,N_3215);
or U6603 (N_6603,N_5588,N_5060);
xor U6604 (N_6604,N_4853,N_3073);
nor U6605 (N_6605,N_3785,N_4745);
or U6606 (N_6606,N_4367,N_5373);
nand U6607 (N_6607,N_4747,N_5866);
or U6608 (N_6608,N_1380,N_1598);
nand U6609 (N_6609,N_2735,N_3380);
or U6610 (N_6610,N_5254,N_4770);
and U6611 (N_6611,N_1663,N_5942);
or U6612 (N_6612,N_4114,N_1926);
nor U6613 (N_6613,N_1153,N_1196);
xnor U6614 (N_6614,N_5650,N_2840);
xor U6615 (N_6615,N_2870,N_5889);
nor U6616 (N_6616,N_2857,N_4978);
xor U6617 (N_6617,N_258,N_4583);
xor U6618 (N_6618,N_380,N_5466);
or U6619 (N_6619,N_5710,N_3204);
nor U6620 (N_6620,N_2859,N_3223);
and U6621 (N_6621,N_1623,N_2539);
nor U6622 (N_6622,N_5783,N_289);
and U6623 (N_6623,N_5963,N_2268);
and U6624 (N_6624,N_2880,N_4611);
nand U6625 (N_6625,N_1942,N_632);
nor U6626 (N_6626,N_1165,N_1364);
nand U6627 (N_6627,N_1158,N_682);
nand U6628 (N_6628,N_2327,N_5575);
nor U6629 (N_6629,N_293,N_3254);
nand U6630 (N_6630,N_4327,N_4615);
xnor U6631 (N_6631,N_3553,N_3748);
xnor U6632 (N_6632,N_4053,N_3923);
and U6633 (N_6633,N_1424,N_168);
xor U6634 (N_6634,N_5897,N_2971);
or U6635 (N_6635,N_5414,N_3653);
nand U6636 (N_6636,N_2217,N_469);
xor U6637 (N_6637,N_1986,N_452);
nand U6638 (N_6638,N_61,N_1130);
xnor U6639 (N_6639,N_3210,N_3502);
nand U6640 (N_6640,N_1914,N_2658);
and U6641 (N_6641,N_476,N_4535);
and U6642 (N_6642,N_2754,N_1929);
xnor U6643 (N_6643,N_5333,N_2954);
nand U6644 (N_6644,N_5762,N_2553);
nor U6645 (N_6645,N_2694,N_1212);
nor U6646 (N_6646,N_3568,N_3382);
nor U6647 (N_6647,N_1128,N_2641);
nand U6648 (N_6648,N_775,N_3751);
nand U6649 (N_6649,N_4644,N_3384);
xor U6650 (N_6650,N_4343,N_4398);
xor U6651 (N_6651,N_4687,N_3585);
nor U6652 (N_6652,N_5881,N_3130);
and U6653 (N_6653,N_5284,N_4340);
nand U6654 (N_6654,N_1953,N_4392);
and U6655 (N_6655,N_5620,N_38);
xnor U6656 (N_6656,N_3212,N_958);
nor U6657 (N_6657,N_5885,N_2983);
or U6658 (N_6658,N_2871,N_3878);
xor U6659 (N_6659,N_5112,N_740);
nand U6660 (N_6660,N_988,N_4169);
nor U6661 (N_6661,N_4266,N_868);
and U6662 (N_6662,N_5809,N_4707);
or U6663 (N_6663,N_4402,N_5171);
or U6664 (N_6664,N_4815,N_4227);
nor U6665 (N_6665,N_2477,N_5050);
or U6666 (N_6666,N_2950,N_2160);
and U6667 (N_6667,N_5061,N_2034);
xnor U6668 (N_6668,N_2850,N_2062);
nor U6669 (N_6669,N_4831,N_852);
nand U6670 (N_6670,N_2437,N_2781);
or U6671 (N_6671,N_931,N_5397);
or U6672 (N_6672,N_3843,N_3709);
xnor U6673 (N_6673,N_2927,N_5277);
and U6674 (N_6674,N_4247,N_3881);
nand U6675 (N_6675,N_3226,N_516);
xnor U6676 (N_6676,N_1308,N_2740);
and U6677 (N_6677,N_3821,N_4856);
and U6678 (N_6678,N_2492,N_5364);
nand U6679 (N_6679,N_5716,N_1541);
nand U6680 (N_6680,N_3253,N_3784);
nand U6681 (N_6681,N_4142,N_1565);
and U6682 (N_6682,N_726,N_1001);
xnor U6683 (N_6683,N_2232,N_2229);
nand U6684 (N_6684,N_1812,N_4833);
nand U6685 (N_6685,N_3887,N_140);
or U6686 (N_6686,N_4490,N_3663);
xnor U6687 (N_6687,N_5302,N_1125);
nor U6688 (N_6688,N_5486,N_59);
nor U6689 (N_6689,N_1799,N_3834);
nand U6690 (N_6690,N_4357,N_3558);
or U6691 (N_6691,N_3261,N_5476);
xnor U6692 (N_6692,N_5204,N_3089);
nor U6693 (N_6693,N_1039,N_1234);
and U6694 (N_6694,N_5909,N_5148);
xnor U6695 (N_6695,N_1873,N_4134);
nor U6696 (N_6696,N_375,N_1850);
xnor U6697 (N_6697,N_1269,N_4334);
or U6698 (N_6698,N_5210,N_2114);
nand U6699 (N_6699,N_781,N_999);
and U6700 (N_6700,N_1486,N_3614);
nor U6701 (N_6701,N_2384,N_5225);
nor U6702 (N_6702,N_4566,N_2581);
nor U6703 (N_6703,N_1415,N_3462);
xor U6704 (N_6704,N_5794,N_2090);
xnor U6705 (N_6705,N_2294,N_5657);
xor U6706 (N_6706,N_4135,N_5547);
nand U6707 (N_6707,N_4281,N_790);
nor U6708 (N_6708,N_695,N_1183);
xnor U6709 (N_6709,N_5632,N_1305);
xnor U6710 (N_6710,N_4740,N_3933);
nor U6711 (N_6711,N_5743,N_3321);
and U6712 (N_6712,N_1523,N_1845);
or U6713 (N_6713,N_4696,N_3026);
or U6714 (N_6714,N_3533,N_5705);
or U6715 (N_6715,N_5303,N_3126);
nor U6716 (N_6716,N_5539,N_4784);
and U6717 (N_6717,N_2725,N_1110);
nand U6718 (N_6718,N_189,N_2495);
and U6719 (N_6719,N_658,N_3953);
nand U6720 (N_6720,N_4165,N_1383);
or U6721 (N_6721,N_5977,N_984);
xnor U6722 (N_6722,N_2805,N_1428);
nor U6723 (N_6723,N_2593,N_3612);
and U6724 (N_6724,N_5534,N_564);
or U6725 (N_6725,N_4237,N_3977);
and U6726 (N_6726,N_3414,N_953);
xor U6727 (N_6727,N_5477,N_4088);
xnor U6728 (N_6728,N_5968,N_1089);
nor U6729 (N_6729,N_211,N_3165);
xnor U6730 (N_6730,N_5869,N_3097);
or U6731 (N_6731,N_5668,N_4880);
xnor U6732 (N_6732,N_1105,N_5970);
and U6733 (N_6733,N_1491,N_71);
nand U6734 (N_6734,N_1829,N_2941);
or U6735 (N_6735,N_5947,N_3284);
nand U6736 (N_6736,N_92,N_1339);
or U6737 (N_6737,N_1073,N_2100);
xnor U6738 (N_6738,N_1904,N_2403);
or U6739 (N_6739,N_1033,N_4898);
nor U6740 (N_6740,N_5063,N_365);
or U6741 (N_6741,N_753,N_2579);
nor U6742 (N_6742,N_1863,N_5052);
and U6743 (N_6743,N_4632,N_3478);
or U6744 (N_6744,N_2454,N_5871);
and U6745 (N_6745,N_2150,N_4285);
nand U6746 (N_6746,N_3755,N_5899);
nor U6747 (N_6747,N_2811,N_783);
nor U6748 (N_6748,N_1375,N_2606);
nor U6749 (N_6749,N_928,N_4965);
nand U6750 (N_6750,N_3055,N_5402);
nand U6751 (N_6751,N_2311,N_335);
xor U6752 (N_6752,N_5223,N_356);
nand U6753 (N_6753,N_3631,N_4080);
and U6754 (N_6754,N_1585,N_4262);
xor U6755 (N_6755,N_3200,N_231);
or U6756 (N_6756,N_78,N_1354);
nand U6757 (N_6757,N_4732,N_2788);
nor U6758 (N_6758,N_725,N_3400);
or U6759 (N_6759,N_2651,N_716);
and U6760 (N_6760,N_1530,N_690);
or U6761 (N_6761,N_1855,N_3670);
or U6762 (N_6762,N_3770,N_2904);
nand U6763 (N_6763,N_3221,N_4872);
xnor U6764 (N_6764,N_3007,N_703);
nand U6765 (N_6765,N_2696,N_4621);
nand U6766 (N_6766,N_1265,N_919);
nor U6767 (N_6767,N_3980,N_318);
and U6768 (N_6768,N_2796,N_1570);
xor U6769 (N_6769,N_1935,N_3230);
nor U6770 (N_6770,N_5828,N_2336);
nor U6771 (N_6771,N_5612,N_1649);
and U6772 (N_6772,N_5280,N_4700);
or U6773 (N_6773,N_4763,N_4021);
nor U6774 (N_6774,N_3303,N_3850);
or U6775 (N_6775,N_5051,N_315);
xnor U6776 (N_6776,N_510,N_196);
or U6777 (N_6777,N_1210,N_2747);
and U6778 (N_6778,N_2596,N_5432);
nand U6779 (N_6779,N_5067,N_2530);
or U6780 (N_6780,N_2032,N_3095);
and U6781 (N_6781,N_4947,N_4654);
nand U6782 (N_6782,N_1546,N_4684);
xnor U6783 (N_6783,N_153,N_137);
or U6784 (N_6784,N_915,N_2293);
or U6785 (N_6785,N_3184,N_1899);
or U6786 (N_6786,N_269,N_2923);
nand U6787 (N_6787,N_389,N_4847);
and U6788 (N_6788,N_2912,N_1620);
nand U6789 (N_6789,N_3662,N_2518);
nor U6790 (N_6790,N_4069,N_4501);
and U6791 (N_6791,N_4744,N_5164);
and U6792 (N_6792,N_608,N_1106);
nor U6793 (N_6793,N_5328,N_173);
nor U6794 (N_6794,N_1767,N_5645);
nand U6795 (N_6795,N_774,N_1794);
and U6796 (N_6796,N_5608,N_5233);
nand U6797 (N_6797,N_3657,N_2881);
and U6798 (N_6798,N_5686,N_2307);
xor U6799 (N_6799,N_4322,N_1247);
nor U6800 (N_6800,N_4125,N_971);
nor U6801 (N_6801,N_1964,N_32);
nand U6802 (N_6802,N_58,N_1771);
nand U6803 (N_6803,N_2888,N_3877);
nand U6804 (N_6804,N_3185,N_4932);
or U6805 (N_6805,N_5434,N_5200);
or U6806 (N_6806,N_853,N_939);
nor U6807 (N_6807,N_3621,N_1898);
or U6808 (N_6808,N_1249,N_4489);
xor U6809 (N_6809,N_4113,N_170);
nor U6810 (N_6810,N_1610,N_2578);
or U6811 (N_6811,N_108,N_195);
and U6812 (N_6812,N_125,N_3556);
nor U6813 (N_6813,N_1818,N_2597);
or U6814 (N_6814,N_2161,N_355);
and U6815 (N_6815,N_480,N_5980);
xor U6816 (N_6816,N_696,N_1282);
and U6817 (N_6817,N_1664,N_5483);
or U6818 (N_6818,N_4913,N_3749);
or U6819 (N_6819,N_4812,N_1695);
or U6820 (N_6820,N_5722,N_5801);
nand U6821 (N_6821,N_2908,N_529);
or U6822 (N_6822,N_4699,N_2340);
or U6823 (N_6823,N_1906,N_4551);
xnor U6824 (N_6824,N_88,N_5967);
nor U6825 (N_6825,N_411,N_5037);
nor U6826 (N_6826,N_2199,N_4428);
or U6827 (N_6827,N_5339,N_191);
xnor U6828 (N_6828,N_5248,N_62);
nor U6829 (N_6829,N_4773,N_2225);
xnor U6830 (N_6830,N_1880,N_247);
xor U6831 (N_6831,N_5825,N_418);
nand U6832 (N_6832,N_1378,N_100);
and U6833 (N_6833,N_4040,N_4588);
and U6834 (N_6834,N_5766,N_3625);
xor U6835 (N_6835,N_5816,N_3496);
and U6836 (N_6836,N_144,N_1427);
and U6837 (N_6837,N_130,N_1342);
or U6838 (N_6838,N_594,N_310);
nand U6839 (N_6839,N_4239,N_5271);
nor U6840 (N_6840,N_5462,N_5335);
nor U6841 (N_6841,N_648,N_5300);
or U6842 (N_6842,N_1322,N_3580);
xor U6843 (N_6843,N_878,N_4497);
or U6844 (N_6844,N_3431,N_2377);
and U6845 (N_6845,N_3757,N_4487);
xor U6846 (N_6846,N_4764,N_2970);
or U6847 (N_6847,N_271,N_3925);
xnor U6848 (N_6848,N_1502,N_4834);
nor U6849 (N_6849,N_1902,N_974);
nand U6850 (N_6850,N_4024,N_91);
xnor U6851 (N_6851,N_5847,N_735);
nor U6852 (N_6852,N_1068,N_1193);
nor U6853 (N_6853,N_697,N_5481);
nor U6854 (N_6854,N_1684,N_1496);
nor U6855 (N_6855,N_5792,N_3139);
xnor U6856 (N_6856,N_4330,N_1175);
and U6857 (N_6857,N_903,N_972);
nor U6858 (N_6858,N_1934,N_1439);
nor U6859 (N_6859,N_1463,N_5540);
nor U6860 (N_6860,N_5229,N_5155);
or U6861 (N_6861,N_550,N_5704);
or U6862 (N_6862,N_1728,N_5163);
or U6863 (N_6863,N_3206,N_3699);
nand U6864 (N_6864,N_5132,N_2107);
xnor U6865 (N_6865,N_4045,N_1251);
nand U6866 (N_6866,N_978,N_4443);
xnor U6867 (N_6867,N_20,N_1749);
and U6868 (N_6868,N_4444,N_490);
and U6869 (N_6869,N_4332,N_5635);
nor U6870 (N_6870,N_1881,N_1206);
or U6871 (N_6871,N_5971,N_4379);
and U6872 (N_6872,N_4804,N_17);
xnor U6873 (N_6873,N_4279,N_693);
xor U6874 (N_6874,N_4749,N_5676);
xnor U6875 (N_6875,N_4194,N_5212);
or U6876 (N_6876,N_3680,N_5948);
nor U6877 (N_6877,N_3076,N_5199);
xnor U6878 (N_6878,N_4779,N_3291);
and U6879 (N_6879,N_5342,N_5045);
xor U6880 (N_6880,N_4225,N_3836);
nor U6881 (N_6881,N_5152,N_2113);
xor U6882 (N_6882,N_4309,N_5641);
and U6883 (N_6883,N_1597,N_1981);
xnor U6884 (N_6884,N_2323,N_3745);
nor U6885 (N_6885,N_4364,N_5446);
nand U6886 (N_6886,N_2098,N_1154);
xor U6887 (N_6887,N_3396,N_3771);
nand U6888 (N_6888,N_2813,N_2527);
and U6889 (N_6889,N_2070,N_1976);
xor U6890 (N_6890,N_3000,N_2470);
or U6891 (N_6891,N_506,N_3285);
xnor U6892 (N_6892,N_2019,N_1639);
and U6893 (N_6893,N_3903,N_3885);
xnor U6894 (N_6894,N_901,N_1493);
nand U6895 (N_6895,N_1451,N_2935);
or U6896 (N_6896,N_3300,N_4505);
and U6897 (N_6897,N_291,N_5844);
and U6898 (N_6898,N_3131,N_1511);
nor U6899 (N_6899,N_1908,N_1572);
nand U6900 (N_6900,N_2352,N_940);
or U6901 (N_6901,N_4715,N_2755);
and U6902 (N_6902,N_1232,N_193);
and U6903 (N_6903,N_2259,N_1041);
and U6904 (N_6904,N_5128,N_1694);
xnor U6905 (N_6905,N_543,N_2087);
nor U6906 (N_6906,N_1271,N_2966);
or U6907 (N_6907,N_445,N_4299);
xor U6908 (N_6908,N_2013,N_649);
xor U6909 (N_6909,N_5526,N_2917);
nor U6910 (N_6910,N_712,N_3429);
nor U6911 (N_6911,N_3010,N_4154);
xor U6912 (N_6912,N_99,N_2521);
and U6913 (N_6913,N_4561,N_2898);
and U6914 (N_6914,N_5503,N_5124);
xor U6915 (N_6915,N_750,N_2589);
nor U6916 (N_6916,N_2863,N_5987);
xor U6917 (N_6917,N_2794,N_2972);
and U6918 (N_6918,N_834,N_3970);
nor U6919 (N_6919,N_3033,N_4519);
nor U6920 (N_6920,N_4083,N_1080);
nor U6921 (N_6921,N_3112,N_1455);
xor U6922 (N_6922,N_2018,N_4087);
and U6923 (N_6923,N_1886,N_3196);
and U6924 (N_6924,N_1608,N_906);
nor U6925 (N_6925,N_5625,N_3586);
xnor U6926 (N_6926,N_4903,N_181);
xnor U6927 (N_6927,N_4275,N_405);
nand U6928 (N_6928,N_5359,N_5640);
nand U6929 (N_6929,N_5505,N_26);
nor U6930 (N_6930,N_1241,N_5266);
or U6931 (N_6931,N_2358,N_993);
xor U6932 (N_6932,N_5886,N_2721);
nand U6933 (N_6933,N_2654,N_5143);
xnor U6934 (N_6934,N_90,N_3677);
xnor U6935 (N_6935,N_3317,N_4437);
nor U6936 (N_6936,N_1468,N_3922);
nor U6937 (N_6937,N_4303,N_2962);
xor U6938 (N_6938,N_5606,N_1482);
nor U6939 (N_6939,N_704,N_2742);
and U6940 (N_6940,N_5845,N_4681);
xor U6941 (N_6941,N_3021,N_1691);
nor U6942 (N_6942,N_344,N_5208);
and U6943 (N_6943,N_1937,N_676);
nor U6944 (N_6944,N_1434,N_5127);
and U6945 (N_6945,N_932,N_5378);
nor U6946 (N_6946,N_5247,N_4337);
and U6947 (N_6947,N_882,N_881);
nor U6948 (N_6948,N_3835,N_687);
nand U6949 (N_6949,N_2419,N_3377);
or U6950 (N_6950,N_4373,N_3628);
xnor U6951 (N_6951,N_3907,N_5105);
and U6952 (N_6952,N_5735,N_4581);
nand U6953 (N_6953,N_5036,N_4986);
nor U6954 (N_6954,N_18,N_1553);
and U6955 (N_6955,N_1216,N_1999);
xor U6956 (N_6956,N_5879,N_5450);
and U6957 (N_6957,N_4229,N_1036);
and U6958 (N_6958,N_2827,N_4597);
nor U6959 (N_6959,N_3693,N_5129);
and U6960 (N_6960,N_4132,N_5214);
nor U6961 (N_6961,N_2167,N_3660);
nor U6962 (N_6962,N_3461,N_5863);
nor U6963 (N_6963,N_512,N_2844);
nand U6964 (N_6964,N_3739,N_1930);
or U6965 (N_6965,N_2685,N_1614);
nand U6966 (N_6966,N_2503,N_2973);
and U6967 (N_6967,N_1187,N_5502);
nand U6968 (N_6968,N_1189,N_1838);
nor U6969 (N_6969,N_527,N_5135);
xor U6970 (N_6970,N_4668,N_4645);
or U6971 (N_6971,N_3259,N_5004);
nor U6972 (N_6972,N_3775,N_4633);
nor U6973 (N_6973,N_2011,N_2471);
xor U6974 (N_6974,N_409,N_4147);
or U6975 (N_6975,N_4046,N_1725);
nand U6976 (N_6976,N_3335,N_1097);
or U6977 (N_6977,N_1798,N_1550);
nor U6978 (N_6978,N_4808,N_135);
and U6979 (N_6979,N_3003,N_1891);
nor U6980 (N_6980,N_3975,N_1472);
xor U6981 (N_6981,N_5482,N_4025);
or U6982 (N_6982,N_5498,N_5541);
xor U6983 (N_6983,N_957,N_2104);
nand U6984 (N_6984,N_5949,N_2494);
nand U6985 (N_6985,N_5348,N_1410);
nor U6986 (N_6986,N_779,N_1515);
and U6987 (N_6987,N_2004,N_4537);
xor U6988 (N_6988,N_1118,N_1395);
nand U6989 (N_6989,N_5545,N_1571);
nand U6990 (N_6990,N_105,N_2500);
xor U6991 (N_6991,N_248,N_561);
or U6992 (N_6992,N_5626,N_3093);
xor U6993 (N_6993,N_4382,N_3408);
and U6994 (N_6994,N_5822,N_2916);
xnor U6995 (N_6995,N_3469,N_276);
or U6996 (N_6996,N_4232,N_1005);
xnor U6997 (N_6997,N_336,N_961);
nor U6998 (N_6998,N_3232,N_4026);
and U6999 (N_6999,N_2772,N_4817);
or U7000 (N_7000,N_3594,N_1270);
or U7001 (N_7001,N_5715,N_5465);
or U7002 (N_7002,N_3002,N_2254);
nor U7003 (N_7003,N_4257,N_637);
and U7004 (N_7004,N_1108,N_1109);
or U7005 (N_7005,N_5639,N_5250);
and U7006 (N_7006,N_2438,N_5853);
xor U7007 (N_7007,N_3762,N_222);
nor U7008 (N_7008,N_692,N_1783);
nand U7009 (N_7009,N_3800,N_2499);
xnor U7010 (N_7010,N_2275,N_5421);
nor U7011 (N_7011,N_4059,N_4235);
nor U7012 (N_7012,N_2257,N_3487);
xnor U7013 (N_7013,N_4339,N_4264);
xor U7014 (N_7014,N_1217,N_1376);
nand U7015 (N_7015,N_899,N_5934);
xor U7016 (N_7016,N_3627,N_838);
nand U7017 (N_7017,N_628,N_1031);
or U7018 (N_7018,N_4677,N_1813);
or U7019 (N_7019,N_5499,N_5141);
xnor U7020 (N_7020,N_2238,N_1648);
nand U7021 (N_7021,N_1277,N_3791);
or U7022 (N_7022,N_5082,N_185);
xor U7023 (N_7023,N_2428,N_599);
nor U7024 (N_7024,N_4825,N_3982);
xnor U7025 (N_7025,N_3974,N_1564);
nand U7026 (N_7026,N_4917,N_793);
or U7027 (N_7027,N_2717,N_3237);
nor U7028 (N_7028,N_1365,N_2900);
xor U7029 (N_7029,N_5901,N_4015);
and U7030 (N_7030,N_3547,N_4950);
nand U7031 (N_7031,N_2524,N_3248);
xnor U7032 (N_7032,N_2140,N_1910);
or U7033 (N_7033,N_37,N_2734);
xor U7034 (N_7034,N_4701,N_1000);
nand U7035 (N_7035,N_1606,N_5316);
nor U7036 (N_7036,N_1536,N_2223);
and U7037 (N_7037,N_5928,N_5393);
or U7038 (N_7038,N_1388,N_4691);
nor U7039 (N_7039,N_5044,N_2911);
xor U7040 (N_7040,N_2689,N_3047);
xnor U7041 (N_7041,N_1084,N_1274);
nand U7042 (N_7042,N_5571,N_1301);
xor U7043 (N_7043,N_407,N_5361);
xor U7044 (N_7044,N_3655,N_4139);
or U7045 (N_7045,N_3788,N_3083);
or U7046 (N_7046,N_4923,N_362);
or U7047 (N_7047,N_4105,N_1280);
or U7048 (N_7048,N_4766,N_5290);
and U7049 (N_7049,N_5098,N_229);
nor U7050 (N_7050,N_4481,N_1933);
and U7051 (N_7051,N_2653,N_5493);
nand U7052 (N_7052,N_2452,N_4265);
or U7053 (N_7053,N_1655,N_113);
nand U7054 (N_7054,N_2473,N_323);
and U7055 (N_7055,N_329,N_672);
or U7056 (N_7056,N_3805,N_4418);
and U7057 (N_7057,N_5929,N_5724);
xnor U7058 (N_7058,N_1734,N_1473);
xnor U7059 (N_7059,N_3481,N_188);
and U7060 (N_7060,N_331,N_1837);
nand U7061 (N_7061,N_5099,N_154);
xor U7062 (N_7062,N_1436,N_5009);
nand U7063 (N_7063,N_3035,N_3551);
nand U7064 (N_7064,N_2637,N_5255);
or U7065 (N_7065,N_2571,N_1370);
and U7066 (N_7066,N_646,N_1622);
nor U7067 (N_7067,N_1346,N_4048);
nor U7068 (N_7068,N_2874,N_4935);
nand U7069 (N_7069,N_2882,N_4719);
nand U7070 (N_7070,N_4344,N_4249);
nand U7071 (N_7071,N_2,N_1479);
nand U7072 (N_7072,N_4741,N_1143);
xnor U7073 (N_7073,N_4879,N_204);
and U7074 (N_7074,N_457,N_3978);
and U7075 (N_7075,N_5805,N_4432);
or U7076 (N_7076,N_1230,N_5331);
and U7077 (N_7077,N_5336,N_1440);
xnor U7078 (N_7078,N_3935,N_4656);
xor U7079 (N_7079,N_4797,N_1198);
xnor U7080 (N_7080,N_769,N_1231);
or U7081 (N_7081,N_3639,N_1276);
nor U7082 (N_7082,N_3034,N_76);
nand U7083 (N_7083,N_1795,N_228);
and U7084 (N_7084,N_1665,N_1025);
or U7085 (N_7085,N_5780,N_5306);
nor U7086 (N_7086,N_2557,N_1149);
xnor U7087 (N_7087,N_5991,N_1787);
nand U7088 (N_7088,N_187,N_3107);
xor U7089 (N_7089,N_373,N_2314);
nor U7090 (N_7090,N_1438,N_3715);
xnor U7091 (N_7091,N_640,N_671);
xnor U7092 (N_7092,N_5609,N_902);
or U7093 (N_7093,N_5595,N_4614);
or U7094 (N_7094,N_2556,N_304);
or U7095 (N_7095,N_1722,N_183);
and U7096 (N_7096,N_2791,N_2975);
nor U7097 (N_7097,N_2967,N_3926);
nand U7098 (N_7098,N_3271,N_3456);
and U7099 (N_7099,N_3637,N_5583);
xnor U7100 (N_7100,N_2035,N_1461);
xnor U7101 (N_7101,N_3772,N_502);
and U7102 (N_7102,N_2261,N_1802);
and U7103 (N_7103,N_1233,N_2349);
xnor U7104 (N_7104,N_3060,N_3354);
xor U7105 (N_7105,N_5567,N_4346);
or U7106 (N_7106,N_5536,N_3525);
or U7107 (N_7107,N_2071,N_3310);
xor U7108 (N_7108,N_244,N_664);
and U7109 (N_7109,N_4280,N_5763);
xor U7110 (N_7110,N_503,N_4420);
and U7111 (N_7111,N_951,N_1897);
xnor U7112 (N_7112,N_555,N_2849);
or U7113 (N_7113,N_1894,N_5352);
nand U7114 (N_7114,N_5803,N_5011);
xnor U7115 (N_7115,N_943,N_4043);
nor U7116 (N_7116,N_3654,N_4906);
and U7117 (N_7117,N_2048,N_4035);
nor U7118 (N_7118,N_4472,N_879);
nor U7119 (N_7119,N_3052,N_3944);
xnor U7120 (N_7120,N_1653,N_5875);
or U7121 (N_7121,N_1499,N_5940);
and U7122 (N_7122,N_1470,N_4985);
or U7123 (N_7123,N_4120,N_254);
xor U7124 (N_7124,N_2990,N_3268);
xnor U7125 (N_7125,N_1992,N_5319);
and U7126 (N_7126,N_5504,N_5382);
or U7127 (N_7127,N_610,N_350);
xor U7128 (N_7128,N_2626,N_5713);
xnor U7129 (N_7129,N_4195,N_5945);
and U7130 (N_7130,N_3552,N_1952);
or U7131 (N_7131,N_2305,N_4624);
nand U7132 (N_7132,N_3611,N_178);
and U7133 (N_7133,N_4002,N_4937);
xnor U7134 (N_7134,N_2414,N_2322);
or U7135 (N_7135,N_1675,N_930);
nand U7136 (N_7136,N_4622,N_5151);
and U7137 (N_7137,N_1129,N_3851);
nand U7138 (N_7138,N_2031,N_4065);
or U7139 (N_7139,N_4820,N_3366);
or U7140 (N_7140,N_3858,N_2378);
nor U7141 (N_7141,N_2219,N_2002);
and U7142 (N_7142,N_4170,N_2668);
and U7143 (N_7143,N_25,N_357);
or U7144 (N_7144,N_3929,N_4292);
and U7145 (N_7145,N_3053,N_3985);
nand U7146 (N_7146,N_4942,N_5167);
and U7147 (N_7147,N_1911,N_337);
or U7148 (N_7148,N_2228,N_3665);
or U7149 (N_7149,N_3588,N_2833);
and U7150 (N_7150,N_5295,N_5246);
nor U7151 (N_7151,N_4304,N_5656);
nor U7152 (N_7152,N_5080,N_4689);
and U7153 (N_7153,N_5294,N_1492);
xnor U7154 (N_7154,N_2007,N_1368);
nor U7155 (N_7155,N_3460,N_5389);
nor U7156 (N_7156,N_4484,N_468);
and U7157 (N_7157,N_3114,N_4380);
xor U7158 (N_7158,N_1542,N_551);
and U7159 (N_7159,N_4928,N_5106);
xnor U7160 (N_7160,N_317,N_3869);
xnor U7161 (N_7161,N_511,N_3348);
and U7162 (N_7162,N_251,N_1819);
nand U7163 (N_7163,N_1641,N_5257);
nand U7164 (N_7164,N_4173,N_4342);
xor U7165 (N_7165,N_106,N_4027);
or U7166 (N_7166,N_1529,N_4548);
and U7167 (N_7167,N_5406,N_2632);
or U7168 (N_7168,N_744,N_575);
xor U7169 (N_7169,N_4191,N_2078);
nand U7170 (N_7170,N_778,N_446);
nor U7171 (N_7171,N_3079,N_3704);
xnor U7172 (N_7172,N_3189,N_3376);
and U7173 (N_7173,N_2688,N_1297);
or U7174 (N_7174,N_1497,N_200);
and U7175 (N_7175,N_3838,N_4987);
or U7176 (N_7176,N_3957,N_545);
or U7177 (N_7177,N_1975,N_5017);
nor U7178 (N_7178,N_2345,N_3900);
xor U7179 (N_7179,N_3963,N_3360);
nand U7180 (N_7180,N_5230,N_1869);
nand U7181 (N_7181,N_491,N_3451);
nand U7182 (N_7182,N_4852,N_257);
and U7183 (N_7183,N_227,N_1494);
and U7184 (N_7184,N_73,N_2274);
and U7185 (N_7185,N_5409,N_4150);
or U7186 (N_7186,N_5721,N_2299);
xnor U7187 (N_7187,N_4792,N_2659);
nor U7188 (N_7188,N_5508,N_994);
and U7189 (N_7189,N_4612,N_2525);
nor U7190 (N_7190,N_3505,N_3081);
nand U7191 (N_7191,N_4746,N_4540);
and U7192 (N_7192,N_700,N_839);
nand U7193 (N_7193,N_4731,N_4761);
nor U7194 (N_7194,N_1925,N_1581);
or U7195 (N_7195,N_245,N_1576);
or U7196 (N_7196,N_5388,N_1384);
xnor U7197 (N_7197,N_2851,N_1343);
or U7198 (N_7198,N_3861,N_1513);
and U7199 (N_7199,N_2504,N_1862);
or U7200 (N_7200,N_5170,N_1534);
or U7201 (N_7201,N_535,N_2860);
nor U7202 (N_7202,N_2484,N_1047);
xnor U7203 (N_7203,N_2829,N_2572);
nor U7204 (N_7204,N_2817,N_1706);
nand U7205 (N_7205,N_2127,N_5956);
xnor U7206 (N_7206,N_886,N_5047);
or U7207 (N_7207,N_5529,N_2380);
or U7208 (N_7208,N_2839,N_578);
nor U7209 (N_7209,N_1290,N_5415);
nor U7210 (N_7210,N_1770,N_3238);
xnor U7211 (N_7211,N_2132,N_1121);
xnor U7212 (N_7212,N_643,N_604);
nor U7213 (N_7213,N_1475,N_4828);
nor U7214 (N_7214,N_4242,N_4293);
nand U7215 (N_7215,N_3652,N_4593);
nand U7216 (N_7216,N_1647,N_4436);
and U7217 (N_7217,N_3,N_4128);
nand U7218 (N_7218,N_2703,N_4555);
and U7219 (N_7219,N_2853,N_4502);
or U7220 (N_7220,N_5984,N_5667);
and U7221 (N_7221,N_3403,N_51);
xnor U7222 (N_7222,N_4901,N_2386);
nor U7223 (N_7223,N_2041,N_880);
and U7224 (N_7224,N_1262,N_4591);
nor U7225 (N_7225,N_1208,N_1884);
nor U7226 (N_7226,N_5850,N_3104);
or U7227 (N_7227,N_4798,N_3090);
or U7228 (N_7228,N_5460,N_5241);
and U7229 (N_7229,N_5380,N_2977);
and U7230 (N_7230,N_1531,N_3776);
and U7231 (N_7231,N_2306,N_844);
xnor U7232 (N_7232,N_5533,N_438);
nor U7233 (N_7233,N_3708,N_4301);
and U7234 (N_7234,N_23,N_5120);
or U7235 (N_7235,N_5175,N_420);
and U7236 (N_7236,N_4777,N_733);
xor U7237 (N_7237,N_1955,N_3318);
xnor U7238 (N_7238,N_47,N_887);
xnor U7239 (N_7239,N_3814,N_3592);
xor U7240 (N_7240,N_2585,N_5086);
or U7241 (N_7241,N_3208,N_4140);
nor U7242 (N_7242,N_2806,N_160);
nand U7243 (N_7243,N_3956,N_5074);
nand U7244 (N_7244,N_4981,N_4401);
and U7245 (N_7245,N_5327,N_2149);
or U7246 (N_7246,N_2339,N_1382);
nand U7247 (N_7247,N_4952,N_2574);
xor U7248 (N_7248,N_5001,N_2955);
nand U7249 (N_7249,N_1225,N_1435);
or U7250 (N_7250,N_11,N_2288);
nand U7251 (N_7251,N_127,N_366);
xor U7252 (N_7252,N_4943,N_2063);
xnor U7253 (N_7253,N_1116,N_3361);
nand U7254 (N_7254,N_4970,N_5849);
or U7255 (N_7255,N_117,N_5178);
and U7256 (N_7256,N_841,N_3442);
xnor U7257 (N_7257,N_5351,N_225);
nand U7258 (N_7258,N_5039,N_5556);
nand U7259 (N_7259,N_4117,N_431);
and U7260 (N_7260,N_849,N_3995);
nor U7261 (N_7261,N_2146,N_2256);
xor U7262 (N_7262,N_4620,N_2625);
nor U7263 (N_7263,N_2397,N_2426);
or U7264 (N_7264,N_635,N_641);
xor U7265 (N_7265,N_5053,N_3837);
nand U7266 (N_7266,N_5261,N_3754);
and U7267 (N_7267,N_3939,N_4854);
xnor U7268 (N_7268,N_2792,N_1822);
nor U7269 (N_7269,N_1441,N_3888);
and U7270 (N_7270,N_2086,N_5244);
and U7271 (N_7271,N_1526,N_3048);
and U7272 (N_7272,N_653,N_4442);
and U7273 (N_7273,N_1013,N_1021);
or U7274 (N_7274,N_3379,N_4794);
nand U7275 (N_7275,N_536,N_2564);
nor U7276 (N_7276,N_5064,N_4938);
nand U7277 (N_7277,N_4867,N_2101);
or U7278 (N_7278,N_221,N_5569);
xnor U7279 (N_7279,N_1215,N_4399);
nor U7280 (N_7280,N_3276,N_5193);
or U7281 (N_7281,N_5912,N_2478);
xor U7282 (N_7282,N_3717,N_152);
nor U7283 (N_7283,N_5671,N_5452);
nand U7284 (N_7284,N_1682,N_2568);
or U7285 (N_7285,N_617,N_4881);
xnor U7286 (N_7286,N_3302,N_4652);
nand U7287 (N_7287,N_2298,N_5096);
xnor U7288 (N_7288,N_2451,N_2300);
nand U7289 (N_7289,N_3597,N_2535);
nand U7290 (N_7290,N_2848,N_157);
xnor U7291 (N_7291,N_5636,N_4860);
and U7292 (N_7292,N_2961,N_3789);
nand U7293 (N_7293,N_1548,N_5054);
and U7294 (N_7294,N_4743,N_399);
xor U7295 (N_7295,N_2997,N_3191);
nand U7296 (N_7296,N_1683,N_2825);
xor U7297 (N_7297,N_155,N_4994);
xor U7298 (N_7298,N_2822,N_4214);
or U7299 (N_7299,N_2650,N_5049);
nor U7300 (N_7300,N_2762,N_3051);
nand U7301 (N_7301,N_4840,N_4184);
and U7302 (N_7302,N_1372,N_5591);
nand U7303 (N_7303,N_5374,N_1969);
nor U7304 (N_7304,N_3077,N_1801);
and U7305 (N_7305,N_371,N_242);
nor U7306 (N_7306,N_5461,N_2577);
nand U7307 (N_7307,N_4336,N_4211);
nor U7308 (N_7308,N_2948,N_4598);
or U7309 (N_7309,N_3410,N_3500);
or U7310 (N_7310,N_4217,N_351);
or U7311 (N_7311,N_1551,N_862);
or U7312 (N_7312,N_2802,N_4238);
nand U7313 (N_7313,N_4570,N_2172);
or U7314 (N_7314,N_2681,N_4816);
nand U7315 (N_7315,N_5160,N_1993);
nor U7316 (N_7316,N_308,N_601);
and U7317 (N_7317,N_2102,N_884);
nor U7318 (N_7318,N_3413,N_334);
nor U7319 (N_7319,N_1865,N_2391);
nand U7320 (N_7320,N_4762,N_4366);
xnor U7321 (N_7321,N_3192,N_995);
nor U7322 (N_7322,N_1458,N_4174);
nand U7323 (N_7323,N_4586,N_5387);
or U7324 (N_7324,N_1456,N_1102);
and U7325 (N_7325,N_3831,N_4294);
nor U7326 (N_7326,N_1878,N_4325);
or U7327 (N_7327,N_5831,N_1432);
or U7328 (N_7328,N_5385,N_2886);
xnor U7329 (N_7329,N_739,N_4842);
nor U7330 (N_7330,N_2334,N_4298);
nor U7331 (N_7331,N_328,N_3735);
nor U7332 (N_7332,N_3565,N_1951);
or U7333 (N_7333,N_796,N_4983);
nor U7334 (N_7334,N_2541,N_2198);
xor U7335 (N_7335,N_102,N_5893);
xnor U7336 (N_7336,N_3557,N_5066);
or U7337 (N_7337,N_4878,N_5898);
and U7338 (N_7338,N_2493,N_3993);
or U7339 (N_7339,N_2877,N_2926);
and U7340 (N_7340,N_5702,N_5237);
or U7341 (N_7341,N_5480,N_1857);
xor U7342 (N_7342,N_1676,N_991);
nand U7343 (N_7343,N_5506,N_67);
xnor U7344 (N_7344,N_5675,N_3543);
xor U7345 (N_7345,N_5586,N_4152);
nand U7346 (N_7346,N_3387,N_1805);
nor U7347 (N_7347,N_5624,N_1558);
or U7348 (N_7348,N_1735,N_4836);
and U7349 (N_7349,N_4604,N_2548);
xor U7350 (N_7350,N_5785,N_5478);
and U7351 (N_7351,N_1755,N_5717);
xnor U7352 (N_7352,N_5925,N_760);
nor U7353 (N_7353,N_2248,N_5439);
nand U7354 (N_7354,N_358,N_4111);
or U7355 (N_7355,N_2580,N_2807);
xnor U7356 (N_7356,N_2357,N_4508);
xor U7357 (N_7357,N_2705,N_1776);
and U7358 (N_7358,N_5727,N_4724);
nor U7359 (N_7359,N_3626,N_4713);
nor U7360 (N_7360,N_5197,N_997);
nor U7361 (N_7361,N_496,N_4526);
xnor U7362 (N_7362,N_1645,N_2047);
and U7363 (N_7363,N_4233,N_4092);
nor U7364 (N_7364,N_2365,N_3536);
or U7365 (N_7365,N_1389,N_3994);
and U7366 (N_7366,N_5719,N_851);
nand U7367 (N_7367,N_3416,N_1310);
xnor U7368 (N_7368,N_2280,N_5553);
xnor U7369 (N_7369,N_3067,N_727);
or U7370 (N_7370,N_3043,N_2836);
or U7371 (N_7371,N_3863,N_1613);
or U7372 (N_7372,N_4453,N_2544);
or U7373 (N_7373,N_3419,N_1248);
nor U7374 (N_7374,N_876,N_4888);
and U7375 (N_7375,N_4486,N_1715);
or U7376 (N_7376,N_1750,N_3509);
or U7377 (N_7377,N_5764,N_945);
nor U7378 (N_7378,N_729,N_3719);
or U7379 (N_7379,N_3229,N_5950);
and U7380 (N_7380,N_1266,N_1353);
or U7381 (N_7381,N_2768,N_2965);
xnor U7382 (N_7382,N_1294,N_5558);
and U7383 (N_7383,N_3698,N_1600);
xor U7384 (N_7384,N_4354,N_2628);
nor U7385 (N_7385,N_84,N_544);
or U7386 (N_7386,N_2993,N_5923);
and U7387 (N_7387,N_1257,N_2629);
or U7388 (N_7388,N_4079,N_4425);
and U7389 (N_7389,N_2342,N_391);
nor U7390 (N_7390,N_5978,N_1174);
and U7391 (N_7391,N_2847,N_1002);
nand U7392 (N_7392,N_3683,N_2155);
or U7393 (N_7393,N_1061,N_656);
nand U7394 (N_7394,N_1412,N_385);
nor U7395 (N_7395,N_2142,N_1604);
nand U7396 (N_7396,N_4312,N_1679);
and U7397 (N_7397,N_2036,N_4491);
nand U7398 (N_7398,N_4572,N_630);
and U7399 (N_7399,N_3465,N_1421);
nand U7400 (N_7400,N_652,N_3044);
nand U7401 (N_7401,N_3066,N_3273);
nor U7402 (N_7402,N_167,N_3293);
xor U7403 (N_7403,N_4209,N_4989);
or U7404 (N_7404,N_115,N_1751);
nor U7405 (N_7405,N_3435,N_624);
and U7406 (N_7406,N_3528,N_5253);
or U7407 (N_7407,N_1786,N_2770);
and U7408 (N_7408,N_4272,N_1796);
xor U7409 (N_7409,N_4635,N_1027);
xor U7410 (N_7410,N_2509,N_5862);
and U7411 (N_7411,N_4094,N_33);
nand U7412 (N_7412,N_3673,N_5638);
xnor U7413 (N_7413,N_2116,N_4871);
and U7414 (N_7414,N_2987,N_677);
or U7415 (N_7415,N_4698,N_5664);
and U7416 (N_7416,N_582,N_3209);
xor U7417 (N_7417,N_3669,N_2175);
or U7418 (N_7418,N_4890,N_590);
or U7419 (N_7419,N_818,N_2759);
or U7420 (N_7420,N_1139,N_577);
nor U7421 (N_7421,N_2646,N_1745);
nor U7422 (N_7422,N_1936,N_3172);
and U7423 (N_7423,N_4899,N_3493);
nor U7424 (N_7424,N_1632,N_4874);
nand U7425 (N_7425,N_3024,N_1035);
xor U7426 (N_7426,N_1092,N_4997);
and U7427 (N_7427,N_499,N_3439);
nor U7428 (N_7428,N_5436,N_5981);
or U7429 (N_7429,N_5062,N_2943);
nor U7430 (N_7430,N_1474,N_2460);
or U7431 (N_7431,N_4356,N_175);
xnor U7432 (N_7432,N_2022,N_3346);
or U7433 (N_7433,N_2241,N_2110);
or U7434 (N_7434,N_5891,N_4116);
or U7435 (N_7435,N_5140,N_613);
or U7436 (N_7436,N_4573,N_4520);
nor U7437 (N_7437,N_683,N_921);
nand U7438 (N_7438,N_2106,N_3839);
nor U7439 (N_7439,N_3595,N_3087);
and U7440 (N_7440,N_3651,N_2105);
nand U7441 (N_7441,N_1689,N_822);
xor U7442 (N_7442,N_3220,N_2395);
and U7443 (N_7443,N_5585,N_5289);
xor U7444 (N_7444,N_5854,N_5602);
nand U7445 (N_7445,N_1315,N_5812);
and U7446 (N_7446,N_2203,N_871);
xor U7447 (N_7447,N_4394,N_5416);
xnor U7448 (N_7448,N_4627,N_2239);
xor U7449 (N_7449,N_5213,N_4137);
or U7450 (N_7450,N_4585,N_4028);
xnor U7451 (N_7451,N_2354,N_2988);
and U7452 (N_7452,N_5357,N_2841);
nand U7453 (N_7453,N_5855,N_5273);
xor U7454 (N_7454,N_1961,N_3707);
and U7455 (N_7455,N_854,N_1619);
and U7456 (N_7456,N_4296,N_3420);
nor U7457 (N_7457,N_1338,N_312);
and U7458 (N_7458,N_2995,N_367);
or U7459 (N_7459,N_2563,N_2046);
or U7460 (N_7460,N_2000,N_492);
nand U7461 (N_7461,N_4776,N_1893);
xor U7462 (N_7462,N_5299,N_4438);
nand U7463 (N_7463,N_4845,N_5058);
nand U7464 (N_7464,N_4115,N_4915);
and U7465 (N_7465,N_2823,N_2714);
or U7466 (N_7466,N_2200,N_5681);
nand U7467 (N_7467,N_1629,N_1429);
xor U7468 (N_7468,N_2600,N_4333);
nand U7469 (N_7469,N_4411,N_1508);
xnor U7470 (N_7470,N_3554,N_4967);
xor U7471 (N_7471,N_3890,N_5516);
and U7472 (N_7472,N_4589,N_4929);
xor U7473 (N_7473,N_4085,N_2054);
xnor U7474 (N_7474,N_416,N_49);
xnor U7475 (N_7475,N_4431,N_2309);
xnor U7476 (N_7476,N_2830,N_2490);
nand U7477 (N_7477,N_3871,N_5690);
xnor U7478 (N_7478,N_27,N_2769);
nor U7479 (N_7479,N_546,N_1971);
or U7480 (N_7480,N_5549,N_4029);
nand U7481 (N_7481,N_1916,N_5726);
nand U7482 (N_7482,N_3061,N_1152);
and U7483 (N_7483,N_898,N_1313);
nor U7484 (N_7484,N_4664,N_1179);
or U7485 (N_7485,N_4931,N_5038);
xnor U7486 (N_7486,N_623,N_281);
nor U7487 (N_7487,N_4063,N_1698);
nand U7488 (N_7488,N_4993,N_383);
or U7489 (N_7489,N_4274,N_2605);
xnor U7490 (N_7490,N_5939,N_525);
nand U7491 (N_7491,N_3058,N_1268);
nor U7492 (N_7492,N_3390,N_2279);
nand U7493 (N_7493,N_1712,N_4823);
and U7494 (N_7494,N_1807,N_3880);
nor U7495 (N_7495,N_1711,N_4538);
xnor U7496 (N_7496,N_893,N_4859);
and U7497 (N_7497,N_1763,N_2076);
and U7498 (N_7498,N_5914,N_5777);
nor U7499 (N_7499,N_5087,N_5296);
nor U7500 (N_7500,N_1505,N_5824);
nor U7501 (N_7501,N_2905,N_1254);
nand U7502 (N_7502,N_855,N_3176);
nor U7503 (N_7503,N_524,N_4186);
xnor U7504 (N_7504,N_1704,N_2885);
or U7505 (N_7505,N_2179,N_846);
nand U7506 (N_7506,N_3472,N_3549);
nand U7507 (N_7507,N_1076,N_2182);
xnor U7508 (N_7508,N_3599,N_5005);
nor U7509 (N_7509,N_5025,N_4255);
nor U7510 (N_7510,N_3175,N_3622);
and U7511 (N_7511,N_4933,N_4671);
xnor U7512 (N_7512,N_2552,N_2540);
or U7513 (N_7513,N_2752,N_376);
and U7514 (N_7514,N_4811,N_2242);
nor U7515 (N_7515,N_1983,N_918);
nor U7516 (N_7516,N_4910,N_3955);
nor U7517 (N_7517,N_4047,N_4596);
xor U7518 (N_7518,N_3609,N_5739);
nand U7519 (N_7519,N_811,N_3450);
or U7520 (N_7520,N_5917,N_5043);
nor U7521 (N_7521,N_241,N_2890);
and U7522 (N_7522,N_1943,N_3718);
and U7523 (N_7523,N_1670,N_809);
nand U7524 (N_7524,N_2315,N_4529);
xor U7525 (N_7525,N_4451,N_5329);
xor U7526 (N_7526,N_4228,N_718);
or U7527 (N_7527,N_2431,N_3070);
or U7528 (N_7528,N_3883,N_5926);
xnor U7529 (N_7529,N_1635,N_3705);
or U7530 (N_7530,N_353,N_4619);
nand U7531 (N_7531,N_5400,N_2119);
or U7532 (N_7532,N_3924,N_4708);
and U7533 (N_7533,N_1004,N_1397);
nor U7534 (N_7534,N_3475,N_840);
nor U7535 (N_7535,N_897,N_765);
nor U7536 (N_7536,N_1008,N_4594);
xnor U7537 (N_7537,N_3912,N_213);
xnor U7538 (N_7538,N_3174,N_1467);
xor U7539 (N_7539,N_2099,N_3548);
nor U7540 (N_7540,N_134,N_4999);
nand U7541 (N_7541,N_3520,N_3031);
nand U7542 (N_7542,N_53,N_4471);
nor U7543 (N_7543,N_5338,N_3965);
and U7544 (N_7544,N_1810,N_447);
nor U7545 (N_7545,N_3132,N_2701);
and U7546 (N_7546,N_72,N_3501);
nand U7547 (N_7547,N_1578,N_3600);
and U7548 (N_7548,N_3515,N_5310);
or U7549 (N_7549,N_324,N_5276);
and U7550 (N_7550,N_3716,N_322);
xnor U7551 (N_7551,N_3983,N_5574);
xnor U7552 (N_7552,N_1199,N_660);
nand U7553 (N_7553,N_5839,N_1844);
or U7554 (N_7554,N_1145,N_866);
nor U7555 (N_7555,N_2304,N_3140);
and U7556 (N_7556,N_5224,N_3793);
xor U7557 (N_7557,N_4,N_3011);
nor U7558 (N_7558,N_5411,N_209);
nand U7559 (N_7559,N_465,N_5467);
or U7560 (N_7560,N_4352,N_539);
or U7561 (N_7561,N_4528,N_1656);
nand U7562 (N_7562,N_2456,N_5611);
or U7563 (N_7563,N_2907,N_3582);
and U7564 (N_7564,N_1117,N_1069);
nand U7565 (N_7565,N_1334,N_5699);
nand U7566 (N_7566,N_5315,N_2513);
xor U7567 (N_7567,N_2940,N_3418);
or U7568 (N_7568,N_4454,N_3084);
and U7569 (N_7569,N_2611,N_1811);
or U7570 (N_7570,N_12,N_4909);
or U7571 (N_7571,N_3799,N_5852);
nor U7572 (N_7572,N_3920,N_4889);
and U7573 (N_7573,N_2321,N_631);
or U7574 (N_7574,N_4758,N_4243);
and U7575 (N_7575,N_1416,N_3572);
nor U7576 (N_7576,N_453,N_5552);
nor U7577 (N_7577,N_2240,N_1883);
and U7578 (N_7578,N_2326,N_2612);
or U7579 (N_7579,N_1053,N_1409);
nand U7580 (N_7580,N_1815,N_808);
and U7581 (N_7581,N_5860,N_2383);
xnor U7582 (N_7582,N_95,N_5815);
nand U7583 (N_7583,N_4647,N_908);
xor U7584 (N_7584,N_799,N_4558);
xor U7585 (N_7585,N_2820,N_3763);
and U7586 (N_7586,N_4896,N_4951);
nor U7587 (N_7587,N_2173,N_5002);
xnor U7588 (N_7588,N_836,N_1240);
or U7589 (N_7589,N_1028,N_5746);
or U7590 (N_7590,N_1178,N_5779);
and U7591 (N_7591,N_3650,N_3485);
xnor U7592 (N_7592,N_2519,N_1259);
and U7593 (N_7593,N_2757,N_966);
nor U7594 (N_7594,N_4984,N_1340);
nor U7595 (N_7595,N_1177,N_5652);
nand U7596 (N_7596,N_5405,N_5930);
and U7597 (N_7597,N_1480,N_397);
or U7598 (N_7598,N_5680,N_2929);
xnor U7599 (N_7599,N_585,N_219);
or U7600 (N_7600,N_1405,N_2014);
and U7601 (N_7601,N_4386,N_4467);
nand U7602 (N_7602,N_2224,N_4075);
or U7603 (N_7603,N_133,N_4507);
nor U7604 (N_7604,N_3796,N_1113);
and U7605 (N_7605,N_4930,N_2607);
and U7606 (N_7606,N_4968,N_832);
nor U7607 (N_7607,N_2180,N_4463);
and U7608 (N_7608,N_5220,N_454);
xor U7609 (N_7609,N_1088,N_2399);
nand U7610 (N_7610,N_1690,N_417);
nand U7611 (N_7611,N_372,N_5396);
nand U7612 (N_7612,N_4305,N_432);
or U7613 (N_7613,N_1779,N_1612);
xor U7614 (N_7614,N_1444,N_4801);
xor U7615 (N_7615,N_5107,N_4010);
nand U7616 (N_7616,N_4190,N_4199);
xor U7617 (N_7617,N_1527,N_4578);
and U7618 (N_7618,N_2084,N_618);
and U7619 (N_7619,N_4512,N_979);
nor U7620 (N_7620,N_1687,N_2763);
and U7621 (N_7621,N_1758,N_3250);
and U7622 (N_7622,N_5999,N_5218);
xor U7623 (N_7623,N_2270,N_2208);
or U7624 (N_7624,N_2837,N_425);
nor U7625 (N_7625,N_2049,N_5820);
and U7626 (N_7626,N_4728,N_747);
nand U7627 (N_7627,N_4539,N_3618);
nor U7628 (N_7628,N_3899,N_5922);
xor U7629 (N_7629,N_3295,N_3897);
nand U7630 (N_7630,N_2894,N_3703);
nor U7631 (N_7631,N_3889,N_2020);
and U7632 (N_7632,N_3643,N_2253);
xnor U7633 (N_7633,N_4220,N_3328);
xor U7634 (N_7634,N_275,N_28);
nor U7635 (N_7635,N_1644,N_1418);
or U7636 (N_7636,N_4106,N_3973);
nand U7637 (N_7637,N_5070,N_4642);
xor U7638 (N_7638,N_5630,N_4158);
and U7639 (N_7639,N_4922,N_4640);
or U7640 (N_7640,N_5767,N_3353);
nand U7641 (N_7641,N_4829,N_4757);
nor U7642 (N_7642,N_2687,N_819);
or U7643 (N_7643,N_2251,N_4076);
nor U7644 (N_7644,N_5311,N_295);
nand U7645 (N_7645,N_2507,N_4091);
and U7646 (N_7646,N_3761,N_5637);
or U7647 (N_7647,N_390,N_1335);
nand U7648 (N_7648,N_3830,N_3758);
nand U7649 (N_7649,N_2920,N_2939);
nor U7650 (N_7650,N_1207,N_2001);
nand U7651 (N_7651,N_1602,N_1772);
nand U7652 (N_7652,N_5454,N_3945);
or U7653 (N_7653,N_5156,N_1723);
xor U7654 (N_7654,N_3804,N_5895);
or U7655 (N_7655,N_2056,N_2404);
nand U7656 (N_7656,N_5920,N_3658);
nor U7657 (N_7657,N_3952,N_379);
and U7658 (N_7658,N_5198,N_5550);
nand U7659 (N_7659,N_3159,N_1107);
xnor U7660 (N_7660,N_1668,N_1074);
nor U7661 (N_7661,N_4318,N_4185);
or U7662 (N_7662,N_5679,N_5772);
or U7663 (N_7663,N_3603,N_1103);
and U7664 (N_7664,N_2523,N_4503);
xor U7665 (N_7665,N_2682,N_1024);
nand U7666 (N_7666,N_3527,N_4822);
nor U7667 (N_7667,N_440,N_2079);
xnor U7668 (N_7668,N_2590,N_1716);
and U7669 (N_7669,N_1669,N_2549);
nor U7670 (N_7670,N_41,N_5102);
nand U7671 (N_7671,N_4721,N_5774);
nand U7672 (N_7672,N_738,N_1006);
xor U7673 (N_7673,N_4908,N_1126);
xnor U7674 (N_7674,N_1003,N_5236);
and U7675 (N_7675,N_2936,N_5507);
xnor U7676 (N_7676,N_1250,N_79);
xor U7677 (N_7677,N_5834,N_485);
or U7678 (N_7678,N_4609,N_2068);
xor U7679 (N_7679,N_2560,N_3615);
xnor U7680 (N_7680,N_2408,N_1072);
and U7681 (N_7681,N_2622,N_4767);
xnor U7682 (N_7682,N_3161,N_2138);
nor U7683 (N_7683,N_101,N_1195);
and U7684 (N_7684,N_2038,N_1591);
or U7685 (N_7685,N_1892,N_730);
nand U7686 (N_7686,N_828,N_2135);
nor U7687 (N_7687,N_4639,N_5243);
and U7688 (N_7688,N_5698,N_1255);
and U7689 (N_7689,N_2202,N_202);
or U7690 (N_7690,N_762,N_3753);
and U7691 (N_7691,N_3512,N_1386);
or U7692 (N_7692,N_4369,N_3701);
xor U7693 (N_7693,N_3943,N_4592);
nor U7694 (N_7694,N_3604,N_4391);
nand U7695 (N_7695,N_2928,N_3101);
xnor U7696 (N_7696,N_4582,N_2423);
and U7697 (N_7697,N_5826,N_3555);
or U7698 (N_7698,N_3790,N_3049);
nor U7699 (N_7699,N_2420,N_2545);
nor U7700 (N_7700,N_3144,N_1038);
nand U7701 (N_7701,N_4959,N_513);
and U7702 (N_7702,N_2670,N_2865);
xnor U7703 (N_7703,N_3567,N_1761);
nand U7704 (N_7704,N_4477,N_2634);
and U7705 (N_7705,N_5995,N_172);
xnor U7706 (N_7706,N_5654,N_1332);
nand U7707 (N_7707,N_5150,N_215);
and U7708 (N_7708,N_352,N_5161);
nor U7709 (N_7709,N_410,N_1927);
xnor U7710 (N_7710,N_428,N_609);
nor U7711 (N_7711,N_4973,N_639);
xnor U7712 (N_7712,N_163,N_4446);
or U7713 (N_7713,N_5142,N_3722);
or U7714 (N_7714,N_517,N_627);
nand U7715 (N_7715,N_284,N_891);
nand U7716 (N_7716,N_5116,N_252);
or U7717 (N_7717,N_2594,N_4659);
nor U7718 (N_7718,N_3272,N_1709);
xor U7719 (N_7719,N_4657,N_378);
xor U7720 (N_7720,N_2164,N_850);
nor U7721 (N_7721,N_2374,N_4329);
and U7722 (N_7722,N_5597,N_238);
nor U7723 (N_7723,N_5081,N_4056);
xor U7724 (N_7724,N_773,N_5598);
or U7725 (N_7725,N_4891,N_2631);
or U7726 (N_7726,N_3085,N_3968);
nand U7727 (N_7727,N_1186,N_5709);
xor U7728 (N_7728,N_1417,N_2550);
and U7729 (N_7729,N_1347,N_1034);
xnor U7730 (N_7730,N_3319,N_1430);
nand U7731 (N_7731,N_3351,N_54);
xor U7732 (N_7732,N_1861,N_4754);
or U7733 (N_7733,N_1082,N_1127);
nor U7734 (N_7734,N_2115,N_1244);
xnor U7735 (N_7735,N_843,N_1122);
nand U7736 (N_7736,N_4155,N_856);
xnor U7737 (N_7737,N_2785,N_1124);
or U7738 (N_7738,N_5663,N_5496);
xor U7739 (N_7739,N_5678,N_5172);
xnor U7740 (N_7740,N_4868,N_1917);
xnor U7741 (N_7741,N_3729,N_820);
xor U7742 (N_7742,N_3236,N_4608);
and U7743 (N_7743,N_4736,N_3915);
and U7744 (N_7744,N_3818,N_2797);
and U7745 (N_7745,N_66,N_4396);
or U7746 (N_7746,N_3581,N_5309);
nor U7747 (N_7747,N_3267,N_2867);
or U7748 (N_7748,N_4245,N_4542);
xnor U7749 (N_7749,N_2845,N_5252);
nand U7750 (N_7750,N_1702,N_1577);
nand U7751 (N_7751,N_1509,N_5646);
xnor U7752 (N_7752,N_4415,N_35);
or U7753 (N_7753,N_3534,N_5770);
nor U7754 (N_7754,N_1086,N_5472);
nand U7755 (N_7755,N_354,N_5974);
nand U7756 (N_7756,N_5162,N_5523);
or U7757 (N_7757,N_5092,N_5267);
xnor U7758 (N_7758,N_5169,N_937);
xnor U7759 (N_7759,N_4404,N_2376);
and U7760 (N_7760,N_3598,N_2573);
xnor U7761 (N_7761,N_4213,N_4034);
nor U7762 (N_7762,N_1309,N_400);
nor U7763 (N_7763,N_741,N_297);
nand U7764 (N_7764,N_2673,N_976);
nor U7765 (N_7765,N_1316,N_4830);
nand U7766 (N_7766,N_1775,N_5787);
xor U7767 (N_7767,N_3728,N_473);
nor U7768 (N_7768,N_4841,N_4826);
nand U7769 (N_7769,N_4785,N_694);
and U7770 (N_7770,N_4423,N_3352);
nand U7771 (N_7771,N_2388,N_9);
nand U7772 (N_7772,N_5959,N_1729);
nor U7773 (N_7773,N_3194,N_1966);
xor U7774 (N_7774,N_4291,N_2683);
and U7775 (N_7775,N_4810,N_5563);
and U7776 (N_7776,N_1197,N_43);
nand U7777 (N_7777,N_4071,N_3113);
and U7778 (N_7778,N_4556,N_459);
and U7779 (N_7779,N_909,N_2715);
nor U7780 (N_7780,N_1256,N_4547);
and U7781 (N_7781,N_4258,N_4465);
nand U7782 (N_7782,N_4409,N_4448);
xnor U7783 (N_7783,N_1381,N_1701);
or U7784 (N_7784,N_489,N_1520);
nor U7785 (N_7785,N_2347,N_230);
and U7786 (N_7786,N_4466,N_5371);
and U7787 (N_7787,N_858,N_483);
and U7788 (N_7788,N_3905,N_1017);
nor U7789 (N_7789,N_3813,N_4496);
and U7790 (N_7790,N_1120,N_2691);
nand U7791 (N_7791,N_369,N_3696);
nor U7792 (N_7792,N_1677,N_5961);
nor U7793 (N_7793,N_2215,N_5360);
nand U7794 (N_7794,N_1628,N_3260);
or U7795 (N_7795,N_2005,N_904);
and U7796 (N_7796,N_1095,N_5108);
or U7797 (N_7797,N_3960,N_3499);
or U7798 (N_7798,N_1872,N_5451);
or U7799 (N_7799,N_935,N_347);
and U7800 (N_7800,N_5186,N_2089);
nand U7801 (N_7801,N_4412,N_3015);
or U7802 (N_7802,N_1662,N_2565);
nor U7803 (N_7803,N_1408,N_708);
nand U7804 (N_7804,N_3438,N_2986);
or U7805 (N_7805,N_5020,N_3468);
nand U7806 (N_7806,N_4449,N_3252);
and U7807 (N_7807,N_3275,N_4753);
xor U7808 (N_7808,N_3492,N_75);
xor U7809 (N_7809,N_5966,N_232);
and U7810 (N_7810,N_3181,N_5749);
or U7811 (N_7811,N_3506,N_4131);
xnor U7812 (N_7812,N_3448,N_3812);
xnor U7813 (N_7813,N_2265,N_3287);
nand U7814 (N_7814,N_5101,N_2739);
and U7815 (N_7815,N_110,N_1793);
xnor U7816 (N_7816,N_182,N_4022);
or U7817 (N_7817,N_3009,N_3404);
nand U7818 (N_7818,N_2302,N_3865);
and U7819 (N_7819,N_785,N_825);
nand U7820 (N_7820,N_1939,N_589);
nor U7821 (N_7821,N_600,N_3298);
and U7822 (N_7822,N_2855,N_3892);
nor U7823 (N_7823,N_2727,N_2117);
nor U7824 (N_7824,N_5649,N_5528);
nand U7825 (N_7825,N_3014,N_4136);
or U7826 (N_7826,N_5740,N_313);
xor U7827 (N_7827,N_4739,N_4727);
and U7828 (N_7828,N_5494,N_2808);
nand U7829 (N_7829,N_13,N_2974);
xor U7830 (N_7830,N_1817,N_2407);
and U7831 (N_7831,N_3459,N_4100);
xor U7832 (N_7832,N_2009,N_1990);
and U7833 (N_7833,N_4948,N_1890);
nor U7834 (N_7834,N_5118,N_497);
xor U7835 (N_7835,N_4651,N_4851);
or U7836 (N_7836,N_647,N_1609);
nor U7837 (N_7837,N_1060,N_2774);
nand U7838 (N_7838,N_2103,N_264);
xnor U7839 (N_7839,N_859,N_4145);
xor U7840 (N_7840,N_4939,N_2095);
and U7841 (N_7841,N_4964,N_5330);
or U7842 (N_7842,N_2698,N_2753);
xnor U7843 (N_7843,N_370,N_567);
or U7844 (N_7844,N_5677,N_5298);
or U7845 (N_7845,N_2866,N_4348);
or U7846 (N_7846,N_4974,N_532);
xnor U7847 (N_7847,N_4149,N_705);
nor U7848 (N_7848,N_1286,N_4223);
and U7849 (N_7849,N_131,N_3193);
and U7850 (N_7850,N_615,N_4480);
xor U7851 (N_7851,N_114,N_1119);
or U7852 (N_7852,N_1291,N_620);
and U7853 (N_7853,N_4926,N_857);
nor U7854 (N_7854,N_689,N_5349);
or U7855 (N_7855,N_2130,N_1720);
or U7856 (N_7856,N_2177,N_5532);
xnor U7857 (N_7857,N_4316,N_4290);
nand U7858 (N_7858,N_5068,N_3466);
xor U7859 (N_7859,N_2702,N_1718);
nand U7860 (N_7860,N_2635,N_4307);
nand U7861 (N_7861,N_1949,N_1261);
nor U7862 (N_7862,N_5292,N_3584);
xnor U7863 (N_7863,N_1094,N_4818);
nand U7864 (N_7864,N_5463,N_2736);
nand U7865 (N_7865,N_4726,N_4384);
xor U7866 (N_7866,N_2109,N_3546);
nor U7867 (N_7867,N_4434,N_3309);
nand U7868 (N_7868,N_4167,N_2371);
xor U7869 (N_7869,N_1298,N_2708);
nor U7870 (N_7870,N_1014,N_3412);
and U7871 (N_7871,N_3898,N_4234);
xor U7872 (N_7872,N_1141,N_2675);
or U7873 (N_7873,N_5194,N_2122);
xnor U7874 (N_7874,N_5095,N_2324);
and U7875 (N_7875,N_3426,N_4807);
nor U7876 (N_7876,N_3798,N_5235);
nand U7877 (N_7877,N_3324,N_4549);
or U7878 (N_7878,N_929,N_5694);
and U7879 (N_7879,N_2237,N_1201);
and U7880 (N_7880,N_5935,N_3179);
nor U7881 (N_7881,N_268,N_282);
xor U7882 (N_7882,N_3490,N_3823);
and U7883 (N_7883,N_359,N_1596);
xnor U7884 (N_7884,N_767,N_3737);
xnor U7885 (N_7885,N_4911,N_4122);
xor U7886 (N_7886,N_1059,N_1764);
nor U7887 (N_7887,N_5287,N_4321);
xnor U7888 (N_7888,N_4074,N_4082);
xor U7889 (N_7889,N_2318,N_1104);
nand U7890 (N_7890,N_5887,N_3909);
or U7891 (N_7891,N_1052,N_3854);
and U7892 (N_7892,N_3304,N_2310);
nor U7893 (N_7893,N_528,N_941);
nor U7894 (N_7894,N_4511,N_1142);
or U7895 (N_7895,N_4011,N_3690);
nand U7896 (N_7896,N_956,N_980);
xnor U7897 (N_7897,N_1481,N_4634);
nand U7898 (N_7898,N_439,N_5490);
and U7899 (N_7899,N_1944,N_3163);
nand U7900 (N_7900,N_2379,N_2766);
xor U7901 (N_7901,N_3228,N_5521);
and U7902 (N_7902,N_2992,N_4992);
or U7903 (N_7903,N_4550,N_3949);
or U7904 (N_7904,N_3091,N_3001);
xor U7905 (N_7905,N_208,N_745);
nor U7906 (N_7906,N_1057,N_665);
nand U7907 (N_7907,N_3443,N_2818);
nand U7908 (N_7908,N_3700,N_1643);
nor U7909 (N_7909,N_288,N_2536);
and U7910 (N_7910,N_1273,N_4286);
nor U7911 (N_7911,N_531,N_1970);
xor U7912 (N_7912,N_3740,N_3825);
nor U7913 (N_7913,N_1449,N_1956);
and U7914 (N_7914,N_1442,N_5075);
xnor U7915 (N_7915,N_3473,N_4723);
nor U7916 (N_7916,N_5685,N_2269);
nand U7917 (N_7917,N_4802,N_4799);
nand U7918 (N_7918,N_3173,N_4579);
nand U7919 (N_7919,N_1661,N_5281);
or U7920 (N_7920,N_434,N_5619);
nand U7921 (N_7921,N_5557,N_2183);
or U7922 (N_7922,N_396,N_3484);
nand U7923 (N_7923,N_2091,N_4883);
and U7924 (N_7924,N_2287,N_5542);
nand U7925 (N_7925,N_619,N_3783);
xnor U7926 (N_7926,N_1045,N_2026);
or U7927 (N_7927,N_2489,N_2440);
nand U7928 (N_7928,N_2475,N_673);
and U7929 (N_7929,N_1923,N_2092);
and U7930 (N_7930,N_3057,N_4648);
or U7931 (N_7931,N_5216,N_569);
xnor U7932 (N_7932,N_3234,N_563);
or U7933 (N_7933,N_4782,N_1462);
and U7934 (N_7934,N_3347,N_2819);
and U7935 (N_7935,N_5653,N_889);
or U7936 (N_7936,N_3006,N_2432);
nand U7937 (N_7937,N_1580,N_1015);
nand U7938 (N_7938,N_4121,N_3833);
nor U7939 (N_7939,N_2166,N_4482);
xor U7940 (N_7940,N_1569,N_2247);
nor U7941 (N_7941,N_526,N_3845);
xnor U7942 (N_7942,N_2218,N_5943);
and U7943 (N_7943,N_1022,N_5769);
or U7944 (N_7944,N_1514,N_10);
or U7945 (N_7945,N_31,N_3911);
xor U7946 (N_7946,N_5320,N_3752);
nand U7947 (N_7947,N_4068,N_2558);
xnor U7948 (N_7948,N_4703,N_4918);
or U7949 (N_7949,N_3950,N_2337);
xor U7950 (N_7950,N_2706,N_5365);
xnor U7951 (N_7951,N_870,N_3040);
xnor U7952 (N_7952,N_3457,N_470);
or U7953 (N_7953,N_1727,N_2902);
or U7954 (N_7954,N_4066,N_5870);
nand U7955 (N_7955,N_1123,N_2190);
and U7956 (N_7956,N_471,N_5765);
nand U7957 (N_7957,N_3180,N_2126);
or U7958 (N_7958,N_1214,N_4426);
nor U7959 (N_7959,N_3337,N_3441);
xnor U7960 (N_7960,N_1605,N_190);
nand U7961 (N_7961,N_5712,N_1835);
or U7962 (N_7962,N_622,N_864);
nor U7963 (N_7963,N_5354,N_2003);
nand U7964 (N_7964,N_797,N_4955);
xor U7965 (N_7965,N_2895,N_2027);
or U7966 (N_7966,N_505,N_3449);
nand U7967 (N_7967,N_4610,N_605);
or U7968 (N_7968,N_659,N_1101);
nor U7969 (N_7969,N_5751,N_3069);
and U7970 (N_7970,N_243,N_4311);
nor U7971 (N_7971,N_3157,N_2434);
xnor U7972 (N_7972,N_395,N_5658);
nor U7973 (N_7973,N_1921,N_4181);
or U7974 (N_7974,N_2583,N_5500);
or U7975 (N_7975,N_3710,N_3810);
xor U7976 (N_7976,N_3746,N_5631);
and U7977 (N_7977,N_1657,N_2235);
nand U7978 (N_7978,N_4832,N_3575);
nand U7979 (N_7979,N_1601,N_2665);
xnor U7980 (N_7980,N_3142,N_3623);
and U7981 (N_7981,N_5000,N_5195);
xnor U7982 (N_7982,N_987,N_3342);
and U7983 (N_7983,N_4387,N_3235);
nor U7984 (N_7984,N_1820,N_3128);
nor U7985 (N_7985,N_3879,N_2197);
and U7986 (N_7986,N_4350,N_4737);
or U7987 (N_7987,N_1318,N_2094);
and U7988 (N_7988,N_3649,N_3444);
nor U7989 (N_7989,N_534,N_3145);
and U7990 (N_7990,N_340,N_4772);
xnor U7991 (N_7991,N_713,N_1721);
nand U7992 (N_7992,N_1518,N_4349);
xor U7993 (N_7993,N_5362,N_3108);
nand U7994 (N_7994,N_5215,N_913);
nand U7995 (N_7995,N_3315,N_1398);
nand U7996 (N_7996,N_802,N_1726);
nand U7997 (N_7997,N_2236,N_4516);
nand U7998 (N_7998,N_1814,N_3106);
nor U7999 (N_7999,N_139,N_4450);
nor U8000 (N_8000,N_4513,N_477);
and U8001 (N_8001,N_2464,N_3148);
or U8002 (N_8002,N_3188,N_1967);
nand U8003 (N_8003,N_1330,N_3727);
and U8004 (N_8004,N_4485,N_5117);
or U8005 (N_8005,N_2466,N_3330);
nor U8006 (N_8006,N_5189,N_6);
nor U8007 (N_8007,N_2591,N_3959);
nand U8008 (N_8008,N_1544,N_3470);
and U8009 (N_8009,N_916,N_4643);
nand U8010 (N_8010,N_164,N_3246);
nor U8011 (N_8011,N_501,N_5222);
and U8012 (N_8012,N_4636,N_3513);
and U8013 (N_8013,N_2913,N_5838);
and U8014 (N_8014,N_2040,N_1575);
nand U8015 (N_8015,N_4494,N_2066);
and U8016 (N_8016,N_5018,N_1696);
xnor U8017 (N_8017,N_1692,N_4459);
or U8018 (N_8018,N_494,N_5149);
or U8019 (N_8019,N_3283,N_150);
xor U8020 (N_8020,N_4302,N_429);
nor U8021 (N_8021,N_2621,N_736);
nor U8022 (N_8022,N_421,N_1848);
xor U8023 (N_8023,N_404,N_3624);
and U8024 (N_8024,N_4159,N_5448);
or U8025 (N_8025,N_2624,N_1808);
nor U8026 (N_8026,N_3992,N_798);
or U8027 (N_8027,N_4419,N_1203);
nand U8028 (N_8028,N_2657,N_4314);
nand U8029 (N_8029,N_1595,N_2810);
xnor U8030 (N_8030,N_3278,N_5600);
or U8031 (N_8031,N_4971,N_998);
or U8032 (N_8032,N_1498,N_3966);
nor U8033 (N_8033,N_3149,N_4153);
nor U8034 (N_8034,N_1524,N_720);
nor U8035 (N_8035,N_1889,N_2639);
nor U8036 (N_8036,N_3012,N_3738);
nand U8037 (N_8037,N_3041,N_1797);
nor U8038 (N_8038,N_3357,N_2758);
or U8039 (N_8039,N_4208,N_812);
or U8040 (N_8040,N_2226,N_914);
or U8041 (N_8041,N_3781,N_63);
xnor U8042 (N_8042,N_784,N_5322);
nand U8043 (N_8043,N_3688,N_2613);
and U8044 (N_8044,N_2301,N_1685);
xor U8045 (N_8045,N_3409,N_1093);
nand U8046 (N_8046,N_1896,N_4725);
or U8047 (N_8047,N_1667,N_3723);
nor U8048 (N_8048,N_5874,N_1387);
and U8049 (N_8049,N_1724,N_865);
or U8050 (N_8050,N_3422,N_5391);
nand U8051 (N_8051,N_4188,N_179);
or U8052 (N_8052,N_5738,N_5819);
nand U8053 (N_8053,N_4788,N_1594);
xnor U8054 (N_8054,N_1528,N_2430);
nor U8055 (N_8055,N_3859,N_3297);
nor U8056 (N_8056,N_4397,N_5441);
and U8057 (N_8057,N_4031,N_1307);
nor U8058 (N_8058,N_1693,N_1826);
xnor U8059 (N_8059,N_3530,N_3482);
and U8060 (N_8060,N_5771,N_119);
xor U8061 (N_8061,N_3964,N_2445);
nand U8062 (N_8062,N_4455,N_5946);
xor U8063 (N_8063,N_4033,N_5375);
and U8064 (N_8064,N_3947,N_4532);
or U8065 (N_8065,N_2459,N_5864);
and U8066 (N_8066,N_752,N_1056);
nor U8067 (N_8067,N_2554,N_3138);
nand U8068 (N_8068,N_955,N_3368);
and U8069 (N_8069,N_669,N_813);
nand U8070 (N_8070,N_4381,N_657);
nor U8071 (N_8071,N_5829,N_688);
and U8072 (N_8072,N_593,N_2463);
or U8073 (N_8073,N_636,N_1537);
nand U8074 (N_8074,N_5880,N_3264);
nor U8075 (N_8075,N_8,N_5442);
xnor U8076 (N_8076,N_5896,N_2392);
xnor U8077 (N_8077,N_2012,N_4575);
nor U8078 (N_8078,N_1806,N_86);
and U8079 (N_8079,N_4858,N_1030);
nand U8080 (N_8080,N_3088,N_5695);
and U8081 (N_8081,N_2660,N_5367);
and U8082 (N_8082,N_4050,N_4479);
and U8083 (N_8083,N_5015,N_177);
and U8084 (N_8084,N_734,N_4389);
and U8085 (N_8085,N_2831,N_668);
xnor U8086 (N_8086,N_5433,N_2960);
and U8087 (N_8087,N_4212,N_1279);
and U8088 (N_8088,N_5293,N_5408);
or U8089 (N_8089,N_2760,N_3997);
nand U8090 (N_8090,N_2096,N_4259);
xor U8091 (N_8091,N_1769,N_4869);
nor U8092 (N_8092,N_2638,N_530);
and U8093 (N_8093,N_1452,N_4099);
and U8094 (N_8094,N_4569,N_522);
or U8095 (N_8095,N_1573,N_2816);
or U8096 (N_8096,N_1272,N_2145);
xnor U8097 (N_8097,N_3028,N_3616);
xnor U8098 (N_8098,N_3359,N_4902);
or U8099 (N_8099,N_2390,N_4523);
and U8100 (N_8100,N_3563,N_5634);
xnor U8101 (N_8101,N_1671,N_3292);
or U8102 (N_8102,N_4693,N_2884);
nor U8103 (N_8103,N_2718,N_4143);
or U8104 (N_8104,N_4912,N_3308);
nor U8105 (N_8105,N_4813,N_4559);
xnor U8106 (N_8106,N_1982,N_4514);
nand U8107 (N_8107,N_3702,N_2676);
xor U8108 (N_8108,N_4101,N_4958);
xnor U8109 (N_8109,N_2854,N_1114);
and U8110 (N_8110,N_1740,N_5417);
nor U8111 (N_8111,N_1090,N_634);
nand U8112 (N_8112,N_5088,N_1223);
and U8113 (N_8113,N_1567,N_4328);
nor U8114 (N_8114,N_4164,N_3981);
nor U8115 (N_8115,N_723,N_3742);
xnor U8116 (N_8116,N_3644,N_5035);
and U8117 (N_8117,N_5603,N_3930);
or U8118 (N_8118,N_1377,N_1062);
nand U8119 (N_8119,N_3891,N_1413);
xnor U8120 (N_8120,N_3147,N_4014);
or U8121 (N_8121,N_4445,N_5958);
nand U8122 (N_8122,N_2351,N_1782);
or U8123 (N_8123,N_1753,N_2289);
or U8124 (N_8124,N_5601,N_548);
or U8125 (N_8125,N_2716,N_486);
or U8126 (N_8126,N_989,N_3205);
nor U8127 (N_8127,N_4894,N_2522);
nand U8128 (N_8128,N_4072,N_3860);
xor U8129 (N_8129,N_1281,N_1555);
nand U8130 (N_8130,N_3164,N_2320);
nand U8131 (N_8131,N_398,N_1660);
or U8132 (N_8132,N_1958,N_5593);
nand U8133 (N_8133,N_1419,N_5594);
nor U8134 (N_8134,N_249,N_467);
and U8135 (N_8135,N_5804,N_22);
and U8136 (N_8136,N_5573,N_4388);
xnor U8137 (N_8137,N_1112,N_5976);
nor U8138 (N_8138,N_5487,N_3227);
or U8139 (N_8139,N_5931,N_5399);
nand U8140 (N_8140,N_2730,N_5345);
nor U8141 (N_8141,N_1414,N_4098);
or U8142 (N_8142,N_1673,N_2207);
or U8143 (N_8143,N_3855,N_3919);
or U8144 (N_8144,N_2576,N_877);
nand U8145 (N_8145,N_217,N_107);
and U8146 (N_8146,N_2834,N_5888);
nor U8147 (N_8147,N_2704,N_5168);
or U8148 (N_8148,N_3240,N_5817);
and U8149 (N_8149,N_2050,N_5535);
nor U8150 (N_8150,N_537,N_5697);
or U8151 (N_8151,N_2512,N_1823);
nand U8152 (N_8152,N_5249,N_5185);
nor U8153 (N_8153,N_5177,N_5431);
xnor U8154 (N_8154,N_2405,N_1356);
nand U8155 (N_8155,N_1243,N_4577);
nand U8156 (N_8156,N_4458,N_1484);
or U8157 (N_8157,N_2777,N_2165);
or U8158 (N_8158,N_1566,N_4378);
or U8159 (N_8159,N_4324,N_3445);
and U8160 (N_8160,N_5427,N_5518);
xor U8161 (N_8161,N_3171,N_4462);
nand U8162 (N_8162,N_3591,N_1792);
nand U8163 (N_8163,N_3233,N_246);
xor U8164 (N_8164,N_5546,N_776);
or U8165 (N_8165,N_1593,N_861);
or U8166 (N_8166,N_5527,N_4476);
nor U8167 (N_8167,N_1674,N_2081);
and U8168 (N_8168,N_1876,N_3030);
or U8169 (N_8169,N_81,N_3100);
and U8170 (N_8170,N_4273,N_5153);
nor U8171 (N_8171,N_5179,N_1401);
xnor U8172 (N_8172,N_3313,N_2861);
nand U8173 (N_8173,N_1224,N_3388);
nor U8174 (N_8174,N_2864,N_5846);
and U8175 (N_8175,N_1137,N_226);
nor U8176 (N_8176,N_2409,N_122);
or U8177 (N_8177,N_4403,N_2531);
nor U8178 (N_8178,N_756,N_1543);
or U8179 (N_8179,N_3801,N_2313);
xor U8180 (N_8180,N_298,N_3029);
nand U8181 (N_8181,N_2297,N_4934);
or U8182 (N_8182,N_4655,N_5873);
nor U8183 (N_8183,N_2776,N_5519);
xnor U8184 (N_8184,N_40,N_1900);
and U8185 (N_8185,N_2891,N_3160);
nand U8186 (N_8186,N_3480,N_1888);
nor U8187 (N_8187,N_5031,N_614);
nand U8188 (N_8188,N_5275,N_1707);
nor U8189 (N_8189,N_5205,N_3154);
nand U8190 (N_8190,N_2616,N_5495);
nand U8191 (N_8191,N_5134,N_1478);
nand U8192 (N_8192,N_2620,N_821);
nand U8193 (N_8193,N_4500,N_2159);
nor U8194 (N_8194,N_4862,N_782);
nand U8195 (N_8195,N_1392,N_5059);
nor U8196 (N_8196,N_2088,N_1760);
or U8197 (N_8197,N_5670,N_1633);
nand U8198 (N_8198,N_3691,N_4355);
nand U8199 (N_8199,N_5814,N_576);
nand U8200 (N_8200,N_3239,N_2285);
xor U8201 (N_8201,N_3133,N_435);
and U8202 (N_8202,N_4315,N_5073);
and U8203 (N_8203,N_5903,N_5628);
nand U8204 (N_8204,N_831,N_3198);
or U8205 (N_8205,N_1652,N_1406);
nor U8206 (N_8206,N_5509,N_4587);
and U8207 (N_8207,N_2931,N_5548);
or U8208 (N_8208,N_2184,N_917);
nand U8209 (N_8209,N_4697,N_5201);
and U8210 (N_8210,N_5621,N_474);
and U8211 (N_8211,N_143,N_5286);
or U8212 (N_8212,N_1148,N_970);
or U8213 (N_8213,N_2801,N_3137);
nor U8214 (N_8214,N_558,N_1453);
xnor U8215 (N_8215,N_4039,N_5960);
or U8216 (N_8216,N_3023,N_2195);
or U8217 (N_8217,N_4067,N_5696);
nand U8218 (N_8218,N_3402,N_2976);
or U8219 (N_8219,N_5184,N_368);
xor U8220 (N_8220,N_3744,N_118);
nand U8221 (N_8221,N_2710,N_3856);
or U8222 (N_8222,N_433,N_3689);
and U8223 (N_8223,N_3020,N_3037);
nand U8224 (N_8224,N_1959,N_5341);
nand U8225 (N_8225,N_4517,N_2246);
or U8226 (N_8226,N_2952,N_2108);
nor U8227 (N_8227,N_2143,N_3686);
xnor U8228 (N_8228,N_3027,N_5511);
nand U8229 (N_8229,N_4440,N_3305);
xnor U8230 (N_8230,N_2319,N_1621);
or U8231 (N_8231,N_5457,N_4319);
nor U8232 (N_8232,N_5867,N_2726);
nor U8233 (N_8233,N_4631,N_2979);
nor U8234 (N_8234,N_3476,N_3350);
nand U8235 (N_8235,N_294,N_1833);
nand U8236 (N_8236,N_3251,N_5760);
nor U8237 (N_8237,N_1140,N_4676);
and U8238 (N_8238,N_1054,N_402);
and U8239 (N_8239,N_907,N_103);
xnor U8240 (N_8240,N_1336,N_1190);
nand U8241 (N_8241,N_2338,N_5544);
xnor U8242 (N_8242,N_65,N_1328);
xnor U8243 (N_8243,N_1146,N_572);
and U8244 (N_8244,N_2151,N_5969);
xor U8245 (N_8245,N_2517,N_1922);
or U8246 (N_8246,N_5347,N_5673);
or U8247 (N_8247,N_2015,N_1646);
nand U8248 (N_8248,N_5643,N_5056);
and U8249 (N_8249,N_412,N_2614);
or U8250 (N_8250,N_48,N_1295);
xnor U8251 (N_8251,N_3075,N_3218);
nand U8252 (N_8252,N_1618,N_5426);
nand U8253 (N_8253,N_3927,N_5665);
xor U8254 (N_8254,N_436,N_4269);
and U8255 (N_8255,N_1205,N_814);
or U8256 (N_8256,N_2366,N_240);
nor U8257 (N_8257,N_1058,N_4363);
nor U8258 (N_8258,N_3135,N_595);
nor U8259 (N_8259,N_1592,N_4679);
or U8260 (N_8260,N_4695,N_2021);
or U8261 (N_8261,N_4341,N_1603);
or U8262 (N_8262,N_4800,N_4456);
or U8263 (N_8263,N_3540,N_3121);
and U8264 (N_8264,N_5744,N_1938);
nand U8265 (N_8265,N_1159,N_586);
xor U8266 (N_8266,N_1789,N_3423);
nor U8267 (N_8267,N_2010,N_2538);
nand U8268 (N_8268,N_1016,N_1525);
or U8269 (N_8269,N_5927,N_5802);
xnor U8270 (N_8270,N_1854,N_339);
nor U8271 (N_8271,N_5647,N_64);
nor U8272 (N_8272,N_3025,N_2838);
and U8273 (N_8273,N_626,N_5965);
nor U8274 (N_8274,N_4297,N_2450);
and U8275 (N_8275,N_158,N_5807);
xnor U8276 (N_8276,N_946,N_2978);
nor U8277 (N_8277,N_1885,N_1043);
or U8278 (N_8278,N_5576,N_3503);
nand U8279 (N_8279,N_5072,N_4768);
nand U8280 (N_8280,N_5951,N_4361);
nor U8281 (N_8281,N_287,N_4998);
nor U8282 (N_8282,N_2308,N_3893);
nor U8283 (N_8283,N_4571,N_14);
and U8284 (N_8284,N_1306,N_1228);
or U8285 (N_8285,N_2400,N_5093);
nand U8286 (N_8286,N_3606,N_5666);
nor U8287 (N_8287,N_5404,N_3876);
nand U8288 (N_8288,N_4694,N_292);
or U8289 (N_8289,N_3697,N_5291);
or U8290 (N_8290,N_1100,N_2994);
xor U8291 (N_8291,N_1390,N_1264);
nor U8292 (N_8292,N_5720,N_2480);
nor U8293 (N_8293,N_3687,N_4414);
or U8294 (N_8294,N_571,N_2125);
xor U8295 (N_8295,N_1681,N_3928);
or U8296 (N_8296,N_4256,N_5731);
nand U8297 (N_8297,N_5827,N_990);
nand U8298 (N_8298,N_4953,N_2133);
and U8299 (N_8299,N_1946,N_823);
nand U8300 (N_8300,N_4110,N_1852);
nor U8301 (N_8301,N_805,N_3668);
xnor U8302 (N_8302,N_5407,N_495);
xor U8303 (N_8303,N_314,N_2957);
nor U8304 (N_8304,N_5988,N_4206);
nand U8305 (N_8305,N_869,N_36);
nand U8306 (N_8306,N_1688,N_1834);
and U8307 (N_8307,N_3986,N_1360);
or U8308 (N_8308,N_387,N_4536);
xor U8309 (N_8309,N_44,N_2227);
nand U8310 (N_8310,N_1736,N_2887);
and U8311 (N_8311,N_3289,N_4278);
or U8312 (N_8312,N_3817,N_3526);
and U8313 (N_8313,N_2584,N_2213);
xnor U8314 (N_8314,N_4180,N_1136);
nand U8315 (N_8315,N_1948,N_5091);
xor U8316 (N_8316,N_5217,N_4073);
nand U8317 (N_8317,N_4524,N_4756);
nor U8318 (N_8318,N_1868,N_1547);
xor U8319 (N_8319,N_3732,N_2174);
xnor U8320 (N_8320,N_667,N_1538);
xor U8321 (N_8321,N_3355,N_2467);
or U8322 (N_8322,N_5617,N_449);
xor U8323 (N_8323,N_3312,N_3279);
xor U8324 (N_8324,N_4626,N_4268);
xnor U8325 (N_8325,N_2067,N_1574);
or U8326 (N_8326,N_1374,N_5918);
nor U8327 (N_8327,N_5584,N_2196);
nand U8328 (N_8328,N_565,N_3032);
or U8329 (N_8329,N_3685,N_1912);
nand U8330 (N_8330,N_3538,N_1563);
and U8331 (N_8331,N_2353,N_1064);
nor U8332 (N_8332,N_220,N_5915);
xor U8333 (N_8333,N_3766,N_923);
or U8334 (N_8334,N_674,N_3610);
nand U8335 (N_8335,N_5308,N_2152);
xor U8336 (N_8336,N_2394,N_845);
or U8337 (N_8337,N_2290,N_691);
and U8338 (N_8338,N_5865,N_4250);
nor U8339 (N_8339,N_892,N_5941);
and U8340 (N_8340,N_4795,N_1996);
xnor U8341 (N_8341,N_4468,N_279);
or U8342 (N_8342,N_5629,N_786);
nand U8343 (N_8343,N_3787,N_223);
or U8344 (N_8344,N_3940,N_4924);
nor U8345 (N_8345,N_3931,N_2141);
xor U8346 (N_8346,N_1226,N_4722);
nand U8347 (N_8347,N_1991,N_4018);
nand U8348 (N_8348,N_3397,N_3306);
or U8349 (N_8349,N_5742,N_5258);
nand U8350 (N_8350,N_481,N_5019);
xnor U8351 (N_8351,N_4954,N_4665);
and U8352 (N_8352,N_1009,N_706);
nand U8353 (N_8353,N_5878,N_4752);
or U8354 (N_8354,N_4126,N_1512);
and U8355 (N_8355,N_5269,N_2171);
and U8356 (N_8356,N_3039,N_1487);
and U8357 (N_8357,N_5324,N_1044);
nand U8358 (N_8358,N_5024,N_3972);
nor U8359 (N_8359,N_3714,N_806);
nor U8360 (N_8360,N_3242,N_4172);
xor U8361 (N_8361,N_719,N_109);
nand U8362 (N_8362,N_4163,N_2077);
nand U8363 (N_8363,N_4877,N_552);
nand U8364 (N_8364,N_749,N_1329);
nand U8365 (N_8365,N_5227,N_1757);
and U8366 (N_8366,N_2370,N_759);
nor U8367 (N_8367,N_4187,N_5094);
nand U8368 (N_8368,N_2245,N_942);
nor U8369 (N_8369,N_4848,N_815);
or U8370 (N_8370,N_3434,N_3364);
and U8371 (N_8371,N_4893,N_3633);
nor U8372 (N_8372,N_5919,N_4554);
and U8373 (N_8373,N_5166,N_5993);
and U8374 (N_8374,N_419,N_2123);
or U8375 (N_8375,N_3358,N_2921);
and U8376 (N_8376,N_151,N_3605);
nand U8377 (N_8377,N_1778,N_1945);
nor U8378 (N_8378,N_4616,N_2588);
nor U8379 (N_8379,N_3504,N_3102);
and U8380 (N_8380,N_509,N_3339);
nand U8381 (N_8381,N_2425,N_5041);
and U8382 (N_8382,N_1744,N_2775);
nand U8383 (N_8383,N_2255,N_4429);
nor U8384 (N_8384,N_5972,N_3150);
xor U8385 (N_8385,N_2741,N_1666);
and U8386 (N_8386,N_2147,N_2566);
nand U8387 (N_8387,N_4300,N_4148);
xnor U8388 (N_8388,N_184,N_2057);
nand U8389 (N_8389,N_4730,N_1425);
nand U8390 (N_8390,N_847,N_3477);
and U8391 (N_8391,N_1590,N_4086);
or U8392 (N_8392,N_3577,N_3802);
nor U8393 (N_8393,N_922,N_1454);
xor U8394 (N_8394,N_5030,N_5109);
nand U8395 (N_8395,N_3951,N_3286);
nand U8396 (N_8396,N_1138,N_4317);
or U8397 (N_8397,N_5226,N_5830);
and U8398 (N_8398,N_5750,N_4855);
and U8399 (N_8399,N_3197,N_2587);
or U8400 (N_8400,N_804,N_4843);
nor U8401 (N_8401,N_1012,N_3322);
nor U8402 (N_8402,N_2389,N_463);
and U8403 (N_8403,N_3721,N_320);
or U8404 (N_8404,N_1156,N_300);
or U8405 (N_8405,N_5596,N_2501);
nor U8406 (N_8406,N_4062,N_2932);
and U8407 (N_8407,N_3256,N_2520);
and U8408 (N_8408,N_5517,N_3792);
nor U8409 (N_8409,N_2481,N_967);
xnor U8410 (N_8410,N_4310,N_5459);
xor U8411 (N_8411,N_472,N_4688);
xor U8412 (N_8412,N_2359,N_3589);
nand U8413 (N_8413,N_584,N_5305);
xor U8414 (N_8414,N_5840,N_3086);
nor U8415 (N_8415,N_5877,N_77);
and U8416 (N_8416,N_301,N_464);
xnor U8417 (N_8417,N_2914,N_5372);
and U8418 (N_8418,N_1903,N_2185);
xor U8419 (N_8419,N_280,N_3225);
or U8420 (N_8420,N_4096,N_2804);
nand U8421 (N_8421,N_581,N_5748);
xor U8422 (N_8422,N_5425,N_1391);
xnor U8423 (N_8423,N_377,N_4210);
xnor U8424 (N_8424,N_4127,N_1292);
and U8425 (N_8425,N_5907,N_5008);
and U8426 (N_8426,N_5759,N_2782);
and U8427 (N_8427,N_1236,N_5791);
nand U8428 (N_8428,N_4584,N_3224);
nand U8429 (N_8429,N_5412,N_3363);
or U8430 (N_8430,N_1359,N_1730);
nand U8431 (N_8431,N_21,N_771);
nor U8432 (N_8432,N_5604,N_4982);
xnor U8433 (N_8433,N_4308,N_644);
nor U8434 (N_8434,N_5424,N_1816);
or U8435 (N_8435,N_968,N_5524);
xnor U8436 (N_8436,N_3333,N_3765);
or U8437 (N_8437,N_5703,N_5028);
nor U8438 (N_8438,N_3340,N_1800);
nor U8439 (N_8439,N_3873,N_5180);
and U8440 (N_8440,N_250,N_1913);
xnor U8441 (N_8441,N_3265,N_4030);
xor U8442 (N_8442,N_4421,N_5810);
xor U8443 (N_8443,N_4599,N_5485);
and U8444 (N_8444,N_2835,N_3288);
nor U8445 (N_8445,N_5818,N_4000);
and U8446 (N_8446,N_346,N_286);
nor U8447 (N_8447,N_4372,N_3214);
nand U8448 (N_8448,N_3574,N_4095);
and U8449 (N_8449,N_146,N_3436);
and U8450 (N_8450,N_455,N_2561);
or U8451 (N_8451,N_4565,N_5147);
nand U8452 (N_8452,N_4678,N_2526);
nand U8453 (N_8453,N_3524,N_3022);
and U8454 (N_8454,N_3656,N_2449);
or U8455 (N_8455,N_3780,N_29);
xnor U8456 (N_8456,N_5900,N_5040);
nor U8457 (N_8457,N_795,N_4407);
xnor U8458 (N_8458,N_5016,N_2663);
xnor U8459 (N_8459,N_5097,N_5554);
nor U8460 (N_8460,N_1396,N_722);
nor U8461 (N_8461,N_1560,N_3593);
and U8462 (N_8462,N_2959,N_1411);
xor U8463 (N_8463,N_5655,N_5990);
nor U8464 (N_8464,N_3056,N_1167);
or U8465 (N_8465,N_1169,N_2129);
and U8466 (N_8466,N_4081,N_4439);
nand U8467 (N_8467,N_2764,N_1131);
xnor U8468 (N_8468,N_4509,N_123);
and U8469 (N_8469,N_1267,N_3794);
and U8470 (N_8470,N_4653,N_3672);
or U8471 (N_8471,N_4157,N_1634);
xor U8472 (N_8472,N_3519,N_1026);
and U8473 (N_8473,N_1870,N_4359);
nand U8474 (N_8474,N_4837,N_1096);
nand U8475 (N_8475,N_3013,N_4231);
and U8476 (N_8476,N_3116,N_5369);
nor U8477 (N_8477,N_1756,N_332);
nand U8478 (N_8478,N_1672,N_2643);
nand U8479 (N_8479,N_5651,N_4545);
nor U8480 (N_8480,N_3602,N_5985);
nand U8481 (N_8481,N_5688,N_4416);
nor U8482 (N_8482,N_4666,N_2292);
nor U8483 (N_8483,N_2487,N_3290);
xnor U8484 (N_8484,N_3262,N_4605);
xnor U8485 (N_8485,N_3334,N_3824);
nor U8486 (N_8486,N_4422,N_1803);
and U8487 (N_8487,N_5355,N_5599);
and U8488 (N_8488,N_1954,N_3421);
and U8489 (N_8489,N_3005,N_3638);
nor U8490 (N_8490,N_4109,N_2869);
and U8491 (N_8491,N_1907,N_3852);
nand U8492 (N_8492,N_4846,N_145);
xor U8493 (N_8493,N_1636,N_5444);
and U8494 (N_8494,N_3323,N_872);
nand U8495 (N_8495,N_737,N_4663);
xor U8496 (N_8496,N_4546,N_2476);
nor U8497 (N_8497,N_94,N_3914);
xnor U8498 (N_8498,N_1283,N_129);
and U8499 (N_8499,N_1972,N_2930);
xnor U8500 (N_8500,N_5551,N_2017);
xor U8501 (N_8501,N_2803,N_5732);
nand U8502 (N_8502,N_992,N_3203);
nand U8503 (N_8503,N_611,N_1989);
nor U8504 (N_8504,N_2610,N_4623);
or U8505 (N_8505,N_4686,N_5858);
nor U8506 (N_8506,N_5297,N_1204);
nor U8507 (N_8507,N_1831,N_2761);
or U8508 (N_8508,N_2515,N_519);
nand U8509 (N_8509,N_2333,N_4051);
or U8510 (N_8510,N_2598,N_1091);
xor U8511 (N_8511,N_5103,N_2562);
nand U8512 (N_8512,N_4395,N_1540);
xor U8513 (N_8513,N_2028,N_5936);
nor U8514 (N_8514,N_2148,N_4907);
or U8515 (N_8515,N_3045,N_5623);
or U8516 (N_8516,N_306,N_663);
xnor U8517 (N_8517,N_3894,N_3078);
xnor U8518 (N_8518,N_5566,N_4897);
nand U8519 (N_8519,N_327,N_5278);
nor U8520 (N_8520,N_3954,N_863);
nand U8521 (N_8521,N_507,N_1446);
and U8522 (N_8522,N_3904,N_5182);
or U8523 (N_8523,N_392,N_5090);
and U8524 (N_8524,N_3497,N_52);
nor U8525 (N_8525,N_985,N_5689);
and U8526 (N_8526,N_4461,N_3857);
and U8527 (N_8527,N_1841,N_2271);
xnor U8528 (N_8528,N_4895,N_3725);
xor U8529 (N_8529,N_2922,N_4637);
nor U8530 (N_8530,N_3988,N_4241);
nand U8531 (N_8531,N_2044,N_1617);
and U8532 (N_8532,N_2505,N_1827);
nand U8533 (N_8533,N_1466,N_2427);
and U8534 (N_8534,N_4370,N_4452);
and U8535 (N_8535,N_487,N_3111);
and U8536 (N_8536,N_5232,N_4601);
or U8537 (N_8537,N_3998,N_770);
nor U8538 (N_8538,N_5240,N_4224);
xor U8539 (N_8539,N_330,N_3768);
nor U8540 (N_8540,N_3958,N_2722);
and U8541 (N_8541,N_70,N_1941);
nor U8542 (N_8542,N_731,N_3832);
nor U8543 (N_8543,N_533,N_141);
nor U8544 (N_8544,N_1399,N_2964);
or U8545 (N_8545,N_4755,N_5165);
nor U8546 (N_8546,N_1557,N_401);
nand U8547 (N_8547,N_1488,N_5687);
xnor U8548 (N_8548,N_1422,N_678);
nand U8549 (N_8549,N_4941,N_5026);
nor U8550 (N_8550,N_4553,N_2679);
nand U8551 (N_8551,N_4972,N_4267);
and U8552 (N_8552,N_670,N_4054);
or U8553 (N_8553,N_1077,N_4492);
and U8554 (N_8554,N_4020,N_1599);
xor U8555 (N_8555,N_4925,N_3695);
or U8556 (N_8556,N_4748,N_4712);
or U8557 (N_8557,N_4944,N_5386);
nor U8558 (N_8558,N_2065,N_514);
or U8559 (N_8559,N_835,N_4590);
nor U8560 (N_8560,N_2488,N_5700);
nor U8561 (N_8561,N_5356,N_46);
nor U8562 (N_8562,N_2748,N_3110);
or U8563 (N_8563,N_816,N_2325);
nor U8564 (N_8564,N_2332,N_4595);
nand U8565 (N_8565,N_2720,N_149);
and U8566 (N_8566,N_2828,N_2956);
nand U8567 (N_8567,N_263,N_2387);
and U8568 (N_8568,N_3207,N_2210);
or U8569 (N_8569,N_2618,N_2567);
nor U8570 (N_8570,N_451,N_3901);
xor U8571 (N_8571,N_4673,N_2812);
or U8572 (N_8572,N_4717,N_2575);
and U8573 (N_8573,N_3050,N_4803);
nand U8574 (N_8574,N_5784,N_2924);
or U8575 (N_8575,N_4775,N_479);
and U8576 (N_8576,N_3329,N_5515);
nand U8577 (N_8577,N_2765,N_4146);
or U8578 (N_8578,N_239,N_96);
nor U8579 (N_8579,N_2824,N_2398);
nand U8580 (N_8580,N_1748,N_5188);
and U8581 (N_8581,N_5835,N_5944);
or U8582 (N_8582,N_2963,N_2169);
nor U8583 (N_8583,N_5501,N_5861);
and U8584 (N_8584,N_5343,N_3367);
or U8585 (N_8585,N_1176,N_5562);
nor U8586 (N_8586,N_2485,N_2316);
or U8587 (N_8587,N_5384,N_261);
nand U8588 (N_8588,N_963,N_3967);
or U8589 (N_8589,N_1423,N_4920);
xor U8590 (N_8590,N_0,N_2291);
or U8591 (N_8591,N_2984,N_4358);
or U8592 (N_8592,N_2162,N_5100);
xnor U8593 (N_8593,N_1624,N_3596);
nand U8594 (N_8594,N_4821,N_960);
nand U8595 (N_8595,N_4765,N_285);
nor U8596 (N_8596,N_5745,N_5420);
nor U8597 (N_8597,N_1507,N_5538);
or U8598 (N_8598,N_3155,N_1504);
or U8599 (N_8599,N_5110,N_3494);
or U8600 (N_8600,N_5003,N_2382);
or U8601 (N_8601,N_5789,N_4990);
xor U8602 (N_8602,N_5083,N_3724);
nand U8603 (N_8603,N_5693,N_2868);
xor U8604 (N_8604,N_1552,N_3430);
nand U8605 (N_8605,N_5691,N_1302);
xor U8606 (N_8606,N_3219,N_174);
or U8607 (N_8607,N_1589,N_873);
and U8608 (N_8608,N_5113,N_5084);
nor U8609 (N_8609,N_2949,N_983);
or U8610 (N_8610,N_4606,N_3365);
xor U8611 (N_8611,N_2157,N_1333);
or U8612 (N_8612,N_5183,N_5265);
nor U8613 (N_8613,N_3373,N_3054);
and U8614 (N_8614,N_3786,N_57);
nor U8615 (N_8615,N_788,N_3636);
nor U8616 (N_8616,N_3201,N_621);
and U8617 (N_8617,N_707,N_933);
nand U8618 (N_8618,N_5798,N_1928);
or U8619 (N_8619,N_5144,N_4374);
and U8620 (N_8620,N_4961,N_588);
and U8621 (N_8621,N_827,N_1968);
or U8622 (N_8622,N_3756,N_2082);
nor U8623 (N_8623,N_2356,N_2296);
nand U8624 (N_8624,N_5737,N_4849);
or U8625 (N_8625,N_5139,N_1637);
or U8626 (N_8626,N_2937,N_1300);
or U8627 (N_8627,N_2193,N_1840);
nor U8628 (N_8628,N_2773,N_5390);
xor U8629 (N_8629,N_4560,N_2156);
nor U8630 (N_8630,N_1522,N_1978);
nor U8631 (N_8631,N_2153,N_321);
or U8632 (N_8632,N_5239,N_259);
nor U8633 (N_8633,N_325,N_5471);
or U8634 (N_8634,N_2118,N_3875);
xnor U8635 (N_8635,N_2649,N_456);
xnor U8636 (N_8636,N_714,N_5032);
nor U8637 (N_8637,N_161,N_5379);
and U8638 (N_8638,N_5474,N_3151);
nor U8639 (N_8639,N_4541,N_5530);
or U8640 (N_8640,N_1517,N_3991);
nand U8641 (N_8641,N_1040,N_3177);
and U8642 (N_8642,N_2498,N_5579);
or U8643 (N_8643,N_1950,N_5260);
nor U8644 (N_8644,N_4733,N_1705);
or U8645 (N_8645,N_1404,N_3630);
nor U8646 (N_8646,N_4680,N_5836);
nand U8647 (N_8647,N_427,N_2058);
nor U8648 (N_8648,N_2348,N_3583);
nor U8649 (N_8649,N_2903,N_2024);
or U8650 (N_8650,N_4742,N_500);
xnor U8651 (N_8651,N_5077,N_602);
xnor U8652 (N_8652,N_2746,N_5672);
and U8653 (N_8653,N_2918,N_717);
or U8654 (N_8654,N_1839,N_4977);
or U8655 (N_8655,N_1071,N_5555);
xnor U8656 (N_8656,N_1135,N_2669);
or U8657 (N_8657,N_5334,N_2051);
nor U8658 (N_8658,N_4791,N_5684);
nor U8659 (N_8659,N_5262,N_5882);
xor U8660 (N_8660,N_3561,N_4078);
and U8661 (N_8661,N_754,N_1965);
xnor U8662 (N_8662,N_4189,N_2286);
or U8663 (N_8663,N_4475,N_4646);
xnor U8664 (N_8664,N_5136,N_5429);
xnor U8665 (N_8665,N_5238,N_5332);
and U8666 (N_8666,N_1842,N_2061);
or U8667 (N_8667,N_751,N_570);
or U8668 (N_8668,N_2074,N_2191);
or U8669 (N_8669,N_4351,N_1253);
nand U8670 (N_8670,N_4061,N_3258);
xnor U8671 (N_8671,N_5708,N_5301);
and U8672 (N_8672,N_2284,N_4168);
and U8673 (N_8673,N_3343,N_3316);
xnor U8674 (N_8674,N_4602,N_2355);
or U8675 (N_8675,N_5857,N_5491);
nand U8676 (N_8676,N_772,N_4945);
xnor U8677 (N_8677,N_2915,N_121);
xor U8678 (N_8678,N_5682,N_826);
or U8679 (N_8679,N_2447,N_3098);
xor U8680 (N_8680,N_1998,N_732);
and U8681 (N_8681,N_234,N_1150);
nand U8682 (N_8682,N_2897,N_2693);
nand U8683 (N_8683,N_3216,N_662);
and U8684 (N_8684,N_4271,N_2037);
nand U8685 (N_8685,N_3849,N_896);
xnor U8686 (N_8686,N_3535,N_1708);
and U8687 (N_8687,N_2128,N_4870);
and U8688 (N_8688,N_789,N_7);
nand U8689 (N_8689,N_2443,N_5916);
xor U8690 (N_8690,N_3720,N_4527);
nor U8691 (N_8691,N_1678,N_2441);
xnor U8692 (N_8692,N_3062,N_1111);
xnor U8693 (N_8693,N_4729,N_5952);
nand U8694 (N_8694,N_3872,N_3666);
xnor U8695 (N_8695,N_3803,N_2415);
xnor U8696 (N_8696,N_1510,N_2170);
nand U8697 (N_8697,N_5892,N_2072);
or U8698 (N_8698,N_4824,N_1516);
nor U8699 (N_8699,N_2787,N_3105);
nor U8700 (N_8700,N_2878,N_1099);
nand U8701 (N_8701,N_2508,N_5006);
nand U8702 (N_8702,N_1358,N_1741);
or U8703 (N_8703,N_430,N_2799);
nand U8704 (N_8704,N_2486,N_1804);
nor U8705 (N_8705,N_709,N_1327);
nor U8706 (N_8706,N_1161,N_4839);
and U8707 (N_8707,N_4946,N_1155);
and U8708 (N_8708,N_3274,N_1980);
and U8709 (N_8709,N_2697,N_4567);
nand U8710 (N_8710,N_2852,N_757);
xnor U8711 (N_8711,N_4219,N_3427);
nand U8712 (N_8712,N_5644,N_4892);
nand U8713 (N_8713,N_5580,N_952);
nand U8714 (N_8714,N_4751,N_1349);
nor U8715 (N_8715,N_2282,N_2537);
nor U8716 (N_8716,N_5138,N_3646);
nand U8717 (N_8717,N_5811,N_3743);
nand U8718 (N_8718,N_3371,N_201);
and U8719 (N_8719,N_4649,N_1229);
xor U8720 (N_8720,N_4049,N_2230);
and U8721 (N_8721,N_2778,N_2137);
or U8722 (N_8722,N_2745,N_1915);
nor U8723 (N_8723,N_5734,N_2751);
or U8724 (N_8724,N_5313,N_1843);
xnor U8725 (N_8725,N_1355,N_3741);
nor U8726 (N_8726,N_1588,N_3186);
nand U8727 (N_8727,N_2680,N_3692);
or U8728 (N_8728,N_5605,N_2281);
or U8729 (N_8729,N_1331,N_5986);
nand U8730 (N_8730,N_1083,N_15);
xnor U8731 (N_8731,N_2482,N_2630);
xnor U8732 (N_8732,N_1221,N_5228);
nand U8733 (N_8733,N_2220,N_2163);
xnor U8734 (N_8734,N_414,N_1539);
xnor U8735 (N_8735,N_3826,N_2121);
nand U8736 (N_8736,N_3560,N_1866);
nand U8737 (N_8737,N_1351,N_3170);
or U8738 (N_8738,N_2448,N_5756);
nand U8739 (N_8739,N_3455,N_424);
nor U8740 (N_8740,N_5121,N_2402);
and U8741 (N_8741,N_3392,N_3407);
and U8742 (N_8742,N_973,N_4251);
and U8743 (N_8743,N_986,N_1326);
nand U8744 (N_8744,N_2809,N_3684);
nor U8745 (N_8745,N_1037,N_2461);
nor U8746 (N_8746,N_2546,N_3769);
nand U8747 (N_8747,N_1710,N_1319);
nand U8748 (N_8748,N_3811,N_1242);
nor U8749 (N_8749,N_4084,N_82);
and U8750 (N_8750,N_1851,N_3474);
nor U8751 (N_8751,N_4544,N_3299);
nor U8752 (N_8752,N_4037,N_3733);
nor U8753 (N_8753,N_3247,N_3989);
xor U8754 (N_8754,N_4393,N_3296);
nand U8755 (N_8755,N_4182,N_1495);
nand U8756 (N_8756,N_3601,N_441);
nand U8757 (N_8757,N_1447,N_2678);
nor U8758 (N_8758,N_2016,N_3996);
xnor U8759 (N_8759,N_5377,N_5196);
nand U8760 (N_8760,N_5363,N_681);
xor U8761 (N_8761,N_1830,N_1519);
nand U8762 (N_8762,N_959,N_3440);
nand U8763 (N_8763,N_1385,N_1754);
or U8764 (N_8764,N_2944,N_2295);
nor U8765 (N_8765,N_4375,N_680);
or U8766 (N_8766,N_4525,N_1746);
or U8767 (N_8767,N_2201,N_1535);
or U8768 (N_8768,N_962,N_1584);
xnor U8769 (N_8769,N_5021,N_1784);
nand U8770 (N_8770,N_3587,N_3629);
nor U8771 (N_8771,N_5206,N_5259);
or U8772 (N_8772,N_4827,N_5119);
nor U8773 (N_8773,N_1559,N_3452);
or U8774 (N_8774,N_5683,N_1686);
nor U8775 (N_8775,N_5130,N_5921);
and U8776 (N_8776,N_5440,N_1742);
xor U8777 (N_8777,N_3634,N_348);
nor U8778 (N_8778,N_777,N_3074);
nand U8779 (N_8779,N_4390,N_1172);
nand U8780 (N_8780,N_4760,N_2364);
nand U8781 (N_8781,N_4093,N_5821);
nand U8782 (N_8782,N_4778,N_5795);
xor U8783 (N_8783,N_2412,N_4783);
xor U8784 (N_8784,N_3183,N_1);
xnor U8785 (N_8785,N_498,N_5662);
or U8786 (N_8786,N_1163,N_319);
or U8787 (N_8787,N_4710,N_2842);
nand U8788 (N_8788,N_1284,N_3122);
nand U8789 (N_8789,N_1607,N_338);
xnor U8790 (N_8790,N_4786,N_2421);
or U8791 (N_8791,N_5256,N_3092);
xnor U8792 (N_8792,N_3118,N_4682);
or U8793 (N_8793,N_3425,N_2547);
nand U8794 (N_8794,N_4218,N_1227);
nand U8795 (N_8795,N_3383,N_549);
and U8796 (N_8796,N_5430,N_2514);
nor U8797 (N_8797,N_1010,N_2381);
nor U8798 (N_8798,N_1263,N_748);
nor U8799 (N_8799,N_3018,N_4198);
xnor U8800 (N_8800,N_5841,N_875);
nor U8801 (N_8801,N_2406,N_3840);
and U8802 (N_8802,N_2989,N_592);
and U8803 (N_8803,N_3341,N_1246);
nor U8804 (N_8804,N_3099,N_3325);
nor U8805 (N_8805,N_3671,N_2250);
nand U8806 (N_8806,N_5245,N_278);
xor U8807 (N_8807,N_3608,N_4716);
and U8808 (N_8808,N_4580,N_2363);
or U8809 (N_8809,N_2144,N_3495);
or U8810 (N_8810,N_482,N_3458);
and U8811 (N_8811,N_5078,N_2996);
nor U8812 (N_8812,N_4661,N_34);
nor U8813 (N_8813,N_1957,N_4193);
nor U8814 (N_8814,N_165,N_5209);
and U8815 (N_8815,N_1847,N_210);
nand U8816 (N_8816,N_1303,N_4963);
nor U8817 (N_8817,N_5353,N_5174);
and U8818 (N_8818,N_5578,N_2542);
nor U8819 (N_8819,N_1616,N_5368);
nand U8820 (N_8820,N_3726,N_920);
xor U8821 (N_8821,N_5876,N_3647);
and U8822 (N_8822,N_364,N_743);
xor U8823 (N_8823,N_1901,N_5033);
xnor U8824 (N_8824,N_270,N_4353);
and U8825 (N_8825,N_5122,N_4650);
xnor U8826 (N_8826,N_1219,N_1184);
xnor U8827 (N_8827,N_1714,N_2783);
xnor U8828 (N_8828,N_2154,N_4863);
xor U8829 (N_8829,N_1485,N_1774);
and U8830 (N_8830,N_461,N_112);
or U8831 (N_8831,N_203,N_2375);
nor U8832 (N_8832,N_523,N_2033);
nand U8833 (N_8833,N_2396,N_3681);
or U8834 (N_8834,N_5711,N_5799);
or U8835 (N_8835,N_3774,N_3607);
nor U8836 (N_8836,N_1824,N_1962);
xor U8837 (N_8837,N_5428,N_3332);
or U8838 (N_8838,N_3842,N_3129);
xor U8839 (N_8839,N_4331,N_4129);
or U8840 (N_8840,N_2194,N_3782);
xor U8841 (N_8841,N_5346,N_5674);
and U8842 (N_8842,N_45,N_746);
or U8843 (N_8843,N_194,N_2206);
and U8844 (N_8844,N_1747,N_305);
xnor U8845 (N_8845,N_4013,N_3795);
nor U8846 (N_8846,N_3008,N_2938);
xor U8847 (N_8847,N_3828,N_3411);
or U8848 (N_8848,N_1501,N_4904);
and U8849 (N_8849,N_2892,N_2655);
xnor U8850 (N_8850,N_938,N_4607);
and U8851 (N_8851,N_3641,N_3734);
nand U8852 (N_8852,N_547,N_948);
nor U8853 (N_8853,N_444,N_4662);
xor U8854 (N_8854,N_5270,N_283);
nand U8855 (N_8855,N_5894,N_675);
nor U8856 (N_8856,N_504,N_5423);
nand U8857 (N_8857,N_5340,N_1051);
or U8858 (N_8858,N_654,N_3162);
or U8859 (N_8859,N_3437,N_3902);
nor U8860 (N_8860,N_212,N_5661);
and U8861 (N_8861,N_224,N_2413);
nand U8862 (N_8862,N_4469,N_1703);
and U8863 (N_8863,N_3916,N_3617);
and U8864 (N_8864,N_2186,N_2533);
nand U8865 (N_8865,N_780,N_382);
nor U8866 (N_8866,N_1995,N_4226);
xor U8867 (N_8867,N_3511,N_4162);
and U8868 (N_8868,N_5793,N_3760);
nand U8869 (N_8869,N_5752,N_2216);
nor U8870 (N_8870,N_5832,N_4156);
nand U8871 (N_8871,N_2424,N_5589);
nor U8872 (N_8872,N_4603,N_1583);
nand U8873 (N_8873,N_4628,N_266);
or U8874 (N_8874,N_5010,N_3464);
nor U8875 (N_8875,N_1932,N_2055);
nand U8876 (N_8876,N_1235,N_911);
and U8877 (N_8877,N_4323,N_1087);
nand U8878 (N_8878,N_1431,N_3613);
nand U8879 (N_8879,N_2985,N_437);
and U8880 (N_8880,N_3369,N_1445);
or U8881 (N_8881,N_277,N_5868);
xor U8882 (N_8882,N_4177,N_2410);
and U8883 (N_8883,N_792,N_2249);
xor U8884 (N_8884,N_2496,N_4563);
or U8885 (N_8885,N_3529,N_3489);
nand U8886 (N_8886,N_728,N_4057);
nor U8887 (N_8887,N_3270,N_3486);
and U8888 (N_8888,N_3522,N_342);
nor U8889 (N_8889,N_4009,N_715);
and U8890 (N_8890,N_2534,N_5449);
or U8891 (N_8891,N_3711,N_1768);
or U8892 (N_8892,N_1984,N_1947);
xor U8893 (N_8893,N_4171,N_462);
nand U8894 (N_8894,N_4704,N_4864);
and U8895 (N_8895,N_4282,N_4510);
nand U8896 (N_8896,N_3398,N_1582);
nand U8897 (N_8897,N_2756,N_5187);
nand U8898 (N_8898,N_5234,N_4244);
nor U8899 (N_8899,N_2052,N_4017);
nand U8900 (N_8900,N_642,N_4919);
nor U8901 (N_8901,N_829,N_162);
nor U8902 (N_8902,N_3127,N_2272);
or U8903 (N_8903,N_5317,N_265);
xor U8904 (N_8904,N_256,N_3134);
and U8905 (N_8905,N_1554,N_5133);
or U8906 (N_8906,N_2233,N_4473);
or U8907 (N_8907,N_5023,N_4979);
nor U8908 (N_8908,N_5046,N_1631);
nand U8909 (N_8909,N_2085,N_207);
or U8910 (N_8910,N_2946,N_4276);
or U8911 (N_8911,N_3211,N_5582);
nor U8912 (N_8912,N_4447,N_540);
or U8913 (N_8913,N_3068,N_74);
or U8914 (N_8914,N_5488,N_233);
and U8915 (N_8915,N_4630,N_4023);
nand U8916 (N_8916,N_4564,N_83);
nor U8917 (N_8917,N_5272,N_4771);
or U8918 (N_8918,N_5761,N_3979);
xor U8919 (N_8919,N_3635,N_2401);
or U8920 (N_8920,N_3694,N_5851);
and U8921 (N_8921,N_5954,N_3399);
and U8922 (N_8922,N_3136,N_686);
or U8923 (N_8923,N_4335,N_1627);
and U8924 (N_8924,N_2724,N_824);
nor U8925 (N_8925,N_5843,N_1181);
xnor U8926 (N_8926,N_2181,N_3984);
and U8927 (N_8927,N_260,N_4417);
and U8928 (N_8928,N_394,N_4576);
and U8929 (N_8929,N_2189,N_5013);
xnor U8930 (N_8930,N_363,N_3896);
nor U8931 (N_8931,N_5146,N_5318);
nand U8932 (N_8932,N_1213,N_508);
or U8933 (N_8933,N_837,N_5823);
and U8934 (N_8934,N_4207,N_5778);
xor U8935 (N_8935,N_2317,N_5797);
nand U8936 (N_8936,N_5181,N_4263);
or U8937 (N_8937,N_4090,N_5203);
xnor U8938 (N_8938,N_5736,N_1352);
xor U8939 (N_8939,N_5366,N_5158);
xnor U8940 (N_8940,N_2457,N_3415);
xor U8941 (N_8941,N_4097,N_890);
xnor U8942 (N_8942,N_5325,N_2999);
and U8943 (N_8943,N_236,N_475);
xor U8944 (N_8944,N_3467,N_981);
xor U8945 (N_8945,N_3119,N_5438);
xor U8946 (N_8946,N_5403,N_1133);
nand U8947 (N_8947,N_1737,N_3143);
xor U8948 (N_8948,N_4875,N_1994);
xor U8949 (N_8949,N_2800,N_4774);
xor U8950 (N_8950,N_4201,N_2601);
nand U8951 (N_8951,N_4008,N_5808);
nand U8952 (N_8952,N_1403,N_4750);
and U8953 (N_8953,N_4160,N_587);
nand U8954 (N_8954,N_1007,N_2469);
or U8955 (N_8955,N_3664,N_87);
or U8956 (N_8956,N_2814,N_5833);
nor U8957 (N_8957,N_4326,N_1314);
or U8958 (N_8958,N_1882,N_925);
nor U8959 (N_8959,N_3886,N_2980);
or U8960 (N_8960,N_2843,N_3659);
nor U8961 (N_8961,N_1973,N_218);
xnor U8962 (N_8962,N_2617,N_5479);
nor U8963 (N_8963,N_3378,N_3158);
or U8964 (N_8964,N_3453,N_874);
and U8965 (N_8965,N_386,N_3064);
nand U8966 (N_8966,N_4012,N_3564);
xor U8967 (N_8967,N_3331,N_3345);
nand U8968 (N_8968,N_5531,N_60);
nand U8969 (N_8969,N_5905,N_1018);
or U8970 (N_8970,N_2474,N_2483);
and U8971 (N_8971,N_4533,N_3166);
and U8972 (N_8972,N_1209,N_1373);
and U8973 (N_8973,N_651,N_3374);
and U8974 (N_8974,N_842,N_4103);
and U8975 (N_8975,N_2728,N_1459);
xnor U8976 (N_8976,N_1287,N_2662);
xor U8977 (N_8977,N_5453,N_4976);
and U8978 (N_8978,N_2951,N_1202);
nor U8979 (N_8979,N_4368,N_574);
nand U8980 (N_8980,N_3109,N_5933);
or U8981 (N_8981,N_1680,N_2846);
or U8982 (N_8982,N_5890,N_156);
nor U8983 (N_8983,N_1856,N_2278);
and U8984 (N_8984,N_4552,N_4005);
or U8985 (N_8985,N_1615,N_5);
nor U8986 (N_8986,N_3962,N_5065);
nor U8987 (N_8987,N_3038,N_2025);
nand U8988 (N_8988,N_888,N_596);
nor U8989 (N_8989,N_4660,N_214);
nand U8990 (N_8990,N_4790,N_5924);
or U8991 (N_8991,N_5455,N_1790);
nand U8992 (N_8992,N_2455,N_466);
and U8993 (N_8993,N_4493,N_3243);
nor U8994 (N_8994,N_206,N_554);
or U8995 (N_8995,N_2429,N_3908);
and U8996 (N_8996,N_5418,N_4203);
nor U8997 (N_8997,N_3082,N_5587);
xor U8998 (N_8998,N_4927,N_1931);
xor U8999 (N_8999,N_3063,N_5975);
and U9000 (N_9000,N_817,N_1815);
xnor U9001 (N_9001,N_5085,N_4131);
or U9002 (N_9002,N_337,N_5312);
nor U9003 (N_9003,N_245,N_5648);
nand U9004 (N_9004,N_2470,N_3341);
or U9005 (N_9005,N_3517,N_1464);
or U9006 (N_9006,N_4139,N_2804);
or U9007 (N_9007,N_3258,N_3098);
or U9008 (N_9008,N_4591,N_3399);
or U9009 (N_9009,N_1497,N_3011);
nand U9010 (N_9010,N_3264,N_3638);
nor U9011 (N_9011,N_1441,N_4988);
nand U9012 (N_9012,N_5129,N_300);
nor U9013 (N_9013,N_3884,N_4384);
and U9014 (N_9014,N_1493,N_4995);
or U9015 (N_9015,N_609,N_3148);
or U9016 (N_9016,N_4878,N_1942);
nand U9017 (N_9017,N_4148,N_1551);
and U9018 (N_9018,N_2767,N_5040);
nand U9019 (N_9019,N_4375,N_2076);
or U9020 (N_9020,N_4739,N_1845);
xnor U9021 (N_9021,N_840,N_4486);
nor U9022 (N_9022,N_1879,N_3771);
nand U9023 (N_9023,N_5841,N_4375);
nand U9024 (N_9024,N_1686,N_2069);
nand U9025 (N_9025,N_4586,N_4426);
and U9026 (N_9026,N_864,N_5713);
nand U9027 (N_9027,N_1484,N_578);
nand U9028 (N_9028,N_2717,N_5775);
nand U9029 (N_9029,N_5438,N_2278);
and U9030 (N_9030,N_5348,N_4114);
or U9031 (N_9031,N_5379,N_3178);
xnor U9032 (N_9032,N_5768,N_3143);
or U9033 (N_9033,N_4903,N_5176);
and U9034 (N_9034,N_2079,N_1839);
nor U9035 (N_9035,N_301,N_3918);
nor U9036 (N_9036,N_1411,N_4096);
nand U9037 (N_9037,N_2756,N_3000);
xnor U9038 (N_9038,N_3010,N_1042);
and U9039 (N_9039,N_3221,N_1440);
nand U9040 (N_9040,N_1658,N_3922);
nand U9041 (N_9041,N_4223,N_174);
or U9042 (N_9042,N_461,N_3952);
or U9043 (N_9043,N_4265,N_836);
nor U9044 (N_9044,N_4518,N_1995);
nor U9045 (N_9045,N_233,N_1128);
nor U9046 (N_9046,N_3054,N_2258);
xor U9047 (N_9047,N_1510,N_984);
or U9048 (N_9048,N_1553,N_1508);
xor U9049 (N_9049,N_4198,N_1943);
nand U9050 (N_9050,N_3572,N_3399);
and U9051 (N_9051,N_4297,N_1266);
and U9052 (N_9052,N_171,N_5254);
and U9053 (N_9053,N_1683,N_3487);
xor U9054 (N_9054,N_73,N_4986);
nor U9055 (N_9055,N_1312,N_1845);
and U9056 (N_9056,N_4806,N_5237);
and U9057 (N_9057,N_3059,N_1709);
or U9058 (N_9058,N_3754,N_743);
and U9059 (N_9059,N_2576,N_5186);
and U9060 (N_9060,N_80,N_1183);
nand U9061 (N_9061,N_1741,N_640);
or U9062 (N_9062,N_1848,N_5915);
and U9063 (N_9063,N_3456,N_5594);
and U9064 (N_9064,N_2949,N_5630);
nand U9065 (N_9065,N_625,N_4342);
or U9066 (N_9066,N_5016,N_1428);
nor U9067 (N_9067,N_606,N_1137);
xnor U9068 (N_9068,N_483,N_4915);
and U9069 (N_9069,N_2537,N_5761);
or U9070 (N_9070,N_2310,N_2241);
nand U9071 (N_9071,N_1599,N_190);
or U9072 (N_9072,N_226,N_1522);
and U9073 (N_9073,N_1995,N_5969);
or U9074 (N_9074,N_1784,N_5126);
nand U9075 (N_9075,N_1390,N_258);
xor U9076 (N_9076,N_2207,N_1370);
or U9077 (N_9077,N_5879,N_2800);
or U9078 (N_9078,N_4291,N_4651);
nand U9079 (N_9079,N_817,N_5685);
xnor U9080 (N_9080,N_3416,N_914);
nor U9081 (N_9081,N_1282,N_5372);
and U9082 (N_9082,N_3430,N_2670);
xnor U9083 (N_9083,N_168,N_2306);
xor U9084 (N_9084,N_945,N_3853);
or U9085 (N_9085,N_1683,N_3506);
nand U9086 (N_9086,N_1937,N_4153);
or U9087 (N_9087,N_4935,N_3850);
and U9088 (N_9088,N_1089,N_1165);
or U9089 (N_9089,N_3413,N_1267);
or U9090 (N_9090,N_2970,N_490);
and U9091 (N_9091,N_2218,N_588);
xnor U9092 (N_9092,N_4641,N_5105);
or U9093 (N_9093,N_1851,N_3399);
or U9094 (N_9094,N_3802,N_4714);
xor U9095 (N_9095,N_4995,N_4376);
nor U9096 (N_9096,N_4864,N_1048);
xor U9097 (N_9097,N_3141,N_4201);
nor U9098 (N_9098,N_2733,N_5940);
or U9099 (N_9099,N_1889,N_4594);
nor U9100 (N_9100,N_4144,N_52);
xor U9101 (N_9101,N_5750,N_5757);
and U9102 (N_9102,N_2921,N_2750);
nor U9103 (N_9103,N_2739,N_394);
or U9104 (N_9104,N_2510,N_1737);
nor U9105 (N_9105,N_1593,N_2832);
and U9106 (N_9106,N_4983,N_3099);
or U9107 (N_9107,N_2775,N_4015);
xor U9108 (N_9108,N_4658,N_1623);
or U9109 (N_9109,N_1646,N_4910);
and U9110 (N_9110,N_3746,N_3072);
xnor U9111 (N_9111,N_2963,N_4459);
nor U9112 (N_9112,N_524,N_4709);
or U9113 (N_9113,N_628,N_421);
and U9114 (N_9114,N_1019,N_3724);
or U9115 (N_9115,N_4072,N_613);
nand U9116 (N_9116,N_5510,N_3492);
xor U9117 (N_9117,N_2973,N_798);
nand U9118 (N_9118,N_5821,N_4314);
nand U9119 (N_9119,N_4013,N_4955);
and U9120 (N_9120,N_627,N_3393);
or U9121 (N_9121,N_3870,N_5998);
nor U9122 (N_9122,N_4842,N_2490);
nor U9123 (N_9123,N_2949,N_2883);
and U9124 (N_9124,N_1450,N_3433);
xnor U9125 (N_9125,N_1516,N_2463);
xnor U9126 (N_9126,N_2895,N_4136);
or U9127 (N_9127,N_5396,N_2770);
or U9128 (N_9128,N_526,N_2903);
xnor U9129 (N_9129,N_5888,N_590);
xor U9130 (N_9130,N_4414,N_5911);
and U9131 (N_9131,N_1227,N_2233);
xnor U9132 (N_9132,N_5338,N_2732);
xor U9133 (N_9133,N_573,N_5199);
xor U9134 (N_9134,N_5439,N_791);
and U9135 (N_9135,N_585,N_364);
nand U9136 (N_9136,N_3703,N_3444);
nand U9137 (N_9137,N_5072,N_1533);
xnor U9138 (N_9138,N_1658,N_2641);
nor U9139 (N_9139,N_831,N_4416);
nor U9140 (N_9140,N_3113,N_438);
nor U9141 (N_9141,N_4150,N_40);
xnor U9142 (N_9142,N_399,N_3294);
nand U9143 (N_9143,N_892,N_1070);
and U9144 (N_9144,N_5384,N_3585);
nor U9145 (N_9145,N_516,N_1431);
and U9146 (N_9146,N_2047,N_4853);
nand U9147 (N_9147,N_4107,N_1887);
nand U9148 (N_9148,N_2282,N_4850);
or U9149 (N_9149,N_2120,N_2793);
and U9150 (N_9150,N_689,N_5309);
or U9151 (N_9151,N_5274,N_4297);
xor U9152 (N_9152,N_245,N_507);
xor U9153 (N_9153,N_4469,N_1731);
and U9154 (N_9154,N_1063,N_5207);
nor U9155 (N_9155,N_2269,N_605);
or U9156 (N_9156,N_4334,N_2711);
and U9157 (N_9157,N_3851,N_3128);
or U9158 (N_9158,N_5613,N_1640);
nor U9159 (N_9159,N_3879,N_3442);
or U9160 (N_9160,N_4425,N_1686);
and U9161 (N_9161,N_1575,N_332);
or U9162 (N_9162,N_4761,N_1315);
and U9163 (N_9163,N_4906,N_4951);
and U9164 (N_9164,N_3080,N_4591);
xnor U9165 (N_9165,N_1475,N_3131);
nor U9166 (N_9166,N_3745,N_4855);
xnor U9167 (N_9167,N_3272,N_2641);
nand U9168 (N_9168,N_2099,N_5170);
xor U9169 (N_9169,N_2154,N_2305);
nor U9170 (N_9170,N_886,N_4318);
nand U9171 (N_9171,N_4018,N_4803);
or U9172 (N_9172,N_1245,N_5525);
nor U9173 (N_9173,N_1275,N_701);
nand U9174 (N_9174,N_5242,N_132);
nor U9175 (N_9175,N_5735,N_4559);
nand U9176 (N_9176,N_4713,N_5429);
xnor U9177 (N_9177,N_991,N_1563);
xor U9178 (N_9178,N_745,N_4143);
nand U9179 (N_9179,N_1372,N_1366);
xor U9180 (N_9180,N_4287,N_673);
nand U9181 (N_9181,N_4244,N_5000);
or U9182 (N_9182,N_5739,N_492);
nand U9183 (N_9183,N_5455,N_5053);
and U9184 (N_9184,N_4341,N_34);
and U9185 (N_9185,N_1613,N_2169);
or U9186 (N_9186,N_4402,N_2151);
or U9187 (N_9187,N_5449,N_2394);
and U9188 (N_9188,N_5358,N_5211);
xor U9189 (N_9189,N_4081,N_2633);
or U9190 (N_9190,N_445,N_3568);
xnor U9191 (N_9191,N_3939,N_4073);
or U9192 (N_9192,N_5280,N_5745);
nand U9193 (N_9193,N_3481,N_4778);
and U9194 (N_9194,N_1446,N_2273);
and U9195 (N_9195,N_1546,N_19);
nor U9196 (N_9196,N_5229,N_271);
nor U9197 (N_9197,N_307,N_3316);
and U9198 (N_9198,N_2195,N_2715);
nand U9199 (N_9199,N_5838,N_3123);
xnor U9200 (N_9200,N_2887,N_5725);
or U9201 (N_9201,N_5297,N_3428);
nor U9202 (N_9202,N_791,N_4290);
and U9203 (N_9203,N_3100,N_3376);
xor U9204 (N_9204,N_3992,N_5965);
xor U9205 (N_9205,N_2316,N_368);
nand U9206 (N_9206,N_4287,N_1677);
or U9207 (N_9207,N_2881,N_633);
and U9208 (N_9208,N_3470,N_4241);
and U9209 (N_9209,N_5445,N_5114);
or U9210 (N_9210,N_5910,N_3367);
xnor U9211 (N_9211,N_2630,N_1060);
and U9212 (N_9212,N_4554,N_2103);
nand U9213 (N_9213,N_4500,N_781);
nor U9214 (N_9214,N_2491,N_4115);
xnor U9215 (N_9215,N_669,N_3565);
xor U9216 (N_9216,N_2657,N_4939);
nand U9217 (N_9217,N_1573,N_4614);
nor U9218 (N_9218,N_310,N_910);
or U9219 (N_9219,N_4400,N_3915);
nand U9220 (N_9220,N_2703,N_845);
or U9221 (N_9221,N_728,N_2103);
and U9222 (N_9222,N_965,N_3604);
or U9223 (N_9223,N_5980,N_2559);
xnor U9224 (N_9224,N_5246,N_3430);
or U9225 (N_9225,N_334,N_3833);
xnor U9226 (N_9226,N_1873,N_4897);
nor U9227 (N_9227,N_4015,N_599);
or U9228 (N_9228,N_3750,N_1590);
nand U9229 (N_9229,N_4100,N_5647);
and U9230 (N_9230,N_3335,N_5506);
nor U9231 (N_9231,N_4204,N_1992);
nor U9232 (N_9232,N_3147,N_4342);
xor U9233 (N_9233,N_3273,N_2283);
xnor U9234 (N_9234,N_3475,N_5041);
nor U9235 (N_9235,N_1536,N_2617);
and U9236 (N_9236,N_68,N_1829);
or U9237 (N_9237,N_1417,N_600);
nor U9238 (N_9238,N_4928,N_5143);
nand U9239 (N_9239,N_3163,N_4861);
nand U9240 (N_9240,N_5318,N_1864);
nor U9241 (N_9241,N_112,N_2168);
nand U9242 (N_9242,N_4624,N_1634);
or U9243 (N_9243,N_2760,N_5551);
nand U9244 (N_9244,N_1097,N_5176);
nand U9245 (N_9245,N_1570,N_2799);
and U9246 (N_9246,N_684,N_4329);
nor U9247 (N_9247,N_4523,N_3154);
xor U9248 (N_9248,N_1305,N_3013);
nor U9249 (N_9249,N_5510,N_3652);
nor U9250 (N_9250,N_1722,N_3806);
and U9251 (N_9251,N_460,N_3411);
or U9252 (N_9252,N_4013,N_4068);
nor U9253 (N_9253,N_1780,N_4517);
or U9254 (N_9254,N_3011,N_84);
or U9255 (N_9255,N_3610,N_1449);
and U9256 (N_9256,N_1621,N_1558);
nand U9257 (N_9257,N_1921,N_172);
or U9258 (N_9258,N_3412,N_5032);
nor U9259 (N_9259,N_5019,N_3288);
nand U9260 (N_9260,N_171,N_759);
nand U9261 (N_9261,N_3041,N_1233);
and U9262 (N_9262,N_4579,N_1531);
xnor U9263 (N_9263,N_2702,N_4224);
nor U9264 (N_9264,N_5643,N_1010);
xor U9265 (N_9265,N_4056,N_559);
nand U9266 (N_9266,N_4032,N_829);
nor U9267 (N_9267,N_1003,N_4465);
xnor U9268 (N_9268,N_915,N_380);
nor U9269 (N_9269,N_4013,N_4072);
or U9270 (N_9270,N_5987,N_3089);
nor U9271 (N_9271,N_3217,N_2693);
nor U9272 (N_9272,N_5288,N_3453);
xor U9273 (N_9273,N_286,N_2914);
nor U9274 (N_9274,N_43,N_4206);
and U9275 (N_9275,N_5660,N_3052);
nor U9276 (N_9276,N_335,N_2217);
and U9277 (N_9277,N_894,N_1505);
nand U9278 (N_9278,N_4314,N_1339);
nand U9279 (N_9279,N_2996,N_1720);
xnor U9280 (N_9280,N_5291,N_812);
nand U9281 (N_9281,N_4127,N_2231);
and U9282 (N_9282,N_3958,N_5791);
or U9283 (N_9283,N_5460,N_1072);
and U9284 (N_9284,N_4721,N_4385);
nand U9285 (N_9285,N_4766,N_650);
xor U9286 (N_9286,N_3823,N_4240);
and U9287 (N_9287,N_1467,N_1963);
nand U9288 (N_9288,N_4676,N_5120);
nor U9289 (N_9289,N_5467,N_2613);
nand U9290 (N_9290,N_215,N_2104);
nand U9291 (N_9291,N_341,N_3818);
nand U9292 (N_9292,N_953,N_5914);
nand U9293 (N_9293,N_2353,N_2579);
and U9294 (N_9294,N_5976,N_1516);
or U9295 (N_9295,N_201,N_5312);
or U9296 (N_9296,N_4020,N_202);
or U9297 (N_9297,N_3735,N_2436);
and U9298 (N_9298,N_2630,N_3070);
nor U9299 (N_9299,N_2111,N_3027);
nor U9300 (N_9300,N_5308,N_1427);
nor U9301 (N_9301,N_1313,N_3084);
and U9302 (N_9302,N_3447,N_2820);
xnor U9303 (N_9303,N_3294,N_4920);
or U9304 (N_9304,N_1404,N_5935);
and U9305 (N_9305,N_5636,N_5138);
and U9306 (N_9306,N_4836,N_2594);
nor U9307 (N_9307,N_4819,N_2652);
or U9308 (N_9308,N_2151,N_5239);
or U9309 (N_9309,N_2538,N_5740);
and U9310 (N_9310,N_3158,N_1200);
nand U9311 (N_9311,N_386,N_2318);
nand U9312 (N_9312,N_5290,N_2585);
nand U9313 (N_9313,N_5463,N_1619);
and U9314 (N_9314,N_3116,N_1315);
xnor U9315 (N_9315,N_3544,N_2340);
nand U9316 (N_9316,N_1023,N_2243);
nor U9317 (N_9317,N_2844,N_2964);
xnor U9318 (N_9318,N_195,N_5755);
and U9319 (N_9319,N_77,N_277);
nor U9320 (N_9320,N_816,N_4214);
nand U9321 (N_9321,N_3514,N_3532);
nor U9322 (N_9322,N_3219,N_4);
nor U9323 (N_9323,N_2536,N_4117);
and U9324 (N_9324,N_2016,N_3787);
nand U9325 (N_9325,N_1636,N_859);
xnor U9326 (N_9326,N_3572,N_851);
or U9327 (N_9327,N_2930,N_2097);
nand U9328 (N_9328,N_5405,N_3636);
nor U9329 (N_9329,N_3763,N_5553);
nand U9330 (N_9330,N_286,N_1945);
nand U9331 (N_9331,N_304,N_4540);
or U9332 (N_9332,N_5360,N_3074);
nor U9333 (N_9333,N_1985,N_3462);
or U9334 (N_9334,N_4134,N_860);
and U9335 (N_9335,N_2812,N_696);
or U9336 (N_9336,N_4716,N_190);
or U9337 (N_9337,N_5369,N_5278);
xnor U9338 (N_9338,N_5330,N_1350);
nand U9339 (N_9339,N_3842,N_5268);
and U9340 (N_9340,N_4579,N_1501);
xor U9341 (N_9341,N_3157,N_2514);
nand U9342 (N_9342,N_1065,N_4333);
or U9343 (N_9343,N_5953,N_4337);
or U9344 (N_9344,N_710,N_4518);
xnor U9345 (N_9345,N_1157,N_2488);
or U9346 (N_9346,N_5166,N_1302);
and U9347 (N_9347,N_1600,N_175);
and U9348 (N_9348,N_678,N_5585);
nor U9349 (N_9349,N_444,N_5976);
or U9350 (N_9350,N_5614,N_146);
and U9351 (N_9351,N_4967,N_1104);
nand U9352 (N_9352,N_4892,N_1603);
and U9353 (N_9353,N_4261,N_4053);
or U9354 (N_9354,N_4190,N_3430);
nand U9355 (N_9355,N_2155,N_3403);
nor U9356 (N_9356,N_5770,N_4637);
or U9357 (N_9357,N_3793,N_5260);
nor U9358 (N_9358,N_181,N_316);
nand U9359 (N_9359,N_4576,N_2905);
xnor U9360 (N_9360,N_5835,N_836);
and U9361 (N_9361,N_1048,N_1885);
and U9362 (N_9362,N_2941,N_3069);
nor U9363 (N_9363,N_3051,N_4514);
xnor U9364 (N_9364,N_3772,N_5823);
xnor U9365 (N_9365,N_1751,N_2020);
or U9366 (N_9366,N_926,N_5540);
and U9367 (N_9367,N_3616,N_1092);
and U9368 (N_9368,N_391,N_3087);
xnor U9369 (N_9369,N_292,N_5558);
nor U9370 (N_9370,N_1723,N_5216);
or U9371 (N_9371,N_4420,N_3186);
nor U9372 (N_9372,N_3360,N_2855);
nand U9373 (N_9373,N_178,N_359);
xor U9374 (N_9374,N_1691,N_4728);
nor U9375 (N_9375,N_674,N_4272);
nand U9376 (N_9376,N_3942,N_5012);
nor U9377 (N_9377,N_5156,N_2519);
xor U9378 (N_9378,N_22,N_4780);
nand U9379 (N_9379,N_1137,N_4333);
nand U9380 (N_9380,N_4106,N_2765);
or U9381 (N_9381,N_844,N_221);
and U9382 (N_9382,N_2186,N_3173);
and U9383 (N_9383,N_3757,N_179);
and U9384 (N_9384,N_986,N_340);
nor U9385 (N_9385,N_3226,N_1334);
and U9386 (N_9386,N_5735,N_3549);
or U9387 (N_9387,N_2335,N_2537);
or U9388 (N_9388,N_2114,N_3946);
and U9389 (N_9389,N_701,N_1849);
or U9390 (N_9390,N_4887,N_3763);
nor U9391 (N_9391,N_4263,N_2684);
xnor U9392 (N_9392,N_4129,N_3907);
nand U9393 (N_9393,N_1412,N_1341);
nand U9394 (N_9394,N_1932,N_3996);
or U9395 (N_9395,N_4823,N_2042);
or U9396 (N_9396,N_413,N_5135);
or U9397 (N_9397,N_5053,N_5844);
or U9398 (N_9398,N_3681,N_4045);
nand U9399 (N_9399,N_1175,N_5252);
nor U9400 (N_9400,N_2155,N_3053);
or U9401 (N_9401,N_4872,N_591);
nand U9402 (N_9402,N_3737,N_5366);
and U9403 (N_9403,N_5587,N_2173);
and U9404 (N_9404,N_2083,N_1157);
nor U9405 (N_9405,N_2541,N_1535);
and U9406 (N_9406,N_5949,N_3395);
nand U9407 (N_9407,N_2266,N_2373);
and U9408 (N_9408,N_867,N_2934);
or U9409 (N_9409,N_2799,N_770);
or U9410 (N_9410,N_2315,N_5587);
nor U9411 (N_9411,N_1941,N_3478);
nand U9412 (N_9412,N_1725,N_4866);
xnor U9413 (N_9413,N_517,N_2255);
xor U9414 (N_9414,N_959,N_3170);
xor U9415 (N_9415,N_4369,N_1334);
and U9416 (N_9416,N_1515,N_1482);
nand U9417 (N_9417,N_5775,N_3854);
xor U9418 (N_9418,N_1585,N_5391);
nor U9419 (N_9419,N_5962,N_750);
xor U9420 (N_9420,N_750,N_4702);
xor U9421 (N_9421,N_4348,N_5871);
xnor U9422 (N_9422,N_4767,N_3314);
and U9423 (N_9423,N_5986,N_4358);
and U9424 (N_9424,N_898,N_4671);
or U9425 (N_9425,N_4338,N_5037);
nand U9426 (N_9426,N_2817,N_4444);
or U9427 (N_9427,N_3775,N_2463);
and U9428 (N_9428,N_4542,N_1309);
xnor U9429 (N_9429,N_1263,N_4884);
and U9430 (N_9430,N_2476,N_2916);
or U9431 (N_9431,N_4117,N_233);
nor U9432 (N_9432,N_1498,N_5428);
nor U9433 (N_9433,N_2915,N_3946);
xnor U9434 (N_9434,N_3140,N_1254);
xnor U9435 (N_9435,N_4710,N_4155);
nor U9436 (N_9436,N_1459,N_1536);
or U9437 (N_9437,N_4971,N_4912);
or U9438 (N_9438,N_4635,N_3000);
xnor U9439 (N_9439,N_168,N_4324);
nor U9440 (N_9440,N_1479,N_5832);
nor U9441 (N_9441,N_2607,N_2857);
xor U9442 (N_9442,N_5303,N_4033);
and U9443 (N_9443,N_940,N_5281);
nand U9444 (N_9444,N_731,N_27);
and U9445 (N_9445,N_2895,N_3945);
xor U9446 (N_9446,N_4093,N_4866);
xor U9447 (N_9447,N_2467,N_2876);
and U9448 (N_9448,N_4026,N_4658);
or U9449 (N_9449,N_1045,N_5484);
and U9450 (N_9450,N_693,N_4914);
or U9451 (N_9451,N_2277,N_4243);
and U9452 (N_9452,N_3111,N_2593);
nand U9453 (N_9453,N_2643,N_2448);
and U9454 (N_9454,N_5980,N_4914);
nor U9455 (N_9455,N_1893,N_3770);
xor U9456 (N_9456,N_206,N_1453);
nand U9457 (N_9457,N_4637,N_5311);
nor U9458 (N_9458,N_3693,N_3124);
xor U9459 (N_9459,N_4044,N_2250);
xor U9460 (N_9460,N_4079,N_3445);
or U9461 (N_9461,N_4972,N_2475);
or U9462 (N_9462,N_1499,N_3132);
nand U9463 (N_9463,N_4418,N_364);
or U9464 (N_9464,N_3330,N_5528);
and U9465 (N_9465,N_1806,N_2884);
xnor U9466 (N_9466,N_3687,N_4039);
or U9467 (N_9467,N_1856,N_3497);
or U9468 (N_9468,N_3298,N_996);
nor U9469 (N_9469,N_1841,N_5758);
or U9470 (N_9470,N_2460,N_3924);
or U9471 (N_9471,N_4662,N_4041);
xor U9472 (N_9472,N_3484,N_993);
nor U9473 (N_9473,N_631,N_420);
or U9474 (N_9474,N_5495,N_1793);
nand U9475 (N_9475,N_3494,N_1247);
nand U9476 (N_9476,N_4101,N_554);
or U9477 (N_9477,N_4865,N_3921);
xor U9478 (N_9478,N_1274,N_3957);
or U9479 (N_9479,N_3884,N_347);
or U9480 (N_9480,N_5392,N_3462);
xnor U9481 (N_9481,N_4367,N_5908);
and U9482 (N_9482,N_5612,N_1072);
nor U9483 (N_9483,N_692,N_5125);
and U9484 (N_9484,N_2853,N_5395);
nand U9485 (N_9485,N_2,N_161);
and U9486 (N_9486,N_1172,N_2471);
xnor U9487 (N_9487,N_1484,N_4232);
xnor U9488 (N_9488,N_4958,N_5594);
nor U9489 (N_9489,N_1889,N_83);
or U9490 (N_9490,N_2489,N_4509);
and U9491 (N_9491,N_3674,N_1644);
and U9492 (N_9492,N_2033,N_4970);
nor U9493 (N_9493,N_3197,N_4082);
and U9494 (N_9494,N_5955,N_3755);
nor U9495 (N_9495,N_1063,N_1152);
nor U9496 (N_9496,N_3053,N_5774);
and U9497 (N_9497,N_5339,N_323);
xor U9498 (N_9498,N_4668,N_4266);
xor U9499 (N_9499,N_5080,N_1601);
nand U9500 (N_9500,N_4892,N_2365);
or U9501 (N_9501,N_3951,N_4647);
nand U9502 (N_9502,N_937,N_927);
and U9503 (N_9503,N_2568,N_386);
and U9504 (N_9504,N_56,N_1440);
nor U9505 (N_9505,N_1301,N_3417);
and U9506 (N_9506,N_5595,N_2414);
nand U9507 (N_9507,N_934,N_4220);
and U9508 (N_9508,N_3116,N_944);
nor U9509 (N_9509,N_3719,N_2157);
nand U9510 (N_9510,N_1738,N_5625);
and U9511 (N_9511,N_338,N_3511);
nand U9512 (N_9512,N_3136,N_2384);
nand U9513 (N_9513,N_3409,N_3524);
nand U9514 (N_9514,N_842,N_220);
xor U9515 (N_9515,N_3577,N_2712);
and U9516 (N_9516,N_2990,N_5565);
or U9517 (N_9517,N_4544,N_5259);
or U9518 (N_9518,N_230,N_1495);
xor U9519 (N_9519,N_2975,N_1428);
nand U9520 (N_9520,N_5412,N_3522);
and U9521 (N_9521,N_344,N_293);
nand U9522 (N_9522,N_5644,N_4195);
nand U9523 (N_9523,N_471,N_5138);
nand U9524 (N_9524,N_4407,N_4450);
or U9525 (N_9525,N_4854,N_5961);
and U9526 (N_9526,N_3383,N_491);
nand U9527 (N_9527,N_1064,N_1276);
nor U9528 (N_9528,N_442,N_4101);
or U9529 (N_9529,N_3915,N_5054);
and U9530 (N_9530,N_811,N_1564);
nor U9531 (N_9531,N_1792,N_5950);
nand U9532 (N_9532,N_3438,N_5410);
nor U9533 (N_9533,N_2664,N_2674);
nor U9534 (N_9534,N_3385,N_3827);
nor U9535 (N_9535,N_2883,N_3403);
nand U9536 (N_9536,N_5464,N_4127);
nand U9537 (N_9537,N_1389,N_4229);
nor U9538 (N_9538,N_5945,N_5986);
nor U9539 (N_9539,N_4608,N_2461);
nor U9540 (N_9540,N_5585,N_1301);
nand U9541 (N_9541,N_385,N_2497);
or U9542 (N_9542,N_4114,N_1356);
or U9543 (N_9543,N_2028,N_2641);
xnor U9544 (N_9544,N_5073,N_2223);
and U9545 (N_9545,N_38,N_2000);
nand U9546 (N_9546,N_2921,N_142);
nand U9547 (N_9547,N_602,N_0);
nand U9548 (N_9548,N_4134,N_2223);
nand U9549 (N_9549,N_2138,N_5128);
and U9550 (N_9550,N_5728,N_3812);
nand U9551 (N_9551,N_3904,N_1835);
nor U9552 (N_9552,N_2504,N_258);
and U9553 (N_9553,N_4891,N_4631);
xor U9554 (N_9554,N_1376,N_5731);
and U9555 (N_9555,N_4132,N_4694);
xnor U9556 (N_9556,N_1207,N_2605);
or U9557 (N_9557,N_4940,N_4972);
nor U9558 (N_9558,N_5425,N_3852);
or U9559 (N_9559,N_4884,N_1913);
nand U9560 (N_9560,N_642,N_1178);
nand U9561 (N_9561,N_1000,N_3420);
nand U9562 (N_9562,N_3047,N_3923);
and U9563 (N_9563,N_578,N_4388);
and U9564 (N_9564,N_4321,N_681);
nand U9565 (N_9565,N_5391,N_2454);
nand U9566 (N_9566,N_1156,N_4310);
nor U9567 (N_9567,N_226,N_4867);
xnor U9568 (N_9568,N_800,N_4969);
or U9569 (N_9569,N_3349,N_4008);
or U9570 (N_9570,N_2790,N_1995);
or U9571 (N_9571,N_1067,N_48);
xor U9572 (N_9572,N_112,N_1878);
and U9573 (N_9573,N_4374,N_1182);
and U9574 (N_9574,N_1431,N_3389);
nand U9575 (N_9575,N_3169,N_1368);
nand U9576 (N_9576,N_3874,N_2102);
xor U9577 (N_9577,N_3409,N_2012);
and U9578 (N_9578,N_3247,N_1315);
xor U9579 (N_9579,N_2296,N_2575);
xor U9580 (N_9580,N_5294,N_3627);
nand U9581 (N_9581,N_4225,N_2421);
nand U9582 (N_9582,N_1476,N_3805);
nor U9583 (N_9583,N_3382,N_3494);
nand U9584 (N_9584,N_1423,N_2728);
xor U9585 (N_9585,N_4770,N_4283);
nor U9586 (N_9586,N_546,N_5186);
and U9587 (N_9587,N_1125,N_530);
and U9588 (N_9588,N_1781,N_103);
nor U9589 (N_9589,N_2371,N_3362);
xnor U9590 (N_9590,N_2941,N_5078);
xor U9591 (N_9591,N_2428,N_1788);
nand U9592 (N_9592,N_5261,N_1808);
and U9593 (N_9593,N_2469,N_1024);
and U9594 (N_9594,N_1332,N_5727);
xor U9595 (N_9595,N_2863,N_3794);
and U9596 (N_9596,N_5391,N_2918);
nand U9597 (N_9597,N_306,N_1086);
or U9598 (N_9598,N_557,N_5990);
and U9599 (N_9599,N_1042,N_2013);
nor U9600 (N_9600,N_2529,N_999);
xor U9601 (N_9601,N_5317,N_972);
or U9602 (N_9602,N_5435,N_4140);
and U9603 (N_9603,N_3124,N_1215);
nor U9604 (N_9604,N_5299,N_2923);
or U9605 (N_9605,N_2764,N_1171);
and U9606 (N_9606,N_497,N_3831);
nand U9607 (N_9607,N_5097,N_4090);
nor U9608 (N_9608,N_3435,N_262);
nor U9609 (N_9609,N_4103,N_2401);
nand U9610 (N_9610,N_848,N_2216);
xor U9611 (N_9611,N_3326,N_2068);
xnor U9612 (N_9612,N_3996,N_5563);
and U9613 (N_9613,N_1224,N_110);
xnor U9614 (N_9614,N_3345,N_2480);
nand U9615 (N_9615,N_3135,N_1083);
nand U9616 (N_9616,N_1435,N_5974);
xor U9617 (N_9617,N_4828,N_41);
or U9618 (N_9618,N_2272,N_4905);
or U9619 (N_9619,N_2681,N_2610);
and U9620 (N_9620,N_3103,N_5507);
xor U9621 (N_9621,N_20,N_4354);
nand U9622 (N_9622,N_726,N_4794);
nand U9623 (N_9623,N_3529,N_5371);
and U9624 (N_9624,N_4817,N_3849);
and U9625 (N_9625,N_5599,N_5398);
or U9626 (N_9626,N_362,N_1017);
nand U9627 (N_9627,N_4394,N_2527);
nor U9628 (N_9628,N_4637,N_2460);
or U9629 (N_9629,N_3468,N_2471);
nand U9630 (N_9630,N_3467,N_5326);
xor U9631 (N_9631,N_3858,N_4138);
nand U9632 (N_9632,N_4131,N_47);
nor U9633 (N_9633,N_4641,N_305);
xor U9634 (N_9634,N_4542,N_952);
or U9635 (N_9635,N_5910,N_3717);
xnor U9636 (N_9636,N_767,N_5626);
nor U9637 (N_9637,N_1813,N_1226);
or U9638 (N_9638,N_3743,N_342);
nor U9639 (N_9639,N_2146,N_2752);
or U9640 (N_9640,N_5381,N_5102);
xor U9641 (N_9641,N_4871,N_2315);
xor U9642 (N_9642,N_1208,N_4000);
and U9643 (N_9643,N_3036,N_2903);
xnor U9644 (N_9644,N_2073,N_2667);
or U9645 (N_9645,N_4643,N_951);
nor U9646 (N_9646,N_3006,N_3186);
or U9647 (N_9647,N_3733,N_5765);
or U9648 (N_9648,N_525,N_640);
nand U9649 (N_9649,N_5024,N_5548);
nor U9650 (N_9650,N_1748,N_4077);
xnor U9651 (N_9651,N_4411,N_5569);
xor U9652 (N_9652,N_2386,N_1053);
or U9653 (N_9653,N_3464,N_5189);
xor U9654 (N_9654,N_1168,N_1815);
xnor U9655 (N_9655,N_2775,N_4241);
nand U9656 (N_9656,N_5744,N_3822);
nand U9657 (N_9657,N_2521,N_4053);
or U9658 (N_9658,N_1707,N_4495);
nor U9659 (N_9659,N_3032,N_187);
nand U9660 (N_9660,N_1682,N_2488);
or U9661 (N_9661,N_1259,N_2995);
xnor U9662 (N_9662,N_4463,N_5832);
or U9663 (N_9663,N_3620,N_1896);
nor U9664 (N_9664,N_573,N_3826);
and U9665 (N_9665,N_460,N_5508);
nand U9666 (N_9666,N_4312,N_2927);
nand U9667 (N_9667,N_197,N_2611);
nor U9668 (N_9668,N_720,N_3562);
and U9669 (N_9669,N_4137,N_3788);
nor U9670 (N_9670,N_2490,N_5312);
or U9671 (N_9671,N_279,N_917);
xor U9672 (N_9672,N_3443,N_2008);
nand U9673 (N_9673,N_2371,N_3522);
xor U9674 (N_9674,N_5577,N_3770);
and U9675 (N_9675,N_5366,N_707);
nand U9676 (N_9676,N_3470,N_1917);
nor U9677 (N_9677,N_4854,N_1420);
or U9678 (N_9678,N_377,N_5111);
and U9679 (N_9679,N_180,N_3604);
or U9680 (N_9680,N_4437,N_2009);
or U9681 (N_9681,N_460,N_3521);
and U9682 (N_9682,N_5923,N_2534);
and U9683 (N_9683,N_5171,N_919);
xor U9684 (N_9684,N_4858,N_5136);
nor U9685 (N_9685,N_4910,N_2617);
or U9686 (N_9686,N_2704,N_790);
nor U9687 (N_9687,N_5084,N_436);
xor U9688 (N_9688,N_2110,N_981);
and U9689 (N_9689,N_1429,N_4453);
nand U9690 (N_9690,N_2132,N_2202);
nor U9691 (N_9691,N_888,N_3903);
nor U9692 (N_9692,N_4242,N_2430);
or U9693 (N_9693,N_1573,N_762);
and U9694 (N_9694,N_3615,N_2299);
nor U9695 (N_9695,N_3692,N_3077);
xnor U9696 (N_9696,N_414,N_5351);
nor U9697 (N_9697,N_5196,N_1105);
or U9698 (N_9698,N_4065,N_228);
nor U9699 (N_9699,N_1834,N_362);
xor U9700 (N_9700,N_2465,N_3519);
nor U9701 (N_9701,N_2967,N_2058);
or U9702 (N_9702,N_3509,N_1154);
nand U9703 (N_9703,N_1993,N_1278);
or U9704 (N_9704,N_1736,N_4524);
or U9705 (N_9705,N_5240,N_3915);
or U9706 (N_9706,N_5280,N_2367);
nand U9707 (N_9707,N_5695,N_2251);
and U9708 (N_9708,N_2665,N_403);
xor U9709 (N_9709,N_2608,N_2771);
nand U9710 (N_9710,N_1588,N_4398);
or U9711 (N_9711,N_4906,N_4205);
or U9712 (N_9712,N_4512,N_3785);
and U9713 (N_9713,N_4978,N_1066);
or U9714 (N_9714,N_1379,N_4924);
nand U9715 (N_9715,N_366,N_1373);
nand U9716 (N_9716,N_325,N_5282);
nand U9717 (N_9717,N_2441,N_4960);
and U9718 (N_9718,N_3058,N_2615);
nor U9719 (N_9719,N_2900,N_3021);
and U9720 (N_9720,N_4222,N_2119);
nand U9721 (N_9721,N_1792,N_3319);
and U9722 (N_9722,N_1807,N_232);
xor U9723 (N_9723,N_5215,N_3331);
and U9724 (N_9724,N_5809,N_5674);
and U9725 (N_9725,N_2797,N_2615);
xnor U9726 (N_9726,N_4192,N_2026);
nand U9727 (N_9727,N_5844,N_209);
and U9728 (N_9728,N_1014,N_4390);
or U9729 (N_9729,N_5803,N_1777);
nand U9730 (N_9730,N_32,N_1355);
or U9731 (N_9731,N_1694,N_5022);
or U9732 (N_9732,N_3856,N_5532);
nand U9733 (N_9733,N_1852,N_3041);
or U9734 (N_9734,N_1415,N_4238);
xnor U9735 (N_9735,N_3651,N_778);
and U9736 (N_9736,N_1792,N_5123);
or U9737 (N_9737,N_2956,N_5807);
or U9738 (N_9738,N_1434,N_2324);
nor U9739 (N_9739,N_5466,N_1917);
or U9740 (N_9740,N_4873,N_642);
or U9741 (N_9741,N_3939,N_1650);
or U9742 (N_9742,N_5679,N_1841);
or U9743 (N_9743,N_2997,N_3137);
and U9744 (N_9744,N_624,N_1987);
nor U9745 (N_9745,N_5373,N_2764);
and U9746 (N_9746,N_2505,N_1738);
xnor U9747 (N_9747,N_812,N_1099);
xnor U9748 (N_9748,N_575,N_1974);
and U9749 (N_9749,N_560,N_3323);
xnor U9750 (N_9750,N_686,N_927);
and U9751 (N_9751,N_1884,N_3293);
nand U9752 (N_9752,N_728,N_3302);
and U9753 (N_9753,N_5462,N_2792);
xnor U9754 (N_9754,N_1093,N_5323);
nor U9755 (N_9755,N_2444,N_1991);
nand U9756 (N_9756,N_2203,N_2206);
or U9757 (N_9757,N_4131,N_5012);
nand U9758 (N_9758,N_4836,N_2675);
and U9759 (N_9759,N_3578,N_2613);
nand U9760 (N_9760,N_628,N_5045);
and U9761 (N_9761,N_4015,N_3359);
xnor U9762 (N_9762,N_4766,N_5244);
xor U9763 (N_9763,N_1962,N_4349);
nand U9764 (N_9764,N_5970,N_3706);
xor U9765 (N_9765,N_3425,N_682);
nand U9766 (N_9766,N_663,N_2427);
and U9767 (N_9767,N_4692,N_5697);
or U9768 (N_9768,N_4495,N_913);
nor U9769 (N_9769,N_3876,N_1776);
nand U9770 (N_9770,N_3915,N_3027);
and U9771 (N_9771,N_5720,N_3940);
or U9772 (N_9772,N_2221,N_2985);
or U9773 (N_9773,N_374,N_3518);
nor U9774 (N_9774,N_11,N_5274);
and U9775 (N_9775,N_5942,N_187);
nand U9776 (N_9776,N_2596,N_4275);
nand U9777 (N_9777,N_1674,N_5856);
xnor U9778 (N_9778,N_5828,N_2481);
or U9779 (N_9779,N_406,N_5180);
or U9780 (N_9780,N_460,N_2980);
nand U9781 (N_9781,N_4638,N_5307);
and U9782 (N_9782,N_1467,N_2536);
nand U9783 (N_9783,N_3456,N_3409);
xnor U9784 (N_9784,N_3884,N_4141);
or U9785 (N_9785,N_1804,N_5217);
and U9786 (N_9786,N_2349,N_5480);
or U9787 (N_9787,N_1497,N_5679);
xor U9788 (N_9788,N_1231,N_677);
or U9789 (N_9789,N_5695,N_4984);
xnor U9790 (N_9790,N_1701,N_989);
and U9791 (N_9791,N_306,N_4007);
nor U9792 (N_9792,N_1631,N_238);
and U9793 (N_9793,N_3197,N_3279);
xor U9794 (N_9794,N_2742,N_4271);
or U9795 (N_9795,N_1349,N_3436);
xnor U9796 (N_9796,N_2453,N_5154);
nor U9797 (N_9797,N_4811,N_63);
nor U9798 (N_9798,N_3664,N_4672);
or U9799 (N_9799,N_3045,N_4464);
xor U9800 (N_9800,N_2108,N_4355);
or U9801 (N_9801,N_2018,N_2368);
and U9802 (N_9802,N_1731,N_4004);
xnor U9803 (N_9803,N_3654,N_2501);
and U9804 (N_9804,N_4372,N_2890);
and U9805 (N_9805,N_3243,N_4764);
xor U9806 (N_9806,N_3559,N_1650);
or U9807 (N_9807,N_1242,N_4189);
nand U9808 (N_9808,N_233,N_3560);
and U9809 (N_9809,N_1146,N_5808);
nand U9810 (N_9810,N_3268,N_1338);
nand U9811 (N_9811,N_296,N_5560);
nand U9812 (N_9812,N_4683,N_4464);
and U9813 (N_9813,N_292,N_5169);
nor U9814 (N_9814,N_1870,N_4991);
xor U9815 (N_9815,N_3651,N_2688);
and U9816 (N_9816,N_2951,N_2853);
nor U9817 (N_9817,N_5716,N_5549);
and U9818 (N_9818,N_993,N_1861);
and U9819 (N_9819,N_889,N_809);
nor U9820 (N_9820,N_1540,N_3841);
and U9821 (N_9821,N_1762,N_5770);
nor U9822 (N_9822,N_897,N_4578);
xor U9823 (N_9823,N_384,N_5144);
and U9824 (N_9824,N_1986,N_4961);
nor U9825 (N_9825,N_4297,N_5564);
and U9826 (N_9826,N_2079,N_3464);
xor U9827 (N_9827,N_2781,N_5230);
xor U9828 (N_9828,N_5225,N_476);
nand U9829 (N_9829,N_2714,N_3653);
nor U9830 (N_9830,N_3811,N_2696);
xor U9831 (N_9831,N_1595,N_981);
and U9832 (N_9832,N_2573,N_2359);
and U9833 (N_9833,N_3948,N_4631);
nand U9834 (N_9834,N_1473,N_3493);
xor U9835 (N_9835,N_782,N_2010);
nor U9836 (N_9836,N_4092,N_2304);
or U9837 (N_9837,N_4367,N_4286);
and U9838 (N_9838,N_2705,N_5577);
and U9839 (N_9839,N_1070,N_371);
or U9840 (N_9840,N_2004,N_5071);
nand U9841 (N_9841,N_4403,N_3940);
and U9842 (N_9842,N_1705,N_5907);
xor U9843 (N_9843,N_220,N_85);
and U9844 (N_9844,N_1936,N_3902);
nor U9845 (N_9845,N_3580,N_777);
and U9846 (N_9846,N_5864,N_3433);
or U9847 (N_9847,N_2603,N_1230);
nand U9848 (N_9848,N_5733,N_2627);
and U9849 (N_9849,N_5493,N_656);
nor U9850 (N_9850,N_2206,N_4766);
nor U9851 (N_9851,N_810,N_4209);
nand U9852 (N_9852,N_4560,N_717);
and U9853 (N_9853,N_3587,N_5074);
nand U9854 (N_9854,N_222,N_5601);
xnor U9855 (N_9855,N_1610,N_3715);
nor U9856 (N_9856,N_5750,N_1974);
or U9857 (N_9857,N_1452,N_4394);
nor U9858 (N_9858,N_5398,N_3442);
nor U9859 (N_9859,N_5970,N_2277);
nand U9860 (N_9860,N_1914,N_2970);
and U9861 (N_9861,N_1154,N_3345);
or U9862 (N_9862,N_5357,N_2907);
nand U9863 (N_9863,N_2842,N_5890);
and U9864 (N_9864,N_4552,N_3398);
nor U9865 (N_9865,N_4403,N_3852);
or U9866 (N_9866,N_5039,N_5378);
and U9867 (N_9867,N_5876,N_3599);
xor U9868 (N_9868,N_2560,N_3916);
nor U9869 (N_9869,N_4985,N_1985);
nor U9870 (N_9870,N_4320,N_3780);
nand U9871 (N_9871,N_651,N_1677);
nor U9872 (N_9872,N_2953,N_1558);
xnor U9873 (N_9873,N_2220,N_5641);
xor U9874 (N_9874,N_2038,N_402);
nor U9875 (N_9875,N_5601,N_3240);
and U9876 (N_9876,N_3046,N_3411);
or U9877 (N_9877,N_3860,N_5713);
and U9878 (N_9878,N_2028,N_1154);
xnor U9879 (N_9879,N_3373,N_5503);
nor U9880 (N_9880,N_3591,N_923);
nand U9881 (N_9881,N_4193,N_3044);
nand U9882 (N_9882,N_1139,N_1533);
and U9883 (N_9883,N_4991,N_500);
or U9884 (N_9884,N_1557,N_2757);
xnor U9885 (N_9885,N_4410,N_2190);
and U9886 (N_9886,N_3462,N_1446);
nand U9887 (N_9887,N_2719,N_5581);
and U9888 (N_9888,N_4795,N_3465);
xor U9889 (N_9889,N_1203,N_407);
nand U9890 (N_9890,N_703,N_2234);
xnor U9891 (N_9891,N_3057,N_2417);
and U9892 (N_9892,N_2545,N_4797);
nand U9893 (N_9893,N_5474,N_2058);
or U9894 (N_9894,N_4580,N_685);
xnor U9895 (N_9895,N_3453,N_2836);
or U9896 (N_9896,N_4471,N_446);
nand U9897 (N_9897,N_3272,N_5206);
nand U9898 (N_9898,N_343,N_5150);
and U9899 (N_9899,N_3991,N_790);
or U9900 (N_9900,N_4210,N_3534);
or U9901 (N_9901,N_5284,N_5753);
xor U9902 (N_9902,N_2275,N_5384);
nor U9903 (N_9903,N_5478,N_4122);
xnor U9904 (N_9904,N_1954,N_3624);
and U9905 (N_9905,N_1849,N_3752);
and U9906 (N_9906,N_3436,N_3405);
and U9907 (N_9907,N_3356,N_5749);
or U9908 (N_9908,N_4297,N_1026);
nand U9909 (N_9909,N_1100,N_4070);
nand U9910 (N_9910,N_1958,N_4190);
nor U9911 (N_9911,N_2311,N_1674);
and U9912 (N_9912,N_1937,N_5082);
xnor U9913 (N_9913,N_5345,N_1391);
or U9914 (N_9914,N_5443,N_2936);
or U9915 (N_9915,N_5953,N_5439);
nand U9916 (N_9916,N_4141,N_3068);
nor U9917 (N_9917,N_5351,N_4860);
and U9918 (N_9918,N_1061,N_1752);
nand U9919 (N_9919,N_195,N_2146);
nor U9920 (N_9920,N_986,N_4242);
or U9921 (N_9921,N_347,N_1949);
xnor U9922 (N_9922,N_1163,N_1824);
nand U9923 (N_9923,N_5038,N_5868);
xor U9924 (N_9924,N_2,N_5949);
nand U9925 (N_9925,N_3599,N_2800);
xnor U9926 (N_9926,N_348,N_932);
xnor U9927 (N_9927,N_4289,N_339);
or U9928 (N_9928,N_2975,N_584);
and U9929 (N_9929,N_1438,N_2943);
xnor U9930 (N_9930,N_4571,N_2488);
xor U9931 (N_9931,N_5271,N_329);
nand U9932 (N_9932,N_3522,N_1893);
and U9933 (N_9933,N_606,N_3915);
and U9934 (N_9934,N_883,N_176);
or U9935 (N_9935,N_1721,N_1251);
and U9936 (N_9936,N_4458,N_4918);
nor U9937 (N_9937,N_810,N_2497);
xor U9938 (N_9938,N_474,N_1153);
and U9939 (N_9939,N_5568,N_3800);
and U9940 (N_9940,N_952,N_4110);
nand U9941 (N_9941,N_5875,N_3387);
and U9942 (N_9942,N_5228,N_382);
xnor U9943 (N_9943,N_4620,N_3838);
xnor U9944 (N_9944,N_2462,N_3772);
nand U9945 (N_9945,N_3706,N_3548);
nand U9946 (N_9946,N_5947,N_976);
xnor U9947 (N_9947,N_1354,N_4002);
nor U9948 (N_9948,N_5659,N_5819);
nand U9949 (N_9949,N_5848,N_510);
xor U9950 (N_9950,N_5041,N_3567);
nand U9951 (N_9951,N_2771,N_5900);
nand U9952 (N_9952,N_5908,N_3154);
or U9953 (N_9953,N_3831,N_3458);
nor U9954 (N_9954,N_2692,N_3198);
nor U9955 (N_9955,N_197,N_4567);
nor U9956 (N_9956,N_3300,N_624);
or U9957 (N_9957,N_5097,N_1750);
xor U9958 (N_9958,N_3158,N_913);
nor U9959 (N_9959,N_586,N_1800);
or U9960 (N_9960,N_5591,N_315);
nor U9961 (N_9961,N_3301,N_4183);
nand U9962 (N_9962,N_5541,N_1067);
and U9963 (N_9963,N_5588,N_4176);
and U9964 (N_9964,N_377,N_2650);
and U9965 (N_9965,N_1784,N_5742);
xnor U9966 (N_9966,N_4323,N_5265);
nand U9967 (N_9967,N_1069,N_403);
or U9968 (N_9968,N_4715,N_542);
or U9969 (N_9969,N_1100,N_2003);
and U9970 (N_9970,N_3480,N_926);
nand U9971 (N_9971,N_231,N_5912);
and U9972 (N_9972,N_3927,N_3072);
nand U9973 (N_9973,N_2413,N_1075);
nand U9974 (N_9974,N_5971,N_4303);
and U9975 (N_9975,N_315,N_1086);
xnor U9976 (N_9976,N_2079,N_5682);
or U9977 (N_9977,N_3444,N_2731);
xnor U9978 (N_9978,N_1485,N_1634);
nand U9979 (N_9979,N_128,N_402);
xnor U9980 (N_9980,N_2055,N_4740);
nand U9981 (N_9981,N_4590,N_1034);
and U9982 (N_9982,N_753,N_1630);
nor U9983 (N_9983,N_821,N_750);
nand U9984 (N_9984,N_3591,N_4940);
or U9985 (N_9985,N_5191,N_5510);
nor U9986 (N_9986,N_3967,N_39);
nand U9987 (N_9987,N_193,N_418);
and U9988 (N_9988,N_2601,N_4491);
nor U9989 (N_9989,N_5746,N_3320);
and U9990 (N_9990,N_3690,N_5695);
xnor U9991 (N_9991,N_5864,N_4168);
xnor U9992 (N_9992,N_3702,N_2463);
xor U9993 (N_9993,N_5384,N_4365);
nor U9994 (N_9994,N_2732,N_3024);
nand U9995 (N_9995,N_3913,N_941);
nor U9996 (N_9996,N_4709,N_459);
xnor U9997 (N_9997,N_4154,N_5789);
or U9998 (N_9998,N_2430,N_4091);
or U9999 (N_9999,N_4245,N_3310);
nand U10000 (N_10000,N_1397,N_3559);
nand U10001 (N_10001,N_3707,N_5518);
xor U10002 (N_10002,N_2198,N_2817);
and U10003 (N_10003,N_3711,N_3820);
or U10004 (N_10004,N_4212,N_1906);
nor U10005 (N_10005,N_3972,N_546);
nor U10006 (N_10006,N_2752,N_4928);
and U10007 (N_10007,N_2686,N_1037);
or U10008 (N_10008,N_4205,N_5493);
or U10009 (N_10009,N_3911,N_3940);
nand U10010 (N_10010,N_3246,N_5513);
and U10011 (N_10011,N_3778,N_1347);
or U10012 (N_10012,N_5109,N_4319);
nor U10013 (N_10013,N_83,N_3222);
xor U10014 (N_10014,N_1542,N_3048);
nand U10015 (N_10015,N_4289,N_1674);
or U10016 (N_10016,N_2863,N_2362);
or U10017 (N_10017,N_5265,N_5345);
nand U10018 (N_10018,N_318,N_737);
nand U10019 (N_10019,N_61,N_2268);
nand U10020 (N_10020,N_2919,N_3523);
nand U10021 (N_10021,N_3350,N_799);
nand U10022 (N_10022,N_1812,N_4356);
and U10023 (N_10023,N_815,N_4490);
nand U10024 (N_10024,N_5340,N_4136);
nor U10025 (N_10025,N_4310,N_1810);
xnor U10026 (N_10026,N_3553,N_4377);
nand U10027 (N_10027,N_4516,N_4144);
and U10028 (N_10028,N_1335,N_2521);
nand U10029 (N_10029,N_3062,N_4935);
and U10030 (N_10030,N_5174,N_3038);
and U10031 (N_10031,N_1713,N_1091);
nand U10032 (N_10032,N_1401,N_5705);
and U10033 (N_10033,N_431,N_2013);
and U10034 (N_10034,N_3425,N_5492);
xnor U10035 (N_10035,N_625,N_1315);
nand U10036 (N_10036,N_1058,N_4390);
xor U10037 (N_10037,N_4385,N_5109);
nand U10038 (N_10038,N_3213,N_1067);
and U10039 (N_10039,N_3591,N_4577);
and U10040 (N_10040,N_4628,N_3152);
nor U10041 (N_10041,N_4782,N_5646);
nor U10042 (N_10042,N_3472,N_1004);
and U10043 (N_10043,N_1446,N_5017);
xnor U10044 (N_10044,N_42,N_3776);
or U10045 (N_10045,N_5316,N_591);
or U10046 (N_10046,N_1923,N_4459);
nand U10047 (N_10047,N_3824,N_1640);
nand U10048 (N_10048,N_5651,N_1171);
nand U10049 (N_10049,N_1387,N_2093);
xor U10050 (N_10050,N_5097,N_4632);
nor U10051 (N_10051,N_5377,N_4987);
xor U10052 (N_10052,N_5371,N_3985);
nor U10053 (N_10053,N_1774,N_2442);
or U10054 (N_10054,N_1472,N_1078);
and U10055 (N_10055,N_2158,N_3597);
xor U10056 (N_10056,N_1357,N_206);
nand U10057 (N_10057,N_2922,N_3101);
nor U10058 (N_10058,N_5960,N_545);
or U10059 (N_10059,N_3297,N_2316);
xnor U10060 (N_10060,N_569,N_5470);
nor U10061 (N_10061,N_119,N_4942);
or U10062 (N_10062,N_3604,N_1694);
xnor U10063 (N_10063,N_481,N_4029);
nand U10064 (N_10064,N_1437,N_3826);
nand U10065 (N_10065,N_697,N_2520);
xor U10066 (N_10066,N_1963,N_3156);
and U10067 (N_10067,N_1927,N_777);
xor U10068 (N_10068,N_2990,N_5161);
nor U10069 (N_10069,N_4764,N_2362);
nand U10070 (N_10070,N_5468,N_90);
nor U10071 (N_10071,N_4650,N_2625);
xor U10072 (N_10072,N_735,N_5338);
and U10073 (N_10073,N_4016,N_1432);
nor U10074 (N_10074,N_5344,N_5267);
and U10075 (N_10075,N_1202,N_2773);
and U10076 (N_10076,N_3285,N_2448);
nor U10077 (N_10077,N_2667,N_1333);
or U10078 (N_10078,N_2450,N_5399);
nor U10079 (N_10079,N_2503,N_5965);
or U10080 (N_10080,N_5622,N_5594);
and U10081 (N_10081,N_3075,N_2759);
xnor U10082 (N_10082,N_1115,N_3807);
xnor U10083 (N_10083,N_407,N_3311);
nand U10084 (N_10084,N_5142,N_176);
xor U10085 (N_10085,N_83,N_215);
nor U10086 (N_10086,N_1620,N_5728);
nand U10087 (N_10087,N_2033,N_3268);
nor U10088 (N_10088,N_4118,N_5603);
nand U10089 (N_10089,N_5248,N_1947);
or U10090 (N_10090,N_3263,N_2689);
nand U10091 (N_10091,N_1039,N_2662);
nor U10092 (N_10092,N_3591,N_1604);
nand U10093 (N_10093,N_3244,N_4721);
and U10094 (N_10094,N_4768,N_5218);
xnor U10095 (N_10095,N_615,N_4188);
and U10096 (N_10096,N_3675,N_1695);
xnor U10097 (N_10097,N_436,N_578);
nand U10098 (N_10098,N_796,N_3860);
nor U10099 (N_10099,N_5670,N_550);
xor U10100 (N_10100,N_4266,N_4964);
and U10101 (N_10101,N_3779,N_2946);
or U10102 (N_10102,N_2830,N_5111);
nor U10103 (N_10103,N_1747,N_844);
and U10104 (N_10104,N_3717,N_1201);
nand U10105 (N_10105,N_5137,N_5587);
and U10106 (N_10106,N_1122,N_1024);
nand U10107 (N_10107,N_2806,N_4819);
or U10108 (N_10108,N_4022,N_2601);
and U10109 (N_10109,N_3106,N_1869);
xnor U10110 (N_10110,N_1277,N_1042);
and U10111 (N_10111,N_4212,N_1530);
and U10112 (N_10112,N_5842,N_246);
xor U10113 (N_10113,N_3670,N_887);
and U10114 (N_10114,N_1521,N_4867);
nand U10115 (N_10115,N_2805,N_5164);
nor U10116 (N_10116,N_5561,N_3989);
xnor U10117 (N_10117,N_4449,N_4171);
xor U10118 (N_10118,N_5636,N_5999);
nor U10119 (N_10119,N_5191,N_4885);
xnor U10120 (N_10120,N_3871,N_4163);
xor U10121 (N_10121,N_4959,N_1159);
xnor U10122 (N_10122,N_354,N_2466);
nor U10123 (N_10123,N_2691,N_215);
nand U10124 (N_10124,N_1866,N_5997);
xor U10125 (N_10125,N_5245,N_4299);
or U10126 (N_10126,N_1850,N_17);
nor U10127 (N_10127,N_4758,N_4181);
and U10128 (N_10128,N_484,N_10);
xnor U10129 (N_10129,N_679,N_434);
and U10130 (N_10130,N_533,N_23);
or U10131 (N_10131,N_5240,N_3410);
xor U10132 (N_10132,N_3893,N_2990);
nor U10133 (N_10133,N_3476,N_3268);
and U10134 (N_10134,N_3834,N_2737);
or U10135 (N_10135,N_4693,N_3099);
nand U10136 (N_10136,N_5329,N_4022);
and U10137 (N_10137,N_1182,N_635);
or U10138 (N_10138,N_1778,N_211);
or U10139 (N_10139,N_767,N_5961);
xor U10140 (N_10140,N_3193,N_5611);
xor U10141 (N_10141,N_4639,N_3261);
xnor U10142 (N_10142,N_5796,N_4698);
xnor U10143 (N_10143,N_474,N_4942);
or U10144 (N_10144,N_5668,N_4773);
and U10145 (N_10145,N_4358,N_359);
xor U10146 (N_10146,N_5013,N_2218);
xor U10147 (N_10147,N_5335,N_4093);
nand U10148 (N_10148,N_526,N_2801);
nor U10149 (N_10149,N_868,N_3012);
and U10150 (N_10150,N_1368,N_865);
or U10151 (N_10151,N_3437,N_4169);
nor U10152 (N_10152,N_3736,N_1429);
or U10153 (N_10153,N_4468,N_1363);
or U10154 (N_10154,N_3843,N_3513);
xor U10155 (N_10155,N_3741,N_4536);
nand U10156 (N_10156,N_1881,N_3803);
or U10157 (N_10157,N_560,N_2419);
or U10158 (N_10158,N_4083,N_2882);
nor U10159 (N_10159,N_1608,N_2663);
and U10160 (N_10160,N_4275,N_5083);
and U10161 (N_10161,N_5317,N_3634);
nand U10162 (N_10162,N_3950,N_5577);
and U10163 (N_10163,N_3041,N_3437);
nor U10164 (N_10164,N_4367,N_5408);
or U10165 (N_10165,N_3676,N_3261);
xnor U10166 (N_10166,N_3077,N_3428);
or U10167 (N_10167,N_4134,N_3975);
and U10168 (N_10168,N_2812,N_787);
and U10169 (N_10169,N_5255,N_4270);
nor U10170 (N_10170,N_730,N_4073);
nor U10171 (N_10171,N_100,N_1279);
nand U10172 (N_10172,N_3630,N_5060);
nand U10173 (N_10173,N_4971,N_381);
nor U10174 (N_10174,N_5317,N_4142);
or U10175 (N_10175,N_216,N_1660);
or U10176 (N_10176,N_624,N_555);
nand U10177 (N_10177,N_1948,N_50);
or U10178 (N_10178,N_462,N_1588);
or U10179 (N_10179,N_3395,N_261);
or U10180 (N_10180,N_4148,N_538);
xor U10181 (N_10181,N_3178,N_2708);
nor U10182 (N_10182,N_5314,N_4956);
nor U10183 (N_10183,N_3387,N_4752);
or U10184 (N_10184,N_3619,N_4160);
and U10185 (N_10185,N_5471,N_5461);
or U10186 (N_10186,N_5344,N_154);
or U10187 (N_10187,N_5600,N_616);
xnor U10188 (N_10188,N_925,N_2079);
nand U10189 (N_10189,N_347,N_1165);
and U10190 (N_10190,N_2252,N_608);
xor U10191 (N_10191,N_585,N_1478);
or U10192 (N_10192,N_3899,N_1542);
and U10193 (N_10193,N_421,N_5079);
and U10194 (N_10194,N_2749,N_5526);
or U10195 (N_10195,N_1089,N_38);
nor U10196 (N_10196,N_5012,N_3947);
nand U10197 (N_10197,N_2318,N_2130);
and U10198 (N_10198,N_3427,N_557);
or U10199 (N_10199,N_2367,N_3470);
nor U10200 (N_10200,N_4960,N_1889);
xnor U10201 (N_10201,N_5202,N_2262);
nor U10202 (N_10202,N_1889,N_4542);
or U10203 (N_10203,N_333,N_3357);
or U10204 (N_10204,N_4680,N_5659);
and U10205 (N_10205,N_2750,N_3044);
xor U10206 (N_10206,N_2264,N_60);
xor U10207 (N_10207,N_3834,N_644);
nor U10208 (N_10208,N_1291,N_5163);
nor U10209 (N_10209,N_3913,N_2288);
xor U10210 (N_10210,N_5276,N_1548);
nor U10211 (N_10211,N_3038,N_4841);
and U10212 (N_10212,N_2145,N_5007);
nand U10213 (N_10213,N_1665,N_5461);
nand U10214 (N_10214,N_2000,N_5713);
nor U10215 (N_10215,N_2348,N_5875);
or U10216 (N_10216,N_3027,N_4177);
and U10217 (N_10217,N_2103,N_455);
and U10218 (N_10218,N_2887,N_1690);
xnor U10219 (N_10219,N_921,N_437);
nand U10220 (N_10220,N_3057,N_602);
nor U10221 (N_10221,N_660,N_481);
xor U10222 (N_10222,N_4674,N_705);
xnor U10223 (N_10223,N_4069,N_2434);
xor U10224 (N_10224,N_1739,N_4100);
or U10225 (N_10225,N_4341,N_992);
or U10226 (N_10226,N_5735,N_180);
xnor U10227 (N_10227,N_2015,N_2520);
and U10228 (N_10228,N_4753,N_2867);
or U10229 (N_10229,N_2853,N_736);
xor U10230 (N_10230,N_1538,N_332);
nor U10231 (N_10231,N_1802,N_62);
or U10232 (N_10232,N_51,N_2834);
xnor U10233 (N_10233,N_5980,N_3843);
or U10234 (N_10234,N_4850,N_5032);
and U10235 (N_10235,N_1860,N_5123);
nor U10236 (N_10236,N_3119,N_5000);
xnor U10237 (N_10237,N_5649,N_4926);
and U10238 (N_10238,N_3504,N_5276);
or U10239 (N_10239,N_1646,N_940);
nand U10240 (N_10240,N_3287,N_2740);
and U10241 (N_10241,N_5188,N_2682);
nand U10242 (N_10242,N_4547,N_426);
or U10243 (N_10243,N_5867,N_2242);
nor U10244 (N_10244,N_5410,N_5521);
nand U10245 (N_10245,N_3776,N_3053);
and U10246 (N_10246,N_687,N_299);
and U10247 (N_10247,N_148,N_5060);
and U10248 (N_10248,N_5367,N_29);
or U10249 (N_10249,N_3740,N_2033);
nor U10250 (N_10250,N_5004,N_2094);
or U10251 (N_10251,N_783,N_5138);
nand U10252 (N_10252,N_1898,N_4678);
or U10253 (N_10253,N_2710,N_3584);
xor U10254 (N_10254,N_5386,N_1764);
and U10255 (N_10255,N_653,N_1196);
nand U10256 (N_10256,N_2427,N_4448);
xor U10257 (N_10257,N_5749,N_5306);
xnor U10258 (N_10258,N_1326,N_1617);
or U10259 (N_10259,N_216,N_1982);
nand U10260 (N_10260,N_1532,N_5410);
and U10261 (N_10261,N_4058,N_1066);
and U10262 (N_10262,N_879,N_2490);
or U10263 (N_10263,N_3515,N_521);
nor U10264 (N_10264,N_4186,N_1052);
nor U10265 (N_10265,N_753,N_1249);
and U10266 (N_10266,N_4703,N_912);
or U10267 (N_10267,N_397,N_5364);
and U10268 (N_10268,N_536,N_3074);
or U10269 (N_10269,N_1701,N_1774);
xnor U10270 (N_10270,N_2938,N_5814);
nor U10271 (N_10271,N_5520,N_2927);
nor U10272 (N_10272,N_708,N_1878);
and U10273 (N_10273,N_2980,N_5351);
xnor U10274 (N_10274,N_1349,N_3202);
nor U10275 (N_10275,N_5945,N_3572);
nand U10276 (N_10276,N_5962,N_3637);
nand U10277 (N_10277,N_1844,N_2703);
nand U10278 (N_10278,N_2741,N_1382);
or U10279 (N_10279,N_1861,N_3554);
or U10280 (N_10280,N_855,N_2156);
or U10281 (N_10281,N_660,N_2055);
xor U10282 (N_10282,N_2495,N_5083);
nor U10283 (N_10283,N_4277,N_100);
nor U10284 (N_10284,N_1707,N_5900);
and U10285 (N_10285,N_2571,N_242);
or U10286 (N_10286,N_2785,N_1279);
nand U10287 (N_10287,N_1527,N_1848);
and U10288 (N_10288,N_3415,N_1496);
and U10289 (N_10289,N_5643,N_5027);
nand U10290 (N_10290,N_2992,N_3054);
nand U10291 (N_10291,N_5240,N_92);
nand U10292 (N_10292,N_4239,N_5091);
or U10293 (N_10293,N_4337,N_5607);
nor U10294 (N_10294,N_2989,N_3011);
or U10295 (N_10295,N_1196,N_4029);
xor U10296 (N_10296,N_924,N_1204);
nand U10297 (N_10297,N_5643,N_5280);
nand U10298 (N_10298,N_3215,N_4912);
or U10299 (N_10299,N_2313,N_2979);
xnor U10300 (N_10300,N_2746,N_4090);
nor U10301 (N_10301,N_5575,N_1543);
nor U10302 (N_10302,N_5729,N_2449);
nand U10303 (N_10303,N_1098,N_4256);
and U10304 (N_10304,N_5656,N_2776);
nand U10305 (N_10305,N_3518,N_127);
nand U10306 (N_10306,N_3599,N_5887);
or U10307 (N_10307,N_3752,N_5399);
or U10308 (N_10308,N_4014,N_5903);
xnor U10309 (N_10309,N_4176,N_1775);
and U10310 (N_10310,N_2713,N_1845);
xnor U10311 (N_10311,N_1195,N_774);
nor U10312 (N_10312,N_785,N_3917);
xnor U10313 (N_10313,N_5717,N_531);
xor U10314 (N_10314,N_2370,N_2710);
nand U10315 (N_10315,N_795,N_1448);
and U10316 (N_10316,N_1972,N_2534);
xor U10317 (N_10317,N_5018,N_4815);
and U10318 (N_10318,N_1666,N_50);
and U10319 (N_10319,N_5192,N_4216);
nand U10320 (N_10320,N_5972,N_5246);
and U10321 (N_10321,N_5117,N_3332);
and U10322 (N_10322,N_4114,N_5219);
and U10323 (N_10323,N_5617,N_2978);
or U10324 (N_10324,N_4754,N_5009);
nand U10325 (N_10325,N_2725,N_3462);
or U10326 (N_10326,N_764,N_4553);
nand U10327 (N_10327,N_2478,N_603);
nand U10328 (N_10328,N_5610,N_1088);
xnor U10329 (N_10329,N_4950,N_567);
xnor U10330 (N_10330,N_3809,N_4763);
and U10331 (N_10331,N_5560,N_1924);
nand U10332 (N_10332,N_5036,N_841);
nor U10333 (N_10333,N_187,N_4214);
nand U10334 (N_10334,N_401,N_1564);
nor U10335 (N_10335,N_3674,N_1315);
xor U10336 (N_10336,N_5847,N_5158);
nor U10337 (N_10337,N_1091,N_717);
nand U10338 (N_10338,N_3296,N_3446);
nand U10339 (N_10339,N_1613,N_764);
nor U10340 (N_10340,N_1018,N_4098);
nand U10341 (N_10341,N_2386,N_3454);
or U10342 (N_10342,N_5329,N_2728);
nand U10343 (N_10343,N_5950,N_2168);
nand U10344 (N_10344,N_4297,N_964);
or U10345 (N_10345,N_4149,N_3751);
nor U10346 (N_10346,N_4464,N_5416);
nand U10347 (N_10347,N_800,N_240);
nand U10348 (N_10348,N_5125,N_5636);
nor U10349 (N_10349,N_2689,N_4421);
nor U10350 (N_10350,N_1580,N_1707);
or U10351 (N_10351,N_2077,N_3455);
and U10352 (N_10352,N_2950,N_5622);
nor U10353 (N_10353,N_1115,N_5953);
nand U10354 (N_10354,N_5053,N_4671);
nand U10355 (N_10355,N_3560,N_3038);
and U10356 (N_10356,N_5585,N_2886);
nor U10357 (N_10357,N_3236,N_285);
nor U10358 (N_10358,N_5516,N_4653);
xor U10359 (N_10359,N_5338,N_1558);
nor U10360 (N_10360,N_3911,N_91);
and U10361 (N_10361,N_5223,N_3505);
nor U10362 (N_10362,N_2191,N_5653);
xor U10363 (N_10363,N_3274,N_5198);
or U10364 (N_10364,N_5374,N_4981);
nor U10365 (N_10365,N_1793,N_5968);
nor U10366 (N_10366,N_4504,N_3776);
or U10367 (N_10367,N_3541,N_3972);
xor U10368 (N_10368,N_2482,N_3552);
nand U10369 (N_10369,N_5801,N_4243);
or U10370 (N_10370,N_1907,N_4331);
nand U10371 (N_10371,N_2453,N_2617);
xor U10372 (N_10372,N_5932,N_709);
and U10373 (N_10373,N_5058,N_2402);
and U10374 (N_10374,N_1643,N_2346);
nand U10375 (N_10375,N_1487,N_1965);
xor U10376 (N_10376,N_4973,N_988);
or U10377 (N_10377,N_683,N_1747);
nand U10378 (N_10378,N_2683,N_4083);
xnor U10379 (N_10379,N_1942,N_4057);
nand U10380 (N_10380,N_1357,N_1621);
and U10381 (N_10381,N_3789,N_3798);
nor U10382 (N_10382,N_4323,N_3560);
or U10383 (N_10383,N_5853,N_4590);
nor U10384 (N_10384,N_2245,N_1355);
nand U10385 (N_10385,N_5855,N_5135);
xor U10386 (N_10386,N_5003,N_4021);
and U10387 (N_10387,N_1033,N_2036);
or U10388 (N_10388,N_2338,N_3365);
or U10389 (N_10389,N_2223,N_3407);
xnor U10390 (N_10390,N_1758,N_3297);
or U10391 (N_10391,N_2624,N_5716);
nor U10392 (N_10392,N_2852,N_5944);
or U10393 (N_10393,N_4153,N_4477);
or U10394 (N_10394,N_372,N_2836);
and U10395 (N_10395,N_5811,N_21);
nor U10396 (N_10396,N_2546,N_2295);
and U10397 (N_10397,N_4151,N_5285);
or U10398 (N_10398,N_5702,N_5761);
nor U10399 (N_10399,N_3189,N_1815);
nand U10400 (N_10400,N_330,N_3002);
xnor U10401 (N_10401,N_4295,N_4867);
nand U10402 (N_10402,N_122,N_1241);
nand U10403 (N_10403,N_1700,N_2851);
nor U10404 (N_10404,N_5624,N_5147);
nor U10405 (N_10405,N_1126,N_1995);
or U10406 (N_10406,N_895,N_3056);
nor U10407 (N_10407,N_2602,N_3494);
and U10408 (N_10408,N_4622,N_204);
nor U10409 (N_10409,N_5232,N_4065);
nand U10410 (N_10410,N_1703,N_3601);
nand U10411 (N_10411,N_2344,N_5543);
nor U10412 (N_10412,N_4823,N_4579);
nand U10413 (N_10413,N_4524,N_4464);
or U10414 (N_10414,N_1918,N_4284);
nor U10415 (N_10415,N_4597,N_114);
nand U10416 (N_10416,N_2306,N_5081);
nand U10417 (N_10417,N_3943,N_3622);
or U10418 (N_10418,N_588,N_5448);
xor U10419 (N_10419,N_4315,N_5175);
or U10420 (N_10420,N_3698,N_3601);
xor U10421 (N_10421,N_577,N_3556);
nand U10422 (N_10422,N_2380,N_596);
and U10423 (N_10423,N_1049,N_1684);
nand U10424 (N_10424,N_4570,N_738);
and U10425 (N_10425,N_4197,N_2277);
and U10426 (N_10426,N_5385,N_5693);
nor U10427 (N_10427,N_3333,N_4125);
nor U10428 (N_10428,N_4342,N_4984);
and U10429 (N_10429,N_1975,N_4852);
nor U10430 (N_10430,N_4048,N_420);
and U10431 (N_10431,N_2217,N_815);
nand U10432 (N_10432,N_3205,N_1262);
or U10433 (N_10433,N_3063,N_1225);
xor U10434 (N_10434,N_991,N_3186);
or U10435 (N_10435,N_1994,N_1068);
or U10436 (N_10436,N_5319,N_4096);
or U10437 (N_10437,N_5732,N_4186);
nand U10438 (N_10438,N_5872,N_490);
xor U10439 (N_10439,N_4910,N_197);
or U10440 (N_10440,N_997,N_1819);
nor U10441 (N_10441,N_5722,N_1747);
nor U10442 (N_10442,N_877,N_5570);
nand U10443 (N_10443,N_3367,N_3604);
xnor U10444 (N_10444,N_4450,N_3750);
xnor U10445 (N_10445,N_1895,N_3684);
nor U10446 (N_10446,N_4494,N_5567);
or U10447 (N_10447,N_1551,N_4243);
xnor U10448 (N_10448,N_2260,N_5187);
nand U10449 (N_10449,N_589,N_4229);
and U10450 (N_10450,N_4242,N_1254);
or U10451 (N_10451,N_5154,N_2242);
nand U10452 (N_10452,N_1197,N_1070);
or U10453 (N_10453,N_4375,N_521);
xor U10454 (N_10454,N_2664,N_2812);
or U10455 (N_10455,N_789,N_1651);
nor U10456 (N_10456,N_788,N_4986);
nand U10457 (N_10457,N_122,N_5697);
nand U10458 (N_10458,N_5840,N_4244);
xor U10459 (N_10459,N_1458,N_4236);
nand U10460 (N_10460,N_2036,N_5147);
xor U10461 (N_10461,N_2620,N_4217);
or U10462 (N_10462,N_3830,N_5626);
nor U10463 (N_10463,N_2146,N_2116);
nand U10464 (N_10464,N_4844,N_4638);
or U10465 (N_10465,N_3733,N_748);
and U10466 (N_10466,N_2159,N_1163);
nor U10467 (N_10467,N_5189,N_3299);
and U10468 (N_10468,N_5947,N_5525);
and U10469 (N_10469,N_3619,N_5377);
and U10470 (N_10470,N_1609,N_5205);
nor U10471 (N_10471,N_5268,N_5719);
xor U10472 (N_10472,N_4901,N_1843);
nand U10473 (N_10473,N_3729,N_172);
nor U10474 (N_10474,N_175,N_2795);
and U10475 (N_10475,N_5722,N_4224);
xor U10476 (N_10476,N_4195,N_5510);
xnor U10477 (N_10477,N_5511,N_310);
xnor U10478 (N_10478,N_2817,N_5056);
and U10479 (N_10479,N_374,N_1778);
and U10480 (N_10480,N_311,N_5376);
and U10481 (N_10481,N_5336,N_5901);
nand U10482 (N_10482,N_2882,N_1969);
or U10483 (N_10483,N_5491,N_2100);
xnor U10484 (N_10484,N_2365,N_1637);
nor U10485 (N_10485,N_1051,N_2334);
xnor U10486 (N_10486,N_91,N_5008);
nand U10487 (N_10487,N_1466,N_4528);
and U10488 (N_10488,N_878,N_5213);
xnor U10489 (N_10489,N_1188,N_5249);
nor U10490 (N_10490,N_1264,N_1522);
or U10491 (N_10491,N_842,N_4051);
nor U10492 (N_10492,N_1295,N_668);
nand U10493 (N_10493,N_2707,N_690);
nand U10494 (N_10494,N_4283,N_3113);
xnor U10495 (N_10495,N_4136,N_2341);
or U10496 (N_10496,N_1505,N_5109);
or U10497 (N_10497,N_2429,N_309);
and U10498 (N_10498,N_2408,N_2800);
nand U10499 (N_10499,N_4327,N_2243);
xnor U10500 (N_10500,N_405,N_5208);
nor U10501 (N_10501,N_5500,N_5006);
or U10502 (N_10502,N_1399,N_670);
and U10503 (N_10503,N_1459,N_4978);
or U10504 (N_10504,N_2828,N_2426);
nand U10505 (N_10505,N_2497,N_4075);
xor U10506 (N_10506,N_995,N_1266);
nand U10507 (N_10507,N_4374,N_1552);
or U10508 (N_10508,N_891,N_1878);
and U10509 (N_10509,N_2899,N_3078);
nor U10510 (N_10510,N_3948,N_2168);
nand U10511 (N_10511,N_5515,N_292);
or U10512 (N_10512,N_3410,N_427);
nand U10513 (N_10513,N_5221,N_4807);
and U10514 (N_10514,N_2292,N_5869);
and U10515 (N_10515,N_943,N_2328);
nor U10516 (N_10516,N_3433,N_699);
nand U10517 (N_10517,N_2593,N_3084);
nand U10518 (N_10518,N_2113,N_4393);
nand U10519 (N_10519,N_1186,N_3059);
nor U10520 (N_10520,N_74,N_5048);
nand U10521 (N_10521,N_3534,N_7);
and U10522 (N_10522,N_2219,N_4192);
nor U10523 (N_10523,N_1289,N_171);
and U10524 (N_10524,N_2290,N_1955);
xnor U10525 (N_10525,N_3215,N_3807);
xor U10526 (N_10526,N_5177,N_1705);
xnor U10527 (N_10527,N_5666,N_2812);
and U10528 (N_10528,N_4540,N_326);
nand U10529 (N_10529,N_2138,N_4094);
and U10530 (N_10530,N_1496,N_1533);
nand U10531 (N_10531,N_2908,N_5844);
nand U10532 (N_10532,N_1968,N_178);
and U10533 (N_10533,N_869,N_1863);
and U10534 (N_10534,N_3969,N_1461);
or U10535 (N_10535,N_2833,N_3799);
and U10536 (N_10536,N_5058,N_5955);
xnor U10537 (N_10537,N_5208,N_2455);
xor U10538 (N_10538,N_5816,N_408);
xor U10539 (N_10539,N_3183,N_4180);
nor U10540 (N_10540,N_828,N_2080);
xnor U10541 (N_10541,N_740,N_5419);
xor U10542 (N_10542,N_1331,N_2140);
and U10543 (N_10543,N_2106,N_5719);
nand U10544 (N_10544,N_3599,N_3379);
xor U10545 (N_10545,N_1255,N_355);
nand U10546 (N_10546,N_4820,N_1312);
or U10547 (N_10547,N_5166,N_2447);
or U10548 (N_10548,N_2741,N_590);
nor U10549 (N_10549,N_4718,N_2255);
and U10550 (N_10550,N_759,N_4093);
xor U10551 (N_10551,N_2272,N_4538);
xor U10552 (N_10552,N_5459,N_5178);
or U10553 (N_10553,N_648,N_5852);
nand U10554 (N_10554,N_1522,N_5706);
nand U10555 (N_10555,N_1595,N_139);
nand U10556 (N_10556,N_3179,N_3976);
and U10557 (N_10557,N_2118,N_807);
and U10558 (N_10558,N_4475,N_222);
or U10559 (N_10559,N_3877,N_4887);
nand U10560 (N_10560,N_5619,N_2848);
nor U10561 (N_10561,N_5503,N_2069);
xnor U10562 (N_10562,N_1372,N_5911);
or U10563 (N_10563,N_496,N_91);
and U10564 (N_10564,N_5579,N_2070);
or U10565 (N_10565,N_4867,N_2766);
xnor U10566 (N_10566,N_1621,N_1576);
xor U10567 (N_10567,N_5033,N_4389);
and U10568 (N_10568,N_4556,N_4299);
nor U10569 (N_10569,N_2194,N_8);
and U10570 (N_10570,N_582,N_5821);
nor U10571 (N_10571,N_1712,N_3270);
and U10572 (N_10572,N_3706,N_1766);
or U10573 (N_10573,N_2770,N_1450);
nor U10574 (N_10574,N_5931,N_19);
nor U10575 (N_10575,N_979,N_2136);
nor U10576 (N_10576,N_3480,N_145);
or U10577 (N_10577,N_3110,N_20);
nor U10578 (N_10578,N_3081,N_1662);
nand U10579 (N_10579,N_3400,N_691);
or U10580 (N_10580,N_564,N_3787);
and U10581 (N_10581,N_1858,N_2634);
xnor U10582 (N_10582,N_4135,N_4152);
and U10583 (N_10583,N_4914,N_2271);
nand U10584 (N_10584,N_1240,N_5656);
xor U10585 (N_10585,N_2327,N_5616);
or U10586 (N_10586,N_1602,N_2424);
nand U10587 (N_10587,N_5113,N_2043);
and U10588 (N_10588,N_4919,N_3173);
and U10589 (N_10589,N_3573,N_2665);
xnor U10590 (N_10590,N_5617,N_5212);
and U10591 (N_10591,N_3619,N_1034);
or U10592 (N_10592,N_5216,N_5853);
xnor U10593 (N_10593,N_2335,N_4868);
xnor U10594 (N_10594,N_2173,N_3575);
or U10595 (N_10595,N_2726,N_948);
nor U10596 (N_10596,N_5431,N_5048);
nand U10597 (N_10597,N_1128,N_3319);
nor U10598 (N_10598,N_3230,N_1338);
or U10599 (N_10599,N_612,N_231);
nand U10600 (N_10600,N_2027,N_2107);
nor U10601 (N_10601,N_4897,N_5512);
or U10602 (N_10602,N_5542,N_2195);
or U10603 (N_10603,N_1077,N_4518);
nand U10604 (N_10604,N_3007,N_1220);
and U10605 (N_10605,N_5415,N_3190);
xnor U10606 (N_10606,N_1250,N_5230);
nand U10607 (N_10607,N_1593,N_3818);
and U10608 (N_10608,N_1899,N_5256);
or U10609 (N_10609,N_4191,N_4852);
and U10610 (N_10610,N_58,N_205);
nand U10611 (N_10611,N_5021,N_5831);
nand U10612 (N_10612,N_1576,N_3209);
nand U10613 (N_10613,N_3398,N_5269);
or U10614 (N_10614,N_261,N_2987);
nand U10615 (N_10615,N_798,N_4531);
and U10616 (N_10616,N_1980,N_5366);
or U10617 (N_10617,N_5807,N_3992);
xnor U10618 (N_10618,N_5124,N_4598);
or U10619 (N_10619,N_5787,N_555);
or U10620 (N_10620,N_2165,N_1073);
and U10621 (N_10621,N_5292,N_3613);
and U10622 (N_10622,N_693,N_754);
xnor U10623 (N_10623,N_749,N_40);
and U10624 (N_10624,N_859,N_2904);
and U10625 (N_10625,N_3852,N_4716);
xor U10626 (N_10626,N_462,N_5268);
nor U10627 (N_10627,N_2555,N_3595);
nor U10628 (N_10628,N_1592,N_3786);
nand U10629 (N_10629,N_4133,N_2740);
and U10630 (N_10630,N_3419,N_3145);
xor U10631 (N_10631,N_3286,N_2968);
and U10632 (N_10632,N_2176,N_581);
or U10633 (N_10633,N_1405,N_4852);
xor U10634 (N_10634,N_5113,N_2601);
or U10635 (N_10635,N_3397,N_1679);
and U10636 (N_10636,N_5047,N_1113);
nor U10637 (N_10637,N_2348,N_2067);
xnor U10638 (N_10638,N_2642,N_4162);
nand U10639 (N_10639,N_228,N_4588);
xnor U10640 (N_10640,N_4801,N_197);
nand U10641 (N_10641,N_4348,N_1234);
xor U10642 (N_10642,N_4565,N_3838);
and U10643 (N_10643,N_3151,N_4608);
xnor U10644 (N_10644,N_2454,N_5981);
and U10645 (N_10645,N_3927,N_4263);
or U10646 (N_10646,N_3470,N_1631);
and U10647 (N_10647,N_1664,N_3983);
nor U10648 (N_10648,N_2190,N_4086);
nand U10649 (N_10649,N_2283,N_5933);
xor U10650 (N_10650,N_4925,N_4789);
and U10651 (N_10651,N_1556,N_5216);
nor U10652 (N_10652,N_2381,N_5076);
and U10653 (N_10653,N_3591,N_3434);
xor U10654 (N_10654,N_738,N_1929);
nor U10655 (N_10655,N_3852,N_4381);
and U10656 (N_10656,N_3258,N_3310);
nand U10657 (N_10657,N_4164,N_5411);
or U10658 (N_10658,N_2978,N_4588);
and U10659 (N_10659,N_5396,N_3718);
or U10660 (N_10660,N_1676,N_4079);
and U10661 (N_10661,N_4476,N_525);
nor U10662 (N_10662,N_1413,N_2877);
xor U10663 (N_10663,N_1324,N_3803);
nand U10664 (N_10664,N_1470,N_2239);
and U10665 (N_10665,N_5295,N_2404);
and U10666 (N_10666,N_3682,N_5615);
nand U10667 (N_10667,N_5320,N_4502);
nor U10668 (N_10668,N_4279,N_970);
nand U10669 (N_10669,N_4602,N_234);
nor U10670 (N_10670,N_4098,N_4858);
xnor U10671 (N_10671,N_3834,N_5163);
or U10672 (N_10672,N_3750,N_3741);
or U10673 (N_10673,N_2743,N_2054);
xnor U10674 (N_10674,N_5827,N_5791);
nor U10675 (N_10675,N_1033,N_1807);
nor U10676 (N_10676,N_5983,N_3333);
nor U10677 (N_10677,N_1808,N_5954);
xor U10678 (N_10678,N_5927,N_304);
nor U10679 (N_10679,N_3812,N_3206);
or U10680 (N_10680,N_18,N_4484);
nand U10681 (N_10681,N_5905,N_3830);
nand U10682 (N_10682,N_3495,N_1669);
and U10683 (N_10683,N_4224,N_4660);
xor U10684 (N_10684,N_1784,N_1207);
nand U10685 (N_10685,N_4070,N_675);
and U10686 (N_10686,N_1464,N_3408);
or U10687 (N_10687,N_1507,N_3922);
and U10688 (N_10688,N_895,N_5996);
nor U10689 (N_10689,N_1865,N_4401);
nand U10690 (N_10690,N_4485,N_5573);
or U10691 (N_10691,N_5139,N_5161);
and U10692 (N_10692,N_5340,N_2913);
xor U10693 (N_10693,N_352,N_4202);
or U10694 (N_10694,N_2460,N_4113);
nand U10695 (N_10695,N_3913,N_1628);
nand U10696 (N_10696,N_3219,N_2002);
nor U10697 (N_10697,N_3159,N_3242);
and U10698 (N_10698,N_3370,N_1218);
or U10699 (N_10699,N_5858,N_4259);
or U10700 (N_10700,N_3847,N_1272);
and U10701 (N_10701,N_3433,N_692);
or U10702 (N_10702,N_3670,N_820);
nand U10703 (N_10703,N_1998,N_4568);
and U10704 (N_10704,N_4092,N_2228);
or U10705 (N_10705,N_3011,N_4351);
nor U10706 (N_10706,N_173,N_2816);
nor U10707 (N_10707,N_1171,N_1530);
nor U10708 (N_10708,N_3999,N_3844);
and U10709 (N_10709,N_3305,N_1750);
and U10710 (N_10710,N_2747,N_3422);
or U10711 (N_10711,N_3899,N_5999);
xnor U10712 (N_10712,N_3204,N_5879);
xor U10713 (N_10713,N_5684,N_2275);
and U10714 (N_10714,N_669,N_2171);
and U10715 (N_10715,N_5661,N_4705);
nand U10716 (N_10716,N_1434,N_351);
or U10717 (N_10717,N_3201,N_5509);
or U10718 (N_10718,N_4982,N_5622);
nand U10719 (N_10719,N_1744,N_3174);
nor U10720 (N_10720,N_3639,N_3451);
or U10721 (N_10721,N_1012,N_504);
and U10722 (N_10722,N_542,N_5394);
and U10723 (N_10723,N_4621,N_4660);
nor U10724 (N_10724,N_4426,N_2640);
nand U10725 (N_10725,N_1465,N_2955);
and U10726 (N_10726,N_5787,N_4000);
xor U10727 (N_10727,N_1719,N_5930);
xnor U10728 (N_10728,N_4944,N_5706);
xor U10729 (N_10729,N_3003,N_4282);
nand U10730 (N_10730,N_2618,N_355);
and U10731 (N_10731,N_4749,N_1062);
nor U10732 (N_10732,N_4162,N_4789);
xnor U10733 (N_10733,N_637,N_3691);
xnor U10734 (N_10734,N_4596,N_152);
xnor U10735 (N_10735,N_4418,N_5693);
and U10736 (N_10736,N_5972,N_4700);
nor U10737 (N_10737,N_4679,N_4151);
or U10738 (N_10738,N_4974,N_3463);
xnor U10739 (N_10739,N_4871,N_75);
nor U10740 (N_10740,N_96,N_3585);
and U10741 (N_10741,N_4235,N_5224);
nor U10742 (N_10742,N_5159,N_4356);
xnor U10743 (N_10743,N_5292,N_3548);
nand U10744 (N_10744,N_3879,N_5922);
nor U10745 (N_10745,N_4167,N_2664);
nand U10746 (N_10746,N_1503,N_3988);
nor U10747 (N_10747,N_445,N_1071);
and U10748 (N_10748,N_4356,N_2634);
and U10749 (N_10749,N_4451,N_427);
and U10750 (N_10750,N_3675,N_2029);
or U10751 (N_10751,N_3941,N_2385);
xnor U10752 (N_10752,N_3637,N_2509);
or U10753 (N_10753,N_1489,N_892);
and U10754 (N_10754,N_2203,N_5712);
xor U10755 (N_10755,N_736,N_1050);
or U10756 (N_10756,N_4091,N_3255);
nand U10757 (N_10757,N_2598,N_113);
and U10758 (N_10758,N_2212,N_3176);
nand U10759 (N_10759,N_5227,N_4983);
xnor U10760 (N_10760,N_5194,N_814);
xnor U10761 (N_10761,N_4808,N_5211);
xnor U10762 (N_10762,N_2215,N_3421);
xor U10763 (N_10763,N_5473,N_5458);
or U10764 (N_10764,N_2482,N_3846);
and U10765 (N_10765,N_3208,N_3881);
nand U10766 (N_10766,N_2626,N_2961);
or U10767 (N_10767,N_4359,N_2939);
or U10768 (N_10768,N_3111,N_404);
and U10769 (N_10769,N_1985,N_489);
nor U10770 (N_10770,N_1181,N_3570);
and U10771 (N_10771,N_3231,N_5411);
nand U10772 (N_10772,N_5246,N_3996);
xnor U10773 (N_10773,N_3660,N_2405);
nor U10774 (N_10774,N_5741,N_2417);
or U10775 (N_10775,N_3389,N_5139);
xor U10776 (N_10776,N_99,N_5492);
and U10777 (N_10777,N_1209,N_3654);
and U10778 (N_10778,N_1162,N_2378);
xnor U10779 (N_10779,N_1759,N_4258);
xor U10780 (N_10780,N_5499,N_3704);
nand U10781 (N_10781,N_5159,N_5082);
or U10782 (N_10782,N_2323,N_5808);
nor U10783 (N_10783,N_2536,N_3088);
nand U10784 (N_10784,N_4816,N_2645);
and U10785 (N_10785,N_4297,N_5502);
xnor U10786 (N_10786,N_4175,N_4962);
and U10787 (N_10787,N_1451,N_5642);
nand U10788 (N_10788,N_738,N_3107);
or U10789 (N_10789,N_5087,N_3514);
and U10790 (N_10790,N_4661,N_3799);
or U10791 (N_10791,N_734,N_2492);
nand U10792 (N_10792,N_2604,N_5153);
or U10793 (N_10793,N_793,N_379);
nor U10794 (N_10794,N_129,N_4964);
or U10795 (N_10795,N_5233,N_1657);
and U10796 (N_10796,N_65,N_5390);
or U10797 (N_10797,N_1135,N_4267);
xnor U10798 (N_10798,N_2905,N_58);
or U10799 (N_10799,N_3594,N_2498);
xor U10800 (N_10800,N_2624,N_741);
or U10801 (N_10801,N_25,N_2710);
or U10802 (N_10802,N_2154,N_5272);
or U10803 (N_10803,N_5399,N_556);
or U10804 (N_10804,N_3539,N_5784);
and U10805 (N_10805,N_5495,N_320);
or U10806 (N_10806,N_3367,N_2540);
or U10807 (N_10807,N_527,N_4341);
or U10808 (N_10808,N_172,N_5940);
nand U10809 (N_10809,N_4647,N_5484);
or U10810 (N_10810,N_5926,N_2625);
xnor U10811 (N_10811,N_5629,N_4016);
nand U10812 (N_10812,N_2891,N_3780);
xnor U10813 (N_10813,N_3760,N_1912);
and U10814 (N_10814,N_640,N_5907);
nor U10815 (N_10815,N_5238,N_3836);
and U10816 (N_10816,N_4796,N_4226);
xnor U10817 (N_10817,N_2221,N_1150);
nand U10818 (N_10818,N_1128,N_4921);
xor U10819 (N_10819,N_3002,N_183);
or U10820 (N_10820,N_1480,N_2329);
xor U10821 (N_10821,N_1771,N_888);
and U10822 (N_10822,N_4379,N_3577);
nand U10823 (N_10823,N_5117,N_2270);
or U10824 (N_10824,N_3050,N_1312);
xor U10825 (N_10825,N_1250,N_4712);
nand U10826 (N_10826,N_3783,N_5888);
and U10827 (N_10827,N_2502,N_5031);
xnor U10828 (N_10828,N_5452,N_343);
nor U10829 (N_10829,N_3303,N_5815);
nor U10830 (N_10830,N_4016,N_1305);
nor U10831 (N_10831,N_753,N_2936);
nor U10832 (N_10832,N_4135,N_4587);
or U10833 (N_10833,N_4854,N_1827);
or U10834 (N_10834,N_5681,N_4985);
nor U10835 (N_10835,N_2001,N_4246);
and U10836 (N_10836,N_2122,N_2433);
nor U10837 (N_10837,N_5348,N_784);
or U10838 (N_10838,N_5238,N_5443);
xor U10839 (N_10839,N_5220,N_4135);
or U10840 (N_10840,N_2598,N_1608);
and U10841 (N_10841,N_2620,N_579);
nor U10842 (N_10842,N_673,N_3274);
nor U10843 (N_10843,N_3145,N_3197);
nand U10844 (N_10844,N_5529,N_3859);
nand U10845 (N_10845,N_2029,N_5693);
nand U10846 (N_10846,N_1625,N_3152);
xor U10847 (N_10847,N_3263,N_688);
nand U10848 (N_10848,N_2436,N_2734);
nor U10849 (N_10849,N_4593,N_1827);
xor U10850 (N_10850,N_3740,N_5936);
or U10851 (N_10851,N_3274,N_493);
and U10852 (N_10852,N_5951,N_5360);
xor U10853 (N_10853,N_5985,N_2038);
nor U10854 (N_10854,N_2455,N_1997);
or U10855 (N_10855,N_4011,N_4205);
nor U10856 (N_10856,N_5745,N_2542);
or U10857 (N_10857,N_2136,N_1018);
nor U10858 (N_10858,N_3915,N_5590);
nor U10859 (N_10859,N_1066,N_2031);
and U10860 (N_10860,N_4328,N_766);
nand U10861 (N_10861,N_4983,N_4435);
nand U10862 (N_10862,N_427,N_4083);
or U10863 (N_10863,N_267,N_3064);
or U10864 (N_10864,N_2739,N_4560);
nor U10865 (N_10865,N_5220,N_3041);
and U10866 (N_10866,N_2991,N_1282);
xor U10867 (N_10867,N_1149,N_924);
nor U10868 (N_10868,N_3353,N_1314);
or U10869 (N_10869,N_2592,N_2857);
or U10870 (N_10870,N_2147,N_888);
nor U10871 (N_10871,N_4350,N_3628);
and U10872 (N_10872,N_5608,N_4878);
or U10873 (N_10873,N_3810,N_636);
and U10874 (N_10874,N_5724,N_2137);
nor U10875 (N_10875,N_4754,N_2948);
nor U10876 (N_10876,N_1565,N_255);
nand U10877 (N_10877,N_3981,N_4762);
or U10878 (N_10878,N_5213,N_379);
and U10879 (N_10879,N_2615,N_1286);
xnor U10880 (N_10880,N_5276,N_1371);
nor U10881 (N_10881,N_983,N_1707);
xor U10882 (N_10882,N_344,N_1613);
xor U10883 (N_10883,N_3720,N_4061);
nor U10884 (N_10884,N_5816,N_2409);
nor U10885 (N_10885,N_4952,N_4099);
nor U10886 (N_10886,N_2721,N_5022);
nor U10887 (N_10887,N_1730,N_372);
xnor U10888 (N_10888,N_1854,N_2426);
xnor U10889 (N_10889,N_3523,N_5113);
nand U10890 (N_10890,N_2917,N_1235);
nor U10891 (N_10891,N_1205,N_4418);
nor U10892 (N_10892,N_1643,N_3732);
or U10893 (N_10893,N_2679,N_569);
nor U10894 (N_10894,N_4965,N_2914);
and U10895 (N_10895,N_3502,N_4141);
and U10896 (N_10896,N_5018,N_374);
or U10897 (N_10897,N_2889,N_1940);
and U10898 (N_10898,N_725,N_5145);
xor U10899 (N_10899,N_994,N_4739);
and U10900 (N_10900,N_1662,N_1511);
nand U10901 (N_10901,N_1233,N_5270);
or U10902 (N_10902,N_4396,N_1917);
nand U10903 (N_10903,N_1500,N_5125);
nor U10904 (N_10904,N_2422,N_5829);
nand U10905 (N_10905,N_2882,N_2382);
nor U10906 (N_10906,N_1632,N_3001);
nor U10907 (N_10907,N_956,N_1282);
or U10908 (N_10908,N_5241,N_1687);
nor U10909 (N_10909,N_1411,N_1978);
and U10910 (N_10910,N_4287,N_2198);
nand U10911 (N_10911,N_2569,N_158);
nor U10912 (N_10912,N_3658,N_5328);
or U10913 (N_10913,N_1204,N_3493);
nor U10914 (N_10914,N_5491,N_5552);
nand U10915 (N_10915,N_337,N_1167);
nor U10916 (N_10916,N_4906,N_3219);
and U10917 (N_10917,N_5433,N_4620);
xnor U10918 (N_10918,N_4067,N_788);
nor U10919 (N_10919,N_1248,N_1148);
nor U10920 (N_10920,N_2954,N_5640);
xor U10921 (N_10921,N_4145,N_3026);
nand U10922 (N_10922,N_1029,N_4461);
nor U10923 (N_10923,N_4422,N_1251);
nor U10924 (N_10924,N_3249,N_5237);
or U10925 (N_10925,N_2747,N_3489);
nor U10926 (N_10926,N_5244,N_747);
xnor U10927 (N_10927,N_2586,N_4394);
or U10928 (N_10928,N_623,N_2105);
or U10929 (N_10929,N_1468,N_242);
or U10930 (N_10930,N_2361,N_3064);
xnor U10931 (N_10931,N_5524,N_1761);
nand U10932 (N_10932,N_385,N_4870);
or U10933 (N_10933,N_1449,N_2023);
xor U10934 (N_10934,N_2111,N_5023);
nand U10935 (N_10935,N_1456,N_4174);
xor U10936 (N_10936,N_3928,N_4712);
nor U10937 (N_10937,N_2559,N_1047);
or U10938 (N_10938,N_2189,N_1214);
and U10939 (N_10939,N_5559,N_5686);
nor U10940 (N_10940,N_5805,N_984);
or U10941 (N_10941,N_4004,N_1258);
nor U10942 (N_10942,N_4747,N_440);
nor U10943 (N_10943,N_648,N_795);
xnor U10944 (N_10944,N_3192,N_2670);
nand U10945 (N_10945,N_536,N_202);
or U10946 (N_10946,N_3154,N_5450);
xnor U10947 (N_10947,N_5559,N_4020);
nand U10948 (N_10948,N_999,N_1241);
nor U10949 (N_10949,N_421,N_916);
nor U10950 (N_10950,N_1049,N_1188);
and U10951 (N_10951,N_4156,N_4176);
and U10952 (N_10952,N_5158,N_5273);
nand U10953 (N_10953,N_1561,N_5980);
nand U10954 (N_10954,N_2959,N_5763);
nand U10955 (N_10955,N_4259,N_1877);
nor U10956 (N_10956,N_5532,N_4116);
and U10957 (N_10957,N_2865,N_3583);
xnor U10958 (N_10958,N_4959,N_5522);
or U10959 (N_10959,N_3867,N_2051);
nor U10960 (N_10960,N_4287,N_1727);
xnor U10961 (N_10961,N_846,N_2270);
or U10962 (N_10962,N_3536,N_3545);
or U10963 (N_10963,N_685,N_914);
and U10964 (N_10964,N_4261,N_1817);
nor U10965 (N_10965,N_3768,N_4361);
nor U10966 (N_10966,N_3480,N_877);
and U10967 (N_10967,N_3034,N_1440);
nor U10968 (N_10968,N_501,N_646);
xor U10969 (N_10969,N_1626,N_5569);
or U10970 (N_10970,N_5843,N_3264);
nor U10971 (N_10971,N_4268,N_4921);
and U10972 (N_10972,N_2389,N_2615);
nor U10973 (N_10973,N_3227,N_2569);
nand U10974 (N_10974,N_5864,N_2987);
nand U10975 (N_10975,N_4729,N_2095);
and U10976 (N_10976,N_170,N_2457);
nand U10977 (N_10977,N_497,N_4976);
xnor U10978 (N_10978,N_3153,N_4561);
nor U10979 (N_10979,N_3684,N_1304);
nand U10980 (N_10980,N_4949,N_3123);
nand U10981 (N_10981,N_3620,N_3589);
nor U10982 (N_10982,N_5686,N_896);
nand U10983 (N_10983,N_2395,N_62);
nand U10984 (N_10984,N_2114,N_3529);
nand U10985 (N_10985,N_2201,N_706);
or U10986 (N_10986,N_1985,N_3567);
nor U10987 (N_10987,N_3999,N_5391);
or U10988 (N_10988,N_97,N_5917);
nor U10989 (N_10989,N_3333,N_4941);
nand U10990 (N_10990,N_3202,N_2108);
or U10991 (N_10991,N_5487,N_3762);
nor U10992 (N_10992,N_5138,N_1749);
nor U10993 (N_10993,N_2859,N_3497);
or U10994 (N_10994,N_703,N_3397);
nor U10995 (N_10995,N_2545,N_4916);
nor U10996 (N_10996,N_3556,N_3121);
xnor U10997 (N_10997,N_523,N_1910);
or U10998 (N_10998,N_409,N_350);
or U10999 (N_10999,N_1324,N_776);
or U11000 (N_11000,N_4834,N_1682);
and U11001 (N_11001,N_4798,N_4956);
xor U11002 (N_11002,N_5788,N_4703);
xnor U11003 (N_11003,N_4794,N_5443);
and U11004 (N_11004,N_1435,N_5597);
xnor U11005 (N_11005,N_1094,N_2159);
xor U11006 (N_11006,N_2141,N_2292);
or U11007 (N_11007,N_293,N_3296);
xnor U11008 (N_11008,N_4245,N_4525);
nand U11009 (N_11009,N_3307,N_2879);
nand U11010 (N_11010,N_3688,N_1611);
nand U11011 (N_11011,N_5693,N_3812);
xor U11012 (N_11012,N_3478,N_2550);
or U11013 (N_11013,N_2516,N_2318);
or U11014 (N_11014,N_4888,N_5397);
nor U11015 (N_11015,N_3574,N_3364);
and U11016 (N_11016,N_688,N_975);
xor U11017 (N_11017,N_2364,N_1543);
nand U11018 (N_11018,N_364,N_1621);
xor U11019 (N_11019,N_2669,N_3496);
xnor U11020 (N_11020,N_4691,N_444);
and U11021 (N_11021,N_5244,N_2082);
xnor U11022 (N_11022,N_1277,N_544);
nand U11023 (N_11023,N_3792,N_1147);
xor U11024 (N_11024,N_1258,N_728);
or U11025 (N_11025,N_329,N_4470);
or U11026 (N_11026,N_2348,N_4244);
nand U11027 (N_11027,N_349,N_2748);
nand U11028 (N_11028,N_3212,N_4665);
and U11029 (N_11029,N_3458,N_5736);
nor U11030 (N_11030,N_1049,N_849);
nor U11031 (N_11031,N_2568,N_1123);
and U11032 (N_11032,N_4825,N_1763);
and U11033 (N_11033,N_4669,N_1929);
or U11034 (N_11034,N_4624,N_1101);
xnor U11035 (N_11035,N_732,N_2583);
xor U11036 (N_11036,N_4822,N_2989);
nand U11037 (N_11037,N_3345,N_3106);
nor U11038 (N_11038,N_4333,N_5038);
nand U11039 (N_11039,N_3599,N_4456);
and U11040 (N_11040,N_3536,N_4062);
nand U11041 (N_11041,N_353,N_4642);
nand U11042 (N_11042,N_5979,N_552);
nand U11043 (N_11043,N_4404,N_3425);
and U11044 (N_11044,N_4785,N_3065);
or U11045 (N_11045,N_3586,N_4559);
or U11046 (N_11046,N_1471,N_889);
nor U11047 (N_11047,N_3710,N_916);
and U11048 (N_11048,N_5555,N_5750);
and U11049 (N_11049,N_3248,N_181);
nor U11050 (N_11050,N_5674,N_2204);
xnor U11051 (N_11051,N_5962,N_1567);
nand U11052 (N_11052,N_1044,N_5395);
or U11053 (N_11053,N_1899,N_1064);
nor U11054 (N_11054,N_1532,N_2095);
xnor U11055 (N_11055,N_3645,N_2971);
or U11056 (N_11056,N_1215,N_5801);
and U11057 (N_11057,N_3407,N_4736);
nor U11058 (N_11058,N_1072,N_5820);
nor U11059 (N_11059,N_1248,N_862);
or U11060 (N_11060,N_140,N_4373);
and U11061 (N_11061,N_4186,N_5046);
and U11062 (N_11062,N_5548,N_3759);
nor U11063 (N_11063,N_1611,N_5852);
nand U11064 (N_11064,N_5483,N_3184);
nor U11065 (N_11065,N_860,N_4789);
nand U11066 (N_11066,N_3211,N_27);
xor U11067 (N_11067,N_989,N_4673);
and U11068 (N_11068,N_4481,N_1048);
nand U11069 (N_11069,N_5481,N_2608);
xnor U11070 (N_11070,N_563,N_1891);
xnor U11071 (N_11071,N_2703,N_831);
and U11072 (N_11072,N_1139,N_3234);
nor U11073 (N_11073,N_1248,N_4883);
nor U11074 (N_11074,N_1561,N_4236);
and U11075 (N_11075,N_4432,N_1596);
xnor U11076 (N_11076,N_5493,N_2960);
xor U11077 (N_11077,N_5174,N_1813);
and U11078 (N_11078,N_486,N_1640);
xnor U11079 (N_11079,N_3377,N_3870);
nand U11080 (N_11080,N_2458,N_4102);
and U11081 (N_11081,N_1975,N_4262);
nor U11082 (N_11082,N_572,N_2890);
nand U11083 (N_11083,N_1580,N_4425);
nand U11084 (N_11084,N_5979,N_4002);
nand U11085 (N_11085,N_5624,N_4895);
nand U11086 (N_11086,N_3139,N_1715);
and U11087 (N_11087,N_1791,N_5007);
and U11088 (N_11088,N_3703,N_3763);
nand U11089 (N_11089,N_4102,N_395);
xnor U11090 (N_11090,N_4590,N_4723);
and U11091 (N_11091,N_4386,N_4492);
nor U11092 (N_11092,N_5826,N_2025);
xor U11093 (N_11093,N_3625,N_4899);
or U11094 (N_11094,N_1766,N_3720);
xnor U11095 (N_11095,N_5639,N_1385);
and U11096 (N_11096,N_3093,N_1346);
xnor U11097 (N_11097,N_5924,N_895);
and U11098 (N_11098,N_3346,N_3695);
or U11099 (N_11099,N_2810,N_317);
nor U11100 (N_11100,N_2728,N_4554);
nor U11101 (N_11101,N_4183,N_5598);
nor U11102 (N_11102,N_3811,N_5646);
nand U11103 (N_11103,N_5628,N_384);
and U11104 (N_11104,N_1530,N_5762);
and U11105 (N_11105,N_363,N_2598);
or U11106 (N_11106,N_915,N_4971);
and U11107 (N_11107,N_2165,N_1703);
nor U11108 (N_11108,N_3381,N_656);
nor U11109 (N_11109,N_4282,N_226);
or U11110 (N_11110,N_1198,N_695);
nand U11111 (N_11111,N_5656,N_12);
xor U11112 (N_11112,N_1753,N_2766);
and U11113 (N_11113,N_4870,N_4076);
nand U11114 (N_11114,N_228,N_5339);
and U11115 (N_11115,N_4962,N_2799);
nor U11116 (N_11116,N_210,N_5752);
nor U11117 (N_11117,N_2012,N_1845);
or U11118 (N_11118,N_3208,N_236);
or U11119 (N_11119,N_5365,N_5724);
nor U11120 (N_11120,N_2951,N_4436);
xor U11121 (N_11121,N_2466,N_586);
or U11122 (N_11122,N_1794,N_6);
nand U11123 (N_11123,N_2008,N_2838);
nand U11124 (N_11124,N_1005,N_5785);
nand U11125 (N_11125,N_1554,N_1685);
xor U11126 (N_11126,N_1369,N_3957);
nor U11127 (N_11127,N_435,N_5506);
nor U11128 (N_11128,N_3855,N_624);
nand U11129 (N_11129,N_608,N_4506);
nor U11130 (N_11130,N_3251,N_779);
or U11131 (N_11131,N_102,N_2634);
and U11132 (N_11132,N_5673,N_4335);
nand U11133 (N_11133,N_3461,N_3646);
nor U11134 (N_11134,N_3799,N_3488);
nor U11135 (N_11135,N_5395,N_2128);
xnor U11136 (N_11136,N_3818,N_348);
nor U11137 (N_11137,N_3566,N_2464);
nor U11138 (N_11138,N_3913,N_5324);
nor U11139 (N_11139,N_3419,N_5138);
nand U11140 (N_11140,N_878,N_1179);
or U11141 (N_11141,N_4485,N_635);
and U11142 (N_11142,N_2456,N_2359);
xor U11143 (N_11143,N_4635,N_2998);
or U11144 (N_11144,N_84,N_5291);
or U11145 (N_11145,N_397,N_3790);
nand U11146 (N_11146,N_5863,N_473);
nor U11147 (N_11147,N_251,N_5552);
nor U11148 (N_11148,N_1656,N_4960);
or U11149 (N_11149,N_5889,N_2962);
nand U11150 (N_11150,N_4898,N_4687);
and U11151 (N_11151,N_71,N_3212);
and U11152 (N_11152,N_184,N_4034);
xor U11153 (N_11153,N_1611,N_1946);
nor U11154 (N_11154,N_5588,N_3835);
nor U11155 (N_11155,N_1271,N_5331);
xnor U11156 (N_11156,N_1948,N_258);
nor U11157 (N_11157,N_4921,N_1459);
nand U11158 (N_11158,N_4121,N_1339);
nand U11159 (N_11159,N_4059,N_2597);
nor U11160 (N_11160,N_1676,N_1682);
and U11161 (N_11161,N_1805,N_3296);
or U11162 (N_11162,N_1742,N_5996);
xor U11163 (N_11163,N_1846,N_3445);
nand U11164 (N_11164,N_3467,N_3493);
and U11165 (N_11165,N_186,N_4541);
and U11166 (N_11166,N_5900,N_3764);
nor U11167 (N_11167,N_1830,N_4383);
or U11168 (N_11168,N_3838,N_3985);
xnor U11169 (N_11169,N_164,N_5798);
xor U11170 (N_11170,N_2962,N_2808);
nand U11171 (N_11171,N_1373,N_661);
or U11172 (N_11172,N_205,N_4933);
or U11173 (N_11173,N_1129,N_3391);
xor U11174 (N_11174,N_3025,N_4694);
xor U11175 (N_11175,N_3790,N_5388);
xor U11176 (N_11176,N_5875,N_3269);
xnor U11177 (N_11177,N_3188,N_1790);
nor U11178 (N_11178,N_5764,N_1271);
xnor U11179 (N_11179,N_5328,N_3550);
xor U11180 (N_11180,N_2488,N_3032);
nand U11181 (N_11181,N_988,N_885);
and U11182 (N_11182,N_4253,N_5285);
xor U11183 (N_11183,N_5532,N_1700);
or U11184 (N_11184,N_1961,N_4446);
nor U11185 (N_11185,N_2493,N_3707);
nand U11186 (N_11186,N_5284,N_2429);
xnor U11187 (N_11187,N_4845,N_948);
nor U11188 (N_11188,N_1847,N_482);
xor U11189 (N_11189,N_1041,N_4273);
nor U11190 (N_11190,N_1821,N_1515);
nor U11191 (N_11191,N_3391,N_318);
xor U11192 (N_11192,N_26,N_791);
nor U11193 (N_11193,N_33,N_4654);
nand U11194 (N_11194,N_3392,N_4033);
or U11195 (N_11195,N_5048,N_1359);
xor U11196 (N_11196,N_5511,N_2087);
nor U11197 (N_11197,N_3541,N_3402);
and U11198 (N_11198,N_4645,N_3360);
and U11199 (N_11199,N_2556,N_952);
or U11200 (N_11200,N_4462,N_4189);
nor U11201 (N_11201,N_1411,N_5495);
or U11202 (N_11202,N_3385,N_2571);
nand U11203 (N_11203,N_2441,N_2468);
nand U11204 (N_11204,N_158,N_318);
or U11205 (N_11205,N_3568,N_1902);
or U11206 (N_11206,N_3287,N_4984);
nor U11207 (N_11207,N_1679,N_1627);
xnor U11208 (N_11208,N_2238,N_843);
and U11209 (N_11209,N_164,N_5065);
xnor U11210 (N_11210,N_1053,N_268);
xor U11211 (N_11211,N_2210,N_1392);
nor U11212 (N_11212,N_2125,N_214);
nand U11213 (N_11213,N_3103,N_2402);
xnor U11214 (N_11214,N_90,N_4289);
and U11215 (N_11215,N_3594,N_3282);
or U11216 (N_11216,N_4831,N_3763);
nor U11217 (N_11217,N_1752,N_2554);
xnor U11218 (N_11218,N_987,N_3162);
and U11219 (N_11219,N_1746,N_515);
nor U11220 (N_11220,N_5641,N_2442);
nor U11221 (N_11221,N_389,N_5009);
and U11222 (N_11222,N_1205,N_8);
nor U11223 (N_11223,N_5491,N_360);
nor U11224 (N_11224,N_3351,N_2899);
nor U11225 (N_11225,N_4763,N_744);
nor U11226 (N_11226,N_4474,N_2443);
or U11227 (N_11227,N_4946,N_3055);
nor U11228 (N_11228,N_518,N_1500);
or U11229 (N_11229,N_3265,N_3186);
or U11230 (N_11230,N_4261,N_3381);
nor U11231 (N_11231,N_2063,N_1872);
or U11232 (N_11232,N_3944,N_2075);
xnor U11233 (N_11233,N_4399,N_919);
or U11234 (N_11234,N_4739,N_1796);
nand U11235 (N_11235,N_2060,N_2054);
and U11236 (N_11236,N_268,N_2923);
nor U11237 (N_11237,N_3897,N_5481);
and U11238 (N_11238,N_3468,N_2241);
xor U11239 (N_11239,N_5558,N_350);
nand U11240 (N_11240,N_5439,N_4500);
or U11241 (N_11241,N_5325,N_3280);
xnor U11242 (N_11242,N_4705,N_3924);
nor U11243 (N_11243,N_1174,N_4155);
xor U11244 (N_11244,N_975,N_912);
nor U11245 (N_11245,N_4974,N_2019);
or U11246 (N_11246,N_3324,N_4416);
and U11247 (N_11247,N_1743,N_1957);
nand U11248 (N_11248,N_2863,N_2734);
nor U11249 (N_11249,N_637,N_5022);
or U11250 (N_11250,N_1032,N_4251);
and U11251 (N_11251,N_3608,N_2591);
nor U11252 (N_11252,N_3592,N_5502);
nor U11253 (N_11253,N_2415,N_1470);
xor U11254 (N_11254,N_3119,N_2561);
xnor U11255 (N_11255,N_4483,N_3620);
nor U11256 (N_11256,N_4787,N_634);
or U11257 (N_11257,N_884,N_4359);
nor U11258 (N_11258,N_685,N_994);
and U11259 (N_11259,N_5978,N_738);
and U11260 (N_11260,N_4089,N_2495);
nand U11261 (N_11261,N_4579,N_3724);
nand U11262 (N_11262,N_1126,N_181);
nand U11263 (N_11263,N_36,N_1912);
or U11264 (N_11264,N_5342,N_5133);
nand U11265 (N_11265,N_5671,N_1128);
nand U11266 (N_11266,N_4068,N_1608);
or U11267 (N_11267,N_3375,N_1322);
nor U11268 (N_11268,N_3125,N_1981);
and U11269 (N_11269,N_3958,N_1143);
xor U11270 (N_11270,N_333,N_3786);
or U11271 (N_11271,N_2516,N_1099);
or U11272 (N_11272,N_5336,N_4852);
and U11273 (N_11273,N_553,N_823);
and U11274 (N_11274,N_987,N_830);
nand U11275 (N_11275,N_4507,N_343);
nand U11276 (N_11276,N_416,N_844);
nand U11277 (N_11277,N_4114,N_3311);
xnor U11278 (N_11278,N_1578,N_4123);
nand U11279 (N_11279,N_2721,N_2209);
nor U11280 (N_11280,N_1012,N_4928);
and U11281 (N_11281,N_5733,N_4779);
nor U11282 (N_11282,N_2467,N_2422);
nand U11283 (N_11283,N_5571,N_2205);
nor U11284 (N_11284,N_3599,N_4484);
or U11285 (N_11285,N_1852,N_1623);
xnor U11286 (N_11286,N_4820,N_1596);
or U11287 (N_11287,N_4879,N_657);
nand U11288 (N_11288,N_4785,N_2496);
and U11289 (N_11289,N_4447,N_2707);
or U11290 (N_11290,N_3972,N_2058);
nor U11291 (N_11291,N_2311,N_5304);
nand U11292 (N_11292,N_2786,N_2044);
nand U11293 (N_11293,N_4696,N_2211);
xnor U11294 (N_11294,N_957,N_2902);
or U11295 (N_11295,N_5825,N_650);
nand U11296 (N_11296,N_4071,N_1451);
and U11297 (N_11297,N_3829,N_5851);
nor U11298 (N_11298,N_1594,N_5648);
nor U11299 (N_11299,N_574,N_4497);
and U11300 (N_11300,N_3825,N_3009);
xnor U11301 (N_11301,N_3310,N_3943);
nand U11302 (N_11302,N_5816,N_658);
and U11303 (N_11303,N_2792,N_5465);
xnor U11304 (N_11304,N_5871,N_4296);
or U11305 (N_11305,N_5178,N_1071);
xor U11306 (N_11306,N_1461,N_66);
or U11307 (N_11307,N_5611,N_3159);
nand U11308 (N_11308,N_2509,N_262);
xnor U11309 (N_11309,N_247,N_4176);
or U11310 (N_11310,N_977,N_2887);
nand U11311 (N_11311,N_4381,N_3232);
nand U11312 (N_11312,N_4460,N_3906);
and U11313 (N_11313,N_5723,N_146);
or U11314 (N_11314,N_4489,N_4594);
or U11315 (N_11315,N_2254,N_4965);
and U11316 (N_11316,N_1400,N_4482);
xnor U11317 (N_11317,N_2857,N_5431);
nor U11318 (N_11318,N_5384,N_2797);
nor U11319 (N_11319,N_4907,N_5887);
or U11320 (N_11320,N_2376,N_5030);
xor U11321 (N_11321,N_573,N_1167);
or U11322 (N_11322,N_105,N_4389);
xnor U11323 (N_11323,N_4335,N_3234);
nor U11324 (N_11324,N_341,N_3365);
nor U11325 (N_11325,N_2088,N_1769);
nand U11326 (N_11326,N_5129,N_2859);
or U11327 (N_11327,N_3938,N_735);
nor U11328 (N_11328,N_5145,N_2732);
and U11329 (N_11329,N_1199,N_5336);
and U11330 (N_11330,N_5933,N_4500);
xor U11331 (N_11331,N_5734,N_4404);
or U11332 (N_11332,N_2665,N_3418);
xnor U11333 (N_11333,N_128,N_1048);
and U11334 (N_11334,N_3173,N_4760);
xor U11335 (N_11335,N_5178,N_3691);
xor U11336 (N_11336,N_1120,N_5168);
nor U11337 (N_11337,N_1958,N_2211);
xor U11338 (N_11338,N_1014,N_2172);
and U11339 (N_11339,N_1854,N_2386);
or U11340 (N_11340,N_3087,N_1963);
nand U11341 (N_11341,N_4506,N_5571);
xnor U11342 (N_11342,N_5629,N_4352);
or U11343 (N_11343,N_539,N_3304);
xor U11344 (N_11344,N_4326,N_1363);
and U11345 (N_11345,N_178,N_1581);
and U11346 (N_11346,N_2973,N_2528);
nand U11347 (N_11347,N_5528,N_1649);
nor U11348 (N_11348,N_1317,N_1307);
or U11349 (N_11349,N_3259,N_4183);
or U11350 (N_11350,N_1986,N_5705);
and U11351 (N_11351,N_5350,N_284);
and U11352 (N_11352,N_5391,N_458);
nor U11353 (N_11353,N_830,N_1578);
nor U11354 (N_11354,N_5885,N_2172);
nand U11355 (N_11355,N_1833,N_1096);
and U11356 (N_11356,N_3194,N_221);
nor U11357 (N_11357,N_5826,N_275);
and U11358 (N_11358,N_2922,N_1320);
or U11359 (N_11359,N_1855,N_1933);
nand U11360 (N_11360,N_3681,N_5825);
and U11361 (N_11361,N_336,N_2400);
nor U11362 (N_11362,N_2702,N_403);
xor U11363 (N_11363,N_5376,N_5550);
xor U11364 (N_11364,N_1941,N_3495);
nand U11365 (N_11365,N_2971,N_5824);
and U11366 (N_11366,N_4303,N_246);
nand U11367 (N_11367,N_3029,N_4931);
nand U11368 (N_11368,N_1682,N_1366);
nor U11369 (N_11369,N_4320,N_5760);
and U11370 (N_11370,N_5827,N_5404);
xor U11371 (N_11371,N_1719,N_5972);
xor U11372 (N_11372,N_1360,N_442);
xnor U11373 (N_11373,N_1886,N_979);
nand U11374 (N_11374,N_1543,N_4016);
xnor U11375 (N_11375,N_3832,N_1290);
nand U11376 (N_11376,N_3885,N_2768);
or U11377 (N_11377,N_3346,N_3354);
nand U11378 (N_11378,N_1728,N_3841);
nor U11379 (N_11379,N_62,N_3452);
or U11380 (N_11380,N_871,N_1460);
or U11381 (N_11381,N_4385,N_5803);
or U11382 (N_11382,N_1510,N_5550);
and U11383 (N_11383,N_736,N_1770);
or U11384 (N_11384,N_5911,N_1483);
xor U11385 (N_11385,N_3421,N_587);
nand U11386 (N_11386,N_4641,N_1488);
or U11387 (N_11387,N_224,N_2264);
or U11388 (N_11388,N_3585,N_4800);
nor U11389 (N_11389,N_4926,N_5737);
nand U11390 (N_11390,N_3806,N_1955);
and U11391 (N_11391,N_2463,N_204);
nand U11392 (N_11392,N_5415,N_4014);
or U11393 (N_11393,N_269,N_3592);
nand U11394 (N_11394,N_2587,N_4917);
xnor U11395 (N_11395,N_168,N_4107);
xor U11396 (N_11396,N_1280,N_2822);
xor U11397 (N_11397,N_2064,N_1001);
nor U11398 (N_11398,N_4001,N_2851);
nand U11399 (N_11399,N_1470,N_5337);
or U11400 (N_11400,N_2428,N_929);
xor U11401 (N_11401,N_5901,N_746);
xnor U11402 (N_11402,N_2505,N_5871);
and U11403 (N_11403,N_3654,N_1457);
nand U11404 (N_11404,N_171,N_295);
and U11405 (N_11405,N_334,N_1836);
nor U11406 (N_11406,N_3096,N_3004);
and U11407 (N_11407,N_4690,N_5663);
nand U11408 (N_11408,N_2563,N_2986);
xnor U11409 (N_11409,N_5054,N_2506);
nand U11410 (N_11410,N_2851,N_5348);
and U11411 (N_11411,N_3761,N_1064);
or U11412 (N_11412,N_3428,N_3148);
or U11413 (N_11413,N_1896,N_4862);
and U11414 (N_11414,N_662,N_4604);
nand U11415 (N_11415,N_525,N_4970);
or U11416 (N_11416,N_3291,N_1907);
nor U11417 (N_11417,N_5768,N_1372);
and U11418 (N_11418,N_2928,N_2193);
and U11419 (N_11419,N_39,N_1234);
nor U11420 (N_11420,N_4410,N_1626);
xor U11421 (N_11421,N_843,N_799);
or U11422 (N_11422,N_2268,N_4095);
xnor U11423 (N_11423,N_241,N_2664);
nor U11424 (N_11424,N_5427,N_1180);
and U11425 (N_11425,N_5051,N_5129);
or U11426 (N_11426,N_1831,N_5785);
nor U11427 (N_11427,N_5851,N_5056);
and U11428 (N_11428,N_5465,N_2534);
or U11429 (N_11429,N_4167,N_1105);
or U11430 (N_11430,N_2236,N_1716);
xor U11431 (N_11431,N_4219,N_1213);
xor U11432 (N_11432,N_3096,N_4654);
and U11433 (N_11433,N_1679,N_3325);
and U11434 (N_11434,N_2282,N_3888);
and U11435 (N_11435,N_2042,N_3936);
and U11436 (N_11436,N_1028,N_5951);
nand U11437 (N_11437,N_4960,N_3608);
or U11438 (N_11438,N_5966,N_4565);
nor U11439 (N_11439,N_74,N_1578);
or U11440 (N_11440,N_228,N_2635);
or U11441 (N_11441,N_2206,N_5822);
xnor U11442 (N_11442,N_5315,N_1760);
nor U11443 (N_11443,N_1041,N_1766);
or U11444 (N_11444,N_4282,N_2175);
xnor U11445 (N_11445,N_1645,N_2581);
xnor U11446 (N_11446,N_5428,N_1143);
nor U11447 (N_11447,N_1376,N_5847);
or U11448 (N_11448,N_4317,N_5332);
nand U11449 (N_11449,N_3514,N_3618);
and U11450 (N_11450,N_2382,N_422);
and U11451 (N_11451,N_1407,N_3437);
nand U11452 (N_11452,N_3092,N_3105);
or U11453 (N_11453,N_394,N_3551);
nand U11454 (N_11454,N_5912,N_3812);
nand U11455 (N_11455,N_2523,N_3697);
or U11456 (N_11456,N_175,N_808);
xor U11457 (N_11457,N_3912,N_561);
nand U11458 (N_11458,N_332,N_3000);
xor U11459 (N_11459,N_3309,N_1234);
nand U11460 (N_11460,N_4524,N_5374);
and U11461 (N_11461,N_1135,N_2353);
or U11462 (N_11462,N_2912,N_1299);
and U11463 (N_11463,N_2269,N_2642);
and U11464 (N_11464,N_3624,N_4754);
or U11465 (N_11465,N_3447,N_3145);
and U11466 (N_11466,N_4207,N_149);
or U11467 (N_11467,N_2217,N_1089);
and U11468 (N_11468,N_3648,N_1697);
xor U11469 (N_11469,N_5985,N_3797);
or U11470 (N_11470,N_971,N_4133);
or U11471 (N_11471,N_2524,N_5671);
or U11472 (N_11472,N_3751,N_976);
xor U11473 (N_11473,N_2144,N_4388);
or U11474 (N_11474,N_5518,N_1225);
or U11475 (N_11475,N_4493,N_3106);
and U11476 (N_11476,N_3438,N_74);
or U11477 (N_11477,N_2111,N_1341);
nor U11478 (N_11478,N_1867,N_2538);
nand U11479 (N_11479,N_4597,N_5542);
xnor U11480 (N_11480,N_3800,N_5492);
nand U11481 (N_11481,N_3482,N_4250);
and U11482 (N_11482,N_5004,N_672);
and U11483 (N_11483,N_2663,N_5192);
or U11484 (N_11484,N_119,N_5974);
nand U11485 (N_11485,N_5581,N_92);
or U11486 (N_11486,N_2366,N_802);
xnor U11487 (N_11487,N_2687,N_5649);
nand U11488 (N_11488,N_528,N_2724);
nand U11489 (N_11489,N_3817,N_5175);
and U11490 (N_11490,N_5781,N_4080);
or U11491 (N_11491,N_4334,N_5376);
nor U11492 (N_11492,N_5255,N_5578);
xnor U11493 (N_11493,N_1801,N_5217);
and U11494 (N_11494,N_4520,N_71);
nand U11495 (N_11495,N_3331,N_2637);
nor U11496 (N_11496,N_686,N_2474);
and U11497 (N_11497,N_4508,N_5081);
xnor U11498 (N_11498,N_3730,N_1209);
and U11499 (N_11499,N_915,N_2431);
nand U11500 (N_11500,N_3635,N_3607);
or U11501 (N_11501,N_4635,N_2294);
nand U11502 (N_11502,N_3189,N_799);
or U11503 (N_11503,N_1400,N_5182);
or U11504 (N_11504,N_967,N_239);
or U11505 (N_11505,N_126,N_1131);
or U11506 (N_11506,N_2589,N_4317);
xor U11507 (N_11507,N_117,N_2237);
xor U11508 (N_11508,N_962,N_1907);
or U11509 (N_11509,N_4134,N_1469);
nor U11510 (N_11510,N_3054,N_5942);
xnor U11511 (N_11511,N_5808,N_3418);
nand U11512 (N_11512,N_3605,N_2671);
xnor U11513 (N_11513,N_241,N_3091);
or U11514 (N_11514,N_4516,N_201);
or U11515 (N_11515,N_2700,N_69);
nor U11516 (N_11516,N_1471,N_4345);
and U11517 (N_11517,N_1956,N_4523);
and U11518 (N_11518,N_4745,N_2264);
nor U11519 (N_11519,N_5510,N_1267);
nor U11520 (N_11520,N_4442,N_3875);
and U11521 (N_11521,N_3378,N_1913);
nand U11522 (N_11522,N_4656,N_2225);
nand U11523 (N_11523,N_2139,N_695);
nor U11524 (N_11524,N_451,N_849);
nand U11525 (N_11525,N_3579,N_1695);
or U11526 (N_11526,N_2108,N_977);
nand U11527 (N_11527,N_811,N_4888);
nor U11528 (N_11528,N_3147,N_1115);
nand U11529 (N_11529,N_1024,N_3736);
or U11530 (N_11530,N_4830,N_5169);
xnor U11531 (N_11531,N_2395,N_610);
nor U11532 (N_11532,N_226,N_3167);
and U11533 (N_11533,N_2146,N_3792);
and U11534 (N_11534,N_3959,N_1385);
or U11535 (N_11535,N_1345,N_5439);
nor U11536 (N_11536,N_2877,N_3458);
nor U11537 (N_11537,N_3368,N_4829);
nor U11538 (N_11538,N_48,N_23);
or U11539 (N_11539,N_3862,N_3494);
xor U11540 (N_11540,N_3933,N_4643);
and U11541 (N_11541,N_4843,N_2896);
xnor U11542 (N_11542,N_420,N_5890);
xor U11543 (N_11543,N_2796,N_4258);
xnor U11544 (N_11544,N_4186,N_580);
and U11545 (N_11545,N_3449,N_5733);
and U11546 (N_11546,N_2581,N_5256);
xnor U11547 (N_11547,N_5681,N_4283);
xor U11548 (N_11548,N_5986,N_3427);
nand U11549 (N_11549,N_5019,N_4732);
or U11550 (N_11550,N_4680,N_426);
xnor U11551 (N_11551,N_5318,N_554);
and U11552 (N_11552,N_5872,N_2395);
nor U11553 (N_11553,N_4507,N_1512);
nand U11554 (N_11554,N_5300,N_3433);
and U11555 (N_11555,N_4160,N_2753);
or U11556 (N_11556,N_3857,N_870);
xnor U11557 (N_11557,N_5621,N_2371);
nor U11558 (N_11558,N_281,N_1510);
xor U11559 (N_11559,N_3393,N_4402);
nand U11560 (N_11560,N_1173,N_478);
xnor U11561 (N_11561,N_1994,N_5874);
and U11562 (N_11562,N_3275,N_5723);
and U11563 (N_11563,N_4086,N_1399);
and U11564 (N_11564,N_3211,N_4036);
or U11565 (N_11565,N_2342,N_4138);
nor U11566 (N_11566,N_5716,N_1370);
xor U11567 (N_11567,N_2232,N_3090);
or U11568 (N_11568,N_3593,N_108);
and U11569 (N_11569,N_1509,N_5473);
xnor U11570 (N_11570,N_3240,N_648);
nand U11571 (N_11571,N_2575,N_3368);
xor U11572 (N_11572,N_4173,N_1952);
or U11573 (N_11573,N_5,N_5596);
xnor U11574 (N_11574,N_2905,N_3719);
or U11575 (N_11575,N_3073,N_5089);
nor U11576 (N_11576,N_4600,N_2025);
or U11577 (N_11577,N_5274,N_5778);
nor U11578 (N_11578,N_5763,N_2941);
and U11579 (N_11579,N_597,N_1990);
or U11580 (N_11580,N_2113,N_1927);
nand U11581 (N_11581,N_3555,N_5107);
or U11582 (N_11582,N_2319,N_1869);
nand U11583 (N_11583,N_1766,N_576);
nor U11584 (N_11584,N_2059,N_4074);
and U11585 (N_11585,N_387,N_63);
nand U11586 (N_11586,N_1204,N_4861);
nor U11587 (N_11587,N_1650,N_1887);
nand U11588 (N_11588,N_186,N_1531);
or U11589 (N_11589,N_1905,N_4800);
nand U11590 (N_11590,N_4035,N_1953);
nand U11591 (N_11591,N_3670,N_602);
nor U11592 (N_11592,N_3188,N_2401);
xor U11593 (N_11593,N_3038,N_5674);
nor U11594 (N_11594,N_2263,N_1219);
or U11595 (N_11595,N_5841,N_207);
nand U11596 (N_11596,N_475,N_2085);
and U11597 (N_11597,N_5003,N_5230);
xnor U11598 (N_11598,N_4276,N_5959);
xor U11599 (N_11599,N_4055,N_2875);
nand U11600 (N_11600,N_312,N_4938);
and U11601 (N_11601,N_5030,N_2015);
or U11602 (N_11602,N_3144,N_2153);
xor U11603 (N_11603,N_5170,N_4891);
or U11604 (N_11604,N_1836,N_1631);
or U11605 (N_11605,N_4323,N_3855);
nor U11606 (N_11606,N_3167,N_4037);
or U11607 (N_11607,N_3307,N_3721);
xnor U11608 (N_11608,N_821,N_3392);
xor U11609 (N_11609,N_4438,N_3119);
and U11610 (N_11610,N_1961,N_4421);
and U11611 (N_11611,N_1254,N_4458);
nor U11612 (N_11612,N_2587,N_1967);
and U11613 (N_11613,N_2320,N_2555);
and U11614 (N_11614,N_432,N_235);
nor U11615 (N_11615,N_1050,N_4150);
and U11616 (N_11616,N_4896,N_4890);
or U11617 (N_11617,N_3988,N_3945);
nand U11618 (N_11618,N_3923,N_3908);
and U11619 (N_11619,N_5766,N_3380);
and U11620 (N_11620,N_909,N_2346);
nand U11621 (N_11621,N_3848,N_4545);
or U11622 (N_11622,N_3781,N_4262);
xnor U11623 (N_11623,N_4771,N_4292);
and U11624 (N_11624,N_637,N_5562);
or U11625 (N_11625,N_1840,N_1087);
nor U11626 (N_11626,N_5072,N_2052);
nand U11627 (N_11627,N_3523,N_1815);
and U11628 (N_11628,N_2096,N_5574);
xor U11629 (N_11629,N_1352,N_799);
xnor U11630 (N_11630,N_262,N_5885);
nand U11631 (N_11631,N_5771,N_499);
nor U11632 (N_11632,N_509,N_5293);
and U11633 (N_11633,N_2402,N_3618);
nand U11634 (N_11634,N_2138,N_5069);
nand U11635 (N_11635,N_4964,N_5750);
nor U11636 (N_11636,N_1108,N_2200);
and U11637 (N_11637,N_5620,N_2851);
xnor U11638 (N_11638,N_4268,N_2542);
nor U11639 (N_11639,N_3054,N_154);
nor U11640 (N_11640,N_1733,N_493);
nor U11641 (N_11641,N_2152,N_5842);
or U11642 (N_11642,N_651,N_866);
nand U11643 (N_11643,N_1200,N_1398);
xor U11644 (N_11644,N_2881,N_3775);
or U11645 (N_11645,N_2506,N_4789);
nor U11646 (N_11646,N_2861,N_2284);
or U11647 (N_11647,N_3675,N_1945);
xor U11648 (N_11648,N_2699,N_1786);
nor U11649 (N_11649,N_3959,N_5826);
xnor U11650 (N_11650,N_1785,N_2236);
xor U11651 (N_11651,N_2237,N_5010);
nand U11652 (N_11652,N_5152,N_5664);
or U11653 (N_11653,N_3179,N_5322);
nand U11654 (N_11654,N_3503,N_2210);
and U11655 (N_11655,N_5850,N_1952);
xnor U11656 (N_11656,N_2944,N_910);
xor U11657 (N_11657,N_3207,N_631);
and U11658 (N_11658,N_3018,N_5792);
nor U11659 (N_11659,N_2614,N_3723);
and U11660 (N_11660,N_1296,N_3698);
nor U11661 (N_11661,N_1263,N_930);
xor U11662 (N_11662,N_3442,N_927);
xor U11663 (N_11663,N_1497,N_2786);
and U11664 (N_11664,N_4672,N_1360);
nand U11665 (N_11665,N_2351,N_4078);
nor U11666 (N_11666,N_165,N_858);
nor U11667 (N_11667,N_5970,N_3069);
nand U11668 (N_11668,N_1924,N_545);
nand U11669 (N_11669,N_1788,N_1975);
nor U11670 (N_11670,N_4702,N_4950);
or U11671 (N_11671,N_1201,N_2615);
nand U11672 (N_11672,N_4046,N_5013);
and U11673 (N_11673,N_436,N_522);
nand U11674 (N_11674,N_3347,N_5496);
or U11675 (N_11675,N_5437,N_2375);
xnor U11676 (N_11676,N_2255,N_4550);
xor U11677 (N_11677,N_2999,N_2313);
nand U11678 (N_11678,N_3338,N_2338);
xor U11679 (N_11679,N_5399,N_4305);
xor U11680 (N_11680,N_3396,N_3309);
and U11681 (N_11681,N_5605,N_4446);
nand U11682 (N_11682,N_5536,N_5817);
xnor U11683 (N_11683,N_4898,N_1705);
nand U11684 (N_11684,N_969,N_5065);
or U11685 (N_11685,N_5753,N_2017);
and U11686 (N_11686,N_3667,N_3045);
xor U11687 (N_11687,N_2245,N_1718);
xor U11688 (N_11688,N_3462,N_5881);
and U11689 (N_11689,N_2587,N_4244);
nor U11690 (N_11690,N_1500,N_4542);
nand U11691 (N_11691,N_5654,N_4377);
nor U11692 (N_11692,N_5261,N_4723);
nand U11693 (N_11693,N_1036,N_1660);
nand U11694 (N_11694,N_146,N_1107);
nand U11695 (N_11695,N_132,N_1008);
nand U11696 (N_11696,N_882,N_2836);
xor U11697 (N_11697,N_2192,N_1600);
xor U11698 (N_11698,N_3693,N_4126);
nand U11699 (N_11699,N_4250,N_3094);
xnor U11700 (N_11700,N_16,N_5179);
nor U11701 (N_11701,N_5779,N_814);
xor U11702 (N_11702,N_5968,N_2320);
nand U11703 (N_11703,N_4780,N_5341);
and U11704 (N_11704,N_4257,N_1089);
and U11705 (N_11705,N_4622,N_3594);
and U11706 (N_11706,N_986,N_882);
or U11707 (N_11707,N_1622,N_376);
nor U11708 (N_11708,N_1687,N_1891);
or U11709 (N_11709,N_5526,N_3780);
or U11710 (N_11710,N_776,N_2185);
xnor U11711 (N_11711,N_4260,N_3900);
nand U11712 (N_11712,N_1731,N_1834);
nor U11713 (N_11713,N_3614,N_5422);
and U11714 (N_11714,N_1464,N_1251);
or U11715 (N_11715,N_5892,N_2010);
and U11716 (N_11716,N_66,N_1612);
nand U11717 (N_11717,N_3222,N_3987);
nand U11718 (N_11718,N_5541,N_933);
or U11719 (N_11719,N_1664,N_3460);
nor U11720 (N_11720,N_103,N_3108);
and U11721 (N_11721,N_1058,N_1071);
nand U11722 (N_11722,N_2806,N_5691);
xnor U11723 (N_11723,N_5827,N_926);
and U11724 (N_11724,N_155,N_2545);
and U11725 (N_11725,N_3241,N_2014);
nand U11726 (N_11726,N_4165,N_3436);
nand U11727 (N_11727,N_2720,N_4071);
and U11728 (N_11728,N_3292,N_488);
and U11729 (N_11729,N_3064,N_3273);
and U11730 (N_11730,N_1728,N_479);
nand U11731 (N_11731,N_2255,N_4796);
or U11732 (N_11732,N_2228,N_1450);
nor U11733 (N_11733,N_4127,N_2);
nand U11734 (N_11734,N_375,N_1245);
xor U11735 (N_11735,N_4038,N_1518);
nand U11736 (N_11736,N_1916,N_716);
nor U11737 (N_11737,N_1917,N_5474);
nand U11738 (N_11738,N_3025,N_5675);
xnor U11739 (N_11739,N_614,N_1645);
or U11740 (N_11740,N_3427,N_1705);
nor U11741 (N_11741,N_1789,N_1278);
nand U11742 (N_11742,N_636,N_534);
nor U11743 (N_11743,N_985,N_2949);
or U11744 (N_11744,N_798,N_4992);
or U11745 (N_11745,N_4872,N_935);
and U11746 (N_11746,N_706,N_380);
or U11747 (N_11747,N_3,N_1469);
nor U11748 (N_11748,N_5084,N_2520);
or U11749 (N_11749,N_1474,N_3869);
xnor U11750 (N_11750,N_80,N_5844);
nor U11751 (N_11751,N_3263,N_4183);
nand U11752 (N_11752,N_2883,N_3124);
and U11753 (N_11753,N_1377,N_110);
nor U11754 (N_11754,N_5026,N_2412);
nand U11755 (N_11755,N_397,N_4909);
or U11756 (N_11756,N_4983,N_5096);
nor U11757 (N_11757,N_2393,N_3979);
nand U11758 (N_11758,N_5978,N_5794);
nand U11759 (N_11759,N_1058,N_5728);
xnor U11760 (N_11760,N_3615,N_5796);
xnor U11761 (N_11761,N_2972,N_1846);
or U11762 (N_11762,N_2367,N_5617);
nor U11763 (N_11763,N_1255,N_1447);
nand U11764 (N_11764,N_7,N_441);
and U11765 (N_11765,N_186,N_1746);
nand U11766 (N_11766,N_4986,N_1856);
nor U11767 (N_11767,N_61,N_1840);
nor U11768 (N_11768,N_2486,N_3668);
nor U11769 (N_11769,N_2799,N_1780);
nor U11770 (N_11770,N_4045,N_966);
nor U11771 (N_11771,N_4132,N_447);
nor U11772 (N_11772,N_1946,N_1422);
and U11773 (N_11773,N_2758,N_804);
nor U11774 (N_11774,N_5746,N_2624);
or U11775 (N_11775,N_2124,N_3309);
xnor U11776 (N_11776,N_5569,N_2134);
or U11777 (N_11777,N_3010,N_2172);
nand U11778 (N_11778,N_4027,N_1817);
nand U11779 (N_11779,N_4755,N_3000);
nor U11780 (N_11780,N_4548,N_807);
and U11781 (N_11781,N_281,N_5140);
or U11782 (N_11782,N_636,N_2852);
nor U11783 (N_11783,N_2342,N_2691);
and U11784 (N_11784,N_3307,N_3261);
xnor U11785 (N_11785,N_1038,N_1984);
xnor U11786 (N_11786,N_4862,N_455);
nor U11787 (N_11787,N_3082,N_2820);
or U11788 (N_11788,N_3823,N_887);
nor U11789 (N_11789,N_222,N_2578);
nor U11790 (N_11790,N_4766,N_5980);
and U11791 (N_11791,N_1841,N_4041);
nand U11792 (N_11792,N_5785,N_3328);
xnor U11793 (N_11793,N_4817,N_1200);
or U11794 (N_11794,N_4453,N_1659);
xor U11795 (N_11795,N_3244,N_4076);
nor U11796 (N_11796,N_2158,N_5790);
xnor U11797 (N_11797,N_1582,N_4707);
xnor U11798 (N_11798,N_2492,N_4141);
or U11799 (N_11799,N_5442,N_1951);
and U11800 (N_11800,N_5169,N_2241);
nand U11801 (N_11801,N_4675,N_1295);
nor U11802 (N_11802,N_3107,N_581);
and U11803 (N_11803,N_2495,N_3852);
and U11804 (N_11804,N_4230,N_2396);
and U11805 (N_11805,N_4215,N_3474);
or U11806 (N_11806,N_5739,N_257);
or U11807 (N_11807,N_675,N_3873);
and U11808 (N_11808,N_2802,N_4473);
xnor U11809 (N_11809,N_1376,N_1395);
xnor U11810 (N_11810,N_1727,N_5500);
or U11811 (N_11811,N_4777,N_3315);
or U11812 (N_11812,N_1297,N_574);
nor U11813 (N_11813,N_3741,N_1690);
nand U11814 (N_11814,N_5972,N_2651);
and U11815 (N_11815,N_5136,N_5173);
nand U11816 (N_11816,N_4413,N_1168);
xnor U11817 (N_11817,N_1598,N_1350);
nor U11818 (N_11818,N_5970,N_1448);
or U11819 (N_11819,N_2120,N_1649);
and U11820 (N_11820,N_4663,N_4130);
nor U11821 (N_11821,N_5545,N_5303);
nor U11822 (N_11822,N_4613,N_2061);
and U11823 (N_11823,N_5617,N_2553);
or U11824 (N_11824,N_2132,N_877);
and U11825 (N_11825,N_4815,N_3673);
nor U11826 (N_11826,N_4607,N_3166);
xnor U11827 (N_11827,N_5840,N_5364);
nand U11828 (N_11828,N_5478,N_1619);
or U11829 (N_11829,N_3526,N_1624);
and U11830 (N_11830,N_3622,N_3751);
nor U11831 (N_11831,N_5162,N_5987);
or U11832 (N_11832,N_3982,N_3777);
nand U11833 (N_11833,N_2899,N_5064);
and U11834 (N_11834,N_3834,N_4696);
or U11835 (N_11835,N_3748,N_1986);
xnor U11836 (N_11836,N_3949,N_2334);
xor U11837 (N_11837,N_1888,N_4624);
or U11838 (N_11838,N_1820,N_1824);
xor U11839 (N_11839,N_30,N_5897);
or U11840 (N_11840,N_4255,N_2723);
and U11841 (N_11841,N_4253,N_1422);
and U11842 (N_11842,N_3609,N_5288);
nand U11843 (N_11843,N_4020,N_2175);
and U11844 (N_11844,N_4751,N_3995);
nor U11845 (N_11845,N_5068,N_1345);
or U11846 (N_11846,N_782,N_4689);
or U11847 (N_11847,N_5822,N_4626);
or U11848 (N_11848,N_1676,N_5152);
xnor U11849 (N_11849,N_1118,N_3183);
and U11850 (N_11850,N_3020,N_1774);
or U11851 (N_11851,N_2760,N_1020);
xor U11852 (N_11852,N_1058,N_3291);
nand U11853 (N_11853,N_3298,N_5286);
or U11854 (N_11854,N_3679,N_3775);
and U11855 (N_11855,N_3751,N_5886);
xor U11856 (N_11856,N_462,N_4423);
nor U11857 (N_11857,N_2139,N_1727);
xnor U11858 (N_11858,N_418,N_3945);
xnor U11859 (N_11859,N_661,N_4449);
nor U11860 (N_11860,N_1170,N_3899);
and U11861 (N_11861,N_905,N_5858);
and U11862 (N_11862,N_3267,N_1741);
nand U11863 (N_11863,N_4350,N_5165);
nand U11864 (N_11864,N_893,N_5587);
xnor U11865 (N_11865,N_560,N_5720);
and U11866 (N_11866,N_1726,N_3162);
or U11867 (N_11867,N_629,N_1815);
and U11868 (N_11868,N_1237,N_2464);
and U11869 (N_11869,N_640,N_4925);
nor U11870 (N_11870,N_2354,N_4325);
nor U11871 (N_11871,N_4162,N_5775);
or U11872 (N_11872,N_2751,N_4649);
and U11873 (N_11873,N_4183,N_3059);
or U11874 (N_11874,N_3653,N_5718);
xor U11875 (N_11875,N_4730,N_3395);
xor U11876 (N_11876,N_3826,N_4055);
and U11877 (N_11877,N_1393,N_2992);
and U11878 (N_11878,N_718,N_5641);
nand U11879 (N_11879,N_1381,N_1361);
xnor U11880 (N_11880,N_985,N_1120);
nand U11881 (N_11881,N_3875,N_43);
and U11882 (N_11882,N_5322,N_5784);
nand U11883 (N_11883,N_658,N_4307);
and U11884 (N_11884,N_1145,N_1060);
xor U11885 (N_11885,N_5866,N_5830);
nand U11886 (N_11886,N_5902,N_594);
or U11887 (N_11887,N_5429,N_4459);
or U11888 (N_11888,N_5267,N_3634);
xor U11889 (N_11889,N_3924,N_2847);
nand U11890 (N_11890,N_3273,N_3017);
nor U11891 (N_11891,N_5902,N_4710);
nand U11892 (N_11892,N_1439,N_1178);
and U11893 (N_11893,N_5483,N_3134);
nor U11894 (N_11894,N_4430,N_5708);
nand U11895 (N_11895,N_4061,N_3244);
xnor U11896 (N_11896,N_545,N_5271);
xor U11897 (N_11897,N_406,N_725);
xnor U11898 (N_11898,N_1927,N_767);
nand U11899 (N_11899,N_2417,N_1371);
xor U11900 (N_11900,N_3168,N_3465);
or U11901 (N_11901,N_2624,N_3806);
nand U11902 (N_11902,N_2389,N_5250);
nor U11903 (N_11903,N_65,N_2689);
and U11904 (N_11904,N_4791,N_3188);
and U11905 (N_11905,N_35,N_5250);
xor U11906 (N_11906,N_2959,N_5311);
nand U11907 (N_11907,N_3257,N_763);
nor U11908 (N_11908,N_4485,N_1564);
xor U11909 (N_11909,N_3584,N_5788);
xnor U11910 (N_11910,N_5895,N_2574);
and U11911 (N_11911,N_1945,N_3144);
and U11912 (N_11912,N_5121,N_3085);
xnor U11913 (N_11913,N_2351,N_2983);
nand U11914 (N_11914,N_1651,N_5821);
xnor U11915 (N_11915,N_4742,N_439);
and U11916 (N_11916,N_3937,N_4403);
nor U11917 (N_11917,N_5160,N_4546);
and U11918 (N_11918,N_59,N_1667);
and U11919 (N_11919,N_4681,N_3907);
nand U11920 (N_11920,N_5382,N_4455);
nand U11921 (N_11921,N_4918,N_707);
xor U11922 (N_11922,N_569,N_1705);
nand U11923 (N_11923,N_804,N_172);
nor U11924 (N_11924,N_4190,N_216);
xnor U11925 (N_11925,N_3567,N_2598);
or U11926 (N_11926,N_2742,N_3666);
or U11927 (N_11927,N_519,N_4604);
nor U11928 (N_11928,N_3317,N_2677);
nor U11929 (N_11929,N_5194,N_2454);
xnor U11930 (N_11930,N_4374,N_3371);
or U11931 (N_11931,N_1386,N_5617);
nand U11932 (N_11932,N_5545,N_5464);
nand U11933 (N_11933,N_2,N_3775);
nor U11934 (N_11934,N_2487,N_4025);
and U11935 (N_11935,N_3296,N_1950);
or U11936 (N_11936,N_3114,N_4490);
and U11937 (N_11937,N_623,N_5967);
xor U11938 (N_11938,N_1931,N_1647);
nor U11939 (N_11939,N_5457,N_3936);
or U11940 (N_11940,N_5353,N_5372);
or U11941 (N_11941,N_1305,N_3684);
and U11942 (N_11942,N_3728,N_501);
and U11943 (N_11943,N_3286,N_689);
or U11944 (N_11944,N_274,N_3286);
nor U11945 (N_11945,N_5658,N_319);
or U11946 (N_11946,N_5984,N_3315);
or U11947 (N_11947,N_5727,N_4989);
or U11948 (N_11948,N_1778,N_2423);
nand U11949 (N_11949,N_1646,N_1220);
or U11950 (N_11950,N_3602,N_1294);
or U11951 (N_11951,N_5689,N_3054);
nand U11952 (N_11952,N_4931,N_5635);
xor U11953 (N_11953,N_1950,N_2991);
nor U11954 (N_11954,N_767,N_2836);
and U11955 (N_11955,N_4521,N_2952);
or U11956 (N_11956,N_5371,N_4375);
nand U11957 (N_11957,N_5982,N_5322);
xnor U11958 (N_11958,N_1492,N_5347);
xnor U11959 (N_11959,N_1575,N_2419);
and U11960 (N_11960,N_224,N_4466);
nor U11961 (N_11961,N_2272,N_4919);
or U11962 (N_11962,N_1638,N_1647);
xor U11963 (N_11963,N_1566,N_2228);
or U11964 (N_11964,N_5017,N_170);
or U11965 (N_11965,N_5093,N_1372);
xnor U11966 (N_11966,N_3600,N_1657);
and U11967 (N_11967,N_2765,N_1914);
xor U11968 (N_11968,N_2976,N_4232);
xor U11969 (N_11969,N_4888,N_3641);
and U11970 (N_11970,N_1362,N_5491);
xnor U11971 (N_11971,N_1449,N_5487);
or U11972 (N_11972,N_3466,N_3335);
nand U11973 (N_11973,N_60,N_3031);
xnor U11974 (N_11974,N_1117,N_860);
nor U11975 (N_11975,N_2605,N_5607);
nor U11976 (N_11976,N_1738,N_1636);
nor U11977 (N_11977,N_1359,N_2692);
and U11978 (N_11978,N_2633,N_4159);
or U11979 (N_11979,N_745,N_666);
nand U11980 (N_11980,N_5352,N_1629);
xnor U11981 (N_11981,N_3504,N_5683);
or U11982 (N_11982,N_5404,N_1919);
xnor U11983 (N_11983,N_4457,N_5434);
xnor U11984 (N_11984,N_3509,N_1703);
or U11985 (N_11985,N_36,N_5831);
nor U11986 (N_11986,N_5701,N_4404);
or U11987 (N_11987,N_3087,N_4029);
or U11988 (N_11988,N_3385,N_1191);
nor U11989 (N_11989,N_3292,N_3594);
xor U11990 (N_11990,N_1620,N_2401);
or U11991 (N_11991,N_5166,N_1479);
or U11992 (N_11992,N_3677,N_5364);
and U11993 (N_11993,N_2941,N_5740);
nand U11994 (N_11994,N_2162,N_2901);
nand U11995 (N_11995,N_5188,N_710);
nor U11996 (N_11996,N_1591,N_1908);
nor U11997 (N_11997,N_1315,N_1313);
nand U11998 (N_11998,N_1871,N_5579);
xnor U11999 (N_11999,N_2602,N_3984);
and U12000 (N_12000,N_8146,N_8516);
nand U12001 (N_12001,N_10922,N_6616);
xor U12002 (N_12002,N_7083,N_6182);
nor U12003 (N_12003,N_10761,N_9375);
or U12004 (N_12004,N_9490,N_7649);
or U12005 (N_12005,N_8561,N_10058);
nand U12006 (N_12006,N_6023,N_9715);
and U12007 (N_12007,N_8399,N_7463);
nor U12008 (N_12008,N_10814,N_9571);
nand U12009 (N_12009,N_10684,N_11087);
nand U12010 (N_12010,N_9338,N_10030);
nor U12011 (N_12011,N_6793,N_11537);
or U12012 (N_12012,N_6375,N_10393);
nand U12013 (N_12013,N_8330,N_7330);
or U12014 (N_12014,N_9155,N_9021);
nand U12015 (N_12015,N_11754,N_8385);
or U12016 (N_12016,N_11008,N_9546);
xor U12017 (N_12017,N_6998,N_7513);
xor U12018 (N_12018,N_9769,N_8938);
or U12019 (N_12019,N_7319,N_7071);
or U12020 (N_12020,N_11112,N_11368);
and U12021 (N_12021,N_10890,N_8735);
and U12022 (N_12022,N_7087,N_7064);
nand U12023 (N_12023,N_10924,N_9753);
nor U12024 (N_12024,N_11733,N_6573);
nand U12025 (N_12025,N_6835,N_9694);
xor U12026 (N_12026,N_6963,N_8960);
nor U12027 (N_12027,N_10698,N_9685);
or U12028 (N_12028,N_11883,N_11435);
nor U12029 (N_12029,N_9859,N_7677);
nor U12030 (N_12030,N_9201,N_7050);
nor U12031 (N_12031,N_7156,N_11329);
nor U12032 (N_12032,N_10448,N_10589);
and U12033 (N_12033,N_6501,N_11571);
or U12034 (N_12034,N_9506,N_11132);
nand U12035 (N_12035,N_6489,N_8693);
nor U12036 (N_12036,N_9582,N_7868);
and U12037 (N_12037,N_9622,N_10450);
xor U12038 (N_12038,N_8916,N_9364);
xor U12039 (N_12039,N_6643,N_6527);
nand U12040 (N_12040,N_9829,N_10179);
and U12041 (N_12041,N_7914,N_11715);
nor U12042 (N_12042,N_9004,N_9600);
xnor U12043 (N_12043,N_10380,N_6220);
xor U12044 (N_12044,N_7538,N_10577);
or U12045 (N_12045,N_10999,N_10488);
or U12046 (N_12046,N_6048,N_8336);
nand U12047 (N_12047,N_7865,N_11876);
and U12048 (N_12048,N_7630,N_9119);
or U12049 (N_12049,N_8768,N_6286);
or U12050 (N_12050,N_7490,N_7522);
nor U12051 (N_12051,N_8535,N_6192);
or U12052 (N_12052,N_7237,N_10257);
xor U12053 (N_12053,N_10797,N_7024);
nand U12054 (N_12054,N_8003,N_7375);
nor U12055 (N_12055,N_6332,N_9505);
nand U12056 (N_12056,N_9325,N_10171);
xnor U12057 (N_12057,N_7235,N_11152);
nand U12058 (N_12058,N_11682,N_11190);
xor U12059 (N_12059,N_10403,N_6629);
and U12060 (N_12060,N_9792,N_10462);
nand U12061 (N_12061,N_8449,N_9232);
nand U12062 (N_12062,N_11014,N_10127);
xnor U12063 (N_12063,N_7027,N_7048);
xnor U12064 (N_12064,N_9326,N_10433);
xnor U12065 (N_12065,N_7858,N_10702);
nor U12066 (N_12066,N_11969,N_7180);
nand U12067 (N_12067,N_6498,N_8346);
or U12068 (N_12068,N_8813,N_10222);
or U12069 (N_12069,N_8817,N_9065);
nand U12070 (N_12070,N_8181,N_9175);
nand U12071 (N_12071,N_7433,N_7898);
nand U12072 (N_12072,N_9118,N_11243);
and U12073 (N_12073,N_9482,N_6738);
and U12074 (N_12074,N_6030,N_7049);
xnor U12075 (N_12075,N_9510,N_11166);
or U12076 (N_12076,N_10697,N_6411);
xnor U12077 (N_12077,N_10156,N_9708);
nand U12078 (N_12078,N_10184,N_6890);
nor U12079 (N_12079,N_9634,N_9768);
nand U12080 (N_12080,N_6709,N_7567);
xnor U12081 (N_12081,N_6370,N_9337);
nand U12082 (N_12082,N_10015,N_8446);
and U12083 (N_12083,N_6311,N_6927);
xor U12084 (N_12084,N_6318,N_9635);
xnor U12085 (N_12085,N_6471,N_9186);
and U12086 (N_12086,N_9152,N_8224);
or U12087 (N_12087,N_11099,N_11489);
nor U12088 (N_12088,N_8404,N_7878);
nand U12089 (N_12089,N_9268,N_7403);
nand U12090 (N_12090,N_6851,N_10266);
and U12091 (N_12091,N_9128,N_10031);
nor U12092 (N_12092,N_10777,N_9327);
nor U12093 (N_12093,N_6455,N_11987);
and U12094 (N_12094,N_8295,N_10636);
nor U12095 (N_12095,N_8176,N_9380);
and U12096 (N_12096,N_10330,N_10224);
xor U12097 (N_12097,N_8485,N_11332);
xor U12098 (N_12098,N_9568,N_7446);
nor U12099 (N_12099,N_8034,N_7933);
or U12100 (N_12100,N_8131,N_9484);
or U12101 (N_12101,N_9242,N_8286);
xnor U12102 (N_12102,N_7352,N_10319);
and U12103 (N_12103,N_11211,N_9609);
nor U12104 (N_12104,N_8673,N_7041);
nor U12105 (N_12105,N_8434,N_7571);
xnor U12106 (N_12106,N_7263,N_9025);
nand U12107 (N_12107,N_10437,N_9725);
nand U12108 (N_12108,N_8808,N_8028);
and U12109 (N_12109,N_7026,N_8431);
nand U12110 (N_12110,N_8806,N_6559);
or U12111 (N_12111,N_7427,N_10677);
nor U12112 (N_12112,N_8284,N_7657);
and U12113 (N_12113,N_10893,N_11017);
nand U12114 (N_12114,N_8581,N_7275);
xor U12115 (N_12115,N_11028,N_10861);
nand U12116 (N_12116,N_6980,N_9028);
xor U12117 (N_12117,N_6625,N_11766);
nor U12118 (N_12118,N_7569,N_8403);
nor U12119 (N_12119,N_11413,N_10857);
or U12120 (N_12120,N_8054,N_10102);
and U12121 (N_12121,N_9778,N_11718);
xor U12122 (N_12122,N_10824,N_6670);
nor U12123 (N_12123,N_7122,N_10440);
nor U12124 (N_12124,N_9504,N_10232);
nand U12125 (N_12125,N_9147,N_7240);
xnor U12126 (N_12126,N_11869,N_10091);
and U12127 (N_12127,N_8700,N_7272);
nor U12128 (N_12128,N_11418,N_10351);
nand U12129 (N_12129,N_11314,N_7756);
nor U12130 (N_12130,N_10788,N_11130);
nand U12131 (N_12131,N_10162,N_6881);
and U12132 (N_12132,N_10167,N_6758);
xor U12133 (N_12133,N_8216,N_8629);
nand U12134 (N_12134,N_10760,N_8958);
and U12135 (N_12135,N_10001,N_9771);
nand U12136 (N_12136,N_8202,N_7553);
xnor U12137 (N_12137,N_10226,N_6033);
nand U12138 (N_12138,N_8745,N_9370);
nand U12139 (N_12139,N_9400,N_7256);
or U12140 (N_12140,N_8245,N_8942);
nand U12141 (N_12141,N_6502,N_6212);
nand U12142 (N_12142,N_7701,N_9717);
or U12143 (N_12143,N_8635,N_7721);
nor U12144 (N_12144,N_8848,N_6968);
and U12145 (N_12145,N_6706,N_9744);
nor U12146 (N_12146,N_8133,N_8225);
nor U12147 (N_12147,N_7036,N_6158);
nand U12148 (N_12148,N_9463,N_11351);
xnor U12149 (N_12149,N_7825,N_7796);
and U12150 (N_12150,N_8513,N_10984);
or U12151 (N_12151,N_11509,N_11444);
xor U12152 (N_12152,N_10988,N_6976);
nand U12153 (N_12153,N_6753,N_11621);
nand U12154 (N_12154,N_8904,N_11086);
and U12155 (N_12155,N_11762,N_8596);
xnor U12156 (N_12156,N_6691,N_11336);
or U12157 (N_12157,N_6729,N_11209);
xnor U12158 (N_12158,N_10856,N_10611);
nor U12159 (N_12159,N_6148,N_9023);
nor U12160 (N_12160,N_8753,N_6909);
and U12161 (N_12161,N_6293,N_8788);
xor U12162 (N_12162,N_11731,N_6591);
and U12163 (N_12163,N_10242,N_8272);
and U12164 (N_12164,N_7264,N_10308);
nand U12165 (N_12165,N_8274,N_7607);
xor U12166 (N_12166,N_10275,N_11390);
and U12167 (N_12167,N_8889,N_10656);
nor U12168 (N_12168,N_11089,N_6662);
xor U12169 (N_12169,N_10818,N_7851);
nand U12170 (N_12170,N_9449,N_7199);
or U12171 (N_12171,N_6693,N_10303);
xnor U12172 (N_12172,N_10635,N_9251);
or U12173 (N_12173,N_11233,N_6154);
or U12174 (N_12174,N_11524,N_9237);
nand U12175 (N_12175,N_11349,N_8876);
and U12176 (N_12176,N_10496,N_9098);
nor U12177 (N_12177,N_8812,N_6389);
xor U12178 (N_12178,N_9150,N_7430);
nor U12179 (N_12179,N_8429,N_9354);
xnor U12180 (N_12180,N_6805,N_8487);
and U12181 (N_12181,N_8572,N_11823);
nand U12182 (N_12182,N_9450,N_11281);
or U12183 (N_12183,N_7231,N_8549);
or U12184 (N_12184,N_9143,N_11931);
or U12185 (N_12185,N_6514,N_11882);
nor U12186 (N_12186,N_11143,N_7273);
nor U12187 (N_12187,N_6407,N_11309);
or U12188 (N_12188,N_10143,N_7932);
xor U12189 (N_12189,N_10871,N_8332);
nor U12190 (N_12190,N_11171,N_10479);
nand U12191 (N_12191,N_10534,N_9094);
or U12192 (N_12192,N_8348,N_7872);
nand U12193 (N_12193,N_10367,N_8379);
xnor U12194 (N_12194,N_11664,N_7722);
and U12195 (N_12195,N_7303,N_8619);
xor U12196 (N_12196,N_10585,N_8577);
and U12197 (N_12197,N_8939,N_6075);
nand U12198 (N_12198,N_6928,N_8398);
nor U12199 (N_12199,N_7092,N_8903);
nor U12200 (N_12200,N_11277,N_6213);
nor U12201 (N_12201,N_7090,N_10352);
or U12202 (N_12202,N_11949,N_9418);
nand U12203 (N_12203,N_10418,N_7012);
xor U12204 (N_12204,N_11051,N_9131);
xor U12205 (N_12205,N_11848,N_7670);
nor U12206 (N_12206,N_8732,N_6701);
nand U12207 (N_12207,N_6045,N_6235);
nand U12208 (N_12208,N_11575,N_8575);
nor U12209 (N_12209,N_8105,N_11486);
nand U12210 (N_12210,N_7008,N_6133);
nand U12211 (N_12211,N_9036,N_7308);
nand U12212 (N_12212,N_8502,N_10630);
nand U12213 (N_12213,N_10100,N_6579);
or U12214 (N_12214,N_6565,N_9979);
and U12215 (N_12215,N_10569,N_11153);
nor U12216 (N_12216,N_7009,N_11915);
or U12217 (N_12217,N_11710,N_9987);
nand U12218 (N_12218,N_10020,N_10620);
and U12219 (N_12219,N_10688,N_6827);
nor U12220 (N_12220,N_8857,N_10685);
nor U12221 (N_12221,N_8068,N_9466);
nor U12222 (N_12222,N_6686,N_8305);
and U12223 (N_12223,N_8165,N_10512);
or U12224 (N_12224,N_8603,N_11124);
or U12225 (N_12225,N_9933,N_11777);
and U12226 (N_12226,N_6530,N_6143);
xnor U12227 (N_12227,N_11021,N_9525);
nor U12228 (N_12228,N_10157,N_10672);
xnor U12229 (N_12229,N_7713,N_7334);
or U12230 (N_12230,N_10757,N_8791);
xnor U12231 (N_12231,N_6683,N_9460);
nor U12232 (N_12232,N_8759,N_11272);
and U12233 (N_12233,N_9730,N_11307);
nor U12234 (N_12234,N_10465,N_8369);
and U12235 (N_12235,N_8175,N_11903);
xor U12236 (N_12236,N_11020,N_6113);
and U12237 (N_12237,N_10798,N_11866);
nand U12238 (N_12238,N_9937,N_6297);
nand U12239 (N_12239,N_9688,N_7007);
or U12240 (N_12240,N_7472,N_11078);
and U12241 (N_12241,N_8643,N_9132);
nand U12242 (N_12242,N_7989,N_9783);
or U12243 (N_12243,N_8443,N_8411);
nand U12244 (N_12244,N_11096,N_7435);
and U12245 (N_12245,N_9573,N_6245);
or U12246 (N_12246,N_6885,N_6145);
nand U12247 (N_12247,N_9897,N_8082);
or U12248 (N_12248,N_8326,N_10305);
and U12249 (N_12249,N_11968,N_10564);
or U12250 (N_12250,N_7848,N_7291);
and U12251 (N_12251,N_11460,N_6380);
and U12252 (N_12252,N_10822,N_7051);
and U12253 (N_12253,N_10557,N_8730);
xor U12254 (N_12254,N_8649,N_7314);
or U12255 (N_12255,N_11414,N_10276);
nor U12256 (N_12256,N_8138,N_7243);
nand U12257 (N_12257,N_8676,N_8183);
or U12258 (N_12258,N_11854,N_11226);
nand U12259 (N_12259,N_11195,N_8554);
or U12260 (N_12260,N_9864,N_11807);
or U12261 (N_12261,N_6634,N_8481);
and U12262 (N_12262,N_8329,N_7525);
nor U12263 (N_12263,N_11775,N_11522);
or U12264 (N_12264,N_8235,N_10599);
xnor U12265 (N_12265,N_10578,N_8041);
or U12266 (N_12266,N_7925,N_9086);
or U12267 (N_12267,N_11716,N_8881);
and U12268 (N_12268,N_7192,N_9154);
or U12269 (N_12269,N_11748,N_11478);
nor U12270 (N_12270,N_11502,N_10912);
xnor U12271 (N_12271,N_11077,N_9133);
xnor U12272 (N_12272,N_11264,N_7945);
nor U12273 (N_12273,N_7593,N_8739);
nor U12274 (N_12274,N_8221,N_8828);
nand U12275 (N_12275,N_10374,N_10144);
and U12276 (N_12276,N_9277,N_7732);
nand U12277 (N_12277,N_9565,N_10742);
nand U12278 (N_12278,N_11137,N_9451);
or U12279 (N_12279,N_7755,N_11518);
nor U12280 (N_12280,N_11007,N_6110);
and U12281 (N_12281,N_7107,N_8821);
nor U12282 (N_12282,N_8835,N_10318);
xor U12283 (N_12283,N_11129,N_6111);
nand U12284 (N_12284,N_8076,N_6458);
nand U12285 (N_12285,N_7327,N_6642);
or U12286 (N_12286,N_10808,N_9913);
nor U12287 (N_12287,N_7703,N_9224);
or U12288 (N_12288,N_11113,N_7961);
xnor U12289 (N_12289,N_6923,N_11410);
nand U12290 (N_12290,N_9555,N_6915);
nand U12291 (N_12291,N_6703,N_6173);
nor U12292 (N_12292,N_10961,N_6977);
xnor U12293 (N_12293,N_10561,N_10172);
or U12294 (N_12294,N_10463,N_11123);
and U12295 (N_12295,N_9584,N_8213);
nor U12296 (N_12296,N_9178,N_7552);
nor U12297 (N_12297,N_6903,N_10401);
or U12298 (N_12298,N_7346,N_10164);
nand U12299 (N_12299,N_10904,N_9229);
nand U12300 (N_12300,N_6050,N_11749);
nor U12301 (N_12301,N_11359,N_7078);
nor U12302 (N_12302,N_10563,N_8112);
nand U12303 (N_12303,N_7310,N_11128);
or U12304 (N_12304,N_7198,N_10573);
or U12305 (N_12305,N_7488,N_8712);
nor U12306 (N_12306,N_7194,N_11594);
nand U12307 (N_12307,N_11764,N_10241);
or U12308 (N_12308,N_11759,N_11040);
and U12309 (N_12309,N_8237,N_9014);
nand U12310 (N_12310,N_8327,N_8921);
xor U12311 (N_12311,N_8609,N_8714);
nand U12312 (N_12312,N_11030,N_11898);
and U12313 (N_12313,N_8683,N_9174);
xor U12314 (N_12314,N_10190,N_10674);
or U12315 (N_12315,N_6441,N_6041);
nand U12316 (N_12316,N_11217,N_6539);
and U12317 (N_12317,N_6021,N_11405);
or U12318 (N_12318,N_9795,N_7819);
nand U12319 (N_12319,N_7603,N_10391);
xnor U12320 (N_12320,N_7658,N_9832);
and U12321 (N_12321,N_7101,N_11284);
nand U12322 (N_12322,N_10938,N_11525);
xor U12323 (N_12323,N_10333,N_8360);
and U12324 (N_12324,N_11494,N_9898);
xor U12325 (N_12325,N_7464,N_9592);
and U12326 (N_12326,N_10926,N_6610);
and U12327 (N_12327,N_11001,N_7145);
nand U12328 (N_12328,N_8962,N_8684);
xor U12329 (N_12329,N_7389,N_9056);
nor U12330 (N_12330,N_9789,N_7710);
or U12331 (N_12331,N_11204,N_10795);
and U12332 (N_12332,N_9714,N_7972);
nand U12333 (N_12333,N_10460,N_8674);
nand U12334 (N_12334,N_6602,N_9233);
xor U12335 (N_12335,N_8040,N_7896);
nand U12336 (N_12336,N_6343,N_10544);
and U12337 (N_12337,N_9379,N_11523);
xor U12338 (N_12338,N_8267,N_7734);
xnor U12339 (N_12339,N_9027,N_9103);
and U12340 (N_12340,N_7568,N_10386);
or U12341 (N_12341,N_9531,N_6681);
or U12342 (N_12342,N_8064,N_9092);
and U12343 (N_12343,N_11273,N_10219);
or U12344 (N_12344,N_10491,N_11322);
or U12345 (N_12345,N_9005,N_11639);
nor U12346 (N_12346,N_9318,N_8707);
or U12347 (N_12347,N_9385,N_9442);
or U12348 (N_12348,N_8617,N_10420);
nand U12349 (N_12349,N_10028,N_8891);
or U12350 (N_12350,N_10216,N_6460);
nand U12351 (N_12351,N_11467,N_11728);
xor U12352 (N_12352,N_10047,N_11690);
nand U12353 (N_12353,N_6027,N_11052);
nand U12354 (N_12354,N_6736,N_7253);
or U12355 (N_12355,N_10415,N_9781);
or U12356 (N_12356,N_11401,N_11758);
or U12357 (N_12357,N_11832,N_10866);
xor U12358 (N_12358,N_9365,N_7025);
or U12359 (N_12359,N_8657,N_6448);
or U12360 (N_12360,N_9307,N_10087);
or U12361 (N_12361,N_10247,N_8877);
and U12362 (N_12362,N_7641,N_9167);
or U12363 (N_12363,N_6777,N_6948);
nor U12364 (N_12364,N_9182,N_11044);
xnor U12365 (N_12365,N_10598,N_9308);
nor U12366 (N_12366,N_8843,N_10382);
nand U12367 (N_12367,N_8620,N_6306);
and U12368 (N_12368,N_10361,N_7884);
and U12369 (N_12369,N_11382,N_7342);
and U12370 (N_12370,N_9498,N_7269);
xnor U12371 (N_12371,N_6038,N_6762);
or U12372 (N_12372,N_6198,N_8762);
nand U12373 (N_12373,N_10992,N_9244);
nor U12374 (N_12374,N_6790,N_9162);
nand U12375 (N_12375,N_10476,N_6649);
or U12376 (N_12376,N_8037,N_8424);
nor U12377 (N_12377,N_7062,N_9079);
nor U12378 (N_12378,N_10586,N_8229);
or U12379 (N_12379,N_6303,N_7663);
or U12380 (N_12380,N_10641,N_6676);
nand U12381 (N_12381,N_8312,N_7528);
and U12382 (N_12382,N_8189,N_11809);
nand U12383 (N_12383,N_11425,N_10312);
and U12384 (N_12384,N_11651,N_8574);
nand U12385 (N_12385,N_6959,N_7072);
xnor U12386 (N_12386,N_8177,N_11330);
nand U12387 (N_12387,N_10033,N_11360);
xnor U12388 (N_12388,N_8994,N_11991);
and U12389 (N_12389,N_6354,N_10451);
or U12390 (N_12390,N_9591,N_6105);
or U12391 (N_12391,N_8556,N_11855);
nand U12392 (N_12392,N_7099,N_6986);
and U12393 (N_12393,N_11162,N_6237);
nor U12394 (N_12394,N_6540,N_6692);
nand U12395 (N_12395,N_7150,N_7377);
xor U12396 (N_12396,N_7395,N_9124);
and U12397 (N_12397,N_6680,N_6508);
nand U12398 (N_12398,N_11097,N_9615);
and U12399 (N_12399,N_6672,N_10836);
nor U12400 (N_12400,N_10354,N_9170);
xnor U12401 (N_12401,N_6926,N_9633);
xor U12402 (N_12402,N_9099,N_9952);
nand U12403 (N_12403,N_7118,N_8970);
or U12404 (N_12404,N_10037,N_8357);
nor U12405 (N_12405,N_6694,N_10900);
nor U12406 (N_12406,N_10273,N_7262);
xor U12407 (N_12407,N_8084,N_8032);
nor U12408 (N_12408,N_11827,N_10583);
or U12409 (N_12409,N_6816,N_7448);
or U12410 (N_12410,N_6752,N_6262);
nor U12411 (N_12411,N_8810,N_11877);
nand U12412 (N_12412,N_9323,N_10840);
xnor U12413 (N_12413,N_11830,N_7178);
nand U12414 (N_12414,N_10634,N_7533);
xnor U12415 (N_12415,N_11505,N_8153);
xnor U12416 (N_12416,N_6079,N_6178);
and U12417 (N_12417,N_10221,N_11784);
and U12418 (N_12418,N_8965,N_9331);
xor U12419 (N_12419,N_8898,N_8966);
and U12420 (N_12420,N_7279,N_6846);
nor U12421 (N_12421,N_6774,N_10414);
and U12422 (N_12422,N_6025,N_11598);
and U12423 (N_12423,N_10103,N_11938);
or U12424 (N_12424,N_11634,N_10071);
and U12425 (N_12425,N_9647,N_8380);
nor U12426 (N_12426,N_6239,N_9724);
and U12427 (N_12427,N_8586,N_9411);
nor U12428 (N_12428,N_7599,N_7977);
nand U12429 (N_12429,N_6697,N_9241);
and U12430 (N_12430,N_6367,N_11899);
xor U12431 (N_12431,N_7632,N_8778);
nor U12432 (N_12432,N_8850,N_9650);
xnor U12433 (N_12433,N_6490,N_8520);
and U12434 (N_12434,N_8887,N_6608);
nand U12435 (N_12435,N_8621,N_9095);
and U12436 (N_12436,N_8280,N_9653);
and U12437 (N_12437,N_9976,N_7614);
or U12438 (N_12438,N_11713,N_8039);
nor U12439 (N_12439,N_11424,N_9807);
or U12440 (N_12440,N_11358,N_7356);
nor U12441 (N_12441,N_6981,N_11047);
or U12442 (N_12442,N_9619,N_6026);
xnor U12443 (N_12443,N_8746,N_9877);
xnor U12444 (N_12444,N_9502,N_10016);
or U12445 (N_12445,N_7134,N_7359);
nor U12446 (N_12446,N_7102,N_11702);
nor U12447 (N_12447,N_6264,N_6383);
xor U12448 (N_12448,N_7594,N_11248);
and U12449 (N_12449,N_11530,N_6080);
or U12450 (N_12450,N_7218,N_6204);
xor U12451 (N_12451,N_10289,N_10088);
or U12452 (N_12452,N_6406,N_7208);
xor U12453 (N_12453,N_7675,N_8462);
or U12454 (N_12454,N_11420,N_10399);
xor U12455 (N_12455,N_7274,N_8646);
or U12456 (N_12456,N_11836,N_7207);
and U12457 (N_12457,N_9966,N_10622);
nor U12458 (N_12458,N_9285,N_10452);
and U12459 (N_12459,N_11274,N_7979);
nor U12460 (N_12460,N_8888,N_9944);
or U12461 (N_12461,N_10271,N_10208);
nor U12462 (N_12462,N_6832,N_10477);
nand U12463 (N_12463,N_7551,N_6272);
nand U12464 (N_12464,N_6537,N_8100);
nor U12465 (N_12465,N_7693,N_11543);
and U12466 (N_12466,N_9999,N_7863);
xor U12467 (N_12467,N_6429,N_11814);
nor U12468 (N_12468,N_6718,N_10657);
or U12469 (N_12469,N_10402,N_9226);
and U12470 (N_12470,N_8906,N_9097);
and U12471 (N_12471,N_6496,N_7596);
xor U12472 (N_12472,N_8299,N_10355);
and U12473 (N_12473,N_7250,N_9472);
and U12474 (N_12474,N_7927,N_7517);
and U12475 (N_12475,N_8014,N_10350);
xnor U12476 (N_12476,N_9289,N_7298);
or U12477 (N_12477,N_10531,N_6872);
nand U12478 (N_12478,N_7137,N_11495);
or U12479 (N_12479,N_6645,N_8704);
nor U12480 (N_12480,N_8439,N_10647);
xnor U12481 (N_12481,N_10036,N_6342);
nor U12482 (N_12482,N_6186,N_7656);
and U12483 (N_12483,N_7196,N_9538);
nand U12484 (N_12484,N_9184,N_9672);
or U12485 (N_12485,N_8292,N_6092);
and U12486 (N_12486,N_11100,N_10724);
nand U12487 (N_12487,N_11158,N_9754);
nand U12488 (N_12488,N_8979,N_6039);
xor U12489 (N_12489,N_8754,N_6163);
xor U12490 (N_12490,N_7852,N_7644);
or U12491 (N_12491,N_8118,N_10061);
xor U12492 (N_12492,N_7339,N_6557);
nand U12493 (N_12493,N_7271,N_8579);
nand U12494 (N_12494,N_9423,N_9928);
nor U12495 (N_12495,N_8314,N_8832);
nand U12496 (N_12496,N_8027,N_8951);
xnor U12497 (N_12497,N_8242,N_11251);
nor U12498 (N_12498,N_9080,N_7128);
and U12499 (N_12499,N_6453,N_11999);
and U12500 (N_12500,N_6515,N_10291);
and U12501 (N_12501,N_9480,N_7918);
nor U12502 (N_12502,N_9286,N_6786);
nor U12503 (N_12503,N_10096,N_7524);
xnor U12504 (N_12504,N_11815,N_6285);
or U12505 (N_12505,N_8220,N_9535);
nor U12506 (N_12506,N_8159,N_7501);
and U12507 (N_12507,N_8974,N_7299);
and U12508 (N_12508,N_10228,N_7789);
nor U12509 (N_12509,N_11189,N_6241);
nor U12510 (N_12510,N_9335,N_7212);
nor U12511 (N_12511,N_6136,N_7365);
or U12512 (N_12512,N_11125,N_9396);
and U12513 (N_12513,N_6538,N_7168);
xor U12514 (N_12514,N_8288,N_10492);
and U12515 (N_12515,N_7795,N_7100);
xor U12516 (N_12516,N_10246,N_9831);
or U12517 (N_12517,N_9298,N_10529);
and U12518 (N_12518,N_7402,N_6391);
or U12519 (N_12519,N_8907,N_11579);
or U12520 (N_12520,N_10195,N_7006);
xor U12521 (N_12521,N_9631,N_11174);
and U12522 (N_12522,N_8308,N_11656);
or U12523 (N_12523,N_6781,N_10515);
nor U12524 (N_12524,N_6864,N_9791);
xnor U12525 (N_12525,N_9853,N_10383);
or U12526 (N_12526,N_10965,N_10043);
or U12527 (N_12527,N_8364,N_7622);
nor U12528 (N_12528,N_8142,N_9405);
and U12529 (N_12529,N_9245,N_9122);
nand U12530 (N_12530,N_11079,N_9545);
nand U12531 (N_12531,N_7705,N_9324);
or U12532 (N_12532,N_6160,N_6950);
nor U12533 (N_12533,N_7297,N_8894);
or U12534 (N_12534,N_8931,N_8913);
nor U12535 (N_12535,N_10484,N_9607);
or U12536 (N_12536,N_7073,N_6583);
xnor U12537 (N_12537,N_10789,N_9599);
xnor U12538 (N_12538,N_7222,N_7532);
and U12539 (N_12539,N_6666,N_8612);
or U12540 (N_12540,N_9749,N_8251);
or U12541 (N_12541,N_11517,N_8414);
nor U12542 (N_12542,N_11147,N_10054);
nand U12543 (N_12543,N_10118,N_11400);
nand U12544 (N_12544,N_10663,N_7067);
nand U12545 (N_12545,N_8797,N_9930);
nand U12546 (N_12546,N_10658,N_9151);
or U12547 (N_12547,N_10626,N_8926);
nor U12548 (N_12548,N_8228,N_10117);
nand U12549 (N_12549,N_8097,N_7733);
nand U12550 (N_12550,N_11948,N_7468);
xnor U12551 (N_12551,N_11327,N_8537);
nand U12552 (N_12552,N_11002,N_8343);
nor U12553 (N_12553,N_11377,N_7258);
nor U12554 (N_12554,N_9367,N_8760);
nor U12555 (N_12555,N_9948,N_7881);
or U12556 (N_12556,N_6492,N_10213);
nand U12557 (N_12557,N_10163,N_7870);
nor U12558 (N_12558,N_8858,N_9508);
nand U12559 (N_12559,N_6229,N_7129);
nor U12560 (N_12560,N_7633,N_9360);
nand U12561 (N_12561,N_6924,N_10729);
or U12562 (N_12562,N_11055,N_11239);
and U12563 (N_12563,N_7003,N_8349);
nor U12564 (N_12564,N_8491,N_10400);
xor U12565 (N_12565,N_11244,N_9895);
nor U12566 (N_12566,N_6556,N_11095);
or U12567 (N_12567,N_7023,N_11753);
nand U12568 (N_12568,N_8370,N_8875);
nand U12569 (N_12569,N_7017,N_9397);
nand U12570 (N_12570,N_10738,N_8710);
or U12571 (N_12571,N_9867,N_11145);
nor U12572 (N_12572,N_10692,N_11626);
nand U12573 (N_12573,N_8738,N_11972);
nor U12574 (N_12574,N_6077,N_7473);
nand U12575 (N_12575,N_9901,N_9275);
nor U12576 (N_12576,N_10412,N_6520);
nand U12577 (N_12577,N_10908,N_9243);
and U12578 (N_12578,N_8307,N_11364);
xnor U12579 (N_12579,N_7289,N_7320);
nor U12580 (N_12580,N_8376,N_10104);
nand U12581 (N_12581,N_8466,N_8134);
xnor U12582 (N_12582,N_6421,N_7595);
xor U12583 (N_12583,N_11298,N_11556);
nor U12584 (N_12584,N_10804,N_7579);
or U12585 (N_12585,N_6531,N_10124);
xnor U12586 (N_12586,N_7787,N_11864);
and U12587 (N_12587,N_7728,N_11920);
and U12588 (N_12588,N_11465,N_8987);
xnor U12589 (N_12589,N_10495,N_9847);
and U12590 (N_12590,N_9932,N_11199);
xnor U12591 (N_12591,N_9117,N_11352);
and U12592 (N_12592,N_11101,N_11813);
nand U12593 (N_12593,N_10292,N_8320);
xnor U12594 (N_12594,N_11873,N_10898);
xnor U12595 (N_12595,N_6408,N_6839);
and U12596 (N_12596,N_10869,N_7204);
nand U12597 (N_12597,N_7992,N_7348);
or U12598 (N_12598,N_6821,N_11778);
or U12599 (N_12599,N_6730,N_6106);
nor U12600 (N_12600,N_7360,N_8792);
or U12601 (N_12601,N_7246,N_9141);
nor U12602 (N_12602,N_9851,N_7456);
xor U12603 (N_12603,N_10097,N_9785);
xor U12604 (N_12604,N_6661,N_9388);
and U12605 (N_12605,N_10302,N_11837);
xnor U12606 (N_12606,N_6290,N_6479);
or U12607 (N_12607,N_9939,N_9804);
nand U12608 (N_12608,N_6255,N_8950);
and U12609 (N_12609,N_10095,N_8772);
nand U12610 (N_12610,N_7077,N_8233);
nand U12611 (N_12611,N_8381,N_10007);
xnor U12612 (N_12612,N_11335,N_9759);
xnor U12613 (N_12613,N_8383,N_9390);
nor U12614 (N_12614,N_9046,N_6260);
nor U12615 (N_12615,N_8615,N_7778);
nor U12616 (N_12616,N_11568,N_11108);
or U12617 (N_12617,N_6197,N_6347);
nand U12618 (N_12618,N_6096,N_9959);
and U12619 (N_12619,N_10205,N_7322);
nor U12620 (N_12620,N_6362,N_11802);
xor U12621 (N_12621,N_9914,N_8086);
xor U12622 (N_12622,N_9891,N_7761);
xnor U12623 (N_12623,N_10769,N_8743);
or U12624 (N_12624,N_10752,N_8154);
and U12625 (N_12625,N_7954,N_10379);
nand U12626 (N_12626,N_8990,N_11681);
nor U12627 (N_12627,N_9641,N_11875);
and U12628 (N_12628,N_7362,N_11735);
or U12629 (N_12629,N_9656,N_6930);
xnor U12630 (N_12630,N_6472,N_10859);
and U12631 (N_12631,N_9648,N_10381);
xnor U12632 (N_12632,N_9697,N_11737);
or U12633 (N_12633,N_11990,N_8063);
xor U12634 (N_12634,N_8971,N_11236);
and U12635 (N_12635,N_8544,N_9580);
xor U12636 (N_12636,N_7056,N_10048);
or U12637 (N_12637,N_6543,N_11472);
or U12638 (N_12638,N_6308,N_8663);
nand U12639 (N_12639,N_8587,N_8666);
xor U12640 (N_12640,N_7542,N_6012);
nor U12641 (N_12641,N_7776,N_7561);
xnor U12642 (N_12642,N_10042,N_9258);
and U12643 (N_12643,N_6918,N_7964);
nor U12644 (N_12644,N_11888,N_8318);
or U12645 (N_12645,N_8293,N_6210);
or U12646 (N_12646,N_8149,N_8243);
or U12647 (N_12647,N_6022,N_10417);
or U12648 (N_12648,N_7496,N_6368);
or U12649 (N_12649,N_7510,N_8169);
nand U12650 (N_12650,N_10678,N_6242);
xnor U12651 (N_12651,N_7393,N_8029);
or U12652 (N_12652,N_7287,N_8048);
nand U12653 (N_12653,N_11527,N_9625);
nor U12654 (N_12654,N_11391,N_6588);
xor U12655 (N_12655,N_7479,N_8981);
nand U12656 (N_12656,N_11648,N_9435);
or U12657 (N_12657,N_8108,N_6234);
nor U12658 (N_12658,N_10750,N_6646);
xnor U12659 (N_12659,N_9674,N_9371);
nor U12660 (N_12660,N_8447,N_7920);
or U12661 (N_12661,N_9602,N_10762);
nand U12662 (N_12662,N_9675,N_10998);
xor U12663 (N_12663,N_11326,N_11463);
nor U12664 (N_12664,N_11511,N_6688);
xnor U12665 (N_12665,N_8697,N_8451);
xnor U12666 (N_12666,N_6165,N_7895);
and U12667 (N_12667,N_9376,N_10606);
and U12668 (N_12668,N_9179,N_7788);
nor U12669 (N_12669,N_10576,N_8928);
nand U12670 (N_12670,N_7164,N_6257);
nor U12671 (N_12671,N_11323,N_6401);
nand U12672 (N_12672,N_10498,N_9257);
nand U12673 (N_12673,N_7904,N_10911);
and U12674 (N_12674,N_6750,N_9317);
or U12675 (N_12675,N_7546,N_10109);
xnor U12676 (N_12676,N_8016,N_9292);
xnor U12677 (N_12677,N_8338,N_7689);
or U12678 (N_12678,N_11526,N_7300);
nor U12679 (N_12679,N_6216,N_8204);
nor U12680 (N_12680,N_6900,N_8661);
nor U12681 (N_12681,N_8626,N_11389);
nor U12682 (N_12682,N_8934,N_9666);
nor U12683 (N_12683,N_10555,N_11538);
and U12684 (N_12684,N_8405,N_8841);
nor U12685 (N_12685,N_8955,N_8150);
or U12686 (N_12686,N_7281,N_8470);
xnor U12687 (N_12687,N_10614,N_7492);
xnor U12688 (N_12688,N_7955,N_7195);
and U12689 (N_12689,N_6994,N_7133);
nand U12690 (N_12690,N_11039,N_7193);
xnor U12691 (N_12691,N_10506,N_10227);
xor U12692 (N_12692,N_8087,N_9761);
nor U12693 (N_12693,N_7309,N_6785);
nand U12694 (N_12694,N_7792,N_6512);
xnor U12695 (N_12695,N_9313,N_9551);
xnor U12696 (N_12696,N_9497,N_6933);
and U12697 (N_12697,N_10306,N_9302);
nor U12698 (N_12698,N_7406,N_10099);
and U12699 (N_12699,N_6265,N_9171);
or U12700 (N_12700,N_9682,N_10875);
nor U12701 (N_12701,N_6913,N_8456);
nor U12702 (N_12702,N_8069,N_9936);
nor U12703 (N_12703,N_6570,N_11691);
or U12704 (N_12704,N_8512,N_11411);
nor U12705 (N_12705,N_10723,N_8935);
nand U12706 (N_12706,N_6201,N_11602);
nand U12707 (N_12707,N_11092,N_6803);
xor U12708 (N_12708,N_9552,N_11295);
or U12709 (N_12709,N_11266,N_8129);
nand U12710 (N_12710,N_7877,N_11859);
nor U12711 (N_12711,N_6576,N_8773);
nand U12712 (N_12712,N_9890,N_7793);
and U12713 (N_12713,N_9392,N_10983);
or U12714 (N_12714,N_8354,N_11041);
nor U12715 (N_12715,N_6118,N_8919);
nand U12716 (N_12716,N_10737,N_10874);
or U12717 (N_12717,N_7481,N_7477);
and U12718 (N_12718,N_9111,N_9283);
or U12719 (N_12719,N_11600,N_10538);
or U12720 (N_12720,N_11671,N_8884);
nor U12721 (N_12721,N_6117,N_7624);
nor U12722 (N_12722,N_8952,N_7968);
nand U12723 (N_12723,N_11934,N_7687);
or U12724 (N_12724,N_6794,N_7763);
or U12725 (N_12725,N_6461,N_7304);
nand U12726 (N_12726,N_6897,N_10605);
nand U12727 (N_12727,N_7414,N_10800);
nand U12728 (N_12728,N_9569,N_10725);
or U12729 (N_12729,N_11259,N_8805);
or U12730 (N_12730,N_8395,N_8834);
nand U12731 (N_12731,N_9422,N_11780);
nor U12732 (N_12732,N_8664,N_10334);
nand U12733 (N_12733,N_10980,N_10664);
nand U12734 (N_12734,N_10159,N_11941);
and U12735 (N_12735,N_8737,N_10323);
and U12736 (N_12736,N_8253,N_9986);
or U12737 (N_12737,N_6153,N_9089);
nor U12738 (N_12738,N_7172,N_10089);
or U12739 (N_12739,N_7167,N_10131);
and U12740 (N_12740,N_7673,N_9398);
or U12741 (N_12741,N_11608,N_10607);
nand U12742 (N_12742,N_11619,N_6764);
or U12743 (N_12743,N_7387,N_7388);
nand U12744 (N_12744,N_6584,N_10870);
and U12745 (N_12745,N_11514,N_7609);
nand U12746 (N_12746,N_6970,N_11084);
nand U12747 (N_12747,N_7521,N_7505);
and U12748 (N_12748,N_7620,N_7943);
nor U12749 (N_12749,N_6742,N_8782);
xnor U12750 (N_12750,N_10771,N_7838);
and U12751 (N_12751,N_9322,N_11160);
xor U12752 (N_12752,N_11114,N_6400);
xor U12753 (N_12753,N_9709,N_11140);
nand U12754 (N_12754,N_8494,N_7519);
nor U12755 (N_12755,N_11618,N_10066);
and U12756 (N_12756,N_11757,N_6085);
and U12757 (N_12757,N_10915,N_9902);
and U12758 (N_12758,N_6253,N_9955);
or U12759 (N_12759,N_10810,N_8441);
nor U12760 (N_12760,N_7200,N_8254);
xnor U12761 (N_12761,N_11304,N_9486);
and U12762 (N_12762,N_8382,N_8623);
nor U12763 (N_12763,N_9949,N_6350);
or U12764 (N_12764,N_8050,N_6831);
nand U12765 (N_12765,N_11297,N_10486);
xor U12766 (N_12766,N_9920,N_7803);
nor U12767 (N_12767,N_11170,N_11957);
xnor U12768 (N_12768,N_7498,N_11826);
nor U12769 (N_12769,N_6908,N_6511);
or U12770 (N_12770,N_9984,N_7185);
or U12771 (N_12771,N_6295,N_11643);
nor U12772 (N_12772,N_11255,N_10435);
or U12773 (N_12773,N_11886,N_11670);
xor U12774 (N_12774,N_9951,N_11820);
nor U12775 (N_12775,N_8501,N_8123);
nor U12776 (N_12776,N_8473,N_7857);
and U12777 (N_12777,N_9344,N_10327);
nand U12778 (N_12778,N_7127,N_11944);
nor U12779 (N_12779,N_9039,N_8721);
nand U12780 (N_12780,N_8377,N_9915);
nand U12781 (N_12781,N_10006,N_9972);
or U12782 (N_12782,N_10682,N_11422);
xnor U12783 (N_12783,N_10895,N_8895);
nand U12784 (N_12784,N_11353,N_6425);
nand U12785 (N_12785,N_11895,N_9537);
nand U12786 (N_12786,N_8306,N_11590);
nor U12787 (N_12787,N_7242,N_9048);
nor U12788 (N_12788,N_6518,N_8933);
and U12789 (N_12789,N_8600,N_6323);
nor U12790 (N_12790,N_7942,N_8294);
xnor U12791 (N_12791,N_7205,N_7465);
xnor U12792 (N_12792,N_8690,N_6603);
and U12793 (N_12793,N_9995,N_10413);
or U12794 (N_12794,N_7854,N_11925);
or U12795 (N_12795,N_7063,N_8499);
and U12796 (N_12796,N_9063,N_6731);
or U12797 (N_12797,N_8961,N_9561);
and U12798 (N_12798,N_11874,N_8347);
nand U12799 (N_12799,N_6856,N_7112);
nand U12800 (N_12800,N_11896,N_9345);
nand U12801 (N_12801,N_6572,N_9764);
and U12802 (N_12802,N_8102,N_10021);
nor U12803 (N_12803,N_8417,N_6600);
nor U12804 (N_12804,N_8319,N_11333);
nor U12805 (N_12805,N_10986,N_8899);
xnor U12806 (N_12806,N_9329,N_11346);
nor U12807 (N_12807,N_11455,N_11705);
nor U12808 (N_12808,N_9616,N_10193);
nor U12809 (N_12809,N_11105,N_7842);
or U12810 (N_12810,N_11117,N_8392);
or U12811 (N_12811,N_9691,N_7093);
nor U12812 (N_12812,N_7431,N_7000);
nand U12813 (N_12813,N_7699,N_6656);
or U12814 (N_12814,N_11881,N_10079);
and U12815 (N_12815,N_10828,N_8388);
nor U12816 (N_12816,N_7627,N_11890);
and U12817 (N_12817,N_10285,N_8304);
and U12818 (N_12818,N_8669,N_9267);
and U12819 (N_12819,N_7450,N_9703);
xor U12820 (N_12820,N_11587,N_7221);
nand U12821 (N_12821,N_6953,N_11439);
or U12822 (N_12822,N_7080,N_9078);
and U12823 (N_12823,N_6863,N_9515);
nand U12824 (N_12824,N_9563,N_8366);
and U12825 (N_12825,N_6858,N_11557);
or U12826 (N_12826,N_8529,N_6637);
and U12827 (N_12827,N_9250,N_7543);
nor U12828 (N_12828,N_8985,N_11994);
or U12829 (N_12829,N_11646,N_6622);
nand U12830 (N_12830,N_11131,N_9518);
nand U12831 (N_12831,N_11269,N_11214);
nand U12832 (N_12832,N_10942,N_10566);
or U12833 (N_12833,N_8065,N_11104);
xor U12834 (N_12834,N_6161,N_7153);
or U12835 (N_12835,N_11788,N_6138);
xor U12836 (N_12836,N_6417,N_8713);
or U12837 (N_12837,N_8656,N_6632);
nand U12838 (N_12838,N_7771,N_11965);
and U12839 (N_12839,N_9389,N_6259);
or U12840 (N_12840,N_9312,N_11122);
or U12841 (N_12841,N_8495,N_6965);
or U12842 (N_12842,N_8226,N_6619);
nor U12843 (N_12843,N_11013,N_8723);
nand U12844 (N_12844,N_7650,N_6008);
and U12845 (N_12845,N_6439,N_8871);
xor U12846 (N_12846,N_7216,N_6058);
and U12847 (N_12847,N_10086,N_6481);
or U12848 (N_12848,N_6219,N_7382);
or U12849 (N_12849,N_10940,N_10137);
nand U12850 (N_12850,N_7236,N_8725);
and U12851 (N_12851,N_7631,N_9087);
nor U12852 (N_12852,N_6139,N_11986);
and U12853 (N_12853,N_8652,N_8557);
and U12854 (N_12854,N_10040,N_8796);
xnor U12855 (N_12855,N_9121,N_10787);
and U12856 (N_12856,N_10045,N_8604);
or U12857 (N_12857,N_11761,N_11479);
nand U12858 (N_12858,N_10821,N_11254);
or U12859 (N_12859,N_10730,N_11916);
nand U12860 (N_12860,N_9000,N_9413);
nor U12861 (N_12861,N_9372,N_11605);
and U12862 (N_12862,N_6733,N_7919);
and U12863 (N_12863,N_7058,N_10150);
nor U12864 (N_12864,N_11768,N_8091);
and U12865 (N_12865,N_8840,N_7610);
nor U12866 (N_12866,N_10584,N_8498);
xor U12867 (N_12867,N_7374,N_8418);
and U12868 (N_12868,N_8264,N_8983);
nand U12869 (N_12869,N_10958,N_11406);
and U12870 (N_12870,N_6905,N_8519);
nand U12871 (N_12871,N_8896,N_11000);
and U12872 (N_12872,N_7223,N_9213);
xnor U12873 (N_12873,N_11238,N_8627);
xnor U12874 (N_12874,N_6782,N_10231);
or U12875 (N_12875,N_8230,N_8185);
nor U12876 (N_12876,N_11937,N_9722);
and U12877 (N_12877,N_11144,N_7985);
and U12878 (N_12878,N_6580,N_9852);
nand U12879 (N_12879,N_9457,N_10480);
or U12880 (N_12880,N_11580,N_6721);
nor U12881 (N_12881,N_6702,N_10180);
nand U12882 (N_12882,N_10268,N_9077);
nor U12883 (N_12883,N_8550,N_9051);
xor U12884 (N_12884,N_11564,N_11378);
or U12885 (N_12885,N_9358,N_10183);
or U12886 (N_12886,N_8208,N_9907);
or U12887 (N_12887,N_8504,N_8043);
and U12888 (N_12888,N_11005,N_11477);
and U12889 (N_12889,N_8964,N_10610);
xnor U12890 (N_12890,N_8505,N_10739);
nand U12891 (N_12891,N_11541,N_8764);
or U12892 (N_12892,N_9989,N_8433);
nor U12893 (N_12893,N_9485,N_9052);
or U12894 (N_12894,N_6107,N_6476);
nand U12895 (N_12895,N_11617,N_11283);
and U12896 (N_12896,N_6387,N_9784);
and U12897 (N_12897,N_10431,N_10715);
nor U12898 (N_12898,N_7830,N_11230);
nand U12899 (N_12899,N_10572,N_9975);
nand U12900 (N_12900,N_6162,N_8436);
and U12901 (N_12901,N_8194,N_11018);
nor U12902 (N_12902,N_10830,N_11009);
or U12903 (N_12903,N_10823,N_11829);
nor U12904 (N_12904,N_8527,N_10909);
or U12905 (N_12905,N_7106,N_7998);
xnor U12906 (N_12906,N_9980,N_9904);
xnor U12907 (N_12907,N_11819,N_10754);
and U12908 (N_12908,N_7081,N_7729);
or U12909 (N_12909,N_6620,N_9738);
nor U12910 (N_12910,N_11701,N_8140);
nand U12911 (N_12911,N_8143,N_10278);
and U12912 (N_12912,N_11911,N_10956);
or U12913 (N_12913,N_7592,N_7823);
and U12914 (N_12914,N_8453,N_9387);
and U12915 (N_12915,N_8248,N_10168);
xor U12916 (N_12916,N_11370,N_10782);
and U12917 (N_12917,N_9339,N_6604);
and U12918 (N_12918,N_10793,N_6098);
or U12919 (N_12919,N_7461,N_8541);
xnor U12920 (N_12920,N_6826,N_7441);
and U12921 (N_12921,N_8196,N_11155);
xor U12922 (N_12922,N_10304,N_11376);
nor U12923 (N_12923,N_10562,N_10632);
and U12924 (N_12924,N_6533,N_6711);
xor U12925 (N_12925,N_11747,N_9031);
nor U12926 (N_12926,N_8659,N_9828);
nor U12927 (N_12927,N_8651,N_6132);
and U12928 (N_12928,N_6633,N_9383);
or U12929 (N_12929,N_9815,N_8679);
and U12930 (N_12930,N_11193,N_11426);
or U12931 (N_12931,N_6878,N_11967);
and U12932 (N_12932,N_10122,N_10661);
nand U12933 (N_12933,N_10733,N_7691);
nor U12934 (N_12934,N_8282,N_11993);
nor U12935 (N_12935,N_10817,N_10835);
nor U12936 (N_12936,N_7442,N_9030);
xnor U12937 (N_12937,N_7454,N_10863);
and U12938 (N_12938,N_9817,N_11631);
nand U12939 (N_12939,N_6862,N_10616);
nor U12940 (N_12940,N_8271,N_9796);
and U12941 (N_12941,N_7621,N_9626);
nand U12942 (N_12942,N_10834,N_10720);
xor U12943 (N_12943,N_8589,N_9043);
xor U12944 (N_12944,N_8477,N_8117);
nor U12945 (N_12945,N_6934,N_8580);
and U12946 (N_12946,N_6477,N_8198);
or U12947 (N_12947,N_8359,N_7398);
and U12948 (N_12948,N_9042,N_7834);
and U12949 (N_12949,N_7239,N_9992);
and U12950 (N_12950,N_10136,N_6628);
or U12951 (N_12951,N_6975,N_9765);
and U12952 (N_12952,N_6788,N_11253);
nand U12953 (N_12953,N_9982,N_6185);
and U12954 (N_12954,N_9355,N_11806);
and U12955 (N_12955,N_7457,N_10806);
and U12956 (N_12956,N_6780,N_7843);
and U12957 (N_12957,N_7978,N_7589);
nor U12958 (N_12958,N_8215,N_11149);
and U12959 (N_12959,N_6855,N_11501);
nand U12960 (N_12960,N_8444,N_10995);
nand U12961 (N_12961,N_8551,N_11858);
and U12962 (N_12962,N_8948,N_9845);
nand U12963 (N_12963,N_6416,N_6267);
xnor U12964 (N_12964,N_7913,N_7762);
nor U12965 (N_12965,N_11507,N_10372);
xnor U12966 (N_12966,N_8374,N_8406);
nor U12967 (N_12967,N_11606,N_8905);
xor U12968 (N_12968,N_9443,N_7737);
or U12969 (N_12969,N_6317,N_9459);
or U12970 (N_12970,N_11071,N_10348);
xnor U12971 (N_12971,N_11050,N_6073);
nor U12972 (N_12972,N_9588,N_10960);
nand U12973 (N_12973,N_11127,N_11240);
nand U12974 (N_12974,N_10691,N_7969);
xnor U12975 (N_12975,N_10467,N_9746);
xor U12976 (N_12976,N_8633,N_7386);
and U12977 (N_12977,N_7751,N_10182);
nand U12978 (N_12978,N_7980,N_6405);
and U12979 (N_12979,N_7815,N_7660);
xnor U12980 (N_12980,N_11892,N_11786);
xnor U12981 (N_12981,N_10847,N_9349);
and U12982 (N_12982,N_11466,N_8310);
xnor U12983 (N_12983,N_9399,N_6888);
and U12984 (N_12984,N_6519,N_11192);
nand U12985 (N_12985,N_6437,N_10517);
xor U12986 (N_12986,N_9630,N_6504);
or U12987 (N_12987,N_9198,N_9054);
nand U12988 (N_12988,N_11252,N_10928);
nor U12989 (N_12989,N_9818,N_9462);
xnor U12990 (N_12990,N_11584,N_8992);
and U12991 (N_12991,N_10322,N_10187);
xor U12992 (N_12992,N_6659,N_10064);
and U12993 (N_12993,N_8463,N_8145);
xnor U12994 (N_12994,N_8234,N_7747);
nor U12995 (N_12995,N_7791,N_11825);
and U12996 (N_12996,N_7890,N_8978);
xor U12997 (N_12997,N_8636,N_9668);
nand U12998 (N_12998,N_7068,N_7731);
nor U12999 (N_12999,N_10056,N_10545);
and U13000 (N_13000,N_9827,N_9314);
and U13001 (N_13001,N_6034,N_6190);
or U13002 (N_13002,N_8923,N_6587);
nand U13003 (N_13003,N_9287,N_7061);
nor U13004 (N_13004,N_11989,N_9820);
nor U13005 (N_13005,N_6298,N_6919);
xor U13006 (N_13006,N_11187,N_9824);
xnor U13007 (N_13007,N_11306,N_6558);
nand U13008 (N_13008,N_11449,N_10317);
nor U13009 (N_13009,N_7635,N_9351);
xor U13010 (N_13010,N_9011,N_11660);
and U13011 (N_13011,N_9810,N_7502);
and U13012 (N_13012,N_11061,N_11212);
and U13013 (N_13013,N_9707,N_7799);
or U13014 (N_13014,N_11141,N_11069);
nand U13015 (N_13015,N_11142,N_11116);
and U13016 (N_13016,N_8897,N_7759);
nand U13017 (N_13017,N_9608,N_10041);
nand U13018 (N_13018,N_7715,N_11203);
and U13019 (N_13019,N_10277,N_8908);
and U13020 (N_13020,N_11235,N_11367);
or U13021 (N_13021,N_11569,N_6035);
xor U13022 (N_13022,N_10948,N_11205);
nor U13023 (N_13023,N_8837,N_11027);
and U13024 (N_13024,N_6802,N_11677);
xor U13025 (N_13025,N_10148,N_9998);
nor U13026 (N_13026,N_11270,N_7052);
nor U13027 (N_13027,N_6754,N_9455);
nor U13028 (N_13028,N_11056,N_9157);
nor U13029 (N_13029,N_8915,N_10721);
nor U13030 (N_13030,N_11225,N_7190);
xnor U13031 (N_13031,N_7783,N_9090);
nor U13032 (N_13032,N_11090,N_10199);
nand U13033 (N_13033,N_11962,N_6225);
xor U13034 (N_13034,N_10500,N_10160);
xnor U13035 (N_13035,N_6181,N_7813);
xor U13036 (N_13036,N_8525,N_8780);
xnor U13037 (N_13037,N_8728,N_8660);
xnor U13038 (N_13038,N_11134,N_6522);
xnor U13039 (N_13039,N_6971,N_8826);
or U13040 (N_13040,N_10204,N_11513);
xnor U13041 (N_13041,N_7353,N_10055);
nand U13042 (N_13042,N_6006,N_8386);
nand U13043 (N_13043,N_9679,N_8394);
xor U13044 (N_13044,N_10676,N_9942);
and U13045 (N_13045,N_9108,N_8004);
xnor U13046 (N_13046,N_8283,N_6435);
or U13047 (N_13047,N_10882,N_6452);
nand U13048 (N_13048,N_9297,N_10181);
nand U13049 (N_13049,N_9854,N_9994);
nor U13050 (N_13050,N_6678,N_8256);
xor U13051 (N_13051,N_8861,N_11924);
nor U13052 (N_13052,N_10978,N_6796);
nand U13053 (N_13053,N_8545,N_10432);
and U13054 (N_13054,N_10811,N_7059);
and U13055 (N_13055,N_10887,N_6638);
nand U13056 (N_13056,N_11228,N_7976);
and U13057 (N_13057,N_7527,N_11073);
nand U13058 (N_13058,N_8042,N_10326);
nand U13059 (N_13059,N_10528,N_10311);
and U13060 (N_13060,N_6301,N_11996);
and U13061 (N_13061,N_6164,N_9126);
or U13062 (N_13062,N_10005,N_8830);
or U13063 (N_13063,N_10772,N_8658);
and U13064 (N_13064,N_9183,N_11966);
nor U13065 (N_13065,N_7438,N_7897);
or U13066 (N_13066,N_10785,N_11698);
nand U13067 (N_13067,N_6459,N_10639);
and U13068 (N_13068,N_7820,N_8783);
nand U13069 (N_13069,N_10341,N_7923);
nand U13070 (N_13070,N_8367,N_6899);
nor U13071 (N_13071,N_8371,N_6867);
nor U13072 (N_13072,N_9263,N_9747);
nand U13073 (N_13073,N_6103,N_9927);
or U13074 (N_13074,N_8777,N_6684);
nand U13075 (N_13075,N_7698,N_6244);
or U13076 (N_13076,N_10210,N_6517);
nor U13077 (N_13077,N_7440,N_10996);
nand U13078 (N_13078,N_9160,N_11573);
and U13079 (N_13079,N_10023,N_9168);
nand U13080 (N_13080,N_10296,N_9921);
xnor U13081 (N_13081,N_11107,N_8410);
and U13082 (N_13082,N_6807,N_10642);
nor U13083 (N_13083,N_11303,N_11918);
and U13084 (N_13084,N_7363,N_6189);
xor U13085 (N_13085,N_8113,N_7822);
xor U13086 (N_13086,N_10907,N_9203);
nand U13087 (N_13087,N_7905,N_9594);
nand U13088 (N_13088,N_10706,N_7850);
and U13089 (N_13089,N_10408,N_7680);
and U13090 (N_13090,N_11200,N_6280);
and U13091 (N_13091,N_6621,N_8120);
xnor U13092 (N_13092,N_9265,N_9008);
nand U13093 (N_13093,N_11072,N_11154);
or U13094 (N_13094,N_7413,N_7494);
or U13095 (N_13095,N_9911,N_7573);
or U13096 (N_13096,N_11862,N_10186);
xnor U13097 (N_13097,N_6935,N_9192);
xnor U13098 (N_13098,N_10394,N_11696);
and U13099 (N_13099,N_6704,N_7130);
and U13100 (N_13100,N_6119,N_7812);
and U13101 (N_13101,N_9742,N_11496);
nand U13102 (N_13102,N_7432,N_8628);
nor U13103 (N_13103,N_9806,N_11637);
or U13104 (N_13104,N_9104,N_6227);
nand U13105 (N_13105,N_11396,N_9542);
xor U13106 (N_13106,N_8262,N_8668);
nand U13107 (N_13107,N_11812,N_10133);
and U13108 (N_13108,N_7123,N_6967);
and U13109 (N_13109,N_11946,N_9020);
xor U13110 (N_13110,N_6562,N_9146);
nor U13111 (N_13111,N_10236,N_9445);
nor U13112 (N_13112,N_6444,N_9088);
or U13113 (N_13113,N_10653,N_10662);
nor U13114 (N_13114,N_10194,N_10776);
and U13115 (N_13115,N_6695,N_10748);
and U13116 (N_13116,N_11529,N_9977);
nor U13117 (N_13117,N_7154,N_9954);
and U13118 (N_13118,N_8893,N_8790);
nand U13119 (N_13119,N_7184,N_11453);
nand U13120 (N_13120,N_10745,N_8325);
and U13121 (N_13121,N_7712,N_10704);
nand U13122 (N_13122,N_8009,N_9687);
and U13123 (N_13123,N_9342,N_11481);
nor U13124 (N_13124,N_8435,N_8696);
nand U13125 (N_13125,N_9846,N_10542);
nor U13126 (N_13126,N_8083,N_7772);
xor U13127 (N_13127,N_6756,N_8925);
xor U13128 (N_13128,N_7990,N_6818);
nand U13129 (N_13129,N_11649,N_6443);
nor U13130 (N_13130,N_10149,N_8476);
nand U13131 (N_13131,N_8767,N_9658);
nor U13132 (N_13132,N_9655,N_10946);
and U13133 (N_13133,N_11487,N_10746);
or U13134 (N_13134,N_10686,N_7619);
xor U13135 (N_13135,N_10854,N_6388);
nand U13136 (N_13136,N_9019,N_10371);
nand U13137 (N_13137,N_10666,N_7217);
nand U13138 (N_13138,N_11708,N_6420);
or U13139 (N_13139,N_7993,N_6617);
or U13140 (N_13140,N_7074,N_6451);
nor U13141 (N_13141,N_10446,N_8820);
nor U13142 (N_13142,N_7034,N_6344);
and U13143 (N_13143,N_9530,N_11172);
nor U13144 (N_13144,N_9888,N_6233);
or U13145 (N_13145,N_10254,N_6393);
nand U13146 (N_13146,N_11572,N_9713);
nor U13147 (N_13147,N_7583,N_9002);
nand U13148 (N_13148,N_11707,N_10541);
and U13149 (N_13149,N_11926,N_9135);
or U13150 (N_13150,N_9664,N_9044);
nor U13151 (N_13151,N_8672,N_9532);
or U13152 (N_13152,N_11810,N_6226);
nor U13153 (N_13153,N_7103,N_8798);
and U13154 (N_13154,N_6223,N_6848);
nor U13155 (N_13155,N_10051,N_11585);
and U13156 (N_13156,N_11910,N_7141);
nand U13157 (N_13157,N_9874,N_11844);
nand U13158 (N_13158,N_7426,N_9067);
xnor U13159 (N_13159,N_10035,N_6349);
or U13160 (N_13160,N_8426,N_6268);
nand U13161 (N_13161,N_9777,N_8632);
and U13162 (N_13162,N_10074,N_6094);
or U13163 (N_13163,N_6377,N_11878);
and U13164 (N_13164,N_8273,N_11325);
or U13165 (N_13165,N_10690,N_9819);
or U13166 (N_13166,N_11023,N_6076);
or U13167 (N_13167,N_9879,N_10766);
xnor U13168 (N_13168,N_6808,N_7839);
or U13169 (N_13169,N_11293,N_10239);
nand U13170 (N_13170,N_8186,N_10851);
nor U13171 (N_13171,N_6741,N_9830);
nand U13172 (N_13172,N_11229,N_7428);
nor U13173 (N_13173,N_7029,N_6252);
or U13174 (N_13174,N_9524,N_7159);
and U13175 (N_13175,N_9038,N_11578);
or U13176 (N_13176,N_8507,N_8546);
nor U13177 (N_13177,N_8249,N_10868);
and U13178 (N_13178,N_8287,N_7284);
nor U13179 (N_13179,N_8500,N_9470);
xnor U13180 (N_13180,N_9776,N_6606);
nand U13181 (N_13181,N_6751,N_9643);
or U13182 (N_13182,N_8538,N_6093);
or U13183 (N_13183,N_8214,N_7189);
nor U13184 (N_13184,N_7939,N_7182);
xnor U13185 (N_13185,N_10974,N_7769);
and U13186 (N_13186,N_10093,N_11563);
xnor U13187 (N_13187,N_7292,N_9756);
or U13188 (N_13188,N_9711,N_9654);
xnor U13189 (N_13189,N_9665,N_9071);
nor U13190 (N_13190,N_7966,N_8540);
and U13191 (N_13191,N_11015,N_10077);
and U13192 (N_13192,N_11138,N_7640);
xor U13193 (N_13193,N_11774,N_11659);
nor U13194 (N_13194,N_10604,N_10546);
or U13195 (N_13195,N_11685,N_7086);
nor U13196 (N_13196,N_6546,N_7044);
or U13197 (N_13197,N_10929,N_11970);
or U13198 (N_13198,N_6560,N_7926);
and U13199 (N_13199,N_6011,N_6532);
or U13200 (N_13200,N_9222,N_7069);
and U13201 (N_13201,N_9394,N_9953);
xnor U13202 (N_13202,N_7807,N_9842);
and U13203 (N_13203,N_9492,N_6665);
nor U13204 (N_13204,N_9598,N_10426);
xnor U13205 (N_13205,N_6129,N_11480);
nor U13206 (N_13206,N_7367,N_8533);
nand U13207 (N_13207,N_8432,N_8396);
and U13208 (N_13208,N_9195,N_6689);
nor U13209 (N_13209,N_8335,N_7165);
or U13210 (N_13210,N_11743,N_10962);
and U13211 (N_13211,N_9590,N_11003);
and U13212 (N_13212,N_6941,N_6059);
xnor U13213 (N_13213,N_7368,N_8099);
and U13214 (N_13214,N_7576,N_8625);
nand U13215 (N_13215,N_10140,N_6351);
nand U13216 (N_13216,N_8571,N_6830);
or U13217 (N_13217,N_6072,N_11719);
and U13218 (N_13218,N_11499,N_6447);
nor U13219 (N_13219,N_11773,N_8508);
and U13220 (N_13220,N_11299,N_11756);
or U13221 (N_13221,N_7958,N_8799);
xnor U13222 (N_13222,N_11434,N_9176);
or U13223 (N_13223,N_11599,N_10331);
or U13224 (N_13224,N_10328,N_11380);
nand U13225 (N_13225,N_10741,N_6099);
or U13226 (N_13226,N_7545,N_11279);
and U13227 (N_13227,N_11818,N_8553);
xor U13228 (N_13228,N_9693,N_11740);
xnor U13229 (N_13229,N_10714,N_8006);
and U13230 (N_13230,N_10613,N_6179);
xnor U13231 (N_13231,N_9391,N_11746);
or U13232 (N_13232,N_8106,N_11997);
xor U13233 (N_13233,N_10017,N_6374);
xor U13234 (N_13234,N_9429,N_10429);
nor U13235 (N_13235,N_9521,N_9947);
xnor U13236 (N_13236,N_7340,N_8867);
nor U13237 (N_13237,N_7973,N_10973);
and U13238 (N_13238,N_9507,N_10934);
or U13239 (N_13239,N_11363,N_11657);
nor U13240 (N_13240,N_7739,N_9006);
nor U13241 (N_13241,N_9434,N_11893);
or U13242 (N_13242,N_6993,N_11687);
nor U13243 (N_13243,N_10963,N_7476);
nand U13244 (N_13244,N_10300,N_11182);
or U13245 (N_13245,N_7871,N_6488);
or U13246 (N_13246,N_11868,N_9456);
and U13247 (N_13247,N_6294,N_7797);
nor U13248 (N_13248,N_6887,N_10363);
and U13249 (N_13249,N_11689,N_6837);
nand U13250 (N_13250,N_10537,N_7847);
xnor U13251 (N_13251,N_7238,N_8701);
and U13252 (N_13252,N_9330,N_9553);
xnor U13253 (N_13253,N_10876,N_6737);
nand U13254 (N_13254,N_7197,N_10468);
or U13255 (N_13255,N_8067,N_10258);
nor U13256 (N_13256,N_6352,N_6358);
nor U13257 (N_13257,N_9757,N_6363);
or U13258 (N_13258,N_11431,N_7449);
xor U13259 (N_13259,N_10553,N_9064);
nor U13260 (N_13260,N_11497,N_9912);
and U13261 (N_13261,N_10829,N_6396);
xor U13262 (N_13262,N_11738,N_9483);
xor U13263 (N_13263,N_6188,N_9116);
xnor U13264 (N_13264,N_11553,N_11959);
or U13265 (N_13265,N_8164,N_8309);
nand U13266 (N_13266,N_11245,N_8132);
or U13267 (N_13267,N_6761,N_7634);
nand U13268 (N_13268,N_10002,N_8088);
and U13269 (N_13269,N_11048,N_8741);
nor U13270 (N_13270,N_8807,N_9669);
nor U13271 (N_13271,N_6605,N_10629);
xnor U13272 (N_13272,N_6353,N_6874);
nor U13273 (N_13273,N_7211,N_11721);
or U13274 (N_13274,N_11744,N_9862);
nor U13275 (N_13275,N_7404,N_8192);
and U13276 (N_13276,N_10581,N_11379);
or U13277 (N_13277,N_7119,N_6772);
xor U13278 (N_13278,N_11672,N_9578);
or U13279 (N_13279,N_8187,N_7810);
nor U13280 (N_13280,N_6426,N_6624);
nand U13281 (N_13281,N_9906,N_8795);
or U13282 (N_13282,N_10796,N_11121);
and U13283 (N_13283,N_10325,N_11133);
xor U13284 (N_13284,N_9001,N_9499);
or U13285 (N_13285,N_6123,N_8608);
xor U13286 (N_13286,N_9085,N_7391);
nor U13287 (N_13287,N_10590,N_7931);
nor U13288 (N_13288,N_9219,N_10736);
nor U13289 (N_13289,N_8428,N_7971);
nand U13290 (N_13290,N_8079,N_10009);
nor U13291 (N_13291,N_11796,N_7136);
xnor U13292 (N_13292,N_9101,N_7421);
nor U13293 (N_13293,N_7014,N_11397);
nor U13294 (N_13294,N_7229,N_10384);
xnor U13295 (N_13295,N_6526,N_6497);
nand U13296 (N_13296,N_8709,N_8914);
nand U13297 (N_13297,N_8836,N_8257);
xor U13298 (N_13298,N_9359,N_6047);
or U13299 (N_13299,N_8757,N_10510);
or U13300 (N_13300,N_6548,N_9766);
nor U13301 (N_13301,N_6078,N_9652);
xor U13302 (N_13302,N_7341,N_9452);
and U13303 (N_13303,N_11515,N_10654);
and U13304 (N_13304,N_9015,N_6956);
nor U13305 (N_13305,N_6712,N_7504);
or U13306 (N_13306,N_9985,N_6500);
nor U13307 (N_13307,N_8531,N_10509);
nor U13308 (N_13308,N_11547,N_11035);
nor U13309 (N_13309,N_7899,N_9567);
or U13310 (N_13310,N_10090,N_7018);
or U13311 (N_13311,N_11311,N_8265);
xnor U13312 (N_13312,N_9284,N_6859);
xnor U13313 (N_13313,N_9259,N_9395);
nor U13314 (N_13314,N_11038,N_7140);
xnor U13315 (N_13315,N_9958,N_9127);
or U13316 (N_13316,N_11908,N_10366);
xnor U13317 (N_13317,N_10112,N_7700);
nor U13318 (N_13318,N_6328,N_7183);
or U13319 (N_13319,N_11983,N_7929);
or U13320 (N_13320,N_7779,N_11354);
nor U13321 (N_13321,N_8752,N_8361);
and U13322 (N_13322,N_7602,N_11907);
nor U13323 (N_13323,N_8103,N_9793);
and U13324 (N_13324,N_9610,N_10189);
nor U13325 (N_13325,N_8800,N_6795);
nor U13326 (N_13326,N_10801,N_10178);
or U13327 (N_13327,N_10234,N_11213);
nor U13328 (N_13328,N_6324,N_8515);
or U13329 (N_13329,N_7241,N_6127);
and U13330 (N_13330,N_9562,N_6937);
nand U13331 (N_13331,N_11318,N_10455);
xnor U13332 (N_13332,N_6513,N_9973);
nor U13333 (N_13333,N_6784,N_8035);
xnor U13334 (N_13334,N_6946,N_10220);
nand U13335 (N_13335,N_11287,N_9758);
and U13336 (N_13336,N_9705,N_9055);
and U13337 (N_13337,N_9223,N_6222);
nor U13338 (N_13338,N_7711,N_8488);
xnor U13339 (N_13339,N_10151,N_6141);
xnor U13340 (N_13340,N_10378,N_6116);
nor U13341 (N_13341,N_8824,N_11765);
nand U13342 (N_13342,N_8080,N_9556);
nand U13343 (N_13343,N_9191,N_11454);
and U13344 (N_13344,N_8872,N_11168);
nor U13345 (N_13345,N_8862,N_7639);
xor U13346 (N_13346,N_9280,N_6857);
and U13347 (N_13347,N_10655,N_6922);
or U13348 (N_13348,N_10373,N_11654);
nor U13349 (N_13349,N_11201,N_6916);
nand U13350 (N_13350,N_8613,N_7053);
nor U13351 (N_13351,N_9032,N_7669);
or U13352 (N_13352,N_6865,N_8786);
xnor U13353 (N_13353,N_10913,N_7697);
nand U13354 (N_13354,N_8423,N_6630);
xor U13355 (N_13355,N_10376,N_9683);
and U13356 (N_13356,N_10892,N_10770);
or U13357 (N_13357,N_8301,N_10805);
nor U13358 (N_13358,N_8815,N_11165);
or U13359 (N_13359,N_10430,N_10780);
and U13360 (N_13360,N_6880,N_6486);
nand U13361 (N_13361,N_8421,N_7824);
nand U13362 (N_13362,N_7415,N_8999);
and U13363 (N_13363,N_6200,N_7176);
nor U13364 (N_13364,N_8478,N_10651);
or U13365 (N_13365,N_11650,N_6082);
xor U13366 (N_13366,N_10891,N_6258);
nor U13367 (N_13367,N_6004,N_11493);
and U13368 (N_13368,N_8631,N_9899);
nand U13369 (N_13369,N_8157,N_9366);
and U13370 (N_13370,N_11512,N_7267);
and U13371 (N_13371,N_11471,N_7115);
nor U13372 (N_13372,N_7944,N_9642);
nor U13373 (N_13373,N_6727,N_8565);
and U13374 (N_13374,N_9033,N_11430);
and U13375 (N_13375,N_11615,N_9433);
xor U13376 (N_13376,N_11010,N_9528);
and U13377 (N_13377,N_8543,N_11109);
nand U13378 (N_13378,N_9415,N_10283);
and U13379 (N_13379,N_11849,N_6534);
and U13380 (N_13380,N_8662,N_11388);
and U13381 (N_13381,N_8458,N_7160);
nor U13382 (N_13382,N_6987,N_9855);
nand U13383 (N_13383,N_9253,N_11482);
nor U13384 (N_13384,N_6765,N_11080);
nor U13385 (N_13385,N_6482,N_11782);
or U13386 (N_13386,N_8205,N_9024);
nor U13387 (N_13387,N_10717,N_11923);
and U13388 (N_13388,N_11870,N_9362);
nor U13389 (N_13389,N_11412,N_8490);
or U13390 (N_13390,N_7209,N_11163);
nor U13391 (N_13391,N_6304,N_6183);
and U13392 (N_13392,N_8430,N_10879);
and U13393 (N_13393,N_6609,N_11544);
and U13394 (N_13394,N_8511,N_9595);
and U13395 (N_13395,N_7152,N_9016);
nand U13396 (N_13396,N_8045,N_6483);
nor U13397 (N_13397,N_9458,N_6215);
xnor U13398 (N_13398,N_11246,N_6450);
xnor U13399 (N_13399,N_6951,N_9721);
xor U13400 (N_13400,N_6134,N_11451);
nand U13401 (N_13401,N_7572,N_9332);
xor U13402 (N_13402,N_10022,N_11922);
nand U13403 (N_13403,N_8135,N_9835);
nand U13404 (N_13404,N_8036,N_10731);
nand U13405 (N_13405,N_6246,N_11752);
and U13406 (N_13406,N_11889,N_10625);
or U13407 (N_13407,N_9704,N_6449);
xnor U13408 (N_13408,N_8765,N_9421);
nor U13409 (N_13409,N_7959,N_10588);
and U13410 (N_13410,N_10214,N_9409);
xor U13411 (N_13411,N_11772,N_10082);
nor U13412 (N_13412,N_7260,N_10844);
nor U13413 (N_13413,N_7833,N_10779);
or U13414 (N_13414,N_8622,N_8393);
and U13415 (N_13415,N_7045,N_10906);
xor U13416 (N_13416,N_7378,N_7930);
nand U13417 (N_13417,N_8492,N_10344);
and U13418 (N_13418,N_6966,N_8528);
or U13419 (N_13419,N_7946,N_10501);
xor U13420 (N_13420,N_7245,N_8568);
xor U13421 (N_13421,N_6929,N_11103);
nor U13422 (N_13422,N_6064,N_10364);
nand U13423 (N_13423,N_10464,N_6271);
xor U13424 (N_13424,N_10526,N_6167);
nand U13425 (N_13425,N_10523,N_6945);
or U13426 (N_13426,N_6221,N_7005);
nor U13427 (N_13427,N_10671,N_10921);
nor U13428 (N_13428,N_9677,N_11049);
or U13429 (N_13429,N_11644,N_11697);
nor U13430 (N_13430,N_11362,N_9670);
and U13431 (N_13431,N_6326,N_7563);
and U13432 (N_13432,N_6014,N_7575);
and U13433 (N_13433,N_6525,N_9662);
and U13434 (N_13434,N_6719,N_7110);
nor U13435 (N_13435,N_6985,N_8049);
and U13436 (N_13436,N_10139,N_6071);
nor U13437 (N_13437,N_11885,N_11984);
xnor U13438 (N_13438,N_8689,N_9856);
nor U13439 (N_13439,N_7934,N_7786);
and U13440 (N_13440,N_7511,N_6849);
xnor U13441 (N_13441,N_6480,N_9739);
and U13442 (N_13442,N_8869,N_6997);
and U13443 (N_13443,N_7462,N_11345);
nor U13444 (N_13444,N_7094,N_6334);
nor U13445 (N_13445,N_11081,N_8779);
xor U13446 (N_13446,N_9809,N_9889);
nand U13447 (N_13447,N_7529,N_10596);
nand U13448 (N_13448,N_8845,N_7350);
or U13449 (N_13449,N_10816,N_9583);
xor U13450 (N_13450,N_9440,N_9593);
and U13451 (N_13451,N_10722,N_11824);
or U13452 (N_13452,N_8258,N_10153);
nand U13453 (N_13453,N_8217,N_8278);
xor U13454 (N_13454,N_8959,N_10860);
or U13455 (N_13455,N_7605,N_6801);
and U13456 (N_13456,N_11419,N_7158);
nor U13457 (N_13457,N_6544,N_7827);
and U13458 (N_13458,N_9803,N_9560);
or U13459 (N_13459,N_7495,N_8947);
nor U13460 (N_13460,N_7412,N_9800);
or U13461 (N_13461,N_11539,N_6809);
nor U13462 (N_13462,N_7296,N_6563);
xor U13463 (N_13463,N_10527,N_9165);
xnor U13464 (N_13464,N_8413,N_9378);
xor U13465 (N_13465,N_8640,N_6427);
and U13466 (N_13466,N_7720,N_8482);
nand U13467 (N_13467,N_8261,N_10885);
nor U13468 (N_13468,N_8787,N_6357);
xnor U13469 (N_13469,N_10597,N_6044);
nand U13470 (N_13470,N_7665,N_7447);
nor U13471 (N_13471,N_10862,N_10427);
and U13472 (N_13472,N_8547,N_9353);
xnor U13473 (N_13473,N_9962,N_10353);
or U13474 (N_13474,N_11094,N_10406);
or U13475 (N_13475,N_11611,N_7856);
or U13476 (N_13476,N_10101,N_6302);
xnor U13477 (N_13477,N_9012,N_8351);
nand U13478 (N_13478,N_11181,N_10825);
and U13479 (N_13479,N_9488,N_7144);
nor U13480 (N_13480,N_6747,N_6995);
or U13481 (N_13481,N_9386,N_11816);
xor U13482 (N_13482,N_7482,N_8052);
xor U13483 (N_13483,N_6053,N_11542);
or U13484 (N_13484,N_8022,N_8909);
xor U13485 (N_13485,N_7888,N_10809);
nand U13486 (N_13486,N_10146,N_11177);
or U13487 (N_13487,N_10899,N_10198);
or U13488 (N_13488,N_7648,N_10994);
nand U13489 (N_13489,N_10987,N_7142);
nand U13490 (N_13490,N_7066,N_11609);
nand U13491 (N_13491,N_8465,N_7373);
nor U13492 (N_13492,N_11851,N_6696);
xor U13493 (N_13493,N_9681,N_6121);
nand U13494 (N_13494,N_8448,N_6746);
xnor U13495 (N_13495,N_8937,N_10612);
xor U13496 (N_13496,N_7709,N_8316);
nand U13497 (N_13497,N_8078,N_8472);
xnor U13498 (N_13498,N_6566,N_8412);
xnor U13499 (N_13499,N_11680,N_10894);
or U13500 (N_13500,N_10683,N_11157);
xnor U13501 (N_13501,N_10068,N_10392);
nand U13502 (N_13502,N_11950,N_6087);
and U13503 (N_13503,N_7116,N_6146);
nor U13504 (N_13504,N_11776,N_10701);
and U13505 (N_13505,N_10357,N_10883);
nor U13506 (N_13506,N_7328,N_8337);
or U13507 (N_13507,N_11369,N_9125);
nand U13508 (N_13508,N_6545,N_10206);
nand U13509 (N_13509,N_6313,N_8074);
xor U13510 (N_13510,N_11632,N_6256);
and U13511 (N_13511,N_11324,N_11723);
and U13512 (N_13512,N_6282,N_11595);
or U13513 (N_13513,N_9790,N_8781);
nor U13514 (N_13514,N_7623,N_10867);
nor U13515 (N_13515,N_9945,N_9428);
xor U13516 (N_13516,N_8168,N_11037);
xnor U13517 (N_13517,N_11415,N_7887);
xnor U13518 (N_13518,N_11797,N_10903);
and U13519 (N_13519,N_11357,N_8749);
or U13520 (N_13520,N_11012,N_9495);
nor U13521 (N_13521,N_6385,N_10191);
or U13522 (N_13522,N_8026,N_9357);
nand U13523 (N_13523,N_8849,N_11088);
and U13524 (N_13524,N_6778,N_11395);
nand U13525 (N_13525,N_11256,N_10525);
or U13526 (N_13526,N_10196,N_10126);
or U13527 (N_13527,N_6036,N_8695);
or U13528 (N_13528,N_10176,N_7455);
and U13529 (N_13529,N_10223,N_10718);
xnor U13530 (N_13530,N_10145,N_6879);
or U13531 (N_13531,N_7261,N_11935);
or U13532 (N_13532,N_11334,N_11603);
nand U13533 (N_13533,N_9113,N_9279);
or U13534 (N_13534,N_9808,N_6542);
xor U13535 (N_13535,N_6369,N_8023);
or U13536 (N_13536,N_8573,N_8151);
nand U13537 (N_13537,N_9702,N_7355);
xnor U13538 (N_13538,N_10765,N_8854);
nand U13539 (N_13539,N_7070,N_6650);
and U13540 (N_13540,N_10848,N_10767);
nor U13541 (N_13541,N_8747,N_11974);
nor U13542 (N_13542,N_6996,N_10505);
nand U13543 (N_13543,N_9217,N_11734);
or U13544 (N_13544,N_8401,N_6668);
nor U13545 (N_13545,N_10508,N_11282);
xor U13546 (N_13546,N_6333,N_8122);
nor U13547 (N_13547,N_7459,N_8152);
and U13548 (N_13548,N_11126,N_8174);
nor U13549 (N_13549,N_6983,N_9863);
and U13550 (N_13550,N_7784,N_11207);
nor U13551 (N_13551,N_6205,N_9519);
xor U13552 (N_13552,N_6175,N_8818);
and U13553 (N_13553,N_6549,N_9575);
xnor U13554 (N_13554,N_10482,N_8769);
nor U13555 (N_13555,N_7560,N_9940);
nand U13556 (N_13556,N_11624,N_7901);
nand U13557 (N_13557,N_9427,N_8058);
or U13558 (N_13558,N_11328,N_7220);
or U13559 (N_13559,N_6473,N_7909);
xor U13560 (N_13560,N_6590,N_7169);
and U13561 (N_13561,N_6218,N_6861);
or U13562 (N_13562,N_6337,N_7326);
and U13563 (N_13563,N_11534,N_9883);
nand U13564 (N_13564,N_8240,N_11464);
or U13565 (N_13565,N_10067,N_10803);
nand U13566 (N_13566,N_9748,N_8081);
xnor U13567 (N_13567,N_10073,N_7912);
nand U13568 (N_13568,N_6381,N_7113);
nand U13569 (N_13569,N_6470,N_9164);
and U13570 (N_13570,N_10459,N_7768);
nor U13571 (N_13571,N_11939,N_7982);
nor U13572 (N_13572,N_8847,N_11833);
nor U13573 (N_13573,N_6611,N_9570);
nor U13574 (N_13574,N_9471,N_11065);
and U13575 (N_13575,N_7257,N_11469);
nor U13576 (N_13576,N_9606,N_11237);
nand U13577 (N_13577,N_10985,N_11082);
xnor U13578 (N_13578,N_6325,N_9603);
nand U13579 (N_13579,N_11288,N_8932);
or U13580 (N_13580,N_7148,N_9627);
nor U13581 (N_13581,N_9917,N_7690);
and U13582 (N_13582,N_7875,N_6112);
and U13583 (N_13583,N_9058,N_8972);
nor U13584 (N_13584,N_10410,N_10648);
or U13585 (N_13585,N_6466,N_6732);
nor U13586 (N_13586,N_8582,N_9134);
nand U13587 (N_13587,N_7956,N_11751);
nand U13588 (N_13588,N_9872,N_11120);
and U13589 (N_13589,N_11392,N_10335);
and U13590 (N_13590,N_9882,N_11929);
or U13591 (N_13591,N_6339,N_11732);
and U13592 (N_13592,N_7004,N_7999);
nand U13593 (N_13593,N_8471,N_8936);
and U13594 (N_13594,N_7420,N_11249);
nand U13595 (N_13595,N_11385,N_10591);
and U13596 (N_13596,N_6266,N_6776);
nand U13597 (N_13597,N_10601,N_11227);
xnor U13598 (N_13598,N_8296,N_9996);
xnor U13599 (N_13599,N_8863,N_6414);
and U13600 (N_13600,N_8809,N_11188);
nor U13601 (N_13601,N_9997,N_7746);
or U13602 (N_13602,N_9513,N_8062);
xor U13603 (N_13603,N_7549,N_10982);
or U13604 (N_13604,N_8263,N_11771);
or U13605 (N_13605,N_9710,N_11576);
nand U13606 (N_13606,N_10255,N_10057);
nand U13607 (N_13607,N_6964,N_8212);
and U13608 (N_13608,N_6390,N_7047);
nor U13609 (N_13609,N_7900,N_10203);
xnor U13610 (N_13610,N_8200,N_10024);
xnor U13611 (N_13611,N_10747,N_9667);
nand U13612 (N_13612,N_7736,N_8827);
or U13613 (N_13613,N_11900,N_10902);
or U13614 (N_13614,N_8973,N_8860);
and U13615 (N_13615,N_6211,N_9034);
xor U13616 (N_13616,N_10502,N_10920);
and U13617 (N_13617,N_9554,N_9425);
nor U13618 (N_13618,N_9923,N_9865);
nor U13619 (N_13619,N_11135,N_9211);
nand U13620 (N_13620,N_9049,N_8755);
xnor U13621 (N_13621,N_9306,N_10072);
nand U13622 (N_13622,N_8751,N_8219);
or U13623 (N_13623,N_10078,N_10975);
nor U13624 (N_13624,N_10645,N_10084);
xor U13625 (N_13625,N_11068,N_10608);
nor U13626 (N_13626,N_7821,N_11531);
xnor U13627 (N_13627,N_7782,N_10158);
and U13628 (N_13628,N_6281,N_6176);
or U13629 (N_13629,N_8618,N_7790);
and U13630 (N_13630,N_11679,N_11403);
nor U13631 (N_13631,N_11548,N_11562);
nand U13632 (N_13632,N_8982,N_6882);
or U13633 (N_13633,N_6541,N_11694);
nand U13634 (N_13634,N_6194,N_10680);
or U13635 (N_13635,N_10229,N_6309);
nor U13636 (N_13636,N_6757,N_9255);
or U13637 (N_13637,N_8594,N_8610);
nand U13638 (N_13638,N_10643,N_10314);
nor U13639 (N_13639,N_7981,N_8682);
nor U13640 (N_13640,N_6415,N_11794);
nor U13641 (N_13641,N_8139,N_11712);
nor U13642 (N_13642,N_9780,N_6594);
nor U13643 (N_13643,N_10274,N_6191);
nand U13644 (N_13644,N_10559,N_7497);
nand U13645 (N_13645,N_7392,N_8954);
nand U13646 (N_13646,N_10536,N_10170);
nor U13647 (N_13647,N_9018,N_10602);
nor U13648 (N_13648,N_7915,N_6238);
nand U13649 (N_13649,N_9252,N_6356);
or U13650 (N_13650,N_6914,N_11091);
nand U13651 (N_13651,N_6142,N_9204);
nand U13652 (N_13652,N_8879,N_7577);
or U13653 (N_13653,N_7740,N_11803);
xor U13654 (N_13654,N_7213,N_10315);
xnor U13655 (N_13655,N_6744,N_6667);
xor U13656 (N_13656,N_8166,N_6278);
nand U13657 (N_13657,N_6952,N_8900);
or U13658 (N_13658,N_10853,N_10901);
xnor U13659 (N_13659,N_7224,N_9873);
nor U13660 (N_13660,N_7518,N_7166);
xnor U13661 (N_13661,N_6705,N_10652);
nor U13662 (N_13662,N_8266,N_7889);
xnor U13663 (N_13663,N_10775,N_10062);
xnor U13664 (N_13664,N_11267,N_6898);
xnor U13665 (N_13665,N_7940,N_8880);
xor U13666 (N_13666,N_8020,N_10425);
and U13667 (N_13667,N_9180,N_6170);
nor U13668 (N_13668,N_8012,N_11347);
or U13669 (N_13669,N_7873,N_10969);
nand U13670 (N_13670,N_11628,N_6921);
xor U13671 (N_13671,N_9881,N_7467);
xnor U13672 (N_13672,N_10799,N_10489);
nand U13673 (N_13673,N_10716,N_10884);
or U13674 (N_13674,N_11263,N_7706);
and U13675 (N_13675,N_7541,N_11956);
nand U13676 (N_13676,N_11913,N_7040);
nand U13677 (N_13677,N_10419,N_6992);
xor U13678 (N_13678,N_10262,N_6892);
nand U13679 (N_13679,N_8521,N_10230);
or U13680 (N_13680,N_7318,N_11711);
or U13681 (N_13681,N_7345,N_8853);
or U13682 (N_13682,N_9589,N_8648);
or U13683 (N_13683,N_11241,N_7766);
xor U13684 (N_13684,N_9910,N_9356);
and U13685 (N_13685,N_11286,N_10081);
xnor U13686 (N_13686,N_8718,N_9741);
nand U13687 (N_13687,N_6873,N_6798);
or U13688 (N_13688,N_9310,N_7754);
or U13689 (N_13689,N_8655,N_8514);
nor U13690 (N_13690,N_6893,N_6647);
and U13691 (N_13691,N_10618,N_10693);
and U13692 (N_13692,N_11800,N_11402);
nand U13693 (N_13693,N_9282,N_10925);
nor U13694 (N_13694,N_9718,N_8702);
xnor U13695 (N_13695,N_10952,N_9755);
and U13696 (N_13696,N_7922,N_10269);
nand U13697 (N_13697,N_7173,N_10705);
nand U13698 (N_13698,N_10640,N_8665);
nor U13699 (N_13699,N_9968,N_10290);
xor U13700 (N_13700,N_11450,N_10758);
or U13701 (N_13701,N_7506,N_11206);
nor U13702 (N_13702,N_6019,N_10359);
nand U13703 (N_13703,N_9811,N_8967);
nor U13704 (N_13704,N_8846,N_6657);
nand U13705 (N_13705,N_8147,N_7399);
or U13706 (N_13706,N_6740,N_7500);
and U13707 (N_13707,N_10864,N_10556);
or U13708 (N_13708,N_11470,N_11535);
and U13709 (N_13709,N_6555,N_7653);
xnor U13710 (N_13710,N_11742,N_11093);
nand U13711 (N_13711,N_11085,N_10886);
nor U13712 (N_13712,N_11022,N_7661);
and U13713 (N_13713,N_11164,N_10548);
nor U13714 (N_13714,N_7131,N_10951);
xor U13715 (N_13715,N_11016,N_8523);
nand U13716 (N_13716,N_6180,N_8708);
nand U13717 (N_13717,N_6759,N_9469);
xor U13718 (N_13718,N_10444,N_11031);
nor U13719 (N_13719,N_6410,N_6251);
nand U13720 (N_13720,N_10441,N_10727);
xnor U13721 (N_13721,N_6168,N_9319);
nor U13722 (N_13722,N_7886,N_11437);
or U13723 (N_13723,N_7410,N_7604);
nand U13724 (N_13724,N_8055,N_6320);
or U13725 (N_13725,N_8193,N_9190);
nand U13726 (N_13726,N_9212,N_8244);
or U13727 (N_13727,N_9273,N_9309);
and U13728 (N_13728,N_11655,N_6618);
and U13729 (N_13729,N_6028,N_11887);
nor U13730 (N_13730,N_6734,N_7798);
nor U13731 (N_13731,N_8607,N_11250);
nand U13732 (N_13732,N_6423,N_7268);
xnor U13733 (N_13733,N_9805,N_10356);
nand U13734 (N_13734,N_8878,N_7613);
nor U13735 (N_13735,N_8137,N_8279);
xor U13736 (N_13736,N_7846,N_9346);
nor U13737 (N_13737,N_7668,N_9481);
nand U13738 (N_13738,N_7390,N_7227);
xnor U13739 (N_13739,N_10063,N_11528);
and U13740 (N_13740,N_6852,N_9009);
xnor U13741 (N_13741,N_10298,N_8644);
nor U13742 (N_13742,N_10115,N_11421);
nand U13743 (N_13743,N_9260,N_6506);
and U13744 (N_13744,N_9334,N_6054);
and U13745 (N_13745,N_9637,N_9639);
xor U13746 (N_13746,N_8416,N_11667);
or U13747 (N_13747,N_11119,N_6932);
or U13748 (N_13748,N_8509,N_11076);
xor U13749 (N_13749,N_11853,N_9731);
nor U13750 (N_13750,N_7247,N_10188);
or U13751 (N_13751,N_6896,N_9295);
nor U13752 (N_13752,N_10332,N_8576);
and U13753 (N_13753,N_7652,N_11620);
nand U13754 (N_13754,N_10000,N_9788);
nand U13755 (N_13755,N_10513,N_11136);
nor U13756 (N_13756,N_8180,N_6895);
nand U13757 (N_13757,N_7419,N_9159);
xor U13758 (N_13758,N_8148,N_6462);
nand U13759 (N_13759,N_10345,N_7265);
nand U13760 (N_13760,N_11973,N_6631);
xor U13761 (N_13761,N_10141,N_9896);
and U13762 (N_13762,N_8890,N_9206);
nand U13763 (N_13763,N_9493,N_7151);
or U13764 (N_13764,N_9215,N_10264);
nand U13765 (N_13765,N_6291,N_9843);
xor U13766 (N_13766,N_10815,N_7149);
xnor U13767 (N_13767,N_10161,N_10889);
xnor U13768 (N_13768,N_7696,N_10025);
or U13769 (N_13769,N_10004,N_6442);
or U13770 (N_13770,N_10233,N_11301);
or U13771 (N_13771,N_8570,N_9514);
nand U13772 (N_13772,N_8163,N_9969);
nor U13773 (N_13773,N_8630,N_10466);
nand U13774 (N_13774,N_9196,N_7752);
and U13775 (N_13775,N_7418,N_7228);
nor U13776 (N_13776,N_6787,N_6135);
nand U13777 (N_13777,N_8047,N_11861);
and U13778 (N_13778,N_6287,N_6708);
and U13779 (N_13779,N_10633,N_7323);
nand U13780 (N_13780,N_9060,N_11736);
nand U13781 (N_13781,N_9239,N_7407);
xnor U13782 (N_13782,N_9719,N_11075);
nor U13783 (N_13783,N_7750,N_6961);
or U13784 (N_13784,N_8071,N_9050);
nor U13785 (N_13785,N_7794,N_9712);
nor U13786 (N_13786,N_8924,N_10397);
nand U13787 (N_13787,N_6886,N_6845);
nand U13788 (N_13788,N_6860,N_11372);
and U13789 (N_13789,N_10535,N_10945);
or U13790 (N_13790,N_11706,N_6000);
xnor U13791 (N_13791,N_9924,N_9410);
and U13792 (N_13792,N_10473,N_11176);
or U13793 (N_13793,N_8002,N_7580);
nand U13794 (N_13794,N_7015,N_11319);
nand U13795 (N_13795,N_11979,N_9938);
or U13796 (N_13796,N_7286,N_9503);
xnor U13797 (N_13797,N_10309,N_11111);
nand U13798 (N_13798,N_9453,N_10337);
or U13799 (N_13799,N_6870,N_8232);
nor U13800 (N_13800,N_6101,N_9581);
or U13801 (N_13801,N_7039,N_10046);
nand U13802 (N_13802,N_9918,N_8111);
xnor U13803 (N_13803,N_9120,N_7885);
and U13804 (N_13804,N_6713,N_11146);
and U13805 (N_13805,N_7146,N_10650);
or U13806 (N_13806,N_8092,N_9526);
nand U13807 (N_13807,N_7233,N_9278);
and U13808 (N_13808,N_7480,N_7829);
nand U13809 (N_13809,N_7042,N_8362);
nand U13810 (N_13810,N_8269,N_7664);
or U13811 (N_13811,N_11275,N_11260);
and U13812 (N_13812,N_8715,N_6484);
nand U13813 (N_13813,N_11662,N_10012);
nand U13814 (N_13814,N_8770,N_8814);
xor U13815 (N_13815,N_10550,N_7019);
nor U13816 (N_13816,N_7666,N_9177);
nor U13817 (N_13817,N_11552,N_11416);
nor U13818 (N_13818,N_10932,N_9148);
xor U13819 (N_13819,N_7928,N_7282);
nand U13820 (N_13820,N_6386,N_7617);
xor U13821 (N_13821,N_6203,N_8352);
or U13822 (N_13822,N_10595,N_6199);
nor U13823 (N_13823,N_9448,N_10668);
or U13824 (N_13824,N_9185,N_10914);
and U13825 (N_13825,N_8077,N_9946);
and U13826 (N_13826,N_10694,N_11674);
xor U13827 (N_13827,N_7333,N_8455);
xnor U13828 (N_13828,N_6819,N_9129);
and U13829 (N_13829,N_8530,N_9447);
and U13830 (N_13830,N_7380,N_6869);
or U13831 (N_13831,N_6063,N_11932);
nand U13832 (N_13832,N_7385,N_6763);
or U13833 (N_13833,N_9377,N_7556);
nor U13834 (N_13834,N_10841,N_8801);
and U13835 (N_13835,N_9587,N_7010);
nor U13836 (N_13836,N_11383,N_11614);
and U13837 (N_13837,N_6902,N_6195);
or U13838 (N_13838,N_11894,N_8699);
nor U13839 (N_13839,N_7629,N_11033);
nand U13840 (N_13840,N_9114,N_6841);
and U13841 (N_13841,N_11348,N_6017);
xor U13842 (N_13842,N_8339,N_11976);
nand U13843 (N_13843,N_11341,N_10833);
or U13844 (N_13844,N_9840,N_6060);
nand U13845 (N_13845,N_6940,N_7764);
and U13846 (N_13846,N_8838,N_8859);
nand U13847 (N_13847,N_9316,N_9636);
nand U13848 (N_13848,N_7637,N_8104);
nor U13849 (N_13849,N_6614,N_6217);
nor U13850 (N_13850,N_6487,N_7785);
nand U13851 (N_13851,N_7434,N_8724);
or U13852 (N_13852,N_6596,N_8184);
nand U13853 (N_13853,N_10487,N_6889);
nor U13854 (N_13854,N_10991,N_10295);
or U13855 (N_13855,N_6463,N_8350);
or U13856 (N_13856,N_10549,N_10954);
or U13857 (N_13857,N_10211,N_6150);
and U13858 (N_13858,N_10732,N_11658);
nor U13859 (N_13859,N_6671,N_8526);
xnor U13860 (N_13860,N_7114,N_9698);
nand U13861 (N_13861,N_10173,N_7307);
nand U13862 (N_13862,N_11613,N_8774);
xor U13863 (N_13863,N_11508,N_9408);
xnor U13864 (N_13864,N_8775,N_6844);
nor U13865 (N_13865,N_11845,N_6768);
nand U13866 (N_13866,N_11373,N_7654);
and U13867 (N_13867,N_11958,N_11838);
xnor U13868 (N_13868,N_8281,N_7636);
nor U13869 (N_13869,N_10931,N_9611);
xnor U13870 (N_13870,N_10734,N_11942);
nor U13871 (N_13871,N_7537,N_10375);
xor U13872 (N_13872,N_9909,N_9660);
nand U13873 (N_13873,N_6070,N_10644);
nand U13874 (N_13874,N_7876,N_11305);
or U13875 (N_13875,N_11760,N_6955);
and U13876 (N_13876,N_8363,N_9137);
or U13877 (N_13877,N_10218,N_10930);
xnor U13878 (N_13878,N_9156,N_8161);
or U13879 (N_13879,N_6615,N_9084);
or U13880 (N_13880,N_6655,N_10543);
xnor U13881 (N_13881,N_6209,N_7361);
nor U13882 (N_13882,N_9770,N_6943);
nand U13883 (N_13883,N_9404,N_11456);
and U13884 (N_13884,N_9199,N_8522);
or U13885 (N_13885,N_6001,N_6840);
or U13886 (N_13886,N_11635,N_8590);
nand U13887 (N_13887,N_7984,N_10447);
and U13888 (N_13888,N_10609,N_11763);
and U13889 (N_13889,N_7804,N_8469);
or U13890 (N_13890,N_10522,N_7826);
or U13891 (N_13891,N_6418,N_9187);
and U13892 (N_13892,N_8803,N_10263);
nand U13893 (N_13893,N_7951,N_8980);
and U13894 (N_13894,N_7383,N_8559);
or U13895 (N_13895,N_10910,N_11375);
xnor U13896 (N_13896,N_10349,N_9062);
or U13897 (N_13897,N_11933,N_11954);
and U13898 (N_13898,N_8667,N_6722);
or U13899 (N_13899,N_10240,N_10076);
and U13900 (N_13900,N_9040,N_11350);
nor U13901 (N_13901,N_6433,N_8171);
or U13902 (N_13902,N_7539,N_8252);
or U13903 (N_13903,N_6037,N_9690);
nor U13904 (N_13904,N_11663,N_9294);
xnor U13905 (N_13905,N_6184,N_10580);
nand U13906 (N_13906,N_6866,N_8425);
and U13907 (N_13907,N_9406,N_9336);
nor U13908 (N_13908,N_10695,N_9579);
nor U13909 (N_13909,N_9478,N_10405);
or U13910 (N_13910,N_6029,N_8085);
nor U13911 (N_13911,N_9053,N_8653);
and U13912 (N_13912,N_11320,N_10069);
or U13913 (N_13913,N_7800,N_7683);
xor U13914 (N_13914,N_10294,N_7001);
or U13915 (N_13915,N_8420,N_7332);
xor U13916 (N_13916,N_9109,N_9517);
xor U13917 (N_13917,N_7841,N_6247);
nor U13918 (N_13918,N_8094,N_10949);
nor U13919 (N_13919,N_10570,N_6651);
or U13920 (N_13920,N_9957,N_8125);
and U13921 (N_13921,N_10751,N_9696);
or U13922 (N_13922,N_7646,N_8584);
nand U13923 (N_13923,N_11423,N_11173);
or U13924 (N_13924,N_10735,N_10813);
xnor U13925 (N_13925,N_8484,N_6046);
and U13926 (N_13926,N_6104,N_9678);
nand U13927 (N_13927,N_10445,N_10085);
or U13928 (N_13928,N_7312,N_6836);
and U13929 (N_13929,N_6081,N_6137);
xor U13930 (N_13930,N_7162,N_6773);
and U13931 (N_13931,N_8387,N_6593);
xor U13932 (N_13932,N_8324,N_6091);
xnor U13933 (N_13933,N_11717,N_6904);
and U13934 (N_13934,N_7507,N_6685);
nor U13935 (N_13935,N_11386,N_11904);
xor U13936 (N_13936,N_7987,N_11577);
xor U13937 (N_13937,N_11688,N_6149);
or U13938 (N_13938,N_11221,N_8005);
and U13939 (N_13939,N_7523,N_7244);
nor U13940 (N_13940,N_11503,N_8917);
or U13941 (N_13941,N_10299,N_10660);
and U13942 (N_13942,N_11506,N_10358);
nand U13943 (N_13943,N_11724,N_10442);
or U13944 (N_13944,N_8868,N_8953);
xnor U13945 (N_13945,N_11156,N_10083);
nand U13946 (N_13946,N_11491,N_9919);
nor U13947 (N_13947,N_10070,N_11285);
and U13948 (N_13948,N_11622,N_9869);
and U13949 (N_13949,N_11787,N_9315);
xnor U13950 (N_13950,N_7562,N_10369);
and U13951 (N_13951,N_9629,N_7109);
nand U13952 (N_13952,N_9105,N_7849);
and U13953 (N_13953,N_11863,N_10933);
and U13954 (N_13954,N_9993,N_8341);
nor U13955 (N_13955,N_6789,N_8823);
and U13956 (N_13956,N_10499,N_9716);
and U13957 (N_13957,N_11978,N_6231);
nor U13958 (N_13958,N_8124,N_7121);
xnor U13959 (N_13959,N_9597,N_9236);
nor U13960 (N_13960,N_11183,N_6109);
or U13961 (N_13961,N_7321,N_6682);
xnor U13962 (N_13962,N_9110,N_7486);
nor U13963 (N_13963,N_6510,N_11831);
nor U13964 (N_13964,N_10280,N_8110);
nand U13965 (N_13965,N_8811,N_9857);
xor U13966 (N_13966,N_11488,N_6083);
xnor U13967 (N_13967,N_7883,N_8182);
nor U13968 (N_13968,N_8654,N_6509);
and U13969 (N_13969,N_8595,N_10699);
and U13970 (N_13970,N_9189,N_7316);
nor U13971 (N_13971,N_11755,N_7835);
and U13972 (N_13972,N_7483,N_11561);
nand U13973 (N_13973,N_10142,N_6939);
nor U13974 (N_13974,N_11940,N_6193);
or U13975 (N_13975,N_11914,N_6040);
or U13976 (N_13976,N_11847,N_6284);
nand U13977 (N_13977,N_6202,N_11884);
or U13978 (N_13978,N_8920,N_6505);
or U13979 (N_13979,N_11597,N_9970);
or U13980 (N_13980,N_10120,N_6360);
and U13981 (N_13981,N_10582,N_6800);
xnor U13982 (N_13982,N_6055,N_10316);
or U13983 (N_13983,N_10279,N_8227);
or U13984 (N_13984,N_11321,N_10106);
or U13985 (N_13985,N_11669,N_10019);
nor U13986 (N_13986,N_10700,N_11462);
xnor U13987 (N_13987,N_7960,N_8011);
and U13988 (N_13988,N_7259,N_9706);
or U13989 (N_13989,N_6552,N_10696);
or U13990 (N_13990,N_10897,N_6010);
nor U13991 (N_13991,N_9673,N_10192);
nand U13992 (N_13992,N_10852,N_7758);
xnor U13993 (N_13993,N_10511,N_6432);
and U13994 (N_13994,N_11436,N_9072);
nor U13995 (N_13995,N_8555,N_10398);
or U13996 (N_13996,N_9102,N_10950);
and U13997 (N_13997,N_7422,N_6925);
xnor U13998 (N_13998,N_10014,N_11196);
xnor U13999 (N_13999,N_8675,N_8044);
or U14000 (N_14000,N_6973,N_8066);
and U14001 (N_14001,N_9695,N_8686);
nor U14002 (N_14002,N_8532,N_7201);
nor U14003 (N_14003,N_6842,N_6043);
nor U14004 (N_14004,N_6822,N_9875);
nor U14005 (N_14005,N_11793,N_10603);
nor U14006 (N_14006,N_8918,N_8922);
and U14007 (N_14007,N_11004,N_6728);
or U14008 (N_14008,N_6917,N_8624);
and U14009 (N_14009,N_8422,N_8552);
xor U14010 (N_14010,N_8489,N_7301);
or U14011 (N_14011,N_8096,N_6261);
xor U14012 (N_14012,N_8650,N_11589);
or U14013 (N_14013,N_11591,N_9145);
xor U14014 (N_14014,N_11223,N_7002);
or U14015 (N_14015,N_7908,N_9438);
and U14016 (N_14016,N_6850,N_7672);
nor U14017 (N_14017,N_9978,N_10225);
nor U14018 (N_14018,N_6875,N_6249);
or U14019 (N_14019,N_8209,N_7554);
or U14020 (N_14020,N_8483,N_6699);
or U14021 (N_14021,N_6300,N_11739);
nand U14022 (N_14022,N_6015,N_9885);
or U14023 (N_14023,N_11337,N_9205);
or U14024 (N_14024,N_11098,N_10519);
xor U14025 (N_14025,N_10389,N_11936);
or U14026 (N_14026,N_6516,N_10458);
nor U14027 (N_14027,N_11652,N_11064);
and U14028 (N_14028,N_9446,N_11545);
xor U14029 (N_14029,N_9274,N_6062);
nand U14030 (N_14030,N_8941,N_7597);
xor U14031 (N_14031,N_11629,N_10837);
xor U14032 (N_14032,N_6068,N_8705);
nand U14033 (N_14033,N_9767,N_7558);
or U14034 (N_14034,N_7453,N_8452);
and U14035 (N_14035,N_8467,N_11399);
xor U14036 (N_14036,N_11257,N_7016);
or U14037 (N_14037,N_6402,N_7874);
and U14038 (N_14038,N_10342,N_6521);
and U14039 (N_14039,N_8599,N_10600);
nor U14040 (N_14040,N_8128,N_10551);
nor U14041 (N_14041,N_10121,N_6825);
or U14042 (N_14042,N_10865,N_10111);
nand U14043 (N_14043,N_10673,N_6906);
or U14044 (N_14044,N_7638,N_11045);
nor U14045 (N_14045,N_8593,N_9106);
or U14046 (N_14046,N_8445,N_8344);
nand U14047 (N_14047,N_9474,N_8611);
xnor U14048 (N_14048,N_6196,N_10719);
nor U14049 (N_14049,N_9733,N_11880);
and U14050 (N_14050,N_9468,N_9061);
xnor U14051 (N_14051,N_7487,N_6340);
xnor U14052 (N_14052,N_11521,N_9247);
xnor U14053 (N_14053,N_10615,N_10759);
and U14054 (N_14054,N_6329,N_7626);
xnor U14055 (N_14055,N_6156,N_6529);
or U14056 (N_14056,N_7667,N_6378);
or U14057 (N_14057,N_10533,N_6920);
xor U14058 (N_14058,N_7616,N_6536);
nor U14059 (N_14059,N_9271,N_8598);
and U14060 (N_14060,N_10524,N_10594);
nand U14061 (N_14061,N_7643,N_8427);
nand U14062 (N_14062,N_11801,N_6749);
or U14063 (N_14063,N_11795,N_8789);
nand U14064 (N_14064,N_8995,N_8353);
nand U14065 (N_14065,N_8241,N_10669);
or U14066 (N_14066,N_8606,N_9363);
or U14067 (N_14067,N_9540,N_8315);
and U14068 (N_14068,N_11208,N_11808);
and U14069 (N_14069,N_9281,N_7037);
or U14070 (N_14070,N_11210,N_9214);
and U14071 (N_14071,N_11727,N_7397);
and U14072 (N_14072,N_8785,N_11151);
xor U14073 (N_14073,N_11822,N_6884);
nand U14074 (N_14074,N_9574,N_6748);
nand U14075 (N_14075,N_9981,N_6413);
or U14076 (N_14076,N_8691,N_10516);
xnor U14077 (N_14077,N_6088,N_6065);
nand U14078 (N_14078,N_7443,N_8748);
xnor U14079 (N_14079,N_6499,N_9614);
and U14080 (N_14080,N_6289,N_11356);
or U14081 (N_14081,N_7364,N_6382);
nand U14082 (N_14082,N_6206,N_10592);
or U14083 (N_14083,N_9751,N_7591);
nor U14084 (N_14084,N_10481,N_8457);
and U14085 (N_14085,N_8172,N_10679);
or U14086 (N_14086,N_10514,N_8601);
xor U14087 (N_14087,N_8098,N_6056);
xnor U14088 (N_14088,N_11799,N_9689);
and U14089 (N_14089,N_9272,N_10753);
or U14090 (N_14090,N_8634,N_10360);
or U14091 (N_14091,N_9934,N_9774);
or U14092 (N_14092,N_6097,N_7757);
or U14093 (N_14093,N_7478,N_9931);
nor U14094 (N_14094,N_10554,N_6627);
xor U14095 (N_14095,N_10286,N_7466);
or U14096 (N_14096,N_6456,N_11271);
or U14097 (N_14097,N_11683,N_11839);
or U14098 (N_14098,N_10259,N_11475);
and U14099 (N_14099,N_7186,N_11601);
xnor U14100 (N_14100,N_10711,N_7674);
xnor U14101 (N_14101,N_9728,N_6949);
nand U14102 (N_14102,N_11441,N_7175);
or U14103 (N_14103,N_6330,N_6715);
and U14104 (N_14104,N_7117,N_6288);
or U14105 (N_14105,N_7313,N_7293);
xnor U14106 (N_14106,N_8761,N_10617);
nand U14107 (N_14107,N_10990,N_6978);
nor U14108 (N_14108,N_9489,N_6797);
nor U14109 (N_14109,N_9858,N_8833);
nand U14110 (N_14110,N_11300,N_11483);
xor U14111 (N_14111,N_10010,N_10881);
nor U14112 (N_14112,N_11684,N_6554);
and U14113 (N_14113,N_9734,N_11586);
nand U14114 (N_14114,N_10003,N_7170);
or U14115 (N_14115,N_8865,N_6275);
or U14116 (N_14116,N_11879,N_8638);
or U14117 (N_14117,N_8408,N_8119);
nand U14118 (N_14118,N_9059,N_11909);
xnor U14119 (N_14119,N_9520,N_11261);
nand U14120 (N_14120,N_8616,N_7547);
nor U14121 (N_14121,N_7460,N_9892);
nand U14122 (N_14122,N_8825,N_6361);
nand U14123 (N_14123,N_7163,N_7828);
nor U14124 (N_14124,N_7469,N_6270);
xnor U14125 (N_14125,N_10878,N_11490);
and U14126 (N_14126,N_11856,N_9070);
nand U14127 (N_14127,N_7191,N_9262);
or U14128 (N_14128,N_9786,N_10108);
nor U14129 (N_14129,N_6474,N_9974);
and U14130 (N_14130,N_11770,N_8602);
or U14131 (N_14131,N_8641,N_10175);
nand U14132 (N_14132,N_7565,N_6009);
xor U14133 (N_14133,N_9604,N_8442);
nor U14134 (N_14134,N_10114,N_9494);
nor U14135 (N_14135,N_11750,N_10152);
or U14136 (N_14136,N_6723,N_9720);
xnor U14137 (N_14137,N_8384,N_7564);
and U14138 (N_14138,N_10128,N_6074);
nand U14139 (N_14139,N_8300,N_11917);
nor U14140 (N_14140,N_6095,N_9628);
nand U14141 (N_14141,N_6771,N_10846);
nor U14142 (N_14142,N_11981,N_8358);
and U14143 (N_14143,N_8378,N_11943);
nand U14144 (N_14144,N_11741,N_7138);
nor U14145 (N_14145,N_9210,N_11835);
or U14146 (N_14146,N_10687,N_10774);
nand U14147 (N_14147,N_11785,N_7684);
and U14148 (N_14148,N_10260,N_6958);
xnor U14149 (N_14149,N_6066,N_11169);
or U14150 (N_14150,N_7452,N_9618);
nand U14151 (N_14151,N_11912,N_9320);
or U14152 (N_14152,N_6894,N_11722);
and U14153 (N_14153,N_9417,N_6669);
nor U14154 (N_14154,N_8195,N_9623);
nand U14155 (N_14155,N_8685,N_9188);
xor U14156 (N_14156,N_9181,N_10845);
nand U14157 (N_14157,N_6335,N_9699);
nor U14158 (N_14158,N_6436,N_11955);
or U14159 (N_14159,N_9772,N_8750);
nor U14160 (N_14160,N_10177,N_7662);
nor U14161 (N_14161,N_11404,N_11581);
and U14162 (N_14162,N_7860,N_10343);
and U14163 (N_14163,N_10244,N_8771);
nand U14164 (N_14164,N_11427,N_7867);
nand U14165 (N_14165,N_6942,N_6409);
or U14166 (N_14166,N_7135,N_11310);
and U14167 (N_14167,N_11331,N_7344);
and U14168 (N_14168,N_10749,N_11846);
nor U14169 (N_14169,N_10029,N_7132);
nand U14170 (N_14170,N_9465,N_11678);
or U14171 (N_14171,N_7503,N_7986);
or U14172 (N_14172,N_6811,N_7707);
or U14173 (N_14173,N_9246,N_6910);
or U14174 (N_14174,N_11550,N_9509);
and U14175 (N_14175,N_6931,N_8883);
or U14176 (N_14176,N_6125,N_11474);
and U14177 (N_14177,N_10456,N_8583);
xnor U14178 (N_14178,N_6187,N_9527);
and U14179 (N_14179,N_10832,N_6597);
xor U14180 (N_14180,N_11139,N_10827);
or U14181 (N_14181,N_6523,N_11627);
xnor U14182 (N_14182,N_11180,N_7615);
nor U14183 (N_14183,N_6679,N_10155);
xor U14184 (N_14184,N_10939,N_11964);
nor U14185 (N_14185,N_6230,N_6208);
or U14186 (N_14186,N_7251,N_7730);
or U14187 (N_14187,N_9424,N_11902);
and U14188 (N_14188,N_7686,N_9073);
nor U14189 (N_14189,N_7126,N_9343);
and U14190 (N_14190,N_9841,N_8059);
and U14191 (N_14191,N_7471,N_6574);
nand U14192 (N_14192,N_8218,N_11725);
nand U14193 (N_14193,N_11790,N_9130);
or U14194 (N_14194,N_7936,N_11308);
or U14195 (N_14195,N_11458,N_6524);
or U14196 (N_14196,N_9671,N_7544);
nor U14197 (N_14197,N_11317,N_10339);
xor U14198 (N_14198,N_9305,N_10850);
nand U14199 (N_14199,N_7489,N_11365);
or U14200 (N_14200,N_10981,N_6493);
xnor U14201 (N_14201,N_6250,N_11215);
and U14202 (N_14202,N_10320,N_6051);
or U14203 (N_14203,N_6564,N_7203);
nand U14204 (N_14204,N_7574,N_10712);
and U14205 (N_14205,N_8681,N_10110);
xnor U14206 (N_14206,N_9866,N_11074);
nor U14207 (N_14207,N_7283,N_11461);
and U14208 (N_14208,N_10483,N_9228);
nor U14209 (N_14209,N_6799,N_10989);
or U14210 (N_14210,N_6319,N_7470);
or U14211 (N_14211,N_9983,N_10470);
nor U14212 (N_14212,N_8912,N_9464);
nand U14213 (N_14213,N_8260,N_10838);
xnor U14214 (N_14214,N_9393,N_9091);
xnor U14215 (N_14215,N_11115,N_11053);
and U14216 (N_14216,N_7401,N_9173);
and U14217 (N_14217,N_6399,N_6299);
or U14218 (N_14218,N_6042,N_11596);
or U14219 (N_14219,N_7315,N_6936);
or U14220 (N_14220,N_11995,N_11897);
or U14221 (N_14221,N_11791,N_8136);
nor U14222 (N_14222,N_8536,N_10627);
nor U14223 (N_14223,N_6989,N_11432);
nor U14224 (N_14224,N_9291,N_9727);
or U14225 (N_14225,N_11219,N_8373);
nor U14226 (N_14226,N_7285,N_9347);
nor U14227 (N_14227,N_7692,N_7832);
and U14228 (N_14228,N_6089,N_9905);
or U14229 (N_14229,N_6640,N_11428);
or U14230 (N_14230,N_9644,N_7060);
nor U14231 (N_14231,N_8988,N_7474);
nand U14232 (N_14232,N_10858,N_10098);
and U14233 (N_14233,N_8943,N_6430);
xnor U14234 (N_14234,N_6725,N_8740);
xnor U14235 (N_14235,N_10530,N_7625);
nor U14236 (N_14236,N_6639,N_10547);
and U14237 (N_14237,N_7174,N_8692);
or U14238 (N_14238,N_8001,N_9407);
nor U14239 (N_14239,N_11167,N_10154);
or U14240 (N_14240,N_11291,N_6126);
xnor U14241 (N_14241,N_7032,N_9558);
or U14242 (N_14242,N_9737,N_8297);
or U14243 (N_14243,N_10237,N_6838);
and U14244 (N_14244,N_9142,N_8440);
xnor U14245 (N_14245,N_10917,N_9017);
nand U14246 (N_14246,N_7124,N_10941);
nand U14247 (N_14247,N_7111,N_10792);
xnor U14248 (N_14248,N_9878,N_6714);
nor U14249 (N_14249,N_9301,N_6644);
nor U14250 (N_14250,N_10454,N_10053);
nor U14251 (N_14251,N_11604,N_9651);
or U14252 (N_14252,N_7076,N_8560);
nor U14253 (N_14253,N_10977,N_9158);
or U14254 (N_14254,N_8645,N_8178);
xnor U14255 (N_14255,N_10049,N_9149);
xor U14256 (N_14256,N_10565,N_10947);
and U14257 (N_14257,N_6147,N_7590);
or U14258 (N_14258,N_9340,N_7753);
and U14259 (N_14259,N_7681,N_6843);
or U14260 (N_14260,N_11473,N_10147);
and U14261 (N_14261,N_11294,N_6236);
nor U14262 (N_14262,N_7608,N_11292);
or U14263 (N_14263,N_8075,N_11220);
nor U14264 (N_14264,N_8211,N_11234);
xnor U14265 (N_14265,N_9123,N_9646);
or U14266 (N_14266,N_11242,N_7248);
xnor U14267 (N_14267,N_10396,N_11675);
xor U14268 (N_14268,N_8719,N_11011);
nor U14269 (N_14269,N_7020,N_6535);
nand U14270 (N_14270,N_11703,N_9971);
and U14271 (N_14271,N_7206,N_8053);
xnor U14272 (N_14272,N_9925,N_8247);
or U14273 (N_14273,N_6115,N_7679);
nor U14274 (N_14274,N_7458,N_6248);
nand U14275 (N_14275,N_10385,N_11960);
and U14276 (N_14276,N_8368,N_9533);
nand U14277 (N_14277,N_8199,N_7671);
or U14278 (N_14278,N_6528,N_6031);
xnor U14279 (N_14279,N_10368,N_9844);
and U14280 (N_14280,N_10209,N_9760);
xnor U14281 (N_14281,N_11559,N_8864);
nor U14282 (N_14282,N_7906,N_7095);
and U14283 (N_14283,N_9956,N_6791);
nand U14284 (N_14284,N_11184,N_10781);
or U14285 (N_14285,N_8534,N_6475);
or U14286 (N_14286,N_10252,N_6891);
xnor U14287 (N_14287,N_6673,N_8419);
nand U14288 (N_14288,N_7949,N_7702);
or U14289 (N_14289,N_11558,N_10784);
or U14290 (N_14290,N_6792,N_6177);
nor U14291 (N_14291,N_8389,N_7294);
or U14292 (N_14292,N_8744,N_6876);
or U14293 (N_14293,N_6648,N_8290);
nor U14294 (N_14294,N_6371,N_6440);
xnor U14295 (N_14295,N_11276,N_9256);
or U14296 (N_14296,N_7409,N_10212);
nand U14297 (N_14297,N_10624,N_7379);
nand U14298 (N_14298,N_10297,N_8021);
nand U14299 (N_14299,N_11185,N_9990);
nor U14300 (N_14300,N_10740,N_11792);
nor U14301 (N_14301,N_8250,N_9348);
and U14302 (N_14302,N_7688,N_7997);
xor U14303 (N_14303,N_7451,N_8115);
xnor U14304 (N_14304,N_10411,N_10471);
and U14305 (N_14305,N_7290,N_8121);
xor U14306 (N_14306,N_9401,N_7033);
or U14307 (N_14307,N_6228,N_7306);
nor U14308 (N_14308,N_8268,N_7947);
xnor U14309 (N_14309,N_7606,N_8839);
xnor U14310 (N_14310,N_11692,N_8173);
xor U14311 (N_14311,N_6032,N_8015);
and U14312 (N_14312,N_10116,N_7035);
xor U14313 (N_14313,N_8731,N_8323);
or U14314 (N_14314,N_6057,N_7941);
and U14315 (N_14315,N_7651,N_9500);
or U14316 (N_14316,N_8345,N_6322);
and U14317 (N_14317,N_11268,N_6991);
xnor U14318 (N_14318,N_6155,N_6674);
nor U14319 (N_14319,N_9454,N_10474);
or U14320 (N_14320,N_6005,N_6561);
or U14321 (N_14321,N_11445,N_9163);
nor U14322 (N_14322,N_9461,N_7818);
nand U14323 (N_14323,N_10261,N_9491);
nor U14324 (N_14324,N_10877,N_6755);
xor U14325 (N_14325,N_6575,N_6578);
and U14326 (N_14326,N_9529,N_7057);
nand U14327 (N_14327,N_6140,N_11029);
and U14328 (N_14328,N_8464,N_7676);
xor U14329 (N_14329,N_6652,N_9361);
xor U14330 (N_14330,N_6457,N_11057);
nand U14331 (N_14331,N_6331,N_8831);
xnor U14332 (N_14332,N_11767,N_8997);
nand U14333 (N_14333,N_8539,N_11693);
nor U14334 (N_14334,N_6207,N_11175);
nor U14335 (N_14335,N_7742,N_7802);
nor U14336 (N_14336,N_7911,N_6020);
nor U14337 (N_14337,N_6372,N_6658);
nand U14338 (N_14338,N_10927,N_8706);
xor U14339 (N_14339,N_9692,N_8277);
xor U14340 (N_14340,N_7965,N_10416);
xnor U14341 (N_14341,N_9596,N_11661);
and U14342 (N_14342,N_11842,N_10490);
xor U14343 (N_14343,N_11988,N_9439);
and U14344 (N_14344,N_11533,N_6296);
xnor U14345 (N_14345,N_6024,N_9821);
xnor U14346 (N_14346,N_7423,N_9368);
xnor U14347 (N_14347,N_8870,N_11429);
nand U14348 (N_14348,N_9083,N_8886);
xor U14349 (N_14349,N_6394,N_11340);
nor U14350 (N_14350,N_8056,N_7727);
xor U14351 (N_14351,N_8585,N_7376);
and U14352 (N_14352,N_6454,N_9161);
or U14353 (N_14353,N_8866,N_8687);
nand U14354 (N_14354,N_10783,N_9207);
nor U14355 (N_14355,N_6346,N_9341);
and U14356 (N_14356,N_8756,N_6269);
nand U14357 (N_14357,N_6717,N_9304);
nor U14358 (N_14358,N_7935,N_11459);
nor U14359 (N_14359,N_6833,N_8179);
or U14360 (N_14360,N_9303,N_8116);
nor U14361 (N_14361,N_7587,N_9823);
nor U14362 (N_14362,N_8109,N_11686);
nor U14363 (N_14363,N_11457,N_10235);
xnor U14364 (N_14364,N_11186,N_6321);
or U14365 (N_14365,N_11110,N_9893);
xnor U14366 (N_14366,N_10248,N_6824);
and U14367 (N_14367,N_10628,N_6770);
nand U14368 (N_14368,N_10768,N_7038);
or U14369 (N_14369,N_6972,N_8929);
nor U14370 (N_14370,N_6467,N_7343);
or U14371 (N_14371,N_7891,N_8402);
xnor U14372 (N_14372,N_11612,N_10659);
nand U14373 (N_14373,N_7337,N_7559);
or U14374 (N_14374,N_9943,N_9479);
or U14375 (N_14375,N_9543,N_11222);
nor U14376 (N_14376,N_10166,N_9432);
and U14377 (N_14377,N_9903,N_7484);
or U14378 (N_14378,N_10880,N_6999);
or U14379 (N_14379,N_7493,N_10478);
nand U14380 (N_14380,N_7177,N_10571);
nor U14381 (N_14381,N_8851,N_6812);
and U14382 (N_14382,N_8856,N_9136);
xnor U14383 (N_14383,N_6157,N_9536);
xor U14384 (N_14384,N_9220,N_10575);
nand U14385 (N_14385,N_7013,N_8144);
and U14386 (N_14386,N_6635,N_6739);
and U14387 (N_14387,N_6434,N_10842);
and U14388 (N_14388,N_9382,N_7219);
nor U14389 (N_14389,N_11216,N_7417);
nand U14390 (N_14390,N_7907,N_6102);
nor U14391 (N_14391,N_6131,N_11817);
xnor U14392 (N_14392,N_11161,N_6814);
nor U14393 (N_14393,N_11640,N_10812);
or U14394 (N_14394,N_10107,N_9550);
xor U14395 (N_14395,N_7515,N_7735);
and U14396 (N_14396,N_7408,N_9779);
or U14397 (N_14397,N_7444,N_7975);
xor U14398 (N_14398,N_6598,N_8342);
nor U14399 (N_14399,N_8070,N_10065);
xnor U14400 (N_14400,N_6336,N_10637);
nand U14401 (N_14401,N_7089,N_9922);
xnor U14402 (N_14402,N_9221,N_7995);
nor U14403 (N_14403,N_8046,N_9169);
nand U14404 (N_14404,N_10094,N_9762);
or U14405 (N_14405,N_7381,N_10646);
nand U14406 (N_14406,N_7043,N_10251);
nand U14407 (N_14407,N_8793,N_7526);
nor U14408 (N_14408,N_11218,N_8991);
or U14409 (N_14409,N_9420,N_9328);
nand U14410 (N_14410,N_10207,N_11641);
or U14411 (N_14411,N_10905,N_8210);
nand U14412 (N_14412,N_10197,N_7277);
nor U14413 (N_14413,N_9617,N_11871);
nand U14414 (N_14414,N_8902,N_11891);
nor U14415 (N_14415,N_6907,N_8882);
or U14416 (N_14416,N_10976,N_7357);
nand U14417 (N_14417,N_7717,N_7801);
nand U14418 (N_14418,N_11560,N_9801);
and U14419 (N_14419,N_8155,N_7394);
and U14420 (N_14420,N_8474,N_10726);
or U14421 (N_14421,N_11043,N_7859);
xnor U14422 (N_14422,N_9557,N_7179);
and U14423 (N_14423,N_10253,N_9585);
xnor U14424 (N_14424,N_11036,N_10623);
and U14425 (N_14425,N_7424,N_7642);
or U14426 (N_14426,N_7924,N_9013);
or U14427 (N_14427,N_10560,N_6675);
or U14428 (N_14428,N_8605,N_11551);
or U14429 (N_14429,N_11720,N_8298);
nand U14430 (N_14430,N_10923,N_9381);
nand U14431 (N_14431,N_7550,N_10034);
nand U14432 (N_14432,N_8493,N_8270);
nor U14433 (N_14433,N_6641,N_11574);
or U14434 (N_14434,N_10052,N_8711);
or U14435 (N_14435,N_8562,N_9564);
xnor U14436 (N_14436,N_9775,N_11860);
xnor U14437 (N_14437,N_8639,N_7957);
nand U14438 (N_14438,N_10011,N_6061);
xor U14439 (N_14439,N_10703,N_9825);
nand U14440 (N_14440,N_11398,N_11872);
or U14441 (N_14441,N_10215,N_6174);
and U14442 (N_14442,N_9900,N_6947);
nand U14443 (N_14443,N_9333,N_6716);
or U14444 (N_14444,N_8188,N_10265);
or U14445 (N_14445,N_6469,N_10449);
or U14446 (N_14446,N_9107,N_9988);
nor U14447 (N_14447,N_10993,N_11224);
and U14448 (N_14448,N_8333,N_7210);
nor U14449 (N_14449,N_9200,N_11769);
or U14450 (N_14450,N_8829,N_10169);
and U14451 (N_14451,N_7598,N_8158);
and U14452 (N_14452,N_9799,N_8203);
nor U14453 (N_14453,N_7445,N_9350);
xor U14454 (N_14454,N_8852,N_8567);
nand U14455 (N_14455,N_8975,N_10843);
or U14456 (N_14456,N_8289,N_8816);
nor U14457 (N_14457,N_7910,N_7416);
nor U14458 (N_14458,N_11811,N_10307);
xnor U14459 (N_14459,N_6404,N_7143);
nor U14460 (N_14460,N_8191,N_9868);
or U14461 (N_14461,N_9680,N_7311);
nor U14462 (N_14462,N_8018,N_11510);
or U14463 (N_14463,N_8670,N_6775);
or U14464 (N_14464,N_9496,N_6626);
or U14465 (N_14465,N_10708,N_8409);
xor U14466 (N_14466,N_7584,N_8008);
nor U14467 (N_14467,N_11638,N_11106);
or U14468 (N_14468,N_8231,N_7996);
xor U14469 (N_14469,N_11714,N_7749);
or U14470 (N_14470,N_11006,N_10568);
nor U14471 (N_14471,N_9812,N_9269);
and U14472 (N_14472,N_9419,N_9929);
or U14473 (N_14473,N_7512,N_6307);
or U14474 (N_14474,N_7021,N_10540);
xor U14475 (N_14475,N_6806,N_7817);
or U14476 (N_14476,N_11296,N_11202);
and U14477 (N_14477,N_11565,N_8564);
nor U14478 (N_14478,N_11546,N_9894);
nand U14479 (N_14479,N_9093,N_9850);
nor U14480 (N_14480,N_11919,N_9814);
xnor U14481 (N_14481,N_8727,N_8201);
or U14482 (N_14482,N_10123,N_6823);
xor U14483 (N_14483,N_10134,N_6607);
and U14484 (N_14484,N_7280,N_10675);
and U14485 (N_14485,N_8614,N_10321);
nor U14486 (N_14486,N_10238,N_9649);
or U14487 (N_14487,N_11433,N_7570);
and U14488 (N_14488,N_6292,N_6144);
nor U14489 (N_14489,N_7372,N_10202);
nor U14490 (N_14490,N_7840,N_8993);
xor U14491 (N_14491,N_6166,N_10113);
and U14492 (N_14492,N_7678,N_8024);
xor U14493 (N_14493,N_10301,N_9621);
xnor U14494 (N_14494,N_10896,N_6013);
nand U14495 (N_14495,N_10336,N_7724);
nand U14496 (N_14496,N_9541,N_10520);
xnor U14497 (N_14497,N_10763,N_8356);
or U14498 (N_14498,N_9373,N_8030);
and U14499 (N_14499,N_6820,N_9701);
and U14500 (N_14500,N_7582,N_10270);
xor U14501 (N_14501,N_9544,N_10281);
xor U14502 (N_14502,N_6018,N_7714);
xor U14503 (N_14503,N_10132,N_9076);
xnor U14504 (N_14504,N_9745,N_11060);
and U14505 (N_14505,N_8038,N_9657);
xor U14506 (N_14506,N_8569,N_8141);
xnor U14507 (N_14507,N_9908,N_11554);
or U14508 (N_14508,N_9836,N_11673);
and U14509 (N_14509,N_9522,N_6494);
and U14510 (N_14510,N_10681,N_9576);
nor U14511 (N_14511,N_8892,N_8729);
and U14512 (N_14512,N_7491,N_8503);
and U14513 (N_14513,N_10728,N_7862);
nand U14514 (N_14514,N_6783,N_8093);
nor U14515 (N_14515,N_11653,N_11821);
xnor U14516 (N_14516,N_11148,N_9700);
and U14517 (N_14517,N_10174,N_10916);
xor U14518 (N_14518,N_7628,N_8167);
nor U14519 (N_14519,N_9075,N_8162);
and U14520 (N_14520,N_6491,N_7530);
or U14521 (N_14521,N_6601,N_7948);
and U14522 (N_14522,N_6769,N_6571);
and U14523 (N_14523,N_6086,N_11699);
xor U14524 (N_14524,N_10744,N_11484);
or U14525 (N_14525,N_8206,N_10217);
or U14526 (N_14526,N_9659,N_9225);
nor U14527 (N_14527,N_8794,N_8397);
xnor U14528 (N_14528,N_9638,N_11384);
nor U14529 (N_14529,N_8496,N_7659);
or U14530 (N_14530,N_6359,N_7585);
xor U14531 (N_14531,N_9276,N_9849);
or U14532 (N_14532,N_10272,N_6364);
or U14533 (N_14533,N_11034,N_10539);
and U14534 (N_14534,N_7336,N_6468);
nand U14535 (N_14535,N_8222,N_7082);
or U14536 (N_14536,N_8734,N_9539);
or U14537 (N_14537,N_6151,N_9577);
xnor U14538 (N_14538,N_9074,N_6550);
xnor U14539 (N_14539,N_7725,N_6341);
nor U14540 (N_14540,N_11852,N_11583);
and U14541 (N_14541,N_9870,N_10284);
xnor U14542 (N_14542,N_10340,N_8334);
or U14543 (N_14543,N_9264,N_9311);
and U14544 (N_14544,N_11452,N_6547);
nor U14545 (N_14545,N_7046,N_6424);
xor U14546 (N_14546,N_8930,N_9886);
nand U14547 (N_14547,N_8592,N_10953);
or U14548 (N_14548,N_11447,N_6310);
xnor U14549 (N_14549,N_9476,N_7249);
xnor U14550 (N_14550,N_8000,N_11118);
or U14551 (N_14551,N_7534,N_8956);
and U14552 (N_14552,N_9750,N_11709);
nand U14553 (N_14553,N_10979,N_8518);
or U14554 (N_14554,N_10293,N_8291);
and U14555 (N_14555,N_8259,N_6314);
or U14556 (N_14556,N_8207,N_8984);
xor U14557 (N_14557,N_10310,N_6877);
xor U14558 (N_14558,N_7708,N_6745);
nor U14559 (N_14559,N_9041,N_8236);
and U14560 (N_14560,N_8060,N_9444);
xor U14561 (N_14561,N_11381,N_7566);
nand U14562 (N_14562,N_6049,N_9194);
nor U14563 (N_14563,N_10873,N_7744);
or U14564 (N_14564,N_9218,N_10439);
and U14565 (N_14565,N_6438,N_7588);
or U14566 (N_14566,N_8716,N_11665);
nand U14567 (N_14567,N_11312,N_6707);
nand U14568 (N_14568,N_11062,N_10485);
nand U14569 (N_14569,N_8506,N_7475);
nor U14570 (N_14570,N_9735,N_9029);
nand U14571 (N_14571,N_10521,N_9037);
xnor U14572 (N_14572,N_9822,N_9066);
or U14573 (N_14573,N_8720,N_6829);
nor U14574 (N_14574,N_9723,N_7780);
and U14575 (N_14575,N_11633,N_6355);
and U14576 (N_14576,N_9441,N_11374);
nand U14577 (N_14577,N_7864,N_8927);
and U14578 (N_14578,N_7331,N_10377);
xor U14579 (N_14579,N_8415,N_8486);
nand U14580 (N_14580,N_7963,N_11828);
or U14581 (N_14581,N_8437,N_7718);
nor U14582 (N_14582,N_7437,N_10820);
nand U14583 (N_14583,N_8588,N_7938);
nand U14584 (N_14584,N_7845,N_7520);
xor U14585 (N_14585,N_9426,N_7893);
nor U14586 (N_14586,N_7097,N_8372);
nand U14587 (N_14587,N_9965,N_7305);
or U14588 (N_14588,N_11178,N_6465);
xnor U14589 (N_14589,N_6503,N_7120);
and U14590 (N_14590,N_11371,N_7805);
nor U14591 (N_14591,N_6379,N_8355);
xnor U14592 (N_14592,N_8246,N_8340);
xor U14593 (N_14593,N_9726,N_8365);
nor U14594 (N_14594,N_9686,N_6677);
xor U14595 (N_14595,N_7695,N_11197);
xor U14596 (N_14596,N_9112,N_6854);
nand U14597 (N_14597,N_10532,N_6403);
or U14598 (N_14598,N_7202,N_10831);
xnor U14599 (N_14599,N_9645,N_6612);
xnor U14600 (N_14600,N_7816,N_6446);
and U14601 (N_14601,N_6384,N_7777);
nor U14602 (N_14602,N_9566,N_7618);
nor U14603 (N_14603,N_9230,N_8726);
xnor U14604 (N_14604,N_8940,N_8480);
nand U14605 (N_14605,N_11647,N_8996);
nor U14606 (N_14606,N_8722,N_9057);
nand U14607 (N_14607,N_6114,N_6954);
and U14608 (N_14608,N_10997,N_6984);
xnor U14609 (N_14609,N_10105,N_11645);
or U14610 (N_14610,N_11366,N_7808);
nor U14611 (N_14611,N_8090,N_11977);
and U14612 (N_14612,N_10370,N_10944);
xor U14613 (N_14613,N_6883,N_11789);
or U14614 (N_14614,N_7147,N_9431);
nor U14615 (N_14615,N_11630,N_9613);
xnor U14616 (N_14616,N_7704,N_8391);
or U14617 (N_14617,N_11342,N_7882);
nand U14618 (N_14618,N_6224,N_9826);
or U14619 (N_14619,N_9227,N_10039);
xnor U14620 (N_14620,N_10855,N_9412);
and U14621 (N_14621,N_11355,N_7105);
and U14622 (N_14622,N_6912,N_10130);
nor U14623 (N_14623,N_8642,N_11440);
nor U14624 (N_14624,N_7366,N_10504);
and U14625 (N_14625,N_11083,N_9964);
nor U14626 (N_14626,N_10443,N_8910);
and U14627 (N_14627,N_7028,N_7600);
and U14628 (N_14628,N_6283,N_7578);
xor U14629 (N_14629,N_7171,N_9941);
nor U14630 (N_14630,N_11798,N_8776);
xnor U14631 (N_14631,N_7555,N_9586);
and U14632 (N_14632,N_11980,N_11394);
or U14633 (N_14633,N_7108,N_11947);
xor U14634 (N_14634,N_8842,N_9238);
or U14635 (N_14635,N_8095,N_7647);
nand U14636 (N_14636,N_10119,N_7836);
nand U14637 (N_14637,N_9436,N_11730);
nor U14638 (N_14638,N_9640,N_9069);
and U14639 (N_14639,N_11952,N_10497);
and U14640 (N_14640,N_7400,N_9290);
nand U14641 (N_14641,N_11468,N_9402);
nor U14642 (N_14642,N_6243,N_6214);
nor U14643 (N_14643,N_9802,N_7338);
and U14644 (N_14644,N_10839,N_10918);
and U14645 (N_14645,N_9007,N_11438);
nor U14646 (N_14646,N_7232,N_10574);
xor U14647 (N_14647,N_10013,N_7266);
and U14648 (N_14648,N_7970,N_9501);
nand U14649 (N_14649,N_11921,N_8548);
and U14650 (N_14650,N_6664,N_6327);
and U14651 (N_14651,N_8694,N_8944);
nor U14652 (N_14652,N_8688,N_8051);
and U14653 (N_14653,N_11504,N_7075);
nor U14654 (N_14654,N_6240,N_7869);
xnor U14655 (N_14655,N_7347,N_11975);
and U14656 (N_14656,N_9838,N_6130);
xnor U14657 (N_14657,N_10955,N_11588);
and U14658 (N_14658,N_6232,N_7531);
or U14659 (N_14659,N_10256,N_7988);
and U14660 (N_14660,N_6263,N_11867);
xor U14661 (N_14661,N_11361,N_11945);
nor U14662 (N_14662,N_9384,N_7773);
nand U14663 (N_14663,N_6428,N_7809);
and U14664 (N_14664,N_11448,N_11067);
xnor U14665 (N_14665,N_8819,N_7011);
xor U14666 (N_14666,N_6422,N_8998);
or U14667 (N_14667,N_8968,N_6938);
or U14668 (N_14668,N_11642,N_10710);
and U14669 (N_14669,N_9202,N_9216);
xor U14670 (N_14670,N_8677,N_11302);
nand U14671 (N_14671,N_7429,N_6366);
or U14672 (N_14672,N_10428,N_9172);
or U14673 (N_14673,N_8671,N_6901);
and U14674 (N_14674,N_11840,N_8945);
or U14675 (N_14675,N_6122,N_9231);
or U14676 (N_14676,N_11961,N_9235);
and U14677 (N_14677,N_7358,N_10365);
nand U14678 (N_14678,N_11850,N_9732);
nand U14679 (N_14679,N_11781,N_7916);
and U14680 (N_14680,N_7811,N_6804);
or U14681 (N_14681,N_6767,N_11729);
or U14682 (N_14682,N_10826,N_9144);
and U14683 (N_14683,N_11700,N_10201);
xnor U14684 (N_14684,N_7276,N_10936);
or U14685 (N_14685,N_8468,N_9153);
nor U14686 (N_14686,N_7726,N_10060);
or U14687 (N_14687,N_11387,N_9477);
nor U14688 (N_14688,N_10872,N_10567);
nand U14689 (N_14689,N_10849,N_10469);
nand U14690 (N_14690,N_8275,N_10346);
and U14691 (N_14691,N_7682,N_7557);
nor U14692 (N_14692,N_6724,N_6569);
and U14693 (N_14693,N_9100,N_8017);
nand U14694 (N_14694,N_11930,N_11232);
nor U14695 (N_14695,N_9261,N_7814);
nand U14696 (N_14696,N_6067,N_8156);
nand U14697 (N_14697,N_7645,N_11549);
and U14698 (N_14698,N_10407,N_6871);
xnor U14699 (N_14699,N_9676,N_7054);
nor U14700 (N_14700,N_9534,N_7738);
nand U14701 (N_14701,N_9967,N_10773);
nor U14702 (N_14702,N_6152,N_9834);
and U14703 (N_14703,N_6990,N_8061);
or U14704 (N_14704,N_10558,N_9763);
xor U14705 (N_14705,N_8986,N_7371);
or U14706 (N_14706,N_6589,N_10044);
or U14707 (N_14707,N_6276,N_9234);
xnor U14708 (N_14708,N_7509,N_10494);
and U14709 (N_14709,N_6911,N_6090);
xor U14710 (N_14710,N_8454,N_6365);
xor U14711 (N_14711,N_7844,N_10631);
xnor U14712 (N_14712,N_8479,N_10267);
or U14713 (N_14713,N_6581,N_11843);
or U14714 (N_14714,N_8989,N_11446);
or U14715 (N_14715,N_9403,N_11058);
or U14716 (N_14716,N_11992,N_11262);
xnor U14717 (N_14717,N_10587,N_11046);
xor U14718 (N_14718,N_11485,N_7861);
or U14719 (N_14719,N_8057,N_8976);
xor U14720 (N_14720,N_9848,N_6585);
nor U14721 (N_14721,N_6815,N_6507);
xnor U14722 (N_14722,N_11258,N_7295);
and U14723 (N_14723,N_7031,N_11582);
nand U14724 (N_14724,N_7255,N_9880);
or U14725 (N_14725,N_9798,N_6279);
nand U14726 (N_14726,N_10472,N_10619);
xnor U14727 (N_14727,N_6274,N_7188);
or U14728 (N_14728,N_11179,N_7586);
xor U14729 (N_14729,N_9752,N_8375);
nor U14730 (N_14730,N_9437,N_11963);
xor U14731 (N_14731,N_8238,N_11026);
nor U14732 (N_14732,N_9022,N_8822);
nor U14733 (N_14733,N_9876,N_11492);
nor U14734 (N_14734,N_11676,N_10390);
and U14735 (N_14735,N_11865,N_8089);
or U14736 (N_14736,N_8390,N_9374);
xor U14737 (N_14737,N_8742,N_10395);
nor U14738 (N_14738,N_6345,N_10802);
and U14739 (N_14739,N_7278,N_9288);
nand U14740 (N_14740,N_11745,N_9839);
nand U14741 (N_14741,N_6553,N_9661);
and U14742 (N_14742,N_7384,N_10503);
nand U14743 (N_14743,N_9193,N_11278);
nand U14744 (N_14744,N_9663,N_11393);
or U14745 (N_14745,N_9081,N_9559);
or U14746 (N_14746,N_10461,N_8461);
xor U14747 (N_14747,N_9887,N_9026);
or U14748 (N_14748,N_7760,N_9871);
or U14749 (N_14749,N_10404,N_10970);
or U14750 (N_14750,N_11607,N_6398);
and U14751 (N_14751,N_8276,N_6171);
or U14752 (N_14752,N_8303,N_8855);
or U14753 (N_14753,N_7022,N_11668);
or U14754 (N_14754,N_9736,N_8013);
nor U14755 (N_14755,N_6868,N_6159);
or U14756 (N_14756,N_10388,N_10971);
or U14757 (N_14757,N_7723,N_7329);
or U14758 (N_14758,N_7535,N_8597);
nor U14759 (N_14759,N_9512,N_11566);
nand U14760 (N_14760,N_8311,N_6779);
or U14761 (N_14761,N_8130,N_8331);
xor U14762 (N_14762,N_10967,N_11059);
and U14763 (N_14763,N_11159,N_7396);
nor U14764 (N_14764,N_6944,N_7741);
nor U14765 (N_14765,N_10080,N_9240);
and U14766 (N_14766,N_7994,N_11289);
nor U14767 (N_14767,N_10689,N_9624);
nand U14768 (N_14768,N_11536,N_11998);
and U14769 (N_14769,N_11191,N_8223);
nor U14770 (N_14770,N_7187,N_7685);
and U14771 (N_14771,N_7765,N_8438);
and U14772 (N_14772,N_11344,N_10743);
and U14773 (N_14773,N_11316,N_6003);
xor U14774 (N_14774,N_10362,N_7349);
or U14775 (N_14775,N_9296,N_6568);
xnor U14776 (N_14776,N_6395,N_6002);
nand U14777 (N_14777,N_9082,N_10424);
or U14778 (N_14778,N_10518,N_9299);
and U14779 (N_14779,N_7088,N_7962);
nand U14780 (N_14780,N_9166,N_10786);
nor U14781 (N_14781,N_10038,N_8302);
xnor U14782 (N_14782,N_11704,N_6069);
xnor U14783 (N_14783,N_10288,N_6700);
or U14784 (N_14784,N_9045,N_7775);
xnor U14785 (N_14785,N_6760,N_7405);
nor U14786 (N_14786,N_7335,N_11519);
or U14787 (N_14787,N_6338,N_9605);
nor U14788 (N_14788,N_7499,N_11338);
nor U14789 (N_14789,N_10972,N_8566);
and U14790 (N_14790,N_9010,N_7806);
or U14791 (N_14791,N_10937,N_8680);
xor U14792 (N_14792,N_7952,N_6690);
and U14793 (N_14793,N_11783,N_9782);
nand U14794 (N_14794,N_8717,N_10050);
xnor U14795 (N_14795,N_10966,N_10018);
and U14796 (N_14796,N_7974,N_10282);
or U14797 (N_14797,N_10791,N_7225);
xnor U14798 (N_14798,N_10475,N_8885);
nand U14799 (N_14799,N_9916,N_10756);
nand U14800 (N_14800,N_10819,N_10409);
nor U14801 (N_14801,N_7485,N_10943);
or U14802 (N_14802,N_6305,N_7065);
xnor U14803 (N_14803,N_8911,N_9475);
xor U14804 (N_14804,N_6743,N_11265);
nand U14805 (N_14805,N_11532,N_8703);
or U14806 (N_14806,N_7317,N_9416);
xnor U14807 (N_14807,N_8497,N_10888);
or U14808 (N_14808,N_11054,N_6108);
and U14809 (N_14809,N_7694,N_6653);
or U14810 (N_14810,N_7091,N_9547);
nand U14811 (N_14811,N_6962,N_11928);
nand U14812 (N_14812,N_8578,N_9197);
and U14813 (N_14813,N_10245,N_10507);
xnor U14814 (N_14814,N_9068,N_6654);
xnor U14815 (N_14815,N_8114,N_6254);
nor U14816 (N_14816,N_8510,N_8766);
nand U14817 (N_14817,N_9601,N_9516);
or U14818 (N_14818,N_10200,N_6464);
or U14819 (N_14819,N_9430,N_7439);
nand U14820 (N_14820,N_10709,N_9138);
and U14821 (N_14821,N_7917,N_8033);
or U14822 (N_14822,N_10135,N_9884);
and U14823 (N_14823,N_6735,N_9321);
nand U14824 (N_14824,N_9523,N_9861);
or U14825 (N_14825,N_8450,N_11520);
nor U14826 (N_14826,N_11443,N_11834);
and U14827 (N_14827,N_8844,N_7774);
xnor U14828 (N_14828,N_6392,N_8733);
xor U14829 (N_14829,N_11804,N_9794);
or U14830 (N_14830,N_6979,N_11247);
nand U14831 (N_14831,N_8736,N_10707);
nand U14832 (N_14832,N_7084,N_6348);
and U14833 (N_14833,N_8073,N_10026);
or U14834 (N_14834,N_8802,N_10552);
nor U14835 (N_14835,N_7214,N_6128);
and U14836 (N_14836,N_7226,N_9266);
or U14837 (N_14837,N_10968,N_11540);
nand U14838 (N_14838,N_7745,N_10453);
or U14839 (N_14839,N_9632,N_9548);
nor U14840 (N_14840,N_7781,N_10329);
xor U14841 (N_14841,N_7351,N_9813);
and U14842 (N_14842,N_10027,N_8107);
nand U14843 (N_14843,N_10249,N_7894);
or U14844 (N_14844,N_8197,N_7880);
nor U14845 (N_14845,N_8804,N_7548);
and U14846 (N_14846,N_7508,N_9773);
nand U14847 (N_14847,N_10313,N_8459);
nor U14848 (N_14848,N_7950,N_7540);
and U14849 (N_14849,N_9787,N_6726);
nand U14850 (N_14850,N_8873,N_6853);
nor U14851 (N_14851,N_7611,N_8007);
xnor U14852 (N_14852,N_10338,N_8591);
and U14853 (N_14853,N_6817,N_9254);
and U14854 (N_14854,N_8517,N_10794);
nor U14855 (N_14855,N_6376,N_7157);
or U14856 (N_14856,N_6698,N_9035);
xor U14857 (N_14857,N_6124,N_9572);
or U14858 (N_14858,N_8963,N_7743);
or U14859 (N_14859,N_8647,N_8285);
nor U14860 (N_14860,N_9833,N_11695);
nor U14861 (N_14861,N_9612,N_9140);
nor U14862 (N_14862,N_7770,N_9860);
nand U14863 (N_14863,N_9961,N_8190);
xor U14864 (N_14864,N_8949,N_9963);
nor U14865 (N_14865,N_6720,N_11623);
nand U14866 (N_14866,N_6828,N_11779);
nand U14867 (N_14867,N_10075,N_8558);
and U14868 (N_14868,N_11063,N_6687);
and U14869 (N_14869,N_10423,N_6551);
nor U14870 (N_14870,N_7125,N_10964);
and U14871 (N_14871,N_10138,N_6084);
or U14872 (N_14872,N_6660,N_11313);
and U14873 (N_14873,N_7215,N_7921);
xor U14874 (N_14874,N_7055,N_7767);
nand U14875 (N_14875,N_6599,N_11198);
xnor U14876 (N_14876,N_9960,N_9096);
or U14877 (N_14877,N_11516,N_9047);
or U14878 (N_14878,N_6016,N_7903);
xnor U14879 (N_14879,N_10129,N_6431);
xnor U14880 (N_14880,N_7953,N_6623);
nor U14881 (N_14881,N_6412,N_7030);
nand U14882 (N_14882,N_11901,N_11636);
xnor U14883 (N_14883,N_9003,N_6813);
or U14884 (N_14884,N_6315,N_6613);
nor U14885 (N_14885,N_7155,N_8170);
nor U14886 (N_14886,N_9950,N_10638);
xor U14887 (N_14887,N_6485,N_7516);
nand U14888 (N_14888,N_11953,N_7104);
or U14889 (N_14889,N_7581,N_6100);
or U14890 (N_14890,N_8322,N_11042);
nand U14891 (N_14891,N_11927,N_7853);
and U14892 (N_14892,N_8313,N_8542);
nor U14893 (N_14893,N_10935,N_11593);
xnor U14894 (N_14894,N_8160,N_7230);
and U14895 (N_14895,N_10125,N_10347);
and U14896 (N_14896,N_11442,N_10387);
and U14897 (N_14897,N_7536,N_7879);
nand U14898 (N_14898,N_7252,N_8874);
nand U14899 (N_14899,N_6273,N_10434);
or U14900 (N_14900,N_8763,N_9209);
xor U14901 (N_14901,N_7748,N_9473);
nand U14902 (N_14902,N_6052,N_9511);
nand U14903 (N_14903,N_11407,N_11625);
and U14904 (N_14904,N_11610,N_10755);
xor U14905 (N_14905,N_10493,N_6988);
nand U14906 (N_14906,N_8126,N_8255);
nor U14907 (N_14907,N_8957,N_6567);
and U14908 (N_14908,N_11417,N_10092);
nand U14909 (N_14909,N_11070,N_10790);
or U14910 (N_14910,N_7079,N_8321);
nor U14911 (N_14911,N_10421,N_11726);
and U14912 (N_14912,N_11982,N_8637);
nor U14913 (N_14913,N_9270,N_6592);
or U14914 (N_14914,N_9139,N_6636);
and U14915 (N_14915,N_10287,N_7855);
nor U14916 (N_14916,N_9684,N_11150);
or U14917 (N_14917,N_11231,N_7139);
or U14918 (N_14918,N_8010,N_7288);
xor U14919 (N_14919,N_8475,N_8784);
and U14920 (N_14920,N_8239,N_8400);
or U14921 (N_14921,N_7161,N_6957);
nor U14922 (N_14922,N_7324,N_7098);
xnor U14923 (N_14923,N_8127,N_9300);
and U14924 (N_14924,N_10667,N_10649);
and U14925 (N_14925,N_11019,N_10165);
and U14926 (N_14926,N_6586,N_9208);
nor U14927 (N_14927,N_7719,N_7655);
nor U14928 (N_14928,N_9487,N_7514);
xnor U14929 (N_14929,N_8407,N_9926);
nor U14930 (N_14930,N_7302,N_7369);
nor U14931 (N_14931,N_11408,N_6007);
nand U14932 (N_14932,N_11592,N_9115);
or U14933 (N_14933,N_11409,N_6960);
and U14934 (N_14934,N_9816,N_11498);
or U14935 (N_14935,N_8317,N_9743);
xor U14936 (N_14936,N_6582,N_6312);
xor U14937 (N_14937,N_6982,N_7181);
nor U14938 (N_14938,N_7937,N_8101);
xnor U14939 (N_14939,N_8025,N_10621);
xor U14940 (N_14940,N_7096,N_7354);
nand U14941 (N_14941,N_6847,N_10185);
and U14942 (N_14942,N_8524,N_9352);
nor U14943 (N_14943,N_7436,N_8969);
and U14944 (N_14944,N_11500,N_9740);
xnor U14945 (N_14945,N_6445,N_6710);
and U14946 (N_14946,N_8678,N_8460);
xnor U14947 (N_14947,N_8019,N_11857);
xor U14948 (N_14948,N_10665,N_11102);
and U14949 (N_14949,N_7967,N_11024);
nand U14950 (N_14950,N_11280,N_7085);
nand U14951 (N_14951,N_10032,N_7411);
xnor U14952 (N_14952,N_6834,N_8977);
nor U14953 (N_14953,N_11032,N_9935);
and U14954 (N_14954,N_7831,N_6120);
or U14955 (N_14955,N_10593,N_11805);
and U14956 (N_14956,N_10324,N_11616);
or U14957 (N_14957,N_6974,N_11841);
and U14958 (N_14958,N_10008,N_10957);
or U14959 (N_14959,N_9549,N_10457);
or U14960 (N_14960,N_11025,N_7991);
nor U14961 (N_14961,N_9797,N_8698);
or U14962 (N_14962,N_9620,N_8072);
nor U14963 (N_14963,N_6169,N_6810);
and U14964 (N_14964,N_6969,N_7866);
nor U14965 (N_14965,N_8901,N_10438);
and U14966 (N_14966,N_11555,N_8946);
nand U14967 (N_14967,N_8328,N_11339);
and U14968 (N_14968,N_11290,N_7234);
nor U14969 (N_14969,N_7325,N_6577);
nor U14970 (N_14970,N_6316,N_7270);
and U14971 (N_14971,N_10436,N_10250);
nand U14972 (N_14972,N_7601,N_11971);
or U14973 (N_14973,N_9991,N_10959);
nor U14974 (N_14974,N_8563,N_6595);
or U14975 (N_14975,N_11315,N_10670);
and U14976 (N_14976,N_9467,N_9249);
and U14977 (N_14977,N_7983,N_11567);
nor U14978 (N_14978,N_6478,N_11985);
nand U14979 (N_14979,N_9369,N_8758);
nand U14980 (N_14980,N_9248,N_10919);
or U14981 (N_14981,N_7892,N_6495);
nand U14982 (N_14982,N_9729,N_10807);
nand U14983 (N_14983,N_6172,N_6766);
and U14984 (N_14984,N_6419,N_7254);
nor U14985 (N_14985,N_11570,N_10579);
nor U14986 (N_14986,N_10243,N_9414);
nand U14987 (N_14987,N_6277,N_7370);
or U14988 (N_14988,N_8031,N_9293);
and U14989 (N_14989,N_6373,N_10764);
nor U14990 (N_14990,N_7425,N_11906);
and U14991 (N_14991,N_6663,N_7837);
xnor U14992 (N_14992,N_11194,N_10778);
nor U14993 (N_14993,N_11476,N_10713);
or U14994 (N_14994,N_11666,N_7612);
xnor U14995 (N_14995,N_11951,N_7716);
or U14996 (N_14996,N_9837,N_7902);
xor U14997 (N_14997,N_11905,N_10059);
xor U14998 (N_14998,N_6397,N_11066);
xor U14999 (N_14999,N_11343,N_10422);
or U15000 (N_15000,N_8564,N_8784);
and U15001 (N_15001,N_6871,N_9561);
nor U15002 (N_15002,N_10789,N_7427);
xor U15003 (N_15003,N_7366,N_6108);
or U15004 (N_15004,N_11097,N_8194);
xnor U15005 (N_15005,N_7347,N_10598);
xnor U15006 (N_15006,N_8706,N_11110);
or U15007 (N_15007,N_6383,N_7493);
xnor U15008 (N_15008,N_8274,N_8588);
xnor U15009 (N_15009,N_6846,N_9577);
or U15010 (N_15010,N_9246,N_7924);
and U15011 (N_15011,N_8983,N_10747);
nand U15012 (N_15012,N_10519,N_8698);
nor U15013 (N_15013,N_7410,N_6360);
nand U15014 (N_15014,N_6602,N_7907);
nand U15015 (N_15015,N_8967,N_9548);
xnor U15016 (N_15016,N_6012,N_9764);
nor U15017 (N_15017,N_10978,N_6128);
nor U15018 (N_15018,N_8708,N_11024);
nand U15019 (N_15019,N_11538,N_9888);
or U15020 (N_15020,N_6226,N_9879);
nand U15021 (N_15021,N_11387,N_8107);
nor U15022 (N_15022,N_8187,N_6680);
nor U15023 (N_15023,N_9174,N_11530);
and U15024 (N_15024,N_11134,N_6637);
nand U15025 (N_15025,N_7181,N_8318);
and U15026 (N_15026,N_11230,N_7148);
xor U15027 (N_15027,N_7879,N_8122);
and U15028 (N_15028,N_11079,N_9441);
xor U15029 (N_15029,N_11190,N_8778);
nand U15030 (N_15030,N_10129,N_6764);
nor U15031 (N_15031,N_11024,N_8063);
and U15032 (N_15032,N_10960,N_9400);
and U15033 (N_15033,N_8364,N_7081);
and U15034 (N_15034,N_6930,N_11733);
nand U15035 (N_15035,N_6563,N_7713);
xnor U15036 (N_15036,N_11707,N_7851);
nor U15037 (N_15037,N_9790,N_10693);
xnor U15038 (N_15038,N_9860,N_11147);
and U15039 (N_15039,N_6100,N_10821);
nor U15040 (N_15040,N_7597,N_7714);
or U15041 (N_15041,N_11260,N_7211);
or U15042 (N_15042,N_6981,N_9853);
nor U15043 (N_15043,N_10422,N_10583);
nand U15044 (N_15044,N_9591,N_11228);
nand U15045 (N_15045,N_7069,N_8281);
xnor U15046 (N_15046,N_11861,N_7748);
and U15047 (N_15047,N_10789,N_8020);
and U15048 (N_15048,N_9867,N_10204);
nor U15049 (N_15049,N_8158,N_11959);
xor U15050 (N_15050,N_11476,N_10015);
nand U15051 (N_15051,N_10068,N_8360);
nor U15052 (N_15052,N_10891,N_9876);
xor U15053 (N_15053,N_9870,N_6162);
xnor U15054 (N_15054,N_9029,N_10289);
nor U15055 (N_15055,N_9026,N_9952);
nand U15056 (N_15056,N_11743,N_8774);
xnor U15057 (N_15057,N_10463,N_10697);
and U15058 (N_15058,N_9220,N_10170);
nor U15059 (N_15059,N_9866,N_7573);
or U15060 (N_15060,N_7868,N_11317);
or U15061 (N_15061,N_8059,N_8391);
nand U15062 (N_15062,N_6715,N_9465);
nor U15063 (N_15063,N_9541,N_10189);
nand U15064 (N_15064,N_7013,N_8695);
or U15065 (N_15065,N_7863,N_8806);
and U15066 (N_15066,N_9035,N_8405);
nor U15067 (N_15067,N_11983,N_6494);
or U15068 (N_15068,N_11445,N_7737);
or U15069 (N_15069,N_9056,N_6249);
nand U15070 (N_15070,N_10352,N_9373);
xor U15071 (N_15071,N_6271,N_6362);
xnor U15072 (N_15072,N_9438,N_10922);
xnor U15073 (N_15073,N_9759,N_7474);
nand U15074 (N_15074,N_10315,N_11728);
and U15075 (N_15075,N_6368,N_6865);
and U15076 (N_15076,N_10612,N_10850);
or U15077 (N_15077,N_9412,N_9703);
nor U15078 (N_15078,N_11684,N_7837);
and U15079 (N_15079,N_10248,N_10777);
xor U15080 (N_15080,N_10439,N_9850);
and U15081 (N_15081,N_10787,N_6436);
nor U15082 (N_15082,N_8549,N_9726);
or U15083 (N_15083,N_8036,N_10572);
nor U15084 (N_15084,N_9783,N_10562);
xor U15085 (N_15085,N_7329,N_9888);
nor U15086 (N_15086,N_7779,N_9327);
nand U15087 (N_15087,N_7512,N_9351);
or U15088 (N_15088,N_8659,N_8550);
or U15089 (N_15089,N_8694,N_9618);
xor U15090 (N_15090,N_8299,N_11038);
and U15091 (N_15091,N_11001,N_9003);
nor U15092 (N_15092,N_7349,N_7443);
nor U15093 (N_15093,N_8273,N_11877);
nor U15094 (N_15094,N_8786,N_10969);
and U15095 (N_15095,N_9306,N_6541);
nand U15096 (N_15096,N_9506,N_11918);
and U15097 (N_15097,N_6277,N_6136);
or U15098 (N_15098,N_10512,N_10522);
or U15099 (N_15099,N_8580,N_11201);
nor U15100 (N_15100,N_9388,N_6369);
or U15101 (N_15101,N_11078,N_9844);
nor U15102 (N_15102,N_11993,N_6398);
nor U15103 (N_15103,N_11354,N_10546);
nand U15104 (N_15104,N_8941,N_11850);
or U15105 (N_15105,N_9547,N_8225);
or U15106 (N_15106,N_9945,N_7773);
nor U15107 (N_15107,N_10171,N_6550);
or U15108 (N_15108,N_7409,N_9170);
and U15109 (N_15109,N_8394,N_8149);
or U15110 (N_15110,N_7098,N_6928);
and U15111 (N_15111,N_6939,N_10889);
xor U15112 (N_15112,N_7619,N_10604);
and U15113 (N_15113,N_9440,N_8759);
nor U15114 (N_15114,N_9637,N_9017);
and U15115 (N_15115,N_11293,N_9936);
and U15116 (N_15116,N_6591,N_7371);
or U15117 (N_15117,N_6240,N_10628);
xnor U15118 (N_15118,N_10085,N_10179);
nor U15119 (N_15119,N_8994,N_10900);
and U15120 (N_15120,N_9738,N_7536);
nor U15121 (N_15121,N_7051,N_11556);
nand U15122 (N_15122,N_9316,N_9438);
and U15123 (N_15123,N_7210,N_7525);
or U15124 (N_15124,N_9592,N_10085);
xnor U15125 (N_15125,N_6037,N_11095);
xnor U15126 (N_15126,N_9083,N_11478);
and U15127 (N_15127,N_11465,N_8642);
or U15128 (N_15128,N_6160,N_7494);
or U15129 (N_15129,N_8542,N_11004);
and U15130 (N_15130,N_9033,N_11669);
and U15131 (N_15131,N_11671,N_7352);
and U15132 (N_15132,N_8426,N_7299);
nand U15133 (N_15133,N_9304,N_11628);
or U15134 (N_15134,N_11134,N_9227);
and U15135 (N_15135,N_7990,N_7767);
or U15136 (N_15136,N_7825,N_7892);
or U15137 (N_15137,N_8693,N_11832);
nand U15138 (N_15138,N_10428,N_8132);
nand U15139 (N_15139,N_7890,N_6755);
xnor U15140 (N_15140,N_9073,N_11902);
or U15141 (N_15141,N_9587,N_10523);
xor U15142 (N_15142,N_10262,N_11477);
nand U15143 (N_15143,N_9794,N_10720);
or U15144 (N_15144,N_8941,N_6134);
nor U15145 (N_15145,N_11288,N_8096);
nor U15146 (N_15146,N_7086,N_9974);
nor U15147 (N_15147,N_6712,N_10098);
or U15148 (N_15148,N_9989,N_8477);
and U15149 (N_15149,N_11386,N_8535);
and U15150 (N_15150,N_8318,N_7309);
and U15151 (N_15151,N_8714,N_9249);
and U15152 (N_15152,N_9698,N_8089);
nor U15153 (N_15153,N_9801,N_8360);
xnor U15154 (N_15154,N_6049,N_10506);
xnor U15155 (N_15155,N_10700,N_8139);
and U15156 (N_15156,N_9933,N_7253);
or U15157 (N_15157,N_8153,N_9483);
or U15158 (N_15158,N_11850,N_6487);
nor U15159 (N_15159,N_11784,N_11704);
nor U15160 (N_15160,N_8540,N_9531);
and U15161 (N_15161,N_6634,N_8478);
nand U15162 (N_15162,N_11110,N_10855);
nor U15163 (N_15163,N_11757,N_8698);
nor U15164 (N_15164,N_9435,N_8473);
xor U15165 (N_15165,N_11658,N_8360);
or U15166 (N_15166,N_7338,N_8139);
or U15167 (N_15167,N_11549,N_7149);
nor U15168 (N_15168,N_7481,N_8067);
and U15169 (N_15169,N_9446,N_11364);
and U15170 (N_15170,N_8094,N_10795);
or U15171 (N_15171,N_7922,N_6951);
nand U15172 (N_15172,N_11147,N_6739);
nor U15173 (N_15173,N_6654,N_11480);
nor U15174 (N_15174,N_10014,N_7655);
nor U15175 (N_15175,N_8214,N_11818);
and U15176 (N_15176,N_9127,N_11955);
nand U15177 (N_15177,N_9815,N_8908);
or U15178 (N_15178,N_7810,N_8737);
nand U15179 (N_15179,N_6355,N_8078);
nand U15180 (N_15180,N_9665,N_8901);
and U15181 (N_15181,N_7115,N_10734);
nand U15182 (N_15182,N_8022,N_6045);
or U15183 (N_15183,N_11663,N_10559);
nand U15184 (N_15184,N_9166,N_6774);
and U15185 (N_15185,N_9702,N_7610);
nand U15186 (N_15186,N_10799,N_8891);
or U15187 (N_15187,N_11252,N_10485);
xor U15188 (N_15188,N_10223,N_8016);
nor U15189 (N_15189,N_6635,N_7511);
xor U15190 (N_15190,N_6847,N_9213);
nor U15191 (N_15191,N_11823,N_9197);
and U15192 (N_15192,N_10647,N_8087);
xnor U15193 (N_15193,N_9388,N_11894);
nor U15194 (N_15194,N_10033,N_8360);
nor U15195 (N_15195,N_11260,N_11345);
nor U15196 (N_15196,N_7702,N_9199);
or U15197 (N_15197,N_10485,N_10151);
xnor U15198 (N_15198,N_7712,N_7343);
nor U15199 (N_15199,N_9008,N_8824);
nand U15200 (N_15200,N_11005,N_11826);
nor U15201 (N_15201,N_8474,N_9245);
nand U15202 (N_15202,N_8980,N_10207);
nor U15203 (N_15203,N_9416,N_7310);
nand U15204 (N_15204,N_9324,N_7462);
nor U15205 (N_15205,N_7259,N_10734);
and U15206 (N_15206,N_6414,N_8547);
nand U15207 (N_15207,N_9253,N_8386);
and U15208 (N_15208,N_7266,N_9744);
nand U15209 (N_15209,N_11534,N_9529);
nand U15210 (N_15210,N_9924,N_7410);
xor U15211 (N_15211,N_7190,N_11411);
nand U15212 (N_15212,N_10600,N_6298);
nor U15213 (N_15213,N_10971,N_10238);
and U15214 (N_15214,N_7194,N_7540);
nor U15215 (N_15215,N_10155,N_11849);
or U15216 (N_15216,N_9198,N_9894);
and U15217 (N_15217,N_10559,N_10518);
nand U15218 (N_15218,N_9209,N_10050);
nor U15219 (N_15219,N_11990,N_10885);
xnor U15220 (N_15220,N_9972,N_6632);
nand U15221 (N_15221,N_10784,N_6403);
xor U15222 (N_15222,N_8955,N_10102);
nand U15223 (N_15223,N_7765,N_11554);
nor U15224 (N_15224,N_6711,N_6464);
nor U15225 (N_15225,N_10835,N_10048);
and U15226 (N_15226,N_6901,N_10681);
and U15227 (N_15227,N_11076,N_11029);
xor U15228 (N_15228,N_10622,N_7837);
xnor U15229 (N_15229,N_6830,N_6087);
nand U15230 (N_15230,N_11318,N_9501);
and U15231 (N_15231,N_9245,N_8035);
nand U15232 (N_15232,N_9719,N_6413);
and U15233 (N_15233,N_10541,N_9843);
nor U15234 (N_15234,N_6081,N_11122);
nor U15235 (N_15235,N_9910,N_9141);
xor U15236 (N_15236,N_7769,N_9545);
nand U15237 (N_15237,N_7322,N_9342);
nand U15238 (N_15238,N_9202,N_8412);
nand U15239 (N_15239,N_7843,N_8484);
nand U15240 (N_15240,N_6478,N_8200);
or U15241 (N_15241,N_11407,N_10506);
and U15242 (N_15242,N_7155,N_10718);
xnor U15243 (N_15243,N_7349,N_8543);
xnor U15244 (N_15244,N_10101,N_8788);
nor U15245 (N_15245,N_10017,N_7012);
nand U15246 (N_15246,N_7509,N_8738);
or U15247 (N_15247,N_11898,N_11997);
xor U15248 (N_15248,N_8004,N_11308);
nor U15249 (N_15249,N_10975,N_8195);
or U15250 (N_15250,N_10385,N_6103);
and U15251 (N_15251,N_8933,N_6081);
and U15252 (N_15252,N_8597,N_10646);
or U15253 (N_15253,N_10856,N_6954);
xnor U15254 (N_15254,N_9752,N_9081);
nand U15255 (N_15255,N_9747,N_7467);
nor U15256 (N_15256,N_9901,N_7253);
xnor U15257 (N_15257,N_10871,N_8581);
or U15258 (N_15258,N_7686,N_7666);
nor U15259 (N_15259,N_6793,N_8432);
nand U15260 (N_15260,N_10295,N_10301);
or U15261 (N_15261,N_10790,N_6931);
xor U15262 (N_15262,N_6576,N_8835);
nor U15263 (N_15263,N_8978,N_10214);
nand U15264 (N_15264,N_9141,N_9835);
and U15265 (N_15265,N_10584,N_10302);
xnor U15266 (N_15266,N_8561,N_8552);
and U15267 (N_15267,N_10127,N_7119);
nor U15268 (N_15268,N_9792,N_8620);
and U15269 (N_15269,N_9539,N_10711);
nor U15270 (N_15270,N_7496,N_6807);
xor U15271 (N_15271,N_11451,N_7401);
or U15272 (N_15272,N_9646,N_8609);
xor U15273 (N_15273,N_7321,N_9622);
and U15274 (N_15274,N_7034,N_10372);
or U15275 (N_15275,N_7141,N_10378);
nor U15276 (N_15276,N_9441,N_7257);
xnor U15277 (N_15277,N_9144,N_9317);
nor U15278 (N_15278,N_10809,N_10750);
nand U15279 (N_15279,N_9788,N_8629);
xor U15280 (N_15280,N_9418,N_8617);
nand U15281 (N_15281,N_7003,N_9140);
nand U15282 (N_15282,N_9467,N_8723);
and U15283 (N_15283,N_8805,N_6744);
xnor U15284 (N_15284,N_7677,N_8989);
and U15285 (N_15285,N_10333,N_7082);
xor U15286 (N_15286,N_6621,N_9728);
nand U15287 (N_15287,N_7694,N_8595);
nor U15288 (N_15288,N_6781,N_10712);
nor U15289 (N_15289,N_10002,N_9784);
and U15290 (N_15290,N_6765,N_7884);
nand U15291 (N_15291,N_11396,N_9981);
nor U15292 (N_15292,N_10147,N_9126);
xnor U15293 (N_15293,N_7193,N_7130);
or U15294 (N_15294,N_11022,N_7410);
or U15295 (N_15295,N_6719,N_8692);
nor U15296 (N_15296,N_7277,N_11419);
nor U15297 (N_15297,N_10246,N_9000);
nor U15298 (N_15298,N_6514,N_6855);
and U15299 (N_15299,N_10086,N_6044);
nand U15300 (N_15300,N_8837,N_8043);
and U15301 (N_15301,N_10634,N_9297);
nor U15302 (N_15302,N_6481,N_8275);
or U15303 (N_15303,N_9838,N_10655);
nor U15304 (N_15304,N_6191,N_9446);
nor U15305 (N_15305,N_10948,N_8880);
or U15306 (N_15306,N_6321,N_10349);
nor U15307 (N_15307,N_7957,N_6901);
nor U15308 (N_15308,N_8650,N_10357);
nand U15309 (N_15309,N_8388,N_8853);
nand U15310 (N_15310,N_10222,N_8664);
nor U15311 (N_15311,N_9157,N_9656);
nor U15312 (N_15312,N_7493,N_9147);
nand U15313 (N_15313,N_7767,N_11872);
xor U15314 (N_15314,N_9697,N_10820);
xor U15315 (N_15315,N_6647,N_6077);
nand U15316 (N_15316,N_10851,N_8656);
nand U15317 (N_15317,N_10367,N_10087);
nand U15318 (N_15318,N_10880,N_8573);
and U15319 (N_15319,N_11323,N_11562);
nor U15320 (N_15320,N_10862,N_8282);
xor U15321 (N_15321,N_7392,N_8299);
xor U15322 (N_15322,N_6583,N_8140);
or U15323 (N_15323,N_8026,N_8396);
nor U15324 (N_15324,N_9811,N_10883);
nor U15325 (N_15325,N_6062,N_9992);
and U15326 (N_15326,N_9419,N_9096);
xnor U15327 (N_15327,N_6209,N_7983);
xor U15328 (N_15328,N_6050,N_7400);
nor U15329 (N_15329,N_6889,N_6572);
and U15330 (N_15330,N_9734,N_9149);
nand U15331 (N_15331,N_7886,N_9416);
nor U15332 (N_15332,N_9613,N_10708);
nor U15333 (N_15333,N_10508,N_9292);
and U15334 (N_15334,N_11220,N_11575);
xnor U15335 (N_15335,N_6312,N_11107);
xnor U15336 (N_15336,N_7732,N_11066);
nor U15337 (N_15337,N_10794,N_8146);
xor U15338 (N_15338,N_8246,N_7724);
nand U15339 (N_15339,N_9300,N_6698);
and U15340 (N_15340,N_9916,N_11070);
nand U15341 (N_15341,N_7757,N_7192);
or U15342 (N_15342,N_6596,N_6972);
nor U15343 (N_15343,N_6403,N_8646);
nand U15344 (N_15344,N_6960,N_10912);
nor U15345 (N_15345,N_10193,N_9290);
nand U15346 (N_15346,N_6341,N_8240);
nand U15347 (N_15347,N_10424,N_6359);
nand U15348 (N_15348,N_9266,N_9398);
xor U15349 (N_15349,N_11515,N_9079);
nand U15350 (N_15350,N_7431,N_6716);
and U15351 (N_15351,N_9521,N_8983);
xor U15352 (N_15352,N_8572,N_6006);
and U15353 (N_15353,N_9001,N_10738);
nand U15354 (N_15354,N_10106,N_6250);
nand U15355 (N_15355,N_8314,N_10493);
xor U15356 (N_15356,N_9284,N_9958);
xnor U15357 (N_15357,N_7617,N_7992);
nand U15358 (N_15358,N_7611,N_7114);
xor U15359 (N_15359,N_10251,N_9197);
or U15360 (N_15360,N_9968,N_8023);
and U15361 (N_15361,N_8259,N_10607);
and U15362 (N_15362,N_10988,N_11024);
nor U15363 (N_15363,N_7650,N_9533);
nor U15364 (N_15364,N_6875,N_9480);
and U15365 (N_15365,N_8005,N_11155);
nand U15366 (N_15366,N_7013,N_8663);
xor U15367 (N_15367,N_6822,N_11108);
xor U15368 (N_15368,N_6439,N_7710);
nor U15369 (N_15369,N_9341,N_8110);
xor U15370 (N_15370,N_9827,N_6982);
and U15371 (N_15371,N_7444,N_10761);
or U15372 (N_15372,N_10675,N_8901);
or U15373 (N_15373,N_10262,N_11844);
and U15374 (N_15374,N_10080,N_6666);
nor U15375 (N_15375,N_10271,N_7356);
xor U15376 (N_15376,N_9575,N_8959);
nor U15377 (N_15377,N_8143,N_7942);
xor U15378 (N_15378,N_10668,N_10847);
or U15379 (N_15379,N_8086,N_7015);
and U15380 (N_15380,N_8962,N_6450);
xnor U15381 (N_15381,N_11112,N_11460);
xor U15382 (N_15382,N_6662,N_9942);
xnor U15383 (N_15383,N_7977,N_11826);
nand U15384 (N_15384,N_9146,N_10694);
nor U15385 (N_15385,N_9202,N_7519);
nand U15386 (N_15386,N_10705,N_8049);
nand U15387 (N_15387,N_8162,N_6314);
and U15388 (N_15388,N_8417,N_11132);
nand U15389 (N_15389,N_10145,N_9660);
nor U15390 (N_15390,N_6067,N_10886);
xor U15391 (N_15391,N_9468,N_9592);
and U15392 (N_15392,N_11828,N_6152);
nand U15393 (N_15393,N_8335,N_7364);
and U15394 (N_15394,N_7744,N_9678);
and U15395 (N_15395,N_10212,N_7718);
nor U15396 (N_15396,N_9068,N_6887);
and U15397 (N_15397,N_8882,N_7836);
and U15398 (N_15398,N_11644,N_6025);
or U15399 (N_15399,N_8405,N_11037);
xor U15400 (N_15400,N_11794,N_10983);
nor U15401 (N_15401,N_11019,N_11492);
and U15402 (N_15402,N_8238,N_7016);
and U15403 (N_15403,N_6110,N_6541);
xnor U15404 (N_15404,N_8351,N_7451);
nor U15405 (N_15405,N_6808,N_9233);
nand U15406 (N_15406,N_6295,N_9774);
nand U15407 (N_15407,N_11008,N_7376);
or U15408 (N_15408,N_9557,N_6052);
and U15409 (N_15409,N_10152,N_11640);
and U15410 (N_15410,N_8238,N_9721);
nand U15411 (N_15411,N_11941,N_11688);
nor U15412 (N_15412,N_6061,N_10536);
or U15413 (N_15413,N_7044,N_7495);
nand U15414 (N_15414,N_9368,N_6010);
and U15415 (N_15415,N_8953,N_8502);
nand U15416 (N_15416,N_10693,N_8940);
nor U15417 (N_15417,N_8662,N_11187);
nor U15418 (N_15418,N_10756,N_8042);
nand U15419 (N_15419,N_8718,N_7194);
and U15420 (N_15420,N_11225,N_11770);
nand U15421 (N_15421,N_11456,N_11704);
or U15422 (N_15422,N_9384,N_8258);
xnor U15423 (N_15423,N_8671,N_6185);
xor U15424 (N_15424,N_11038,N_11000);
xor U15425 (N_15425,N_8376,N_7458);
and U15426 (N_15426,N_9212,N_9676);
nand U15427 (N_15427,N_10347,N_10259);
nand U15428 (N_15428,N_10004,N_9344);
and U15429 (N_15429,N_11113,N_9456);
nand U15430 (N_15430,N_7402,N_8994);
nor U15431 (N_15431,N_8345,N_7473);
nand U15432 (N_15432,N_8890,N_9992);
xnor U15433 (N_15433,N_6766,N_6121);
nor U15434 (N_15434,N_6528,N_9141);
nor U15435 (N_15435,N_8349,N_9860);
xnor U15436 (N_15436,N_10421,N_11886);
and U15437 (N_15437,N_11718,N_7042);
and U15438 (N_15438,N_11138,N_6981);
or U15439 (N_15439,N_6032,N_11935);
nor U15440 (N_15440,N_6939,N_11457);
or U15441 (N_15441,N_6580,N_11382);
nor U15442 (N_15442,N_10501,N_9614);
or U15443 (N_15443,N_6112,N_11925);
xor U15444 (N_15444,N_8271,N_11226);
nand U15445 (N_15445,N_11325,N_8000);
xnor U15446 (N_15446,N_8357,N_8833);
xnor U15447 (N_15447,N_9841,N_9969);
nand U15448 (N_15448,N_9462,N_9751);
nor U15449 (N_15449,N_11918,N_11424);
nor U15450 (N_15450,N_6019,N_6264);
nor U15451 (N_15451,N_10738,N_6213);
xor U15452 (N_15452,N_8670,N_6608);
xor U15453 (N_15453,N_11381,N_8146);
or U15454 (N_15454,N_10525,N_6199);
nor U15455 (N_15455,N_7272,N_11983);
nand U15456 (N_15456,N_10326,N_8295);
and U15457 (N_15457,N_7929,N_9136);
or U15458 (N_15458,N_8170,N_6327);
and U15459 (N_15459,N_7905,N_11663);
xor U15460 (N_15460,N_7837,N_11928);
nand U15461 (N_15461,N_9919,N_7076);
nor U15462 (N_15462,N_8821,N_6544);
xor U15463 (N_15463,N_9699,N_8896);
nand U15464 (N_15464,N_9781,N_8635);
nand U15465 (N_15465,N_11550,N_6200);
nor U15466 (N_15466,N_11414,N_9267);
nand U15467 (N_15467,N_9592,N_8505);
xnor U15468 (N_15468,N_7093,N_9272);
and U15469 (N_15469,N_7280,N_8503);
nor U15470 (N_15470,N_11345,N_9896);
nand U15471 (N_15471,N_9365,N_7922);
xor U15472 (N_15472,N_6467,N_10977);
xor U15473 (N_15473,N_6059,N_9929);
and U15474 (N_15474,N_7407,N_11854);
nand U15475 (N_15475,N_9926,N_6685);
nand U15476 (N_15476,N_7155,N_8369);
and U15477 (N_15477,N_7368,N_7301);
nor U15478 (N_15478,N_10490,N_10314);
and U15479 (N_15479,N_8097,N_8295);
or U15480 (N_15480,N_10667,N_7939);
or U15481 (N_15481,N_7855,N_11825);
and U15482 (N_15482,N_9185,N_7798);
and U15483 (N_15483,N_7620,N_6606);
nor U15484 (N_15484,N_8768,N_9096);
nand U15485 (N_15485,N_11489,N_9261);
nor U15486 (N_15486,N_9547,N_7630);
xor U15487 (N_15487,N_10889,N_6047);
or U15488 (N_15488,N_11457,N_9739);
xnor U15489 (N_15489,N_9307,N_11997);
nand U15490 (N_15490,N_6643,N_8613);
and U15491 (N_15491,N_11539,N_10023);
xor U15492 (N_15492,N_7973,N_10393);
or U15493 (N_15493,N_7189,N_6868);
and U15494 (N_15494,N_11084,N_8838);
nor U15495 (N_15495,N_8655,N_8854);
nand U15496 (N_15496,N_8791,N_10872);
or U15497 (N_15497,N_8654,N_11363);
nand U15498 (N_15498,N_8005,N_10004);
xor U15499 (N_15499,N_8037,N_9879);
xor U15500 (N_15500,N_7864,N_8992);
or U15501 (N_15501,N_10055,N_8854);
nand U15502 (N_15502,N_6048,N_11742);
xnor U15503 (N_15503,N_9120,N_7170);
and U15504 (N_15504,N_10551,N_8806);
nor U15505 (N_15505,N_9802,N_11490);
nor U15506 (N_15506,N_6241,N_11604);
and U15507 (N_15507,N_6553,N_8099);
xnor U15508 (N_15508,N_9342,N_7583);
nand U15509 (N_15509,N_7756,N_11819);
nand U15510 (N_15510,N_9667,N_6392);
and U15511 (N_15511,N_10891,N_8924);
or U15512 (N_15512,N_7996,N_9697);
nor U15513 (N_15513,N_9411,N_8725);
xnor U15514 (N_15514,N_10941,N_9094);
nor U15515 (N_15515,N_9217,N_9583);
or U15516 (N_15516,N_8855,N_8548);
nand U15517 (N_15517,N_6848,N_7127);
and U15518 (N_15518,N_11686,N_6604);
nand U15519 (N_15519,N_6215,N_10607);
and U15520 (N_15520,N_8045,N_11202);
xor U15521 (N_15521,N_7251,N_8053);
nor U15522 (N_15522,N_9054,N_8296);
nand U15523 (N_15523,N_6715,N_9133);
and U15524 (N_15524,N_8180,N_9301);
nor U15525 (N_15525,N_6047,N_9606);
or U15526 (N_15526,N_10695,N_6336);
nand U15527 (N_15527,N_9355,N_8737);
nor U15528 (N_15528,N_7618,N_10214);
nor U15529 (N_15529,N_7964,N_9091);
nor U15530 (N_15530,N_10988,N_10658);
and U15531 (N_15531,N_7391,N_9389);
nand U15532 (N_15532,N_9225,N_9190);
nand U15533 (N_15533,N_7834,N_8868);
xor U15534 (N_15534,N_10434,N_8785);
nand U15535 (N_15535,N_11590,N_10507);
xnor U15536 (N_15536,N_8029,N_6539);
and U15537 (N_15537,N_10767,N_8588);
xor U15538 (N_15538,N_10316,N_9319);
xnor U15539 (N_15539,N_6557,N_9652);
and U15540 (N_15540,N_8928,N_9828);
and U15541 (N_15541,N_6592,N_10105);
nor U15542 (N_15542,N_7942,N_10046);
xnor U15543 (N_15543,N_10005,N_7523);
and U15544 (N_15544,N_10964,N_9092);
and U15545 (N_15545,N_6749,N_9510);
nand U15546 (N_15546,N_11597,N_6266);
or U15547 (N_15547,N_11176,N_9759);
or U15548 (N_15548,N_11567,N_9574);
xnor U15549 (N_15549,N_11598,N_11925);
xor U15550 (N_15550,N_8658,N_7418);
nor U15551 (N_15551,N_11572,N_8190);
nand U15552 (N_15552,N_7413,N_9951);
nor U15553 (N_15553,N_9507,N_10392);
nor U15554 (N_15554,N_9826,N_7347);
nand U15555 (N_15555,N_9943,N_10898);
nor U15556 (N_15556,N_11596,N_10775);
nand U15557 (N_15557,N_10899,N_11250);
xnor U15558 (N_15558,N_11728,N_11027);
and U15559 (N_15559,N_7647,N_6249);
nor U15560 (N_15560,N_9189,N_9743);
and U15561 (N_15561,N_11317,N_8167);
xor U15562 (N_15562,N_6669,N_10053);
or U15563 (N_15563,N_10205,N_8606);
xnor U15564 (N_15564,N_11401,N_8767);
nor U15565 (N_15565,N_9255,N_8396);
nor U15566 (N_15566,N_8280,N_11997);
xor U15567 (N_15567,N_8441,N_8586);
xnor U15568 (N_15568,N_7873,N_8216);
xor U15569 (N_15569,N_11150,N_8435);
nor U15570 (N_15570,N_10303,N_6004);
or U15571 (N_15571,N_11661,N_6893);
and U15572 (N_15572,N_8617,N_10059);
and U15573 (N_15573,N_10776,N_8074);
nand U15574 (N_15574,N_10203,N_11172);
and U15575 (N_15575,N_6657,N_8481);
and U15576 (N_15576,N_8160,N_8852);
and U15577 (N_15577,N_8062,N_8964);
xor U15578 (N_15578,N_8772,N_6994);
and U15579 (N_15579,N_10251,N_6209);
or U15580 (N_15580,N_7423,N_10583);
and U15581 (N_15581,N_10253,N_8561);
xnor U15582 (N_15582,N_10653,N_9151);
nor U15583 (N_15583,N_6209,N_11357);
or U15584 (N_15584,N_6389,N_11683);
nand U15585 (N_15585,N_7203,N_7279);
nor U15586 (N_15586,N_10630,N_10858);
and U15587 (N_15587,N_10072,N_6359);
or U15588 (N_15588,N_9409,N_8149);
xor U15589 (N_15589,N_9104,N_11019);
nand U15590 (N_15590,N_7652,N_8819);
xor U15591 (N_15591,N_7447,N_9989);
and U15592 (N_15592,N_9916,N_6044);
or U15593 (N_15593,N_8828,N_8349);
nand U15594 (N_15594,N_6993,N_6946);
or U15595 (N_15595,N_7860,N_8269);
nand U15596 (N_15596,N_6196,N_9758);
xor U15597 (N_15597,N_9907,N_6236);
nor U15598 (N_15598,N_11804,N_8492);
nor U15599 (N_15599,N_6282,N_10103);
and U15600 (N_15600,N_7076,N_6933);
and U15601 (N_15601,N_8327,N_7423);
xnor U15602 (N_15602,N_8155,N_9072);
xor U15603 (N_15603,N_7620,N_8529);
xnor U15604 (N_15604,N_7178,N_7424);
and U15605 (N_15605,N_6890,N_7913);
nand U15606 (N_15606,N_6731,N_9243);
nand U15607 (N_15607,N_10855,N_10584);
nand U15608 (N_15608,N_7211,N_11910);
or U15609 (N_15609,N_6321,N_9418);
nor U15610 (N_15610,N_8622,N_9804);
and U15611 (N_15611,N_10260,N_6233);
and U15612 (N_15612,N_7823,N_11316);
nand U15613 (N_15613,N_8515,N_9009);
xor U15614 (N_15614,N_6630,N_10197);
nand U15615 (N_15615,N_7933,N_11777);
nor U15616 (N_15616,N_8031,N_11676);
nand U15617 (N_15617,N_9879,N_9551);
nand U15618 (N_15618,N_9111,N_9921);
nor U15619 (N_15619,N_7722,N_9783);
and U15620 (N_15620,N_11971,N_7029);
and U15621 (N_15621,N_8494,N_8403);
or U15622 (N_15622,N_6084,N_9035);
nor U15623 (N_15623,N_9038,N_7360);
xor U15624 (N_15624,N_11030,N_6843);
xnor U15625 (N_15625,N_10770,N_9189);
nand U15626 (N_15626,N_7509,N_7483);
or U15627 (N_15627,N_7537,N_7452);
nor U15628 (N_15628,N_11131,N_10088);
xnor U15629 (N_15629,N_10156,N_8894);
nor U15630 (N_15630,N_11194,N_9858);
nand U15631 (N_15631,N_9792,N_9522);
nand U15632 (N_15632,N_7928,N_9410);
and U15633 (N_15633,N_11068,N_8268);
and U15634 (N_15634,N_8045,N_8866);
nand U15635 (N_15635,N_7191,N_8668);
xor U15636 (N_15636,N_7955,N_11491);
xnor U15637 (N_15637,N_9852,N_7016);
nor U15638 (N_15638,N_8696,N_9865);
xnor U15639 (N_15639,N_8003,N_7905);
and U15640 (N_15640,N_11152,N_9830);
or U15641 (N_15641,N_7240,N_9392);
nand U15642 (N_15642,N_9313,N_9303);
xor U15643 (N_15643,N_9696,N_11445);
nand U15644 (N_15644,N_9904,N_9189);
nand U15645 (N_15645,N_9885,N_8581);
xor U15646 (N_15646,N_8258,N_9239);
or U15647 (N_15647,N_11802,N_10099);
nand U15648 (N_15648,N_11739,N_6766);
or U15649 (N_15649,N_10145,N_6450);
xnor U15650 (N_15650,N_6542,N_7032);
xor U15651 (N_15651,N_10428,N_11887);
nor U15652 (N_15652,N_8106,N_6906);
and U15653 (N_15653,N_11226,N_10858);
or U15654 (N_15654,N_11179,N_11853);
xor U15655 (N_15655,N_8608,N_10106);
nand U15656 (N_15656,N_8751,N_7986);
and U15657 (N_15657,N_9875,N_10700);
or U15658 (N_15658,N_11983,N_6782);
xnor U15659 (N_15659,N_8376,N_11950);
xnor U15660 (N_15660,N_9316,N_7258);
and U15661 (N_15661,N_9255,N_8903);
or U15662 (N_15662,N_7727,N_6057);
nand U15663 (N_15663,N_7608,N_6104);
and U15664 (N_15664,N_6594,N_9274);
and U15665 (N_15665,N_6367,N_9701);
or U15666 (N_15666,N_6669,N_7422);
or U15667 (N_15667,N_7665,N_7105);
xnor U15668 (N_15668,N_11404,N_11014);
or U15669 (N_15669,N_6486,N_10276);
nand U15670 (N_15670,N_10161,N_6432);
and U15671 (N_15671,N_6312,N_6962);
nor U15672 (N_15672,N_9169,N_11343);
nand U15673 (N_15673,N_11406,N_10139);
nand U15674 (N_15674,N_6726,N_7210);
xnor U15675 (N_15675,N_9414,N_7963);
and U15676 (N_15676,N_11979,N_11048);
nor U15677 (N_15677,N_10889,N_8823);
and U15678 (N_15678,N_7478,N_11515);
nor U15679 (N_15679,N_10734,N_9973);
xnor U15680 (N_15680,N_9746,N_7997);
nand U15681 (N_15681,N_9689,N_7604);
xor U15682 (N_15682,N_6452,N_9602);
and U15683 (N_15683,N_7027,N_9427);
xor U15684 (N_15684,N_10310,N_8801);
or U15685 (N_15685,N_7125,N_8178);
nand U15686 (N_15686,N_6679,N_8317);
nand U15687 (N_15687,N_7545,N_6778);
nor U15688 (N_15688,N_11512,N_11966);
or U15689 (N_15689,N_6108,N_10416);
and U15690 (N_15690,N_6054,N_11697);
or U15691 (N_15691,N_7601,N_10277);
nor U15692 (N_15692,N_6739,N_6097);
or U15693 (N_15693,N_10375,N_11759);
xor U15694 (N_15694,N_11401,N_9341);
nor U15695 (N_15695,N_11608,N_7053);
nor U15696 (N_15696,N_8419,N_11864);
nand U15697 (N_15697,N_8366,N_9376);
xor U15698 (N_15698,N_11362,N_8539);
or U15699 (N_15699,N_7138,N_8382);
and U15700 (N_15700,N_6042,N_7429);
nand U15701 (N_15701,N_9047,N_11484);
and U15702 (N_15702,N_11108,N_10239);
and U15703 (N_15703,N_9609,N_7650);
or U15704 (N_15704,N_11058,N_11227);
and U15705 (N_15705,N_7916,N_6362);
xnor U15706 (N_15706,N_8530,N_9367);
and U15707 (N_15707,N_11499,N_8520);
xor U15708 (N_15708,N_6986,N_9333);
and U15709 (N_15709,N_9563,N_10390);
xor U15710 (N_15710,N_9145,N_10567);
or U15711 (N_15711,N_7332,N_7092);
xnor U15712 (N_15712,N_9792,N_10141);
nand U15713 (N_15713,N_7441,N_9884);
nor U15714 (N_15714,N_11468,N_8037);
or U15715 (N_15715,N_6175,N_8083);
nor U15716 (N_15716,N_10043,N_8815);
nand U15717 (N_15717,N_7202,N_11646);
xnor U15718 (N_15718,N_10003,N_10127);
or U15719 (N_15719,N_6522,N_6476);
xnor U15720 (N_15720,N_8805,N_7967);
and U15721 (N_15721,N_9035,N_8533);
or U15722 (N_15722,N_6338,N_6401);
xnor U15723 (N_15723,N_8834,N_6212);
and U15724 (N_15724,N_10792,N_6522);
or U15725 (N_15725,N_7868,N_10483);
xor U15726 (N_15726,N_8657,N_8489);
and U15727 (N_15727,N_6325,N_8943);
xor U15728 (N_15728,N_8035,N_11233);
xor U15729 (N_15729,N_7875,N_8804);
or U15730 (N_15730,N_8775,N_6620);
and U15731 (N_15731,N_10229,N_7760);
nand U15732 (N_15732,N_8046,N_7532);
nor U15733 (N_15733,N_6337,N_11323);
and U15734 (N_15734,N_10055,N_6485);
or U15735 (N_15735,N_7684,N_11013);
nor U15736 (N_15736,N_7024,N_7376);
or U15737 (N_15737,N_8653,N_9388);
nand U15738 (N_15738,N_10101,N_6977);
and U15739 (N_15739,N_11680,N_9241);
and U15740 (N_15740,N_8375,N_11329);
and U15741 (N_15741,N_9145,N_11859);
and U15742 (N_15742,N_11245,N_8940);
nor U15743 (N_15743,N_7360,N_9928);
or U15744 (N_15744,N_10589,N_9590);
or U15745 (N_15745,N_8999,N_9323);
and U15746 (N_15746,N_11647,N_9715);
nand U15747 (N_15747,N_7013,N_11059);
or U15748 (N_15748,N_7687,N_6197);
or U15749 (N_15749,N_11736,N_8562);
nor U15750 (N_15750,N_7085,N_8561);
nand U15751 (N_15751,N_6010,N_7211);
nor U15752 (N_15752,N_11897,N_9587);
nor U15753 (N_15753,N_7954,N_9684);
nand U15754 (N_15754,N_6130,N_6932);
or U15755 (N_15755,N_7718,N_7288);
or U15756 (N_15756,N_7363,N_8874);
or U15757 (N_15757,N_7436,N_8007);
nand U15758 (N_15758,N_8065,N_8603);
and U15759 (N_15759,N_9628,N_6048);
xor U15760 (N_15760,N_10498,N_10270);
nor U15761 (N_15761,N_6433,N_9785);
and U15762 (N_15762,N_7674,N_10231);
nor U15763 (N_15763,N_8907,N_10967);
xnor U15764 (N_15764,N_10481,N_6655);
xor U15765 (N_15765,N_6216,N_8297);
nand U15766 (N_15766,N_6218,N_7469);
nand U15767 (N_15767,N_10134,N_7736);
xnor U15768 (N_15768,N_9715,N_6008);
and U15769 (N_15769,N_7411,N_7426);
or U15770 (N_15770,N_6499,N_11811);
or U15771 (N_15771,N_10753,N_11430);
nand U15772 (N_15772,N_7941,N_9569);
xor U15773 (N_15773,N_7474,N_11487);
xnor U15774 (N_15774,N_10379,N_9997);
or U15775 (N_15775,N_8873,N_8552);
or U15776 (N_15776,N_6686,N_6978);
nand U15777 (N_15777,N_6302,N_9814);
or U15778 (N_15778,N_8020,N_6599);
nand U15779 (N_15779,N_6188,N_6205);
nor U15780 (N_15780,N_6877,N_9374);
nor U15781 (N_15781,N_10388,N_8066);
and U15782 (N_15782,N_10677,N_10588);
xnor U15783 (N_15783,N_7368,N_7399);
or U15784 (N_15784,N_11442,N_10480);
xnor U15785 (N_15785,N_11176,N_7152);
nor U15786 (N_15786,N_10423,N_11529);
nor U15787 (N_15787,N_8160,N_8440);
nand U15788 (N_15788,N_7363,N_7313);
or U15789 (N_15789,N_8153,N_8625);
and U15790 (N_15790,N_6921,N_11503);
nor U15791 (N_15791,N_11167,N_7266);
xnor U15792 (N_15792,N_10241,N_11811);
or U15793 (N_15793,N_6172,N_7233);
nor U15794 (N_15794,N_8191,N_9297);
xnor U15795 (N_15795,N_8564,N_11425);
and U15796 (N_15796,N_9374,N_8001);
nand U15797 (N_15797,N_10157,N_6090);
or U15798 (N_15798,N_7724,N_11985);
or U15799 (N_15799,N_11606,N_10934);
and U15800 (N_15800,N_11406,N_7719);
xnor U15801 (N_15801,N_8202,N_9663);
or U15802 (N_15802,N_8497,N_7187);
nand U15803 (N_15803,N_7626,N_10512);
nand U15804 (N_15804,N_7998,N_9037);
nor U15805 (N_15805,N_7311,N_9117);
nor U15806 (N_15806,N_8103,N_6840);
or U15807 (N_15807,N_11768,N_8249);
or U15808 (N_15808,N_7751,N_10139);
xor U15809 (N_15809,N_9037,N_7631);
and U15810 (N_15810,N_7321,N_10921);
and U15811 (N_15811,N_10188,N_10279);
xor U15812 (N_15812,N_9842,N_7339);
nor U15813 (N_15813,N_7846,N_7442);
and U15814 (N_15814,N_10372,N_10229);
nand U15815 (N_15815,N_11306,N_10256);
and U15816 (N_15816,N_9052,N_6548);
nand U15817 (N_15817,N_8860,N_7829);
nor U15818 (N_15818,N_10365,N_6939);
or U15819 (N_15819,N_8942,N_10943);
and U15820 (N_15820,N_7696,N_9139);
nor U15821 (N_15821,N_11142,N_6212);
nor U15822 (N_15822,N_7711,N_10549);
xor U15823 (N_15823,N_11696,N_9682);
nor U15824 (N_15824,N_7401,N_8937);
xnor U15825 (N_15825,N_10032,N_10625);
nor U15826 (N_15826,N_7491,N_11324);
and U15827 (N_15827,N_9003,N_9179);
xor U15828 (N_15828,N_7869,N_9066);
nor U15829 (N_15829,N_7906,N_9151);
nand U15830 (N_15830,N_6738,N_8376);
xnor U15831 (N_15831,N_6921,N_11812);
xor U15832 (N_15832,N_6639,N_8495);
and U15833 (N_15833,N_10783,N_7619);
or U15834 (N_15834,N_6526,N_8192);
nor U15835 (N_15835,N_11472,N_11155);
and U15836 (N_15836,N_10893,N_10924);
nor U15837 (N_15837,N_11598,N_8144);
nor U15838 (N_15838,N_11337,N_10013);
nor U15839 (N_15839,N_10845,N_10237);
nand U15840 (N_15840,N_9201,N_8011);
or U15841 (N_15841,N_10414,N_7179);
xor U15842 (N_15842,N_8698,N_11566);
xnor U15843 (N_15843,N_6756,N_6966);
or U15844 (N_15844,N_10784,N_8990);
or U15845 (N_15845,N_9262,N_8045);
and U15846 (N_15846,N_7800,N_10746);
or U15847 (N_15847,N_10827,N_8523);
or U15848 (N_15848,N_11097,N_10146);
or U15849 (N_15849,N_10464,N_8777);
nor U15850 (N_15850,N_11817,N_10299);
or U15851 (N_15851,N_9158,N_10610);
nor U15852 (N_15852,N_6692,N_7349);
nor U15853 (N_15853,N_9116,N_7532);
nor U15854 (N_15854,N_11432,N_6689);
and U15855 (N_15855,N_6575,N_8907);
or U15856 (N_15856,N_8367,N_9327);
nor U15857 (N_15857,N_8023,N_8741);
nor U15858 (N_15858,N_8049,N_10211);
or U15859 (N_15859,N_10508,N_9792);
or U15860 (N_15860,N_11926,N_6693);
or U15861 (N_15861,N_10771,N_9882);
xor U15862 (N_15862,N_8699,N_10683);
and U15863 (N_15863,N_6235,N_9915);
xnor U15864 (N_15864,N_11603,N_8046);
xor U15865 (N_15865,N_9863,N_11241);
nor U15866 (N_15866,N_10970,N_7546);
and U15867 (N_15867,N_9143,N_8652);
and U15868 (N_15868,N_8206,N_11303);
nand U15869 (N_15869,N_8313,N_8767);
nand U15870 (N_15870,N_8910,N_7974);
nor U15871 (N_15871,N_11759,N_9248);
or U15872 (N_15872,N_6085,N_7925);
and U15873 (N_15873,N_8456,N_6315);
and U15874 (N_15874,N_11234,N_6250);
xor U15875 (N_15875,N_6834,N_11755);
or U15876 (N_15876,N_6453,N_6100);
xnor U15877 (N_15877,N_6519,N_8971);
nor U15878 (N_15878,N_9628,N_10731);
and U15879 (N_15879,N_11864,N_7502);
or U15880 (N_15880,N_10115,N_10834);
or U15881 (N_15881,N_6257,N_10115);
nor U15882 (N_15882,N_8140,N_9941);
xnor U15883 (N_15883,N_9159,N_9498);
xor U15884 (N_15884,N_8469,N_7097);
xnor U15885 (N_15885,N_9063,N_8647);
nor U15886 (N_15886,N_9868,N_10920);
or U15887 (N_15887,N_9654,N_10864);
or U15888 (N_15888,N_6137,N_10341);
nor U15889 (N_15889,N_8394,N_9330);
or U15890 (N_15890,N_8019,N_11663);
nand U15891 (N_15891,N_10446,N_6602);
nand U15892 (N_15892,N_7999,N_11789);
xor U15893 (N_15893,N_10712,N_8971);
and U15894 (N_15894,N_8353,N_7700);
or U15895 (N_15895,N_6584,N_9884);
and U15896 (N_15896,N_6919,N_11625);
and U15897 (N_15897,N_7555,N_7641);
and U15898 (N_15898,N_11024,N_9264);
and U15899 (N_15899,N_11519,N_8480);
nand U15900 (N_15900,N_7365,N_6004);
nor U15901 (N_15901,N_7480,N_8901);
nor U15902 (N_15902,N_7324,N_7881);
and U15903 (N_15903,N_10069,N_7240);
and U15904 (N_15904,N_7277,N_7229);
nand U15905 (N_15905,N_8572,N_9579);
or U15906 (N_15906,N_9079,N_7531);
or U15907 (N_15907,N_11933,N_10914);
or U15908 (N_15908,N_10720,N_8597);
xnor U15909 (N_15909,N_8308,N_7699);
nand U15910 (N_15910,N_7723,N_11581);
and U15911 (N_15911,N_11808,N_6360);
xor U15912 (N_15912,N_11615,N_8506);
nor U15913 (N_15913,N_6049,N_8551);
or U15914 (N_15914,N_8886,N_6496);
and U15915 (N_15915,N_7368,N_9425);
nor U15916 (N_15916,N_7460,N_9683);
nand U15917 (N_15917,N_11586,N_11916);
xor U15918 (N_15918,N_11715,N_7197);
nor U15919 (N_15919,N_11165,N_9391);
nand U15920 (N_15920,N_8890,N_6490);
or U15921 (N_15921,N_8330,N_8809);
or U15922 (N_15922,N_8719,N_9210);
or U15923 (N_15923,N_8340,N_8227);
nand U15924 (N_15924,N_9005,N_6416);
and U15925 (N_15925,N_6793,N_9691);
or U15926 (N_15926,N_10780,N_10912);
or U15927 (N_15927,N_10265,N_11062);
xnor U15928 (N_15928,N_9110,N_6887);
or U15929 (N_15929,N_10749,N_7965);
nand U15930 (N_15930,N_9264,N_6166);
xor U15931 (N_15931,N_8264,N_11940);
or U15932 (N_15932,N_11633,N_7817);
and U15933 (N_15933,N_6474,N_7746);
and U15934 (N_15934,N_8927,N_10590);
and U15935 (N_15935,N_6790,N_10448);
nor U15936 (N_15936,N_10567,N_7422);
nor U15937 (N_15937,N_9971,N_11570);
and U15938 (N_15938,N_9787,N_7682);
nor U15939 (N_15939,N_8167,N_11581);
nor U15940 (N_15940,N_10794,N_10349);
nand U15941 (N_15941,N_9899,N_11014);
and U15942 (N_15942,N_10597,N_8146);
nand U15943 (N_15943,N_10132,N_9959);
and U15944 (N_15944,N_7789,N_11969);
or U15945 (N_15945,N_9524,N_6329);
xor U15946 (N_15946,N_9634,N_10008);
nand U15947 (N_15947,N_8828,N_10974);
nand U15948 (N_15948,N_9682,N_10322);
xor U15949 (N_15949,N_6019,N_7749);
xor U15950 (N_15950,N_9814,N_9091);
nor U15951 (N_15951,N_9542,N_9414);
nand U15952 (N_15952,N_9619,N_10270);
nor U15953 (N_15953,N_9074,N_6599);
and U15954 (N_15954,N_11213,N_8637);
or U15955 (N_15955,N_10580,N_11980);
and U15956 (N_15956,N_10574,N_9441);
nand U15957 (N_15957,N_7900,N_6623);
xnor U15958 (N_15958,N_11286,N_6906);
and U15959 (N_15959,N_10616,N_6002);
nand U15960 (N_15960,N_10018,N_7845);
and U15961 (N_15961,N_6007,N_10193);
nor U15962 (N_15962,N_11729,N_6819);
xor U15963 (N_15963,N_10700,N_9165);
nor U15964 (N_15964,N_11581,N_9303);
xor U15965 (N_15965,N_10674,N_7813);
or U15966 (N_15966,N_11215,N_6009);
nor U15967 (N_15967,N_10574,N_10873);
nand U15968 (N_15968,N_10726,N_10115);
nand U15969 (N_15969,N_9343,N_9482);
or U15970 (N_15970,N_8866,N_8554);
nand U15971 (N_15971,N_9743,N_10463);
and U15972 (N_15972,N_9669,N_10462);
and U15973 (N_15973,N_6828,N_6254);
xnor U15974 (N_15974,N_9451,N_7807);
nand U15975 (N_15975,N_10774,N_10008);
and U15976 (N_15976,N_10316,N_10933);
xor U15977 (N_15977,N_7143,N_11955);
xor U15978 (N_15978,N_6700,N_7076);
and U15979 (N_15979,N_8462,N_11879);
nor U15980 (N_15980,N_11402,N_7473);
xor U15981 (N_15981,N_9985,N_7420);
nand U15982 (N_15982,N_6986,N_7264);
xor U15983 (N_15983,N_7242,N_6485);
nand U15984 (N_15984,N_8565,N_9098);
and U15985 (N_15985,N_8126,N_6396);
or U15986 (N_15986,N_9308,N_10475);
and U15987 (N_15987,N_10470,N_6521);
xor U15988 (N_15988,N_8423,N_8458);
or U15989 (N_15989,N_6141,N_9173);
nor U15990 (N_15990,N_9284,N_10426);
or U15991 (N_15991,N_11847,N_7052);
nand U15992 (N_15992,N_6275,N_8249);
nand U15993 (N_15993,N_8136,N_8870);
and U15994 (N_15994,N_8877,N_10271);
or U15995 (N_15995,N_8087,N_8058);
nor U15996 (N_15996,N_11064,N_6700);
and U15997 (N_15997,N_10730,N_6669);
and U15998 (N_15998,N_11390,N_10174);
nand U15999 (N_15999,N_7038,N_6627);
or U16000 (N_16000,N_8027,N_8608);
or U16001 (N_16001,N_9450,N_8850);
xnor U16002 (N_16002,N_9682,N_7998);
or U16003 (N_16003,N_8174,N_11669);
nand U16004 (N_16004,N_11412,N_7385);
nand U16005 (N_16005,N_10705,N_11111);
and U16006 (N_16006,N_7125,N_8383);
and U16007 (N_16007,N_11146,N_8805);
and U16008 (N_16008,N_10436,N_8796);
xnor U16009 (N_16009,N_9338,N_6557);
xnor U16010 (N_16010,N_11575,N_6073);
and U16011 (N_16011,N_11724,N_6199);
nor U16012 (N_16012,N_7151,N_7762);
nor U16013 (N_16013,N_8307,N_10497);
or U16014 (N_16014,N_6731,N_9881);
xor U16015 (N_16015,N_7022,N_7553);
or U16016 (N_16016,N_6374,N_11886);
nand U16017 (N_16017,N_7878,N_11525);
or U16018 (N_16018,N_11894,N_9987);
nand U16019 (N_16019,N_6134,N_9993);
nand U16020 (N_16020,N_10683,N_7808);
nand U16021 (N_16021,N_8463,N_9892);
xnor U16022 (N_16022,N_6108,N_9141);
and U16023 (N_16023,N_6551,N_10123);
or U16024 (N_16024,N_11225,N_9591);
nor U16025 (N_16025,N_7004,N_6877);
and U16026 (N_16026,N_6881,N_9748);
and U16027 (N_16027,N_11481,N_8628);
xnor U16028 (N_16028,N_7491,N_6644);
and U16029 (N_16029,N_7441,N_10222);
nand U16030 (N_16030,N_6362,N_7977);
or U16031 (N_16031,N_9917,N_11075);
and U16032 (N_16032,N_6890,N_8412);
or U16033 (N_16033,N_10483,N_9533);
or U16034 (N_16034,N_10007,N_11712);
nor U16035 (N_16035,N_6067,N_10210);
xor U16036 (N_16036,N_7573,N_9004);
or U16037 (N_16037,N_10252,N_8433);
nand U16038 (N_16038,N_9369,N_7501);
and U16039 (N_16039,N_7251,N_11182);
or U16040 (N_16040,N_9229,N_6221);
and U16041 (N_16041,N_11412,N_10027);
xnor U16042 (N_16042,N_6660,N_11249);
xnor U16043 (N_16043,N_8916,N_10153);
and U16044 (N_16044,N_10536,N_11140);
or U16045 (N_16045,N_7052,N_6767);
or U16046 (N_16046,N_7422,N_11836);
nand U16047 (N_16047,N_8965,N_9579);
nor U16048 (N_16048,N_11866,N_6611);
xnor U16049 (N_16049,N_10678,N_10312);
xnor U16050 (N_16050,N_7627,N_10382);
nor U16051 (N_16051,N_6796,N_7673);
xor U16052 (N_16052,N_7492,N_9472);
and U16053 (N_16053,N_6407,N_10258);
nand U16054 (N_16054,N_9539,N_6792);
nand U16055 (N_16055,N_8504,N_6894);
or U16056 (N_16056,N_11028,N_10115);
or U16057 (N_16057,N_9980,N_8808);
xor U16058 (N_16058,N_7739,N_6601);
xor U16059 (N_16059,N_7421,N_10483);
nand U16060 (N_16060,N_7846,N_7554);
nand U16061 (N_16061,N_10318,N_8170);
and U16062 (N_16062,N_8603,N_6244);
nand U16063 (N_16063,N_9780,N_11784);
nor U16064 (N_16064,N_6527,N_9464);
nor U16065 (N_16065,N_11255,N_8676);
or U16066 (N_16066,N_6960,N_7762);
or U16067 (N_16067,N_9846,N_11111);
xor U16068 (N_16068,N_7153,N_7172);
and U16069 (N_16069,N_10022,N_9221);
and U16070 (N_16070,N_6259,N_9005);
xor U16071 (N_16071,N_10547,N_10415);
xor U16072 (N_16072,N_8114,N_10908);
nand U16073 (N_16073,N_8937,N_6617);
nor U16074 (N_16074,N_7603,N_6650);
or U16075 (N_16075,N_9047,N_8634);
nand U16076 (N_16076,N_8813,N_7935);
nor U16077 (N_16077,N_9512,N_10363);
nand U16078 (N_16078,N_9142,N_9294);
xnor U16079 (N_16079,N_9497,N_6790);
and U16080 (N_16080,N_7059,N_7166);
and U16081 (N_16081,N_7881,N_8334);
xnor U16082 (N_16082,N_11062,N_8272);
nor U16083 (N_16083,N_11542,N_7967);
xor U16084 (N_16084,N_11591,N_10005);
and U16085 (N_16085,N_11826,N_11641);
or U16086 (N_16086,N_6818,N_9879);
nand U16087 (N_16087,N_7666,N_6224);
nand U16088 (N_16088,N_7061,N_9879);
xnor U16089 (N_16089,N_8031,N_8762);
nor U16090 (N_16090,N_8441,N_10358);
nand U16091 (N_16091,N_9091,N_7422);
or U16092 (N_16092,N_9488,N_7042);
or U16093 (N_16093,N_9894,N_11171);
or U16094 (N_16094,N_6149,N_9832);
or U16095 (N_16095,N_11576,N_8044);
nor U16096 (N_16096,N_9611,N_9891);
or U16097 (N_16097,N_6348,N_10977);
xnor U16098 (N_16098,N_6774,N_6142);
or U16099 (N_16099,N_10976,N_9216);
nand U16100 (N_16100,N_8371,N_11504);
and U16101 (N_16101,N_6449,N_6175);
nand U16102 (N_16102,N_6071,N_11294);
nand U16103 (N_16103,N_9089,N_7065);
xor U16104 (N_16104,N_10542,N_7722);
or U16105 (N_16105,N_11492,N_9844);
xnor U16106 (N_16106,N_8146,N_10077);
and U16107 (N_16107,N_7904,N_6444);
nor U16108 (N_16108,N_10258,N_10123);
or U16109 (N_16109,N_8593,N_7249);
nand U16110 (N_16110,N_8189,N_11472);
nand U16111 (N_16111,N_9279,N_7150);
and U16112 (N_16112,N_9919,N_10157);
or U16113 (N_16113,N_7790,N_7162);
nor U16114 (N_16114,N_7021,N_8399);
xnor U16115 (N_16115,N_11886,N_6776);
nand U16116 (N_16116,N_7429,N_6789);
nand U16117 (N_16117,N_7721,N_6628);
and U16118 (N_16118,N_11394,N_8173);
or U16119 (N_16119,N_10178,N_11562);
nor U16120 (N_16120,N_7359,N_7718);
or U16121 (N_16121,N_9875,N_9626);
and U16122 (N_16122,N_10531,N_9525);
nand U16123 (N_16123,N_8299,N_11646);
xnor U16124 (N_16124,N_6188,N_11124);
nand U16125 (N_16125,N_7844,N_11122);
or U16126 (N_16126,N_10619,N_7003);
and U16127 (N_16127,N_7690,N_7469);
or U16128 (N_16128,N_6388,N_11478);
and U16129 (N_16129,N_8612,N_8555);
or U16130 (N_16130,N_7940,N_6987);
xor U16131 (N_16131,N_9489,N_9307);
or U16132 (N_16132,N_8167,N_8811);
xnor U16133 (N_16133,N_11421,N_9241);
nor U16134 (N_16134,N_9244,N_11664);
and U16135 (N_16135,N_7084,N_9581);
nand U16136 (N_16136,N_7488,N_9733);
and U16137 (N_16137,N_6651,N_8599);
and U16138 (N_16138,N_6458,N_6139);
and U16139 (N_16139,N_8959,N_11183);
nand U16140 (N_16140,N_6194,N_9794);
nor U16141 (N_16141,N_8208,N_10817);
xor U16142 (N_16142,N_7483,N_11417);
and U16143 (N_16143,N_9069,N_11908);
nor U16144 (N_16144,N_8194,N_8172);
nand U16145 (N_16145,N_6856,N_8611);
and U16146 (N_16146,N_10279,N_9661);
and U16147 (N_16147,N_6551,N_9382);
and U16148 (N_16148,N_9621,N_11878);
nand U16149 (N_16149,N_9195,N_11313);
nand U16150 (N_16150,N_7358,N_9044);
xor U16151 (N_16151,N_7217,N_6823);
nor U16152 (N_16152,N_6494,N_10501);
nand U16153 (N_16153,N_10002,N_8064);
and U16154 (N_16154,N_10669,N_11880);
or U16155 (N_16155,N_9335,N_8444);
and U16156 (N_16156,N_8491,N_10264);
nor U16157 (N_16157,N_6409,N_11505);
nor U16158 (N_16158,N_7508,N_6366);
nand U16159 (N_16159,N_9947,N_9866);
or U16160 (N_16160,N_11015,N_7021);
or U16161 (N_16161,N_6066,N_11589);
nand U16162 (N_16162,N_8272,N_11183);
nand U16163 (N_16163,N_6889,N_7145);
nand U16164 (N_16164,N_10406,N_9671);
and U16165 (N_16165,N_7741,N_9658);
or U16166 (N_16166,N_9138,N_7402);
nor U16167 (N_16167,N_9929,N_9869);
or U16168 (N_16168,N_11204,N_8391);
nand U16169 (N_16169,N_11657,N_10743);
nor U16170 (N_16170,N_9505,N_6585);
xnor U16171 (N_16171,N_8279,N_11302);
and U16172 (N_16172,N_6787,N_11326);
or U16173 (N_16173,N_10222,N_6797);
nor U16174 (N_16174,N_11668,N_9062);
nand U16175 (N_16175,N_10529,N_8440);
nor U16176 (N_16176,N_6440,N_9119);
nand U16177 (N_16177,N_7217,N_8973);
or U16178 (N_16178,N_7536,N_6241);
and U16179 (N_16179,N_9109,N_8134);
or U16180 (N_16180,N_11729,N_10101);
nand U16181 (N_16181,N_6738,N_6227);
or U16182 (N_16182,N_7816,N_6304);
nand U16183 (N_16183,N_7857,N_11276);
and U16184 (N_16184,N_11071,N_8966);
and U16185 (N_16185,N_6865,N_7240);
nor U16186 (N_16186,N_7735,N_6761);
or U16187 (N_16187,N_7988,N_6557);
and U16188 (N_16188,N_8170,N_7710);
nor U16189 (N_16189,N_6685,N_6034);
or U16190 (N_16190,N_10035,N_9106);
nand U16191 (N_16191,N_11230,N_10035);
xor U16192 (N_16192,N_11941,N_11845);
and U16193 (N_16193,N_9655,N_11661);
and U16194 (N_16194,N_9767,N_9921);
nor U16195 (N_16195,N_8351,N_11634);
and U16196 (N_16196,N_9623,N_9384);
xnor U16197 (N_16197,N_10202,N_10483);
xor U16198 (N_16198,N_10912,N_8820);
nand U16199 (N_16199,N_6223,N_9905);
nor U16200 (N_16200,N_7132,N_10222);
nor U16201 (N_16201,N_10467,N_9854);
nand U16202 (N_16202,N_8334,N_9937);
nor U16203 (N_16203,N_6729,N_7723);
xor U16204 (N_16204,N_8258,N_10131);
nand U16205 (N_16205,N_7557,N_10275);
nand U16206 (N_16206,N_8137,N_6675);
nand U16207 (N_16207,N_7036,N_9603);
or U16208 (N_16208,N_8503,N_6639);
or U16209 (N_16209,N_6769,N_8557);
nand U16210 (N_16210,N_11318,N_9435);
or U16211 (N_16211,N_8262,N_9373);
nand U16212 (N_16212,N_11605,N_11625);
nand U16213 (N_16213,N_6240,N_8850);
nor U16214 (N_16214,N_6835,N_6257);
nand U16215 (N_16215,N_6885,N_8782);
nor U16216 (N_16216,N_11003,N_10678);
and U16217 (N_16217,N_8222,N_10122);
nand U16218 (N_16218,N_8897,N_10703);
nand U16219 (N_16219,N_6656,N_7115);
nand U16220 (N_16220,N_6404,N_6780);
or U16221 (N_16221,N_8349,N_9197);
nand U16222 (N_16222,N_7923,N_7681);
nor U16223 (N_16223,N_6291,N_11734);
nor U16224 (N_16224,N_11960,N_9533);
and U16225 (N_16225,N_6507,N_8267);
xnor U16226 (N_16226,N_9661,N_10984);
xnor U16227 (N_16227,N_10510,N_6589);
nor U16228 (N_16228,N_9790,N_10853);
and U16229 (N_16229,N_9175,N_11305);
or U16230 (N_16230,N_9212,N_8777);
nor U16231 (N_16231,N_9185,N_11058);
nand U16232 (N_16232,N_7329,N_8830);
or U16233 (N_16233,N_9467,N_6372);
and U16234 (N_16234,N_9390,N_7630);
nor U16235 (N_16235,N_7541,N_7563);
nand U16236 (N_16236,N_7278,N_7169);
xnor U16237 (N_16237,N_10113,N_9979);
nor U16238 (N_16238,N_8219,N_9802);
and U16239 (N_16239,N_11904,N_6435);
xor U16240 (N_16240,N_7567,N_9734);
and U16241 (N_16241,N_9945,N_9529);
or U16242 (N_16242,N_10618,N_6355);
xnor U16243 (N_16243,N_9725,N_9625);
nand U16244 (N_16244,N_11531,N_10798);
nor U16245 (N_16245,N_10740,N_8095);
xor U16246 (N_16246,N_6896,N_9903);
nand U16247 (N_16247,N_10331,N_8956);
or U16248 (N_16248,N_10643,N_10493);
and U16249 (N_16249,N_6363,N_8394);
nor U16250 (N_16250,N_8761,N_8283);
nor U16251 (N_16251,N_7166,N_10636);
or U16252 (N_16252,N_6535,N_10376);
nand U16253 (N_16253,N_9169,N_9014);
and U16254 (N_16254,N_8495,N_9275);
nor U16255 (N_16255,N_11925,N_6543);
nand U16256 (N_16256,N_7389,N_11679);
nand U16257 (N_16257,N_8295,N_6331);
and U16258 (N_16258,N_6412,N_9386);
nand U16259 (N_16259,N_9391,N_11511);
xor U16260 (N_16260,N_11827,N_11817);
nand U16261 (N_16261,N_10766,N_8317);
nand U16262 (N_16262,N_9496,N_11056);
xor U16263 (N_16263,N_6151,N_8141);
and U16264 (N_16264,N_9101,N_9947);
xor U16265 (N_16265,N_10081,N_11846);
xnor U16266 (N_16266,N_9489,N_6122);
xnor U16267 (N_16267,N_11543,N_6124);
nand U16268 (N_16268,N_8942,N_7879);
xor U16269 (N_16269,N_10078,N_8949);
or U16270 (N_16270,N_8527,N_9377);
xnor U16271 (N_16271,N_7050,N_6503);
nor U16272 (N_16272,N_6166,N_6026);
nor U16273 (N_16273,N_11867,N_7558);
nor U16274 (N_16274,N_10483,N_9665);
or U16275 (N_16275,N_8742,N_8925);
nand U16276 (N_16276,N_11991,N_11947);
xor U16277 (N_16277,N_8839,N_11659);
nand U16278 (N_16278,N_7609,N_7667);
nor U16279 (N_16279,N_11246,N_7172);
and U16280 (N_16280,N_7313,N_8900);
and U16281 (N_16281,N_7735,N_11092);
or U16282 (N_16282,N_8080,N_8971);
and U16283 (N_16283,N_8688,N_10117);
xor U16284 (N_16284,N_11703,N_10386);
or U16285 (N_16285,N_11419,N_8295);
xor U16286 (N_16286,N_6736,N_6734);
or U16287 (N_16287,N_7636,N_7228);
and U16288 (N_16288,N_10716,N_10280);
xnor U16289 (N_16289,N_6068,N_6795);
and U16290 (N_16290,N_9616,N_8996);
nand U16291 (N_16291,N_7950,N_6494);
or U16292 (N_16292,N_10920,N_9528);
nand U16293 (N_16293,N_8479,N_9120);
and U16294 (N_16294,N_11287,N_6324);
xnor U16295 (N_16295,N_8846,N_10888);
xnor U16296 (N_16296,N_7570,N_10919);
nor U16297 (N_16297,N_8860,N_6048);
and U16298 (N_16298,N_8474,N_11291);
or U16299 (N_16299,N_6969,N_11135);
nand U16300 (N_16300,N_10470,N_11541);
or U16301 (N_16301,N_7251,N_8114);
nand U16302 (N_16302,N_10333,N_11064);
and U16303 (N_16303,N_10089,N_9875);
or U16304 (N_16304,N_11449,N_10822);
or U16305 (N_16305,N_11900,N_7147);
xnor U16306 (N_16306,N_9859,N_10926);
and U16307 (N_16307,N_7727,N_8431);
or U16308 (N_16308,N_9717,N_9471);
and U16309 (N_16309,N_9138,N_7020);
nand U16310 (N_16310,N_9473,N_10419);
nor U16311 (N_16311,N_9278,N_8794);
or U16312 (N_16312,N_9988,N_9678);
nand U16313 (N_16313,N_10901,N_6701);
xnor U16314 (N_16314,N_11432,N_9402);
xor U16315 (N_16315,N_8873,N_11742);
and U16316 (N_16316,N_8804,N_8559);
nand U16317 (N_16317,N_11319,N_11667);
and U16318 (N_16318,N_9869,N_9432);
and U16319 (N_16319,N_6993,N_8785);
nor U16320 (N_16320,N_6520,N_11967);
or U16321 (N_16321,N_10284,N_10416);
or U16322 (N_16322,N_8608,N_7899);
and U16323 (N_16323,N_9573,N_7189);
xor U16324 (N_16324,N_7918,N_11558);
nand U16325 (N_16325,N_8704,N_6587);
or U16326 (N_16326,N_6535,N_10614);
nor U16327 (N_16327,N_9317,N_7062);
xor U16328 (N_16328,N_6557,N_6336);
or U16329 (N_16329,N_8807,N_8036);
or U16330 (N_16330,N_6039,N_8913);
or U16331 (N_16331,N_7832,N_7202);
xnor U16332 (N_16332,N_6877,N_10287);
nor U16333 (N_16333,N_10616,N_6284);
nand U16334 (N_16334,N_7662,N_7313);
xor U16335 (N_16335,N_11810,N_10559);
nand U16336 (N_16336,N_11140,N_9502);
and U16337 (N_16337,N_8166,N_9142);
nor U16338 (N_16338,N_6895,N_8241);
xor U16339 (N_16339,N_11035,N_8328);
nor U16340 (N_16340,N_9378,N_7434);
or U16341 (N_16341,N_8280,N_8898);
and U16342 (N_16342,N_6280,N_11312);
and U16343 (N_16343,N_6480,N_7032);
nor U16344 (N_16344,N_10031,N_6349);
nand U16345 (N_16345,N_7238,N_10025);
nand U16346 (N_16346,N_7526,N_9555);
or U16347 (N_16347,N_9513,N_6143);
and U16348 (N_16348,N_8251,N_9441);
xor U16349 (N_16349,N_7304,N_6591);
nand U16350 (N_16350,N_11143,N_10165);
nand U16351 (N_16351,N_9134,N_8550);
and U16352 (N_16352,N_10938,N_6016);
or U16353 (N_16353,N_8524,N_9589);
xnor U16354 (N_16354,N_6513,N_6631);
nand U16355 (N_16355,N_7538,N_11300);
or U16356 (N_16356,N_10578,N_7138);
nand U16357 (N_16357,N_6373,N_10178);
or U16358 (N_16358,N_10036,N_8893);
nand U16359 (N_16359,N_11764,N_10632);
and U16360 (N_16360,N_7541,N_9804);
xor U16361 (N_16361,N_11491,N_8469);
and U16362 (N_16362,N_11650,N_8002);
or U16363 (N_16363,N_7742,N_8554);
xnor U16364 (N_16364,N_9605,N_9867);
or U16365 (N_16365,N_8975,N_6246);
nand U16366 (N_16366,N_7706,N_6294);
nand U16367 (N_16367,N_7128,N_6891);
or U16368 (N_16368,N_8385,N_11978);
xor U16369 (N_16369,N_8333,N_8074);
or U16370 (N_16370,N_6319,N_7552);
nand U16371 (N_16371,N_9248,N_11165);
nand U16372 (N_16372,N_9163,N_11152);
nor U16373 (N_16373,N_11213,N_11228);
nand U16374 (N_16374,N_8126,N_6437);
nor U16375 (N_16375,N_7197,N_6702);
and U16376 (N_16376,N_11265,N_11814);
nand U16377 (N_16377,N_9633,N_9048);
nor U16378 (N_16378,N_11734,N_10441);
or U16379 (N_16379,N_6268,N_10805);
or U16380 (N_16380,N_11025,N_6829);
nor U16381 (N_16381,N_10424,N_7040);
nor U16382 (N_16382,N_10924,N_7683);
nor U16383 (N_16383,N_11034,N_9687);
or U16384 (N_16384,N_8611,N_7901);
nor U16385 (N_16385,N_6878,N_10141);
or U16386 (N_16386,N_9726,N_9545);
xnor U16387 (N_16387,N_10358,N_9906);
or U16388 (N_16388,N_7715,N_8261);
nor U16389 (N_16389,N_10705,N_6145);
nand U16390 (N_16390,N_8236,N_10726);
xor U16391 (N_16391,N_8214,N_11082);
xor U16392 (N_16392,N_7386,N_11780);
nand U16393 (N_16393,N_9810,N_8764);
xnor U16394 (N_16394,N_10237,N_8550);
and U16395 (N_16395,N_8040,N_7589);
xnor U16396 (N_16396,N_10298,N_8838);
xor U16397 (N_16397,N_11815,N_7990);
and U16398 (N_16398,N_7582,N_7206);
nand U16399 (N_16399,N_7683,N_6342);
nor U16400 (N_16400,N_9264,N_7011);
xor U16401 (N_16401,N_9310,N_8774);
nand U16402 (N_16402,N_7089,N_6094);
nor U16403 (N_16403,N_7892,N_10296);
xor U16404 (N_16404,N_11083,N_10364);
and U16405 (N_16405,N_10046,N_9519);
nor U16406 (N_16406,N_11270,N_10246);
and U16407 (N_16407,N_11184,N_7599);
xor U16408 (N_16408,N_7522,N_9640);
xnor U16409 (N_16409,N_6214,N_8656);
nor U16410 (N_16410,N_9155,N_10878);
nand U16411 (N_16411,N_7059,N_10300);
or U16412 (N_16412,N_9880,N_6055);
xnor U16413 (N_16413,N_8976,N_11595);
xor U16414 (N_16414,N_11648,N_8140);
or U16415 (N_16415,N_7002,N_11564);
xnor U16416 (N_16416,N_6269,N_9499);
xnor U16417 (N_16417,N_11769,N_9557);
xor U16418 (N_16418,N_6265,N_10342);
and U16419 (N_16419,N_7177,N_8785);
xnor U16420 (N_16420,N_6621,N_8945);
nor U16421 (N_16421,N_9615,N_8760);
xnor U16422 (N_16422,N_7768,N_11856);
and U16423 (N_16423,N_7155,N_7492);
or U16424 (N_16424,N_11524,N_9724);
xnor U16425 (N_16425,N_10942,N_9185);
nor U16426 (N_16426,N_6167,N_6812);
xnor U16427 (N_16427,N_6981,N_9692);
xnor U16428 (N_16428,N_8534,N_11793);
xnor U16429 (N_16429,N_6940,N_11812);
or U16430 (N_16430,N_6665,N_7338);
nor U16431 (N_16431,N_6095,N_7704);
nor U16432 (N_16432,N_6970,N_10304);
xor U16433 (N_16433,N_6700,N_8602);
nand U16434 (N_16434,N_11084,N_7239);
or U16435 (N_16435,N_8165,N_11779);
and U16436 (N_16436,N_7175,N_9899);
or U16437 (N_16437,N_6116,N_6430);
and U16438 (N_16438,N_9389,N_9410);
nand U16439 (N_16439,N_11637,N_9979);
and U16440 (N_16440,N_7741,N_9298);
and U16441 (N_16441,N_8513,N_9439);
nand U16442 (N_16442,N_10706,N_8559);
nand U16443 (N_16443,N_6393,N_10345);
and U16444 (N_16444,N_6566,N_10906);
xnor U16445 (N_16445,N_10570,N_10488);
nor U16446 (N_16446,N_9856,N_7314);
xnor U16447 (N_16447,N_8072,N_10570);
xor U16448 (N_16448,N_7953,N_6039);
nand U16449 (N_16449,N_11921,N_7357);
xor U16450 (N_16450,N_10049,N_6067);
xnor U16451 (N_16451,N_8979,N_6043);
xnor U16452 (N_16452,N_7086,N_10159);
and U16453 (N_16453,N_10805,N_10590);
or U16454 (N_16454,N_6944,N_7656);
xor U16455 (N_16455,N_11696,N_7300);
and U16456 (N_16456,N_7952,N_6974);
xnor U16457 (N_16457,N_6587,N_7668);
nand U16458 (N_16458,N_8006,N_7247);
nand U16459 (N_16459,N_8178,N_9821);
xnor U16460 (N_16460,N_11129,N_9840);
xor U16461 (N_16461,N_6934,N_6834);
nand U16462 (N_16462,N_10749,N_6866);
xor U16463 (N_16463,N_8558,N_10399);
nor U16464 (N_16464,N_6432,N_6301);
nand U16465 (N_16465,N_9180,N_9860);
nand U16466 (N_16466,N_11523,N_7341);
xnor U16467 (N_16467,N_7214,N_8794);
or U16468 (N_16468,N_11185,N_9263);
and U16469 (N_16469,N_11374,N_11043);
nand U16470 (N_16470,N_9526,N_8470);
xnor U16471 (N_16471,N_9795,N_11768);
nor U16472 (N_16472,N_10523,N_10855);
nand U16473 (N_16473,N_10690,N_8162);
or U16474 (N_16474,N_7467,N_11924);
xor U16475 (N_16475,N_10799,N_6626);
nand U16476 (N_16476,N_9766,N_7712);
nor U16477 (N_16477,N_6329,N_10429);
xor U16478 (N_16478,N_9234,N_11877);
and U16479 (N_16479,N_6466,N_11645);
nand U16480 (N_16480,N_6488,N_11968);
and U16481 (N_16481,N_7718,N_11949);
xnor U16482 (N_16482,N_7935,N_6558);
and U16483 (N_16483,N_9085,N_9771);
xor U16484 (N_16484,N_8105,N_10567);
and U16485 (N_16485,N_7974,N_6914);
xor U16486 (N_16486,N_7577,N_11605);
or U16487 (N_16487,N_8839,N_10972);
nor U16488 (N_16488,N_6396,N_9318);
nand U16489 (N_16489,N_6697,N_7152);
or U16490 (N_16490,N_6419,N_6544);
and U16491 (N_16491,N_6167,N_11677);
nor U16492 (N_16492,N_7929,N_7915);
or U16493 (N_16493,N_10377,N_10109);
nand U16494 (N_16494,N_8958,N_10516);
or U16495 (N_16495,N_6263,N_6217);
and U16496 (N_16496,N_11831,N_8510);
or U16497 (N_16497,N_10869,N_7767);
and U16498 (N_16498,N_11325,N_10504);
nor U16499 (N_16499,N_8373,N_11523);
or U16500 (N_16500,N_7272,N_9766);
nand U16501 (N_16501,N_8902,N_7833);
or U16502 (N_16502,N_8605,N_10976);
xnor U16503 (N_16503,N_11240,N_8810);
nand U16504 (N_16504,N_8754,N_9932);
and U16505 (N_16505,N_6739,N_10466);
nand U16506 (N_16506,N_10554,N_11088);
nor U16507 (N_16507,N_9336,N_11564);
or U16508 (N_16508,N_11047,N_11501);
nand U16509 (N_16509,N_8522,N_9100);
xor U16510 (N_16510,N_9924,N_11344);
or U16511 (N_16511,N_6008,N_8252);
nor U16512 (N_16512,N_11716,N_6527);
or U16513 (N_16513,N_8075,N_8512);
nor U16514 (N_16514,N_10059,N_7354);
nand U16515 (N_16515,N_6949,N_6760);
xor U16516 (N_16516,N_9713,N_10169);
nor U16517 (N_16517,N_11241,N_11408);
or U16518 (N_16518,N_6800,N_6012);
nor U16519 (N_16519,N_10694,N_8880);
and U16520 (N_16520,N_11321,N_6556);
nor U16521 (N_16521,N_8829,N_6318);
nor U16522 (N_16522,N_9751,N_6862);
or U16523 (N_16523,N_6452,N_11494);
or U16524 (N_16524,N_9311,N_7983);
and U16525 (N_16525,N_6033,N_10399);
nand U16526 (N_16526,N_7264,N_11056);
nor U16527 (N_16527,N_11000,N_11249);
and U16528 (N_16528,N_11855,N_6380);
or U16529 (N_16529,N_11935,N_11133);
and U16530 (N_16530,N_10952,N_10028);
or U16531 (N_16531,N_8447,N_7530);
nor U16532 (N_16532,N_8143,N_10298);
xor U16533 (N_16533,N_10578,N_6273);
or U16534 (N_16534,N_7832,N_10670);
and U16535 (N_16535,N_7275,N_7147);
nor U16536 (N_16536,N_6332,N_11754);
nor U16537 (N_16537,N_9962,N_6460);
and U16538 (N_16538,N_6775,N_6138);
nor U16539 (N_16539,N_9231,N_6716);
xnor U16540 (N_16540,N_6324,N_11019);
nor U16541 (N_16541,N_9928,N_7843);
xnor U16542 (N_16542,N_8531,N_6818);
nor U16543 (N_16543,N_9950,N_8025);
xor U16544 (N_16544,N_8046,N_9339);
or U16545 (N_16545,N_11717,N_6178);
or U16546 (N_16546,N_6035,N_6447);
nor U16547 (N_16547,N_9325,N_10432);
or U16548 (N_16548,N_10549,N_6338);
and U16549 (N_16549,N_9952,N_11869);
and U16550 (N_16550,N_11384,N_7074);
or U16551 (N_16551,N_7675,N_10423);
and U16552 (N_16552,N_7077,N_8767);
nand U16553 (N_16553,N_6848,N_10504);
xor U16554 (N_16554,N_9765,N_10011);
xor U16555 (N_16555,N_9219,N_11943);
and U16556 (N_16556,N_10692,N_7910);
nor U16557 (N_16557,N_9166,N_6501);
nand U16558 (N_16558,N_6791,N_11080);
nor U16559 (N_16559,N_7466,N_7225);
and U16560 (N_16560,N_9394,N_11138);
nand U16561 (N_16561,N_9057,N_6989);
nand U16562 (N_16562,N_8773,N_7036);
nand U16563 (N_16563,N_9039,N_6569);
or U16564 (N_16564,N_7371,N_11954);
nor U16565 (N_16565,N_8241,N_6718);
nand U16566 (N_16566,N_9968,N_7911);
or U16567 (N_16567,N_7092,N_10934);
and U16568 (N_16568,N_7677,N_11534);
nor U16569 (N_16569,N_9138,N_11294);
xnor U16570 (N_16570,N_8480,N_10374);
nor U16571 (N_16571,N_8926,N_11984);
and U16572 (N_16572,N_7629,N_6758);
nor U16573 (N_16573,N_6412,N_7605);
nor U16574 (N_16574,N_9032,N_7200);
and U16575 (N_16575,N_7427,N_10488);
and U16576 (N_16576,N_9204,N_7638);
nand U16577 (N_16577,N_9784,N_6677);
nor U16578 (N_16578,N_9838,N_9362);
nand U16579 (N_16579,N_7339,N_7573);
and U16580 (N_16580,N_7317,N_9427);
and U16581 (N_16581,N_10948,N_11557);
and U16582 (N_16582,N_7801,N_6250);
and U16583 (N_16583,N_7058,N_8012);
and U16584 (N_16584,N_7625,N_8518);
nor U16585 (N_16585,N_11666,N_10114);
and U16586 (N_16586,N_9267,N_6593);
nor U16587 (N_16587,N_8126,N_10924);
and U16588 (N_16588,N_9617,N_8761);
nand U16589 (N_16589,N_8172,N_8458);
and U16590 (N_16590,N_10021,N_8657);
and U16591 (N_16591,N_9831,N_10718);
nand U16592 (N_16592,N_7186,N_10783);
nor U16593 (N_16593,N_10256,N_8425);
nor U16594 (N_16594,N_11987,N_11881);
nand U16595 (N_16595,N_8257,N_6210);
and U16596 (N_16596,N_11064,N_8797);
nand U16597 (N_16597,N_11115,N_8631);
or U16598 (N_16598,N_10573,N_10841);
xor U16599 (N_16599,N_9357,N_9103);
and U16600 (N_16600,N_9777,N_11970);
or U16601 (N_16601,N_7764,N_8707);
xnor U16602 (N_16602,N_6118,N_9959);
nand U16603 (N_16603,N_9838,N_9891);
or U16604 (N_16604,N_7903,N_10784);
and U16605 (N_16605,N_7122,N_8176);
or U16606 (N_16606,N_10586,N_11512);
xor U16607 (N_16607,N_10367,N_6974);
and U16608 (N_16608,N_7055,N_9744);
nor U16609 (N_16609,N_9742,N_8650);
xnor U16610 (N_16610,N_9721,N_8672);
nor U16611 (N_16611,N_6839,N_8022);
and U16612 (N_16612,N_8585,N_8536);
and U16613 (N_16613,N_9206,N_8602);
nand U16614 (N_16614,N_6478,N_7820);
nor U16615 (N_16615,N_11413,N_7077);
nand U16616 (N_16616,N_6724,N_9944);
nor U16617 (N_16617,N_9077,N_8041);
nand U16618 (N_16618,N_8663,N_8956);
nand U16619 (N_16619,N_11924,N_6662);
or U16620 (N_16620,N_11749,N_7432);
and U16621 (N_16621,N_11439,N_8329);
nor U16622 (N_16622,N_10744,N_10285);
xor U16623 (N_16623,N_7563,N_7458);
nor U16624 (N_16624,N_6283,N_9949);
nor U16625 (N_16625,N_8720,N_9370);
xor U16626 (N_16626,N_10960,N_9356);
and U16627 (N_16627,N_10158,N_6101);
or U16628 (N_16628,N_6056,N_6053);
nor U16629 (N_16629,N_6227,N_8016);
or U16630 (N_16630,N_9631,N_9123);
nor U16631 (N_16631,N_7056,N_10310);
nor U16632 (N_16632,N_10450,N_11232);
nand U16633 (N_16633,N_6215,N_11691);
or U16634 (N_16634,N_9810,N_7487);
nand U16635 (N_16635,N_8327,N_8232);
or U16636 (N_16636,N_11134,N_10618);
nand U16637 (N_16637,N_6577,N_10265);
and U16638 (N_16638,N_10938,N_8250);
and U16639 (N_16639,N_6860,N_8754);
xnor U16640 (N_16640,N_8799,N_10443);
or U16641 (N_16641,N_6789,N_9469);
or U16642 (N_16642,N_8618,N_9768);
xor U16643 (N_16643,N_8620,N_10051);
nor U16644 (N_16644,N_11473,N_6927);
nand U16645 (N_16645,N_9470,N_6886);
and U16646 (N_16646,N_11779,N_8912);
xnor U16647 (N_16647,N_9952,N_11926);
nand U16648 (N_16648,N_8624,N_6895);
xor U16649 (N_16649,N_10291,N_8159);
nand U16650 (N_16650,N_8243,N_7372);
or U16651 (N_16651,N_8655,N_11848);
or U16652 (N_16652,N_6010,N_10759);
or U16653 (N_16653,N_9365,N_8637);
nand U16654 (N_16654,N_8709,N_10289);
nor U16655 (N_16655,N_7913,N_11937);
and U16656 (N_16656,N_8756,N_9533);
xor U16657 (N_16657,N_7161,N_8449);
and U16658 (N_16658,N_11965,N_7242);
or U16659 (N_16659,N_11218,N_6854);
nor U16660 (N_16660,N_9382,N_10484);
or U16661 (N_16661,N_11813,N_10075);
and U16662 (N_16662,N_10297,N_8451);
xnor U16663 (N_16663,N_6311,N_9311);
nand U16664 (N_16664,N_10195,N_11073);
nand U16665 (N_16665,N_7010,N_9850);
and U16666 (N_16666,N_9075,N_7176);
nor U16667 (N_16667,N_8036,N_6280);
nor U16668 (N_16668,N_9068,N_6824);
or U16669 (N_16669,N_11343,N_11928);
or U16670 (N_16670,N_6820,N_7080);
xnor U16671 (N_16671,N_6723,N_8105);
nor U16672 (N_16672,N_9640,N_6246);
or U16673 (N_16673,N_8534,N_11408);
or U16674 (N_16674,N_11623,N_10086);
xor U16675 (N_16675,N_11392,N_7545);
xnor U16676 (N_16676,N_7041,N_10744);
or U16677 (N_16677,N_9426,N_7255);
nor U16678 (N_16678,N_10520,N_7678);
xor U16679 (N_16679,N_8276,N_11693);
nand U16680 (N_16680,N_7011,N_7399);
and U16681 (N_16681,N_8154,N_11599);
and U16682 (N_16682,N_9910,N_6091);
and U16683 (N_16683,N_6983,N_11780);
and U16684 (N_16684,N_6730,N_6766);
nand U16685 (N_16685,N_7951,N_10552);
nor U16686 (N_16686,N_11528,N_10074);
xor U16687 (N_16687,N_6685,N_9116);
xnor U16688 (N_16688,N_8350,N_11584);
xnor U16689 (N_16689,N_9616,N_9380);
or U16690 (N_16690,N_8101,N_8759);
nor U16691 (N_16691,N_11773,N_9371);
or U16692 (N_16692,N_9670,N_11489);
nor U16693 (N_16693,N_11587,N_9423);
xnor U16694 (N_16694,N_11427,N_8324);
or U16695 (N_16695,N_10863,N_6922);
xor U16696 (N_16696,N_10109,N_10777);
nor U16697 (N_16697,N_10076,N_8029);
and U16698 (N_16698,N_8984,N_7825);
nor U16699 (N_16699,N_7171,N_7691);
and U16700 (N_16700,N_9290,N_7452);
nor U16701 (N_16701,N_7775,N_9164);
nand U16702 (N_16702,N_10937,N_8378);
xor U16703 (N_16703,N_7758,N_10090);
or U16704 (N_16704,N_8263,N_8612);
nor U16705 (N_16705,N_9863,N_6916);
and U16706 (N_16706,N_8363,N_8337);
xnor U16707 (N_16707,N_11680,N_6760);
or U16708 (N_16708,N_7715,N_9743);
nand U16709 (N_16709,N_7171,N_8480);
xnor U16710 (N_16710,N_6579,N_8159);
or U16711 (N_16711,N_6788,N_8773);
and U16712 (N_16712,N_7318,N_7076);
nor U16713 (N_16713,N_10044,N_10404);
and U16714 (N_16714,N_8944,N_8842);
and U16715 (N_16715,N_9400,N_11389);
nand U16716 (N_16716,N_6756,N_8299);
xor U16717 (N_16717,N_10056,N_6094);
xnor U16718 (N_16718,N_6728,N_6950);
xnor U16719 (N_16719,N_7432,N_9964);
xor U16720 (N_16720,N_7928,N_6625);
and U16721 (N_16721,N_9340,N_11749);
nand U16722 (N_16722,N_9668,N_6678);
xnor U16723 (N_16723,N_10396,N_7853);
or U16724 (N_16724,N_11563,N_9141);
and U16725 (N_16725,N_10029,N_11883);
or U16726 (N_16726,N_9786,N_6123);
nand U16727 (N_16727,N_7685,N_7487);
or U16728 (N_16728,N_10714,N_8678);
nand U16729 (N_16729,N_6329,N_9270);
nand U16730 (N_16730,N_8681,N_11961);
or U16731 (N_16731,N_10387,N_10513);
nand U16732 (N_16732,N_8574,N_11177);
xnor U16733 (N_16733,N_7134,N_6431);
xor U16734 (N_16734,N_6819,N_7971);
nor U16735 (N_16735,N_8464,N_6176);
nor U16736 (N_16736,N_7750,N_10566);
or U16737 (N_16737,N_6141,N_8405);
xnor U16738 (N_16738,N_8474,N_6356);
xor U16739 (N_16739,N_8566,N_11189);
nand U16740 (N_16740,N_10327,N_6884);
nor U16741 (N_16741,N_7925,N_6466);
nand U16742 (N_16742,N_10528,N_9567);
or U16743 (N_16743,N_11448,N_9317);
and U16744 (N_16744,N_7773,N_6137);
xnor U16745 (N_16745,N_11097,N_9739);
and U16746 (N_16746,N_8875,N_6551);
nor U16747 (N_16747,N_11820,N_7981);
xnor U16748 (N_16748,N_11622,N_7561);
xnor U16749 (N_16749,N_11018,N_8802);
and U16750 (N_16750,N_11902,N_10964);
xnor U16751 (N_16751,N_8719,N_9084);
xnor U16752 (N_16752,N_7673,N_7394);
nor U16753 (N_16753,N_6387,N_7672);
and U16754 (N_16754,N_10380,N_7998);
nand U16755 (N_16755,N_6810,N_7957);
nor U16756 (N_16756,N_7980,N_7365);
nor U16757 (N_16757,N_11813,N_8264);
and U16758 (N_16758,N_7783,N_7101);
nand U16759 (N_16759,N_8521,N_11875);
xnor U16760 (N_16760,N_7591,N_8170);
and U16761 (N_16761,N_10286,N_6119);
nand U16762 (N_16762,N_11811,N_8940);
or U16763 (N_16763,N_6433,N_11113);
and U16764 (N_16764,N_10615,N_10850);
xor U16765 (N_16765,N_7744,N_9067);
or U16766 (N_16766,N_11343,N_11581);
and U16767 (N_16767,N_9955,N_10328);
and U16768 (N_16768,N_9183,N_11693);
or U16769 (N_16769,N_8070,N_6278);
xor U16770 (N_16770,N_7293,N_10156);
xor U16771 (N_16771,N_10003,N_8059);
nor U16772 (N_16772,N_9092,N_10440);
and U16773 (N_16773,N_8699,N_10085);
nor U16774 (N_16774,N_6566,N_7975);
and U16775 (N_16775,N_9693,N_9415);
nand U16776 (N_16776,N_9304,N_9974);
and U16777 (N_16777,N_7479,N_10675);
nor U16778 (N_16778,N_11269,N_11895);
xor U16779 (N_16779,N_6367,N_9480);
and U16780 (N_16780,N_10706,N_7308);
and U16781 (N_16781,N_9518,N_11117);
and U16782 (N_16782,N_6322,N_10658);
nor U16783 (N_16783,N_7452,N_9119);
and U16784 (N_16784,N_9237,N_9685);
xor U16785 (N_16785,N_6052,N_6022);
nand U16786 (N_16786,N_10963,N_11450);
and U16787 (N_16787,N_9853,N_6676);
nor U16788 (N_16788,N_10716,N_11406);
or U16789 (N_16789,N_8132,N_10861);
xor U16790 (N_16790,N_6176,N_11327);
or U16791 (N_16791,N_9109,N_6075);
nor U16792 (N_16792,N_7548,N_8528);
nor U16793 (N_16793,N_9973,N_9933);
nor U16794 (N_16794,N_8626,N_10094);
xnor U16795 (N_16795,N_11810,N_11889);
xnor U16796 (N_16796,N_7434,N_7056);
nand U16797 (N_16797,N_11464,N_9695);
xor U16798 (N_16798,N_9277,N_6586);
nand U16799 (N_16799,N_9798,N_10164);
nand U16800 (N_16800,N_9614,N_9404);
or U16801 (N_16801,N_11912,N_8873);
xnor U16802 (N_16802,N_10873,N_7147);
xor U16803 (N_16803,N_9841,N_10371);
xor U16804 (N_16804,N_11614,N_6129);
nand U16805 (N_16805,N_10546,N_8902);
xor U16806 (N_16806,N_7791,N_10511);
xor U16807 (N_16807,N_7269,N_9693);
nor U16808 (N_16808,N_11481,N_11639);
nand U16809 (N_16809,N_7834,N_8349);
xor U16810 (N_16810,N_6764,N_6648);
and U16811 (N_16811,N_10842,N_9985);
or U16812 (N_16812,N_6835,N_11429);
nand U16813 (N_16813,N_8762,N_8045);
and U16814 (N_16814,N_9451,N_7569);
or U16815 (N_16815,N_7090,N_10351);
nor U16816 (N_16816,N_8376,N_8668);
xor U16817 (N_16817,N_7667,N_7631);
xor U16818 (N_16818,N_9038,N_11582);
nand U16819 (N_16819,N_7978,N_8124);
nor U16820 (N_16820,N_6333,N_7775);
or U16821 (N_16821,N_8289,N_7459);
and U16822 (N_16822,N_11802,N_10650);
or U16823 (N_16823,N_11525,N_7342);
nor U16824 (N_16824,N_10590,N_10222);
nand U16825 (N_16825,N_8191,N_11507);
or U16826 (N_16826,N_8214,N_8507);
and U16827 (N_16827,N_6505,N_6769);
nor U16828 (N_16828,N_6123,N_11006);
nand U16829 (N_16829,N_6829,N_10122);
xnor U16830 (N_16830,N_11590,N_10865);
nand U16831 (N_16831,N_8218,N_9686);
nand U16832 (N_16832,N_6961,N_6087);
or U16833 (N_16833,N_8619,N_9072);
or U16834 (N_16834,N_8854,N_8665);
or U16835 (N_16835,N_6375,N_6086);
nor U16836 (N_16836,N_7401,N_8541);
and U16837 (N_16837,N_6842,N_10955);
or U16838 (N_16838,N_9582,N_7732);
nor U16839 (N_16839,N_10494,N_9497);
nand U16840 (N_16840,N_6221,N_8029);
and U16841 (N_16841,N_8972,N_9275);
xor U16842 (N_16842,N_10991,N_11000);
xor U16843 (N_16843,N_8316,N_10585);
and U16844 (N_16844,N_10714,N_8701);
or U16845 (N_16845,N_7417,N_10896);
nor U16846 (N_16846,N_7034,N_6243);
nor U16847 (N_16847,N_7554,N_10488);
and U16848 (N_16848,N_11203,N_11343);
and U16849 (N_16849,N_9882,N_7262);
or U16850 (N_16850,N_9729,N_10478);
or U16851 (N_16851,N_9661,N_6454);
nor U16852 (N_16852,N_8637,N_7379);
and U16853 (N_16853,N_6714,N_10239);
and U16854 (N_16854,N_6258,N_8694);
nand U16855 (N_16855,N_8943,N_6941);
and U16856 (N_16856,N_10955,N_8415);
xnor U16857 (N_16857,N_10718,N_8982);
or U16858 (N_16858,N_7667,N_10834);
and U16859 (N_16859,N_10881,N_9759);
xnor U16860 (N_16860,N_6356,N_11767);
and U16861 (N_16861,N_8819,N_10362);
nor U16862 (N_16862,N_8323,N_8725);
nor U16863 (N_16863,N_6995,N_10936);
or U16864 (N_16864,N_8677,N_9799);
xnor U16865 (N_16865,N_6352,N_8697);
xnor U16866 (N_16866,N_10114,N_7404);
nor U16867 (N_16867,N_6088,N_9999);
nor U16868 (N_16868,N_7286,N_9598);
or U16869 (N_16869,N_10192,N_10433);
and U16870 (N_16870,N_9150,N_6559);
and U16871 (N_16871,N_9310,N_9484);
xor U16872 (N_16872,N_11832,N_7319);
nor U16873 (N_16873,N_10340,N_9562);
or U16874 (N_16874,N_11755,N_10890);
or U16875 (N_16875,N_8599,N_11050);
xnor U16876 (N_16876,N_7148,N_8136);
or U16877 (N_16877,N_7996,N_8488);
or U16878 (N_16878,N_8023,N_7751);
xnor U16879 (N_16879,N_7830,N_11889);
and U16880 (N_16880,N_6521,N_7725);
nand U16881 (N_16881,N_11742,N_7890);
or U16882 (N_16882,N_6943,N_10477);
or U16883 (N_16883,N_6947,N_11225);
or U16884 (N_16884,N_11321,N_10118);
nor U16885 (N_16885,N_8777,N_8642);
nand U16886 (N_16886,N_6379,N_10288);
nor U16887 (N_16887,N_11914,N_7619);
or U16888 (N_16888,N_10886,N_9919);
or U16889 (N_16889,N_11857,N_7058);
xor U16890 (N_16890,N_10587,N_9474);
and U16891 (N_16891,N_9990,N_11211);
nand U16892 (N_16892,N_10167,N_7770);
and U16893 (N_16893,N_7510,N_6037);
and U16894 (N_16894,N_11868,N_7028);
nor U16895 (N_16895,N_9830,N_11512);
and U16896 (N_16896,N_10909,N_10784);
xor U16897 (N_16897,N_9386,N_9428);
nor U16898 (N_16898,N_8826,N_9321);
and U16899 (N_16899,N_6104,N_9446);
nor U16900 (N_16900,N_10850,N_7948);
and U16901 (N_16901,N_7760,N_11428);
nand U16902 (N_16902,N_7196,N_10599);
nand U16903 (N_16903,N_11059,N_7767);
xnor U16904 (N_16904,N_8848,N_10980);
nand U16905 (N_16905,N_11525,N_11268);
or U16906 (N_16906,N_9077,N_10898);
and U16907 (N_16907,N_9656,N_6734);
nand U16908 (N_16908,N_11275,N_6159);
or U16909 (N_16909,N_9817,N_9691);
and U16910 (N_16910,N_11387,N_8997);
or U16911 (N_16911,N_9448,N_9322);
nor U16912 (N_16912,N_10731,N_7458);
nand U16913 (N_16913,N_11766,N_6144);
xor U16914 (N_16914,N_7369,N_7951);
xnor U16915 (N_16915,N_11758,N_8679);
nor U16916 (N_16916,N_10392,N_11557);
nand U16917 (N_16917,N_8549,N_11106);
xnor U16918 (N_16918,N_9897,N_8312);
nand U16919 (N_16919,N_10285,N_9692);
or U16920 (N_16920,N_8003,N_11108);
nor U16921 (N_16921,N_8644,N_11732);
nand U16922 (N_16922,N_8412,N_10585);
nand U16923 (N_16923,N_7174,N_7744);
xor U16924 (N_16924,N_8028,N_8562);
nand U16925 (N_16925,N_8228,N_11293);
nor U16926 (N_16926,N_7561,N_10195);
nor U16927 (N_16927,N_7046,N_10748);
or U16928 (N_16928,N_10027,N_8970);
nand U16929 (N_16929,N_7244,N_6098);
or U16930 (N_16930,N_7493,N_6483);
nor U16931 (N_16931,N_6465,N_10359);
and U16932 (N_16932,N_6657,N_9220);
nor U16933 (N_16933,N_9132,N_8775);
nand U16934 (N_16934,N_11401,N_11115);
xor U16935 (N_16935,N_11338,N_8599);
xnor U16936 (N_16936,N_11779,N_6135);
nand U16937 (N_16937,N_10120,N_9792);
or U16938 (N_16938,N_7614,N_9319);
or U16939 (N_16939,N_10177,N_8181);
and U16940 (N_16940,N_6761,N_9330);
and U16941 (N_16941,N_7941,N_10690);
and U16942 (N_16942,N_8138,N_7385);
nor U16943 (N_16943,N_10393,N_8483);
or U16944 (N_16944,N_11100,N_9902);
nor U16945 (N_16945,N_9948,N_6036);
and U16946 (N_16946,N_10506,N_7154);
nor U16947 (N_16947,N_6272,N_11061);
nor U16948 (N_16948,N_8255,N_7135);
nor U16949 (N_16949,N_7495,N_7690);
and U16950 (N_16950,N_7227,N_7321);
nand U16951 (N_16951,N_9661,N_10032);
or U16952 (N_16952,N_7975,N_11158);
or U16953 (N_16953,N_8620,N_11900);
nor U16954 (N_16954,N_6062,N_9480);
nor U16955 (N_16955,N_8178,N_9717);
and U16956 (N_16956,N_11716,N_6188);
and U16957 (N_16957,N_8803,N_10425);
xnor U16958 (N_16958,N_9349,N_10476);
nor U16959 (N_16959,N_9946,N_6670);
or U16960 (N_16960,N_8887,N_8220);
and U16961 (N_16961,N_6479,N_9047);
and U16962 (N_16962,N_6473,N_10526);
nor U16963 (N_16963,N_11266,N_8239);
or U16964 (N_16964,N_7175,N_11445);
nand U16965 (N_16965,N_8071,N_8939);
nand U16966 (N_16966,N_10599,N_8619);
or U16967 (N_16967,N_6441,N_7974);
nand U16968 (N_16968,N_7767,N_7572);
xnor U16969 (N_16969,N_10393,N_8863);
and U16970 (N_16970,N_8769,N_10462);
nand U16971 (N_16971,N_10878,N_7905);
nand U16972 (N_16972,N_7391,N_11724);
and U16973 (N_16973,N_10136,N_6299);
xnor U16974 (N_16974,N_10771,N_9104);
or U16975 (N_16975,N_8875,N_10841);
and U16976 (N_16976,N_6437,N_6982);
and U16977 (N_16977,N_9492,N_7067);
nor U16978 (N_16978,N_6672,N_9589);
and U16979 (N_16979,N_10327,N_11098);
and U16980 (N_16980,N_10794,N_10433);
nand U16981 (N_16981,N_11998,N_10017);
nor U16982 (N_16982,N_6464,N_11286);
nor U16983 (N_16983,N_8444,N_9253);
xor U16984 (N_16984,N_11370,N_7375);
or U16985 (N_16985,N_11226,N_10386);
nor U16986 (N_16986,N_10709,N_7799);
and U16987 (N_16987,N_8458,N_7503);
and U16988 (N_16988,N_9891,N_10705);
nand U16989 (N_16989,N_7938,N_6561);
nor U16990 (N_16990,N_9073,N_10850);
and U16991 (N_16991,N_6321,N_7222);
nand U16992 (N_16992,N_8313,N_10769);
or U16993 (N_16993,N_7536,N_6752);
or U16994 (N_16994,N_11679,N_10543);
xor U16995 (N_16995,N_11384,N_6721);
xnor U16996 (N_16996,N_11400,N_10325);
nor U16997 (N_16997,N_10308,N_8546);
or U16998 (N_16998,N_10194,N_7494);
nor U16999 (N_16999,N_11135,N_7228);
xnor U17000 (N_17000,N_11545,N_7536);
and U17001 (N_17001,N_10418,N_7561);
nand U17002 (N_17002,N_11914,N_9768);
xor U17003 (N_17003,N_10947,N_9394);
and U17004 (N_17004,N_6492,N_11411);
nand U17005 (N_17005,N_9339,N_11529);
and U17006 (N_17006,N_9969,N_11031);
and U17007 (N_17007,N_6852,N_10647);
nand U17008 (N_17008,N_7297,N_9456);
nand U17009 (N_17009,N_9441,N_11108);
and U17010 (N_17010,N_11759,N_11095);
or U17011 (N_17011,N_10548,N_11193);
nand U17012 (N_17012,N_8056,N_11824);
and U17013 (N_17013,N_10402,N_6396);
and U17014 (N_17014,N_11898,N_9023);
or U17015 (N_17015,N_6210,N_11089);
xnor U17016 (N_17016,N_10844,N_11585);
xor U17017 (N_17017,N_8405,N_11088);
nor U17018 (N_17018,N_10405,N_7794);
or U17019 (N_17019,N_11109,N_11351);
xnor U17020 (N_17020,N_8963,N_9112);
nand U17021 (N_17021,N_11433,N_6970);
nand U17022 (N_17022,N_11297,N_6355);
xnor U17023 (N_17023,N_10678,N_7513);
nand U17024 (N_17024,N_6888,N_9549);
nor U17025 (N_17025,N_9567,N_10031);
xnor U17026 (N_17026,N_9073,N_11704);
xor U17027 (N_17027,N_6799,N_6009);
and U17028 (N_17028,N_7385,N_9681);
and U17029 (N_17029,N_6058,N_11264);
or U17030 (N_17030,N_8545,N_7989);
or U17031 (N_17031,N_7300,N_8437);
nor U17032 (N_17032,N_6413,N_11916);
nor U17033 (N_17033,N_10487,N_8647);
and U17034 (N_17034,N_7402,N_9109);
or U17035 (N_17035,N_6712,N_6662);
nand U17036 (N_17036,N_8920,N_7871);
nor U17037 (N_17037,N_7598,N_7232);
nor U17038 (N_17038,N_7712,N_10859);
xor U17039 (N_17039,N_7642,N_11161);
xnor U17040 (N_17040,N_11400,N_10772);
or U17041 (N_17041,N_9371,N_10540);
xor U17042 (N_17042,N_11708,N_6974);
or U17043 (N_17043,N_11694,N_7967);
or U17044 (N_17044,N_7191,N_7104);
xnor U17045 (N_17045,N_9512,N_11816);
and U17046 (N_17046,N_11654,N_6757);
nand U17047 (N_17047,N_6324,N_7324);
and U17048 (N_17048,N_8473,N_11172);
and U17049 (N_17049,N_10004,N_8349);
xor U17050 (N_17050,N_9679,N_6460);
xor U17051 (N_17051,N_6252,N_11883);
or U17052 (N_17052,N_10379,N_8963);
nand U17053 (N_17053,N_11469,N_10307);
nor U17054 (N_17054,N_6435,N_6120);
nand U17055 (N_17055,N_11495,N_10212);
or U17056 (N_17056,N_10645,N_9923);
and U17057 (N_17057,N_11466,N_10488);
nor U17058 (N_17058,N_6488,N_6721);
and U17059 (N_17059,N_11625,N_8715);
xnor U17060 (N_17060,N_8755,N_8503);
and U17061 (N_17061,N_10481,N_9165);
or U17062 (N_17062,N_7567,N_8365);
and U17063 (N_17063,N_9962,N_9901);
nand U17064 (N_17064,N_8173,N_8707);
or U17065 (N_17065,N_10060,N_11128);
or U17066 (N_17066,N_9247,N_8149);
nor U17067 (N_17067,N_9220,N_11144);
nand U17068 (N_17068,N_7112,N_7194);
and U17069 (N_17069,N_7516,N_10452);
xor U17070 (N_17070,N_10800,N_10544);
nand U17071 (N_17071,N_8776,N_9331);
nand U17072 (N_17072,N_10511,N_7597);
nand U17073 (N_17073,N_10809,N_8918);
nor U17074 (N_17074,N_9450,N_9184);
or U17075 (N_17075,N_7224,N_10188);
nand U17076 (N_17076,N_6493,N_6517);
nor U17077 (N_17077,N_7897,N_6089);
nand U17078 (N_17078,N_11578,N_9135);
xor U17079 (N_17079,N_11154,N_11841);
nand U17080 (N_17080,N_8039,N_6302);
xnor U17081 (N_17081,N_10679,N_6617);
and U17082 (N_17082,N_6393,N_11802);
nor U17083 (N_17083,N_8395,N_9850);
nand U17084 (N_17084,N_10112,N_10237);
nand U17085 (N_17085,N_11191,N_6762);
and U17086 (N_17086,N_8889,N_6086);
xor U17087 (N_17087,N_8936,N_11188);
and U17088 (N_17088,N_11669,N_7139);
and U17089 (N_17089,N_7534,N_6258);
and U17090 (N_17090,N_11831,N_9805);
xnor U17091 (N_17091,N_9001,N_9797);
nand U17092 (N_17092,N_6374,N_6601);
nor U17093 (N_17093,N_9096,N_8363);
nor U17094 (N_17094,N_11075,N_9296);
xnor U17095 (N_17095,N_10489,N_9856);
xnor U17096 (N_17096,N_8184,N_8549);
nor U17097 (N_17097,N_8412,N_11058);
xnor U17098 (N_17098,N_6626,N_6951);
and U17099 (N_17099,N_10684,N_9134);
or U17100 (N_17100,N_7248,N_11449);
and U17101 (N_17101,N_6511,N_10216);
nor U17102 (N_17102,N_7547,N_7467);
nand U17103 (N_17103,N_7191,N_9205);
nand U17104 (N_17104,N_6163,N_8836);
xor U17105 (N_17105,N_8455,N_11509);
and U17106 (N_17106,N_10472,N_11623);
xor U17107 (N_17107,N_7128,N_9036);
or U17108 (N_17108,N_10718,N_6339);
nor U17109 (N_17109,N_7427,N_11731);
nand U17110 (N_17110,N_8041,N_10914);
nand U17111 (N_17111,N_10372,N_8812);
and U17112 (N_17112,N_10781,N_11094);
nand U17113 (N_17113,N_9908,N_8897);
xnor U17114 (N_17114,N_9512,N_7240);
xnor U17115 (N_17115,N_6925,N_10980);
and U17116 (N_17116,N_6436,N_11220);
nand U17117 (N_17117,N_8107,N_9392);
or U17118 (N_17118,N_11964,N_10863);
xor U17119 (N_17119,N_10527,N_7740);
and U17120 (N_17120,N_10016,N_10716);
or U17121 (N_17121,N_8185,N_10902);
and U17122 (N_17122,N_6770,N_10105);
xnor U17123 (N_17123,N_10176,N_8571);
or U17124 (N_17124,N_10644,N_9860);
nand U17125 (N_17125,N_10942,N_6931);
xor U17126 (N_17126,N_6816,N_7663);
nor U17127 (N_17127,N_10453,N_10803);
nor U17128 (N_17128,N_10582,N_11353);
and U17129 (N_17129,N_8605,N_10361);
nor U17130 (N_17130,N_10191,N_7004);
nand U17131 (N_17131,N_9161,N_9835);
xor U17132 (N_17132,N_9491,N_7499);
nand U17133 (N_17133,N_11494,N_8230);
xor U17134 (N_17134,N_11048,N_8379);
or U17135 (N_17135,N_10047,N_11014);
or U17136 (N_17136,N_7968,N_10183);
nor U17137 (N_17137,N_6292,N_6966);
nand U17138 (N_17138,N_11825,N_8870);
xor U17139 (N_17139,N_8904,N_8679);
or U17140 (N_17140,N_6319,N_8359);
nand U17141 (N_17141,N_10009,N_10199);
or U17142 (N_17142,N_10303,N_7900);
and U17143 (N_17143,N_6162,N_10322);
nand U17144 (N_17144,N_8450,N_9590);
xor U17145 (N_17145,N_7587,N_9197);
or U17146 (N_17146,N_8763,N_6285);
nand U17147 (N_17147,N_10959,N_6892);
xor U17148 (N_17148,N_7429,N_8946);
and U17149 (N_17149,N_8880,N_8051);
nand U17150 (N_17150,N_9725,N_11009);
and U17151 (N_17151,N_7648,N_9429);
nand U17152 (N_17152,N_9546,N_9335);
or U17153 (N_17153,N_6242,N_10991);
or U17154 (N_17154,N_10189,N_7643);
or U17155 (N_17155,N_8886,N_8387);
xnor U17156 (N_17156,N_11976,N_6685);
or U17157 (N_17157,N_11476,N_9690);
or U17158 (N_17158,N_7237,N_6485);
and U17159 (N_17159,N_8045,N_8859);
and U17160 (N_17160,N_9416,N_10525);
and U17161 (N_17161,N_7774,N_8130);
nand U17162 (N_17162,N_7439,N_10245);
and U17163 (N_17163,N_6120,N_6427);
nand U17164 (N_17164,N_9683,N_6370);
xor U17165 (N_17165,N_7387,N_9266);
and U17166 (N_17166,N_9695,N_10439);
and U17167 (N_17167,N_9654,N_9389);
or U17168 (N_17168,N_10363,N_11226);
nand U17169 (N_17169,N_6088,N_10253);
or U17170 (N_17170,N_9498,N_8640);
and U17171 (N_17171,N_8199,N_9288);
xor U17172 (N_17172,N_11081,N_7741);
and U17173 (N_17173,N_9182,N_7593);
nor U17174 (N_17174,N_7024,N_7915);
nor U17175 (N_17175,N_10142,N_10197);
xor U17176 (N_17176,N_11435,N_7278);
or U17177 (N_17177,N_8799,N_8577);
and U17178 (N_17178,N_8071,N_8912);
nand U17179 (N_17179,N_6401,N_7312);
xnor U17180 (N_17180,N_8070,N_8958);
xor U17181 (N_17181,N_7472,N_9263);
or U17182 (N_17182,N_7852,N_11957);
xor U17183 (N_17183,N_11286,N_9320);
nand U17184 (N_17184,N_11836,N_9201);
nand U17185 (N_17185,N_8808,N_7556);
nor U17186 (N_17186,N_10710,N_8369);
nand U17187 (N_17187,N_10877,N_11301);
nor U17188 (N_17188,N_10761,N_8882);
nand U17189 (N_17189,N_11923,N_8758);
nor U17190 (N_17190,N_10772,N_11685);
and U17191 (N_17191,N_7995,N_7406);
nor U17192 (N_17192,N_6564,N_11236);
xnor U17193 (N_17193,N_9499,N_11906);
nand U17194 (N_17194,N_6879,N_6589);
and U17195 (N_17195,N_10335,N_9715);
and U17196 (N_17196,N_9695,N_11094);
or U17197 (N_17197,N_7433,N_6236);
xor U17198 (N_17198,N_9315,N_7057);
xor U17199 (N_17199,N_9897,N_11592);
nor U17200 (N_17200,N_7919,N_11707);
and U17201 (N_17201,N_8229,N_6184);
nor U17202 (N_17202,N_10651,N_8353);
and U17203 (N_17203,N_8903,N_8630);
nand U17204 (N_17204,N_9906,N_8857);
nand U17205 (N_17205,N_9339,N_8493);
and U17206 (N_17206,N_9810,N_11442);
nand U17207 (N_17207,N_9457,N_7104);
nor U17208 (N_17208,N_7955,N_9421);
nor U17209 (N_17209,N_11276,N_6890);
nor U17210 (N_17210,N_10468,N_7310);
or U17211 (N_17211,N_6376,N_6757);
nor U17212 (N_17212,N_8946,N_7616);
nand U17213 (N_17213,N_7246,N_10008);
and U17214 (N_17214,N_10393,N_9599);
nor U17215 (N_17215,N_11370,N_9188);
nand U17216 (N_17216,N_7051,N_7957);
nor U17217 (N_17217,N_10019,N_10334);
xor U17218 (N_17218,N_9299,N_6083);
nand U17219 (N_17219,N_6233,N_11085);
xnor U17220 (N_17220,N_10214,N_10110);
or U17221 (N_17221,N_6738,N_11331);
or U17222 (N_17222,N_10737,N_8796);
and U17223 (N_17223,N_9068,N_7073);
or U17224 (N_17224,N_11189,N_9946);
or U17225 (N_17225,N_6406,N_7042);
nand U17226 (N_17226,N_6181,N_10591);
nor U17227 (N_17227,N_6775,N_8592);
and U17228 (N_17228,N_9631,N_8553);
nand U17229 (N_17229,N_7342,N_11718);
nor U17230 (N_17230,N_6693,N_7139);
nor U17231 (N_17231,N_9050,N_10753);
and U17232 (N_17232,N_6146,N_8219);
or U17233 (N_17233,N_7484,N_8518);
xor U17234 (N_17234,N_6590,N_7689);
xor U17235 (N_17235,N_10795,N_6636);
or U17236 (N_17236,N_6130,N_11455);
nor U17237 (N_17237,N_8324,N_9410);
xor U17238 (N_17238,N_6263,N_11951);
or U17239 (N_17239,N_7675,N_6062);
or U17240 (N_17240,N_11288,N_11975);
and U17241 (N_17241,N_6534,N_9281);
and U17242 (N_17242,N_7007,N_8953);
nor U17243 (N_17243,N_10100,N_11697);
nor U17244 (N_17244,N_10588,N_11030);
or U17245 (N_17245,N_8526,N_6743);
nor U17246 (N_17246,N_7123,N_10608);
nor U17247 (N_17247,N_7481,N_10368);
xor U17248 (N_17248,N_6198,N_7882);
xor U17249 (N_17249,N_8366,N_10952);
and U17250 (N_17250,N_10776,N_11119);
or U17251 (N_17251,N_10739,N_10881);
and U17252 (N_17252,N_6213,N_6768);
xor U17253 (N_17253,N_10003,N_11109);
or U17254 (N_17254,N_9064,N_7112);
nand U17255 (N_17255,N_8513,N_11001);
nor U17256 (N_17256,N_6204,N_8588);
and U17257 (N_17257,N_11000,N_8772);
nor U17258 (N_17258,N_6306,N_8872);
nor U17259 (N_17259,N_6276,N_8939);
or U17260 (N_17260,N_9683,N_8642);
or U17261 (N_17261,N_10543,N_11902);
or U17262 (N_17262,N_6412,N_9385);
nor U17263 (N_17263,N_6689,N_7879);
or U17264 (N_17264,N_9607,N_8179);
or U17265 (N_17265,N_7691,N_7800);
nand U17266 (N_17266,N_6582,N_6091);
nor U17267 (N_17267,N_8815,N_7366);
or U17268 (N_17268,N_6910,N_6760);
xor U17269 (N_17269,N_7904,N_7076);
xnor U17270 (N_17270,N_7389,N_9315);
xor U17271 (N_17271,N_10699,N_7663);
and U17272 (N_17272,N_8991,N_9316);
xnor U17273 (N_17273,N_11014,N_10700);
and U17274 (N_17274,N_11954,N_8534);
xnor U17275 (N_17275,N_11903,N_6204);
xor U17276 (N_17276,N_7772,N_8992);
or U17277 (N_17277,N_7515,N_8500);
nand U17278 (N_17278,N_10021,N_8445);
xor U17279 (N_17279,N_9374,N_7122);
and U17280 (N_17280,N_10133,N_6719);
nand U17281 (N_17281,N_6409,N_11786);
and U17282 (N_17282,N_7122,N_6557);
xor U17283 (N_17283,N_8032,N_8560);
xnor U17284 (N_17284,N_9049,N_7483);
and U17285 (N_17285,N_9999,N_7661);
or U17286 (N_17286,N_10324,N_7942);
and U17287 (N_17287,N_8098,N_7207);
or U17288 (N_17288,N_10672,N_9885);
xnor U17289 (N_17289,N_11998,N_11144);
nand U17290 (N_17290,N_8542,N_8221);
nand U17291 (N_17291,N_7689,N_9999);
nand U17292 (N_17292,N_10978,N_11726);
xnor U17293 (N_17293,N_8356,N_9513);
and U17294 (N_17294,N_9952,N_10077);
xor U17295 (N_17295,N_10286,N_9216);
nor U17296 (N_17296,N_8940,N_10109);
or U17297 (N_17297,N_8634,N_10398);
nand U17298 (N_17298,N_7314,N_11250);
or U17299 (N_17299,N_11923,N_6335);
nand U17300 (N_17300,N_6456,N_10017);
or U17301 (N_17301,N_8624,N_7214);
and U17302 (N_17302,N_11581,N_6823);
nand U17303 (N_17303,N_7830,N_8743);
nand U17304 (N_17304,N_10728,N_10001);
nand U17305 (N_17305,N_6726,N_8191);
nand U17306 (N_17306,N_10838,N_6672);
and U17307 (N_17307,N_7779,N_8355);
and U17308 (N_17308,N_6809,N_10775);
nand U17309 (N_17309,N_11481,N_9438);
or U17310 (N_17310,N_8431,N_9040);
xor U17311 (N_17311,N_8047,N_10996);
xnor U17312 (N_17312,N_6156,N_9054);
xor U17313 (N_17313,N_7354,N_8653);
or U17314 (N_17314,N_7006,N_8403);
and U17315 (N_17315,N_6309,N_9724);
xnor U17316 (N_17316,N_6924,N_10956);
nor U17317 (N_17317,N_6405,N_9476);
or U17318 (N_17318,N_7031,N_6997);
or U17319 (N_17319,N_9373,N_9089);
xnor U17320 (N_17320,N_7434,N_7323);
and U17321 (N_17321,N_10252,N_11973);
xnor U17322 (N_17322,N_6072,N_8637);
nand U17323 (N_17323,N_9249,N_9650);
nor U17324 (N_17324,N_8738,N_8881);
xor U17325 (N_17325,N_8109,N_10223);
nand U17326 (N_17326,N_10979,N_10095);
or U17327 (N_17327,N_7123,N_9940);
nand U17328 (N_17328,N_7930,N_9048);
nor U17329 (N_17329,N_8177,N_6739);
or U17330 (N_17330,N_6835,N_7851);
and U17331 (N_17331,N_6498,N_10807);
and U17332 (N_17332,N_10072,N_11472);
nand U17333 (N_17333,N_8950,N_8288);
nand U17334 (N_17334,N_8455,N_7731);
nor U17335 (N_17335,N_8808,N_7664);
nor U17336 (N_17336,N_10206,N_9149);
or U17337 (N_17337,N_11292,N_8404);
xnor U17338 (N_17338,N_10946,N_10001);
and U17339 (N_17339,N_6567,N_9899);
xnor U17340 (N_17340,N_11539,N_7805);
xnor U17341 (N_17341,N_8683,N_6315);
xnor U17342 (N_17342,N_6448,N_7579);
nor U17343 (N_17343,N_11795,N_8624);
nand U17344 (N_17344,N_7775,N_6420);
xnor U17345 (N_17345,N_8125,N_6192);
xnor U17346 (N_17346,N_7383,N_8495);
or U17347 (N_17347,N_11474,N_10156);
or U17348 (N_17348,N_6545,N_6818);
nand U17349 (N_17349,N_8604,N_6366);
and U17350 (N_17350,N_11546,N_9941);
xnor U17351 (N_17351,N_11844,N_10451);
nand U17352 (N_17352,N_7813,N_8235);
and U17353 (N_17353,N_7507,N_9686);
or U17354 (N_17354,N_9031,N_10401);
and U17355 (N_17355,N_11939,N_9653);
nor U17356 (N_17356,N_7441,N_11860);
xor U17357 (N_17357,N_6053,N_11186);
xor U17358 (N_17358,N_9255,N_8843);
and U17359 (N_17359,N_10761,N_9566);
nor U17360 (N_17360,N_8273,N_10022);
and U17361 (N_17361,N_7294,N_7041);
and U17362 (N_17362,N_10917,N_9031);
nand U17363 (N_17363,N_9852,N_6885);
xor U17364 (N_17364,N_9925,N_10075);
or U17365 (N_17365,N_6226,N_9637);
xor U17366 (N_17366,N_6495,N_9350);
and U17367 (N_17367,N_6500,N_10064);
xnor U17368 (N_17368,N_7517,N_8566);
nor U17369 (N_17369,N_10342,N_10778);
nor U17370 (N_17370,N_10170,N_9155);
xnor U17371 (N_17371,N_10395,N_10584);
and U17372 (N_17372,N_9129,N_8268);
nor U17373 (N_17373,N_9030,N_9904);
xnor U17374 (N_17374,N_8476,N_10621);
nand U17375 (N_17375,N_9488,N_6226);
nand U17376 (N_17376,N_8022,N_11114);
or U17377 (N_17377,N_6495,N_9586);
and U17378 (N_17378,N_9510,N_8578);
nor U17379 (N_17379,N_9638,N_8377);
nand U17380 (N_17380,N_7031,N_9377);
nand U17381 (N_17381,N_10684,N_8089);
nand U17382 (N_17382,N_9876,N_9442);
xnor U17383 (N_17383,N_8813,N_6200);
nand U17384 (N_17384,N_7198,N_7257);
xnor U17385 (N_17385,N_10905,N_8863);
and U17386 (N_17386,N_11190,N_8117);
nand U17387 (N_17387,N_9373,N_8850);
nor U17388 (N_17388,N_9748,N_7051);
or U17389 (N_17389,N_8824,N_8353);
nor U17390 (N_17390,N_8699,N_6251);
or U17391 (N_17391,N_7523,N_11701);
nor U17392 (N_17392,N_6926,N_9201);
nand U17393 (N_17393,N_7079,N_8945);
and U17394 (N_17394,N_11773,N_10294);
nand U17395 (N_17395,N_10619,N_6519);
nand U17396 (N_17396,N_8317,N_8410);
nand U17397 (N_17397,N_8390,N_11823);
and U17398 (N_17398,N_7206,N_6359);
nand U17399 (N_17399,N_8899,N_9617);
nand U17400 (N_17400,N_9883,N_7076);
nor U17401 (N_17401,N_10512,N_6994);
and U17402 (N_17402,N_9193,N_7366);
nor U17403 (N_17403,N_7686,N_10893);
or U17404 (N_17404,N_8334,N_9129);
nor U17405 (N_17405,N_9984,N_6713);
nand U17406 (N_17406,N_8773,N_7909);
nand U17407 (N_17407,N_8011,N_7502);
or U17408 (N_17408,N_8348,N_6022);
or U17409 (N_17409,N_6858,N_10760);
nor U17410 (N_17410,N_11912,N_10089);
nor U17411 (N_17411,N_8431,N_10738);
or U17412 (N_17412,N_10665,N_10605);
and U17413 (N_17413,N_9815,N_8440);
nor U17414 (N_17414,N_11492,N_7640);
or U17415 (N_17415,N_11787,N_11752);
and U17416 (N_17416,N_9093,N_9910);
or U17417 (N_17417,N_6676,N_7868);
nand U17418 (N_17418,N_7285,N_9061);
nand U17419 (N_17419,N_8224,N_10498);
or U17420 (N_17420,N_6102,N_10736);
xnor U17421 (N_17421,N_6277,N_9710);
xor U17422 (N_17422,N_9514,N_10008);
or U17423 (N_17423,N_11179,N_8305);
nor U17424 (N_17424,N_10363,N_10650);
or U17425 (N_17425,N_10725,N_6516);
and U17426 (N_17426,N_8835,N_8541);
nand U17427 (N_17427,N_10339,N_9278);
nand U17428 (N_17428,N_11785,N_10509);
nor U17429 (N_17429,N_10755,N_11993);
nand U17430 (N_17430,N_6459,N_9923);
and U17431 (N_17431,N_8918,N_8585);
xor U17432 (N_17432,N_6663,N_9683);
nor U17433 (N_17433,N_6580,N_9487);
xor U17434 (N_17434,N_7100,N_8106);
xor U17435 (N_17435,N_6296,N_7462);
nand U17436 (N_17436,N_11741,N_7220);
and U17437 (N_17437,N_6493,N_7899);
and U17438 (N_17438,N_10522,N_8535);
nor U17439 (N_17439,N_10921,N_8986);
nand U17440 (N_17440,N_6589,N_8557);
and U17441 (N_17441,N_8630,N_7658);
xnor U17442 (N_17442,N_10596,N_7873);
or U17443 (N_17443,N_11743,N_7902);
nor U17444 (N_17444,N_10983,N_8127);
or U17445 (N_17445,N_8711,N_7648);
nor U17446 (N_17446,N_7088,N_8518);
nor U17447 (N_17447,N_7293,N_11416);
nand U17448 (N_17448,N_10617,N_6137);
or U17449 (N_17449,N_7489,N_10463);
nand U17450 (N_17450,N_8307,N_10354);
nand U17451 (N_17451,N_9365,N_10630);
and U17452 (N_17452,N_6287,N_7835);
nor U17453 (N_17453,N_8846,N_11623);
or U17454 (N_17454,N_10012,N_10331);
nand U17455 (N_17455,N_10132,N_7681);
xor U17456 (N_17456,N_7788,N_10647);
xor U17457 (N_17457,N_9096,N_6122);
xor U17458 (N_17458,N_9314,N_10344);
or U17459 (N_17459,N_8462,N_7562);
or U17460 (N_17460,N_8247,N_11886);
nor U17461 (N_17461,N_11619,N_7847);
nand U17462 (N_17462,N_10125,N_8976);
and U17463 (N_17463,N_11681,N_6855);
and U17464 (N_17464,N_6745,N_6537);
and U17465 (N_17465,N_10779,N_9248);
and U17466 (N_17466,N_6848,N_8515);
and U17467 (N_17467,N_6972,N_8846);
and U17468 (N_17468,N_8587,N_7056);
nor U17469 (N_17469,N_7796,N_6668);
nand U17470 (N_17470,N_9644,N_6681);
and U17471 (N_17471,N_7077,N_6372);
nand U17472 (N_17472,N_11456,N_7770);
nor U17473 (N_17473,N_9924,N_11777);
or U17474 (N_17474,N_10658,N_7095);
nand U17475 (N_17475,N_9289,N_10834);
nand U17476 (N_17476,N_11601,N_6564);
or U17477 (N_17477,N_6218,N_8594);
and U17478 (N_17478,N_11323,N_11378);
or U17479 (N_17479,N_9524,N_7772);
and U17480 (N_17480,N_10357,N_9048);
or U17481 (N_17481,N_9675,N_6363);
or U17482 (N_17482,N_9658,N_6086);
xor U17483 (N_17483,N_11938,N_10254);
nor U17484 (N_17484,N_6815,N_6491);
or U17485 (N_17485,N_6597,N_11508);
or U17486 (N_17486,N_7230,N_7350);
or U17487 (N_17487,N_10295,N_11913);
xnor U17488 (N_17488,N_7923,N_8099);
xnor U17489 (N_17489,N_8975,N_10936);
nor U17490 (N_17490,N_9308,N_7579);
xor U17491 (N_17491,N_11250,N_9593);
nand U17492 (N_17492,N_6365,N_7637);
and U17493 (N_17493,N_8328,N_11729);
nor U17494 (N_17494,N_10103,N_6374);
and U17495 (N_17495,N_6196,N_6723);
xor U17496 (N_17496,N_9297,N_7196);
xor U17497 (N_17497,N_11320,N_9460);
and U17498 (N_17498,N_8516,N_8870);
nand U17499 (N_17499,N_9667,N_9670);
xor U17500 (N_17500,N_8015,N_6386);
nor U17501 (N_17501,N_8527,N_9976);
or U17502 (N_17502,N_10943,N_6880);
xor U17503 (N_17503,N_6379,N_6262);
nor U17504 (N_17504,N_6490,N_9645);
xnor U17505 (N_17505,N_7139,N_11904);
nor U17506 (N_17506,N_9304,N_8184);
nand U17507 (N_17507,N_9825,N_11989);
or U17508 (N_17508,N_10350,N_10419);
nand U17509 (N_17509,N_6809,N_11066);
and U17510 (N_17510,N_7335,N_10244);
xnor U17511 (N_17511,N_6211,N_8270);
nand U17512 (N_17512,N_9622,N_6693);
and U17513 (N_17513,N_10676,N_7559);
xor U17514 (N_17514,N_9762,N_9281);
or U17515 (N_17515,N_11184,N_9451);
or U17516 (N_17516,N_10183,N_8467);
xnor U17517 (N_17517,N_7022,N_9133);
or U17518 (N_17518,N_6008,N_6309);
xnor U17519 (N_17519,N_6829,N_7566);
nor U17520 (N_17520,N_8635,N_6658);
and U17521 (N_17521,N_9013,N_9319);
nor U17522 (N_17522,N_6324,N_10580);
or U17523 (N_17523,N_6613,N_10902);
xnor U17524 (N_17524,N_7868,N_9356);
xnor U17525 (N_17525,N_11276,N_10236);
nand U17526 (N_17526,N_7003,N_10434);
nand U17527 (N_17527,N_8418,N_10038);
xor U17528 (N_17528,N_9739,N_6897);
or U17529 (N_17529,N_11626,N_10388);
and U17530 (N_17530,N_6025,N_8191);
nor U17531 (N_17531,N_6587,N_8402);
nand U17532 (N_17532,N_10275,N_6758);
nand U17533 (N_17533,N_6705,N_7853);
nand U17534 (N_17534,N_6232,N_8451);
xor U17535 (N_17535,N_7677,N_11377);
nor U17536 (N_17536,N_10394,N_8431);
xor U17537 (N_17537,N_10275,N_11008);
and U17538 (N_17538,N_11178,N_8529);
xnor U17539 (N_17539,N_11502,N_7500);
nand U17540 (N_17540,N_8021,N_9449);
and U17541 (N_17541,N_10375,N_6730);
nor U17542 (N_17542,N_10327,N_8703);
nor U17543 (N_17543,N_9995,N_7053);
nand U17544 (N_17544,N_8164,N_7124);
or U17545 (N_17545,N_10784,N_10961);
and U17546 (N_17546,N_8307,N_9323);
xor U17547 (N_17547,N_7965,N_11759);
and U17548 (N_17548,N_6293,N_9428);
nand U17549 (N_17549,N_8252,N_7003);
nor U17550 (N_17550,N_11140,N_9446);
or U17551 (N_17551,N_8745,N_7274);
or U17552 (N_17552,N_7285,N_7229);
and U17553 (N_17553,N_11857,N_10653);
xnor U17554 (N_17554,N_7666,N_9089);
or U17555 (N_17555,N_6134,N_8629);
or U17556 (N_17556,N_11352,N_11603);
and U17557 (N_17557,N_9362,N_7539);
nor U17558 (N_17558,N_6978,N_6715);
xor U17559 (N_17559,N_9216,N_9207);
or U17560 (N_17560,N_6626,N_11611);
nor U17561 (N_17561,N_11882,N_9502);
and U17562 (N_17562,N_10368,N_8983);
or U17563 (N_17563,N_9056,N_6252);
xor U17564 (N_17564,N_8556,N_6689);
nor U17565 (N_17565,N_8817,N_7860);
and U17566 (N_17566,N_6516,N_8711);
nand U17567 (N_17567,N_10268,N_9624);
nand U17568 (N_17568,N_10251,N_8049);
nor U17569 (N_17569,N_11855,N_11430);
and U17570 (N_17570,N_7823,N_7045);
xnor U17571 (N_17571,N_8380,N_8812);
xor U17572 (N_17572,N_10106,N_9477);
nand U17573 (N_17573,N_10369,N_11071);
nand U17574 (N_17574,N_6670,N_6028);
and U17575 (N_17575,N_6331,N_9324);
or U17576 (N_17576,N_8888,N_6179);
and U17577 (N_17577,N_6730,N_6665);
nor U17578 (N_17578,N_7724,N_6684);
or U17579 (N_17579,N_6956,N_7818);
and U17580 (N_17580,N_11958,N_8955);
xnor U17581 (N_17581,N_10229,N_9173);
or U17582 (N_17582,N_8463,N_7943);
or U17583 (N_17583,N_10041,N_6059);
and U17584 (N_17584,N_10396,N_11881);
xnor U17585 (N_17585,N_6424,N_6413);
nor U17586 (N_17586,N_10835,N_8606);
nand U17587 (N_17587,N_6452,N_6219);
nand U17588 (N_17588,N_10433,N_9428);
nor U17589 (N_17589,N_9862,N_10254);
or U17590 (N_17590,N_11555,N_10565);
nand U17591 (N_17591,N_8244,N_8813);
nand U17592 (N_17592,N_10233,N_10862);
nand U17593 (N_17593,N_9549,N_9848);
nor U17594 (N_17594,N_6572,N_11379);
xnor U17595 (N_17595,N_11188,N_7457);
or U17596 (N_17596,N_10039,N_8192);
nor U17597 (N_17597,N_6039,N_8065);
nand U17598 (N_17598,N_11171,N_11563);
and U17599 (N_17599,N_7332,N_8058);
nor U17600 (N_17600,N_6011,N_7469);
and U17601 (N_17601,N_8279,N_8373);
nand U17602 (N_17602,N_7452,N_7899);
or U17603 (N_17603,N_10138,N_10555);
nand U17604 (N_17604,N_6625,N_8611);
and U17605 (N_17605,N_6339,N_6282);
and U17606 (N_17606,N_6329,N_11575);
xor U17607 (N_17607,N_10731,N_10442);
nand U17608 (N_17608,N_7339,N_7538);
xnor U17609 (N_17609,N_10541,N_10858);
xnor U17610 (N_17610,N_6952,N_8213);
and U17611 (N_17611,N_11347,N_7064);
xor U17612 (N_17612,N_10392,N_9964);
nor U17613 (N_17613,N_7328,N_11119);
nand U17614 (N_17614,N_7386,N_6960);
or U17615 (N_17615,N_9100,N_9237);
nand U17616 (N_17616,N_10639,N_9083);
and U17617 (N_17617,N_10737,N_6030);
nand U17618 (N_17618,N_9480,N_11977);
or U17619 (N_17619,N_6917,N_8653);
xor U17620 (N_17620,N_8963,N_6301);
xor U17621 (N_17621,N_7278,N_11197);
nand U17622 (N_17622,N_8176,N_9439);
and U17623 (N_17623,N_6769,N_9328);
nor U17624 (N_17624,N_7651,N_9368);
xnor U17625 (N_17625,N_11548,N_8175);
and U17626 (N_17626,N_7675,N_9573);
and U17627 (N_17627,N_7496,N_9491);
nand U17628 (N_17628,N_8015,N_10248);
nor U17629 (N_17629,N_10744,N_11443);
nor U17630 (N_17630,N_10621,N_9025);
nor U17631 (N_17631,N_8522,N_8216);
nand U17632 (N_17632,N_11090,N_8303);
and U17633 (N_17633,N_6242,N_10212);
nor U17634 (N_17634,N_10421,N_11801);
and U17635 (N_17635,N_7946,N_9593);
and U17636 (N_17636,N_11469,N_9872);
xor U17637 (N_17637,N_7528,N_10742);
or U17638 (N_17638,N_8972,N_7574);
xnor U17639 (N_17639,N_11058,N_6670);
nand U17640 (N_17640,N_6057,N_8695);
or U17641 (N_17641,N_7688,N_9010);
xor U17642 (N_17642,N_10986,N_11127);
and U17643 (N_17643,N_8647,N_8315);
xnor U17644 (N_17644,N_8628,N_7264);
or U17645 (N_17645,N_6450,N_8938);
nor U17646 (N_17646,N_9595,N_7255);
or U17647 (N_17647,N_7827,N_6384);
and U17648 (N_17648,N_6344,N_8677);
nand U17649 (N_17649,N_6295,N_10986);
nor U17650 (N_17650,N_8853,N_11141);
and U17651 (N_17651,N_10018,N_11967);
or U17652 (N_17652,N_6523,N_11560);
or U17653 (N_17653,N_6983,N_6973);
nand U17654 (N_17654,N_9280,N_9719);
nor U17655 (N_17655,N_8123,N_11467);
xnor U17656 (N_17656,N_9581,N_9239);
or U17657 (N_17657,N_10348,N_11212);
or U17658 (N_17658,N_8519,N_9750);
nand U17659 (N_17659,N_8223,N_10238);
and U17660 (N_17660,N_11529,N_9073);
xor U17661 (N_17661,N_6981,N_11306);
xnor U17662 (N_17662,N_11299,N_10263);
or U17663 (N_17663,N_6260,N_8394);
and U17664 (N_17664,N_10239,N_11143);
nand U17665 (N_17665,N_6179,N_10909);
and U17666 (N_17666,N_6257,N_9253);
nand U17667 (N_17667,N_9861,N_8184);
and U17668 (N_17668,N_10560,N_9854);
nand U17669 (N_17669,N_10527,N_8069);
and U17670 (N_17670,N_10909,N_6824);
or U17671 (N_17671,N_6274,N_9242);
nor U17672 (N_17672,N_6440,N_8404);
and U17673 (N_17673,N_9249,N_7437);
xnor U17674 (N_17674,N_6255,N_7926);
or U17675 (N_17675,N_11428,N_11826);
nor U17676 (N_17676,N_7996,N_7677);
and U17677 (N_17677,N_9459,N_10850);
nand U17678 (N_17678,N_11040,N_6762);
and U17679 (N_17679,N_9065,N_9451);
nor U17680 (N_17680,N_6405,N_6292);
or U17681 (N_17681,N_10846,N_8168);
or U17682 (N_17682,N_9178,N_7058);
or U17683 (N_17683,N_11208,N_10061);
xor U17684 (N_17684,N_11020,N_6365);
nand U17685 (N_17685,N_6615,N_7090);
or U17686 (N_17686,N_6747,N_7028);
nor U17687 (N_17687,N_10616,N_11157);
nand U17688 (N_17688,N_9801,N_7977);
or U17689 (N_17689,N_7859,N_9003);
nand U17690 (N_17690,N_11266,N_7767);
xor U17691 (N_17691,N_8015,N_10191);
nor U17692 (N_17692,N_7417,N_7258);
xor U17693 (N_17693,N_7986,N_7241);
xor U17694 (N_17694,N_9306,N_9240);
xor U17695 (N_17695,N_7314,N_9121);
xnor U17696 (N_17696,N_10827,N_8266);
nand U17697 (N_17697,N_7965,N_11231);
or U17698 (N_17698,N_6422,N_8012);
nand U17699 (N_17699,N_6025,N_7664);
xnor U17700 (N_17700,N_6456,N_6119);
or U17701 (N_17701,N_8212,N_8117);
nor U17702 (N_17702,N_9723,N_8420);
and U17703 (N_17703,N_8116,N_8547);
and U17704 (N_17704,N_8076,N_8170);
xnor U17705 (N_17705,N_11242,N_8496);
xor U17706 (N_17706,N_7828,N_8184);
xnor U17707 (N_17707,N_7699,N_11955);
nor U17708 (N_17708,N_11667,N_6973);
or U17709 (N_17709,N_8988,N_7288);
and U17710 (N_17710,N_6822,N_10342);
xor U17711 (N_17711,N_10843,N_6525);
and U17712 (N_17712,N_9103,N_10847);
xnor U17713 (N_17713,N_9376,N_10488);
and U17714 (N_17714,N_10597,N_9746);
and U17715 (N_17715,N_11844,N_7061);
or U17716 (N_17716,N_6698,N_9480);
or U17717 (N_17717,N_9612,N_10813);
or U17718 (N_17718,N_7645,N_6557);
xor U17719 (N_17719,N_9786,N_8255);
or U17720 (N_17720,N_11570,N_11910);
nand U17721 (N_17721,N_8779,N_9763);
nand U17722 (N_17722,N_10834,N_6715);
nor U17723 (N_17723,N_9139,N_11777);
and U17724 (N_17724,N_7521,N_6801);
nor U17725 (N_17725,N_9667,N_11878);
nand U17726 (N_17726,N_7743,N_11975);
xor U17727 (N_17727,N_7378,N_6048);
and U17728 (N_17728,N_8220,N_11515);
xnor U17729 (N_17729,N_7414,N_7966);
xor U17730 (N_17730,N_8805,N_8385);
or U17731 (N_17731,N_7064,N_7464);
and U17732 (N_17732,N_11632,N_11234);
or U17733 (N_17733,N_6592,N_10302);
xor U17734 (N_17734,N_6730,N_8986);
or U17735 (N_17735,N_8559,N_10132);
nor U17736 (N_17736,N_10038,N_8086);
xor U17737 (N_17737,N_7892,N_11841);
or U17738 (N_17738,N_10453,N_10950);
nor U17739 (N_17739,N_7862,N_9310);
or U17740 (N_17740,N_6250,N_11539);
nor U17741 (N_17741,N_11751,N_6191);
or U17742 (N_17742,N_6735,N_7986);
and U17743 (N_17743,N_11549,N_9591);
and U17744 (N_17744,N_7309,N_8642);
and U17745 (N_17745,N_6082,N_11456);
and U17746 (N_17746,N_6178,N_8442);
nand U17747 (N_17747,N_10881,N_7928);
and U17748 (N_17748,N_10461,N_10472);
nor U17749 (N_17749,N_7445,N_9278);
nor U17750 (N_17750,N_8359,N_8230);
and U17751 (N_17751,N_6202,N_6517);
nor U17752 (N_17752,N_8231,N_7850);
nor U17753 (N_17753,N_11191,N_6680);
or U17754 (N_17754,N_11974,N_11007);
or U17755 (N_17755,N_8421,N_8952);
nand U17756 (N_17756,N_7300,N_8200);
and U17757 (N_17757,N_8004,N_8203);
and U17758 (N_17758,N_7004,N_6026);
xnor U17759 (N_17759,N_8843,N_8355);
and U17760 (N_17760,N_6467,N_10767);
nor U17761 (N_17761,N_10510,N_6674);
nand U17762 (N_17762,N_11130,N_11707);
nor U17763 (N_17763,N_7106,N_11714);
nand U17764 (N_17764,N_7963,N_11974);
nor U17765 (N_17765,N_6379,N_8295);
nand U17766 (N_17766,N_10720,N_9467);
nor U17767 (N_17767,N_6243,N_11414);
or U17768 (N_17768,N_11377,N_11160);
nor U17769 (N_17769,N_9609,N_8230);
and U17770 (N_17770,N_9409,N_6344);
nor U17771 (N_17771,N_6417,N_11235);
and U17772 (N_17772,N_10014,N_7308);
nand U17773 (N_17773,N_8173,N_7554);
nand U17774 (N_17774,N_6683,N_9185);
nor U17775 (N_17775,N_9686,N_6552);
nor U17776 (N_17776,N_8804,N_6291);
and U17777 (N_17777,N_11111,N_6476);
nand U17778 (N_17778,N_9459,N_8785);
and U17779 (N_17779,N_6153,N_7241);
nand U17780 (N_17780,N_9142,N_6371);
or U17781 (N_17781,N_9090,N_9339);
nor U17782 (N_17782,N_7882,N_10741);
and U17783 (N_17783,N_7023,N_11748);
nor U17784 (N_17784,N_6375,N_7888);
or U17785 (N_17785,N_6915,N_11175);
nor U17786 (N_17786,N_8116,N_11851);
xor U17787 (N_17787,N_8449,N_7751);
xor U17788 (N_17788,N_11190,N_9195);
xor U17789 (N_17789,N_6822,N_9586);
and U17790 (N_17790,N_8407,N_10026);
nor U17791 (N_17791,N_8631,N_8361);
nor U17792 (N_17792,N_8231,N_10472);
xnor U17793 (N_17793,N_7975,N_7996);
and U17794 (N_17794,N_7559,N_11658);
or U17795 (N_17795,N_9972,N_9327);
nand U17796 (N_17796,N_9805,N_7847);
xor U17797 (N_17797,N_11975,N_6780);
nand U17798 (N_17798,N_8898,N_9145);
nor U17799 (N_17799,N_7419,N_6016);
and U17800 (N_17800,N_8436,N_7393);
or U17801 (N_17801,N_7738,N_9155);
or U17802 (N_17802,N_11579,N_7996);
xor U17803 (N_17803,N_9844,N_8862);
or U17804 (N_17804,N_9183,N_10205);
nand U17805 (N_17805,N_7780,N_10716);
or U17806 (N_17806,N_6470,N_8917);
and U17807 (N_17807,N_11342,N_10838);
or U17808 (N_17808,N_8270,N_10347);
nor U17809 (N_17809,N_8874,N_6521);
or U17810 (N_17810,N_10441,N_6938);
nor U17811 (N_17811,N_8483,N_7434);
nand U17812 (N_17812,N_6139,N_9803);
nor U17813 (N_17813,N_6096,N_7436);
and U17814 (N_17814,N_7789,N_8956);
and U17815 (N_17815,N_6387,N_6105);
nand U17816 (N_17816,N_9073,N_8078);
or U17817 (N_17817,N_10159,N_6759);
or U17818 (N_17818,N_7633,N_10770);
nor U17819 (N_17819,N_8252,N_10665);
and U17820 (N_17820,N_8850,N_7730);
xnor U17821 (N_17821,N_9329,N_11919);
and U17822 (N_17822,N_11350,N_9187);
xnor U17823 (N_17823,N_6312,N_10610);
and U17824 (N_17824,N_11909,N_10232);
nand U17825 (N_17825,N_7893,N_9636);
xor U17826 (N_17826,N_6899,N_9613);
or U17827 (N_17827,N_10983,N_10703);
and U17828 (N_17828,N_6154,N_8703);
xor U17829 (N_17829,N_6648,N_9094);
nand U17830 (N_17830,N_11925,N_9135);
xor U17831 (N_17831,N_11111,N_11432);
and U17832 (N_17832,N_10488,N_10477);
and U17833 (N_17833,N_6391,N_8978);
xnor U17834 (N_17834,N_8260,N_6933);
nor U17835 (N_17835,N_9753,N_10386);
and U17836 (N_17836,N_10566,N_6234);
or U17837 (N_17837,N_7914,N_7714);
or U17838 (N_17838,N_8054,N_9547);
nor U17839 (N_17839,N_6839,N_10750);
xnor U17840 (N_17840,N_8337,N_10275);
nor U17841 (N_17841,N_6404,N_11845);
xnor U17842 (N_17842,N_7094,N_6614);
xor U17843 (N_17843,N_7308,N_8140);
xor U17844 (N_17844,N_7703,N_9563);
nand U17845 (N_17845,N_8359,N_8026);
nand U17846 (N_17846,N_11032,N_7997);
xnor U17847 (N_17847,N_6606,N_6161);
or U17848 (N_17848,N_8188,N_7365);
xnor U17849 (N_17849,N_9421,N_8323);
and U17850 (N_17850,N_10541,N_9430);
and U17851 (N_17851,N_7532,N_7491);
xor U17852 (N_17852,N_10135,N_9209);
nand U17853 (N_17853,N_7323,N_11311);
and U17854 (N_17854,N_11677,N_10285);
xnor U17855 (N_17855,N_10346,N_8351);
xor U17856 (N_17856,N_7955,N_7627);
xor U17857 (N_17857,N_6492,N_10060);
nor U17858 (N_17858,N_10913,N_6629);
and U17859 (N_17859,N_9142,N_11928);
xor U17860 (N_17860,N_11074,N_11242);
or U17861 (N_17861,N_6843,N_9172);
nand U17862 (N_17862,N_6518,N_8749);
or U17863 (N_17863,N_10842,N_8505);
nand U17864 (N_17864,N_7719,N_8064);
nand U17865 (N_17865,N_10648,N_10722);
xnor U17866 (N_17866,N_11888,N_8920);
nand U17867 (N_17867,N_7128,N_11072);
nand U17868 (N_17868,N_8324,N_7508);
and U17869 (N_17869,N_6259,N_8563);
nand U17870 (N_17870,N_10836,N_8126);
and U17871 (N_17871,N_10753,N_6643);
xnor U17872 (N_17872,N_7297,N_10217);
xor U17873 (N_17873,N_8756,N_6384);
xor U17874 (N_17874,N_10010,N_9660);
and U17875 (N_17875,N_8055,N_10294);
xor U17876 (N_17876,N_11001,N_7468);
xor U17877 (N_17877,N_8974,N_8859);
and U17878 (N_17878,N_8408,N_7746);
and U17879 (N_17879,N_10771,N_10862);
nor U17880 (N_17880,N_9042,N_11114);
nand U17881 (N_17881,N_9526,N_11375);
xor U17882 (N_17882,N_6234,N_6818);
nor U17883 (N_17883,N_6764,N_8265);
or U17884 (N_17884,N_10769,N_9209);
or U17885 (N_17885,N_9571,N_8744);
and U17886 (N_17886,N_11806,N_8224);
nor U17887 (N_17887,N_10395,N_8815);
nor U17888 (N_17888,N_8148,N_9775);
xor U17889 (N_17889,N_9676,N_7163);
nand U17890 (N_17890,N_10416,N_10438);
xor U17891 (N_17891,N_6464,N_11674);
xnor U17892 (N_17892,N_10039,N_6924);
xnor U17893 (N_17893,N_10325,N_11589);
nor U17894 (N_17894,N_11807,N_7835);
nand U17895 (N_17895,N_10507,N_11079);
xnor U17896 (N_17896,N_8636,N_11471);
xnor U17897 (N_17897,N_10955,N_11361);
and U17898 (N_17898,N_9711,N_7680);
and U17899 (N_17899,N_11643,N_7631);
xor U17900 (N_17900,N_11160,N_7732);
nand U17901 (N_17901,N_6285,N_9122);
and U17902 (N_17902,N_9560,N_6205);
or U17903 (N_17903,N_10190,N_11786);
nor U17904 (N_17904,N_8824,N_8867);
nand U17905 (N_17905,N_7238,N_6291);
and U17906 (N_17906,N_9294,N_8469);
or U17907 (N_17907,N_11282,N_6566);
nand U17908 (N_17908,N_8752,N_7039);
xnor U17909 (N_17909,N_6434,N_9792);
nand U17910 (N_17910,N_9535,N_11006);
nor U17911 (N_17911,N_7597,N_11977);
or U17912 (N_17912,N_7227,N_6066);
nand U17913 (N_17913,N_11471,N_8795);
nor U17914 (N_17914,N_6413,N_7068);
xor U17915 (N_17915,N_10566,N_7638);
xor U17916 (N_17916,N_9899,N_9927);
xor U17917 (N_17917,N_8796,N_11063);
or U17918 (N_17918,N_6315,N_8362);
nand U17919 (N_17919,N_7807,N_7632);
xnor U17920 (N_17920,N_10088,N_8667);
xnor U17921 (N_17921,N_10724,N_7310);
nor U17922 (N_17922,N_9915,N_9225);
nand U17923 (N_17923,N_7275,N_10122);
or U17924 (N_17924,N_11249,N_9813);
xor U17925 (N_17925,N_10553,N_11504);
nor U17926 (N_17926,N_6999,N_6514);
nand U17927 (N_17927,N_6875,N_8826);
or U17928 (N_17928,N_8528,N_9289);
xor U17929 (N_17929,N_10847,N_10963);
and U17930 (N_17930,N_10938,N_8008);
and U17931 (N_17931,N_6527,N_7540);
or U17932 (N_17932,N_11440,N_7384);
and U17933 (N_17933,N_9905,N_6760);
nand U17934 (N_17934,N_6844,N_7991);
and U17935 (N_17935,N_11288,N_7091);
xnor U17936 (N_17936,N_7526,N_11927);
nor U17937 (N_17937,N_7814,N_10767);
or U17938 (N_17938,N_11674,N_9261);
nor U17939 (N_17939,N_9973,N_11492);
nor U17940 (N_17940,N_7792,N_11058);
nand U17941 (N_17941,N_7545,N_10238);
nand U17942 (N_17942,N_7079,N_10682);
nand U17943 (N_17943,N_9271,N_8143);
or U17944 (N_17944,N_11191,N_11488);
nor U17945 (N_17945,N_7019,N_7235);
nand U17946 (N_17946,N_10382,N_10662);
and U17947 (N_17947,N_8541,N_7273);
or U17948 (N_17948,N_6504,N_11792);
nand U17949 (N_17949,N_10044,N_11781);
or U17950 (N_17950,N_9039,N_9419);
or U17951 (N_17951,N_8887,N_9297);
nand U17952 (N_17952,N_11288,N_11378);
nand U17953 (N_17953,N_9166,N_9569);
nand U17954 (N_17954,N_9144,N_11431);
nand U17955 (N_17955,N_9070,N_11644);
and U17956 (N_17956,N_7537,N_9235);
and U17957 (N_17957,N_7168,N_7616);
nor U17958 (N_17958,N_6351,N_7871);
xor U17959 (N_17959,N_10639,N_7575);
nand U17960 (N_17960,N_7320,N_10857);
or U17961 (N_17961,N_6974,N_7419);
nand U17962 (N_17962,N_9726,N_9271);
nor U17963 (N_17963,N_10102,N_6981);
nor U17964 (N_17964,N_7346,N_10403);
and U17965 (N_17965,N_10236,N_9205);
or U17966 (N_17966,N_8676,N_10565);
or U17967 (N_17967,N_11351,N_11635);
xnor U17968 (N_17968,N_11011,N_9322);
and U17969 (N_17969,N_6819,N_7057);
nand U17970 (N_17970,N_10361,N_6227);
or U17971 (N_17971,N_8552,N_11517);
xor U17972 (N_17972,N_8527,N_7561);
xor U17973 (N_17973,N_9186,N_7817);
nand U17974 (N_17974,N_6852,N_7505);
and U17975 (N_17975,N_11311,N_11910);
xnor U17976 (N_17976,N_11751,N_8415);
and U17977 (N_17977,N_10389,N_6564);
or U17978 (N_17978,N_11471,N_7931);
nand U17979 (N_17979,N_7446,N_8806);
nand U17980 (N_17980,N_7985,N_11870);
xnor U17981 (N_17981,N_11786,N_9713);
and U17982 (N_17982,N_11904,N_8678);
nor U17983 (N_17983,N_9429,N_8412);
or U17984 (N_17984,N_7888,N_9305);
xnor U17985 (N_17985,N_8215,N_10602);
or U17986 (N_17986,N_10221,N_10529);
xor U17987 (N_17987,N_9337,N_7618);
nand U17988 (N_17988,N_8930,N_8856);
nand U17989 (N_17989,N_6289,N_7375);
nor U17990 (N_17990,N_10618,N_9526);
or U17991 (N_17991,N_11198,N_9006);
or U17992 (N_17992,N_6798,N_11223);
nor U17993 (N_17993,N_8913,N_6739);
nor U17994 (N_17994,N_6730,N_7956);
xnor U17995 (N_17995,N_10039,N_9865);
or U17996 (N_17996,N_6027,N_7009);
or U17997 (N_17997,N_7176,N_6954);
xor U17998 (N_17998,N_9148,N_10439);
or U17999 (N_17999,N_9039,N_10510);
xor U18000 (N_18000,N_12580,N_14700);
or U18001 (N_18001,N_16099,N_12329);
or U18002 (N_18002,N_14436,N_17578);
nor U18003 (N_18003,N_14874,N_14721);
nand U18004 (N_18004,N_17681,N_14279);
xnor U18005 (N_18005,N_14510,N_17141);
nor U18006 (N_18006,N_17403,N_14878);
xnor U18007 (N_18007,N_14785,N_13222);
nor U18008 (N_18008,N_13633,N_12237);
nor U18009 (N_18009,N_17039,N_12036);
and U18010 (N_18010,N_15333,N_16675);
and U18011 (N_18011,N_15982,N_14630);
xnor U18012 (N_18012,N_17267,N_14895);
xor U18013 (N_18013,N_15086,N_17268);
nor U18014 (N_18014,N_14343,N_17646);
and U18015 (N_18015,N_15037,N_16894);
nand U18016 (N_18016,N_16420,N_15466);
and U18017 (N_18017,N_15379,N_16118);
or U18018 (N_18018,N_17044,N_16710);
and U18019 (N_18019,N_12046,N_16867);
nor U18020 (N_18020,N_15815,N_16276);
nor U18021 (N_18021,N_14003,N_13388);
and U18022 (N_18022,N_12570,N_13022);
xor U18023 (N_18023,N_14983,N_17003);
nand U18024 (N_18024,N_14586,N_17256);
or U18025 (N_18025,N_17189,N_13260);
nand U18026 (N_18026,N_13587,N_13722);
or U18027 (N_18027,N_17532,N_15433);
nand U18028 (N_18028,N_16608,N_14398);
xnor U18029 (N_18029,N_16011,N_13870);
nor U18030 (N_18030,N_13818,N_17880);
and U18031 (N_18031,N_12886,N_13049);
xor U18032 (N_18032,N_13750,N_13980);
and U18033 (N_18033,N_16264,N_13615);
xnor U18034 (N_18034,N_15285,N_16392);
or U18035 (N_18035,N_12736,N_16226);
or U18036 (N_18036,N_15422,N_13531);
and U18037 (N_18037,N_16804,N_13868);
and U18038 (N_18038,N_15762,N_14024);
or U18039 (N_18039,N_14697,N_15563);
or U18040 (N_18040,N_16525,N_15432);
and U18041 (N_18041,N_16881,N_17414);
and U18042 (N_18042,N_13618,N_16468);
and U18043 (N_18043,N_14318,N_15358);
nor U18044 (N_18044,N_13788,N_16232);
or U18045 (N_18045,N_15720,N_13895);
nand U18046 (N_18046,N_12400,N_14396);
xnor U18047 (N_18047,N_14876,N_14899);
nand U18048 (N_18048,N_13632,N_17778);
nand U18049 (N_18049,N_16559,N_17989);
and U18050 (N_18050,N_16012,N_16170);
or U18051 (N_18051,N_14189,N_14817);
nor U18052 (N_18052,N_12838,N_17126);
or U18053 (N_18053,N_17294,N_16152);
nor U18054 (N_18054,N_12070,N_17672);
or U18055 (N_18055,N_12725,N_15420);
xnor U18056 (N_18056,N_13440,N_15146);
nand U18057 (N_18057,N_15745,N_13014);
xnor U18058 (N_18058,N_13904,N_16518);
or U18059 (N_18059,N_13240,N_16641);
nor U18060 (N_18060,N_13918,N_13626);
or U18061 (N_18061,N_14506,N_12303);
nor U18062 (N_18062,N_12941,N_13664);
or U18063 (N_18063,N_16906,N_16619);
and U18064 (N_18064,N_14654,N_15095);
xnor U18065 (N_18065,N_14159,N_15766);
nand U18066 (N_18066,N_13566,N_16854);
xnor U18067 (N_18067,N_17412,N_16485);
xor U18068 (N_18068,N_14511,N_17786);
xor U18069 (N_18069,N_16108,N_17645);
xnor U18070 (N_18070,N_12388,N_16741);
or U18071 (N_18071,N_13371,N_15131);
or U18072 (N_18072,N_13408,N_14245);
xor U18073 (N_18073,N_12948,N_16610);
or U18074 (N_18074,N_14968,N_15518);
nor U18075 (N_18075,N_14941,N_15243);
nand U18076 (N_18076,N_14681,N_12463);
nor U18077 (N_18077,N_16959,N_16960);
or U18078 (N_18078,N_13699,N_12998);
nand U18079 (N_18079,N_14080,N_17378);
xnor U18080 (N_18080,N_15010,N_16127);
nor U18081 (N_18081,N_12245,N_17840);
xnor U18082 (N_18082,N_16712,N_14629);
or U18083 (N_18083,N_13537,N_12997);
or U18084 (N_18084,N_16687,N_12233);
nand U18085 (N_18085,N_13840,N_15625);
nor U18086 (N_18086,N_16928,N_16647);
nor U18087 (N_18087,N_13842,N_12806);
nor U18088 (N_18088,N_15942,N_14621);
and U18089 (N_18089,N_17619,N_17607);
nor U18090 (N_18090,N_17022,N_12839);
or U18091 (N_18091,N_13161,N_12354);
and U18092 (N_18092,N_13053,N_16972);
or U18093 (N_18093,N_13561,N_13469);
xnor U18094 (N_18094,N_13090,N_16387);
or U18095 (N_18095,N_12113,N_14139);
nand U18096 (N_18096,N_17517,N_16184);
nand U18097 (N_18097,N_12572,N_14787);
xnor U18098 (N_18098,N_15101,N_16351);
and U18099 (N_18099,N_15620,N_14407);
and U18100 (N_18100,N_12430,N_12207);
or U18101 (N_18101,N_15427,N_12334);
xnor U18102 (N_18102,N_12232,N_12539);
xnor U18103 (N_18103,N_13644,N_13267);
and U18104 (N_18104,N_16173,N_12314);
or U18105 (N_18105,N_13019,N_16775);
or U18106 (N_18106,N_16103,N_15393);
nor U18107 (N_18107,N_14091,N_13326);
xor U18108 (N_18108,N_17207,N_16191);
and U18109 (N_18109,N_16990,N_14496);
nor U18110 (N_18110,N_12493,N_17703);
xnor U18111 (N_18111,N_13315,N_14831);
and U18112 (N_18112,N_12755,N_13712);
nand U18113 (N_18113,N_14838,N_13927);
nor U18114 (N_18114,N_13684,N_17183);
or U18115 (N_18115,N_16379,N_15287);
or U18116 (N_18116,N_17782,N_12290);
xnor U18117 (N_18117,N_16145,N_17317);
nor U18118 (N_18118,N_16218,N_12045);
nand U18119 (N_18119,N_17376,N_12834);
or U18120 (N_18120,N_17425,N_16797);
and U18121 (N_18121,N_17457,N_16984);
nand U18122 (N_18122,N_12618,N_15861);
or U18123 (N_18123,N_12883,N_14062);
and U18124 (N_18124,N_12435,N_13157);
nor U18125 (N_18125,N_17754,N_16862);
nand U18126 (N_18126,N_16800,N_14584);
and U18127 (N_18127,N_16788,N_13277);
and U18128 (N_18128,N_12379,N_17747);
or U18129 (N_18129,N_13040,N_16878);
and U18130 (N_18130,N_17897,N_17247);
xor U18131 (N_18131,N_12196,N_17010);
and U18132 (N_18132,N_17745,N_16895);
nand U18133 (N_18133,N_16968,N_15821);
xnor U18134 (N_18134,N_17369,N_14829);
nor U18135 (N_18135,N_12035,N_13319);
xor U18136 (N_18136,N_13551,N_13777);
nor U18137 (N_18137,N_14479,N_14355);
nor U18138 (N_18138,N_14944,N_12881);
and U18139 (N_18139,N_12532,N_15520);
xor U18140 (N_18140,N_15853,N_14816);
or U18141 (N_18141,N_13882,N_17445);
xnor U18142 (N_18142,N_13292,N_17174);
and U18143 (N_18143,N_14069,N_16902);
nor U18144 (N_18144,N_16488,N_14628);
nor U18145 (N_18145,N_15675,N_17102);
nor U18146 (N_18146,N_13138,N_14791);
nor U18147 (N_18147,N_13447,N_17854);
or U18148 (N_18148,N_14514,N_12773);
and U18149 (N_18149,N_13489,N_17329);
nand U18150 (N_18150,N_17451,N_16740);
nor U18151 (N_18151,N_14333,N_15538);
and U18152 (N_18152,N_15836,N_16231);
nor U18153 (N_18153,N_13955,N_12407);
xnor U18154 (N_18154,N_17070,N_17934);
xnor U18155 (N_18155,N_15141,N_13742);
or U18156 (N_18156,N_12895,N_15477);
nand U18157 (N_18157,N_16270,N_15841);
and U18158 (N_18158,N_14018,N_13210);
nand U18159 (N_18159,N_16780,N_16460);
nor U18160 (N_18160,N_12300,N_14214);
or U18161 (N_18161,N_15594,N_15939);
or U18162 (N_18162,N_12712,N_17073);
nand U18163 (N_18163,N_13480,N_12537);
or U18164 (N_18164,N_16418,N_14004);
and U18165 (N_18165,N_12221,N_16097);
or U18166 (N_18166,N_16492,N_15715);
xor U18167 (N_18167,N_13805,N_15845);
and U18168 (N_18168,N_15345,N_16642);
nor U18169 (N_18169,N_15318,N_16290);
nand U18170 (N_18170,N_15761,N_17395);
xor U18171 (N_18171,N_16126,N_14197);
nand U18172 (N_18172,N_17889,N_17863);
nand U18173 (N_18173,N_12898,N_12382);
or U18174 (N_18174,N_14712,N_14248);
xnor U18175 (N_18175,N_16803,N_13530);
or U18176 (N_18176,N_15512,N_14172);
and U18177 (N_18177,N_15769,N_16434);
nand U18178 (N_18178,N_12713,N_12648);
and U18179 (N_18179,N_16784,N_17135);
nor U18180 (N_18180,N_13180,N_14653);
or U18181 (N_18181,N_17920,N_14277);
nor U18182 (N_18182,N_13795,N_13442);
nor U18183 (N_18183,N_14076,N_17740);
and U18184 (N_18184,N_14338,N_13875);
or U18185 (N_18185,N_15211,N_13650);
nand U18186 (N_18186,N_13392,N_14695);
and U18187 (N_18187,N_17641,N_13071);
nand U18188 (N_18188,N_14233,N_17752);
nand U18189 (N_18189,N_17583,N_12687);
nor U18190 (N_18190,N_16828,N_14381);
nand U18191 (N_18191,N_16820,N_14786);
xnor U18192 (N_18192,N_14111,N_15820);
nor U18193 (N_18193,N_14567,N_12625);
and U18194 (N_18194,N_14771,N_16429);
and U18195 (N_18195,N_16092,N_15618);
nand U18196 (N_18196,N_14464,N_13596);
or U18197 (N_18197,N_15316,N_14268);
and U18198 (N_18198,N_13784,N_13379);
or U18199 (N_18199,N_13457,N_16472);
xnor U18200 (N_18200,N_13984,N_12542);
and U18201 (N_18201,N_12330,N_16844);
nor U18202 (N_18202,N_16545,N_13485);
and U18203 (N_18203,N_17773,N_15634);
nor U18204 (N_18204,N_14775,N_13852);
or U18205 (N_18205,N_17476,N_13359);
xor U18206 (N_18206,N_13592,N_17760);
nand U18207 (N_18207,N_16386,N_15868);
nor U18208 (N_18208,N_15256,N_13865);
nand U18209 (N_18209,N_14870,N_16432);
and U18210 (N_18210,N_12802,N_17699);
nand U18211 (N_18211,N_14843,N_12208);
nand U18212 (N_18212,N_12538,N_17492);
and U18213 (N_18213,N_13535,N_14369);
and U18214 (N_18214,N_17898,N_12993);
nor U18215 (N_18215,N_13806,N_15572);
xnor U18216 (N_18216,N_13076,N_12964);
and U18217 (N_18217,N_17684,N_16439);
nor U18218 (N_18218,N_12944,N_15478);
xor U18219 (N_18219,N_17439,N_14752);
and U18220 (N_18220,N_16914,N_14422);
or U18221 (N_18221,N_15353,N_14203);
or U18222 (N_18222,N_14038,N_12677);
and U18223 (N_18223,N_16321,N_14296);
or U18224 (N_18224,N_17482,N_15678);
and U18225 (N_18225,N_15689,N_12705);
or U18226 (N_18226,N_16411,N_14860);
and U18227 (N_18227,N_12507,N_12664);
and U18228 (N_18228,N_16363,N_15760);
xor U18229 (N_18229,N_12633,N_16573);
nand U18230 (N_18230,N_15314,N_12868);
and U18231 (N_18231,N_12962,N_16932);
nand U18232 (N_18232,N_16683,N_16723);
and U18233 (N_18233,N_14052,N_16536);
nand U18234 (N_18234,N_13781,N_17364);
xor U18235 (N_18235,N_13741,N_14147);
or U18236 (N_18236,N_15826,N_16738);
and U18237 (N_18237,N_15707,N_17363);
nand U18238 (N_18238,N_16591,N_16565);
nor U18239 (N_18239,N_14557,N_12541);
xnor U18240 (N_18240,N_14662,N_14886);
and U18241 (N_18241,N_14755,N_14702);
or U18242 (N_18242,N_15908,N_14300);
xnor U18243 (N_18243,N_14191,N_15215);
or U18244 (N_18244,N_13082,N_15986);
nand U18245 (N_18245,N_12771,N_13339);
or U18246 (N_18246,N_13060,N_17657);
or U18247 (N_18247,N_17503,N_17366);
nor U18248 (N_18248,N_15952,N_12871);
nor U18249 (N_18249,N_12332,N_14949);
or U18250 (N_18250,N_13380,N_15081);
nand U18251 (N_18251,N_16531,N_12955);
nand U18252 (N_18252,N_17527,N_12905);
xor U18253 (N_18253,N_14015,N_17749);
xnor U18254 (N_18254,N_13009,N_14284);
nor U18255 (N_18255,N_16002,N_16717);
xor U18256 (N_18256,N_13296,N_14358);
or U18257 (N_18257,N_15371,N_15968);
nor U18258 (N_18258,N_14166,N_14352);
and U18259 (N_18259,N_16426,N_15615);
xnor U18260 (N_18260,N_12127,N_13740);
xor U18261 (N_18261,N_17926,N_12082);
nor U18262 (N_18262,N_12470,N_14994);
and U18263 (N_18263,N_14719,N_13581);
xnor U18264 (N_18264,N_17812,N_12885);
or U18265 (N_18265,N_14064,N_12935);
xor U18266 (N_18266,N_15473,N_17980);
or U18267 (N_18267,N_13417,N_17690);
xor U18268 (N_18268,N_16739,N_13929);
nor U18269 (N_18269,N_14118,N_15164);
xor U18270 (N_18270,N_13998,N_14933);
or U18271 (N_18271,N_12823,N_15929);
nor U18272 (N_18272,N_17246,N_15007);
nand U18273 (N_18273,N_17322,N_17049);
nor U18274 (N_18274,N_14760,N_17596);
or U18275 (N_18275,N_16627,N_13027);
xor U18276 (N_18276,N_13900,N_15028);
nor U18277 (N_18277,N_15824,N_17730);
nand U18278 (N_18278,N_15451,N_13560);
and U18279 (N_18279,N_14100,N_14754);
nor U18280 (N_18280,N_17530,N_13878);
nor U18281 (N_18281,N_17082,N_16301);
nor U18282 (N_18282,N_12704,N_13252);
xnor U18283 (N_18283,N_16281,N_12981);
xor U18284 (N_18284,N_16632,N_12292);
nor U18285 (N_18285,N_17558,N_17098);
or U18286 (N_18286,N_16953,N_17396);
nand U18287 (N_18287,N_16572,N_12767);
nor U18288 (N_18288,N_15737,N_13765);
nand U18289 (N_18289,N_12187,N_17144);
nand U18290 (N_18290,N_17581,N_17241);
nand U18291 (N_18291,N_13819,N_14651);
nand U18292 (N_18292,N_14953,N_16725);
and U18293 (N_18293,N_12774,N_12293);
and U18294 (N_18294,N_14193,N_16149);
nand U18295 (N_18295,N_14202,N_17516);
nor U18296 (N_18296,N_13340,N_12462);
or U18297 (N_18297,N_12428,N_16450);
xnor U18298 (N_18298,N_14866,N_16088);
and U18299 (N_18299,N_16155,N_15203);
or U18300 (N_18300,N_15644,N_15811);
or U18301 (N_18301,N_17979,N_16000);
xnor U18302 (N_18302,N_16868,N_15698);
nand U18303 (N_18303,N_16234,N_14302);
or U18304 (N_18304,N_16403,N_16574);
nand U18305 (N_18305,N_16004,N_17836);
and U18306 (N_18306,N_12983,N_14920);
or U18307 (N_18307,N_15126,N_17348);
xnor U18308 (N_18308,N_15343,N_13258);
nor U18309 (N_18309,N_17556,N_12924);
xnor U18310 (N_18310,N_15568,N_12161);
nand U18311 (N_18311,N_12986,N_14414);
or U18312 (N_18312,N_16292,N_15515);
nor U18313 (N_18313,N_17041,N_14609);
and U18314 (N_18314,N_15109,N_13652);
xor U18315 (N_18315,N_15247,N_12138);
and U18316 (N_18316,N_15405,N_13764);
or U18317 (N_18317,N_12236,N_13993);
nand U18318 (N_18318,N_14152,N_17795);
or U18319 (N_18319,N_15921,N_12499);
nor U18320 (N_18320,N_15980,N_15503);
or U18321 (N_18321,N_16700,N_14859);
nor U18322 (N_18322,N_16167,N_13609);
or U18323 (N_18323,N_16793,N_14312);
or U18324 (N_18324,N_17303,N_14849);
nor U18325 (N_18325,N_13310,N_12272);
and U18326 (N_18326,N_15508,N_12423);
and U18327 (N_18327,N_17687,N_15711);
nand U18328 (N_18328,N_17882,N_13235);
nand U18329 (N_18329,N_14360,N_14747);
or U18330 (N_18330,N_17814,N_16356);
nor U18331 (N_18331,N_12162,N_12639);
nor U18332 (N_18332,N_13322,N_14098);
and U18333 (N_18333,N_14703,N_15115);
and U18334 (N_18334,N_12356,N_13568);
nand U18335 (N_18335,N_14385,N_16831);
or U18336 (N_18336,N_16698,N_14986);
and U18337 (N_18337,N_17874,N_13952);
and U18338 (N_18338,N_12882,N_15828);
nand U18339 (N_18339,N_13648,N_15570);
and U18340 (N_18340,N_12321,N_12970);
or U18341 (N_18341,N_14741,N_13317);
and U18342 (N_18342,N_15593,N_15245);
nor U18343 (N_18343,N_17628,N_14243);
xor U18344 (N_18344,N_15495,N_12666);
or U18345 (N_18345,N_16343,N_13896);
nand U18346 (N_18346,N_15143,N_15238);
nand U18347 (N_18347,N_15057,N_13038);
nand U18348 (N_18348,N_15036,N_15017);
or U18349 (N_18349,N_15940,N_17319);
and U18350 (N_18350,N_16731,N_15680);
nor U18351 (N_18351,N_16091,N_17158);
and U18352 (N_18352,N_16703,N_12146);
or U18353 (N_18353,N_14725,N_12027);
nand U18354 (N_18354,N_13483,N_13088);
nor U18355 (N_18355,N_14547,N_13624);
and U18356 (N_18356,N_17604,N_14704);
or U18357 (N_18357,N_17326,N_15053);
nor U18358 (N_18358,N_14581,N_12546);
xor U18359 (N_18359,N_17759,N_15799);
nor U18360 (N_18360,N_17486,N_16307);
or U18361 (N_18361,N_14823,N_12794);
nor U18362 (N_18362,N_13833,N_14819);
nand U18363 (N_18363,N_16063,N_13276);
or U18364 (N_18364,N_15282,N_12131);
nor U18365 (N_18365,N_13314,N_13163);
nand U18366 (N_18366,N_15964,N_13055);
nand U18367 (N_18367,N_16111,N_16613);
nor U18368 (N_18368,N_13406,N_17567);
nand U18369 (N_18369,N_13649,N_16971);
and U18370 (N_18370,N_12500,N_15562);
nor U18371 (N_18371,N_13179,N_13323);
xnor U18372 (N_18372,N_17872,N_15363);
nor U18373 (N_18373,N_12183,N_17998);
xor U18374 (N_18374,N_13982,N_15509);
and U18375 (N_18375,N_12925,N_16874);
xnor U18376 (N_18376,N_14097,N_14445);
nand U18377 (N_18377,N_14117,N_12787);
and U18378 (N_18378,N_15887,N_14865);
and U18379 (N_18379,N_13901,N_17973);
nand U18380 (N_18380,N_13037,N_14813);
and U18381 (N_18381,N_15924,N_14067);
and U18382 (N_18382,N_15795,N_15628);
and U18383 (N_18383,N_17588,N_17499);
xnor U18384 (N_18384,N_15416,N_13183);
xor U18385 (N_18385,N_17169,N_17912);
nor U18386 (N_18386,N_17565,N_17231);
and U18387 (N_18387,N_12012,N_14826);
or U18388 (N_18388,N_15575,N_12482);
nand U18389 (N_18389,N_12912,N_13284);
nand U18390 (N_18390,N_16332,N_12296);
and U18391 (N_18391,N_13119,N_17661);
or U18392 (N_18392,N_12852,N_12847);
or U18393 (N_18393,N_15151,N_14634);
or U18394 (N_18394,N_14985,N_17332);
nor U18395 (N_18395,N_17810,N_12875);
or U18396 (N_18396,N_17716,N_13390);
nand U18397 (N_18397,N_14131,N_14690);
xnor U18398 (N_18398,N_17625,N_12433);
nor U18399 (N_18399,N_16714,N_15901);
and U18400 (N_18400,N_14241,N_16237);
nor U18401 (N_18401,N_16728,N_12768);
nor U18402 (N_18402,N_13543,N_16983);
nand U18403 (N_18403,N_12571,N_17895);
or U18404 (N_18404,N_17523,N_14808);
xnor U18405 (N_18405,N_17184,N_16327);
nor U18406 (N_18406,N_14071,N_17693);
and U18407 (N_18407,N_17368,N_17847);
nand U18408 (N_18408,N_17916,N_14145);
xnor U18409 (N_18409,N_15663,N_16677);
or U18410 (N_18410,N_14575,N_15055);
or U18411 (N_18411,N_17127,N_17869);
nand U18412 (N_18412,N_16481,N_14649);
xnor U18413 (N_18413,N_14850,N_16796);
nor U18414 (N_18414,N_13526,N_17611);
xnor U18415 (N_18415,N_17340,N_12217);
xnor U18416 (N_18416,N_15919,N_16799);
nor U18417 (N_18417,N_12281,N_13482);
or U18418 (N_18418,N_12475,N_12988);
nor U18419 (N_18419,N_15588,N_15277);
or U18420 (N_18420,N_14615,N_17913);
nand U18421 (N_18421,N_17034,N_17248);
nand U18422 (N_18422,N_15886,N_16832);
or U18423 (N_18423,N_13433,N_15903);
and U18424 (N_18424,N_17660,N_17351);
xor U18425 (N_18425,N_17281,N_16020);
nand U18426 (N_18426,N_16143,N_12204);
nand U18427 (N_18427,N_15105,N_13289);
xor U18428 (N_18428,N_14750,N_12449);
nor U18429 (N_18429,N_17411,N_15873);
and U18430 (N_18430,N_14637,N_12312);
nand U18431 (N_18431,N_16751,N_14620);
nand U18432 (N_18432,N_15673,N_17809);
or U18433 (N_18433,N_16277,N_13963);
nand U18434 (N_18434,N_12730,N_12368);
nand U18435 (N_18435,N_12497,N_15557);
nand U18436 (N_18436,N_12809,N_13225);
or U18437 (N_18437,N_16904,N_16124);
xnor U18438 (N_18438,N_16634,N_17494);
or U18439 (N_18439,N_16477,N_12756);
and U18440 (N_18440,N_12394,N_13894);
nand U18441 (N_18441,N_16207,N_17261);
xor U18442 (N_18442,N_16909,N_12927);
xor U18443 (N_18443,N_17334,N_16388);
nand U18444 (N_18444,N_12319,N_15746);
nand U18445 (N_18445,N_17459,N_17388);
nand U18446 (N_18446,N_15082,N_16065);
nand U18447 (N_18447,N_17584,N_12398);
nand U18448 (N_18448,N_14077,N_15208);
nor U18449 (N_18449,N_13961,N_13367);
or U18450 (N_18450,N_13723,N_17839);
nor U18451 (N_18451,N_13773,N_13355);
or U18452 (N_18452,N_14028,N_14665);
nor U18453 (N_18453,N_16414,N_13763);
xor U18454 (N_18454,N_12651,N_15241);
nand U18455 (N_18455,N_16835,N_17471);
nand U18456 (N_18456,N_16724,N_12128);
and U18457 (N_18457,N_17914,N_12489);
nand U18458 (N_18458,N_16678,N_17591);
nand U18459 (N_18459,N_16105,N_12377);
and U18460 (N_18460,N_16034,N_14317);
nand U18461 (N_18461,N_12317,N_14462);
and U18462 (N_18462,N_16760,N_12991);
or U18463 (N_18463,N_15442,N_14321);
and U18464 (N_18464,N_15487,N_12088);
xor U18465 (N_18465,N_15590,N_15573);
xor U18466 (N_18466,N_15201,N_16732);
nand U18467 (N_18467,N_14632,N_15857);
nand U18468 (N_18468,N_17894,N_17013);
nand U18469 (N_18469,N_15564,N_12120);
and U18470 (N_18470,N_12785,N_12355);
nor U18471 (N_18471,N_15870,N_12008);
nor U18472 (N_18472,N_12222,N_17502);
xnor U18473 (N_18473,N_16541,N_17978);
nand U18474 (N_18474,N_16858,N_16402);
nor U18475 (N_18475,N_12455,N_12833);
nor U18476 (N_18476,N_12568,N_17549);
or U18477 (N_18477,N_12308,N_15200);
nand U18478 (N_18478,N_16812,N_16036);
xor U18479 (N_18479,N_16537,N_17715);
and U18480 (N_18480,N_13395,N_16368);
xor U18481 (N_18481,N_15989,N_15790);
or U18482 (N_18482,N_14574,N_12157);
xnor U18483 (N_18483,N_15336,N_16412);
nor U18484 (N_18484,N_15350,N_12911);
or U18485 (N_18485,N_17418,N_16947);
or U18486 (N_18486,N_16033,N_15781);
nand U18487 (N_18487,N_14066,N_17120);
or U18488 (N_18488,N_13979,N_12697);
and U18489 (N_18489,N_15535,N_13746);
nand U18490 (N_18490,N_13548,N_13272);
or U18491 (N_18491,N_14415,N_17548);
nor U18492 (N_18492,N_17290,N_13011);
nand U18493 (N_18493,N_14187,N_13724);
xnor U18494 (N_18494,N_12728,N_16066);
or U18495 (N_18495,N_14938,N_17091);
nor U18496 (N_18496,N_12555,N_13815);
or U18497 (N_18497,N_13470,N_16031);
xor U18498 (N_18498,N_14982,N_13504);
nand U18499 (N_18499,N_14979,N_16093);
and U18500 (N_18500,N_13690,N_16667);
or U18501 (N_18501,N_14151,N_13848);
nor U18502 (N_18502,N_14042,N_16830);
or U18503 (N_18503,N_15054,N_12936);
nand U18504 (N_18504,N_14045,N_16208);
xnor U18505 (N_18505,N_13691,N_16801);
nand U18506 (N_18506,N_15484,N_14995);
and U18507 (N_18507,N_16736,N_12751);
nor U18508 (N_18508,N_14877,N_12411);
and U18509 (N_18509,N_15884,N_15169);
and U18510 (N_18510,N_16229,N_17540);
and U18511 (N_18511,N_12715,N_15462);
and U18512 (N_18512,N_17104,N_13992);
nand U18513 (N_18513,N_14494,N_17791);
xnor U18514 (N_18514,N_12866,N_15695);
nand U18515 (N_18515,N_15452,N_16982);
or U18516 (N_18516,N_14326,N_13135);
and U18517 (N_18517,N_12416,N_13597);
nor U18518 (N_18518,N_13556,N_17036);
xor U18519 (N_18519,N_14387,N_17383);
or U18520 (N_18520,N_13944,N_14240);
and U18521 (N_18521,N_16783,N_12469);
and U18522 (N_18522,N_14955,N_13399);
nand U18523 (N_18523,N_17313,N_12451);
nor U18524 (N_18524,N_15138,N_12897);
nand U18525 (N_18525,N_15339,N_17559);
xor U18526 (N_18526,N_15972,N_17896);
xor U18527 (N_18527,N_13144,N_15875);
and U18528 (N_18528,N_12680,N_14590);
or U18529 (N_18529,N_13219,N_13410);
xnor U18530 (N_18530,N_14086,N_13580);
or U18531 (N_18531,N_16822,N_12425);
xnor U18532 (N_18532,N_14114,N_14664);
nand U18533 (N_18533,N_14684,N_15087);
and U18534 (N_18534,N_12409,N_13676);
or U18535 (N_18535,N_14308,N_14323);
nand U18536 (N_18536,N_17713,N_15645);
nor U18537 (N_18537,N_16258,N_13174);
nand U18538 (N_18538,N_17831,N_13801);
or U18539 (N_18539,N_13342,N_13689);
or U18540 (N_18540,N_13782,N_12361);
nand U18541 (N_18541,N_13559,N_12707);
and U18542 (N_18542,N_16006,N_14297);
xnor U18543 (N_18543,N_13344,N_14359);
and U18544 (N_18544,N_13814,N_16104);
xnor U18545 (N_18545,N_13389,N_17574);
nor U18546 (N_18546,N_15946,N_16315);
nor U18547 (N_18547,N_17473,N_16657);
nor U18548 (N_18548,N_16913,N_13373);
nand U18549 (N_18549,N_15450,N_15822);
and U18550 (N_18550,N_16364,N_16713);
xnor U18551 (N_18551,N_17085,N_16295);
and U18552 (N_18552,N_12069,N_12933);
xor U18553 (N_18553,N_16053,N_13021);
or U18554 (N_18554,N_15531,N_13287);
nand U18555 (N_18555,N_13320,N_16252);
nand U18556 (N_18556,N_16915,N_12478);
nor U18557 (N_18557,N_14576,N_14545);
xnor U18558 (N_18558,N_14606,N_15390);
or U18559 (N_18559,N_12066,N_14427);
or U18560 (N_18560,N_12793,N_14503);
or U18561 (N_18561,N_16544,N_15040);
or U18562 (N_18562,N_16744,N_14970);
nor U18563 (N_18563,N_16061,N_15440);
nor U18564 (N_18564,N_14453,N_12932);
nor U18565 (N_18565,N_14560,N_13738);
nor U18566 (N_18566,N_12173,N_15794);
nand U18567 (N_18567,N_17707,N_13419);
or U18568 (N_18568,N_16090,N_13725);
nor U18569 (N_18569,N_16578,N_15444);
and U18570 (N_18570,N_17479,N_12005);
or U18571 (N_18571,N_15768,N_14729);
xnor U18572 (N_18572,N_12930,N_15724);
or U18573 (N_18573,N_13012,N_12874);
or U18574 (N_18574,N_17629,N_13623);
nand U18575 (N_18575,N_13945,N_16519);
and U18576 (N_18576,N_16493,N_12752);
xor U18577 (N_18577,N_15307,N_14799);
nand U18578 (N_18578,N_15183,N_13431);
xor U18579 (N_18579,N_17834,N_17564);
xnor U18580 (N_18580,N_16349,N_17710);
and U18581 (N_18581,N_15376,N_17284);
and U18582 (N_18582,N_16370,N_12657);
xor U18583 (N_18583,N_13972,N_17933);
xnor U18584 (N_18584,N_15166,N_15199);
nand U18585 (N_18585,N_16702,N_13108);
nand U18586 (N_18586,N_12907,N_12892);
nor U18587 (N_18587,N_12013,N_12363);
xnor U18588 (N_18588,N_16504,N_16203);
nand U18589 (N_18589,N_13377,N_14599);
nand U18590 (N_18590,N_15602,N_16758);
xor U18591 (N_18591,N_13280,N_16176);
nand U18592 (N_18592,N_15013,N_14341);
and U18593 (N_18593,N_12769,N_16567);
and U18594 (N_18594,N_16142,N_15536);
or U18595 (N_18595,N_13813,N_17904);
nand U18596 (N_18596,N_12872,N_13885);
nor U18597 (N_18597,N_13278,N_14679);
nand U18598 (N_18598,N_13593,N_13270);
xnor U18599 (N_18599,N_13321,N_13804);
or U18600 (N_18600,N_16141,N_14987);
nor U18601 (N_18601,N_17006,N_15490);
or U18602 (N_18602,N_14789,N_12609);
and U18603 (N_18603,N_16864,N_14181);
or U18604 (N_18604,N_17531,N_17667);
nand U18605 (N_18605,N_13637,N_12679);
nand U18606 (N_18606,N_13710,N_12086);
nor U18607 (N_18607,N_12077,N_14171);
nand U18608 (N_18608,N_15597,N_15691);
xor U18609 (N_18609,N_14978,N_17288);
or U18610 (N_18610,N_14716,N_15851);
xnor U18611 (N_18611,N_13575,N_15889);
nand U18612 (N_18612,N_12512,N_13295);
xor U18613 (N_18613,N_16287,N_13578);
xor U18614 (N_18614,N_14686,N_13981);
nor U18615 (N_18615,N_13312,N_13673);
or U18616 (N_18616,N_14773,N_16856);
xor U18617 (N_18617,N_17300,N_14509);
or U18618 (N_18618,N_13198,N_17063);
and U18619 (N_18619,N_16267,N_17024);
nor U18620 (N_18620,N_17019,N_13120);
and U18621 (N_18621,N_16309,N_17433);
or U18622 (N_18622,N_12185,N_12498);
and U18623 (N_18623,N_12861,N_16499);
nand U18624 (N_18624,N_13035,N_15823);
and U18625 (N_18625,N_13975,N_17390);
xnor U18626 (N_18626,N_16458,N_17047);
and U18627 (N_18627,N_17195,N_14582);
and U18628 (N_18628,N_14431,N_12089);
or U18629 (N_18629,N_15481,N_15793);
xnor U18630 (N_18630,N_13382,N_15159);
xor U18631 (N_18631,N_15688,N_14794);
xnor U18632 (N_18632,N_17743,N_15402);
and U18633 (N_18633,N_13909,N_13487);
nand U18634 (N_18634,N_16581,N_14861);
nand U18635 (N_18635,N_14573,N_15954);
nor U18636 (N_18636,N_13366,N_13524);
nand U18637 (N_18637,N_17201,N_17407);
nand U18638 (N_18638,N_17617,N_15906);
or U18639 (N_18639,N_17078,N_15471);
and U18640 (N_18640,N_14513,N_16666);
nand U18641 (N_18641,N_13547,N_17446);
nand U18642 (N_18642,N_14037,N_16680);
nor U18643 (N_18643,N_12543,N_16688);
and U18644 (N_18644,N_16837,N_16456);
nor U18645 (N_18645,N_14502,N_12223);
xnor U18646 (N_18646,N_13588,N_12514);
nand U18647 (N_18647,N_14329,N_17188);
xnor U18648 (N_18648,N_12155,N_17415);
nand U18649 (N_18649,N_12610,N_12890);
and U18650 (N_18650,N_16707,N_15843);
and U18651 (N_18651,N_13861,N_12408);
nand U18652 (N_18652,N_12265,N_16210);
nor U18653 (N_18653,N_17995,N_13767);
nand U18654 (N_18654,N_17696,N_12814);
or U18655 (N_18655,N_15780,N_16465);
nand U18656 (N_18656,N_14734,N_15430);
or U18657 (N_18657,N_14597,N_12143);
xor U18658 (N_18658,N_13639,N_14600);
nand U18659 (N_18659,N_14085,N_13350);
and U18660 (N_18660,N_17297,N_14883);
and U18661 (N_18661,N_12782,N_15324);
or U18662 (N_18662,N_12519,N_12176);
or U18663 (N_18663,N_16079,N_15300);
nor U18664 (N_18664,N_12711,N_17084);
nand U18665 (N_18665,N_17107,N_17802);
nand U18666 (N_18666,N_17219,N_12153);
xor U18667 (N_18667,N_12804,N_13351);
nor U18668 (N_18668,N_15008,N_16869);
or U18669 (N_18669,N_12386,N_17491);
xor U18670 (N_18670,N_16255,N_16086);
xnor U18671 (N_18671,N_14926,N_14090);
xnor U18672 (N_18672,N_12968,N_12040);
nor U18673 (N_18673,N_13698,N_17211);
and U18674 (N_18674,N_12853,N_17113);
and U18675 (N_18675,N_13988,N_17352);
nand U18676 (N_18676,N_14180,N_17037);
nor U18677 (N_18677,N_14265,N_12850);
xnor U18678 (N_18678,N_14340,N_17200);
nand U18679 (N_18679,N_16484,N_17515);
xor U18680 (N_18680,N_17148,N_12345);
or U18681 (N_18681,N_15984,N_12401);
xor U18682 (N_18682,N_12240,N_13147);
and U18683 (N_18683,N_14570,N_12765);
and U18684 (N_18684,N_16197,N_16767);
or U18685 (N_18685,N_15107,N_14095);
and U18686 (N_18686,N_13491,N_16926);
nand U18687 (N_18687,N_17321,N_17997);
and U18688 (N_18688,N_17631,N_16785);
nor U18689 (N_18689,N_12797,N_16289);
nand U18690 (N_18690,N_14824,N_12336);
or U18691 (N_18691,N_12828,N_14210);
nand U18692 (N_18692,N_15206,N_14121);
and U18693 (N_18693,N_17197,N_15482);
nor U18694 (N_18694,N_17555,N_16892);
or U18695 (N_18695,N_13678,N_16873);
xor U18696 (N_18696,N_14517,N_16601);
nor U18697 (N_18697,N_15587,N_12766);
xnor U18698 (N_18698,N_15391,N_16540);
nor U18699 (N_18699,N_17996,N_14383);
nand U18700 (N_18700,N_17140,N_16489);
xor U18701 (N_18701,N_12028,N_13434);
and U18702 (N_18702,N_14019,N_16181);
or U18703 (N_18703,N_15401,N_13338);
nand U18704 (N_18704,N_14178,N_12582);
and U18705 (N_18705,N_17057,N_14012);
nor U18706 (N_18706,N_17826,N_13872);
nor U18707 (N_18707,N_17589,N_15519);
or U18708 (N_18708,N_15264,N_13950);
or U18709 (N_18709,N_14314,N_14208);
xor U18710 (N_18710,N_14299,N_12006);
nand U18711 (N_18711,N_15776,N_14235);
xor U18712 (N_18712,N_17016,N_13020);
nor U18713 (N_18713,N_15739,N_16094);
or U18714 (N_18714,N_17963,N_15294);
or U18715 (N_18715,N_15829,N_13205);
nor U18716 (N_18716,N_15825,N_14109);
nor U18717 (N_18717,N_12387,N_16733);
nor U18718 (N_18718,N_14138,N_13685);
or U18719 (N_18719,N_15457,N_16900);
or U18720 (N_18720,N_12205,N_12763);
and U18721 (N_18721,N_13250,N_13472);
xnor U18722 (N_18722,N_15049,N_15226);
nor U18723 (N_18723,N_15816,N_16923);
xor U18724 (N_18724,N_13863,N_15753);
and U18725 (N_18725,N_12214,N_12603);
nand U18726 (N_18726,N_12316,N_14050);
nor U18727 (N_18727,N_12928,N_12010);
or U18728 (N_18728,N_16271,N_12926);
or U18729 (N_18729,N_13445,N_17232);
nor U18730 (N_18730,N_17893,N_14175);
or U18731 (N_18731,N_14136,N_17903);
nor U18732 (N_18732,N_13938,N_16549);
and U18733 (N_18733,N_14693,N_17346);
or U18734 (N_18734,N_14225,N_13743);
nor U18735 (N_18735,N_15607,N_13915);
and U18736 (N_18736,N_15272,N_15566);
or U18737 (N_18737,N_14984,N_16146);
nand U18738 (N_18738,N_17551,N_14677);
nand U18739 (N_18739,N_15777,N_13564);
or U18740 (N_18740,N_17023,N_15110);
and U18741 (N_18741,N_13333,N_16221);
nor U18742 (N_18742,N_17849,N_15348);
and U18743 (N_18743,N_16942,N_14515);
and U18744 (N_18744,N_16058,N_12643);
and U18745 (N_18745,N_15408,N_12829);
or U18746 (N_18746,N_14743,N_16030);
xnor U18747 (N_18747,N_14643,N_17977);
nor U18748 (N_18748,N_12661,N_16169);
or U18749 (N_18749,N_15718,N_15063);
and U18750 (N_18750,N_17137,N_17386);
nand U18751 (N_18751,N_12843,N_13444);
xor U18752 (N_18752,N_17698,N_16845);
xor U18753 (N_18753,N_16278,N_17477);
and U18754 (N_18754,N_14740,N_12702);
and U18755 (N_18755,N_16390,N_14364);
nor U18756 (N_18756,N_16116,N_14007);
or U18757 (N_18757,N_14602,N_15386);
nand U18758 (N_18758,N_14527,N_17289);
xor U18759 (N_18759,N_16161,N_12243);
nor U18760 (N_18760,N_16202,N_15445);
nand U18761 (N_18761,N_17355,N_16437);
or U18762 (N_18762,N_13329,N_17301);
and U18763 (N_18763,N_16377,N_14564);
or U18764 (N_18764,N_14652,N_12781);
or U18765 (N_18765,N_15920,N_12899);
and U18766 (N_18766,N_17115,N_14480);
and U18767 (N_18767,N_14989,N_15709);
nor U18768 (N_18768,N_16125,N_16509);
xnor U18769 (N_18769,N_13110,N_14875);
and U18770 (N_18770,N_17438,N_13577);
nand U18771 (N_18771,N_12139,N_16109);
xnor U18772 (N_18772,N_12599,N_12257);
nor U18773 (N_18773,N_17649,N_12586);
or U18774 (N_18774,N_17714,N_12307);
and U18775 (N_18775,N_15099,N_14939);
nor U18776 (N_18776,N_13134,N_15849);
and U18777 (N_18777,N_13095,N_16839);
and U18778 (N_18778,N_15532,N_15158);
nand U18779 (N_18779,N_14872,N_16206);
xor U18780 (N_18780,N_17264,N_17108);
xor U18781 (N_18781,N_16639,N_15418);
or U18782 (N_18782,N_15658,N_16877);
nand U18783 (N_18783,N_14937,N_17338);
nand U18784 (N_18784,N_16967,N_14688);
xnor U18785 (N_18785,N_12468,N_15204);
and U18786 (N_18786,N_14908,N_17522);
and U18787 (N_18787,N_16298,N_13595);
nand U18788 (N_18788,N_12951,N_17900);
nand U18789 (N_18789,N_12987,N_17506);
and U18790 (N_18790,N_13150,N_13331);
nor U18791 (N_18791,N_14887,N_16344);
nand U18792 (N_18792,N_12004,N_13747);
xor U18793 (N_18793,N_17315,N_17089);
xor U18794 (N_18794,N_12662,N_12057);
or U18795 (N_18795,N_13481,N_15486);
nor U18796 (N_18796,N_17462,N_12150);
and U18797 (N_18797,N_16296,N_14676);
xnor U18798 (N_18798,N_16048,N_15589);
xor U18799 (N_18799,N_12887,N_16697);
xor U18800 (N_18800,N_13864,N_15543);
and U18801 (N_18801,N_14334,N_14348);
xor U18802 (N_18802,N_15608,N_17621);
nand U18803 (N_18803,N_15446,N_16122);
and U18804 (N_18804,N_15084,N_13004);
xnor U18805 (N_18805,N_17941,N_17970);
or U18806 (N_18806,N_17450,N_17676);
or U18807 (N_18807,N_15725,N_12671);
nand U18808 (N_18808,N_17460,N_15356);
nand U18809 (N_18809,N_15510,N_17058);
and U18810 (N_18810,N_12686,N_14660);
nor U18811 (N_18811,N_12339,N_12445);
and U18812 (N_18812,N_13663,N_16095);
or U18813 (N_18813,N_15411,N_12952);
and U18814 (N_18814,N_17888,N_12101);
and U18815 (N_18815,N_12518,N_13511);
xnor U18816 (N_18816,N_14439,N_13299);
nor U18817 (N_18817,N_14552,N_14647);
xnor U18818 (N_18818,N_14542,N_16763);
or U18819 (N_18819,N_12524,N_15627);
and U18820 (N_18820,N_16380,N_17608);
and U18821 (N_18821,N_13500,N_13512);
nand U18822 (N_18822,N_13221,N_13274);
nand U18823 (N_18823,N_16951,N_15775);
nor U18824 (N_18824,N_16433,N_17216);
or U18825 (N_18825,N_14914,N_12526);
xnor U18826 (N_18826,N_13086,N_14732);
xor U18827 (N_18827,N_15896,N_14433);
xor U18828 (N_18828,N_12140,N_16378);
nor U18829 (N_18829,N_14833,N_13523);
nand U18830 (N_18830,N_17767,N_13257);
xor U18831 (N_18831,N_16715,N_16908);
nor U18832 (N_18832,N_15872,N_12020);
or U18833 (N_18833,N_15497,N_12179);
xnor U18834 (N_18834,N_17259,N_14529);
nor U18835 (N_18835,N_14778,N_16888);
or U18836 (N_18836,N_14405,N_14965);
or U18837 (N_18837,N_16135,N_13772);
xor U18838 (N_18838,N_16661,N_12288);
xor U18839 (N_18839,N_16085,N_16186);
xor U18840 (N_18840,N_14701,N_16557);
or U18841 (N_18841,N_15419,N_16013);
nand U18842 (N_18842,N_15156,N_16384);
nor U18843 (N_18843,N_17335,N_17312);
nand U18844 (N_18844,N_13572,N_17076);
nand U18845 (N_18845,N_13249,N_12698);
nand U18846 (N_18846,N_15502,N_14423);
nor U18847 (N_18847,N_16497,N_13488);
xor U18848 (N_18848,N_16043,N_15132);
xnor U18849 (N_18849,N_16986,N_13655);
or U18850 (N_18850,N_13707,N_17722);
nor U18851 (N_18851,N_17570,N_17419);
xnor U18852 (N_18852,N_16483,N_13152);
nand U18853 (N_18853,N_13545,N_15180);
or U18854 (N_18854,N_13942,N_17337);
xnor U18855 (N_18855,N_13974,N_17665);
nand U18856 (N_18856,N_16165,N_14869);
and U18857 (N_18857,N_16664,N_12733);
xor U18858 (N_18858,N_13749,N_17274);
xnor U18859 (N_18859,N_14579,N_15097);
nor U18860 (N_18860,N_14471,N_14337);
and U18861 (N_18861,N_17844,N_12720);
nor U18862 (N_18862,N_17170,N_13450);
nor U18863 (N_18863,N_16849,N_16096);
nand U18864 (N_18864,N_17815,N_14492);
xnor U18865 (N_18865,N_16051,N_12965);
and U18866 (N_18866,N_14781,N_12830);
or U18867 (N_18867,N_12579,N_13549);
or U18868 (N_18868,N_17787,N_14543);
nand U18869 (N_18869,N_17275,N_13248);
xnor U18870 (N_18870,N_17985,N_16653);
nor U18871 (N_18871,N_14685,N_16663);
or U18872 (N_18872,N_14497,N_15424);
and U18873 (N_18873,N_15525,N_15186);
nor U18874 (N_18874,N_16745,N_13256);
nand U18875 (N_18875,N_14105,N_13834);
or U18876 (N_18876,N_17656,N_17133);
nand U18877 (N_18877,N_14650,N_16624);
and U18878 (N_18878,N_13584,N_13922);
nand U18879 (N_18879,N_15346,N_13059);
xor U18880 (N_18880,N_17397,N_14476);
nand U18881 (N_18881,N_17938,N_16994);
xor U18882 (N_18882,N_17606,N_14370);
nor U18883 (N_18883,N_17751,N_16246);
or U18884 (N_18884,N_15630,N_12050);
xor U18885 (N_18885,N_12121,N_13303);
and U18886 (N_18886,N_16046,N_15223);
and U18887 (N_18887,N_15959,N_14252);
nand U18888 (N_18888,N_17712,N_15071);
nand U18889 (N_18889,N_17389,N_14925);
nand U18890 (N_18890,N_12761,N_12835);
nand U18891 (N_18891,N_14762,N_12167);
nor U18892 (N_18892,N_13181,N_15224);
nor U18893 (N_18893,N_14093,N_16297);
nand U18894 (N_18894,N_14837,N_17474);
and U18895 (N_18895,N_17484,N_16580);
or U18896 (N_18896,N_13072,N_15696);
and U18897 (N_18897,N_12522,N_13067);
xnor U18898 (N_18898,N_13149,N_15740);
nand U18899 (N_18899,N_15342,N_17238);
xor U18900 (N_18900,N_12919,N_14853);
and U18901 (N_18901,N_14350,N_12716);
nand U18902 (N_18902,N_14974,N_17097);
xnor U18903 (N_18903,N_15325,N_14963);
or U18904 (N_18904,N_15734,N_14640);
nand U18905 (N_18905,N_17449,N_13361);
nand U18906 (N_18906,N_15913,N_16952);
xor U18907 (N_18907,N_13953,N_16534);
xnor U18908 (N_18908,N_15417,N_15434);
and U18909 (N_18909,N_14940,N_17925);
and U18910 (N_18910,N_15530,N_13372);
or U18911 (N_18911,N_12701,N_14950);
nor U18912 (N_18912,N_14551,N_17221);
nor U18913 (N_18913,N_14541,N_13025);
nand U18914 (N_18914,N_15683,N_17318);
nand U18915 (N_18915,N_13396,N_14531);
nor U18916 (N_18916,N_13398,N_17513);
and U18917 (N_18917,N_13162,N_13094);
or U18918 (N_18918,N_15291,N_15882);
and U18919 (N_18919,N_12811,N_12488);
nand U18920 (N_18920,N_16177,N_12311);
xor U18921 (N_18921,N_12920,N_16670);
nand U18922 (N_18922,N_17966,N_17504);
nand U18923 (N_18923,N_12737,N_15548);
or U18924 (N_18924,N_13744,N_14418);
and U18925 (N_18925,N_12684,N_12800);
and U18926 (N_18926,N_14412,N_17465);
nand U18927 (N_18927,N_15897,N_13496);
and U18928 (N_18928,N_16134,N_17820);
or U18929 (N_18929,N_13204,N_12958);
nor U18930 (N_18930,N_13672,N_13214);
or U18931 (N_18931,N_17420,N_17495);
nor U18932 (N_18932,N_14231,N_12977);
nor U18933 (N_18933,N_14033,N_13991);
or U18934 (N_18934,N_15528,N_15865);
and U18935 (N_18935,N_12277,N_14103);
or U18936 (N_18936,N_16284,N_14182);
or U18937 (N_18937,N_12123,N_17829);
or U18938 (N_18938,N_12674,N_12181);
nand U18939 (N_18939,N_16422,N_13711);
nand U18940 (N_18940,N_12061,N_12271);
nand U18941 (N_18941,N_12495,N_15061);
and U18942 (N_18942,N_13155,N_14537);
nor U18943 (N_18943,N_16113,N_14782);
xnor U18944 (N_18944,N_13130,N_13873);
nand U18945 (N_18945,N_12058,N_16428);
xor U18946 (N_18946,N_13202,N_16988);
nor U18947 (N_18947,N_15207,N_16253);
nor U18948 (N_18948,N_16768,N_14089);
or U18949 (N_18949,N_15425,N_14400);
and U18950 (N_18950,N_14472,N_13462);
xor U18951 (N_18951,N_15142,N_13478);
nand U18952 (N_18952,N_14244,N_15614);
xnor U18953 (N_18953,N_12275,N_15240);
or U18954 (N_18954,N_16310,N_12904);
xnor U18955 (N_18955,N_15842,N_15951);
nand U18956 (N_18956,N_15910,N_13520);
nor U18957 (N_18957,N_15957,N_14889);
xnor U18958 (N_18958,N_14099,N_13057);
xnor U18959 (N_18959,N_13416,N_15782);
and U18960 (N_18960,N_13803,N_13704);
and U18961 (N_18961,N_14604,N_13527);
or U18962 (N_18962,N_16503,N_17422);
xor U18963 (N_18963,N_12612,N_17921);
nor U18964 (N_18964,N_13237,N_17612);
or U18965 (N_18965,N_13065,N_15580);
or U18966 (N_18966,N_14571,N_12552);
nand U18967 (N_18967,N_12735,N_12535);
or U18968 (N_18968,N_13786,N_15830);
nand U18969 (N_18969,N_17788,N_14905);
or U18970 (N_18970,N_13586,N_17121);
nand U18971 (N_18971,N_16782,N_15869);
nor U18972 (N_18972,N_13064,N_16747);
nor U18973 (N_18973,N_13384,N_17145);
nor U18974 (N_18974,N_13041,N_15041);
nor U18975 (N_18975,N_13695,N_13172);
nand U18976 (N_18976,N_14211,N_13855);
or U18977 (N_18977,N_17072,N_12026);
or U18978 (N_18978,N_13118,N_15895);
or U18979 (N_18979,N_16937,N_16220);
or U18980 (N_18980,N_13737,N_15757);
nand U18981 (N_18981,N_14113,N_17043);
nor U18982 (N_18982,N_16676,N_16486);
xnor U18983 (N_18983,N_12553,N_13928);
xnor U18984 (N_18984,N_14409,N_13877);
nor U18985 (N_18985,N_17028,N_15121);
xnor U18986 (N_18986,N_16502,N_12018);
and U18987 (N_18987,N_12349,N_15426);
xnor U18988 (N_18988,N_15571,N_15834);
xor U18989 (N_18989,N_15218,N_14764);
or U18990 (N_18990,N_17639,N_17790);
nor U18991 (N_18991,N_14026,N_13843);
xnor U18992 (N_18992,N_14058,N_16522);
or U18993 (N_18993,N_16811,N_17164);
or U18994 (N_18994,N_15978,N_12778);
and U18995 (N_18995,N_14342,N_12341);
nand U18996 (N_18996,N_12194,N_16174);
nand U18997 (N_18997,N_16352,N_17601);
xnor U18998 (N_18998,N_17528,N_14406);
xor U18999 (N_18999,N_14283,N_16692);
nor U19000 (N_19000,N_16335,N_13264);
and U19001 (N_19001,N_14104,N_17736);
nor U19002 (N_19002,N_14967,N_17737);
or U19003 (N_19003,N_14927,N_16025);
nor U19004 (N_19004,N_13084,N_14389);
and U19005 (N_19005,N_17413,N_14236);
and U19006 (N_19006,N_16425,N_15948);
nor U19007 (N_19007,N_13890,N_13383);
or U19008 (N_19008,N_15463,N_15060);
or U19009 (N_19009,N_14999,N_15859);
nand U19010 (N_19010,N_15246,N_14993);
xnor U19011 (N_19011,N_14000,N_13048);
nand U19012 (N_19012,N_12191,N_12073);
or U19013 (N_19013,N_13031,N_16721);
xnor U19014 (N_19014,N_12864,N_16323);
nor U19015 (N_19015,N_14960,N_16866);
and U19016 (N_19016,N_16922,N_14040);
nor U19017 (N_19017,N_12364,N_12068);
and U19018 (N_19018,N_17750,N_16201);
or U19019 (N_19019,N_15396,N_12758);
and U19020 (N_19020,N_16930,N_14306);
and U19021 (N_19021,N_13600,N_12459);
nand U19022 (N_19022,N_14380,N_15328);
and U19023 (N_19023,N_13334,N_17270);
nor U19024 (N_19024,N_16515,N_15456);
nor U19025 (N_19025,N_15527,N_16787);
xnor U19026 (N_19026,N_17190,N_17553);
and U19027 (N_19027,N_12473,N_13467);
xor U19028 (N_19028,N_14656,N_13006);
and U19029 (N_19029,N_13576,N_15894);
xor U19030 (N_19030,N_15773,N_17956);
xor U19031 (N_19031,N_12485,N_17080);
and U19032 (N_19032,N_13761,N_13158);
or U19033 (N_19033,N_13273,N_15605);
and U19034 (N_19034,N_13394,N_15176);
nor U19035 (N_19035,N_17286,N_15421);
xnor U19036 (N_19036,N_12098,N_14549);
xor U19037 (N_19037,N_12151,N_12627);
xor U19038 (N_19038,N_16443,N_14435);
and U19039 (N_19039,N_12492,N_16781);
nand U19040 (N_19040,N_12940,N_13851);
xnor U19041 (N_19041,N_14683,N_17253);
nor U19042 (N_19042,N_17557,N_14868);
or U19043 (N_19043,N_17432,N_17278);
and U19044 (N_19044,N_15067,N_15961);
nand U19045 (N_19045,N_15283,N_15254);
nand U19046 (N_19046,N_12044,N_12536);
xnor U19047 (N_19047,N_13236,N_13290);
nor U19048 (N_19048,N_12805,N_16194);
and U19049 (N_19049,N_17576,N_17138);
or U19050 (N_19050,N_16024,N_13768);
xnor U19051 (N_19051,N_16319,N_12503);
xor U19052 (N_19052,N_12688,N_17951);
nand U19053 (N_19053,N_12392,N_12071);
xnor U19054 (N_19054,N_12741,N_12371);
nand U19055 (N_19055,N_14417,N_12966);
or U19056 (N_19056,N_16016,N_13168);
nand U19057 (N_19057,N_12949,N_15029);
or U19058 (N_19058,N_17046,N_12180);
xnor U19059 (N_19059,N_15838,N_13241);
nand U19060 (N_19060,N_12483,N_14270);
xnor U19061 (N_19061,N_17030,N_15221);
or U19062 (N_19062,N_16590,N_15073);
and U19063 (N_19063,N_16132,N_14276);
or U19064 (N_19064,N_14013,N_16595);
xor U19065 (N_19065,N_16824,N_15349);
or U19066 (N_19066,N_14293,N_16407);
nor U19067 (N_19067,N_16543,N_14467);
and U19068 (N_19068,N_13719,N_14952);
nor U19069 (N_19069,N_14867,N_14237);
nor U19070 (N_19070,N_12206,N_14657);
xnor U19071 (N_19071,N_16743,N_14563);
nor U19072 (N_19072,N_12280,N_12569);
nor U19073 (N_19073,N_14671,N_12502);
or U19074 (N_19074,N_12790,N_13414);
nor U19075 (N_19075,N_12304,N_17659);
or U19076 (N_19076,N_17074,N_15260);
xnor U19077 (N_19077,N_17785,N_15723);
and U19078 (N_19078,N_15306,N_15187);
or U19079 (N_19079,N_16825,N_14207);
nor U19080 (N_19080,N_15289,N_15559);
or U19081 (N_19081,N_12244,N_16038);
xor U19082 (N_19082,N_13430,N_16929);
or U19083 (N_19083,N_16139,N_15706);
xnor U19084 (N_19084,N_12372,N_14301);
or U19085 (N_19085,N_17994,N_15377);
and U19086 (N_19086,N_16172,N_14331);
nand U19087 (N_19087,N_17071,N_17509);
nor U19088 (N_19088,N_15475,N_15892);
nand U19089 (N_19089,N_13962,N_16106);
nor U19090 (N_19090,N_14680,N_13628);
and U19091 (N_19091,N_13544,N_14378);
and U19092 (N_19092,N_17196,N_12863);
nand U19093 (N_19093,N_16375,N_13370);
nor U19094 (N_19094,N_15955,N_14307);
or U19095 (N_19095,N_17255,N_16791);
xnor U19096 (N_19096,N_14658,N_15464);
xnor U19097 (N_19097,N_14956,N_13617);
nand U19098 (N_19098,N_13642,N_14209);
or U19099 (N_19099,N_12396,N_12262);
nor U19100 (N_19100,N_12906,N_15713);
or U19101 (N_19101,N_13005,N_15694);
nand U19102 (N_19102,N_13733,N_16242);
nor U19103 (N_19103,N_17960,N_14124);
and U19104 (N_19104,N_13223,N_17817);
or U19105 (N_19105,N_16348,N_13679);
or U19106 (N_19106,N_17299,N_14798);
nor U19107 (N_19107,N_15717,N_15684);
xor U19108 (N_19108,N_13886,N_14533);
nand U19109 (N_19109,N_13074,N_16399);
xnor U19110 (N_19110,N_17582,N_12650);
nor U19111 (N_19111,N_16539,N_15565);
or U19112 (N_19112,N_17279,N_15397);
nand U19113 (N_19113,N_12264,N_16035);
nand U19114 (N_19114,N_13003,N_13468);
or U19115 (N_19115,N_17501,N_13352);
xnor U19116 (N_19116,N_15372,N_13627);
nand U19117 (N_19117,N_17209,N_14411);
nand U19118 (N_19118,N_17781,N_17623);
xor U19119 (N_19119,N_15470,N_15414);
xor U19120 (N_19120,N_14774,N_12792);
nor U19121 (N_19121,N_13056,N_14612);
nor U19122 (N_19122,N_16617,N_14206);
or U19123 (N_19123,N_12938,N_15152);
and U19124 (N_19124,N_16623,N_16505);
nor U19125 (N_19125,N_17362,N_16772);
nor U19126 (N_19126,N_17227,N_14487);
xnor U19127 (N_19127,N_13538,N_13362);
nand U19128 (N_19128,N_16305,N_12601);
or U19129 (N_19129,N_12110,N_17139);
xnor U19130 (N_19130,N_12700,N_12528);
or U19131 (N_19131,N_15966,N_14753);
nor U19132 (N_19132,N_12132,N_12723);
xnor U19133 (N_19133,N_17852,N_16654);
xnor U19134 (N_19134,N_15364,N_16950);
nand U19135 (N_19135,N_17359,N_12783);
xnor U19136 (N_19136,N_17086,N_16935);
and U19137 (N_19137,N_15116,N_14120);
xnor U19138 (N_19138,N_13131,N_17262);
xor U19139 (N_19139,N_14096,N_14521);
or U19140 (N_19140,N_13242,N_12200);
or U19141 (N_19141,N_15225,N_15114);
nand U19142 (N_19142,N_15756,N_16897);
xnor U19143 (N_19143,N_16131,N_13681);
and U19144 (N_19144,N_13989,N_13089);
or U19145 (N_19145,N_12880,N_15687);
nor U19146 (N_19146,N_14264,N_12375);
nand U19147 (N_19147,N_15269,N_14696);
xnor U19148 (N_19148,N_13418,N_14578);
nor U19149 (N_19149,N_17671,N_17816);
and U19150 (N_19150,N_12186,N_15676);
nand U19151 (N_19151,N_12309,N_13045);
or U19152 (N_19152,N_17172,N_13613);
xor U19153 (N_19153,N_13466,N_16339);
or U19154 (N_19154,N_16991,N_14935);
or U19155 (N_19155,N_17283,N_14254);
or U19156 (N_19156,N_14212,N_14484);
nor U19157 (N_19157,N_13073,N_16047);
xor U19158 (N_19158,N_12432,N_14610);
xnor U19159 (N_19159,N_13203,N_16734);
nand U19160 (N_19160,N_16028,N_16338);
or U19161 (N_19161,N_16958,N_12107);
nand U19162 (N_19162,N_13898,N_12706);
nor U19163 (N_19163,N_13476,N_16080);
and U19164 (N_19164,N_17011,N_14051);
and U19165 (N_19165,N_16254,N_13790);
xnor U19166 (N_19166,N_17416,N_14561);
nand U19167 (N_19167,N_15958,N_16637);
or U19168 (N_19168,N_16180,N_17571);
nor U19169 (N_19169,N_16137,N_12971);
and U19170 (N_19170,N_14499,N_14616);
nand U19171 (N_19171,N_16185,N_12460);
xnor U19172 (N_19172,N_16939,N_15047);
nand U19173 (N_19173,N_17095,N_15833);
nor U19174 (N_19174,N_14127,N_16395);
nand U19175 (N_19175,N_14553,N_16512);
xnor U19176 (N_19176,N_17929,N_12350);
nand U19177 (N_19177,N_17891,N_14463);
nand U19178 (N_19178,N_14717,N_16166);
nand U19179 (N_19179,N_16067,N_17339);
and U19180 (N_19180,N_12791,N_17877);
or U19181 (N_19181,N_14446,N_13484);
and U19182 (N_19182,N_14046,N_17409);
and U19183 (N_19183,N_12041,N_12675);
and U19184 (N_19184,N_12857,N_16100);
xnor U19185 (N_19185,N_17866,N_15365);
and U19186 (N_19186,N_14936,N_17647);
and U19187 (N_19187,N_13702,N_15340);
xor U19188 (N_19188,N_17824,N_16156);
nand U19189 (N_19189,N_14092,N_16649);
and U19190 (N_19190,N_13170,N_17090);
nor U19191 (N_19191,N_15598,N_13606);
nand U19192 (N_19192,N_16628,N_17128);
and U19193 (N_19193,N_12731,N_16709);
and U19194 (N_19194,N_16317,N_15112);
or U19195 (N_19195,N_13220,N_17068);
nand U19196 (N_19196,N_12626,N_12347);
nand U19197 (N_19197,N_17485,N_14432);
or U19198 (N_19198,N_13357,N_14160);
nand U19199 (N_19199,N_16823,N_12947);
or U19200 (N_19200,N_14539,N_16795);
and U19201 (N_19201,N_17907,N_17159);
nand U19202 (N_19202,N_13471,N_13305);
xor U19203 (N_19203,N_15974,N_14336);
xor U19204 (N_19204,N_16032,N_12644);
nor U19205 (N_19205,N_15219,N_13866);
xnor U19206 (N_19206,N_16245,N_16737);
nor U19207 (N_19207,N_12125,N_15637);
nor U19208 (N_19208,N_14804,N_15922);
nand U19209 (N_19209,N_16834,N_13660);
nor U19210 (N_19210,N_16527,N_14345);
nor U19211 (N_19211,N_13176,N_13293);
xor U19212 (N_19212,N_14916,N_13651);
nor U19213 (N_19213,N_15846,N_17198);
nand U19214 (N_19214,N_12438,N_14714);
nand U19215 (N_19215,N_12592,N_15303);
or U19216 (N_19216,N_14137,N_16808);
nor U19217 (N_19217,N_15205,N_15195);
nand U19218 (N_19218,N_16396,N_17910);
nor U19219 (N_19219,N_13910,N_16482);
xor U19220 (N_19220,N_13846,N_14698);
or U19221 (N_19221,N_15249,N_13629);
xor U19222 (N_19222,N_12119,N_16269);
nor U19223 (N_19223,N_14227,N_16022);
or U19224 (N_19224,N_16644,N_17027);
nand U19225 (N_19225,N_16607,N_17117);
nor U19226 (N_19226,N_15898,N_13335);
or U19227 (N_19227,N_14977,N_12285);
and U19228 (N_19228,N_13589,N_13823);
and U19229 (N_19229,N_13709,N_17861);
and U19230 (N_19230,N_17392,N_17292);
or U19231 (N_19231,N_14371,N_16236);
nor U19232 (N_19232,N_17428,N_13115);
nor U19233 (N_19233,N_14413,N_12945);
xnor U19234 (N_19234,N_15075,N_12760);
nor U19235 (N_19235,N_12683,N_13075);
nor U19236 (N_19236,N_14059,N_14304);
nor U19237 (N_19237,N_13825,N_16979);
xor U19238 (N_19238,N_15192,N_12002);
xor U19239 (N_19239,N_12510,N_17592);
nand U19240 (N_19240,N_12340,N_14770);
xnor U19241 (N_19241,N_14809,N_13667);
nor U19242 (N_19242,N_16530,N_17178);
nor U19243 (N_19243,N_15600,N_15540);
or U19244 (N_19244,N_16303,N_16954);
nand U19245 (N_19245,N_16423,N_12747);
xor U19246 (N_19246,N_15403,N_12562);
or U19247 (N_19247,N_15330,N_16943);
and U19248 (N_19248,N_15059,N_12049);
nor U19249 (N_19249,N_14149,N_17534);
xnor U19250 (N_19250,N_12929,N_13736);
xor U19251 (N_19251,N_17992,N_14659);
and U19252 (N_19252,N_17004,N_14891);
and U19253 (N_19253,N_16899,N_15936);
or U19254 (N_19254,N_14601,N_15380);
or U19255 (N_19255,N_17026,N_15934);
nor U19256 (N_19256,N_12812,N_13435);
nor U19257 (N_19257,N_16148,N_16454);
xor U19258 (N_19258,N_16523,N_14904);
nand U19259 (N_19259,N_17727,N_12511);
nand U19260 (N_19260,N_12249,N_17911);
and U19261 (N_19261,N_12727,N_17489);
xnor U19262 (N_19262,N_15253,N_16381);
nand U19263 (N_19263,N_17040,N_12239);
nor U19264 (N_19264,N_13199,N_15969);
nand U19265 (N_19265,N_14025,N_17724);
nand U19266 (N_19266,N_15522,N_14216);
nor U19267 (N_19267,N_17381,N_15096);
nand U19268 (N_19268,N_14613,N_14668);
xnor U19269 (N_19269,N_15472,N_17613);
nand U19270 (N_19270,N_17154,N_16147);
nor U19271 (N_19271,N_13940,N_17602);
nand U19272 (N_19272,N_12064,N_13611);
or U19273 (N_19273,N_15025,N_14184);
xor U19274 (N_19274,N_12836,N_14319);
and U19275 (N_19275,N_12529,N_15103);
nor U19276 (N_19276,N_13254,N_14470);
and U19277 (N_19277,N_17101,N_12225);
or U19278 (N_19278,N_12630,N_12780);
nand U19279 (N_19279,N_14806,N_15742);
or U19280 (N_19280,N_13460,N_12458);
nand U19281 (N_19281,N_12282,N_12619);
nand U19282 (N_19282,N_16345,N_17968);
xnor U19283 (N_19283,N_13093,N_15864);
nor U19284 (N_19284,N_16673,N_13034);
or U19285 (N_19285,N_17272,N_14242);
nand U19286 (N_19286,N_12424,N_16241);
and U19287 (N_19287,N_15373,N_16882);
xor U19288 (N_19288,N_15366,N_17105);
xnor U19289 (N_19289,N_12192,N_12227);
xnor U19290 (N_19290,N_16620,N_14802);
xor U19291 (N_19291,N_14273,N_16962);
or U19292 (N_19292,N_15524,N_12417);
nand U19293 (N_19293,N_16759,N_15858);
nor U19294 (N_19294,N_15334,N_12663);
and U19295 (N_19295,N_17149,N_13224);
nand U19296 (N_19296,N_16794,N_17066);
and U19297 (N_19297,N_13756,N_14339);
or U19298 (N_19298,N_14249,N_15545);
nor U19299 (N_19299,N_12351,N_17822);
xnor U19300 (N_19300,N_12685,N_13906);
nand U19301 (N_19301,N_15731,N_12323);
or U19302 (N_19302,N_15521,N_14320);
nand U19303 (N_19303,N_13085,N_13859);
xor U19304 (N_19304,N_15995,N_15004);
and U19305 (N_19305,N_15659,N_14715);
and U19306 (N_19306,N_17991,N_17600);
nor U19307 (N_19307,N_13080,N_12081);
nor U19308 (N_19308,N_13811,N_15137);
and U19309 (N_19309,N_15874,N_14253);
xor U19310 (N_19310,N_16334,N_12870);
nor U19311 (N_19311,N_16372,N_13033);
nand U19312 (N_19312,N_14133,N_12659);
and U19313 (N_19313,N_14223,N_12509);
or U19314 (N_19314,N_13215,N_16890);
nand U19315 (N_19315,N_12320,N_15549);
nor U19316 (N_19316,N_15222,N_12365);
and U19317 (N_19317,N_13123,N_15798);
nand U19318 (N_19318,N_14224,N_12287);
nor U19319 (N_19319,N_17225,N_17056);
nand U19320 (N_19320,N_13562,N_14021);
nand U19321 (N_19321,N_12115,N_16719);
nor U19322 (N_19322,N_12531,N_12496);
nand U19323 (N_19323,N_14858,N_17775);
or U19324 (N_19324,N_12270,N_16560);
nand U19325 (N_19325,N_16112,N_16358);
nand U19326 (N_19326,N_14177,N_15428);
or U19327 (N_19327,N_15817,N_15767);
xnor U19328 (N_19328,N_12796,N_12825);
and U19329 (N_19329,N_17915,N_16513);
nand U19330 (N_19330,N_14486,N_17405);
nor U19331 (N_19331,N_14122,N_17638);
xor U19332 (N_19332,N_16547,N_15554);
nor U19333 (N_19333,N_13196,N_15488);
or U19334 (N_19334,N_15899,N_17726);
or U19335 (N_19335,N_17806,N_13438);
and U19336 (N_19336,N_16992,N_15682);
and U19337 (N_19337,N_13930,N_17167);
or U19338 (N_19338,N_14188,N_13907);
and U19339 (N_19339,N_17793,N_17763);
or U19340 (N_19340,N_13050,N_12597);
nor U19341 (N_19341,N_16329,N_14924);
and U19342 (N_19342,N_12654,N_17701);
nor U19343 (N_19343,N_14783,N_15111);
nor U19344 (N_19344,N_14144,N_16769);
nand U19345 (N_19345,N_14148,N_15347);
xnor U19346 (N_19346,N_12118,N_14800);
or U19347 (N_19347,N_14713,N_13010);
xnor U19348 (N_19348,N_13132,N_12159);
nor U19349 (N_19349,N_15640,N_12465);
nor U19350 (N_19350,N_16082,N_17945);
or U19351 (N_19351,N_14063,N_16480);
xor U19352 (N_19352,N_15474,N_12147);
nand U19353 (N_19353,N_16936,N_16766);
xor U19354 (N_19354,N_17307,N_14395);
nand U19355 (N_19355,N_16851,N_15077);
nor U19356 (N_19356,N_17525,N_12267);
or U19357 (N_19357,N_16222,N_14005);
xor U19358 (N_19358,N_16598,N_17430);
and U19359 (N_19359,N_15449,N_14332);
xnor U19360 (N_19360,N_14260,N_12996);
nand U19361 (N_19361,N_12631,N_14186);
and U19362 (N_19362,N_16071,N_17177);
and U19363 (N_19363,N_15392,N_13862);
nand U19364 (N_19364,N_17391,N_15802);
xor U19365 (N_19365,N_17067,N_12638);
nand U19366 (N_19366,N_15783,N_17215);
xnor U19367 (N_19367,N_17770,N_12015);
and U19368 (N_19368,N_14745,N_15983);
or U19369 (N_19369,N_15960,N_12718);
or U19370 (N_19370,N_12934,N_15031);
and U19371 (N_19371,N_15636,N_17521);
nand U19372 (N_19372,N_15026,N_16158);
nor U19373 (N_19373,N_14365,N_14857);
xor U19374 (N_19374,N_17733,N_12055);
nand U19375 (N_19375,N_13405,N_17222);
or U19376 (N_19376,N_13046,N_13509);
nor U19377 (N_19377,N_17858,N_12415);
nor U19378 (N_19378,N_17636,N_13550);
and U19379 (N_19379,N_17928,N_15248);
xnor U19380 (N_19380,N_12743,N_12816);
or U19381 (N_19381,N_16618,N_17799);
and U19382 (N_19382,N_14735,N_14766);
nand U19383 (N_19383,N_14996,N_16633);
xor U19384 (N_19384,N_12034,N_14441);
and U19385 (N_19385,N_15850,N_14888);
xor U19386 (N_19386,N_14598,N_17000);
nor U19387 (N_19387,N_15893,N_16651);
and U19388 (N_19388,N_14954,N_17735);
nor U19389 (N_19389,N_12052,N_13327);
xor U19390 (N_19390,N_12567,N_16235);
xor U19391 (N_19391,N_17731,N_12750);
nor U19392 (N_19392,N_13536,N_15729);
or U19393 (N_19393,N_13680,N_15938);
nor U19394 (N_19394,N_12641,N_14739);
nor U19395 (N_19395,N_13427,N_15992);
or U19396 (N_19396,N_15567,N_14569);
xnor U19397 (N_19397,N_17224,N_17131);
nand U19398 (N_19398,N_13369,N_14110);
and U19399 (N_19399,N_17467,N_16891);
or U19400 (N_19400,N_12376,N_12090);
and U19401 (N_19401,N_12594,N_13265);
nand U19402 (N_19402,N_13579,N_16008);
xnor U19403 (N_19403,N_13424,N_12367);
nor U19404 (N_19404,N_15304,N_15155);
and U19405 (N_19405,N_16819,N_13495);
nand U19406 (N_19406,N_14666,N_12362);
and U19407 (N_19407,N_14591,N_13432);
and U19408 (N_19408,N_14508,N_16209);
nor U19409 (N_19409,N_13047,N_17986);
and U19410 (N_19410,N_14777,N_15185);
nand U19411 (N_19411,N_14913,N_17481);
xnor U19412 (N_19412,N_16949,N_13889);
nand U19413 (N_19413,N_13313,N_15681);
xor U19414 (N_19414,N_17764,N_17655);
or U19415 (N_19415,N_13734,N_15019);
and U19416 (N_19416,N_16359,N_13821);
or U19417 (N_19417,N_15652,N_15190);
and U19418 (N_19418,N_15308,N_16325);
and U19419 (N_19419,N_17218,N_14349);
xor U19420 (N_19420,N_14532,N_14481);
xor U19421 (N_19421,N_17152,N_12007);
and U19422 (N_19422,N_12393,N_15280);
xor U19423 (N_19423,N_13515,N_14661);
nand U19424 (N_19424,N_14367,N_14167);
xnor U19425 (N_19425,N_15914,N_15552);
xor U19426 (N_19426,N_13603,N_15128);
nand U19427 (N_19427,N_12746,N_15738);
or U19428 (N_19428,N_14801,N_14682);
or U19429 (N_19429,N_15006,N_16792);
and U19430 (N_19430,N_12959,N_16040);
xor U19431 (N_19431,N_12389,N_12105);
nand U19432 (N_19432,N_12673,N_12818);
or U19433 (N_19433,N_12560,N_12279);
nor U19434 (N_19434,N_15539,N_16542);
xor U19435 (N_19435,N_12910,N_16469);
or U19436 (N_19436,N_17870,N_15809);
or U19437 (N_19437,N_15355,N_15173);
nor U19438 (N_19438,N_14556,N_13967);
and U19439 (N_19439,N_17061,N_13760);
nor U19440 (N_19440,N_13058,N_15455);
xor U19441 (N_19441,N_16243,N_16300);
nor U19442 (N_19442,N_15098,N_15622);
and U19443 (N_19443,N_15056,N_12346);
nand U19444 (N_19444,N_15154,N_14483);
xnor U19445 (N_19445,N_16730,N_14756);
nor U19446 (N_19446,N_14466,N_17518);
nand U19447 (N_19447,N_16596,N_15193);
xor U19448 (N_19448,N_16535,N_14263);
or U19449 (N_19449,N_14642,N_13307);
and U19450 (N_19450,N_16995,N_13601);
xnor U19451 (N_19451,N_14667,N_14461);
and U19452 (N_19452,N_17633,N_14335);
xnor U19453 (N_19453,N_12577,N_17402);
nand U19454 (N_19454,N_12170,N_17808);
xor U19455 (N_19455,N_12690,N_12978);
nor U19456 (N_19456,N_14966,N_15507);
nand U19457 (N_19457,N_17599,N_16720);
and U19458 (N_19458,N_12975,N_17109);
and U19459 (N_19459,N_17685,N_16860);
nor U19460 (N_19460,N_16863,N_15730);
and U19461 (N_19461,N_17032,N_12596);
xor U19462 (N_19462,N_15170,N_16974);
or U19463 (N_19463,N_15429,N_14135);
and U19464 (N_19464,N_15483,N_17226);
nand U19465 (N_19465,N_16326,N_15979);
nand U19466 (N_19466,N_17964,N_17372);
xor U19467 (N_19467,N_12566,N_12357);
and U19468 (N_19468,N_17114,N_15700);
or U19469 (N_19469,N_15860,N_14101);
xnor U19470 (N_19470,N_16138,N_17678);
and U19471 (N_19471,N_17330,N_14010);
xor U19472 (N_19472,N_13026,N_14767);
or U19473 (N_19473,N_14769,N_12278);
nand U19474 (N_19474,N_14930,N_13255);
nor U19475 (N_19475,N_14027,N_14442);
nand U19476 (N_19476,N_14797,N_17353);
and U19477 (N_19477,N_15194,N_14851);
nor U19478 (N_19478,N_13752,N_16341);
nand U19479 (N_19479,N_14006,N_13714);
and U19480 (N_19480,N_13671,N_16199);
xnor U19481 (N_19481,N_15912,N_13598);
xor U19482 (N_19482,N_15239,N_13413);
nor U19483 (N_19483,N_12172,N_14811);
or U19484 (N_19484,N_17993,N_17541);
and U19485 (N_19485,N_17851,N_16459);
nor U19486 (N_19486,N_15814,N_13730);
nor U19487 (N_19487,N_14596,N_16599);
xor U19488 (N_19488,N_16021,N_13539);
or U19489 (N_19489,N_14577,N_12344);
nor U19490 (N_19490,N_16884,N_15288);
nor U19491 (N_19491,N_12859,N_12645);
xnor U19492 (N_19492,N_12286,N_14044);
or U19493 (N_19493,N_13775,N_16981);
nor U19494 (N_19494,N_16546,N_14452);
and U19495 (N_19495,N_14991,N_15321);
nand U19496 (N_19496,N_12724,N_16342);
nand U19497 (N_19497,N_15127,N_13364);
nor U19498 (N_19498,N_14351,N_17529);
nand U19499 (N_19499,N_16843,N_16859);
nor U19500 (N_19500,N_15883,N_14828);
or U19501 (N_19501,N_12879,N_15278);
and U19502 (N_19502,N_12860,N_17257);
xnor U19503 (N_19503,N_17620,N_14220);
nor U19504 (N_19504,N_16977,N_12865);
xor U19505 (N_19505,N_17981,N_12402);
or U19506 (N_19506,N_14495,N_16213);
or U19507 (N_19507,N_14065,N_14060);
xnor U19508 (N_19508,N_14646,N_14073);
or U19509 (N_19509,N_15990,N_15022);
nand U19510 (N_19510,N_17552,N_13528);
xor U19511 (N_19511,N_13653,N_15657);
nor U19512 (N_19512,N_12795,N_14856);
nor U19513 (N_19513,N_15704,N_13683);
or U19514 (N_19514,N_16401,N_15702);
nor U19515 (N_19515,N_17597,N_14898);
and U19516 (N_19516,N_15744,N_16405);
nand U19517 (N_19517,N_14305,N_16846);
and U19518 (N_19518,N_16708,N_14834);
nor U19519 (N_19519,N_15120,N_15633);
or U19520 (N_19520,N_12457,N_16761);
xnor U19521 (N_19521,N_12672,N_12404);
or U19522 (N_19522,N_14403,N_13958);
nand U19523 (N_19523,N_13207,N_16875);
nor U19524 (N_19524,N_16643,N_17079);
nor U19525 (N_19525,N_13829,N_17794);
xor U19526 (N_19526,N_15963,N_16879);
and U19527 (N_19527,N_14818,N_12348);
nor U19528 (N_19528,N_13091,N_15461);
nor U19529 (N_19529,N_16216,N_16548);
and U19530 (N_19530,N_15410,N_14286);
or U19531 (N_19531,N_15094,N_15273);
nand U19532 (N_19532,N_12302,N_15867);
nand U19533 (N_19533,N_12075,N_16508);
and U19534 (N_19534,N_13343,N_15174);
xor U19535 (N_19535,N_17901,N_16514);
nand U19536 (N_19536,N_16802,N_13391);
nand U19537 (N_19537,N_15569,N_14311);
xor U19538 (N_19538,N_15558,N_13853);
nand U19539 (N_19539,N_17652,N_16652);
and U19540 (N_19540,N_12154,N_17092);
and U19541 (N_19541,N_15124,N_15139);
or U19542 (N_19542,N_12093,N_14884);
xnor U19543 (N_19543,N_13867,N_16840);
xnor U19544 (N_19544,N_12014,N_13669);
nand U19545 (N_19545,N_15905,N_13251);
or U19546 (N_19546,N_13762,N_13218);
or U19547 (N_19547,N_13845,N_13828);
nand U19548 (N_19548,N_14287,N_17853);
nand U19549 (N_19549,N_15436,N_13971);
nand U19550 (N_19550,N_15329,N_16312);
nor U19551 (N_19551,N_13133,N_15642);
or U19552 (N_19552,N_12030,N_16306);
nand U19553 (N_19553,N_13517,N_17310);
xnor U19554 (N_19554,N_13700,N_12291);
and U19555 (N_19555,N_14692,N_14002);
nor U19556 (N_19556,N_16283,N_17060);
nand U19557 (N_19557,N_14032,N_13990);
nor U19558 (N_19558,N_14493,N_17936);
nor U19559 (N_19559,N_15310,N_13880);
or U19560 (N_19560,N_17323,N_13188);
or U19561 (N_19561,N_13558,N_17680);
nand U19562 (N_19562,N_15732,N_15771);
xor U19563 (N_19563,N_12869,N_17214);
or U19564 (N_19564,N_12273,N_15835);
nand U19565 (N_19565,N_15317,N_12856);
nor U19566 (N_19566,N_14969,N_12916);
xor U19567 (N_19567,N_12466,N_15175);
xnor U19568 (N_19568,N_15891,N_15750);
nor U19569 (N_19569,N_15544,N_13770);
xnor U19570 (N_19570,N_15189,N_13142);
or U19571 (N_19571,N_12418,N_16576);
xor U19572 (N_19572,N_14454,N_17547);
and U19573 (N_19573,N_15881,N_14129);
xnor U19574 (N_19574,N_16374,N_15626);
and U19575 (N_19575,N_14540,N_12197);
nand U19576 (N_19576,N_14294,N_17774);
nand U19577 (N_19577,N_14434,N_15276);
xor U19578 (N_19578,N_12152,N_17239);
and U19579 (N_19579,N_17930,N_14232);
nor U19580 (N_19580,N_16479,N_15032);
xor U19581 (N_19581,N_15721,N_15136);
nor U19582 (N_19582,N_15480,N_17717);
xor U19583 (N_19583,N_16976,N_17776);
and U19584 (N_19584,N_15035,N_12624);
nor U19585 (N_19585,N_13213,N_13908);
nor U19586 (N_19586,N_12640,N_13715);
nand U19587 (N_19587,N_13159,N_15182);
nor U19588 (N_19588,N_17668,N_14525);
nor U19589 (N_19589,N_12413,N_13099);
nand U19590 (N_19590,N_13751,N_15855);
nor U19591 (N_19591,N_12283,N_15250);
xor U19592 (N_19592,N_15489,N_16041);
or U19593 (N_19593,N_12378,N_14706);
and U19594 (N_19594,N_14669,N_17605);
nor U19595 (N_19595,N_12366,N_14009);
nor U19596 (N_19596,N_12824,N_17421);
nor U19597 (N_19597,N_15135,N_14255);
nand U19598 (N_19598,N_16506,N_16200);
xnor U19599 (N_19599,N_16674,N_15400);
xor U19600 (N_19600,N_16009,N_17959);
nand U19601 (N_19601,N_14588,N_12447);
nand U19602 (N_19602,N_16294,N_13675);
and U19603 (N_19603,N_12595,N_12556);
nand U19604 (N_19604,N_16806,N_16406);
xor U19605 (N_19605,N_13830,N_12053);
nor U19606 (N_19606,N_13546,N_13439);
or U19607 (N_19607,N_15267,N_12373);
and U19608 (N_19608,N_13899,N_14846);
and U19609 (N_19609,N_15923,N_14589);
and U19610 (N_19610,N_13883,N_14522);
or U19611 (N_19611,N_17974,N_13605);
nand U19612 (N_19612,N_15296,N_12722);
xor U19613 (N_19613,N_16838,N_13105);
nor U19614 (N_19614,N_15529,N_13098);
or U19615 (N_19615,N_14675,N_13941);
and U19616 (N_19616,N_12219,N_14565);
xor U19617 (N_19617,N_12807,N_16178);
and U19618 (N_19618,N_12708,N_17512);
nor U19619 (N_19619,N_14568,N_12374);
nor U19620 (N_19620,N_16594,N_14112);
nand U19621 (N_19621,N_14222,N_12000);
or U19622 (N_19622,N_15911,N_14068);
nor U19623 (N_19623,N_15234,N_14758);
or U19624 (N_19624,N_13153,N_13177);
xor U19625 (N_19625,N_12917,N_13375);
nor U19626 (N_19626,N_15378,N_14228);
nor U19627 (N_19627,N_13454,N_17112);
nand U19628 (N_19628,N_12188,N_14474);
or U19629 (N_19629,N_16219,N_12033);
xnor U19630 (N_19630,N_15679,N_16409);
nor U19631 (N_19631,N_14605,N_14074);
nor U19632 (N_19632,N_13553,N_13759);
xnor U19633 (N_19633,N_13916,N_13905);
nand U19634 (N_19634,N_17358,N_16656);
nor U19635 (N_19635,N_15388,N_12956);
nand U19636 (N_19636,N_17045,N_12810);
nand U19637 (N_19637,N_14457,N_13490);
or U19638 (N_19638,N_14392,N_14932);
and U19639 (N_19639,N_15902,N_12421);
and U19640 (N_19640,N_13402,N_13876);
nand U19641 (N_19641,N_17622,N_12759);
or U19642 (N_19642,N_16164,N_15542);
and U19643 (N_19643,N_12549,N_13178);
and U19644 (N_19644,N_15435,N_17168);
and U19645 (N_19645,N_12678,N_14291);
and U19646 (N_19646,N_13622,N_12452);
nand U19647 (N_19647,N_17940,N_13169);
nor U19648 (N_19648,N_14430,N_13140);
nor U19649 (N_19649,N_15331,N_17429);
or U19650 (N_19650,N_17924,N_15479);
xnor U19651 (N_19651,N_16916,N_16918);
nor U19652 (N_19652,N_13238,N_13452);
or U19653 (N_19653,N_12422,N_12369);
xnor U19654 (N_19654,N_13103,N_13540);
xnor U19655 (N_19655,N_12266,N_16102);
or U19656 (N_19656,N_13044,N_16603);
and U19657 (N_19657,N_14221,N_12611);
xnor U19658 (N_19658,N_17130,N_17083);
xnor U19659 (N_19659,N_17370,N_13688);
nand U19660 (N_19660,N_13463,N_13996);
nor U19661 (N_19661,N_15467,N_14815);
and U19662 (N_19662,N_14674,N_12894);
or U19663 (N_19663,N_14324,N_14376);
xnor U19664 (N_19664,N_16551,N_13052);
xnor U19665 (N_19665,N_13838,N_17967);
xnor U19666 (N_19666,N_12103,N_15093);
nor U19667 (N_19667,N_12590,N_12431);
or U19668 (N_19668,N_16130,N_17295);
nand U19669 (N_19669,N_14393,N_14041);
and U19670 (N_19670,N_12841,N_17308);
xor U19671 (N_19671,N_14437,N_17265);
and U19672 (N_19672,N_16970,N_16083);
and U19673 (N_19673,N_15062,N_15547);
xor U19674 (N_19674,N_16019,N_15423);
nand U19675 (N_19675,N_14123,N_13936);
nand U19676 (N_19676,N_14325,N_16055);
xor U19677 (N_19677,N_17242,N_12331);
nor U19678 (N_19678,N_16214,N_14885);
nor U19679 (N_19679,N_13525,N_15237);
nor U19680 (N_19680,N_15012,N_17417);
and U19681 (N_19681,N_13492,N_16029);
nor U19682 (N_19682,N_15690,N_12699);
or U19683 (N_19683,N_16383,N_14931);
nand U19684 (N_19684,N_15661,N_16579);
and U19685 (N_19685,N_13192,N_15705);
or U19686 (N_19686,N_12563,N_15555);
and U19687 (N_19687,N_14730,N_16660);
nand U19688 (N_19688,N_12253,N_13640);
nor U19689 (N_19689,N_13195,N_14278);
or U19690 (N_19690,N_16896,N_15030);
or U19691 (N_19691,N_12646,N_17111);
xnor U19692 (N_19692,N_15476,N_14218);
and U19693 (N_19693,N_16756,N_12558);
or U19694 (N_19694,N_16431,N_15977);
or U19695 (N_19695,N_15045,N_14303);
and U19696 (N_19696,N_15647,N_17536);
nand U19697 (N_19697,N_13999,N_13662);
xor U19698 (N_19698,N_12914,N_17192);
nand U19699 (N_19699,N_14776,N_17282);
and U19700 (N_19700,N_16015,N_17035);
nor U19701 (N_19701,N_12322,N_17729);
or U19702 (N_19702,N_15697,N_17464);
xor U19703 (N_19703,N_14429,N_17732);
or U19704 (N_19704,N_16248,N_12918);
or U19705 (N_19705,N_17573,N_15214);
and U19706 (N_19706,N_14742,N_16413);
and U19707 (N_19707,N_15370,N_12083);
or U19708 (N_19708,N_15213,N_12772);
nand U19709 (N_19709,N_16777,N_13154);
xnor U19710 (N_19710,N_16026,N_14251);
or U19711 (N_19711,N_17615,N_17663);
or U19712 (N_19712,N_13923,N_16371);
nor U19713 (N_19713,N_17106,N_13716);
and U19714 (N_19714,N_13666,N_12241);
xnor U19715 (N_19715,N_15765,N_12213);
and U19716 (N_19716,N_16626,N_12444);
nor U19717 (N_19717,N_16183,N_17099);
xor U19718 (N_19718,N_13507,N_13288);
or U19719 (N_19719,N_15937,N_16198);
nor U19720 (N_19720,N_13931,N_17230);
or U19721 (N_19721,N_15917,N_17850);
nor U19722 (N_19722,N_12974,N_12135);
and U19723 (N_19723,N_12635,N_16159);
nand U19724 (N_19724,N_16969,N_12097);
nor U19725 (N_19725,N_16789,N_17875);
nand U19726 (N_19726,N_12888,N_14473);
xnor U19727 (N_19727,N_16247,N_13062);
or U19728 (N_19728,N_15797,N_17263);
and U19729 (N_19729,N_17304,N_16911);
and U19730 (N_19730,N_12559,N_17497);
nor U19731 (N_19731,N_17053,N_13285);
nand U19732 (N_19732,N_12903,N_12709);
xor U19733 (N_19733,N_14523,N_16288);
nand U19734 (N_19734,N_14973,N_16056);
nor U19735 (N_19735,N_17803,N_15967);
and U19736 (N_19736,N_15653,N_13884);
and U19737 (N_19737,N_15786,N_15784);
or U19738 (N_19738,N_15085,N_15147);
and U19739 (N_19739,N_17472,N_13937);
nor U19740 (N_19740,N_13817,N_15643);
or U19741 (N_19741,N_16754,N_16123);
nor U19742 (N_19742,N_12175,N_14192);
nand U19743 (N_19743,N_16291,N_14266);
nand U19744 (N_19744,N_15293,N_17103);
nand U19745 (N_19745,N_12565,N_15714);
or U19746 (N_19746,N_15596,N_15915);
nor U19747 (N_19747,N_15819,N_14530);
and U19748 (N_19748,N_13753,N_16282);
and U19749 (N_19749,N_12557,N_16898);
and U19750 (N_19750,N_17739,N_15327);
or U19751 (N_19751,N_13421,N_16360);
nor U19752 (N_19752,N_14535,N_16600);
xor U19753 (N_19753,N_12078,N_12464);
nand U19754 (N_19754,N_13985,N_17932);
xor U19755 (N_19755,N_15374,N_14386);
and U19756 (N_19756,N_17935,N_14150);
xor U19757 (N_19757,N_12065,N_15079);
and U19758 (N_19758,N_17380,N_15381);
nor U19759 (N_19759,N_15384,N_13229);
nor U19760 (N_19760,N_13656,N_15927);
xor U19761 (N_19761,N_17276,N_13778);
and U19762 (N_19762,N_17431,N_17367);
nor U19763 (N_19763,N_14023,N_16996);
or U19764 (N_19764,N_16018,N_14855);
xor U19765 (N_19765,N_13565,N_16496);
nand U19766 (N_19766,N_12284,N_16336);
and U19767 (N_19767,N_12729,N_16809);
xnor U19768 (N_19768,N_16475,N_12775);
nand U19769 (N_19769,N_17881,N_16467);
or U19770 (N_19770,N_13634,N_14163);
nor U19771 (N_19771,N_17042,N_15160);
and U19772 (N_19772,N_13641,N_15069);
and U19773 (N_19773,N_14444,N_17333);
nand U19774 (N_19774,N_13506,N_14126);
and U19775 (N_19775,N_17478,N_15885);
and U19776 (N_19776,N_17356,N_12031);
nand U19777 (N_19777,N_15550,N_16934);
and U19778 (N_19778,N_15617,N_14825);
xor U19779 (N_19779,N_12174,N_12943);
nand U19780 (N_19780,N_14544,N_12048);
and U19781 (N_19781,N_17240,N_17673);
or U19782 (N_19782,N_13943,N_16615);
nand U19783 (N_19783,N_16239,N_15576);
and U19784 (N_19784,N_15024,N_12637);
and U19785 (N_19785,N_14917,N_13858);
nor U19786 (N_19786,N_14670,N_13771);
or U19787 (N_19787,N_15382,N_12096);
or U19788 (N_19788,N_15406,N_15796);
nor U19789 (N_19789,N_16073,N_12734);
and U19790 (N_19790,N_16098,N_16228);
xnor U19791 (N_19791,N_17175,N_12182);
and U19792 (N_19792,N_12142,N_16044);
and U19793 (N_19793,N_13960,N_17838);
nor U19794 (N_19794,N_15629,N_14426);
nand U19795 (N_19795,N_17841,N_13529);
xor U19796 (N_19796,N_15665,N_17594);
and U19797 (N_19797,N_14079,N_17014);
nand U19798 (N_19798,N_16807,N_16853);
and U19799 (N_19799,N_17725,N_14410);
xnor U19800 (N_19800,N_14820,N_13887);
or U19801 (N_19801,N_16592,N_14623);
nand U19802 (N_19802,N_16593,N_12133);
nor U19803 (N_19803,N_14399,N_13732);
nand U19804 (N_19804,N_12544,N_12583);
and U19805 (N_19805,N_13911,N_12840);
nand U19806 (N_19806,N_12092,N_13822);
nand U19807 (N_19807,N_12023,N_17744);
xnor U19808 (N_19808,N_15516,N_16313);
xnor U19809 (N_19809,N_14633,N_12513);
nor U19810 (N_19810,N_16129,N_13164);
nand U19811 (N_19811,N_13298,N_17805);
nand U19812 (N_19812,N_16361,N_17176);
and U19813 (N_19813,N_13247,N_16659);
nand U19814 (N_19814,N_13464,N_17598);
nand U19815 (N_19815,N_17640,N_12501);
or U19816 (N_19816,N_16762,N_14258);
and U19817 (N_19817,N_17958,N_17160);
nand U19818 (N_19818,N_17590,N_16435);
nand U19819 (N_19819,N_15650,N_15197);
and U19820 (N_19820,N_16119,N_14845);
or U19821 (N_19821,N_12789,N_17075);
nand U19822 (N_19822,N_15228,N_12184);
xnor U19823 (N_19823,N_14839,N_16037);
nor U19824 (N_19824,N_14751,N_17885);
xor U19825 (N_19825,N_15727,N_16993);
or U19826 (N_19826,N_13096,N_14456);
and U19827 (N_19827,N_17683,N_14882);
nor U19828 (N_19828,N_15803,N_14491);
and U19829 (N_19829,N_14196,N_14377);
nor U19830 (N_19830,N_13347,N_13473);
nor U19831 (N_19831,N_17962,N_17650);
nand U19832 (N_19832,N_14871,N_15118);
xor U19833 (N_19833,N_13498,N_17982);
nand U19834 (N_19834,N_15162,N_15582);
nand U19835 (N_19835,N_17798,N_12328);
nand U19836 (N_19836,N_12251,N_13332);
and U19837 (N_19837,N_12622,N_17002);
nand U19838 (N_19838,N_13505,N_13368);
xnor U19839 (N_19839,N_13703,N_14140);
nand U19840 (N_19840,N_12141,N_17987);
nor U19841 (N_19841,N_12202,N_12297);
nand U19842 (N_19842,N_17524,N_12397);
or U19843 (N_19843,N_17228,N_12298);
and U19844 (N_19844,N_17260,N_13061);
xnor U19845 (N_19845,N_12937,N_14115);
nand U19846 (N_19846,N_14678,N_14170);
or U19847 (N_19847,N_13514,N_17306);
nand U19848 (N_19848,N_14614,N_13429);
nor U19849 (N_19849,N_16941,N_16955);
or U19850 (N_19850,N_17711,N_15312);
or U19851 (N_19851,N_14500,N_13608);
nand U19852 (N_19852,N_17059,N_15581);
xor U19853 (N_19853,N_12961,N_15848);
nor U19854 (N_19854,N_13643,N_15904);
or U19855 (N_19855,N_17723,N_15439);
xor U19856 (N_19856,N_15407,N_17320);
nand U19857 (N_19857,N_13557,N_13328);
xor U19858 (N_19858,N_14501,N_13116);
nand U19859 (N_19859,N_16273,N_16997);
and U19860 (N_19860,N_17624,N_16550);
nand U19861 (N_19861,N_15916,N_15005);
xnor U19862 (N_19862,N_17818,N_16299);
or U19863 (N_19863,N_14512,N_14907);
or U19864 (N_19864,N_12352,N_16553);
or U19865 (N_19865,N_14546,N_16668);
and U19866 (N_19866,N_15606,N_13776);
nand U19867 (N_19867,N_17314,N_12703);
nor U19868 (N_19868,N_13946,N_12072);
nor U19869 (N_19869,N_13185,N_17245);
nand U19870 (N_19870,N_14841,N_17586);
nor U19871 (N_19871,N_17048,N_15788);
nor U19872 (N_19872,N_14215,N_14239);
and U19873 (N_19873,N_14001,N_15941);
and U19874 (N_19874,N_15149,N_15877);
nor U19875 (N_19875,N_16912,N_17350);
nand U19876 (N_19876,N_12259,N_14372);
xnor U19877 (N_19877,N_16686,N_15947);
nand U19878 (N_19878,N_17539,N_17535);
nor U19879 (N_19879,N_16876,N_16886);
or U19880 (N_19880,N_14281,N_12693);
or U19881 (N_19881,N_12803,N_13346);
and U19882 (N_19882,N_14179,N_15656);
nand U19883 (N_19883,N_17906,N_12649);
nor U19884 (N_19884,N_15023,N_17618);
nor U19885 (N_19885,N_13847,N_16446);
or U19886 (N_19886,N_17927,N_15699);
and U19887 (N_19887,N_12248,N_12667);
or U19888 (N_19888,N_14961,N_12160);
and U19889 (N_19889,N_17490,N_15179);
nand U19890 (N_19890,N_17800,N_14796);
nand U19891 (N_19891,N_16189,N_12632);
and U19892 (N_19892,N_16695,N_16645);
or U19893 (N_19893,N_16689,N_17990);
nor U19894 (N_19894,N_12100,N_16726);
and U19895 (N_19895,N_16362,N_16017);
xor U19896 (N_19896,N_12837,N_16821);
nor U19897 (N_19897,N_14737,N_15499);
or U19898 (N_19898,N_15624,N_12620);
nor U19899 (N_19899,N_13620,N_13209);
and U19900 (N_19900,N_15639,N_14836);
or U19901 (N_19901,N_15257,N_13128);
nand U19902 (N_19902,N_14848,N_16672);
nand U19903 (N_19903,N_13261,N_13513);
xnor U19904 (N_19904,N_13766,N_16829);
nor U19905 (N_19905,N_17021,N_14290);
xor U19906 (N_19906,N_16304,N_15813);
xnor U19907 (N_19907,N_14309,N_17293);
xnor U19908 (N_19908,N_15999,N_13970);
xor U19909 (N_19909,N_12989,N_15722);
or U19910 (N_19910,N_15743,N_14636);
nand U19911 (N_19911,N_13428,N_14315);
nor U19912 (N_19912,N_16568,N_16706);
xor U19913 (N_19913,N_12294,N_14468);
or U19914 (N_19914,N_13796,N_13687);
and U19915 (N_19915,N_14757,N_15177);
xor U19916 (N_19916,N_13914,N_16636);
nor U19917 (N_19917,N_12913,N_17856);
and U19918 (N_19918,N_17738,N_16331);
and U19919 (N_19919,N_14998,N_16771);
and U19920 (N_19920,N_17679,N_12450);
or U19921 (N_19921,N_13353,N_17142);
or U19922 (N_19922,N_14672,N_14275);
nand U19923 (N_19923,N_14903,N_17587);
xnor U19924 (N_19924,N_13291,N_15604);
and U19925 (N_19925,N_13668,N_14183);
or U19926 (N_19926,N_13791,N_12258);
nor U19927 (N_19927,N_15871,N_15693);
nand U19928 (N_19928,N_16223,N_13713);
xnor U19929 (N_19929,N_13308,N_14881);
nor U19930 (N_19930,N_15878,N_15229);
nor U19931 (N_19931,N_16430,N_15404);
or U19932 (N_19932,N_17864,N_16117);
and U19933 (N_19933,N_15140,N_14176);
nand U19934 (N_19934,N_14011,N_14897);
xor U19935 (N_19935,N_14316,N_14047);
nor U19936 (N_19936,N_17251,N_17720);
nand U19937 (N_19937,N_17171,N_13857);
xor U19938 (N_19938,N_17017,N_14298);
xnor U19939 (N_19939,N_13701,N_12490);
xnor U19940 (N_19940,N_12676,N_15827);
xor U19941 (N_19941,N_17161,N_16050);
and U19942 (N_19942,N_16704,N_15415);
nor U19943 (N_19943,N_14964,N_14488);
xor U19944 (N_19944,N_16280,N_16457);
nor U19945 (N_19945,N_17691,N_14107);
xnor U19946 (N_19946,N_17922,N_15338);
nor U19947 (N_19947,N_17843,N_16648);
or U19948 (N_19948,N_13810,N_13015);
xor U19949 (N_19949,N_12479,N_15266);
or U19950 (N_19950,N_17387,N_13387);
xnor U19951 (N_19951,N_16999,N_15375);
or U19952 (N_19952,N_17748,N_12436);
or U19953 (N_19953,N_17173,N_15560);
nor U19954 (N_19954,N_15385,N_17480);
and U19955 (N_19955,N_12276,N_17835);
nor U19956 (N_19956,N_13554,N_16852);
nor U19957 (N_19957,N_14205,N_12623);
and U19958 (N_19958,N_17561,N_12426);
xor U19959 (N_19959,N_17029,N_16448);
and U19960 (N_19960,N_17118,N_14029);
nor U19961 (N_19961,N_12732,N_12326);
xor U19962 (N_19962,N_14720,N_13802);
nand U19963 (N_19963,N_14635,N_13039);
nor U19964 (N_19964,N_15134,N_17285);
nor U19965 (N_19965,N_13499,N_17008);
nand U19966 (N_19966,N_16268,N_16355);
nand U19967 (N_19967,N_16583,N_14972);
nand U19968 (N_19968,N_17033,N_16682);
nor U19969 (N_19969,N_15708,N_17269);
and U19970 (N_19970,N_16790,N_12024);
or U19971 (N_19971,N_16391,N_15976);
xor U19972 (N_19972,N_17373,N_13233);
and U19973 (N_19973,N_15710,N_14194);
or U19974 (N_19974,N_16998,N_15051);
nand U19975 (N_19975,N_12979,N_16773);
and U19976 (N_19976,N_15844,N_16314);
or U19977 (N_19977,N_17361,N_17538);
nor U19978 (N_19978,N_14030,N_17166);
and U19979 (N_19979,N_12842,N_15674);
or U19980 (N_19980,N_17018,N_17012);
nand U19981 (N_19981,N_16588,N_12574);
and U19982 (N_19982,N_17254,N_15042);
xor U19983 (N_19983,N_13087,N_13926);
xor U19984 (N_19984,N_14035,N_15281);
xor U19985 (N_19985,N_12476,N_13948);
xor U19986 (N_19986,N_16752,N_17876);
xor U19987 (N_19987,N_14449,N_12384);
and U19988 (N_19988,N_13269,N_16240);
nor U19989 (N_19989,N_17562,N_13189);
xor U19990 (N_19990,N_14519,N_13216);
nand U19991 (N_19991,N_16451,N_12134);
or U19992 (N_19992,N_14738,N_16885);
xor U19993 (N_19993,N_13077,N_12079);
xor U19994 (N_19994,N_17249,N_15052);
xnor U19995 (N_19995,N_12211,N_17972);
or U19996 (N_19996,N_12960,N_17354);
or U19997 (N_19997,N_15981,N_14915);
or U19998 (N_19998,N_17081,N_13774);
xor U19999 (N_19999,N_13239,N_17664);
nor U20000 (N_20000,N_15262,N_15933);
and U20001 (N_20001,N_12169,N_15001);
and U20002 (N_20002,N_12799,N_12877);
xor U20003 (N_20003,N_17187,N_16049);
or U20004 (N_20004,N_14125,N_12832);
nand U20005 (N_20005,N_13739,N_12108);
or U20006 (N_20006,N_12136,N_17382);
or U20007 (N_20007,N_14951,N_17975);
or U20008 (N_20008,N_14425,N_15018);
xor U20009 (N_20009,N_15800,N_16685);
nor U20010 (N_20010,N_13735,N_14723);
or U20011 (N_20011,N_17742,N_13146);
nand U20012 (N_20012,N_12976,N_15971);
nor U20013 (N_20013,N_12486,N_13824);
nand U20014 (N_20014,N_13028,N_14518);
and U20015 (N_20015,N_14807,N_15302);
xor U20016 (N_20016,N_14548,N_16973);
and U20017 (N_20017,N_15469,N_13582);
nand U20018 (N_20018,N_17871,N_14892);
nor U20019 (N_20019,N_16753,N_14707);
xnor U20020 (N_20020,N_13920,N_16179);
xor U20021 (N_20021,N_13356,N_17444);
or U20022 (N_20022,N_12963,N_17507);
nand U20023 (N_20023,N_16398,N_14054);
nand U20024 (N_20024,N_16193,N_15748);
nand U20025 (N_20025,N_15181,N_12621);
or U20026 (N_20026,N_17344,N_16410);
and U20027 (N_20027,N_12067,N_16907);
nand U20028 (N_20028,N_13785,N_13677);
or U20029 (N_20029,N_14053,N_13518);
nand U20030 (N_20030,N_15930,N_13032);
nand U20031 (N_20031,N_15123,N_17569);
nor U20032 (N_20032,N_14292,N_15599);
and U20033 (N_20033,N_15027,N_14992);
and U20034 (N_20034,N_16865,N_16445);
nand U20035 (N_20035,N_14673,N_16956);
xnor U20036 (N_20036,N_15117,N_15242);
nand U20037 (N_20037,N_17859,N_16931);
or U20038 (N_20038,N_17365,N_13127);
nand U20039 (N_20039,N_15601,N_15965);
or U20040 (N_20040,N_13069,N_13502);
nand U20041 (N_20041,N_16735,N_14102);
nor U20042 (N_20042,N_13386,N_17399);
or U20043 (N_20043,N_16393,N_13104);
and U20044 (N_20044,N_12753,N_16964);
nand U20045 (N_20045,N_15387,N_13234);
nand U20046 (N_20046,N_15395,N_16669);
or U20047 (N_20047,N_15357,N_12116);
or U20048 (N_20048,N_17837,N_17931);
and U20049 (N_20049,N_14896,N_16215);
or U20050 (N_20050,N_15716,N_14447);
or U20051 (N_20051,N_17426,N_15856);
nor U20052 (N_20052,N_12104,N_16005);
or U20053 (N_20053,N_16764,N_17704);
or U20054 (N_20054,N_15163,N_14772);
nand U20055 (N_20055,N_15962,N_13423);
xnor U20056 (N_20056,N_17277,N_13706);
or U20057 (N_20057,N_14593,N_13951);
and U20058 (N_20058,N_17349,N_13827);
xor U20059 (N_20059,N_16924,N_14641);
and U20060 (N_20060,N_14280,N_12598);
and U20061 (N_20061,N_13283,N_16389);
and U20062 (N_20062,N_14627,N_12946);
xor U20063 (N_20063,N_16366,N_16324);
and U20064 (N_20064,N_17702,N_16779);
nor U20065 (N_20065,N_13117,N_14440);
xnor U20066 (N_20066,N_13826,N_17483);
or U20067 (N_20067,N_13893,N_13854);
or U20068 (N_20068,N_12525,N_17692);
or U20069 (N_20069,N_12427,N_15523);
xor U20070 (N_20070,N_12385,N_17182);
and U20071 (N_20071,N_14524,N_14559);
nor U20072 (N_20072,N_17305,N_13070);
xnor U20073 (N_20073,N_17203,N_14765);
nor U20074 (N_20074,N_12908,N_12739);
and U20075 (N_20075,N_15368,N_15792);
and U20076 (N_20076,N_17697,N_12454);
and U20077 (N_20077,N_17610,N_15996);
or U20078 (N_20078,N_16880,N_12749);
nand U20079 (N_20079,N_15398,N_13148);
or U20080 (N_20080,N_14128,N_13674);
nand U20081 (N_20081,N_13266,N_15352);
xor U20082 (N_20082,N_15337,N_17593);
or U20083 (N_20083,N_15448,N_14262);
or U20084 (N_20084,N_16328,N_17575);
nand U20085 (N_20085,N_17185,N_14049);
xnor U20086 (N_20086,N_16070,N_12201);
nand U20087 (N_20087,N_12614,N_17447);
nand U20088 (N_20088,N_17237,N_13461);
and U20089 (N_20089,N_16850,N_17942);
or U20090 (N_20090,N_12056,N_13171);
nor U20091 (N_20091,N_15320,N_12517);
or U20092 (N_20092,N_15685,N_17705);
nand U20093 (N_20093,N_17498,N_17658);
and U20094 (N_20094,N_16571,N_14812);
xnor U20095 (N_20095,N_13324,N_15880);
and U20096 (N_20096,N_16150,N_16494);
xnor U20097 (N_20097,N_13879,N_13102);
or U20098 (N_20098,N_15907,N_12246);
and U20099 (N_20099,N_17025,N_14357);
nor U20100 (N_20100,N_14382,N_13571);
and U20101 (N_20101,N_14057,N_13001);
and U20102 (N_20102,N_14959,N_17511);
nand U20103 (N_20103,N_17637,N_15000);
nor U20104 (N_20104,N_13630,N_17461);
and U20105 (N_20105,N_17448,N_13954);
xnor U20106 (N_20106,N_15468,N_14894);
and U20107 (N_20107,N_15805,N_14173);
and U20108 (N_20108,N_14645,N_13616);
and U20109 (N_20109,N_15326,N_16478);
nand U20110 (N_20110,N_15009,N_13831);
xor U20111 (N_20111,N_16495,N_13661);
xnor U20112 (N_20112,N_14465,N_16511);
xnor U20113 (N_20113,N_16755,N_17243);
xnor U20114 (N_20114,N_15153,N_13166);
xnor U20115 (N_20115,N_12777,N_12822);
nor U20116 (N_20116,N_17813,N_13837);
or U20117 (N_20117,N_13692,N_12038);
and U20118 (N_20118,N_17855,N_13294);
or U20119 (N_20119,N_16447,N_13888);
or U20120 (N_20120,N_13474,N_15651);
or U20121 (N_20121,N_16350,N_15888);
nor U20122 (N_20122,N_14200,N_16487);
xor U20123 (N_20123,N_17514,N_16570);
and U20124 (N_20124,N_17324,N_17758);
and U20125 (N_20125,N_17908,N_17694);
or U20126 (N_20126,N_13051,N_17905);
nand U20127 (N_20127,N_17846,N_12878);
and U20128 (N_20128,N_16975,N_15361);
xnor U20129 (N_20129,N_17434,N_12798);
nor U20130 (N_20130,N_12238,N_12820);
nor U20131 (N_20131,N_17404,N_17487);
xnor U20132 (N_20132,N_17345,N_16400);
and U20133 (N_20133,N_17595,N_17193);
xnor U20134 (N_20134,N_15635,N_12647);
nor U20135 (N_20135,N_14793,N_12299);
or U20136 (N_20136,N_14075,N_17923);
nor U20137 (N_20137,N_15909,N_17229);
or U20138 (N_20138,N_17950,N_14943);
and U20139 (N_20139,N_16417,N_13798);
xor U20140 (N_20140,N_14394,N_12342);
and U20141 (N_20141,N_12815,N_14016);
nand U20142 (N_20142,N_13812,N_13455);
nor U20143 (N_20143,N_16120,N_14934);
nand U20144 (N_20144,N_12613,N_13917);
and U20145 (N_20145,N_13486,N_14346);
xnor U20146 (N_20146,N_16693,N_13956);
xor U20147 (N_20147,N_16462,N_12784);
and U20148 (N_20148,N_15259,N_12189);
and U20149 (N_20149,N_13186,N_14195);
xnor U20150 (N_20150,N_14919,N_15068);
nand U20151 (N_20151,N_17635,N_14958);
nor U20152 (N_20152,N_15772,N_15351);
and U20153 (N_20153,N_15807,N_14736);
and U20154 (N_20154,N_13023,N_14034);
and U20155 (N_20155,N_16045,N_14295);
nand U20156 (N_20156,N_15613,N_13311);
nor U20157 (N_20157,N_17772,N_13947);
nand U20158 (N_20158,N_13275,N_14217);
nor U20159 (N_20159,N_13808,N_13124);
xnor U20160 (N_20160,N_17542,N_17050);
or U20161 (N_20161,N_16274,N_15533);
xor U20162 (N_20162,N_17873,N_15551);
xnor U20163 (N_20163,N_17537,N_17440);
xor U20164 (N_20164,N_17007,N_12573);
nor U20165 (N_20165,N_13836,N_14852);
nor U20166 (N_20166,N_17648,N_16963);
and U20167 (N_20167,N_15517,N_14731);
xnor U20168 (N_20168,N_14269,N_16238);
nor U20169 (N_20169,N_17644,N_12891);
xor U20170 (N_20170,N_14404,N_16308);
or U20171 (N_20171,N_17563,N_16490);
nand U20172 (N_20172,N_14822,N_16917);
nor U20173 (N_20173,N_16007,N_14592);
xor U20174 (N_20174,N_15108,N_17757);
or U20175 (N_20175,N_13190,N_12318);
xnor U20176 (N_20176,N_15413,N_16871);
and U20177 (N_20177,N_16251,N_13731);
or U20178 (N_20178,N_16938,N_13184);
or U20179 (N_20179,N_14795,N_13420);
or U20180 (N_20180,N_13245,N_15985);
and U20181 (N_20181,N_17886,N_12605);
nor U20182 (N_20182,N_14780,N_13552);
nand U20183 (N_20183,N_13263,N_15129);
and U20184 (N_20184,N_12548,N_12726);
nor U20185 (N_20185,N_16262,N_16813);
xnor U20186 (N_20186,N_12022,N_16946);
xnor U20187 (N_20187,N_17500,N_17374);
nand U20188 (N_20188,N_13619,N_13092);
xnor U20189 (N_20189,N_16631,N_13903);
nand U20190 (N_20190,N_12471,N_13978);
and U20191 (N_20191,N_15251,N_15295);
nand U20192 (N_20192,N_16920,N_12441);
nand U20193 (N_20193,N_17250,N_16279);
and U20194 (N_20194,N_15216,N_13625);
or U20195 (N_20195,N_14585,N_12551);
xnor U20196 (N_20196,N_12504,N_15130);
and U20197 (N_20197,N_13533,N_13816);
or U20198 (N_20198,N_13965,N_13809);
nand U20199 (N_20199,N_12313,N_16404);
nand U20200 (N_20200,N_13849,N_14185);
and U20201 (N_20201,N_12380,N_16171);
xnor U20202 (N_20202,N_12102,N_14459);
and U20203 (N_20203,N_12137,N_12391);
xor U20204 (N_20204,N_15161,N_17005);
or U20205 (N_20205,N_17984,N_16749);
xnor U20206 (N_20206,N_12481,N_17311);
nor U20207 (N_20207,N_13066,N_16498);
nand U20208 (N_20208,N_13259,N_12889);
or U20209 (N_20209,N_14603,N_14844);
nor U20210 (N_20210,N_13193,N_12215);
xor U20211 (N_20211,N_17801,N_16265);
nor U20212 (N_20212,N_12972,N_13913);
or U20213 (N_20213,N_14048,N_14310);
nand U20214 (N_20214,N_12744,N_15631);
or U20215 (N_20215,N_17094,N_14450);
or U20216 (N_20216,N_15747,N_15212);
xnor U20217 (N_20217,N_14528,N_15362);
or U20218 (N_20218,N_17325,N_15171);
nand U20219 (N_20219,N_12494,N_15987);
xnor U20220 (N_20220,N_14906,N_12060);
nand U20221 (N_20221,N_12109,N_13297);
or U20222 (N_20222,N_12854,N_15900);
or U20223 (N_20223,N_13268,N_14728);
nor U20224 (N_20224,N_15236,N_16655);
xor U20225 (N_20225,N_15210,N_14458);
or U20226 (N_20226,N_15367,N_14948);
nor U20227 (N_20227,N_12656,N_13206);
and U20228 (N_20228,N_15592,N_13358);
and U20229 (N_20229,N_13573,N_15670);
nor U20230 (N_20230,N_16346,N_12234);
or U20231 (N_20231,N_12973,N_12412);
nor U20232 (N_20232,N_17273,N_17009);
and U20233 (N_20233,N_17909,N_12210);
xor U20234 (N_20234,N_12395,N_15148);
xor U20235 (N_20235,N_12954,N_13079);
or U20236 (N_20236,N_14072,N_12851);
nand U20237 (N_20237,N_17134,N_15932);
nand U20238 (N_20238,N_12434,N_17918);
and U20239 (N_20239,N_14617,N_13459);
xnor U20240 (N_20240,N_14722,N_16582);
or U20241 (N_20241,N_15646,N_15437);
and U20242 (N_20242,N_13282,N_13365);
nand U20243 (N_20243,N_16569,N_13363);
xnor U20244 (N_20244,N_16690,N_17568);
xnor U20245 (N_20245,N_14070,N_12269);
nand U20246 (N_20246,N_13874,N_13374);
nand U20247 (N_20247,N_16746,N_13995);
and U20248 (N_20248,N_17520,N_14942);
xor U20249 (N_20249,N_16564,N_17630);
and U20250 (N_20250,N_17879,N_15774);
and U20251 (N_20251,N_16230,N_12042);
xnor U20252 (N_20252,N_16556,N_12231);
nor U20253 (N_20253,N_17452,N_12209);
nand U20254 (N_20254,N_13401,N_16261);
nand U20255 (N_20255,N_12681,N_13563);
nor U20256 (N_20256,N_16563,N_12037);
and U20257 (N_20257,N_16614,N_17943);
nand U20258 (N_20258,N_17064,N_16847);
and U20259 (N_20259,N_14267,N_14257);
nor U20260 (N_20260,N_13376,N_17077);
and U20261 (N_20261,N_17384,N_16855);
nor U20262 (N_20262,N_13126,N_14893);
xor U20263 (N_20263,N_16233,N_13165);
or U20264 (N_20264,N_14689,N_12813);
and U20265 (N_20265,N_17123,N_15504);
or U20266 (N_20266,N_15648,N_14477);
or U20267 (N_20267,N_16059,N_13727);
and U20268 (N_20268,N_14330,N_12931);
xor U20269 (N_20269,N_12472,N_17580);
nand U20270 (N_20270,N_12124,N_17331);
nor U20271 (N_20271,N_14288,N_14161);
and U20272 (N_20272,N_17519,N_13013);
or U20273 (N_20273,N_16427,N_14130);
and U20274 (N_20274,N_14271,N_12602);
nor U20275 (N_20275,N_14356,N_13614);
or U20276 (N_20276,N_16039,N_16778);
nor U20277 (N_20277,N_15165,N_12255);
xnor U20278 (N_20278,N_15918,N_16003);
nor U20279 (N_20279,N_16192,N_15070);
nor U20280 (N_20280,N_16589,N_16516);
xor U20281 (N_20281,N_13631,N_12491);
nand U20282 (N_20282,N_13145,N_17777);
xor U20283 (N_20283,N_17983,N_13337);
nor U20284 (N_20284,N_17626,N_16815);
and U20285 (N_20285,N_16286,N_16293);
or U20286 (N_20286,N_16042,N_12682);
nor U20287 (N_20287,N_16064,N_15505);
or U20288 (N_20288,N_16357,N_15831);
and U20289 (N_20289,N_15801,N_13449);
or U20290 (N_20290,N_15808,N_12902);
nand U20291 (N_20291,N_15660,N_12268);
nor U20292 (N_20292,N_17093,N_14748);
nand U20293 (N_20293,N_17883,N_13304);
xnor U20294 (N_20294,N_14375,N_14827);
nor U20295 (N_20295,N_17155,N_12957);
nand U20296 (N_20296,N_17132,N_17784);
nor U20297 (N_20297,N_12043,N_14055);
or U20298 (N_20298,N_12383,N_15090);
and U20299 (N_20299,N_12448,N_13599);
nor U20300 (N_20300,N_17252,N_14328);
xnor U20301 (N_20301,N_14520,N_15763);
nand U20302 (N_20302,N_13230,N_12893);
and U20303 (N_20303,N_13018,N_15104);
xnor U20304 (N_20304,N_13100,N_12738);
nand U20305 (N_20305,N_14036,N_14805);
xnor U20306 (N_20306,N_13779,N_14687);
xnor U20307 (N_20307,N_16151,N_14595);
and U20308 (N_20308,N_12446,N_13068);
nor U20309 (N_20309,N_12695,N_15785);
nor U20310 (N_20310,N_15002,N_12604);
nor U20311 (N_20311,N_13211,N_17442);
xnor U20312 (N_20312,N_13645,N_12982);
and U20313 (N_20313,N_15583,N_16612);
or U20314 (N_20314,N_13437,N_17181);
xor U20315 (N_20315,N_17223,N_12305);
or U20316 (N_20316,N_17191,N_16285);
nand U20317 (N_20317,N_12289,N_12719);
and U20318 (N_20318,N_13850,N_16415);
xor U20319 (N_20319,N_16554,N_17210);
and U20320 (N_20320,N_14165,N_16528);
or U20321 (N_20321,N_12063,N_15810);
nand U20322 (N_20322,N_15235,N_13925);
nor U20323 (N_20323,N_12230,N_13594);
xor U20324 (N_20324,N_15021,N_15271);
xnor U20325 (N_20325,N_12149,N_13793);
or U20326 (N_20326,N_13008,N_12229);
nand U20327 (N_20327,N_17686,N_15133);
nand U20328 (N_20328,N_16382,N_16069);
or U20329 (N_20329,N_15973,N_17441);
xnor U20330 (N_20330,N_15852,N_15950);
or U20331 (N_20331,N_15465,N_12443);
xor U20332 (N_20332,N_13769,N_15106);
xnor U20333 (N_20333,N_17887,N_16701);
nand U20334 (N_20334,N_13244,N_13729);
nand U20335 (N_20335,N_16461,N_12710);
or U20336 (N_20336,N_14322,N_16903);
nor U20337 (N_20337,N_14132,N_14289);
nand U20338 (N_20338,N_17890,N_16217);
nor U20339 (N_20339,N_16476,N_15064);
and U20340 (N_20340,N_15787,N_17385);
xnor U20341 (N_20341,N_12554,N_12985);
or U20342 (N_20342,N_12896,N_13591);
or U20343 (N_20343,N_13107,N_13933);
nand U20344 (N_20344,N_13654,N_12405);
or U20345 (N_20345,N_12074,N_13112);
nand U20346 (N_20346,N_15619,N_13794);
and U20347 (N_20347,N_17976,N_12717);
or U20348 (N_20348,N_13934,N_16440);
and U20349 (N_20349,N_12051,N_12788);
nor U20350 (N_20350,N_16416,N_12844);
or U20351 (N_20351,N_14746,N_14388);
or U20352 (N_20352,N_12762,N_17627);
nand U20353 (N_20353,N_16205,N_16507);
nand U20354 (N_20354,N_16765,N_15935);
nand U20355 (N_20355,N_15789,N_12406);
xor U20356 (N_20356,N_13856,N_13717);
or U20357 (N_20357,N_17917,N_14119);
xor U20358 (N_20358,N_12629,N_14550);
xnor U20359 (N_20359,N_12480,N_16727);
or U20360 (N_20360,N_16114,N_12358);
nand U20361 (N_20361,N_13718,N_12390);
or U20362 (N_20362,N_16068,N_17206);
or U20363 (N_20363,N_15431,N_13381);
or U20364 (N_20364,N_16629,N_13570);
or U20365 (N_20365,N_16340,N_17437);
nand U20366 (N_20366,N_14169,N_17709);
nor U20367 (N_20367,N_16893,N_15623);
xnor U20368 (N_20368,N_15072,N_16944);
nor U20369 (N_20369,N_17199,N_17833);
and U20370 (N_20370,N_17830,N_12177);
and U20371 (N_20371,N_13458,N_15585);
and U20372 (N_20372,N_13167,N_14572);
xnor U20373 (N_20373,N_12984,N_13043);
and U20374 (N_20374,N_14911,N_16965);
nand U20375 (N_20375,N_15994,N_12826);
and U20376 (N_20376,N_14862,N_17899);
xor U20377 (N_20377,N_16833,N_12224);
nand U20378 (N_20378,N_12087,N_14879);
or U20379 (N_20379,N_13121,N_16501);
nor U20380 (N_20380,N_13493,N_17453);
nand U20381 (N_20381,N_16635,N_15301);
xnor U20382 (N_20382,N_12527,N_12440);
nor U20383 (N_20383,N_12819,N_16062);
xnor U20384 (N_20384,N_17156,N_16805);
or U20385 (N_20385,N_16272,N_12786);
nor U20386 (N_20386,N_17762,N_16658);
nand U20387 (N_20387,N_15279,N_12487);
or U20388 (N_20388,N_15926,N_14832);
and U20389 (N_20389,N_12846,N_16266);
nor U20390 (N_20390,N_14639,N_17792);
and U20391 (N_20391,N_14401,N_16204);
xnor U20392 (N_20392,N_15441,N_16925);
nand U20393 (N_20393,N_17842,N_14648);
nand U20394 (N_20394,N_13030,N_16748);
xnor U20395 (N_20395,N_12062,N_14814);
nor U20396 (N_20396,N_17616,N_17408);
xnor U20397 (N_20397,N_16473,N_12129);
xor U20398 (N_20398,N_13519,N_15534);
and U20399 (N_20399,N_14726,N_17780);
and U20400 (N_20400,N_12636,N_12437);
and U20401 (N_20401,N_15014,N_16441);
xor U20402 (N_20402,N_17116,N_14611);
and U20403 (N_20403,N_16948,N_14162);
and U20404 (N_20404,N_15943,N_17746);
or U20405 (N_20405,N_15322,N_14997);
xor U20406 (N_20406,N_15020,N_12576);
xor U20407 (N_20407,N_14727,N_12669);
nand U20408 (N_20408,N_16195,N_15537);
nand U20409 (N_20409,N_14864,N_15044);
or U20410 (N_20410,N_15577,N_15033);
and U20411 (N_20411,N_17180,N_17651);
xor U20412 (N_20412,N_15496,N_17454);
nand U20413 (N_20413,N_13349,N_14230);
and U20414 (N_20414,N_12660,N_15443);
nor U20415 (N_20415,N_17955,N_17937);
xnor U20416 (N_20416,N_14347,N_17865);
or U20417 (N_20417,N_13318,N_17328);
nand U20418 (N_20418,N_14428,N_12779);
and U20419 (N_20419,N_16168,N_17377);
or U20420 (N_20420,N_12360,N_14084);
nor U20421 (N_20421,N_17756,N_16449);
and U20422 (N_20422,N_15039,N_17213);
and U20423 (N_20423,N_12901,N_13412);
or U20424 (N_20424,N_12653,N_14923);
nand U20425 (N_20425,N_15043,N_15083);
nand U20426 (N_20426,N_15359,N_16474);
or U20427 (N_20427,N_13721,N_17001);
or U20428 (N_20428,N_14088,N_17543);
xnor U20429 (N_20429,N_14779,N_14362);
and U20430 (N_20430,N_12867,N_13407);
or U20431 (N_20431,N_15611,N_14516);
and U20432 (N_20432,N_17827,N_17266);
nor U20433 (N_20433,N_14971,N_16160);
xor U20434 (N_20434,N_16691,N_16883);
or U20435 (N_20435,N_13696,N_16621);
or U20436 (N_20436,N_12032,N_17796);
or U20437 (N_20437,N_15157,N_13964);
nor U20438 (N_20438,N_16587,N_12250);
xor U20439 (N_20439,N_17470,N_17609);
and U20440 (N_20440,N_12295,N_16072);
or U20441 (N_20441,N_16367,N_12327);
and U20442 (N_20442,N_15168,N_16524);
xnor U20443 (N_20443,N_14946,N_16980);
or U20444 (N_20444,N_13397,N_16662);
and U20445 (N_20445,N_17823,N_16696);
or U20446 (N_20446,N_17508,N_17258);
nand U20447 (N_20447,N_14043,N_15839);
and U20448 (N_20448,N_14142,N_16532);
nor U20449 (N_20449,N_13451,N_13585);
xor U20450 (N_20450,N_14749,N_13281);
and U20451 (N_20451,N_12076,N_17783);
nor U20452 (N_20452,N_12831,N_13924);
or U20453 (N_20453,N_17695,N_17309);
xor U20454 (N_20454,N_16575,N_12216);
xor U20455 (N_20455,N_15703,N_15286);
nand U20456 (N_20456,N_12845,N_13636);
nand U20457 (N_20457,N_16436,N_15712);
xnor U20458 (N_20458,N_13555,N_15275);
and U20459 (N_20459,N_14087,N_12235);
nand U20460 (N_20460,N_16826,N_13403);
and U20461 (N_20461,N_14724,N_16311);
or U20462 (N_20462,N_12950,N_14313);
and U20463 (N_20463,N_15840,N_16424);
xnor U20464 (N_20464,N_12691,N_17957);
and U20465 (N_20465,N_15863,N_14485);
xor U20466 (N_20466,N_12506,N_17845);
or U20467 (N_20467,N_13590,N_13501);
or U20468 (N_20468,N_15719,N_12343);
and U20469 (N_20469,N_17550,N_13173);
and U20470 (N_20470,N_16921,N_17761);
xnor U20471 (N_20471,N_13986,N_16562);
xor U20472 (N_20472,N_17186,N_12505);
or U20473 (N_20473,N_15866,N_15188);
nand U20474 (N_20474,N_15621,N_12515);
xnor U20475 (N_20475,N_17689,N_12817);
nand U20476 (N_20476,N_17545,N_17510);
nor U20477 (N_20477,N_14061,N_13726);
xor U20478 (N_20478,N_13987,N_12521);
nand U20479 (N_20479,N_17136,N_17952);
and U20480 (N_20480,N_15997,N_16330);
or U20481 (N_20481,N_16718,N_13521);
and U20482 (N_20482,N_16602,N_16385);
xnor U20483 (N_20483,N_16750,N_13341);
nand U20484 (N_20484,N_13336,N_17577);
nor U20485 (N_20485,N_17065,N_14424);
xnor U20486 (N_20486,N_13686,N_15975);
xnor U20487 (N_20487,N_17666,N_14708);
or U20488 (N_20488,N_15735,N_13400);
and U20489 (N_20489,N_16842,N_14108);
nor U20490 (N_20490,N_16857,N_17055);
nand U20491 (N_20491,N_14976,N_14554);
xnor U20492 (N_20492,N_16442,N_13345);
and U20493 (N_20493,N_16605,N_14788);
xor U20494 (N_20494,N_12862,N_16110);
and U20495 (N_20495,N_15876,N_16609);
nand U20496 (N_20496,N_16625,N_17670);
or U20497 (N_20497,N_14478,N_17862);
xor U20498 (N_20498,N_17179,N_16140);
nor U20499 (N_20499,N_12589,N_16302);
nor U20500 (N_20500,N_13063,N_17129);
nand U20501 (N_20501,N_15038,N_16263);
xnor U20502 (N_20502,N_13426,N_14014);
xnor U20503 (N_20503,N_16394,N_15058);
or U20504 (N_20504,N_12461,N_15654);
nand U20505 (N_20505,N_13226,N_17544);
and U20506 (N_20506,N_14912,N_13754);
nor U20507 (N_20507,N_12337,N_15252);
nand U20508 (N_20508,N_14536,N_15641);
nor U20509 (N_20509,N_16027,N_13302);
or U20510 (N_20510,N_14285,N_14840);
and U20511 (N_20511,N_16910,N_16188);
nand U20512 (N_20512,N_14008,N_16322);
and U20513 (N_20513,N_13078,N_16162);
nand U20514 (N_20514,N_13919,N_12757);
nand U20515 (N_20515,N_13436,N_12333);
nor U20516 (N_20516,N_15579,N_13253);
xnor U20517 (N_20517,N_15341,N_14562);
xnor U20518 (N_20518,N_15779,N_16681);
or U20519 (N_20519,N_17410,N_16933);
nor U20520 (N_20520,N_14947,N_14022);
xor U20521 (N_20521,N_12111,N_17766);
or U20522 (N_20522,N_16558,N_17944);
and U20523 (N_20523,N_12776,N_12442);
xnor U20524 (N_20524,N_13516,N_13228);
nand U20525 (N_20525,N_17821,N_14945);
nand U20526 (N_20526,N_14106,N_14691);
or U20527 (N_20527,N_12578,N_12017);
xnor U20528 (N_20528,N_15931,N_15493);
or U20529 (N_20529,N_13787,N_12808);
xor U20530 (N_20530,N_12001,N_15227);
nor U20531 (N_20531,N_13959,N_15290);
nand U20532 (N_20532,N_12694,N_15125);
nand U20533 (N_20533,N_17291,N_12658);
and U20534 (N_20534,N_14733,N_14624);
nor U20535 (N_20535,N_16985,N_13139);
or U20536 (N_20536,N_17878,N_15454);
nand U20537 (N_20537,N_16453,N_13994);
nand U20538 (N_20538,N_15233,N_15167);
and U20539 (N_20539,N_15812,N_14353);
or U20540 (N_20540,N_17734,N_17884);
and U20541 (N_20541,N_13404,N_12909);
xnor U20542 (N_20542,N_14261,N_13279);
or U20543 (N_20543,N_16244,N_13300);
and U20544 (N_20544,N_17147,N_16711);
nand U20545 (N_20545,N_15754,N_14710);
nor U20546 (N_20546,N_13160,N_17868);
xnor U20547 (N_20547,N_13446,N_17718);
and U20548 (N_20548,N_16694,N_15751);
or U20549 (N_20549,N_13330,N_13939);
or U20550 (N_20550,N_14583,N_17463);
xnor U20551 (N_20551,N_15574,N_13503);
or U20552 (N_20552,N_12130,N_13682);
and U20553 (N_20553,N_13232,N_14363);
nor U20554 (N_20554,N_15945,N_14141);
or U20555 (N_20555,N_15270,N_12156);
or U20556 (N_20556,N_16757,N_16611);
nor U20557 (N_20557,N_14504,N_16087);
xor U20558 (N_20558,N_13114,N_17828);
nand U20559 (N_20559,N_16817,N_13708);
nor U20560 (N_20560,N_14929,N_15546);
nor U20561 (N_20561,N_12261,N_14158);
and U20562 (N_20562,N_15485,N_12158);
nor U20563 (N_20563,N_15091,N_14116);
nand U20564 (N_20564,N_16776,N_17892);
nor U20565 (N_20565,N_17954,N_12114);
xnor U20566 (N_20566,N_17015,N_12587);
xnor U20567 (N_20567,N_12414,N_14157);
nor U20568 (N_20568,N_14366,N_12550);
and U20569 (N_20569,N_12029,N_16471);
nor U20570 (N_20570,N_15255,N_14168);
nand U20571 (N_20571,N_16584,N_13081);
nor U20572 (N_20572,N_13477,N_14082);
and U20573 (N_20573,N_15879,N_13497);
xor U20574 (N_20574,N_15113,N_12085);
nand U20575 (N_20575,N_17755,N_14909);
or U20576 (N_20576,N_16889,N_17423);
xnor U20577 (N_20577,N_15667,N_16075);
and U20578 (N_20578,N_14990,N_14626);
xnor U20579 (N_20579,N_12508,N_17643);
xnor U20580 (N_20580,N_17122,N_14847);
xnor U20581 (N_20581,N_12520,N_15500);
and U20582 (N_20582,N_16224,N_14384);
xor U20583 (N_20583,N_13262,N_16421);
or U20584 (N_20584,N_15360,N_15759);
xnor U20585 (N_20585,N_15369,N_15258);
or U20586 (N_20586,N_15832,N_12748);
nor U20587 (N_20587,N_17143,N_12199);
nand U20588 (N_20588,N_15076,N_15770);
nor U20589 (N_20589,N_14448,N_12420);
or U20590 (N_20590,N_17458,N_14534);
or U20591 (N_20591,N_13869,N_17632);
nor U20592 (N_20592,N_14327,N_14234);
nand U20593 (N_20593,N_13465,N_17096);
and U20594 (N_20594,N_12714,N_17505);
nor U20595 (N_20595,N_12256,N_12999);
nand U20596 (N_20596,N_14056,N_14489);
nand U20597 (N_20597,N_13200,N_15655);
xnor U20598 (N_20598,N_13007,N_17357);
nor U20599 (N_20599,N_15394,N_16187);
nor U20600 (N_20600,N_15669,N_17700);
and U20601 (N_20601,N_15612,N_15119);
and U20602 (N_20602,N_12606,N_16510);
nor U20603 (N_20603,N_13949,N_15791);
or U20604 (N_20604,N_13212,N_15438);
nor U20605 (N_20605,N_15664,N_13935);
xnor U20606 (N_20606,N_15847,N_14020);
xnor U20607 (N_20607,N_15284,N_17546);
and U20608 (N_20608,N_17674,N_15491);
or U20609 (N_20609,N_16770,N_12884);
or U20610 (N_20610,N_15389,N_17566);
and U20611 (N_20611,N_15818,N_12922);
and U20612 (N_20612,N_16520,N_13441);
or U20613 (N_20613,N_12190,N_17069);
and U20614 (N_20614,N_13748,N_15692);
and U20615 (N_20615,N_12939,N_14622);
or U20616 (N_20616,N_14694,N_13231);
nand U20617 (N_20617,N_13659,N_15541);
xor U20618 (N_20618,N_12608,N_12025);
xnor U20619 (N_20619,N_14922,N_12827);
xor U20620 (N_20620,N_17051,N_15632);
nand U20621 (N_20621,N_15412,N_13604);
or U20622 (N_20622,N_13475,N_17235);
nand U20623 (N_20623,N_17771,N_16354);
nand U20624 (N_20624,N_15609,N_17220);
nor U20625 (N_20625,N_16538,N_16561);
nor U20626 (N_20626,N_16077,N_16989);
xor U20627 (N_20627,N_13839,N_13607);
or U20628 (N_20628,N_16827,N_16604);
and U20629 (N_20629,N_17614,N_17488);
nor U20630 (N_20630,N_16060,N_15409);
and U20631 (N_20631,N_15513,N_17204);
xor U20632 (N_20632,N_12095,N_13271);
nand U20633 (N_20633,N_13638,N_14638);
xnor U20634 (N_20634,N_13792,N_15145);
xnor U20635 (N_20635,N_15383,N_12252);
xnor U20636 (N_20636,N_16444,N_14587);
nor U20637 (N_20637,N_12696,N_16196);
nand U20638 (N_20638,N_15311,N_16115);
and U20639 (N_20639,N_12994,N_16872);
nand U20640 (N_20640,N_17493,N_17719);
xor U20641 (N_20641,N_13301,N_13448);
nor U20642 (N_20642,N_17708,N_17811);
or U20643 (N_20643,N_16365,N_13881);
nand U20644 (N_20644,N_17398,N_13101);
nor U20645 (N_20645,N_14174,N_15949);
nor U20646 (N_20646,N_12410,N_17953);
nor U20647 (N_20647,N_14538,N_14655);
nor U20648 (N_20648,N_14344,N_12923);
and U20649 (N_20649,N_12670,N_16463);
and U20650 (N_20650,N_12453,N_12315);
xnor U20651 (N_20651,N_12585,N_16175);
or U20652 (N_20652,N_17728,N_16054);
xor U20653 (N_20653,N_13612,N_14975);
nor U20654 (N_20654,N_13755,N_13325);
nor U20655 (N_20655,N_13745,N_16814);
or U20656 (N_20656,N_16128,N_14259);
nand U20657 (N_20657,N_13532,N_12942);
and U20658 (N_20658,N_14980,N_17706);
or U20659 (N_20659,N_17721,N_15603);
or U20660 (N_20660,N_12112,N_16023);
and U20661 (N_20661,N_15231,N_14219);
xnor U20662 (N_20662,N_17110,N_13658);
nor U20663 (N_20663,N_12242,N_17087);
or U20664 (N_20664,N_15011,N_14619);
nand U20665 (N_20665,N_17662,N_13453);
and U20666 (N_20666,N_13246,N_17436);
or U20667 (N_20667,N_14373,N_15048);
nor U20668 (N_20668,N_16529,N_17062);
or U20669 (N_20669,N_17020,N_12054);
nor U20670 (N_20670,N_15074,N_13106);
nor U20671 (N_20671,N_15298,N_15335);
and U20672 (N_20672,N_16320,N_13897);
xnor U20673 (N_20673,N_12564,N_15928);
xnor U20674 (N_20674,N_16211,N_13137);
or U20675 (N_20675,N_12530,N_16369);
nand U20676 (N_20676,N_17971,N_17088);
and U20677 (N_20677,N_16927,N_14156);
nor U20678 (N_20678,N_17234,N_15292);
and U20679 (N_20679,N_17946,N_13316);
nor U20680 (N_20680,N_15862,N_13921);
and U20681 (N_20681,N_14374,N_16333);
and U20682 (N_20682,N_12325,N_12324);
and U20683 (N_20683,N_14256,N_14625);
and U20684 (N_20684,N_17208,N_12990);
or U20685 (N_20685,N_12039,N_15610);
and U20686 (N_20686,N_16227,N_17832);
nand U20687 (N_20687,N_13378,N_14390);
or U20688 (N_20688,N_15202,N_17677);
nor U20689 (N_20689,N_14146,N_17124);
xnor U20690 (N_20690,N_12094,N_16250);
or U20691 (N_20691,N_13125,N_15268);
and U20692 (N_20692,N_14274,N_12166);
nor U20693 (N_20693,N_15244,N_12195);
and U20694 (N_20694,N_17347,N_14663);
or U20695 (N_20695,N_12429,N_16397);
or U20696 (N_20696,N_12301,N_12260);
xnor U20697 (N_20697,N_13799,N_12740);
nand U20698 (N_20698,N_12547,N_15804);
xor U20699 (N_20699,N_16347,N_17947);
xnor U20700 (N_20700,N_12665,N_16630);
and U20701 (N_20701,N_14880,N_17287);
and U20702 (N_20702,N_12915,N_13129);
or U20703 (N_20703,N_13042,N_16517);
nand U20704 (N_20704,N_12617,N_13016);
nand U20705 (N_20705,N_13728,N_12848);
nand U20706 (N_20706,N_15263,N_17769);
and U20707 (N_20707,N_14247,N_15498);
and U20708 (N_20708,N_14962,N_15399);
or U20709 (N_20709,N_15323,N_17867);
or U20710 (N_20710,N_16810,N_14443);
and U20711 (N_20711,N_14505,N_16157);
nor U20712 (N_20712,N_13932,N_13036);
or U20713 (N_20713,N_17768,N_13111);
xor U20714 (N_20714,N_14918,N_14631);
xnor U20715 (N_20715,N_12821,N_15305);
or U20716 (N_20716,N_17153,N_16905);
or U20717 (N_20717,N_14618,N_17316);
nand U20718 (N_20718,N_12921,N_14507);
xnor U20719 (N_20719,N_12263,N_15230);
nor U20720 (N_20720,N_16014,N_17949);
nor U20721 (N_20721,N_15078,N_16076);
nor U20722 (N_20722,N_13610,N_13635);
nand U20723 (N_20723,N_14154,N_14711);
nor U20724 (N_20724,N_12228,N_13780);
nand U20725 (N_20725,N_16353,N_17244);
xnor U20726 (N_20726,N_16101,N_17939);
nor U20727 (N_20727,N_13912,N_13122);
nand U20728 (N_20728,N_14594,N_12163);
nor U20729 (N_20729,N_13757,N_13820);
nor U20730 (N_20730,N_17054,N_15701);
or U20731 (N_20731,N_17779,N_13844);
xnor U20732 (N_20732,N_13697,N_16945);
or U20733 (N_20733,N_15102,N_12306);
xor U20734 (N_20734,N_16373,N_16052);
and U20735 (N_20735,N_17150,N_16940);
xor U20736 (N_20736,N_16616,N_16491);
and U20737 (N_20737,N_17789,N_13187);
nor U20738 (N_20738,N_13243,N_13024);
or U20739 (N_20739,N_15184,N_17804);
and U20740 (N_20740,N_15150,N_14873);
nand U20741 (N_20741,N_15806,N_16722);
nor U20742 (N_20742,N_12588,N_16212);
nand U20743 (N_20743,N_15616,N_13997);
xor U20744 (N_20744,N_14759,N_15953);
nor U20745 (N_20745,N_17653,N_13156);
xor U20746 (N_20746,N_15089,N_12992);
xnor U20747 (N_20747,N_17162,N_17807);
nand U20748 (N_20748,N_12178,N_13456);
nor U20749 (N_20749,N_14709,N_14988);
or U20750 (N_20750,N_17475,N_12084);
xor U20751 (N_20751,N_13227,N_16684);
and U20752 (N_20752,N_16861,N_16555);
or U20753 (N_20753,N_17217,N_17298);
nand U20754 (N_20754,N_15511,N_14039);
or U20755 (N_20755,N_12668,N_12876);
and U20756 (N_20756,N_16438,N_15677);
or U20757 (N_20757,N_16798,N_17468);
nand U20758 (N_20758,N_13973,N_15662);
nand U20759 (N_20759,N_16074,N_12969);
nor U20760 (N_20760,N_13968,N_15016);
and U20761 (N_20761,N_17682,N_14213);
or U20762 (N_20762,N_17560,N_15319);
nand U20763 (N_20763,N_16640,N_16716);
or U20764 (N_20764,N_13136,N_15749);
nor U20765 (N_20765,N_16699,N_15332);
or U20766 (N_20766,N_14580,N_13360);
nor U20767 (N_20767,N_14083,N_15638);
or U20768 (N_20768,N_16057,N_12419);
nand U20769 (N_20769,N_12533,N_17342);
and U20770 (N_20770,N_13976,N_12474);
or U20771 (N_20771,N_15993,N_12770);
xor U20772 (N_20772,N_16464,N_14081);
or U20773 (N_20773,N_13411,N_13966);
and U20774 (N_20774,N_14490,N_16887);
and U20775 (N_20775,N_16597,N_16966);
xnor U20776 (N_20776,N_16225,N_14792);
nor U20777 (N_20777,N_12967,N_14498);
xnor U20778 (N_20778,N_15447,N_14229);
or U20779 (N_20779,N_14250,N_16337);
or U20780 (N_20780,N_12059,N_13522);
and U20781 (N_20781,N_13425,N_13194);
xnor U20782 (N_20782,N_17741,N_15453);
or U20783 (N_20783,N_15726,N_17797);
nand U20784 (N_20784,N_14803,N_13665);
or U20785 (N_20785,N_17603,N_13541);
or U20786 (N_20786,N_16978,N_15837);
and U20787 (N_20787,N_12607,N_15459);
and U20788 (N_20788,N_15274,N_15209);
nor U20789 (N_20789,N_14705,N_16121);
xor U20790 (N_20790,N_12011,N_14201);
xnor U20791 (N_20791,N_17194,N_14017);
nor U20792 (N_20792,N_13029,N_12003);
nor U20793 (N_20793,N_16153,N_15998);
nand U20794 (N_20794,N_16901,N_14199);
and U20795 (N_20795,N_16260,N_12254);
and U20796 (N_20796,N_13841,N_13569);
nor U20797 (N_20797,N_14143,N_13720);
xnor U20798 (N_20798,N_17296,N_12591);
xnor U20799 (N_20799,N_16987,N_16256);
xor U20800 (N_20800,N_12581,N_15297);
xor U20801 (N_20801,N_16133,N_13705);
and U20802 (N_20802,N_12009,N_13693);
or U20803 (N_20803,N_12106,N_16466);
xor U20804 (N_20804,N_13208,N_13835);
nor U20805 (N_20805,N_13694,N_17343);
xor U20806 (N_20806,N_16705,N_16408);
nor U20807 (N_20807,N_15003,N_12381);
or U20808 (N_20808,N_16089,N_17052);
and U20809 (N_20809,N_12616,N_17585);
or U20810 (N_20810,N_17554,N_16729);
xnor U20811 (N_20811,N_16679,N_13542);
xor U20812 (N_20812,N_17163,N_14761);
xnor U20813 (N_20813,N_17341,N_15046);
and U20814 (N_20814,N_15764,N_16742);
and U20815 (N_20815,N_13534,N_12689);
and U20816 (N_20816,N_13348,N_15925);
or U20817 (N_20817,N_17336,N_14526);
and U20818 (N_20818,N_15066,N_15261);
nand U20819 (N_20819,N_12212,N_12165);
xnor U20820 (N_20820,N_14475,N_14420);
nand U20821 (N_20821,N_15315,N_14718);
or U20822 (N_20822,N_17031,N_14361);
nand U20823 (N_20823,N_12634,N_15584);
nor U20824 (N_20824,N_17435,N_16257);
or U20825 (N_20825,N_17202,N_13602);
and U20826 (N_20826,N_16671,N_13508);
nand U20827 (N_20827,N_16078,N_17146);
nand U20828 (N_20828,N_15736,N_16419);
nand U20829 (N_20829,N_17466,N_17100);
nor U20830 (N_20830,N_16318,N_15015);
xor U20831 (N_20831,N_13797,N_12953);
xor U20832 (N_20832,N_13182,N_13443);
xnor U20833 (N_20833,N_16774,N_14921);
and U20834 (N_20834,N_17857,N_15265);
or U20835 (N_20835,N_13977,N_15578);
xor U20836 (N_20836,N_13191,N_14031);
and U20837 (N_20837,N_12615,N_15758);
nor U20838 (N_20838,N_16566,N_13309);
nand U20839 (N_20839,N_12047,N_13510);
or U20840 (N_20840,N_16552,N_17212);
nand U20841 (N_20841,N_13017,N_14226);
or U20842 (N_20842,N_14272,N_14910);
nor U20843 (N_20843,N_16870,N_17401);
nor U20844 (N_20844,N_15668,N_13871);
and U20845 (N_20845,N_17205,N_12523);
xor U20846 (N_20846,N_13354,N_13783);
or U20847 (N_20847,N_16526,N_16001);
or U20848 (N_20848,N_13217,N_17371);
nand U20849 (N_20849,N_13409,N_15309);
nor U20850 (N_20850,N_14699,N_15050);
and U20851 (N_20851,N_12655,N_17456);
or U20852 (N_20852,N_15752,N_15122);
and U20853 (N_20853,N_12652,N_17753);
xor U20854 (N_20854,N_17654,N_15034);
nand U20855 (N_20855,N_14451,N_15988);
and U20856 (N_20856,N_17961,N_15970);
nand U20857 (N_20857,N_15313,N_13151);
nor U20858 (N_20858,N_12467,N_13567);
and U20859 (N_20859,N_15088,N_15196);
or U20860 (N_20860,N_17233,N_12099);
nor U20861 (N_20861,N_14981,N_14902);
nor U20862 (N_20862,N_14469,N_16182);
xor U20863 (N_20863,N_14416,N_16533);
xor U20864 (N_20864,N_16816,N_12117);
xor U20865 (N_20865,N_17572,N_15492);
and U20866 (N_20866,N_13393,N_17302);
or U20867 (N_20867,N_15991,N_14900);
or U20868 (N_20868,N_17969,N_12091);
nand U20869 (N_20869,N_15666,N_14482);
nand U20870 (N_20870,N_15556,N_13143);
and U20871 (N_20871,N_13800,N_13758);
and U20872 (N_20872,N_16841,N_13141);
nor U20873 (N_20873,N_17819,N_13054);
and U20874 (N_20874,N_16606,N_12193);
and U20875 (N_20875,N_17634,N_16316);
and U20876 (N_20876,N_14419,N_16638);
or U20877 (N_20877,N_12692,N_13479);
nand U20878 (N_20878,N_12561,N_12019);
and U20879 (N_20879,N_17675,N_14155);
and U20880 (N_20880,N_12126,N_12855);
nor U20881 (N_20881,N_13385,N_14164);
and U20882 (N_20882,N_15220,N_17038);
nand U20883 (N_20883,N_12600,N_12144);
nor U20884 (N_20884,N_14379,N_16376);
and U20885 (N_20885,N_14558,N_16107);
xnor U20886 (N_20886,N_16249,N_16144);
and U20887 (N_20887,N_15514,N_15092);
nor U20888 (N_20888,N_14901,N_13574);
and U20889 (N_20889,N_15956,N_12742);
or U20890 (N_20890,N_16622,N_13415);
or U20891 (N_20891,N_16646,N_13002);
or U20892 (N_20892,N_12593,N_12274);
and U20893 (N_20893,N_12338,N_13113);
nand U20894 (N_20894,N_13097,N_14246);
xnor U20895 (N_20895,N_13891,N_17125);
nor U20896 (N_20896,N_16521,N_12456);
xnor U20897 (N_20897,N_14204,N_13201);
nand U20898 (N_20898,N_14790,N_14460);
and U20899 (N_20899,N_17948,N_12220);
and U20900 (N_20900,N_15591,N_16190);
nand U20901 (N_20901,N_17455,N_13647);
or U20902 (N_20902,N_12171,N_13807);
xnor U20903 (N_20903,N_15232,N_17360);
xnor U20904 (N_20904,N_14835,N_14830);
xnor U20905 (N_20905,N_12353,N_14368);
xor U20906 (N_20906,N_17669,N_12545);
nor U20907 (N_20907,N_15778,N_15890);
or U20908 (N_20908,N_17119,N_12203);
or U20909 (N_20909,N_15526,N_13306);
xnor U20910 (N_20910,N_14744,N_15733);
nand U20911 (N_20911,N_15144,N_17400);
and U20912 (N_20912,N_12540,N_17642);
nor U20913 (N_20913,N_12745,N_17999);
nor U20914 (N_20914,N_14763,N_14608);
or U20915 (N_20915,N_15561,N_16848);
and U20916 (N_20916,N_14198,N_14438);
or U20917 (N_20917,N_14282,N_17902);
xor U20918 (N_20918,N_13175,N_13646);
nor U20919 (N_20919,N_12721,N_15191);
and U20920 (N_20920,N_14153,N_12198);
and U20921 (N_20921,N_14408,N_14391);
and U20922 (N_20922,N_17236,N_12484);
and U20923 (N_20923,N_17496,N_16919);
xor U20924 (N_20924,N_16081,N_12335);
nand U20925 (N_20925,N_14397,N_12764);
or U20926 (N_20926,N_13902,N_14863);
or U20927 (N_20927,N_15741,N_13789);
nor U20928 (N_20928,N_13957,N_17280);
nor U20929 (N_20929,N_16665,N_17394);
or U20930 (N_20930,N_13000,N_12403);
and U20931 (N_20931,N_13657,N_15586);
or U20932 (N_20932,N_16010,N_12080);
and U20933 (N_20933,N_15460,N_12477);
nor U20934 (N_20934,N_12642,N_16586);
and U20935 (N_20935,N_12399,N_12226);
and U20936 (N_20936,N_12122,N_12584);
xor U20937 (N_20937,N_17848,N_15671);
xnor U20938 (N_20938,N_14354,N_12145);
nand U20939 (N_20939,N_13286,N_16470);
xnor U20940 (N_20940,N_17579,N_15299);
nand U20941 (N_20941,N_14821,N_17157);
or U20942 (N_20942,N_14455,N_16084);
nor U20943 (N_20943,N_14784,N_15672);
nor U20944 (N_20944,N_13083,N_16259);
xor U20945 (N_20945,N_17765,N_16500);
and U20946 (N_20946,N_14134,N_15354);
nor U20947 (N_20947,N_12900,N_12628);
nor U20948 (N_20948,N_13621,N_15728);
or U20949 (N_20949,N_15595,N_17533);
and U20950 (N_20950,N_17965,N_17526);
xor U20951 (N_20951,N_14607,N_16650);
nand U20952 (N_20952,N_15553,N_13494);
nand U20953 (N_20953,N_12516,N_15217);
or U20954 (N_20954,N_16275,N_12310);
or U20955 (N_20955,N_14957,N_15344);
and U20956 (N_20956,N_15100,N_17825);
or U20957 (N_20957,N_17988,N_12534);
nand U20958 (N_20958,N_13197,N_15506);
and U20959 (N_20959,N_13422,N_12980);
and U20960 (N_20960,N_16577,N_12016);
xnor U20961 (N_20961,N_16836,N_12575);
nor U20962 (N_20962,N_17165,N_15065);
nor U20963 (N_20963,N_12439,N_17393);
nand U20964 (N_20964,N_15649,N_15686);
or U20965 (N_20965,N_17406,N_17327);
xnor U20966 (N_20966,N_13109,N_12247);
xnor U20967 (N_20967,N_17688,N_15198);
and U20968 (N_20968,N_16957,N_17379);
xor U20969 (N_20969,N_16163,N_14094);
or U20970 (N_20970,N_15172,N_16154);
nor U20971 (N_20971,N_13583,N_12218);
or U20972 (N_20972,N_17919,N_14566);
xor U20973 (N_20973,N_17375,N_13983);
nor U20974 (N_20974,N_12164,N_12995);
and U20975 (N_20975,N_12754,N_15178);
xnor U20976 (N_20976,N_14402,N_17151);
nand U20977 (N_20977,N_12858,N_17469);
xnor U20978 (N_20978,N_16136,N_17860);
xnor U20979 (N_20979,N_12359,N_15494);
nand U20980 (N_20980,N_14421,N_17271);
nor U20981 (N_20981,N_13832,N_16961);
nand U20982 (N_20982,N_12873,N_14644);
xnor U20983 (N_20983,N_12168,N_14238);
nand U20984 (N_20984,N_16455,N_14842);
and U20985 (N_20985,N_15458,N_15501);
or U20986 (N_20986,N_15854,N_13670);
nor U20987 (N_20987,N_17427,N_12148);
xor U20988 (N_20988,N_16818,N_16585);
nand U20989 (N_20989,N_17424,N_15080);
nor U20990 (N_20990,N_14928,N_12849);
or U20991 (N_20991,N_14768,N_14078);
nand U20992 (N_20992,N_13892,N_12370);
nor U20993 (N_20993,N_14190,N_14854);
xnor U20994 (N_20994,N_17443,N_14555);
xor U20995 (N_20995,N_14810,N_16452);
and U20996 (N_20996,N_14890,N_12021);
nor U20997 (N_20997,N_16786,N_13860);
nand U20998 (N_20998,N_15944,N_13969);
and U20999 (N_20999,N_12801,N_15755);
nor U21000 (N_21000,N_17670,N_16325);
or U21001 (N_21001,N_12297,N_13898);
nand U21002 (N_21002,N_16909,N_14078);
and U21003 (N_21003,N_15825,N_13152);
and U21004 (N_21004,N_16075,N_13717);
or U21005 (N_21005,N_16954,N_14157);
or U21006 (N_21006,N_17334,N_17273);
or U21007 (N_21007,N_14434,N_16078);
nand U21008 (N_21008,N_16979,N_15864);
nor U21009 (N_21009,N_13268,N_14010);
nor U21010 (N_21010,N_17060,N_15148);
nand U21011 (N_21011,N_17375,N_12459);
nand U21012 (N_21012,N_12173,N_13130);
xnor U21013 (N_21013,N_14496,N_15660);
nand U21014 (N_21014,N_13049,N_16451);
nand U21015 (N_21015,N_12908,N_14575);
or U21016 (N_21016,N_17624,N_15131);
and U21017 (N_21017,N_15493,N_15913);
nand U21018 (N_21018,N_13888,N_16644);
xor U21019 (N_21019,N_13298,N_17107);
nor U21020 (N_21020,N_12642,N_16425);
xor U21021 (N_21021,N_12711,N_17078);
nor U21022 (N_21022,N_16181,N_15690);
or U21023 (N_21023,N_17541,N_15899);
or U21024 (N_21024,N_15086,N_16444);
xnor U21025 (N_21025,N_15905,N_12285);
nand U21026 (N_21026,N_12206,N_17948);
or U21027 (N_21027,N_14224,N_13474);
nor U21028 (N_21028,N_14438,N_12552);
or U21029 (N_21029,N_16655,N_14047);
and U21030 (N_21030,N_17762,N_15804);
and U21031 (N_21031,N_17667,N_15504);
nand U21032 (N_21032,N_14187,N_16663);
nor U21033 (N_21033,N_16952,N_15790);
nand U21034 (N_21034,N_12313,N_16554);
nand U21035 (N_21035,N_16410,N_12752);
nor U21036 (N_21036,N_13051,N_13589);
nand U21037 (N_21037,N_12202,N_16353);
nor U21038 (N_21038,N_14505,N_13282);
nor U21039 (N_21039,N_17703,N_12947);
xnor U21040 (N_21040,N_16490,N_13877);
xnor U21041 (N_21041,N_17500,N_14775);
xnor U21042 (N_21042,N_14967,N_13841);
xor U21043 (N_21043,N_17601,N_16293);
xnor U21044 (N_21044,N_14617,N_16907);
nand U21045 (N_21045,N_14194,N_16289);
nor U21046 (N_21046,N_16732,N_12904);
nand U21047 (N_21047,N_13394,N_13321);
or U21048 (N_21048,N_17145,N_13192);
and U21049 (N_21049,N_13732,N_15715);
or U21050 (N_21050,N_14112,N_15416);
xnor U21051 (N_21051,N_16954,N_15486);
xnor U21052 (N_21052,N_14424,N_15673);
and U21053 (N_21053,N_17036,N_12705);
or U21054 (N_21054,N_15879,N_13901);
xor U21055 (N_21055,N_17175,N_15819);
nand U21056 (N_21056,N_17215,N_15983);
nor U21057 (N_21057,N_17255,N_14734);
xnor U21058 (N_21058,N_12220,N_15587);
and U21059 (N_21059,N_17574,N_13114);
nor U21060 (N_21060,N_17950,N_13956);
or U21061 (N_21061,N_13646,N_13933);
xor U21062 (N_21062,N_17110,N_12374);
nor U21063 (N_21063,N_15588,N_14504);
xor U21064 (N_21064,N_16277,N_15610);
and U21065 (N_21065,N_13473,N_15340);
nand U21066 (N_21066,N_17483,N_15415);
and U21067 (N_21067,N_17538,N_17622);
xnor U21068 (N_21068,N_16624,N_14681);
nor U21069 (N_21069,N_17249,N_15998);
or U21070 (N_21070,N_12091,N_14093);
or U21071 (N_21071,N_16191,N_17390);
nor U21072 (N_21072,N_13063,N_17006);
nand U21073 (N_21073,N_13103,N_15625);
xnor U21074 (N_21074,N_13440,N_12925);
and U21075 (N_21075,N_17189,N_17332);
nand U21076 (N_21076,N_16950,N_17522);
nand U21077 (N_21077,N_12545,N_12541);
and U21078 (N_21078,N_14443,N_12900);
nand U21079 (N_21079,N_15739,N_17639);
nand U21080 (N_21080,N_14230,N_16018);
and U21081 (N_21081,N_13054,N_13096);
nor U21082 (N_21082,N_16108,N_12833);
nand U21083 (N_21083,N_15080,N_12836);
and U21084 (N_21084,N_14721,N_12633);
or U21085 (N_21085,N_13194,N_15511);
nand U21086 (N_21086,N_16003,N_17119);
and U21087 (N_21087,N_14759,N_14728);
and U21088 (N_21088,N_14561,N_16222);
nor U21089 (N_21089,N_16058,N_16762);
or U21090 (N_21090,N_15757,N_14775);
nor U21091 (N_21091,N_15717,N_13197);
nand U21092 (N_21092,N_14050,N_15516);
nor U21093 (N_21093,N_14757,N_17852);
xnor U21094 (N_21094,N_16761,N_12777);
nand U21095 (N_21095,N_16565,N_14906);
nor U21096 (N_21096,N_16400,N_16709);
xor U21097 (N_21097,N_15945,N_16122);
and U21098 (N_21098,N_16660,N_16390);
xor U21099 (N_21099,N_14518,N_13065);
or U21100 (N_21100,N_17481,N_13256);
nor U21101 (N_21101,N_12140,N_13316);
or U21102 (N_21102,N_15589,N_13750);
nand U21103 (N_21103,N_12305,N_16631);
nand U21104 (N_21104,N_13068,N_12601);
nand U21105 (N_21105,N_15607,N_14795);
xnor U21106 (N_21106,N_15244,N_15631);
nor U21107 (N_21107,N_12636,N_12074);
and U21108 (N_21108,N_13295,N_12131);
nand U21109 (N_21109,N_13753,N_13847);
nor U21110 (N_21110,N_16598,N_12789);
nor U21111 (N_21111,N_15724,N_12254);
nand U21112 (N_21112,N_12517,N_17010);
nand U21113 (N_21113,N_15061,N_12763);
or U21114 (N_21114,N_16417,N_15208);
or U21115 (N_21115,N_12925,N_16136);
and U21116 (N_21116,N_12760,N_12113);
nand U21117 (N_21117,N_14760,N_13472);
and U21118 (N_21118,N_13888,N_17404);
or U21119 (N_21119,N_16686,N_12828);
nor U21120 (N_21120,N_17679,N_16761);
and U21121 (N_21121,N_12010,N_13730);
nor U21122 (N_21122,N_13639,N_15170);
xnor U21123 (N_21123,N_13372,N_15771);
xor U21124 (N_21124,N_16510,N_15490);
or U21125 (N_21125,N_16656,N_14981);
nor U21126 (N_21126,N_12830,N_12925);
xnor U21127 (N_21127,N_16014,N_13476);
nor U21128 (N_21128,N_13290,N_14895);
xor U21129 (N_21129,N_13460,N_15966);
nand U21130 (N_21130,N_16506,N_16899);
nand U21131 (N_21131,N_14111,N_12301);
and U21132 (N_21132,N_17325,N_17274);
or U21133 (N_21133,N_13453,N_16594);
nand U21134 (N_21134,N_17492,N_12754);
nor U21135 (N_21135,N_14906,N_15391);
or U21136 (N_21136,N_12991,N_14120);
or U21137 (N_21137,N_12534,N_13778);
nor U21138 (N_21138,N_14806,N_12446);
or U21139 (N_21139,N_15761,N_16534);
nor U21140 (N_21140,N_13678,N_15397);
xor U21141 (N_21141,N_14445,N_14274);
xor U21142 (N_21142,N_13541,N_14668);
xnor U21143 (N_21143,N_12185,N_14311);
or U21144 (N_21144,N_16487,N_17098);
or U21145 (N_21145,N_16053,N_12274);
and U21146 (N_21146,N_12563,N_17901);
or U21147 (N_21147,N_15402,N_15294);
nor U21148 (N_21148,N_14887,N_17944);
and U21149 (N_21149,N_15705,N_14986);
nor U21150 (N_21150,N_12260,N_12846);
or U21151 (N_21151,N_14155,N_12782);
xnor U21152 (N_21152,N_12872,N_13063);
xnor U21153 (N_21153,N_13642,N_15030);
nand U21154 (N_21154,N_12874,N_12244);
nand U21155 (N_21155,N_13789,N_17367);
or U21156 (N_21156,N_14748,N_13063);
nand U21157 (N_21157,N_13675,N_17178);
xnor U21158 (N_21158,N_14396,N_12575);
nand U21159 (N_21159,N_12672,N_14703);
nor U21160 (N_21160,N_15212,N_14420);
or U21161 (N_21161,N_16089,N_14923);
and U21162 (N_21162,N_12048,N_16522);
xor U21163 (N_21163,N_13657,N_13502);
nor U21164 (N_21164,N_13532,N_15463);
and U21165 (N_21165,N_15225,N_14250);
xnor U21166 (N_21166,N_16955,N_17039);
xor U21167 (N_21167,N_13515,N_16651);
or U21168 (N_21168,N_17475,N_17178);
and U21169 (N_21169,N_17796,N_13199);
or U21170 (N_21170,N_17519,N_15580);
xor U21171 (N_21171,N_15725,N_16426);
or U21172 (N_21172,N_17120,N_13658);
xnor U21173 (N_21173,N_13639,N_16048);
nand U21174 (N_21174,N_16208,N_12715);
nor U21175 (N_21175,N_12412,N_17460);
xor U21176 (N_21176,N_16340,N_14209);
nor U21177 (N_21177,N_16144,N_12000);
and U21178 (N_21178,N_14587,N_16675);
xor U21179 (N_21179,N_12066,N_14287);
or U21180 (N_21180,N_13289,N_16672);
nor U21181 (N_21181,N_14246,N_14335);
and U21182 (N_21182,N_13945,N_13858);
and U21183 (N_21183,N_12391,N_15351);
nand U21184 (N_21184,N_16495,N_15001);
or U21185 (N_21185,N_14979,N_16284);
or U21186 (N_21186,N_12620,N_17508);
nand U21187 (N_21187,N_12777,N_14645);
nor U21188 (N_21188,N_13519,N_15505);
nand U21189 (N_21189,N_14751,N_17530);
nand U21190 (N_21190,N_14015,N_12203);
nand U21191 (N_21191,N_13888,N_13414);
xor U21192 (N_21192,N_15134,N_16352);
and U21193 (N_21193,N_14214,N_13115);
or U21194 (N_21194,N_15573,N_12204);
nand U21195 (N_21195,N_17905,N_16245);
nor U21196 (N_21196,N_15717,N_13703);
or U21197 (N_21197,N_12972,N_12347);
xnor U21198 (N_21198,N_15051,N_14704);
nor U21199 (N_21199,N_17848,N_17600);
xor U21200 (N_21200,N_15305,N_16370);
and U21201 (N_21201,N_15519,N_14252);
and U21202 (N_21202,N_13588,N_12588);
or U21203 (N_21203,N_17414,N_17916);
nand U21204 (N_21204,N_14787,N_13801);
and U21205 (N_21205,N_16817,N_15802);
and U21206 (N_21206,N_13183,N_13529);
xor U21207 (N_21207,N_16474,N_12030);
or U21208 (N_21208,N_16681,N_13924);
and U21209 (N_21209,N_17202,N_13430);
or U21210 (N_21210,N_12092,N_16917);
nor U21211 (N_21211,N_13789,N_15084);
nand U21212 (N_21212,N_16502,N_15360);
nand U21213 (N_21213,N_14872,N_17662);
and U21214 (N_21214,N_13093,N_13214);
or U21215 (N_21215,N_12019,N_14304);
xnor U21216 (N_21216,N_16985,N_14392);
or U21217 (N_21217,N_16780,N_16694);
nand U21218 (N_21218,N_13835,N_12343);
nor U21219 (N_21219,N_14384,N_15661);
nand U21220 (N_21220,N_15557,N_12019);
nand U21221 (N_21221,N_15976,N_17283);
nor U21222 (N_21222,N_12209,N_13014);
xor U21223 (N_21223,N_13869,N_17772);
and U21224 (N_21224,N_16306,N_14976);
xnor U21225 (N_21225,N_12650,N_13430);
or U21226 (N_21226,N_15691,N_16663);
nand U21227 (N_21227,N_15057,N_14726);
or U21228 (N_21228,N_16777,N_14722);
or U21229 (N_21229,N_17713,N_13508);
and U21230 (N_21230,N_17532,N_15609);
nor U21231 (N_21231,N_13137,N_15731);
xor U21232 (N_21232,N_14700,N_15727);
or U21233 (N_21233,N_14818,N_13153);
xnor U21234 (N_21234,N_17961,N_14496);
nor U21235 (N_21235,N_17958,N_14480);
nor U21236 (N_21236,N_13673,N_13863);
xor U21237 (N_21237,N_17746,N_15477);
nor U21238 (N_21238,N_15618,N_16401);
or U21239 (N_21239,N_17482,N_12085);
or U21240 (N_21240,N_16349,N_14716);
xor U21241 (N_21241,N_15269,N_16199);
xor U21242 (N_21242,N_15364,N_15811);
nand U21243 (N_21243,N_14003,N_12359);
or U21244 (N_21244,N_16924,N_15554);
nor U21245 (N_21245,N_16279,N_16615);
or U21246 (N_21246,N_17193,N_14653);
nand U21247 (N_21247,N_16350,N_16726);
nand U21248 (N_21248,N_12603,N_17856);
or U21249 (N_21249,N_15983,N_15149);
and U21250 (N_21250,N_12035,N_14765);
or U21251 (N_21251,N_14334,N_16856);
or U21252 (N_21252,N_13739,N_14652);
and U21253 (N_21253,N_16806,N_17047);
or U21254 (N_21254,N_12024,N_16532);
nor U21255 (N_21255,N_16114,N_12485);
xor U21256 (N_21256,N_15418,N_17289);
or U21257 (N_21257,N_17515,N_17639);
and U21258 (N_21258,N_17348,N_13162);
nor U21259 (N_21259,N_13924,N_12001);
or U21260 (N_21260,N_15644,N_16364);
or U21261 (N_21261,N_14600,N_17273);
nor U21262 (N_21262,N_17971,N_12981);
nor U21263 (N_21263,N_17862,N_15547);
or U21264 (N_21264,N_17140,N_14708);
nand U21265 (N_21265,N_17695,N_13882);
xnor U21266 (N_21266,N_17337,N_17816);
xor U21267 (N_21267,N_16125,N_16554);
xnor U21268 (N_21268,N_15453,N_17897);
nand U21269 (N_21269,N_17991,N_12244);
or U21270 (N_21270,N_12422,N_16217);
xnor U21271 (N_21271,N_16029,N_15351);
or U21272 (N_21272,N_14862,N_17246);
xor U21273 (N_21273,N_14695,N_12402);
or U21274 (N_21274,N_13647,N_13139);
nor U21275 (N_21275,N_14442,N_13036);
nor U21276 (N_21276,N_17054,N_12594);
nor U21277 (N_21277,N_14874,N_14810);
and U21278 (N_21278,N_12289,N_17297);
nand U21279 (N_21279,N_13809,N_15317);
nor U21280 (N_21280,N_12162,N_12849);
nor U21281 (N_21281,N_13780,N_16531);
nand U21282 (N_21282,N_17555,N_14724);
or U21283 (N_21283,N_16455,N_16506);
nand U21284 (N_21284,N_13605,N_12868);
nor U21285 (N_21285,N_13365,N_17919);
nor U21286 (N_21286,N_12606,N_16817);
nand U21287 (N_21287,N_17397,N_16999);
nor U21288 (N_21288,N_14932,N_12937);
and U21289 (N_21289,N_13605,N_13815);
xor U21290 (N_21290,N_14441,N_12506);
nor U21291 (N_21291,N_15530,N_12383);
and U21292 (N_21292,N_13313,N_15938);
nor U21293 (N_21293,N_14936,N_12358);
or U21294 (N_21294,N_15548,N_14590);
nand U21295 (N_21295,N_14250,N_13674);
and U21296 (N_21296,N_12955,N_14825);
nor U21297 (N_21297,N_15654,N_13949);
xor U21298 (N_21298,N_17381,N_12544);
nand U21299 (N_21299,N_14841,N_12698);
xnor U21300 (N_21300,N_15542,N_16641);
and U21301 (N_21301,N_15538,N_15819);
xor U21302 (N_21302,N_13140,N_13897);
or U21303 (N_21303,N_17336,N_13128);
and U21304 (N_21304,N_14286,N_15863);
nand U21305 (N_21305,N_17767,N_12736);
nand U21306 (N_21306,N_12147,N_16938);
nand U21307 (N_21307,N_15531,N_17282);
or U21308 (N_21308,N_13598,N_17799);
or U21309 (N_21309,N_12092,N_17588);
nand U21310 (N_21310,N_16932,N_15443);
xnor U21311 (N_21311,N_12821,N_13222);
nor U21312 (N_21312,N_15028,N_16877);
xnor U21313 (N_21313,N_16329,N_17773);
nor U21314 (N_21314,N_12411,N_16014);
nor U21315 (N_21315,N_13528,N_14880);
and U21316 (N_21316,N_17600,N_16579);
nor U21317 (N_21317,N_17466,N_13920);
xnor U21318 (N_21318,N_16759,N_17816);
nor U21319 (N_21319,N_15959,N_16744);
or U21320 (N_21320,N_12764,N_16405);
nand U21321 (N_21321,N_17749,N_17273);
nor U21322 (N_21322,N_12796,N_14897);
or U21323 (N_21323,N_16005,N_15716);
or U21324 (N_21324,N_17679,N_16046);
nor U21325 (N_21325,N_15482,N_14087);
xnor U21326 (N_21326,N_15391,N_15746);
or U21327 (N_21327,N_12076,N_13727);
or U21328 (N_21328,N_12682,N_16130);
or U21329 (N_21329,N_17238,N_13147);
and U21330 (N_21330,N_15644,N_14481);
xnor U21331 (N_21331,N_13012,N_13659);
or U21332 (N_21332,N_16384,N_13265);
xor U21333 (N_21333,N_12304,N_12252);
nand U21334 (N_21334,N_16561,N_17015);
nor U21335 (N_21335,N_17365,N_13975);
xor U21336 (N_21336,N_15521,N_13015);
and U21337 (N_21337,N_15537,N_15521);
or U21338 (N_21338,N_14344,N_12619);
xnor U21339 (N_21339,N_15071,N_15729);
and U21340 (N_21340,N_17816,N_16378);
and U21341 (N_21341,N_16522,N_16557);
and U21342 (N_21342,N_15249,N_14685);
nor U21343 (N_21343,N_12670,N_12775);
or U21344 (N_21344,N_13659,N_14902);
nand U21345 (N_21345,N_16880,N_15008);
xor U21346 (N_21346,N_15392,N_17302);
and U21347 (N_21347,N_15467,N_16238);
or U21348 (N_21348,N_17095,N_15600);
or U21349 (N_21349,N_13051,N_14567);
and U21350 (N_21350,N_13509,N_17941);
nor U21351 (N_21351,N_12110,N_15162);
xor U21352 (N_21352,N_15348,N_14545);
and U21353 (N_21353,N_17721,N_17455);
nor U21354 (N_21354,N_17111,N_12575);
xor U21355 (N_21355,N_13163,N_14246);
nand U21356 (N_21356,N_16865,N_12910);
xnor U21357 (N_21357,N_12259,N_13087);
nand U21358 (N_21358,N_12724,N_13626);
or U21359 (N_21359,N_16520,N_13426);
and U21360 (N_21360,N_13437,N_14323);
or U21361 (N_21361,N_17659,N_14531);
or U21362 (N_21362,N_14619,N_13196);
nand U21363 (N_21363,N_15915,N_17182);
xor U21364 (N_21364,N_17599,N_16645);
xor U21365 (N_21365,N_15298,N_17467);
nand U21366 (N_21366,N_16659,N_14271);
and U21367 (N_21367,N_15018,N_12939);
xnor U21368 (N_21368,N_15154,N_12282);
or U21369 (N_21369,N_15222,N_15755);
and U21370 (N_21370,N_17346,N_15952);
and U21371 (N_21371,N_12792,N_16071);
xor U21372 (N_21372,N_15889,N_13039);
nand U21373 (N_21373,N_15947,N_16420);
or U21374 (N_21374,N_12383,N_12304);
and U21375 (N_21375,N_12419,N_13245);
nor U21376 (N_21376,N_15848,N_15101);
and U21377 (N_21377,N_17947,N_17650);
or U21378 (N_21378,N_13211,N_14815);
nor U21379 (N_21379,N_17952,N_12334);
nand U21380 (N_21380,N_13878,N_15713);
and U21381 (N_21381,N_17637,N_12459);
or U21382 (N_21382,N_15490,N_13373);
xor U21383 (N_21383,N_12942,N_16628);
nor U21384 (N_21384,N_14718,N_13973);
xnor U21385 (N_21385,N_17852,N_16286);
nor U21386 (N_21386,N_12247,N_15271);
or U21387 (N_21387,N_14326,N_14161);
xor U21388 (N_21388,N_14005,N_12638);
xor U21389 (N_21389,N_12032,N_13843);
xnor U21390 (N_21390,N_17674,N_17857);
nor U21391 (N_21391,N_15228,N_13615);
nor U21392 (N_21392,N_17068,N_14163);
nand U21393 (N_21393,N_13570,N_13589);
and U21394 (N_21394,N_13533,N_14134);
nand U21395 (N_21395,N_16265,N_13069);
xnor U21396 (N_21396,N_16858,N_14842);
xnor U21397 (N_21397,N_16753,N_15594);
nor U21398 (N_21398,N_13734,N_15324);
or U21399 (N_21399,N_16191,N_14970);
nor U21400 (N_21400,N_12049,N_12563);
nand U21401 (N_21401,N_15966,N_13247);
or U21402 (N_21402,N_16733,N_14350);
and U21403 (N_21403,N_15432,N_13342);
and U21404 (N_21404,N_15915,N_14168);
and U21405 (N_21405,N_12918,N_13023);
nor U21406 (N_21406,N_17400,N_14741);
and U21407 (N_21407,N_14167,N_12200);
xor U21408 (N_21408,N_12366,N_15642);
xor U21409 (N_21409,N_13132,N_17059);
xnor U21410 (N_21410,N_15693,N_14154);
or U21411 (N_21411,N_15979,N_16428);
or U21412 (N_21412,N_17037,N_16893);
nor U21413 (N_21413,N_14763,N_15931);
or U21414 (N_21414,N_13594,N_12967);
or U21415 (N_21415,N_13915,N_14216);
xnor U21416 (N_21416,N_15034,N_15019);
and U21417 (N_21417,N_13241,N_17940);
or U21418 (N_21418,N_12022,N_15827);
xnor U21419 (N_21419,N_17571,N_17144);
nor U21420 (N_21420,N_12145,N_16383);
and U21421 (N_21421,N_17387,N_17541);
or U21422 (N_21422,N_12432,N_15299);
and U21423 (N_21423,N_13222,N_15653);
nand U21424 (N_21424,N_16874,N_15179);
xor U21425 (N_21425,N_17686,N_16126);
xnor U21426 (N_21426,N_12633,N_14325);
and U21427 (N_21427,N_15228,N_15234);
and U21428 (N_21428,N_16677,N_13898);
nand U21429 (N_21429,N_16289,N_15097);
nor U21430 (N_21430,N_14910,N_16534);
nor U21431 (N_21431,N_12420,N_13679);
nor U21432 (N_21432,N_12487,N_14621);
nor U21433 (N_21433,N_12567,N_13031);
or U21434 (N_21434,N_14355,N_14795);
xor U21435 (N_21435,N_15865,N_16554);
nor U21436 (N_21436,N_17296,N_13563);
nand U21437 (N_21437,N_13148,N_14604);
and U21438 (N_21438,N_15240,N_14795);
or U21439 (N_21439,N_12499,N_13812);
or U21440 (N_21440,N_14084,N_14677);
xor U21441 (N_21441,N_17136,N_16502);
nor U21442 (N_21442,N_17404,N_16220);
nand U21443 (N_21443,N_12741,N_16940);
xnor U21444 (N_21444,N_12536,N_16619);
nand U21445 (N_21445,N_16764,N_14281);
xor U21446 (N_21446,N_12132,N_13932);
or U21447 (N_21447,N_13888,N_17361);
xor U21448 (N_21448,N_14609,N_12343);
or U21449 (N_21449,N_13045,N_14115);
nor U21450 (N_21450,N_15616,N_16599);
nand U21451 (N_21451,N_12198,N_14167);
nor U21452 (N_21452,N_16475,N_15238);
xor U21453 (N_21453,N_16063,N_17658);
nand U21454 (N_21454,N_13716,N_13155);
nand U21455 (N_21455,N_13801,N_14269);
nand U21456 (N_21456,N_12391,N_13274);
and U21457 (N_21457,N_14617,N_17066);
nand U21458 (N_21458,N_14478,N_12482);
nand U21459 (N_21459,N_12848,N_16079);
or U21460 (N_21460,N_12464,N_16361);
nor U21461 (N_21461,N_16066,N_12997);
xnor U21462 (N_21462,N_16291,N_15918);
nor U21463 (N_21463,N_12047,N_16078);
or U21464 (N_21464,N_16156,N_14020);
xnor U21465 (N_21465,N_16338,N_13131);
or U21466 (N_21466,N_12707,N_15732);
and U21467 (N_21467,N_14194,N_17115);
nand U21468 (N_21468,N_15294,N_13899);
or U21469 (N_21469,N_14533,N_14034);
nand U21470 (N_21470,N_16244,N_17215);
or U21471 (N_21471,N_15992,N_13046);
nand U21472 (N_21472,N_16627,N_16104);
or U21473 (N_21473,N_15426,N_14079);
nor U21474 (N_21474,N_12708,N_13235);
nand U21475 (N_21475,N_12589,N_16735);
and U21476 (N_21476,N_12914,N_12462);
and U21477 (N_21477,N_16297,N_16622);
xnor U21478 (N_21478,N_12741,N_16670);
and U21479 (N_21479,N_13211,N_12051);
nand U21480 (N_21480,N_17141,N_14980);
xor U21481 (N_21481,N_15907,N_12977);
xor U21482 (N_21482,N_12689,N_15339);
nor U21483 (N_21483,N_13722,N_17235);
xor U21484 (N_21484,N_14050,N_14048);
or U21485 (N_21485,N_15267,N_17466);
nor U21486 (N_21486,N_13399,N_14395);
or U21487 (N_21487,N_16156,N_17175);
xor U21488 (N_21488,N_17719,N_15121);
xor U21489 (N_21489,N_13500,N_16128);
or U21490 (N_21490,N_14059,N_16678);
nand U21491 (N_21491,N_13631,N_15807);
nand U21492 (N_21492,N_15119,N_13335);
xnor U21493 (N_21493,N_12241,N_13695);
or U21494 (N_21494,N_14595,N_16635);
nand U21495 (N_21495,N_12243,N_12715);
or U21496 (N_21496,N_12341,N_17433);
or U21497 (N_21497,N_13045,N_15415);
nor U21498 (N_21498,N_17210,N_13816);
xor U21499 (N_21499,N_17258,N_17227);
or U21500 (N_21500,N_12232,N_12678);
and U21501 (N_21501,N_14063,N_13634);
and U21502 (N_21502,N_13868,N_12393);
and U21503 (N_21503,N_15524,N_15526);
xnor U21504 (N_21504,N_16361,N_16593);
nor U21505 (N_21505,N_16519,N_17815);
nor U21506 (N_21506,N_17567,N_13264);
and U21507 (N_21507,N_15368,N_14970);
or U21508 (N_21508,N_14530,N_16048);
or U21509 (N_21509,N_13275,N_12462);
and U21510 (N_21510,N_13684,N_15101);
nand U21511 (N_21511,N_15738,N_13971);
xor U21512 (N_21512,N_14366,N_13147);
nor U21513 (N_21513,N_15137,N_16911);
nor U21514 (N_21514,N_12252,N_12585);
xor U21515 (N_21515,N_16871,N_12156);
nand U21516 (N_21516,N_16060,N_12066);
xnor U21517 (N_21517,N_16343,N_16020);
nor U21518 (N_21518,N_16897,N_14558);
or U21519 (N_21519,N_15334,N_12233);
xnor U21520 (N_21520,N_16531,N_14699);
nor U21521 (N_21521,N_14298,N_14735);
or U21522 (N_21522,N_16539,N_12192);
nor U21523 (N_21523,N_14078,N_15219);
and U21524 (N_21524,N_13611,N_17571);
or U21525 (N_21525,N_15093,N_15043);
or U21526 (N_21526,N_14656,N_16375);
nor U21527 (N_21527,N_12653,N_17066);
and U21528 (N_21528,N_13807,N_14247);
or U21529 (N_21529,N_16019,N_14242);
or U21530 (N_21530,N_13877,N_12516);
xor U21531 (N_21531,N_13320,N_12349);
or U21532 (N_21532,N_14865,N_12493);
and U21533 (N_21533,N_15389,N_12482);
nor U21534 (N_21534,N_13295,N_12576);
nand U21535 (N_21535,N_16899,N_12113);
or U21536 (N_21536,N_14574,N_16896);
nand U21537 (N_21537,N_16952,N_15582);
and U21538 (N_21538,N_15335,N_15834);
or U21539 (N_21539,N_14558,N_17721);
xor U21540 (N_21540,N_13218,N_14230);
and U21541 (N_21541,N_16102,N_12525);
nand U21542 (N_21542,N_12501,N_12165);
or U21543 (N_21543,N_13757,N_15118);
or U21544 (N_21544,N_17799,N_17005);
or U21545 (N_21545,N_12836,N_14040);
or U21546 (N_21546,N_16421,N_13841);
nor U21547 (N_21547,N_12123,N_13951);
nor U21548 (N_21548,N_16703,N_14977);
and U21549 (N_21549,N_12480,N_12760);
or U21550 (N_21550,N_13249,N_14884);
xnor U21551 (N_21551,N_15284,N_17941);
xnor U21552 (N_21552,N_14156,N_15385);
nor U21553 (N_21553,N_17107,N_15884);
and U21554 (N_21554,N_14468,N_12391);
nand U21555 (N_21555,N_13848,N_12532);
xor U21556 (N_21556,N_13117,N_15826);
nand U21557 (N_21557,N_15928,N_15731);
nand U21558 (N_21558,N_14960,N_13945);
nor U21559 (N_21559,N_15621,N_12833);
and U21560 (N_21560,N_15141,N_14660);
and U21561 (N_21561,N_15699,N_13532);
and U21562 (N_21562,N_13878,N_16380);
or U21563 (N_21563,N_12219,N_14802);
xor U21564 (N_21564,N_16424,N_13269);
and U21565 (N_21565,N_12856,N_15041);
or U21566 (N_21566,N_12496,N_12007);
xnor U21567 (N_21567,N_16872,N_17419);
xor U21568 (N_21568,N_16875,N_17083);
or U21569 (N_21569,N_16796,N_15533);
nand U21570 (N_21570,N_13064,N_12532);
xnor U21571 (N_21571,N_16759,N_12937);
nor U21572 (N_21572,N_13041,N_16277);
nand U21573 (N_21573,N_12430,N_15637);
xor U21574 (N_21574,N_12300,N_16991);
nand U21575 (N_21575,N_13758,N_17323);
or U21576 (N_21576,N_12516,N_17767);
nand U21577 (N_21577,N_12221,N_14522);
nor U21578 (N_21578,N_15112,N_12509);
and U21579 (N_21579,N_16275,N_17607);
nor U21580 (N_21580,N_15577,N_14023);
and U21581 (N_21581,N_13489,N_16804);
nor U21582 (N_21582,N_15072,N_12171);
and U21583 (N_21583,N_17532,N_12833);
or U21584 (N_21584,N_15558,N_16427);
xnor U21585 (N_21585,N_16347,N_17616);
and U21586 (N_21586,N_16770,N_16437);
xnor U21587 (N_21587,N_17788,N_12926);
nand U21588 (N_21588,N_13808,N_14846);
nor U21589 (N_21589,N_16658,N_12225);
xnor U21590 (N_21590,N_17734,N_12202);
and U21591 (N_21591,N_17224,N_14630);
nor U21592 (N_21592,N_14753,N_15881);
or U21593 (N_21593,N_14342,N_14733);
and U21594 (N_21594,N_12077,N_14949);
nand U21595 (N_21595,N_12426,N_12947);
and U21596 (N_21596,N_17744,N_15089);
and U21597 (N_21597,N_14019,N_14587);
nand U21598 (N_21598,N_14195,N_14457);
and U21599 (N_21599,N_15542,N_12692);
nor U21600 (N_21600,N_17245,N_15979);
nor U21601 (N_21601,N_13099,N_13669);
nor U21602 (N_21602,N_16439,N_14835);
or U21603 (N_21603,N_13341,N_15036);
or U21604 (N_21604,N_16928,N_16328);
and U21605 (N_21605,N_16084,N_14235);
or U21606 (N_21606,N_12282,N_12444);
nor U21607 (N_21607,N_16670,N_13335);
nand U21608 (N_21608,N_14360,N_13147);
nand U21609 (N_21609,N_17224,N_13433);
nand U21610 (N_21610,N_17043,N_12587);
xnor U21611 (N_21611,N_12552,N_17907);
nor U21612 (N_21612,N_13394,N_16333);
xor U21613 (N_21613,N_16280,N_16346);
xor U21614 (N_21614,N_15486,N_12014);
xnor U21615 (N_21615,N_12060,N_15748);
or U21616 (N_21616,N_14061,N_15249);
xor U21617 (N_21617,N_13770,N_14623);
nor U21618 (N_21618,N_13459,N_16858);
nand U21619 (N_21619,N_17245,N_13133);
xor U21620 (N_21620,N_13065,N_17849);
nand U21621 (N_21621,N_17812,N_16039);
nand U21622 (N_21622,N_15913,N_15238);
and U21623 (N_21623,N_17193,N_16707);
or U21624 (N_21624,N_12601,N_13314);
nand U21625 (N_21625,N_14272,N_12721);
xnor U21626 (N_21626,N_17480,N_17717);
nand U21627 (N_21627,N_16119,N_15109);
and U21628 (N_21628,N_15648,N_15517);
nor U21629 (N_21629,N_12023,N_17828);
or U21630 (N_21630,N_16946,N_13645);
and U21631 (N_21631,N_14413,N_15307);
nor U21632 (N_21632,N_17893,N_12602);
nand U21633 (N_21633,N_16052,N_16428);
nand U21634 (N_21634,N_14144,N_17909);
nand U21635 (N_21635,N_15764,N_14631);
xnor U21636 (N_21636,N_14255,N_16823);
nor U21637 (N_21637,N_17350,N_13865);
nand U21638 (N_21638,N_15596,N_15005);
and U21639 (N_21639,N_13720,N_14357);
nor U21640 (N_21640,N_12927,N_13339);
or U21641 (N_21641,N_12267,N_14480);
nand U21642 (N_21642,N_16484,N_16425);
xnor U21643 (N_21643,N_12985,N_15350);
xnor U21644 (N_21644,N_16096,N_17781);
nand U21645 (N_21645,N_15936,N_15544);
nand U21646 (N_21646,N_13976,N_13348);
or U21647 (N_21647,N_12656,N_17140);
xor U21648 (N_21648,N_13654,N_16948);
or U21649 (N_21649,N_12971,N_12143);
and U21650 (N_21650,N_15495,N_12525);
nand U21651 (N_21651,N_16163,N_17351);
nand U21652 (N_21652,N_14742,N_12562);
or U21653 (N_21653,N_16386,N_16634);
or U21654 (N_21654,N_16382,N_12344);
nand U21655 (N_21655,N_12695,N_12738);
and U21656 (N_21656,N_13328,N_17524);
xnor U21657 (N_21657,N_15945,N_16328);
nand U21658 (N_21658,N_16331,N_12119);
nand U21659 (N_21659,N_17462,N_15265);
nand U21660 (N_21660,N_13082,N_15783);
nand U21661 (N_21661,N_17396,N_16233);
nand U21662 (N_21662,N_16012,N_12683);
nand U21663 (N_21663,N_14077,N_12083);
or U21664 (N_21664,N_16968,N_17454);
and U21665 (N_21665,N_12330,N_13357);
and U21666 (N_21666,N_17564,N_16861);
and U21667 (N_21667,N_13034,N_15355);
or U21668 (N_21668,N_15600,N_14557);
xor U21669 (N_21669,N_12824,N_16271);
or U21670 (N_21670,N_16664,N_12086);
or U21671 (N_21671,N_13020,N_14384);
nand U21672 (N_21672,N_12848,N_14317);
or U21673 (N_21673,N_12313,N_16312);
or U21674 (N_21674,N_17901,N_14918);
or U21675 (N_21675,N_13978,N_13479);
or U21676 (N_21676,N_14948,N_17092);
and U21677 (N_21677,N_15934,N_14101);
and U21678 (N_21678,N_17163,N_14796);
and U21679 (N_21679,N_16035,N_16592);
xnor U21680 (N_21680,N_16581,N_12183);
nand U21681 (N_21681,N_17118,N_17097);
xnor U21682 (N_21682,N_12356,N_15850);
or U21683 (N_21683,N_15287,N_16370);
nand U21684 (N_21684,N_13266,N_14384);
nand U21685 (N_21685,N_13042,N_15914);
nand U21686 (N_21686,N_15669,N_15764);
and U21687 (N_21687,N_13356,N_15138);
xor U21688 (N_21688,N_16618,N_13385);
and U21689 (N_21689,N_16768,N_14325);
nor U21690 (N_21690,N_12121,N_14364);
or U21691 (N_21691,N_16960,N_13021);
xnor U21692 (N_21692,N_15288,N_13099);
or U21693 (N_21693,N_16963,N_15989);
or U21694 (N_21694,N_15734,N_14569);
nand U21695 (N_21695,N_16808,N_14341);
and U21696 (N_21696,N_16608,N_14928);
or U21697 (N_21697,N_13539,N_12269);
nand U21698 (N_21698,N_13294,N_17245);
xnor U21699 (N_21699,N_13424,N_12125);
nor U21700 (N_21700,N_16148,N_12872);
or U21701 (N_21701,N_15746,N_13301);
nor U21702 (N_21702,N_17948,N_17054);
and U21703 (N_21703,N_16498,N_15179);
nor U21704 (N_21704,N_17247,N_14755);
nand U21705 (N_21705,N_17050,N_16790);
and U21706 (N_21706,N_16734,N_13594);
and U21707 (N_21707,N_13394,N_15167);
xnor U21708 (N_21708,N_16084,N_16408);
nand U21709 (N_21709,N_12211,N_15036);
nand U21710 (N_21710,N_14194,N_17059);
nand U21711 (N_21711,N_13445,N_14079);
nor U21712 (N_21712,N_14042,N_12200);
nand U21713 (N_21713,N_15097,N_15656);
nor U21714 (N_21714,N_13145,N_13977);
and U21715 (N_21715,N_14336,N_17045);
or U21716 (N_21716,N_16800,N_14355);
or U21717 (N_21717,N_12391,N_17490);
and U21718 (N_21718,N_12421,N_17732);
or U21719 (N_21719,N_15778,N_12819);
xor U21720 (N_21720,N_17136,N_13773);
or U21721 (N_21721,N_17369,N_12757);
and U21722 (N_21722,N_14889,N_17373);
nor U21723 (N_21723,N_12067,N_12644);
nand U21724 (N_21724,N_14889,N_14262);
nand U21725 (N_21725,N_12450,N_13424);
or U21726 (N_21726,N_17172,N_13529);
nor U21727 (N_21727,N_15166,N_16233);
or U21728 (N_21728,N_14923,N_16960);
nand U21729 (N_21729,N_17321,N_14307);
and U21730 (N_21730,N_14073,N_15602);
nand U21731 (N_21731,N_16783,N_12080);
and U21732 (N_21732,N_15855,N_12798);
nand U21733 (N_21733,N_13940,N_16633);
and U21734 (N_21734,N_16576,N_16416);
nand U21735 (N_21735,N_13181,N_15845);
nor U21736 (N_21736,N_12008,N_12323);
nor U21737 (N_21737,N_16770,N_17856);
xnor U21738 (N_21738,N_14194,N_16096);
and U21739 (N_21739,N_14561,N_14814);
or U21740 (N_21740,N_14694,N_12029);
or U21741 (N_21741,N_17219,N_13479);
xnor U21742 (N_21742,N_17995,N_14871);
xor U21743 (N_21743,N_13524,N_13927);
nand U21744 (N_21744,N_14280,N_15307);
or U21745 (N_21745,N_15615,N_17812);
and U21746 (N_21746,N_13017,N_15959);
or U21747 (N_21747,N_17166,N_17640);
and U21748 (N_21748,N_14130,N_14518);
or U21749 (N_21749,N_14845,N_13337);
xor U21750 (N_21750,N_14303,N_13756);
xnor U21751 (N_21751,N_14324,N_14676);
nor U21752 (N_21752,N_15425,N_16595);
nand U21753 (N_21753,N_15744,N_17681);
nand U21754 (N_21754,N_17028,N_13494);
nand U21755 (N_21755,N_15903,N_16437);
or U21756 (N_21756,N_15734,N_16593);
or U21757 (N_21757,N_17532,N_12351);
xnor U21758 (N_21758,N_14600,N_12316);
or U21759 (N_21759,N_13766,N_12928);
nor U21760 (N_21760,N_12116,N_17957);
nand U21761 (N_21761,N_15564,N_16488);
xor U21762 (N_21762,N_12708,N_15538);
xor U21763 (N_21763,N_13564,N_16327);
nor U21764 (N_21764,N_12495,N_12947);
or U21765 (N_21765,N_13065,N_14034);
nor U21766 (N_21766,N_13306,N_16107);
or U21767 (N_21767,N_15180,N_16626);
nand U21768 (N_21768,N_17448,N_16263);
nor U21769 (N_21769,N_12657,N_17372);
or U21770 (N_21770,N_16551,N_15515);
xnor U21771 (N_21771,N_13792,N_16681);
nand U21772 (N_21772,N_13201,N_12252);
or U21773 (N_21773,N_13896,N_16727);
nand U21774 (N_21774,N_17079,N_14360);
or U21775 (N_21775,N_17380,N_12792);
nand U21776 (N_21776,N_15512,N_12205);
nand U21777 (N_21777,N_12169,N_17935);
xnor U21778 (N_21778,N_15690,N_12593);
nand U21779 (N_21779,N_15151,N_17038);
nand U21780 (N_21780,N_16582,N_13547);
nand U21781 (N_21781,N_17364,N_17770);
xnor U21782 (N_21782,N_12436,N_12197);
and U21783 (N_21783,N_13400,N_12844);
xor U21784 (N_21784,N_13616,N_13147);
nand U21785 (N_21785,N_13861,N_16111);
nor U21786 (N_21786,N_17989,N_17750);
nor U21787 (N_21787,N_14822,N_16031);
nand U21788 (N_21788,N_12402,N_14552);
xnor U21789 (N_21789,N_12947,N_12412);
or U21790 (N_21790,N_15792,N_14801);
xor U21791 (N_21791,N_14101,N_12712);
nor U21792 (N_21792,N_15404,N_12530);
nand U21793 (N_21793,N_12685,N_14428);
or U21794 (N_21794,N_13046,N_17648);
xnor U21795 (N_21795,N_15077,N_12815);
nand U21796 (N_21796,N_13667,N_13180);
nand U21797 (N_21797,N_13726,N_14481);
or U21798 (N_21798,N_14161,N_12323);
nor U21799 (N_21799,N_12723,N_17287);
xnor U21800 (N_21800,N_16432,N_14794);
nor U21801 (N_21801,N_14097,N_15438);
and U21802 (N_21802,N_15041,N_17559);
nor U21803 (N_21803,N_13385,N_14439);
xnor U21804 (N_21804,N_16845,N_12495);
or U21805 (N_21805,N_17259,N_12218);
xnor U21806 (N_21806,N_14077,N_13893);
nor U21807 (N_21807,N_15341,N_15945);
nand U21808 (N_21808,N_12232,N_16003);
nand U21809 (N_21809,N_14489,N_17304);
xnor U21810 (N_21810,N_17010,N_15285);
nand U21811 (N_21811,N_14447,N_12450);
and U21812 (N_21812,N_14291,N_14333);
and U21813 (N_21813,N_17218,N_14576);
nor U21814 (N_21814,N_16674,N_16653);
nor U21815 (N_21815,N_17793,N_14506);
nand U21816 (N_21816,N_14277,N_14143);
xnor U21817 (N_21817,N_16374,N_12806);
nand U21818 (N_21818,N_17125,N_13959);
or U21819 (N_21819,N_13435,N_17932);
and U21820 (N_21820,N_13497,N_17083);
or U21821 (N_21821,N_17084,N_14491);
nand U21822 (N_21822,N_15557,N_13808);
and U21823 (N_21823,N_15820,N_15873);
and U21824 (N_21824,N_13286,N_13125);
or U21825 (N_21825,N_16098,N_14814);
and U21826 (N_21826,N_16537,N_17426);
nand U21827 (N_21827,N_15794,N_12506);
and U21828 (N_21828,N_17833,N_13716);
nor U21829 (N_21829,N_12745,N_13254);
xor U21830 (N_21830,N_14964,N_13895);
nand U21831 (N_21831,N_16598,N_17324);
nand U21832 (N_21832,N_17022,N_17258);
or U21833 (N_21833,N_17057,N_17464);
xnor U21834 (N_21834,N_12916,N_13687);
or U21835 (N_21835,N_14892,N_15096);
and U21836 (N_21836,N_16200,N_13125);
nand U21837 (N_21837,N_13389,N_15094);
nand U21838 (N_21838,N_15857,N_13621);
and U21839 (N_21839,N_15352,N_16546);
and U21840 (N_21840,N_14019,N_16350);
or U21841 (N_21841,N_16731,N_14099);
and U21842 (N_21842,N_15920,N_17520);
and U21843 (N_21843,N_17026,N_13078);
nor U21844 (N_21844,N_17775,N_13602);
or U21845 (N_21845,N_12157,N_15462);
nor U21846 (N_21846,N_14614,N_13449);
nand U21847 (N_21847,N_16742,N_16514);
and U21848 (N_21848,N_14758,N_14951);
nand U21849 (N_21849,N_15807,N_17886);
nor U21850 (N_21850,N_17743,N_12155);
nand U21851 (N_21851,N_16644,N_13103);
xnor U21852 (N_21852,N_13132,N_16128);
and U21853 (N_21853,N_12838,N_12816);
and U21854 (N_21854,N_14305,N_12890);
and U21855 (N_21855,N_16564,N_12655);
nor U21856 (N_21856,N_17828,N_12221);
or U21857 (N_21857,N_17640,N_16029);
and U21858 (N_21858,N_16382,N_16336);
nand U21859 (N_21859,N_15382,N_14898);
xor U21860 (N_21860,N_12354,N_17615);
nand U21861 (N_21861,N_16683,N_17864);
or U21862 (N_21862,N_16686,N_13055);
xnor U21863 (N_21863,N_14350,N_16975);
or U21864 (N_21864,N_16086,N_15660);
nand U21865 (N_21865,N_13076,N_13694);
or U21866 (N_21866,N_14703,N_12787);
nor U21867 (N_21867,N_14344,N_13041);
xnor U21868 (N_21868,N_16142,N_17856);
and U21869 (N_21869,N_14915,N_17072);
xor U21870 (N_21870,N_16395,N_13872);
nand U21871 (N_21871,N_14967,N_14556);
nor U21872 (N_21872,N_16792,N_17922);
xor U21873 (N_21873,N_14054,N_16659);
or U21874 (N_21874,N_16258,N_17480);
xor U21875 (N_21875,N_15521,N_17098);
or U21876 (N_21876,N_13895,N_15235);
and U21877 (N_21877,N_14130,N_15708);
nand U21878 (N_21878,N_17182,N_12271);
nand U21879 (N_21879,N_14586,N_14952);
and U21880 (N_21880,N_15581,N_16837);
or U21881 (N_21881,N_14225,N_15209);
nor U21882 (N_21882,N_17057,N_14140);
and U21883 (N_21883,N_17993,N_14947);
xor U21884 (N_21884,N_17512,N_12962);
nor U21885 (N_21885,N_12852,N_13148);
or U21886 (N_21886,N_17765,N_17405);
nand U21887 (N_21887,N_15095,N_16411);
and U21888 (N_21888,N_17423,N_13273);
or U21889 (N_21889,N_12018,N_16560);
and U21890 (N_21890,N_13274,N_12204);
or U21891 (N_21891,N_13081,N_16984);
xor U21892 (N_21892,N_12021,N_12870);
and U21893 (N_21893,N_14121,N_17489);
nor U21894 (N_21894,N_13320,N_12562);
nand U21895 (N_21895,N_13103,N_14184);
xnor U21896 (N_21896,N_12301,N_15293);
or U21897 (N_21897,N_14726,N_16424);
and U21898 (N_21898,N_16369,N_13963);
nor U21899 (N_21899,N_17193,N_13906);
xor U21900 (N_21900,N_12000,N_13276);
or U21901 (N_21901,N_16931,N_13821);
xnor U21902 (N_21902,N_14221,N_12155);
or U21903 (N_21903,N_16472,N_14390);
xor U21904 (N_21904,N_12766,N_14902);
and U21905 (N_21905,N_12336,N_13672);
nand U21906 (N_21906,N_15162,N_17312);
and U21907 (N_21907,N_13626,N_17829);
or U21908 (N_21908,N_15624,N_13002);
nor U21909 (N_21909,N_13618,N_16260);
xor U21910 (N_21910,N_13352,N_16681);
nor U21911 (N_21911,N_13250,N_15997);
xor U21912 (N_21912,N_12619,N_15270);
or U21913 (N_21913,N_16044,N_17769);
nor U21914 (N_21914,N_12977,N_16310);
nand U21915 (N_21915,N_12837,N_14076);
or U21916 (N_21916,N_17311,N_17357);
or U21917 (N_21917,N_17211,N_13338);
nand U21918 (N_21918,N_17996,N_14326);
or U21919 (N_21919,N_15148,N_17385);
or U21920 (N_21920,N_17584,N_14377);
or U21921 (N_21921,N_14384,N_17549);
xnor U21922 (N_21922,N_12321,N_13964);
nor U21923 (N_21923,N_13868,N_14035);
nor U21924 (N_21924,N_12645,N_14400);
nor U21925 (N_21925,N_14164,N_13934);
nand U21926 (N_21926,N_16316,N_16197);
xnor U21927 (N_21927,N_13216,N_15066);
nor U21928 (N_21928,N_15192,N_14766);
nand U21929 (N_21929,N_15081,N_17269);
xor U21930 (N_21930,N_17919,N_17616);
and U21931 (N_21931,N_14656,N_12429);
xnor U21932 (N_21932,N_12945,N_17764);
and U21933 (N_21933,N_15447,N_16362);
xnor U21934 (N_21934,N_15078,N_16608);
xnor U21935 (N_21935,N_17142,N_12170);
or U21936 (N_21936,N_13094,N_14978);
and U21937 (N_21937,N_16698,N_12186);
xor U21938 (N_21938,N_16180,N_12208);
xor U21939 (N_21939,N_12896,N_16343);
and U21940 (N_21940,N_14448,N_16500);
xor U21941 (N_21941,N_13661,N_14903);
nand U21942 (N_21942,N_15562,N_16608);
or U21943 (N_21943,N_12738,N_14809);
xor U21944 (N_21944,N_16897,N_13143);
or U21945 (N_21945,N_14241,N_14004);
and U21946 (N_21946,N_13665,N_16450);
xor U21947 (N_21947,N_17270,N_16210);
nor U21948 (N_21948,N_12982,N_17093);
xor U21949 (N_21949,N_13034,N_15544);
nor U21950 (N_21950,N_16213,N_16105);
nor U21951 (N_21951,N_16177,N_16210);
or U21952 (N_21952,N_15129,N_12776);
and U21953 (N_21953,N_15200,N_16303);
nor U21954 (N_21954,N_16450,N_15864);
nand U21955 (N_21955,N_16355,N_14711);
or U21956 (N_21956,N_14702,N_13253);
or U21957 (N_21957,N_17421,N_13094);
and U21958 (N_21958,N_17821,N_15118);
or U21959 (N_21959,N_17165,N_13571);
or U21960 (N_21960,N_12121,N_13230);
nor U21961 (N_21961,N_12485,N_16556);
or U21962 (N_21962,N_14276,N_13589);
and U21963 (N_21963,N_17225,N_16592);
nand U21964 (N_21964,N_12292,N_12016);
nand U21965 (N_21965,N_12170,N_15809);
or U21966 (N_21966,N_12064,N_15611);
nor U21967 (N_21967,N_15122,N_13700);
nor U21968 (N_21968,N_14843,N_15984);
xnor U21969 (N_21969,N_12538,N_14610);
and U21970 (N_21970,N_16882,N_13961);
nor U21971 (N_21971,N_12258,N_12484);
and U21972 (N_21972,N_14146,N_15404);
xor U21973 (N_21973,N_17867,N_17530);
xnor U21974 (N_21974,N_17840,N_12937);
nand U21975 (N_21975,N_15770,N_12601);
nand U21976 (N_21976,N_16751,N_17763);
nand U21977 (N_21977,N_15040,N_16477);
or U21978 (N_21978,N_15814,N_17548);
nand U21979 (N_21979,N_16192,N_15819);
nand U21980 (N_21980,N_12759,N_15095);
nor U21981 (N_21981,N_13499,N_16795);
nor U21982 (N_21982,N_16622,N_17717);
and U21983 (N_21983,N_17077,N_12159);
and U21984 (N_21984,N_15762,N_14283);
and U21985 (N_21985,N_17840,N_16531);
nor U21986 (N_21986,N_14995,N_12173);
nor U21987 (N_21987,N_14906,N_16618);
nor U21988 (N_21988,N_16125,N_12400);
or U21989 (N_21989,N_12691,N_15591);
nand U21990 (N_21990,N_15494,N_13305);
nand U21991 (N_21991,N_12363,N_16880);
nor U21992 (N_21992,N_14577,N_14189);
nand U21993 (N_21993,N_15413,N_15229);
xnor U21994 (N_21994,N_13417,N_17612);
nand U21995 (N_21995,N_17817,N_16119);
or U21996 (N_21996,N_12266,N_16138);
nand U21997 (N_21997,N_16576,N_12891);
or U21998 (N_21998,N_17390,N_15137);
and U21999 (N_21999,N_12475,N_12520);
and U22000 (N_22000,N_16858,N_13769);
xnor U22001 (N_22001,N_15320,N_15338);
nand U22002 (N_22002,N_12068,N_15248);
nand U22003 (N_22003,N_14460,N_16399);
nand U22004 (N_22004,N_17693,N_17845);
nor U22005 (N_22005,N_16152,N_13128);
and U22006 (N_22006,N_15854,N_17933);
nand U22007 (N_22007,N_17078,N_13248);
and U22008 (N_22008,N_15033,N_17031);
xnor U22009 (N_22009,N_13828,N_17727);
and U22010 (N_22010,N_17906,N_12303);
xor U22011 (N_22011,N_14204,N_12045);
or U22012 (N_22012,N_16507,N_17138);
nand U22013 (N_22013,N_17225,N_16354);
nor U22014 (N_22014,N_14180,N_13731);
nor U22015 (N_22015,N_16207,N_15565);
nand U22016 (N_22016,N_17634,N_13511);
xnor U22017 (N_22017,N_15420,N_17053);
and U22018 (N_22018,N_16698,N_13722);
or U22019 (N_22019,N_17062,N_17975);
nand U22020 (N_22020,N_17145,N_14672);
or U22021 (N_22021,N_14090,N_14613);
nor U22022 (N_22022,N_17100,N_12809);
and U22023 (N_22023,N_16955,N_15082);
xor U22024 (N_22024,N_17924,N_12014);
nand U22025 (N_22025,N_12295,N_15019);
nor U22026 (N_22026,N_15414,N_17099);
nand U22027 (N_22027,N_12256,N_12528);
nor U22028 (N_22028,N_12991,N_13555);
or U22029 (N_22029,N_14904,N_13566);
nand U22030 (N_22030,N_15437,N_14773);
nand U22031 (N_22031,N_12699,N_13987);
xor U22032 (N_22032,N_13307,N_14901);
nor U22033 (N_22033,N_15866,N_16021);
nor U22034 (N_22034,N_16191,N_14470);
nand U22035 (N_22035,N_14806,N_14210);
or U22036 (N_22036,N_12890,N_17631);
nor U22037 (N_22037,N_16923,N_13634);
or U22038 (N_22038,N_15876,N_12326);
and U22039 (N_22039,N_14479,N_12695);
nand U22040 (N_22040,N_14059,N_16322);
xor U22041 (N_22041,N_17731,N_13516);
nor U22042 (N_22042,N_14535,N_14875);
and U22043 (N_22043,N_17133,N_16549);
nand U22044 (N_22044,N_16073,N_16150);
xor U22045 (N_22045,N_15787,N_13827);
xor U22046 (N_22046,N_12109,N_16965);
nor U22047 (N_22047,N_12406,N_14717);
nor U22048 (N_22048,N_12603,N_14506);
nor U22049 (N_22049,N_12642,N_16745);
xnor U22050 (N_22050,N_12848,N_17785);
nor U22051 (N_22051,N_13142,N_12504);
and U22052 (N_22052,N_12959,N_17929);
nand U22053 (N_22053,N_12507,N_13211);
or U22054 (N_22054,N_16095,N_13353);
nand U22055 (N_22055,N_14485,N_16731);
nand U22056 (N_22056,N_17969,N_12773);
or U22057 (N_22057,N_15451,N_15176);
nor U22058 (N_22058,N_12039,N_16973);
or U22059 (N_22059,N_15403,N_17131);
nand U22060 (N_22060,N_16521,N_13723);
nor U22061 (N_22061,N_12878,N_12708);
xor U22062 (N_22062,N_14760,N_14008);
nor U22063 (N_22063,N_17099,N_15316);
nor U22064 (N_22064,N_15580,N_14434);
and U22065 (N_22065,N_17033,N_13003);
nor U22066 (N_22066,N_13942,N_15470);
nor U22067 (N_22067,N_17244,N_14103);
nand U22068 (N_22068,N_15713,N_15839);
xor U22069 (N_22069,N_17833,N_16811);
and U22070 (N_22070,N_12224,N_12845);
nand U22071 (N_22071,N_12713,N_14682);
and U22072 (N_22072,N_13751,N_12505);
and U22073 (N_22073,N_13349,N_17594);
and U22074 (N_22074,N_17206,N_13543);
and U22075 (N_22075,N_15206,N_13103);
or U22076 (N_22076,N_12238,N_12104);
and U22077 (N_22077,N_13819,N_14968);
or U22078 (N_22078,N_15676,N_15690);
and U22079 (N_22079,N_12743,N_14830);
nand U22080 (N_22080,N_15154,N_12174);
nor U22081 (N_22081,N_17333,N_12300);
and U22082 (N_22082,N_13672,N_17644);
and U22083 (N_22083,N_14250,N_16809);
and U22084 (N_22084,N_16539,N_17907);
xor U22085 (N_22085,N_12767,N_17102);
xnor U22086 (N_22086,N_15022,N_15385);
or U22087 (N_22087,N_13185,N_14450);
or U22088 (N_22088,N_13297,N_14631);
nand U22089 (N_22089,N_17661,N_15326);
nand U22090 (N_22090,N_17152,N_15013);
or U22091 (N_22091,N_17608,N_16868);
xnor U22092 (N_22092,N_17630,N_17935);
nand U22093 (N_22093,N_16381,N_16798);
or U22094 (N_22094,N_15503,N_15574);
and U22095 (N_22095,N_14773,N_15563);
and U22096 (N_22096,N_13644,N_13492);
or U22097 (N_22097,N_16619,N_16942);
and U22098 (N_22098,N_17012,N_14068);
or U22099 (N_22099,N_12300,N_16426);
and U22100 (N_22100,N_16351,N_14740);
or U22101 (N_22101,N_17137,N_17529);
nand U22102 (N_22102,N_16073,N_13932);
and U22103 (N_22103,N_13201,N_16811);
xor U22104 (N_22104,N_14660,N_17786);
nor U22105 (N_22105,N_15717,N_13013);
nand U22106 (N_22106,N_16968,N_15286);
nor U22107 (N_22107,N_14528,N_16173);
and U22108 (N_22108,N_14641,N_15764);
or U22109 (N_22109,N_13124,N_13775);
or U22110 (N_22110,N_12854,N_15216);
and U22111 (N_22111,N_16985,N_13839);
nor U22112 (N_22112,N_17522,N_17519);
xor U22113 (N_22113,N_16253,N_14080);
nand U22114 (N_22114,N_17826,N_15375);
xor U22115 (N_22115,N_16555,N_14134);
nor U22116 (N_22116,N_16452,N_13389);
and U22117 (N_22117,N_16095,N_12927);
or U22118 (N_22118,N_13438,N_13813);
xnor U22119 (N_22119,N_14221,N_17496);
or U22120 (N_22120,N_14150,N_17040);
or U22121 (N_22121,N_12293,N_12673);
and U22122 (N_22122,N_12665,N_15415);
nor U22123 (N_22123,N_15482,N_14037);
and U22124 (N_22124,N_12244,N_12450);
and U22125 (N_22125,N_16538,N_12112);
nor U22126 (N_22126,N_17336,N_14497);
nor U22127 (N_22127,N_13727,N_12704);
nand U22128 (N_22128,N_12680,N_17437);
nand U22129 (N_22129,N_16701,N_16343);
and U22130 (N_22130,N_13425,N_14570);
nand U22131 (N_22131,N_15180,N_14101);
nand U22132 (N_22132,N_14302,N_15476);
xnor U22133 (N_22133,N_16982,N_12543);
or U22134 (N_22134,N_16095,N_17755);
or U22135 (N_22135,N_16183,N_15490);
or U22136 (N_22136,N_17617,N_12561);
or U22137 (N_22137,N_12517,N_17395);
nor U22138 (N_22138,N_14516,N_15502);
or U22139 (N_22139,N_14534,N_14928);
and U22140 (N_22140,N_17666,N_16025);
xnor U22141 (N_22141,N_16578,N_17598);
or U22142 (N_22142,N_16047,N_12272);
xor U22143 (N_22143,N_16352,N_15248);
nand U22144 (N_22144,N_16196,N_12525);
xor U22145 (N_22145,N_16514,N_17212);
or U22146 (N_22146,N_16078,N_12083);
and U22147 (N_22147,N_14905,N_17426);
or U22148 (N_22148,N_15353,N_13497);
nand U22149 (N_22149,N_15961,N_16606);
and U22150 (N_22150,N_12722,N_16850);
nand U22151 (N_22151,N_14505,N_14108);
nor U22152 (N_22152,N_15098,N_16336);
nand U22153 (N_22153,N_16917,N_17119);
nor U22154 (N_22154,N_12998,N_16570);
nand U22155 (N_22155,N_15338,N_13107);
nor U22156 (N_22156,N_15443,N_13119);
xnor U22157 (N_22157,N_15035,N_15447);
nor U22158 (N_22158,N_16533,N_15043);
nor U22159 (N_22159,N_13550,N_14003);
or U22160 (N_22160,N_14968,N_17888);
and U22161 (N_22161,N_17211,N_15095);
or U22162 (N_22162,N_13625,N_13526);
nand U22163 (N_22163,N_17395,N_16343);
or U22164 (N_22164,N_12711,N_14386);
or U22165 (N_22165,N_12686,N_13934);
nand U22166 (N_22166,N_15354,N_17376);
xor U22167 (N_22167,N_12984,N_16201);
or U22168 (N_22168,N_12533,N_14954);
nor U22169 (N_22169,N_15451,N_17124);
xor U22170 (N_22170,N_17535,N_12180);
xor U22171 (N_22171,N_17424,N_13241);
or U22172 (N_22172,N_13632,N_12266);
or U22173 (N_22173,N_17195,N_14727);
nor U22174 (N_22174,N_16653,N_15231);
xor U22175 (N_22175,N_12524,N_14860);
nand U22176 (N_22176,N_13062,N_13831);
nor U22177 (N_22177,N_13423,N_15945);
and U22178 (N_22178,N_14822,N_12505);
nand U22179 (N_22179,N_12028,N_16055);
xor U22180 (N_22180,N_13842,N_12854);
nor U22181 (N_22181,N_17721,N_15588);
and U22182 (N_22182,N_15002,N_17103);
xnor U22183 (N_22183,N_14060,N_17256);
nor U22184 (N_22184,N_13523,N_16297);
nor U22185 (N_22185,N_16781,N_15412);
or U22186 (N_22186,N_15839,N_13290);
and U22187 (N_22187,N_16317,N_17326);
or U22188 (N_22188,N_13576,N_17953);
nand U22189 (N_22189,N_15055,N_14531);
xor U22190 (N_22190,N_15252,N_17559);
nor U22191 (N_22191,N_13751,N_15402);
nand U22192 (N_22192,N_17504,N_17309);
nand U22193 (N_22193,N_13359,N_16439);
nor U22194 (N_22194,N_17273,N_13950);
nor U22195 (N_22195,N_15117,N_14707);
and U22196 (N_22196,N_13403,N_14744);
nand U22197 (N_22197,N_16693,N_15567);
nand U22198 (N_22198,N_15085,N_15067);
nor U22199 (N_22199,N_14611,N_16512);
nand U22200 (N_22200,N_15805,N_16855);
xor U22201 (N_22201,N_17211,N_16925);
and U22202 (N_22202,N_15902,N_15406);
nand U22203 (N_22203,N_15679,N_16149);
and U22204 (N_22204,N_12085,N_14183);
xnor U22205 (N_22205,N_12924,N_12159);
nand U22206 (N_22206,N_12111,N_16791);
nand U22207 (N_22207,N_14803,N_13578);
xor U22208 (N_22208,N_14906,N_16992);
and U22209 (N_22209,N_12779,N_17673);
and U22210 (N_22210,N_13155,N_15441);
and U22211 (N_22211,N_14348,N_17490);
nand U22212 (N_22212,N_12450,N_13177);
nand U22213 (N_22213,N_17782,N_17895);
and U22214 (N_22214,N_14857,N_14331);
and U22215 (N_22215,N_12410,N_17787);
or U22216 (N_22216,N_12894,N_13596);
nand U22217 (N_22217,N_14134,N_12876);
and U22218 (N_22218,N_13212,N_17432);
xnor U22219 (N_22219,N_14067,N_13768);
nand U22220 (N_22220,N_16891,N_16883);
nor U22221 (N_22221,N_14784,N_17469);
and U22222 (N_22222,N_16260,N_14339);
nand U22223 (N_22223,N_13048,N_14839);
nor U22224 (N_22224,N_13716,N_14708);
or U22225 (N_22225,N_15331,N_17741);
xor U22226 (N_22226,N_12996,N_14649);
nand U22227 (N_22227,N_15372,N_17490);
xnor U22228 (N_22228,N_16305,N_13241);
nand U22229 (N_22229,N_17404,N_17895);
and U22230 (N_22230,N_14451,N_12992);
and U22231 (N_22231,N_14330,N_15899);
nor U22232 (N_22232,N_13565,N_17072);
nor U22233 (N_22233,N_13021,N_13999);
or U22234 (N_22234,N_13597,N_16177);
or U22235 (N_22235,N_12495,N_17763);
nand U22236 (N_22236,N_14964,N_13217);
xnor U22237 (N_22237,N_13798,N_12374);
xor U22238 (N_22238,N_12088,N_16170);
and U22239 (N_22239,N_16639,N_14383);
or U22240 (N_22240,N_17434,N_17560);
xor U22241 (N_22241,N_16273,N_15513);
and U22242 (N_22242,N_12951,N_13008);
nand U22243 (N_22243,N_12768,N_12311);
nand U22244 (N_22244,N_13579,N_13135);
and U22245 (N_22245,N_15207,N_13702);
and U22246 (N_22246,N_13299,N_14744);
or U22247 (N_22247,N_14062,N_16912);
or U22248 (N_22248,N_15472,N_14173);
xnor U22249 (N_22249,N_12472,N_14030);
xor U22250 (N_22250,N_15190,N_12381);
nor U22251 (N_22251,N_12891,N_16726);
nand U22252 (N_22252,N_16404,N_12956);
nor U22253 (N_22253,N_15930,N_14492);
nand U22254 (N_22254,N_16437,N_13491);
xnor U22255 (N_22255,N_17252,N_13528);
xnor U22256 (N_22256,N_12280,N_17946);
xnor U22257 (N_22257,N_16493,N_12460);
nand U22258 (N_22258,N_16761,N_13731);
and U22259 (N_22259,N_15068,N_16508);
and U22260 (N_22260,N_17483,N_12357);
and U22261 (N_22261,N_14884,N_15588);
and U22262 (N_22262,N_16114,N_17661);
or U22263 (N_22263,N_16504,N_12890);
nand U22264 (N_22264,N_14044,N_16209);
or U22265 (N_22265,N_17328,N_17217);
xor U22266 (N_22266,N_15581,N_12205);
and U22267 (N_22267,N_15546,N_12727);
xnor U22268 (N_22268,N_13872,N_15280);
or U22269 (N_22269,N_17362,N_14574);
xnor U22270 (N_22270,N_14487,N_16168);
nor U22271 (N_22271,N_14799,N_12997);
xnor U22272 (N_22272,N_15950,N_16672);
nand U22273 (N_22273,N_17267,N_17806);
or U22274 (N_22274,N_14208,N_13681);
nand U22275 (N_22275,N_13699,N_14410);
nor U22276 (N_22276,N_14770,N_16242);
nor U22277 (N_22277,N_16060,N_12155);
and U22278 (N_22278,N_15732,N_12471);
nand U22279 (N_22279,N_17669,N_12416);
nor U22280 (N_22280,N_14572,N_16196);
nand U22281 (N_22281,N_14700,N_16202);
and U22282 (N_22282,N_14085,N_17319);
nand U22283 (N_22283,N_13805,N_12747);
xnor U22284 (N_22284,N_13854,N_13785);
nand U22285 (N_22285,N_17640,N_14608);
and U22286 (N_22286,N_14718,N_16008);
nor U22287 (N_22287,N_16300,N_12966);
and U22288 (N_22288,N_17800,N_12411);
nor U22289 (N_22289,N_14515,N_14569);
nor U22290 (N_22290,N_17643,N_14059);
nor U22291 (N_22291,N_17296,N_13259);
nor U22292 (N_22292,N_15096,N_17606);
or U22293 (N_22293,N_13686,N_17700);
xor U22294 (N_22294,N_14872,N_13680);
nand U22295 (N_22295,N_17076,N_12368);
xor U22296 (N_22296,N_16090,N_16433);
nor U22297 (N_22297,N_15185,N_15366);
nand U22298 (N_22298,N_15934,N_16239);
or U22299 (N_22299,N_15863,N_14058);
nand U22300 (N_22300,N_13104,N_13585);
and U22301 (N_22301,N_12347,N_14865);
nand U22302 (N_22302,N_13482,N_16692);
nor U22303 (N_22303,N_14390,N_16874);
and U22304 (N_22304,N_15788,N_17979);
nor U22305 (N_22305,N_13382,N_15004);
nand U22306 (N_22306,N_12438,N_15105);
or U22307 (N_22307,N_16787,N_17874);
or U22308 (N_22308,N_13337,N_12978);
nand U22309 (N_22309,N_14588,N_16342);
or U22310 (N_22310,N_13215,N_14976);
or U22311 (N_22311,N_13332,N_12289);
nand U22312 (N_22312,N_13100,N_14569);
nand U22313 (N_22313,N_12585,N_13882);
or U22314 (N_22314,N_12488,N_15122);
nand U22315 (N_22315,N_13717,N_13019);
nand U22316 (N_22316,N_17574,N_15962);
xnor U22317 (N_22317,N_14724,N_15967);
or U22318 (N_22318,N_13626,N_13866);
nand U22319 (N_22319,N_13910,N_14256);
xor U22320 (N_22320,N_13415,N_15207);
or U22321 (N_22321,N_14501,N_13948);
nor U22322 (N_22322,N_12652,N_12794);
and U22323 (N_22323,N_16936,N_17408);
nor U22324 (N_22324,N_16910,N_14421);
nor U22325 (N_22325,N_12242,N_14142);
nand U22326 (N_22326,N_15516,N_14899);
or U22327 (N_22327,N_15043,N_17586);
nor U22328 (N_22328,N_16935,N_14769);
and U22329 (N_22329,N_16823,N_15698);
or U22330 (N_22330,N_12821,N_13631);
and U22331 (N_22331,N_14642,N_17446);
or U22332 (N_22332,N_12781,N_15303);
nand U22333 (N_22333,N_17419,N_17840);
or U22334 (N_22334,N_12793,N_13729);
xor U22335 (N_22335,N_13573,N_16912);
and U22336 (N_22336,N_17849,N_14719);
nand U22337 (N_22337,N_17116,N_16024);
nor U22338 (N_22338,N_17748,N_12467);
and U22339 (N_22339,N_12697,N_12489);
xnor U22340 (N_22340,N_17252,N_12861);
nor U22341 (N_22341,N_12530,N_13480);
or U22342 (N_22342,N_14358,N_13095);
and U22343 (N_22343,N_17223,N_13268);
xnor U22344 (N_22344,N_14078,N_13645);
nand U22345 (N_22345,N_13955,N_15145);
or U22346 (N_22346,N_12787,N_13212);
xor U22347 (N_22347,N_15381,N_14954);
or U22348 (N_22348,N_16376,N_17654);
nand U22349 (N_22349,N_13056,N_16133);
or U22350 (N_22350,N_13444,N_14269);
and U22351 (N_22351,N_12682,N_12705);
nand U22352 (N_22352,N_13870,N_16426);
xor U22353 (N_22353,N_15557,N_15572);
xor U22354 (N_22354,N_13563,N_16560);
nand U22355 (N_22355,N_15283,N_12294);
xor U22356 (N_22356,N_14288,N_14924);
nand U22357 (N_22357,N_14366,N_14594);
and U22358 (N_22358,N_15760,N_15918);
nand U22359 (N_22359,N_16936,N_13448);
and U22360 (N_22360,N_17253,N_16831);
and U22361 (N_22361,N_13020,N_15391);
xnor U22362 (N_22362,N_12287,N_16407);
xnor U22363 (N_22363,N_16318,N_16972);
or U22364 (N_22364,N_12022,N_16208);
and U22365 (N_22365,N_17899,N_12460);
nor U22366 (N_22366,N_13599,N_13385);
nand U22367 (N_22367,N_12271,N_14578);
and U22368 (N_22368,N_13757,N_14107);
and U22369 (N_22369,N_12095,N_13632);
or U22370 (N_22370,N_13876,N_12384);
or U22371 (N_22371,N_16978,N_14467);
and U22372 (N_22372,N_15664,N_14559);
nor U22373 (N_22373,N_13519,N_14971);
xnor U22374 (N_22374,N_15197,N_13627);
xnor U22375 (N_22375,N_12455,N_15119);
xnor U22376 (N_22376,N_13441,N_16040);
xnor U22377 (N_22377,N_13153,N_13756);
nand U22378 (N_22378,N_12008,N_15709);
nand U22379 (N_22379,N_16783,N_15378);
xor U22380 (N_22380,N_16704,N_14400);
nor U22381 (N_22381,N_16898,N_13034);
or U22382 (N_22382,N_17608,N_13954);
nor U22383 (N_22383,N_14157,N_14962);
xnor U22384 (N_22384,N_12558,N_14823);
or U22385 (N_22385,N_15183,N_14787);
nand U22386 (N_22386,N_16473,N_17074);
or U22387 (N_22387,N_14662,N_12301);
or U22388 (N_22388,N_16413,N_14991);
xnor U22389 (N_22389,N_13056,N_17283);
or U22390 (N_22390,N_12453,N_17860);
xor U22391 (N_22391,N_15188,N_14270);
xnor U22392 (N_22392,N_14484,N_12165);
and U22393 (N_22393,N_14152,N_13093);
nand U22394 (N_22394,N_13128,N_16437);
nor U22395 (N_22395,N_16600,N_16314);
or U22396 (N_22396,N_17492,N_16012);
xnor U22397 (N_22397,N_15714,N_14370);
and U22398 (N_22398,N_12823,N_12455);
xor U22399 (N_22399,N_13655,N_14512);
and U22400 (N_22400,N_12401,N_14363);
or U22401 (N_22401,N_15521,N_14089);
nand U22402 (N_22402,N_15172,N_15805);
or U22403 (N_22403,N_13252,N_17154);
or U22404 (N_22404,N_14736,N_12301);
xnor U22405 (N_22405,N_12595,N_13917);
nand U22406 (N_22406,N_17474,N_16410);
nor U22407 (N_22407,N_12547,N_17739);
or U22408 (N_22408,N_17099,N_14446);
xor U22409 (N_22409,N_12733,N_13924);
and U22410 (N_22410,N_13368,N_13913);
and U22411 (N_22411,N_13478,N_15251);
or U22412 (N_22412,N_16476,N_16569);
or U22413 (N_22413,N_14519,N_14074);
or U22414 (N_22414,N_15245,N_15410);
and U22415 (N_22415,N_15902,N_14441);
and U22416 (N_22416,N_14470,N_13977);
and U22417 (N_22417,N_17680,N_16739);
xnor U22418 (N_22418,N_13434,N_16250);
nand U22419 (N_22419,N_16667,N_15806);
or U22420 (N_22420,N_14348,N_16418);
or U22421 (N_22421,N_17366,N_16570);
nand U22422 (N_22422,N_15315,N_12807);
xnor U22423 (N_22423,N_16158,N_15617);
xor U22424 (N_22424,N_17426,N_16879);
xnor U22425 (N_22425,N_17466,N_17991);
nor U22426 (N_22426,N_17003,N_12725);
and U22427 (N_22427,N_15115,N_15257);
nor U22428 (N_22428,N_14489,N_12147);
xnor U22429 (N_22429,N_15728,N_17236);
nand U22430 (N_22430,N_13639,N_15290);
xor U22431 (N_22431,N_17245,N_12231);
xor U22432 (N_22432,N_16144,N_13248);
and U22433 (N_22433,N_14190,N_15432);
xnor U22434 (N_22434,N_14539,N_14925);
nor U22435 (N_22435,N_15481,N_16697);
xor U22436 (N_22436,N_16128,N_16706);
or U22437 (N_22437,N_15234,N_12041);
xnor U22438 (N_22438,N_12074,N_16885);
or U22439 (N_22439,N_16666,N_14692);
xnor U22440 (N_22440,N_17982,N_16552);
or U22441 (N_22441,N_16504,N_14681);
nand U22442 (N_22442,N_12346,N_14709);
xnor U22443 (N_22443,N_12275,N_15261);
xor U22444 (N_22444,N_15721,N_12338);
nand U22445 (N_22445,N_14392,N_14448);
nor U22446 (N_22446,N_14738,N_13239);
nand U22447 (N_22447,N_13501,N_14711);
or U22448 (N_22448,N_15890,N_12581);
or U22449 (N_22449,N_13568,N_17016);
nor U22450 (N_22450,N_12079,N_12746);
xor U22451 (N_22451,N_15139,N_14023);
nor U22452 (N_22452,N_15906,N_16253);
nor U22453 (N_22453,N_16849,N_16651);
nor U22454 (N_22454,N_16998,N_14843);
nand U22455 (N_22455,N_13540,N_13284);
xor U22456 (N_22456,N_12781,N_15668);
nand U22457 (N_22457,N_16551,N_15342);
and U22458 (N_22458,N_17061,N_17085);
and U22459 (N_22459,N_17137,N_17378);
or U22460 (N_22460,N_13653,N_15727);
nand U22461 (N_22461,N_12566,N_17702);
and U22462 (N_22462,N_16130,N_13796);
and U22463 (N_22463,N_14295,N_14511);
nand U22464 (N_22464,N_16107,N_17530);
nand U22465 (N_22465,N_14758,N_16356);
or U22466 (N_22466,N_14321,N_12213);
xor U22467 (N_22467,N_17852,N_17324);
nand U22468 (N_22468,N_13875,N_15115);
xnor U22469 (N_22469,N_14488,N_14045);
and U22470 (N_22470,N_14770,N_16863);
xnor U22471 (N_22471,N_17411,N_13023);
or U22472 (N_22472,N_12675,N_15815);
nand U22473 (N_22473,N_16081,N_14618);
nor U22474 (N_22474,N_16404,N_17226);
xor U22475 (N_22475,N_12942,N_16967);
or U22476 (N_22476,N_14074,N_12873);
xor U22477 (N_22477,N_16123,N_13241);
nor U22478 (N_22478,N_14767,N_13569);
or U22479 (N_22479,N_17965,N_14129);
or U22480 (N_22480,N_14726,N_17948);
nor U22481 (N_22481,N_12544,N_14968);
nor U22482 (N_22482,N_12583,N_16125);
nor U22483 (N_22483,N_16528,N_15354);
nor U22484 (N_22484,N_13164,N_14368);
nor U22485 (N_22485,N_16317,N_13166);
or U22486 (N_22486,N_13394,N_14930);
and U22487 (N_22487,N_17940,N_15298);
nor U22488 (N_22488,N_13207,N_15567);
nor U22489 (N_22489,N_15951,N_17355);
nand U22490 (N_22490,N_17032,N_16034);
nor U22491 (N_22491,N_12368,N_13348);
nand U22492 (N_22492,N_17553,N_12332);
and U22493 (N_22493,N_16848,N_12504);
nor U22494 (N_22494,N_13137,N_15595);
nor U22495 (N_22495,N_14999,N_16938);
nor U22496 (N_22496,N_17555,N_14965);
nand U22497 (N_22497,N_17741,N_13379);
and U22498 (N_22498,N_16154,N_16260);
nor U22499 (N_22499,N_12668,N_15325);
nor U22500 (N_22500,N_17512,N_12964);
nor U22501 (N_22501,N_14138,N_15042);
nor U22502 (N_22502,N_15009,N_17004);
or U22503 (N_22503,N_15232,N_15460);
or U22504 (N_22504,N_15827,N_17548);
nand U22505 (N_22505,N_16904,N_17053);
nand U22506 (N_22506,N_13808,N_13246);
and U22507 (N_22507,N_12443,N_12969);
xnor U22508 (N_22508,N_12805,N_15998);
xor U22509 (N_22509,N_16157,N_12534);
xor U22510 (N_22510,N_15347,N_15248);
xor U22511 (N_22511,N_16576,N_15561);
nand U22512 (N_22512,N_17997,N_14870);
or U22513 (N_22513,N_17988,N_14653);
xor U22514 (N_22514,N_17848,N_14082);
or U22515 (N_22515,N_17891,N_13783);
xor U22516 (N_22516,N_14608,N_13682);
and U22517 (N_22517,N_13920,N_14754);
xnor U22518 (N_22518,N_16139,N_12528);
nand U22519 (N_22519,N_17902,N_14587);
nor U22520 (N_22520,N_16641,N_17056);
and U22521 (N_22521,N_17433,N_17247);
or U22522 (N_22522,N_15088,N_17248);
or U22523 (N_22523,N_15410,N_17989);
nand U22524 (N_22524,N_14822,N_16226);
or U22525 (N_22525,N_12293,N_14515);
nor U22526 (N_22526,N_16381,N_15539);
xnor U22527 (N_22527,N_14809,N_16697);
and U22528 (N_22528,N_16089,N_17930);
nand U22529 (N_22529,N_16335,N_12449);
xnor U22530 (N_22530,N_16638,N_13646);
and U22531 (N_22531,N_16718,N_15179);
xnor U22532 (N_22532,N_14470,N_17363);
and U22533 (N_22533,N_16854,N_14339);
xor U22534 (N_22534,N_13281,N_13886);
nor U22535 (N_22535,N_14949,N_16838);
or U22536 (N_22536,N_14771,N_15465);
or U22537 (N_22537,N_12007,N_13337);
xor U22538 (N_22538,N_15071,N_17658);
or U22539 (N_22539,N_16164,N_13960);
nor U22540 (N_22540,N_13848,N_16423);
nor U22541 (N_22541,N_17578,N_12409);
and U22542 (N_22542,N_14305,N_14153);
nand U22543 (N_22543,N_13875,N_15336);
nand U22544 (N_22544,N_12816,N_14276);
or U22545 (N_22545,N_17492,N_16773);
and U22546 (N_22546,N_13079,N_17826);
xor U22547 (N_22547,N_17388,N_14749);
or U22548 (N_22548,N_16366,N_15843);
nand U22549 (N_22549,N_13369,N_17985);
nor U22550 (N_22550,N_16568,N_12372);
nand U22551 (N_22551,N_12205,N_15544);
and U22552 (N_22552,N_13723,N_12106);
nand U22553 (N_22553,N_17696,N_15395);
xor U22554 (N_22554,N_17687,N_16503);
and U22555 (N_22555,N_15643,N_13610);
and U22556 (N_22556,N_12628,N_16355);
nand U22557 (N_22557,N_13321,N_17807);
nand U22558 (N_22558,N_17979,N_15171);
and U22559 (N_22559,N_12510,N_12081);
xor U22560 (N_22560,N_16800,N_14075);
nand U22561 (N_22561,N_14432,N_17343);
nor U22562 (N_22562,N_17931,N_16880);
nand U22563 (N_22563,N_12948,N_16607);
nor U22564 (N_22564,N_16207,N_17654);
nor U22565 (N_22565,N_14524,N_16967);
and U22566 (N_22566,N_16512,N_17303);
nand U22567 (N_22567,N_17499,N_13175);
xnor U22568 (N_22568,N_15069,N_14693);
xnor U22569 (N_22569,N_15246,N_16250);
or U22570 (N_22570,N_12624,N_12412);
nor U22571 (N_22571,N_16742,N_12742);
or U22572 (N_22572,N_17676,N_13142);
nor U22573 (N_22573,N_12241,N_16766);
and U22574 (N_22574,N_16428,N_13898);
xor U22575 (N_22575,N_12807,N_16074);
nor U22576 (N_22576,N_15782,N_15661);
nor U22577 (N_22577,N_13543,N_12398);
and U22578 (N_22578,N_14730,N_17571);
xnor U22579 (N_22579,N_16950,N_17955);
and U22580 (N_22580,N_12935,N_16368);
or U22581 (N_22581,N_12170,N_15104);
or U22582 (N_22582,N_17215,N_15664);
or U22583 (N_22583,N_16886,N_17182);
xor U22584 (N_22584,N_15116,N_16720);
xor U22585 (N_22585,N_17362,N_12246);
nand U22586 (N_22586,N_12897,N_17841);
nor U22587 (N_22587,N_14853,N_17643);
xor U22588 (N_22588,N_12441,N_15415);
nand U22589 (N_22589,N_13782,N_13137);
nor U22590 (N_22590,N_13274,N_12063);
nor U22591 (N_22591,N_15589,N_15643);
and U22592 (N_22592,N_17335,N_15210);
nor U22593 (N_22593,N_13188,N_14815);
xnor U22594 (N_22594,N_17197,N_17851);
nand U22595 (N_22595,N_17223,N_15391);
or U22596 (N_22596,N_13364,N_13161);
nor U22597 (N_22597,N_17002,N_13808);
nand U22598 (N_22598,N_14284,N_16699);
xnor U22599 (N_22599,N_14854,N_17153);
nor U22600 (N_22600,N_17930,N_12402);
nor U22601 (N_22601,N_17195,N_16877);
and U22602 (N_22602,N_16664,N_14434);
xnor U22603 (N_22603,N_17596,N_13950);
nand U22604 (N_22604,N_16823,N_14687);
nand U22605 (N_22605,N_12666,N_12023);
and U22606 (N_22606,N_14863,N_16426);
nor U22607 (N_22607,N_13423,N_14918);
nor U22608 (N_22608,N_12851,N_17815);
nor U22609 (N_22609,N_16421,N_15248);
xor U22610 (N_22610,N_14237,N_13044);
and U22611 (N_22611,N_17897,N_17943);
nand U22612 (N_22612,N_17873,N_16726);
xor U22613 (N_22613,N_13090,N_13079);
or U22614 (N_22614,N_12952,N_15180);
xor U22615 (N_22615,N_13367,N_14680);
nor U22616 (N_22616,N_13885,N_17805);
and U22617 (N_22617,N_16498,N_15900);
and U22618 (N_22618,N_16870,N_16564);
or U22619 (N_22619,N_17068,N_15091);
and U22620 (N_22620,N_16002,N_12538);
or U22621 (N_22621,N_14778,N_12388);
nor U22622 (N_22622,N_17476,N_16195);
nand U22623 (N_22623,N_13961,N_16932);
nand U22624 (N_22624,N_14407,N_15498);
and U22625 (N_22625,N_12427,N_12813);
xnor U22626 (N_22626,N_17135,N_17095);
and U22627 (N_22627,N_12931,N_12968);
nand U22628 (N_22628,N_14228,N_13457);
or U22629 (N_22629,N_15267,N_15907);
xor U22630 (N_22630,N_14684,N_13362);
nor U22631 (N_22631,N_15043,N_15754);
and U22632 (N_22632,N_13039,N_15572);
xnor U22633 (N_22633,N_15288,N_17093);
or U22634 (N_22634,N_13531,N_13450);
nor U22635 (N_22635,N_15496,N_14737);
and U22636 (N_22636,N_12135,N_16838);
nor U22637 (N_22637,N_15087,N_17383);
nor U22638 (N_22638,N_15682,N_16941);
or U22639 (N_22639,N_15479,N_14595);
and U22640 (N_22640,N_12668,N_13682);
and U22641 (N_22641,N_15822,N_12662);
nor U22642 (N_22642,N_16046,N_12328);
xnor U22643 (N_22643,N_16973,N_14389);
or U22644 (N_22644,N_16882,N_17163);
xor U22645 (N_22645,N_17857,N_15118);
nor U22646 (N_22646,N_16424,N_17676);
or U22647 (N_22647,N_14390,N_14856);
xnor U22648 (N_22648,N_13935,N_13491);
and U22649 (N_22649,N_17641,N_12383);
nor U22650 (N_22650,N_12956,N_16491);
xnor U22651 (N_22651,N_13182,N_14992);
nor U22652 (N_22652,N_12895,N_14573);
or U22653 (N_22653,N_12145,N_13286);
or U22654 (N_22654,N_16438,N_14499);
or U22655 (N_22655,N_17330,N_14062);
and U22656 (N_22656,N_16378,N_13388);
and U22657 (N_22657,N_13797,N_14777);
or U22658 (N_22658,N_14795,N_14285);
nand U22659 (N_22659,N_12988,N_17737);
nand U22660 (N_22660,N_12594,N_14488);
and U22661 (N_22661,N_15897,N_12587);
nor U22662 (N_22662,N_14566,N_12797);
nor U22663 (N_22663,N_16189,N_17501);
and U22664 (N_22664,N_16037,N_12455);
xnor U22665 (N_22665,N_14809,N_12538);
nand U22666 (N_22666,N_16260,N_15065);
nand U22667 (N_22667,N_16185,N_16144);
nor U22668 (N_22668,N_15872,N_13974);
nand U22669 (N_22669,N_17755,N_14500);
and U22670 (N_22670,N_14797,N_17422);
or U22671 (N_22671,N_17844,N_15259);
or U22672 (N_22672,N_13327,N_14266);
nor U22673 (N_22673,N_13220,N_15005);
nor U22674 (N_22674,N_16251,N_13766);
xnor U22675 (N_22675,N_12559,N_12387);
nor U22676 (N_22676,N_15460,N_13672);
nand U22677 (N_22677,N_17396,N_15973);
xnor U22678 (N_22678,N_15299,N_13340);
nand U22679 (N_22679,N_15184,N_15585);
nand U22680 (N_22680,N_13379,N_14619);
nor U22681 (N_22681,N_15611,N_14683);
and U22682 (N_22682,N_17321,N_16232);
or U22683 (N_22683,N_12986,N_13495);
nor U22684 (N_22684,N_17947,N_15286);
nand U22685 (N_22685,N_15225,N_13963);
xnor U22686 (N_22686,N_14061,N_16953);
xor U22687 (N_22687,N_13932,N_15063);
nand U22688 (N_22688,N_16533,N_16865);
nand U22689 (N_22689,N_17710,N_14533);
nor U22690 (N_22690,N_15004,N_15444);
nor U22691 (N_22691,N_15731,N_12681);
nor U22692 (N_22692,N_14490,N_17232);
nand U22693 (N_22693,N_12754,N_16921);
nor U22694 (N_22694,N_12346,N_12124);
xor U22695 (N_22695,N_13033,N_12344);
xnor U22696 (N_22696,N_13844,N_13552);
nor U22697 (N_22697,N_17304,N_12100);
xnor U22698 (N_22698,N_17680,N_13837);
nand U22699 (N_22699,N_16671,N_15337);
nor U22700 (N_22700,N_13071,N_12864);
and U22701 (N_22701,N_14782,N_15267);
nor U22702 (N_22702,N_13317,N_14041);
xnor U22703 (N_22703,N_12653,N_14819);
xnor U22704 (N_22704,N_13002,N_14732);
nand U22705 (N_22705,N_12296,N_13141);
or U22706 (N_22706,N_14171,N_16985);
xor U22707 (N_22707,N_14472,N_12696);
xnor U22708 (N_22708,N_17536,N_16663);
or U22709 (N_22709,N_13160,N_13994);
nand U22710 (N_22710,N_13335,N_13426);
nand U22711 (N_22711,N_17175,N_14862);
nor U22712 (N_22712,N_15179,N_14884);
and U22713 (N_22713,N_14585,N_13651);
nand U22714 (N_22714,N_15329,N_17462);
nand U22715 (N_22715,N_14712,N_13927);
or U22716 (N_22716,N_12691,N_13678);
or U22717 (N_22717,N_16217,N_13116);
nor U22718 (N_22718,N_17964,N_13299);
nor U22719 (N_22719,N_13379,N_15941);
nor U22720 (N_22720,N_15255,N_16863);
or U22721 (N_22721,N_15802,N_16663);
or U22722 (N_22722,N_12158,N_16117);
nor U22723 (N_22723,N_13728,N_14236);
or U22724 (N_22724,N_17030,N_12644);
xnor U22725 (N_22725,N_15344,N_17379);
and U22726 (N_22726,N_15760,N_13901);
xor U22727 (N_22727,N_14698,N_13639);
or U22728 (N_22728,N_17748,N_13047);
or U22729 (N_22729,N_12710,N_15585);
xnor U22730 (N_22730,N_16844,N_17996);
and U22731 (N_22731,N_16102,N_15787);
xnor U22732 (N_22732,N_16159,N_15817);
and U22733 (N_22733,N_13481,N_14755);
or U22734 (N_22734,N_13423,N_16854);
nor U22735 (N_22735,N_13248,N_12723);
and U22736 (N_22736,N_16203,N_16773);
xor U22737 (N_22737,N_17117,N_13168);
xnor U22738 (N_22738,N_17525,N_13522);
nor U22739 (N_22739,N_13657,N_14499);
and U22740 (N_22740,N_15275,N_15155);
nor U22741 (N_22741,N_14466,N_14144);
nand U22742 (N_22742,N_17601,N_12426);
and U22743 (N_22743,N_14089,N_13652);
and U22744 (N_22744,N_15490,N_12515);
xnor U22745 (N_22745,N_13147,N_12867);
or U22746 (N_22746,N_15877,N_15355);
or U22747 (N_22747,N_12849,N_14557);
nand U22748 (N_22748,N_15816,N_13149);
xnor U22749 (N_22749,N_12378,N_14414);
or U22750 (N_22750,N_15260,N_12744);
xor U22751 (N_22751,N_13107,N_17049);
xor U22752 (N_22752,N_16575,N_14886);
and U22753 (N_22753,N_12662,N_17270);
nor U22754 (N_22754,N_17077,N_14630);
xnor U22755 (N_22755,N_13628,N_16811);
nor U22756 (N_22756,N_16203,N_13960);
nor U22757 (N_22757,N_14890,N_17021);
nor U22758 (N_22758,N_16290,N_13665);
nor U22759 (N_22759,N_14180,N_12841);
xnor U22760 (N_22760,N_13313,N_16009);
xnor U22761 (N_22761,N_14774,N_13764);
and U22762 (N_22762,N_13861,N_17381);
nand U22763 (N_22763,N_16837,N_12747);
xor U22764 (N_22764,N_12533,N_13505);
nand U22765 (N_22765,N_13706,N_12604);
and U22766 (N_22766,N_17659,N_16510);
and U22767 (N_22767,N_12578,N_14098);
nor U22768 (N_22768,N_14139,N_14380);
nand U22769 (N_22769,N_14514,N_13675);
nor U22770 (N_22770,N_16277,N_16052);
nor U22771 (N_22771,N_13464,N_14539);
xor U22772 (N_22772,N_17503,N_13320);
nand U22773 (N_22773,N_13596,N_17262);
nor U22774 (N_22774,N_14948,N_14083);
and U22775 (N_22775,N_17186,N_17625);
and U22776 (N_22776,N_16464,N_13994);
nand U22777 (N_22777,N_12529,N_13018);
nor U22778 (N_22778,N_17605,N_16245);
or U22779 (N_22779,N_13798,N_12717);
nand U22780 (N_22780,N_15626,N_15813);
or U22781 (N_22781,N_16162,N_14113);
nor U22782 (N_22782,N_16894,N_13179);
nor U22783 (N_22783,N_13118,N_15203);
and U22784 (N_22784,N_13309,N_17069);
nor U22785 (N_22785,N_12315,N_12690);
nand U22786 (N_22786,N_13894,N_13587);
or U22787 (N_22787,N_16614,N_15345);
nand U22788 (N_22788,N_17030,N_14090);
xnor U22789 (N_22789,N_14189,N_16002);
nor U22790 (N_22790,N_13127,N_12318);
or U22791 (N_22791,N_16261,N_14978);
xor U22792 (N_22792,N_17854,N_17623);
xnor U22793 (N_22793,N_14275,N_16878);
and U22794 (N_22794,N_13818,N_13361);
xnor U22795 (N_22795,N_17302,N_15314);
nand U22796 (N_22796,N_13641,N_12571);
and U22797 (N_22797,N_16635,N_16737);
nand U22798 (N_22798,N_17738,N_13410);
nor U22799 (N_22799,N_16293,N_13602);
and U22800 (N_22800,N_13501,N_14987);
nand U22801 (N_22801,N_17646,N_13884);
or U22802 (N_22802,N_14554,N_13134);
nor U22803 (N_22803,N_13020,N_12415);
nor U22804 (N_22804,N_17971,N_12743);
and U22805 (N_22805,N_14513,N_15701);
or U22806 (N_22806,N_14623,N_15882);
nor U22807 (N_22807,N_15125,N_12962);
or U22808 (N_22808,N_15060,N_13965);
or U22809 (N_22809,N_12519,N_14480);
nand U22810 (N_22810,N_15855,N_12295);
or U22811 (N_22811,N_14757,N_13800);
xnor U22812 (N_22812,N_16429,N_14223);
or U22813 (N_22813,N_12432,N_14361);
or U22814 (N_22814,N_16603,N_12122);
or U22815 (N_22815,N_15636,N_14644);
xor U22816 (N_22816,N_14810,N_12246);
nor U22817 (N_22817,N_16029,N_17638);
xor U22818 (N_22818,N_13515,N_17407);
nor U22819 (N_22819,N_12425,N_14524);
nand U22820 (N_22820,N_14742,N_13663);
xnor U22821 (N_22821,N_13789,N_15585);
or U22822 (N_22822,N_12151,N_13082);
xor U22823 (N_22823,N_17526,N_17629);
nand U22824 (N_22824,N_12052,N_12656);
or U22825 (N_22825,N_12216,N_15889);
nor U22826 (N_22826,N_17239,N_12180);
and U22827 (N_22827,N_15284,N_14254);
and U22828 (N_22828,N_12280,N_13546);
nor U22829 (N_22829,N_13010,N_14394);
and U22830 (N_22830,N_15547,N_17725);
or U22831 (N_22831,N_12006,N_12972);
nor U22832 (N_22832,N_15074,N_12031);
or U22833 (N_22833,N_14395,N_15145);
and U22834 (N_22834,N_15985,N_15193);
nand U22835 (N_22835,N_13810,N_13303);
or U22836 (N_22836,N_17721,N_13449);
and U22837 (N_22837,N_16975,N_12415);
xor U22838 (N_22838,N_14667,N_15748);
nor U22839 (N_22839,N_12215,N_13467);
nand U22840 (N_22840,N_14302,N_14834);
xnor U22841 (N_22841,N_14607,N_15887);
nand U22842 (N_22842,N_12662,N_13764);
nand U22843 (N_22843,N_16725,N_15192);
or U22844 (N_22844,N_12058,N_14493);
nand U22845 (N_22845,N_16803,N_16387);
xnor U22846 (N_22846,N_17949,N_14441);
and U22847 (N_22847,N_17726,N_13081);
nand U22848 (N_22848,N_16809,N_15821);
and U22849 (N_22849,N_15907,N_15125);
and U22850 (N_22850,N_13815,N_17453);
xnor U22851 (N_22851,N_16327,N_13862);
or U22852 (N_22852,N_15522,N_16080);
and U22853 (N_22853,N_17877,N_12402);
and U22854 (N_22854,N_17565,N_14475);
or U22855 (N_22855,N_17559,N_15815);
and U22856 (N_22856,N_15239,N_13862);
nand U22857 (N_22857,N_17741,N_16397);
xnor U22858 (N_22858,N_17323,N_14984);
and U22859 (N_22859,N_14435,N_16621);
nand U22860 (N_22860,N_14403,N_14069);
nand U22861 (N_22861,N_17836,N_15495);
nand U22862 (N_22862,N_14483,N_16875);
xnor U22863 (N_22863,N_16603,N_17173);
nor U22864 (N_22864,N_13581,N_16659);
xor U22865 (N_22865,N_13477,N_13106);
or U22866 (N_22866,N_17794,N_17581);
nor U22867 (N_22867,N_13628,N_15919);
xor U22868 (N_22868,N_14931,N_16969);
nor U22869 (N_22869,N_17618,N_16943);
or U22870 (N_22870,N_15111,N_15146);
nor U22871 (N_22871,N_14332,N_17536);
xor U22872 (N_22872,N_13445,N_17669);
and U22873 (N_22873,N_13093,N_13275);
nand U22874 (N_22874,N_16910,N_13298);
nor U22875 (N_22875,N_15302,N_16846);
and U22876 (N_22876,N_12719,N_14882);
and U22877 (N_22877,N_17666,N_15047);
and U22878 (N_22878,N_17509,N_16878);
nand U22879 (N_22879,N_12446,N_14331);
nor U22880 (N_22880,N_17427,N_14473);
xnor U22881 (N_22881,N_16283,N_16596);
xor U22882 (N_22882,N_14234,N_12270);
xnor U22883 (N_22883,N_14063,N_16669);
and U22884 (N_22884,N_13977,N_12919);
nand U22885 (N_22885,N_16611,N_12997);
nand U22886 (N_22886,N_14672,N_14352);
nand U22887 (N_22887,N_17520,N_15466);
or U22888 (N_22888,N_15953,N_17605);
and U22889 (N_22889,N_17207,N_17446);
nor U22890 (N_22890,N_15850,N_17857);
and U22891 (N_22891,N_13615,N_12419);
and U22892 (N_22892,N_12489,N_17778);
or U22893 (N_22893,N_17521,N_13533);
nor U22894 (N_22894,N_14620,N_13345);
nor U22895 (N_22895,N_15062,N_13489);
and U22896 (N_22896,N_13571,N_17761);
or U22897 (N_22897,N_15636,N_16773);
nand U22898 (N_22898,N_13737,N_12993);
or U22899 (N_22899,N_13183,N_12017);
nand U22900 (N_22900,N_16216,N_13983);
and U22901 (N_22901,N_15008,N_16532);
xnor U22902 (N_22902,N_17135,N_12057);
and U22903 (N_22903,N_13025,N_12026);
nand U22904 (N_22904,N_13760,N_16700);
and U22905 (N_22905,N_13861,N_12166);
or U22906 (N_22906,N_16693,N_12820);
or U22907 (N_22907,N_16632,N_13772);
and U22908 (N_22908,N_17994,N_13436);
nor U22909 (N_22909,N_15209,N_14502);
and U22910 (N_22910,N_14157,N_12243);
nor U22911 (N_22911,N_12745,N_12085);
xor U22912 (N_22912,N_15379,N_14022);
xor U22913 (N_22913,N_12478,N_12952);
xnor U22914 (N_22914,N_15511,N_16191);
xor U22915 (N_22915,N_14332,N_12863);
nor U22916 (N_22916,N_17086,N_13313);
and U22917 (N_22917,N_17491,N_14347);
or U22918 (N_22918,N_16395,N_12763);
and U22919 (N_22919,N_14438,N_15954);
xnor U22920 (N_22920,N_14290,N_17001);
or U22921 (N_22921,N_13806,N_12958);
or U22922 (N_22922,N_14383,N_12550);
nand U22923 (N_22923,N_17325,N_12293);
or U22924 (N_22924,N_13747,N_15952);
and U22925 (N_22925,N_16788,N_17508);
nor U22926 (N_22926,N_16539,N_17923);
xnor U22927 (N_22927,N_13006,N_17858);
and U22928 (N_22928,N_15942,N_14920);
or U22929 (N_22929,N_15710,N_16246);
and U22930 (N_22930,N_15310,N_17695);
or U22931 (N_22931,N_13462,N_15039);
and U22932 (N_22932,N_13337,N_14404);
nand U22933 (N_22933,N_16503,N_13604);
nand U22934 (N_22934,N_14504,N_14376);
or U22935 (N_22935,N_17654,N_12969);
nand U22936 (N_22936,N_14163,N_13430);
and U22937 (N_22937,N_15749,N_16101);
nand U22938 (N_22938,N_13717,N_12421);
nand U22939 (N_22939,N_14388,N_17685);
and U22940 (N_22940,N_14111,N_16502);
or U22941 (N_22941,N_14861,N_14236);
nand U22942 (N_22942,N_17867,N_12138);
nand U22943 (N_22943,N_17139,N_14469);
nor U22944 (N_22944,N_12861,N_13349);
nor U22945 (N_22945,N_16185,N_15679);
nor U22946 (N_22946,N_13943,N_16540);
xor U22947 (N_22947,N_13028,N_17787);
or U22948 (N_22948,N_15222,N_17157);
xor U22949 (N_22949,N_16917,N_12433);
or U22950 (N_22950,N_12428,N_16850);
nor U22951 (N_22951,N_15000,N_15506);
or U22952 (N_22952,N_13840,N_16174);
nor U22953 (N_22953,N_14350,N_12853);
nand U22954 (N_22954,N_17450,N_17090);
xnor U22955 (N_22955,N_15078,N_15503);
or U22956 (N_22956,N_15688,N_14369);
nand U22957 (N_22957,N_12859,N_15236);
and U22958 (N_22958,N_16481,N_17889);
xor U22959 (N_22959,N_15069,N_15008);
and U22960 (N_22960,N_14536,N_14916);
nand U22961 (N_22961,N_15887,N_15632);
nand U22962 (N_22962,N_16456,N_12596);
and U22963 (N_22963,N_17070,N_12683);
or U22964 (N_22964,N_15204,N_14915);
and U22965 (N_22965,N_13327,N_15499);
and U22966 (N_22966,N_16705,N_17400);
and U22967 (N_22967,N_14445,N_17122);
or U22968 (N_22968,N_17505,N_16436);
nor U22969 (N_22969,N_12187,N_13220);
or U22970 (N_22970,N_13805,N_15949);
nor U22971 (N_22971,N_14498,N_13523);
nor U22972 (N_22972,N_12349,N_12718);
or U22973 (N_22973,N_15916,N_16439);
or U22974 (N_22974,N_15430,N_17315);
and U22975 (N_22975,N_17271,N_12338);
or U22976 (N_22976,N_14373,N_17985);
or U22977 (N_22977,N_12930,N_15512);
and U22978 (N_22978,N_15727,N_12551);
and U22979 (N_22979,N_15291,N_15703);
and U22980 (N_22980,N_12679,N_16404);
nand U22981 (N_22981,N_14821,N_15721);
or U22982 (N_22982,N_16970,N_13306);
nor U22983 (N_22983,N_13591,N_16552);
xnor U22984 (N_22984,N_12963,N_17334);
nor U22985 (N_22985,N_13189,N_12673);
and U22986 (N_22986,N_12374,N_17617);
xnor U22987 (N_22987,N_15905,N_17802);
xor U22988 (N_22988,N_15546,N_13881);
or U22989 (N_22989,N_13750,N_15679);
xnor U22990 (N_22990,N_16575,N_17932);
nor U22991 (N_22991,N_13295,N_15648);
or U22992 (N_22992,N_12741,N_13323);
or U22993 (N_22993,N_14285,N_13218);
nand U22994 (N_22994,N_16175,N_15586);
nand U22995 (N_22995,N_16187,N_14124);
or U22996 (N_22996,N_17355,N_12790);
nand U22997 (N_22997,N_17470,N_13731);
or U22998 (N_22998,N_15663,N_14007);
nor U22999 (N_22999,N_16835,N_15588);
nand U23000 (N_23000,N_16353,N_16562);
nand U23001 (N_23001,N_14553,N_13084);
nand U23002 (N_23002,N_15913,N_16710);
or U23003 (N_23003,N_16728,N_15025);
nand U23004 (N_23004,N_14900,N_15965);
nand U23005 (N_23005,N_14105,N_15005);
or U23006 (N_23006,N_16844,N_12997);
nand U23007 (N_23007,N_13101,N_13901);
nand U23008 (N_23008,N_17611,N_15523);
nand U23009 (N_23009,N_17481,N_17757);
and U23010 (N_23010,N_15432,N_15291);
or U23011 (N_23011,N_17748,N_12056);
and U23012 (N_23012,N_16736,N_13349);
nor U23013 (N_23013,N_16028,N_14281);
nor U23014 (N_23014,N_16533,N_14641);
nand U23015 (N_23015,N_12814,N_13805);
and U23016 (N_23016,N_15534,N_15409);
and U23017 (N_23017,N_13956,N_15723);
and U23018 (N_23018,N_17087,N_14603);
or U23019 (N_23019,N_14360,N_15690);
xnor U23020 (N_23020,N_12965,N_14572);
and U23021 (N_23021,N_13663,N_17143);
nor U23022 (N_23022,N_12824,N_16084);
or U23023 (N_23023,N_16608,N_14919);
or U23024 (N_23024,N_16527,N_17506);
nor U23025 (N_23025,N_17266,N_12515);
nand U23026 (N_23026,N_16271,N_17222);
and U23027 (N_23027,N_14894,N_12229);
nand U23028 (N_23028,N_16636,N_14662);
or U23029 (N_23029,N_12661,N_17015);
nor U23030 (N_23030,N_16109,N_13455);
and U23031 (N_23031,N_16138,N_12417);
or U23032 (N_23032,N_16880,N_13128);
and U23033 (N_23033,N_14342,N_14853);
xor U23034 (N_23034,N_12937,N_14320);
or U23035 (N_23035,N_15730,N_13292);
nand U23036 (N_23036,N_13552,N_16584);
xnor U23037 (N_23037,N_17778,N_14344);
or U23038 (N_23038,N_14599,N_12573);
or U23039 (N_23039,N_14144,N_13044);
nand U23040 (N_23040,N_16000,N_13846);
nand U23041 (N_23041,N_12530,N_17568);
nor U23042 (N_23042,N_12002,N_15299);
or U23043 (N_23043,N_12660,N_15434);
or U23044 (N_23044,N_17807,N_13227);
nor U23045 (N_23045,N_12771,N_17327);
or U23046 (N_23046,N_16531,N_14587);
xor U23047 (N_23047,N_15572,N_17918);
xnor U23048 (N_23048,N_14411,N_15585);
or U23049 (N_23049,N_14121,N_12890);
or U23050 (N_23050,N_15186,N_17306);
nand U23051 (N_23051,N_14472,N_12060);
and U23052 (N_23052,N_12985,N_12322);
or U23053 (N_23053,N_14593,N_15004);
and U23054 (N_23054,N_13781,N_17249);
nand U23055 (N_23055,N_17188,N_13077);
nor U23056 (N_23056,N_15164,N_14481);
xnor U23057 (N_23057,N_15520,N_16386);
or U23058 (N_23058,N_13310,N_17821);
or U23059 (N_23059,N_15350,N_13956);
nor U23060 (N_23060,N_13851,N_15263);
and U23061 (N_23061,N_12703,N_14444);
and U23062 (N_23062,N_13101,N_12889);
and U23063 (N_23063,N_14608,N_16048);
and U23064 (N_23064,N_17236,N_13265);
or U23065 (N_23065,N_17004,N_12255);
nand U23066 (N_23066,N_17114,N_13047);
xor U23067 (N_23067,N_15182,N_12722);
nor U23068 (N_23068,N_13461,N_13736);
or U23069 (N_23069,N_12225,N_17887);
nor U23070 (N_23070,N_16359,N_13329);
nor U23071 (N_23071,N_13480,N_12473);
and U23072 (N_23072,N_15777,N_14109);
or U23073 (N_23073,N_15782,N_16195);
or U23074 (N_23074,N_13025,N_14540);
xnor U23075 (N_23075,N_17610,N_16188);
or U23076 (N_23076,N_17450,N_13190);
or U23077 (N_23077,N_12843,N_12910);
or U23078 (N_23078,N_15296,N_12349);
nand U23079 (N_23079,N_14968,N_12512);
xor U23080 (N_23080,N_16776,N_16041);
nand U23081 (N_23081,N_13238,N_16532);
and U23082 (N_23082,N_17870,N_14129);
and U23083 (N_23083,N_17586,N_13475);
and U23084 (N_23084,N_15637,N_12362);
nor U23085 (N_23085,N_13215,N_13769);
nor U23086 (N_23086,N_17328,N_13451);
nor U23087 (N_23087,N_13340,N_16108);
nand U23088 (N_23088,N_14721,N_16161);
xnor U23089 (N_23089,N_16079,N_13554);
and U23090 (N_23090,N_16190,N_15716);
nand U23091 (N_23091,N_16428,N_14654);
xor U23092 (N_23092,N_13849,N_14643);
or U23093 (N_23093,N_12613,N_16072);
xnor U23094 (N_23094,N_12547,N_16218);
and U23095 (N_23095,N_16522,N_16949);
and U23096 (N_23096,N_16677,N_16481);
nor U23097 (N_23097,N_15313,N_15772);
nor U23098 (N_23098,N_16930,N_12029);
and U23099 (N_23099,N_15722,N_15153);
xnor U23100 (N_23100,N_14895,N_14010);
or U23101 (N_23101,N_16380,N_16000);
nand U23102 (N_23102,N_16473,N_15225);
or U23103 (N_23103,N_13014,N_13922);
and U23104 (N_23104,N_17767,N_14354);
xor U23105 (N_23105,N_12700,N_14438);
nand U23106 (N_23106,N_14584,N_13911);
xnor U23107 (N_23107,N_12273,N_14522);
and U23108 (N_23108,N_12979,N_17801);
nor U23109 (N_23109,N_14616,N_13989);
or U23110 (N_23110,N_15573,N_12690);
xor U23111 (N_23111,N_17748,N_17444);
or U23112 (N_23112,N_14785,N_14462);
and U23113 (N_23113,N_16178,N_13532);
and U23114 (N_23114,N_13633,N_15527);
nor U23115 (N_23115,N_14573,N_17826);
nor U23116 (N_23116,N_16541,N_15057);
nor U23117 (N_23117,N_12212,N_17500);
xnor U23118 (N_23118,N_15610,N_17323);
nand U23119 (N_23119,N_15583,N_16481);
and U23120 (N_23120,N_16017,N_16960);
nor U23121 (N_23121,N_12699,N_13718);
xor U23122 (N_23122,N_17935,N_14027);
or U23123 (N_23123,N_12956,N_17491);
or U23124 (N_23124,N_12220,N_16148);
and U23125 (N_23125,N_17519,N_14920);
xor U23126 (N_23126,N_14758,N_16803);
and U23127 (N_23127,N_15881,N_13694);
xnor U23128 (N_23128,N_17907,N_14459);
or U23129 (N_23129,N_17547,N_12771);
nand U23130 (N_23130,N_16344,N_12902);
nand U23131 (N_23131,N_12287,N_17328);
nor U23132 (N_23132,N_13692,N_15985);
or U23133 (N_23133,N_15554,N_17077);
or U23134 (N_23134,N_16827,N_17661);
and U23135 (N_23135,N_17431,N_12911);
and U23136 (N_23136,N_13628,N_14031);
xor U23137 (N_23137,N_14998,N_14571);
xnor U23138 (N_23138,N_14562,N_16879);
or U23139 (N_23139,N_16829,N_17572);
xnor U23140 (N_23140,N_15547,N_15618);
nand U23141 (N_23141,N_17246,N_17434);
nand U23142 (N_23142,N_12786,N_12742);
and U23143 (N_23143,N_13986,N_14873);
and U23144 (N_23144,N_17642,N_15420);
nor U23145 (N_23145,N_15328,N_17594);
nor U23146 (N_23146,N_16174,N_13230);
nor U23147 (N_23147,N_13137,N_16498);
nand U23148 (N_23148,N_14679,N_12766);
xor U23149 (N_23149,N_17249,N_14556);
and U23150 (N_23150,N_13067,N_14246);
nor U23151 (N_23151,N_16200,N_16524);
nand U23152 (N_23152,N_16590,N_14512);
nand U23153 (N_23153,N_13122,N_17130);
xor U23154 (N_23154,N_14733,N_13833);
nand U23155 (N_23155,N_13003,N_14520);
or U23156 (N_23156,N_13438,N_16365);
and U23157 (N_23157,N_16191,N_12523);
or U23158 (N_23158,N_12264,N_12982);
xnor U23159 (N_23159,N_14718,N_17330);
or U23160 (N_23160,N_14624,N_13118);
or U23161 (N_23161,N_17607,N_13246);
or U23162 (N_23162,N_13002,N_13600);
nor U23163 (N_23163,N_17526,N_15526);
nand U23164 (N_23164,N_16273,N_17079);
or U23165 (N_23165,N_15208,N_12269);
nand U23166 (N_23166,N_16278,N_12168);
or U23167 (N_23167,N_13806,N_12961);
nor U23168 (N_23168,N_12614,N_14748);
xor U23169 (N_23169,N_13075,N_17610);
xnor U23170 (N_23170,N_12940,N_13931);
nor U23171 (N_23171,N_15202,N_15108);
xor U23172 (N_23172,N_14786,N_17823);
xnor U23173 (N_23173,N_12310,N_13073);
or U23174 (N_23174,N_15253,N_15790);
or U23175 (N_23175,N_12376,N_12260);
and U23176 (N_23176,N_12199,N_12670);
or U23177 (N_23177,N_12886,N_17742);
xnor U23178 (N_23178,N_14012,N_12548);
nor U23179 (N_23179,N_13341,N_14032);
and U23180 (N_23180,N_15865,N_12752);
nand U23181 (N_23181,N_16910,N_12551);
and U23182 (N_23182,N_15968,N_15893);
or U23183 (N_23183,N_16188,N_14674);
xor U23184 (N_23184,N_13699,N_17597);
or U23185 (N_23185,N_15914,N_16335);
xnor U23186 (N_23186,N_15506,N_16533);
and U23187 (N_23187,N_16313,N_16927);
or U23188 (N_23188,N_12118,N_12665);
and U23189 (N_23189,N_12163,N_17017);
and U23190 (N_23190,N_13987,N_12933);
nand U23191 (N_23191,N_13827,N_16905);
xnor U23192 (N_23192,N_16422,N_13269);
and U23193 (N_23193,N_17811,N_15895);
and U23194 (N_23194,N_14301,N_17348);
nor U23195 (N_23195,N_16928,N_15696);
nor U23196 (N_23196,N_15258,N_15256);
or U23197 (N_23197,N_13206,N_15585);
xor U23198 (N_23198,N_14307,N_14229);
nor U23199 (N_23199,N_13160,N_17237);
nand U23200 (N_23200,N_17217,N_13216);
xnor U23201 (N_23201,N_16260,N_15249);
and U23202 (N_23202,N_15529,N_14362);
xor U23203 (N_23203,N_12943,N_15413);
or U23204 (N_23204,N_17901,N_14699);
xnor U23205 (N_23205,N_17381,N_12495);
and U23206 (N_23206,N_14289,N_13140);
or U23207 (N_23207,N_13246,N_17776);
and U23208 (N_23208,N_15827,N_12187);
nand U23209 (N_23209,N_17978,N_12199);
xnor U23210 (N_23210,N_14399,N_17597);
and U23211 (N_23211,N_13374,N_12608);
xnor U23212 (N_23212,N_12472,N_14021);
and U23213 (N_23213,N_13003,N_13351);
and U23214 (N_23214,N_14000,N_14722);
or U23215 (N_23215,N_13737,N_16713);
xor U23216 (N_23216,N_14974,N_17479);
and U23217 (N_23217,N_15875,N_17720);
nor U23218 (N_23218,N_14554,N_14077);
or U23219 (N_23219,N_14383,N_16320);
xor U23220 (N_23220,N_17684,N_17534);
xnor U23221 (N_23221,N_12512,N_14440);
and U23222 (N_23222,N_17672,N_16391);
nand U23223 (N_23223,N_16955,N_17730);
nand U23224 (N_23224,N_16658,N_17556);
nor U23225 (N_23225,N_16653,N_17422);
and U23226 (N_23226,N_13454,N_12373);
and U23227 (N_23227,N_15390,N_12124);
nor U23228 (N_23228,N_15694,N_14896);
nor U23229 (N_23229,N_17493,N_14147);
nor U23230 (N_23230,N_17176,N_15132);
or U23231 (N_23231,N_17851,N_16446);
nand U23232 (N_23232,N_14829,N_13367);
xor U23233 (N_23233,N_13206,N_13771);
nand U23234 (N_23234,N_16041,N_12834);
nand U23235 (N_23235,N_14950,N_17056);
or U23236 (N_23236,N_15763,N_14348);
nor U23237 (N_23237,N_13537,N_13325);
and U23238 (N_23238,N_14926,N_14903);
or U23239 (N_23239,N_12270,N_17546);
nand U23240 (N_23240,N_15932,N_12439);
nor U23241 (N_23241,N_17415,N_13817);
and U23242 (N_23242,N_16608,N_13834);
nor U23243 (N_23243,N_12971,N_15462);
nand U23244 (N_23244,N_17975,N_17791);
or U23245 (N_23245,N_14360,N_12235);
and U23246 (N_23246,N_13715,N_15726);
nor U23247 (N_23247,N_13925,N_12173);
nand U23248 (N_23248,N_14632,N_17216);
nand U23249 (N_23249,N_12249,N_12338);
and U23250 (N_23250,N_17249,N_16167);
nor U23251 (N_23251,N_12509,N_14911);
nand U23252 (N_23252,N_17646,N_16318);
nand U23253 (N_23253,N_12096,N_12673);
xor U23254 (N_23254,N_17150,N_15803);
nor U23255 (N_23255,N_15341,N_12628);
or U23256 (N_23256,N_15555,N_14143);
nand U23257 (N_23257,N_17030,N_17265);
and U23258 (N_23258,N_13969,N_12181);
nor U23259 (N_23259,N_17018,N_16854);
nor U23260 (N_23260,N_14368,N_12565);
nand U23261 (N_23261,N_13738,N_15217);
nand U23262 (N_23262,N_16419,N_13431);
or U23263 (N_23263,N_17172,N_17354);
and U23264 (N_23264,N_15081,N_16538);
xnor U23265 (N_23265,N_15514,N_17695);
nand U23266 (N_23266,N_16795,N_13168);
xor U23267 (N_23267,N_12975,N_17753);
nand U23268 (N_23268,N_15011,N_17648);
nand U23269 (N_23269,N_15297,N_17395);
nor U23270 (N_23270,N_17628,N_14121);
nand U23271 (N_23271,N_12587,N_15899);
or U23272 (N_23272,N_17207,N_15974);
nand U23273 (N_23273,N_17774,N_14715);
xnor U23274 (N_23274,N_12725,N_14909);
xor U23275 (N_23275,N_12667,N_16433);
nand U23276 (N_23276,N_16041,N_17884);
or U23277 (N_23277,N_14543,N_15979);
and U23278 (N_23278,N_15322,N_14126);
nor U23279 (N_23279,N_13051,N_14877);
xor U23280 (N_23280,N_17462,N_16742);
xor U23281 (N_23281,N_16727,N_14864);
or U23282 (N_23282,N_17779,N_12232);
nor U23283 (N_23283,N_14147,N_13165);
xor U23284 (N_23284,N_16656,N_12998);
or U23285 (N_23285,N_15693,N_15339);
and U23286 (N_23286,N_17970,N_13487);
or U23287 (N_23287,N_15893,N_13622);
xnor U23288 (N_23288,N_17999,N_12629);
and U23289 (N_23289,N_12359,N_12001);
xnor U23290 (N_23290,N_12327,N_14633);
or U23291 (N_23291,N_16204,N_16694);
xor U23292 (N_23292,N_14523,N_17794);
xnor U23293 (N_23293,N_15355,N_12716);
nand U23294 (N_23294,N_16088,N_14639);
nand U23295 (N_23295,N_16323,N_15880);
nand U23296 (N_23296,N_15688,N_16454);
xnor U23297 (N_23297,N_12926,N_15783);
or U23298 (N_23298,N_12026,N_12541);
and U23299 (N_23299,N_14230,N_14551);
and U23300 (N_23300,N_14781,N_13999);
and U23301 (N_23301,N_17956,N_12144);
nor U23302 (N_23302,N_17332,N_15826);
and U23303 (N_23303,N_16099,N_14605);
xnor U23304 (N_23304,N_12111,N_14257);
nand U23305 (N_23305,N_13380,N_12246);
nand U23306 (N_23306,N_16045,N_16378);
nand U23307 (N_23307,N_17768,N_15594);
and U23308 (N_23308,N_17251,N_14514);
or U23309 (N_23309,N_12041,N_17415);
xor U23310 (N_23310,N_14760,N_13935);
or U23311 (N_23311,N_17547,N_17128);
nand U23312 (N_23312,N_13116,N_12721);
or U23313 (N_23313,N_16709,N_12290);
nor U23314 (N_23314,N_15783,N_14312);
nand U23315 (N_23315,N_12256,N_15510);
nor U23316 (N_23316,N_12733,N_15561);
nand U23317 (N_23317,N_16405,N_17381);
xor U23318 (N_23318,N_17152,N_17510);
nor U23319 (N_23319,N_16561,N_13544);
or U23320 (N_23320,N_13275,N_14241);
xor U23321 (N_23321,N_17149,N_14365);
xnor U23322 (N_23322,N_14995,N_17598);
xnor U23323 (N_23323,N_12760,N_13327);
nor U23324 (N_23324,N_13084,N_16036);
nand U23325 (N_23325,N_13537,N_16199);
nand U23326 (N_23326,N_13654,N_13379);
nand U23327 (N_23327,N_12916,N_16347);
and U23328 (N_23328,N_13730,N_17523);
and U23329 (N_23329,N_15542,N_15296);
nand U23330 (N_23330,N_14675,N_16003);
xor U23331 (N_23331,N_13709,N_17726);
or U23332 (N_23332,N_16853,N_13132);
and U23333 (N_23333,N_16875,N_13982);
nand U23334 (N_23334,N_12672,N_15976);
and U23335 (N_23335,N_16349,N_12957);
and U23336 (N_23336,N_17240,N_15578);
xnor U23337 (N_23337,N_17462,N_12821);
nand U23338 (N_23338,N_14672,N_14714);
and U23339 (N_23339,N_15035,N_15186);
or U23340 (N_23340,N_15823,N_12278);
nor U23341 (N_23341,N_13318,N_12126);
nand U23342 (N_23342,N_16239,N_17412);
xnor U23343 (N_23343,N_17139,N_17715);
nand U23344 (N_23344,N_16199,N_15003);
nor U23345 (N_23345,N_16903,N_15499);
and U23346 (N_23346,N_17209,N_13631);
nand U23347 (N_23347,N_17558,N_16523);
or U23348 (N_23348,N_12618,N_15636);
or U23349 (N_23349,N_12368,N_15301);
nand U23350 (N_23350,N_16028,N_12863);
and U23351 (N_23351,N_12839,N_13566);
nand U23352 (N_23352,N_16641,N_12757);
nor U23353 (N_23353,N_14402,N_14748);
nor U23354 (N_23354,N_12327,N_17370);
or U23355 (N_23355,N_16817,N_13483);
and U23356 (N_23356,N_12640,N_15263);
or U23357 (N_23357,N_12610,N_13115);
nand U23358 (N_23358,N_12227,N_16069);
nand U23359 (N_23359,N_17087,N_15910);
and U23360 (N_23360,N_14892,N_16672);
or U23361 (N_23361,N_17886,N_12415);
nor U23362 (N_23362,N_14332,N_14814);
nand U23363 (N_23363,N_16749,N_12499);
xor U23364 (N_23364,N_14982,N_14766);
xnor U23365 (N_23365,N_14049,N_16841);
nand U23366 (N_23366,N_17563,N_16250);
or U23367 (N_23367,N_14653,N_12998);
nor U23368 (N_23368,N_14444,N_14429);
nor U23369 (N_23369,N_12995,N_16827);
nand U23370 (N_23370,N_15999,N_12695);
nor U23371 (N_23371,N_15219,N_12026);
nor U23372 (N_23372,N_14695,N_15804);
and U23373 (N_23373,N_15615,N_15471);
nor U23374 (N_23374,N_13677,N_17014);
or U23375 (N_23375,N_17743,N_16311);
or U23376 (N_23376,N_16398,N_12368);
nand U23377 (N_23377,N_13002,N_16139);
or U23378 (N_23378,N_12512,N_17436);
and U23379 (N_23379,N_16783,N_12084);
nand U23380 (N_23380,N_17732,N_12389);
or U23381 (N_23381,N_15593,N_12269);
xnor U23382 (N_23382,N_17610,N_15055);
and U23383 (N_23383,N_16436,N_15323);
nor U23384 (N_23384,N_15130,N_16590);
or U23385 (N_23385,N_12397,N_16084);
and U23386 (N_23386,N_13494,N_13939);
or U23387 (N_23387,N_16690,N_16687);
or U23388 (N_23388,N_15663,N_15580);
nor U23389 (N_23389,N_12499,N_16675);
or U23390 (N_23390,N_12519,N_17365);
nand U23391 (N_23391,N_16444,N_12583);
and U23392 (N_23392,N_13374,N_12308);
and U23393 (N_23393,N_13726,N_13676);
xnor U23394 (N_23394,N_14021,N_17957);
or U23395 (N_23395,N_15590,N_16416);
nor U23396 (N_23396,N_13821,N_17609);
and U23397 (N_23397,N_16897,N_12183);
nand U23398 (N_23398,N_17171,N_13517);
xnor U23399 (N_23399,N_15566,N_17512);
nand U23400 (N_23400,N_15372,N_15219);
nand U23401 (N_23401,N_12314,N_13165);
xor U23402 (N_23402,N_17739,N_15799);
nand U23403 (N_23403,N_15065,N_14963);
nand U23404 (N_23404,N_13910,N_15321);
or U23405 (N_23405,N_16783,N_12101);
and U23406 (N_23406,N_15201,N_13477);
and U23407 (N_23407,N_15868,N_16204);
or U23408 (N_23408,N_17053,N_17279);
or U23409 (N_23409,N_12599,N_12319);
and U23410 (N_23410,N_14672,N_13166);
or U23411 (N_23411,N_14179,N_16873);
and U23412 (N_23412,N_13311,N_12336);
or U23413 (N_23413,N_15097,N_17605);
and U23414 (N_23414,N_15283,N_12165);
xor U23415 (N_23415,N_16192,N_13749);
or U23416 (N_23416,N_17960,N_12860);
nor U23417 (N_23417,N_13477,N_16847);
nor U23418 (N_23418,N_14869,N_17750);
nand U23419 (N_23419,N_13281,N_16154);
nor U23420 (N_23420,N_13767,N_15732);
and U23421 (N_23421,N_16603,N_13228);
xnor U23422 (N_23422,N_12326,N_16067);
nand U23423 (N_23423,N_15080,N_15609);
nor U23424 (N_23424,N_13910,N_14258);
nand U23425 (N_23425,N_16303,N_15971);
and U23426 (N_23426,N_13599,N_17716);
nor U23427 (N_23427,N_12926,N_16296);
or U23428 (N_23428,N_16343,N_14939);
or U23429 (N_23429,N_12066,N_15754);
or U23430 (N_23430,N_13347,N_12434);
or U23431 (N_23431,N_16826,N_13645);
nor U23432 (N_23432,N_13202,N_14902);
and U23433 (N_23433,N_14934,N_15607);
xnor U23434 (N_23434,N_12645,N_13433);
and U23435 (N_23435,N_17447,N_13557);
nor U23436 (N_23436,N_16036,N_12298);
xnor U23437 (N_23437,N_15602,N_13899);
or U23438 (N_23438,N_13066,N_17254);
or U23439 (N_23439,N_13140,N_14370);
nor U23440 (N_23440,N_14344,N_15012);
nor U23441 (N_23441,N_17258,N_14726);
nor U23442 (N_23442,N_15445,N_14149);
and U23443 (N_23443,N_14365,N_17626);
and U23444 (N_23444,N_14831,N_15592);
or U23445 (N_23445,N_13265,N_17620);
xnor U23446 (N_23446,N_14577,N_17895);
xor U23447 (N_23447,N_16659,N_12793);
nand U23448 (N_23448,N_14377,N_17278);
and U23449 (N_23449,N_14762,N_15372);
nand U23450 (N_23450,N_16168,N_17690);
xor U23451 (N_23451,N_15102,N_13922);
nand U23452 (N_23452,N_14614,N_17407);
nor U23453 (N_23453,N_15253,N_15659);
nor U23454 (N_23454,N_15336,N_14354);
nor U23455 (N_23455,N_13096,N_15736);
or U23456 (N_23456,N_15132,N_14500);
xnor U23457 (N_23457,N_17441,N_14849);
nand U23458 (N_23458,N_15892,N_17205);
nor U23459 (N_23459,N_12227,N_14234);
xnor U23460 (N_23460,N_17834,N_17427);
or U23461 (N_23461,N_13084,N_13899);
or U23462 (N_23462,N_16510,N_12013);
xnor U23463 (N_23463,N_12646,N_17589);
nor U23464 (N_23464,N_12185,N_13663);
xor U23465 (N_23465,N_16534,N_14673);
nor U23466 (N_23466,N_15517,N_13711);
and U23467 (N_23467,N_15205,N_16968);
and U23468 (N_23468,N_14162,N_13567);
or U23469 (N_23469,N_16858,N_15864);
xnor U23470 (N_23470,N_14745,N_14670);
xnor U23471 (N_23471,N_15977,N_13473);
or U23472 (N_23472,N_13945,N_15783);
nor U23473 (N_23473,N_14211,N_16403);
and U23474 (N_23474,N_14314,N_16664);
nand U23475 (N_23475,N_14005,N_16445);
nand U23476 (N_23476,N_16256,N_14616);
nand U23477 (N_23477,N_15688,N_16222);
or U23478 (N_23478,N_14059,N_12576);
xnor U23479 (N_23479,N_15822,N_14146);
nor U23480 (N_23480,N_13816,N_12044);
nor U23481 (N_23481,N_17794,N_15049);
nor U23482 (N_23482,N_12585,N_16640);
or U23483 (N_23483,N_14597,N_12862);
xnor U23484 (N_23484,N_16476,N_17204);
and U23485 (N_23485,N_14511,N_17855);
or U23486 (N_23486,N_14663,N_15674);
nand U23487 (N_23487,N_16828,N_13229);
and U23488 (N_23488,N_17252,N_13005);
and U23489 (N_23489,N_15518,N_13639);
xnor U23490 (N_23490,N_13211,N_14911);
nor U23491 (N_23491,N_14221,N_14609);
nor U23492 (N_23492,N_16154,N_15637);
and U23493 (N_23493,N_16430,N_14382);
and U23494 (N_23494,N_14675,N_13784);
nand U23495 (N_23495,N_14443,N_12399);
nand U23496 (N_23496,N_14842,N_16428);
nand U23497 (N_23497,N_13466,N_13046);
nand U23498 (N_23498,N_12130,N_14234);
nor U23499 (N_23499,N_12240,N_14074);
or U23500 (N_23500,N_14536,N_13175);
or U23501 (N_23501,N_16592,N_17210);
and U23502 (N_23502,N_14817,N_13401);
or U23503 (N_23503,N_12540,N_15474);
xnor U23504 (N_23504,N_17682,N_15041);
xnor U23505 (N_23505,N_13756,N_15344);
nand U23506 (N_23506,N_15399,N_14522);
nor U23507 (N_23507,N_15416,N_16868);
nor U23508 (N_23508,N_12814,N_13848);
and U23509 (N_23509,N_15081,N_12019);
xnor U23510 (N_23510,N_15687,N_15811);
or U23511 (N_23511,N_14930,N_17153);
nand U23512 (N_23512,N_13490,N_13472);
xnor U23513 (N_23513,N_17173,N_17995);
nor U23514 (N_23514,N_13560,N_16670);
nor U23515 (N_23515,N_12217,N_14750);
nor U23516 (N_23516,N_12090,N_14449);
xor U23517 (N_23517,N_16583,N_14458);
or U23518 (N_23518,N_14316,N_14720);
nor U23519 (N_23519,N_15519,N_16185);
xnor U23520 (N_23520,N_13877,N_16794);
nor U23521 (N_23521,N_15632,N_13655);
nand U23522 (N_23522,N_12406,N_13708);
nor U23523 (N_23523,N_16243,N_16521);
and U23524 (N_23524,N_12847,N_14864);
and U23525 (N_23525,N_12232,N_14441);
nor U23526 (N_23526,N_17278,N_15676);
xnor U23527 (N_23527,N_14897,N_17248);
and U23528 (N_23528,N_14307,N_13477);
or U23529 (N_23529,N_12746,N_16036);
and U23530 (N_23530,N_16810,N_13981);
nand U23531 (N_23531,N_15741,N_17724);
and U23532 (N_23532,N_12082,N_17920);
and U23533 (N_23533,N_16668,N_12120);
nor U23534 (N_23534,N_13800,N_13961);
xnor U23535 (N_23535,N_17799,N_12525);
or U23536 (N_23536,N_12951,N_16582);
nor U23537 (N_23537,N_14085,N_16945);
and U23538 (N_23538,N_17080,N_12304);
xor U23539 (N_23539,N_13121,N_14552);
or U23540 (N_23540,N_12377,N_13072);
or U23541 (N_23541,N_13867,N_15393);
xnor U23542 (N_23542,N_13130,N_14279);
nor U23543 (N_23543,N_17417,N_16048);
xnor U23544 (N_23544,N_14644,N_12128);
or U23545 (N_23545,N_16348,N_15113);
nor U23546 (N_23546,N_13397,N_15477);
or U23547 (N_23547,N_16465,N_16202);
nand U23548 (N_23548,N_13112,N_16302);
nand U23549 (N_23549,N_17914,N_12979);
and U23550 (N_23550,N_17348,N_15219);
nor U23551 (N_23551,N_15166,N_16528);
nand U23552 (N_23552,N_13565,N_12235);
or U23553 (N_23553,N_17728,N_13157);
and U23554 (N_23554,N_13257,N_17522);
or U23555 (N_23555,N_15703,N_14422);
xor U23556 (N_23556,N_12093,N_16371);
and U23557 (N_23557,N_17217,N_16788);
or U23558 (N_23558,N_16383,N_17803);
nor U23559 (N_23559,N_17864,N_14706);
or U23560 (N_23560,N_16861,N_16148);
nor U23561 (N_23561,N_16257,N_16987);
and U23562 (N_23562,N_13498,N_13767);
nand U23563 (N_23563,N_15696,N_12588);
xnor U23564 (N_23564,N_12090,N_15224);
and U23565 (N_23565,N_13642,N_15499);
nand U23566 (N_23566,N_12330,N_14990);
and U23567 (N_23567,N_13445,N_13520);
and U23568 (N_23568,N_12904,N_13258);
xnor U23569 (N_23569,N_12305,N_12773);
nor U23570 (N_23570,N_14055,N_12017);
nor U23571 (N_23571,N_17597,N_12371);
nor U23572 (N_23572,N_17057,N_13989);
xnor U23573 (N_23573,N_15838,N_12688);
nor U23574 (N_23574,N_13760,N_13906);
xnor U23575 (N_23575,N_15275,N_14755);
nor U23576 (N_23576,N_15842,N_13095);
nand U23577 (N_23577,N_16877,N_17164);
xor U23578 (N_23578,N_16092,N_16003);
nor U23579 (N_23579,N_15959,N_15639);
nand U23580 (N_23580,N_13298,N_14889);
and U23581 (N_23581,N_17775,N_14256);
xor U23582 (N_23582,N_13018,N_15575);
nand U23583 (N_23583,N_17092,N_13042);
or U23584 (N_23584,N_15815,N_13977);
or U23585 (N_23585,N_17978,N_14450);
xor U23586 (N_23586,N_12920,N_15068);
and U23587 (N_23587,N_15952,N_13927);
nand U23588 (N_23588,N_15961,N_16131);
or U23589 (N_23589,N_15646,N_17763);
nand U23590 (N_23590,N_16876,N_13594);
or U23591 (N_23591,N_15665,N_12081);
nand U23592 (N_23592,N_12097,N_15761);
and U23593 (N_23593,N_14482,N_14066);
nand U23594 (N_23594,N_12096,N_12668);
or U23595 (N_23595,N_17252,N_15750);
and U23596 (N_23596,N_16731,N_14601);
nor U23597 (N_23597,N_15765,N_13408);
and U23598 (N_23598,N_17697,N_15106);
or U23599 (N_23599,N_13161,N_17467);
or U23600 (N_23600,N_14771,N_17569);
xnor U23601 (N_23601,N_17805,N_16258);
nand U23602 (N_23602,N_13461,N_17227);
xnor U23603 (N_23603,N_14026,N_17203);
or U23604 (N_23604,N_14278,N_12427);
nand U23605 (N_23605,N_15144,N_15694);
nor U23606 (N_23606,N_13549,N_15112);
xnor U23607 (N_23607,N_16977,N_14090);
xnor U23608 (N_23608,N_15065,N_14261);
nand U23609 (N_23609,N_17384,N_16492);
and U23610 (N_23610,N_14692,N_15878);
and U23611 (N_23611,N_15265,N_13138);
and U23612 (N_23612,N_12009,N_13314);
nand U23613 (N_23613,N_17886,N_16333);
xor U23614 (N_23614,N_16359,N_15121);
nor U23615 (N_23615,N_12902,N_14300);
and U23616 (N_23616,N_17753,N_16910);
nor U23617 (N_23617,N_16912,N_12824);
or U23618 (N_23618,N_13135,N_15473);
xor U23619 (N_23619,N_14170,N_15272);
and U23620 (N_23620,N_16381,N_13565);
and U23621 (N_23621,N_17925,N_15528);
nor U23622 (N_23622,N_12666,N_14796);
nand U23623 (N_23623,N_14567,N_14154);
or U23624 (N_23624,N_13803,N_17110);
nor U23625 (N_23625,N_17018,N_17264);
nand U23626 (N_23626,N_15706,N_13192);
or U23627 (N_23627,N_15676,N_12916);
or U23628 (N_23628,N_13713,N_14233);
and U23629 (N_23629,N_15932,N_16399);
and U23630 (N_23630,N_14976,N_16800);
nor U23631 (N_23631,N_16235,N_17359);
nand U23632 (N_23632,N_14438,N_14256);
nor U23633 (N_23633,N_17631,N_13650);
nor U23634 (N_23634,N_14643,N_12022);
nor U23635 (N_23635,N_12692,N_12754);
and U23636 (N_23636,N_16828,N_14800);
nor U23637 (N_23637,N_15060,N_14853);
nand U23638 (N_23638,N_13105,N_15483);
xor U23639 (N_23639,N_17335,N_15555);
nor U23640 (N_23640,N_13843,N_16273);
and U23641 (N_23641,N_17473,N_13775);
nor U23642 (N_23642,N_12047,N_13131);
nor U23643 (N_23643,N_15532,N_14784);
nand U23644 (N_23644,N_14299,N_12826);
xor U23645 (N_23645,N_14060,N_12903);
xnor U23646 (N_23646,N_14900,N_17673);
or U23647 (N_23647,N_15609,N_14177);
or U23648 (N_23648,N_15996,N_15847);
nand U23649 (N_23649,N_14376,N_15337);
or U23650 (N_23650,N_15335,N_16446);
xnor U23651 (N_23651,N_15517,N_14060);
and U23652 (N_23652,N_13710,N_12546);
and U23653 (N_23653,N_12426,N_16623);
and U23654 (N_23654,N_14629,N_14541);
xnor U23655 (N_23655,N_15447,N_16679);
or U23656 (N_23656,N_13931,N_15588);
or U23657 (N_23657,N_16474,N_15884);
nand U23658 (N_23658,N_12287,N_14246);
and U23659 (N_23659,N_17130,N_12200);
or U23660 (N_23660,N_17576,N_14121);
nor U23661 (N_23661,N_12209,N_14944);
nand U23662 (N_23662,N_14214,N_16180);
and U23663 (N_23663,N_12403,N_14904);
or U23664 (N_23664,N_15511,N_15570);
or U23665 (N_23665,N_17289,N_14164);
and U23666 (N_23666,N_14999,N_12582);
xnor U23667 (N_23667,N_16051,N_15832);
and U23668 (N_23668,N_12599,N_12906);
and U23669 (N_23669,N_13878,N_14086);
and U23670 (N_23670,N_15173,N_15548);
or U23671 (N_23671,N_15509,N_12141);
nand U23672 (N_23672,N_15205,N_13545);
or U23673 (N_23673,N_16811,N_17870);
or U23674 (N_23674,N_13889,N_17169);
or U23675 (N_23675,N_15727,N_17407);
nand U23676 (N_23676,N_12821,N_17477);
or U23677 (N_23677,N_12947,N_14170);
xor U23678 (N_23678,N_14244,N_17325);
or U23679 (N_23679,N_17984,N_14933);
nand U23680 (N_23680,N_15247,N_13022);
nand U23681 (N_23681,N_14216,N_17820);
nand U23682 (N_23682,N_14381,N_17869);
or U23683 (N_23683,N_12626,N_15966);
nand U23684 (N_23684,N_12006,N_15292);
and U23685 (N_23685,N_16030,N_14687);
and U23686 (N_23686,N_17648,N_14427);
nand U23687 (N_23687,N_12347,N_16400);
or U23688 (N_23688,N_16309,N_15678);
nand U23689 (N_23689,N_13565,N_12848);
and U23690 (N_23690,N_14822,N_13308);
nand U23691 (N_23691,N_15082,N_14244);
and U23692 (N_23692,N_15027,N_17527);
nand U23693 (N_23693,N_16136,N_14258);
and U23694 (N_23694,N_15235,N_16688);
nor U23695 (N_23695,N_13856,N_17609);
or U23696 (N_23696,N_15445,N_13625);
and U23697 (N_23697,N_12606,N_17179);
or U23698 (N_23698,N_15041,N_13146);
and U23699 (N_23699,N_13422,N_14039);
nand U23700 (N_23700,N_14114,N_13378);
nor U23701 (N_23701,N_16028,N_14346);
nor U23702 (N_23702,N_16123,N_14132);
and U23703 (N_23703,N_13352,N_16600);
nand U23704 (N_23704,N_17527,N_16628);
nand U23705 (N_23705,N_15113,N_16672);
and U23706 (N_23706,N_16902,N_17650);
or U23707 (N_23707,N_17664,N_16131);
xnor U23708 (N_23708,N_14728,N_16590);
nor U23709 (N_23709,N_15670,N_15037);
nand U23710 (N_23710,N_16557,N_13036);
xor U23711 (N_23711,N_14894,N_13982);
nand U23712 (N_23712,N_14768,N_12045);
nor U23713 (N_23713,N_13385,N_17621);
xnor U23714 (N_23714,N_15292,N_16903);
nor U23715 (N_23715,N_12716,N_16385);
xor U23716 (N_23716,N_14219,N_15736);
nand U23717 (N_23717,N_15459,N_16743);
or U23718 (N_23718,N_15103,N_14611);
or U23719 (N_23719,N_14234,N_14026);
and U23720 (N_23720,N_14712,N_15813);
xor U23721 (N_23721,N_17512,N_15351);
and U23722 (N_23722,N_16624,N_16497);
or U23723 (N_23723,N_12854,N_16268);
nor U23724 (N_23724,N_17251,N_15118);
nand U23725 (N_23725,N_17045,N_12318);
xnor U23726 (N_23726,N_14021,N_12735);
or U23727 (N_23727,N_16000,N_12141);
nor U23728 (N_23728,N_13939,N_13794);
xor U23729 (N_23729,N_14463,N_14565);
xnor U23730 (N_23730,N_13669,N_15041);
nand U23731 (N_23731,N_13211,N_12773);
nor U23732 (N_23732,N_12367,N_16620);
nand U23733 (N_23733,N_14409,N_12935);
xor U23734 (N_23734,N_15270,N_16979);
xnor U23735 (N_23735,N_16623,N_13104);
nand U23736 (N_23736,N_17520,N_12510);
or U23737 (N_23737,N_13344,N_17521);
nor U23738 (N_23738,N_14955,N_12106);
nand U23739 (N_23739,N_12271,N_13085);
or U23740 (N_23740,N_17750,N_15166);
or U23741 (N_23741,N_14598,N_16965);
or U23742 (N_23742,N_14651,N_12722);
nand U23743 (N_23743,N_14658,N_12394);
nand U23744 (N_23744,N_14352,N_13463);
and U23745 (N_23745,N_16248,N_14384);
and U23746 (N_23746,N_14837,N_12473);
xor U23747 (N_23747,N_17257,N_16002);
nor U23748 (N_23748,N_13494,N_17567);
and U23749 (N_23749,N_16033,N_13447);
nand U23750 (N_23750,N_16243,N_14018);
or U23751 (N_23751,N_12202,N_17914);
nand U23752 (N_23752,N_14631,N_12232);
xnor U23753 (N_23753,N_13623,N_16066);
nand U23754 (N_23754,N_13619,N_16466);
or U23755 (N_23755,N_14546,N_12808);
nand U23756 (N_23756,N_17762,N_13782);
nor U23757 (N_23757,N_15756,N_12204);
or U23758 (N_23758,N_13705,N_13753);
xor U23759 (N_23759,N_12553,N_12635);
nand U23760 (N_23760,N_13676,N_15323);
nand U23761 (N_23761,N_14576,N_16386);
and U23762 (N_23762,N_14630,N_15820);
nand U23763 (N_23763,N_15704,N_12094);
nor U23764 (N_23764,N_13282,N_16577);
xnor U23765 (N_23765,N_17001,N_13411);
nand U23766 (N_23766,N_13789,N_17798);
and U23767 (N_23767,N_16512,N_16504);
xnor U23768 (N_23768,N_12225,N_17108);
and U23769 (N_23769,N_17327,N_13129);
xor U23770 (N_23770,N_17713,N_12017);
xor U23771 (N_23771,N_12512,N_15771);
xor U23772 (N_23772,N_13994,N_16786);
and U23773 (N_23773,N_14226,N_13980);
or U23774 (N_23774,N_16775,N_15416);
xnor U23775 (N_23775,N_14412,N_13470);
nor U23776 (N_23776,N_14360,N_14419);
nand U23777 (N_23777,N_17595,N_12940);
xnor U23778 (N_23778,N_12602,N_16847);
or U23779 (N_23779,N_16089,N_17852);
and U23780 (N_23780,N_17126,N_13914);
and U23781 (N_23781,N_12694,N_14449);
and U23782 (N_23782,N_16124,N_14465);
and U23783 (N_23783,N_12929,N_13326);
xnor U23784 (N_23784,N_15051,N_13330);
nor U23785 (N_23785,N_12526,N_16825);
xor U23786 (N_23786,N_12999,N_14726);
nand U23787 (N_23787,N_13390,N_12806);
nand U23788 (N_23788,N_12270,N_12991);
xor U23789 (N_23789,N_14149,N_15333);
and U23790 (N_23790,N_15159,N_12787);
and U23791 (N_23791,N_12114,N_15284);
nor U23792 (N_23792,N_14779,N_15146);
and U23793 (N_23793,N_15603,N_14513);
nor U23794 (N_23794,N_13943,N_14632);
nand U23795 (N_23795,N_17636,N_17772);
or U23796 (N_23796,N_15293,N_15153);
or U23797 (N_23797,N_12066,N_15675);
nand U23798 (N_23798,N_13292,N_15676);
and U23799 (N_23799,N_13423,N_17781);
xor U23800 (N_23800,N_12640,N_13053);
xnor U23801 (N_23801,N_13866,N_17477);
nand U23802 (N_23802,N_12122,N_15020);
nand U23803 (N_23803,N_15879,N_16609);
xor U23804 (N_23804,N_13122,N_12476);
or U23805 (N_23805,N_12135,N_17809);
and U23806 (N_23806,N_16385,N_14737);
and U23807 (N_23807,N_16702,N_16514);
and U23808 (N_23808,N_16765,N_12445);
and U23809 (N_23809,N_17441,N_14041);
xor U23810 (N_23810,N_14537,N_14165);
or U23811 (N_23811,N_16073,N_16476);
and U23812 (N_23812,N_16927,N_15318);
and U23813 (N_23813,N_17878,N_13906);
xnor U23814 (N_23814,N_14562,N_13150);
nor U23815 (N_23815,N_12095,N_13908);
or U23816 (N_23816,N_16630,N_12318);
xor U23817 (N_23817,N_16134,N_13251);
or U23818 (N_23818,N_12067,N_14254);
or U23819 (N_23819,N_14039,N_13294);
xnor U23820 (N_23820,N_14481,N_17628);
nor U23821 (N_23821,N_15667,N_16879);
or U23822 (N_23822,N_14460,N_17390);
xnor U23823 (N_23823,N_16755,N_13621);
and U23824 (N_23824,N_16491,N_12633);
or U23825 (N_23825,N_14143,N_15006);
or U23826 (N_23826,N_15176,N_15033);
xor U23827 (N_23827,N_17828,N_15463);
and U23828 (N_23828,N_13295,N_17698);
and U23829 (N_23829,N_13926,N_16400);
and U23830 (N_23830,N_14483,N_12037);
nor U23831 (N_23831,N_17480,N_14595);
nor U23832 (N_23832,N_16099,N_15853);
xor U23833 (N_23833,N_14709,N_17086);
xnor U23834 (N_23834,N_15406,N_15307);
and U23835 (N_23835,N_13311,N_14140);
xor U23836 (N_23836,N_13989,N_17247);
nand U23837 (N_23837,N_12776,N_12813);
or U23838 (N_23838,N_15530,N_12357);
xnor U23839 (N_23839,N_15844,N_14525);
xor U23840 (N_23840,N_12249,N_13019);
xor U23841 (N_23841,N_12098,N_15540);
and U23842 (N_23842,N_17199,N_12085);
nand U23843 (N_23843,N_16278,N_14821);
or U23844 (N_23844,N_16770,N_14485);
nand U23845 (N_23845,N_16152,N_13141);
nand U23846 (N_23846,N_12971,N_12609);
nor U23847 (N_23847,N_14102,N_15792);
and U23848 (N_23848,N_13392,N_12841);
nand U23849 (N_23849,N_15499,N_16403);
or U23850 (N_23850,N_14414,N_14129);
or U23851 (N_23851,N_13306,N_13736);
xor U23852 (N_23852,N_12052,N_13765);
or U23853 (N_23853,N_13449,N_15932);
nor U23854 (N_23854,N_16596,N_12089);
or U23855 (N_23855,N_17355,N_15403);
xnor U23856 (N_23856,N_16937,N_12861);
and U23857 (N_23857,N_12802,N_15573);
nand U23858 (N_23858,N_12513,N_14499);
and U23859 (N_23859,N_14660,N_12551);
xor U23860 (N_23860,N_13713,N_16520);
and U23861 (N_23861,N_17858,N_17359);
or U23862 (N_23862,N_14523,N_14309);
nand U23863 (N_23863,N_14365,N_15399);
nor U23864 (N_23864,N_16411,N_16946);
nor U23865 (N_23865,N_14889,N_17604);
or U23866 (N_23866,N_16719,N_13751);
nor U23867 (N_23867,N_17743,N_16522);
xor U23868 (N_23868,N_12432,N_14159);
xor U23869 (N_23869,N_14513,N_14437);
nor U23870 (N_23870,N_14936,N_14819);
nor U23871 (N_23871,N_16772,N_17275);
xor U23872 (N_23872,N_13186,N_16721);
nand U23873 (N_23873,N_16027,N_14023);
xnor U23874 (N_23874,N_12926,N_16328);
nor U23875 (N_23875,N_13551,N_14329);
nor U23876 (N_23876,N_17318,N_17151);
nand U23877 (N_23877,N_12247,N_12650);
nor U23878 (N_23878,N_14594,N_17232);
or U23879 (N_23879,N_17976,N_15119);
nand U23880 (N_23880,N_16651,N_15643);
or U23881 (N_23881,N_14768,N_14839);
nand U23882 (N_23882,N_16466,N_16506);
or U23883 (N_23883,N_12881,N_14234);
xor U23884 (N_23884,N_13145,N_13163);
nor U23885 (N_23885,N_12774,N_14895);
nand U23886 (N_23886,N_12006,N_14083);
xnor U23887 (N_23887,N_17663,N_13347);
and U23888 (N_23888,N_16973,N_17245);
and U23889 (N_23889,N_12773,N_15015);
and U23890 (N_23890,N_14740,N_15770);
or U23891 (N_23891,N_15281,N_12967);
nand U23892 (N_23892,N_14269,N_15901);
nand U23893 (N_23893,N_16058,N_17815);
xor U23894 (N_23894,N_12572,N_13150);
and U23895 (N_23895,N_17088,N_12057);
xor U23896 (N_23896,N_13877,N_17895);
xnor U23897 (N_23897,N_17997,N_14710);
nand U23898 (N_23898,N_12786,N_16234);
or U23899 (N_23899,N_13358,N_15114);
or U23900 (N_23900,N_15870,N_15146);
or U23901 (N_23901,N_14659,N_12550);
nor U23902 (N_23902,N_13959,N_13553);
nand U23903 (N_23903,N_17766,N_12664);
nor U23904 (N_23904,N_17208,N_15121);
and U23905 (N_23905,N_12694,N_12603);
or U23906 (N_23906,N_15193,N_14099);
xor U23907 (N_23907,N_13612,N_16406);
xnor U23908 (N_23908,N_14696,N_14838);
nand U23909 (N_23909,N_13126,N_15135);
nor U23910 (N_23910,N_13233,N_17632);
nor U23911 (N_23911,N_16592,N_16800);
xnor U23912 (N_23912,N_16950,N_12483);
nor U23913 (N_23913,N_15777,N_17506);
and U23914 (N_23914,N_14554,N_17077);
and U23915 (N_23915,N_15543,N_14257);
xor U23916 (N_23916,N_14745,N_13652);
nor U23917 (N_23917,N_13327,N_15261);
and U23918 (N_23918,N_12219,N_14452);
and U23919 (N_23919,N_14599,N_17817);
nor U23920 (N_23920,N_14803,N_15756);
nor U23921 (N_23921,N_14915,N_15520);
and U23922 (N_23922,N_17118,N_13561);
nor U23923 (N_23923,N_17350,N_14348);
nor U23924 (N_23924,N_12669,N_16620);
xor U23925 (N_23925,N_12073,N_16589);
nor U23926 (N_23926,N_12711,N_16959);
xnor U23927 (N_23927,N_16943,N_13749);
nand U23928 (N_23928,N_12562,N_13331);
or U23929 (N_23929,N_14354,N_13499);
nand U23930 (N_23930,N_14048,N_14516);
or U23931 (N_23931,N_12124,N_15435);
xor U23932 (N_23932,N_15892,N_14508);
and U23933 (N_23933,N_15319,N_12479);
or U23934 (N_23934,N_16162,N_13132);
and U23935 (N_23935,N_12190,N_14046);
or U23936 (N_23936,N_13634,N_13421);
xnor U23937 (N_23937,N_12990,N_13366);
nand U23938 (N_23938,N_13504,N_16771);
or U23939 (N_23939,N_14771,N_12753);
and U23940 (N_23940,N_12786,N_15114);
xor U23941 (N_23941,N_13749,N_14912);
xnor U23942 (N_23942,N_16911,N_15330);
nor U23943 (N_23943,N_17671,N_12851);
xnor U23944 (N_23944,N_12099,N_12148);
xnor U23945 (N_23945,N_15495,N_13586);
xor U23946 (N_23946,N_13069,N_16572);
and U23947 (N_23947,N_13532,N_17241);
xnor U23948 (N_23948,N_17454,N_17948);
and U23949 (N_23949,N_17505,N_13188);
or U23950 (N_23950,N_17641,N_14703);
and U23951 (N_23951,N_14548,N_15469);
xor U23952 (N_23952,N_12274,N_13047);
nand U23953 (N_23953,N_12578,N_12922);
or U23954 (N_23954,N_15271,N_14554);
and U23955 (N_23955,N_14727,N_14520);
or U23956 (N_23956,N_15455,N_16498);
xnor U23957 (N_23957,N_14666,N_17090);
nand U23958 (N_23958,N_15067,N_15994);
or U23959 (N_23959,N_12987,N_16268);
and U23960 (N_23960,N_17327,N_13309);
nor U23961 (N_23961,N_16928,N_14709);
and U23962 (N_23962,N_12468,N_17752);
nand U23963 (N_23963,N_16622,N_15935);
or U23964 (N_23964,N_16557,N_15270);
and U23965 (N_23965,N_13586,N_17934);
nor U23966 (N_23966,N_16557,N_14873);
or U23967 (N_23967,N_15173,N_15879);
xor U23968 (N_23968,N_13442,N_13770);
xor U23969 (N_23969,N_15121,N_12635);
nor U23970 (N_23970,N_12089,N_15352);
nand U23971 (N_23971,N_17970,N_15933);
nor U23972 (N_23972,N_17156,N_16795);
xnor U23973 (N_23973,N_13165,N_17243);
or U23974 (N_23974,N_15487,N_17884);
and U23975 (N_23975,N_14110,N_13087);
and U23976 (N_23976,N_17984,N_12587);
xor U23977 (N_23977,N_12429,N_12104);
and U23978 (N_23978,N_12324,N_17888);
and U23979 (N_23979,N_15943,N_13562);
nor U23980 (N_23980,N_17650,N_13813);
nor U23981 (N_23981,N_13130,N_15845);
and U23982 (N_23982,N_15438,N_13782);
nand U23983 (N_23983,N_15890,N_12052);
xnor U23984 (N_23984,N_16700,N_17950);
or U23985 (N_23985,N_15492,N_13628);
or U23986 (N_23986,N_13414,N_14754);
or U23987 (N_23987,N_14492,N_14868);
and U23988 (N_23988,N_13934,N_14010);
nor U23989 (N_23989,N_16308,N_12203);
nand U23990 (N_23990,N_14394,N_15556);
and U23991 (N_23991,N_17234,N_15537);
nand U23992 (N_23992,N_15045,N_13591);
or U23993 (N_23993,N_16939,N_16990);
nand U23994 (N_23994,N_13476,N_12162);
xor U23995 (N_23995,N_17045,N_15539);
nand U23996 (N_23996,N_17315,N_15039);
nor U23997 (N_23997,N_15335,N_13905);
and U23998 (N_23998,N_12453,N_12474);
or U23999 (N_23999,N_12832,N_14813);
nor U24000 (N_24000,N_19564,N_23399);
nor U24001 (N_24001,N_21166,N_21237);
nand U24002 (N_24002,N_20427,N_20835);
and U24003 (N_24003,N_19918,N_20606);
nand U24004 (N_24004,N_23970,N_18180);
nor U24005 (N_24005,N_21854,N_22041);
nor U24006 (N_24006,N_21786,N_19230);
nor U24007 (N_24007,N_18395,N_21336);
and U24008 (N_24008,N_19605,N_20627);
and U24009 (N_24009,N_23649,N_21094);
xnor U24010 (N_24010,N_22387,N_23595);
nand U24011 (N_24011,N_20203,N_22992);
nor U24012 (N_24012,N_23190,N_18499);
or U24013 (N_24013,N_23237,N_21218);
xnor U24014 (N_24014,N_20008,N_23340);
and U24015 (N_24015,N_22325,N_21012);
and U24016 (N_24016,N_22292,N_21546);
xor U24017 (N_24017,N_23884,N_23570);
nand U24018 (N_24018,N_19124,N_21531);
nor U24019 (N_24019,N_20936,N_18422);
and U24020 (N_24020,N_19917,N_19031);
nor U24021 (N_24021,N_23529,N_18935);
or U24022 (N_24022,N_18910,N_20505);
nor U24023 (N_24023,N_21517,N_20320);
nand U24024 (N_24024,N_18457,N_20634);
nand U24025 (N_24025,N_19509,N_19270);
nand U24026 (N_24026,N_19075,N_23087);
nor U24027 (N_24027,N_23413,N_20115);
nand U24028 (N_24028,N_18654,N_18617);
nand U24029 (N_24029,N_21378,N_22967);
and U24030 (N_24030,N_18397,N_23184);
nand U24031 (N_24031,N_20804,N_22432);
or U24032 (N_24032,N_21911,N_23779);
or U24033 (N_24033,N_20228,N_18951);
and U24034 (N_24034,N_19303,N_18193);
or U24035 (N_24035,N_18791,N_21916);
nand U24036 (N_24036,N_19851,N_21945);
and U24037 (N_24037,N_18950,N_19544);
or U24038 (N_24038,N_20418,N_23060);
and U24039 (N_24039,N_20177,N_18043);
or U24040 (N_24040,N_23989,N_22035);
and U24041 (N_24041,N_18414,N_19915);
or U24042 (N_24042,N_23279,N_18773);
or U24043 (N_24043,N_21329,N_21678);
xor U24044 (N_24044,N_20692,N_22364);
and U24045 (N_24045,N_20886,N_21015);
nor U24046 (N_24046,N_19956,N_18735);
or U24047 (N_24047,N_19870,N_22481);
or U24048 (N_24048,N_23180,N_23376);
nor U24049 (N_24049,N_19937,N_19485);
or U24050 (N_24050,N_22268,N_21668);
nand U24051 (N_24051,N_23611,N_18251);
nor U24052 (N_24052,N_22779,N_19638);
or U24053 (N_24053,N_23941,N_23113);
or U24054 (N_24054,N_18530,N_22100);
xnor U24055 (N_24055,N_19041,N_19855);
and U24056 (N_24056,N_23815,N_20545);
nand U24057 (N_24057,N_23912,N_18974);
nand U24058 (N_24058,N_23211,N_20376);
nand U24059 (N_24059,N_22142,N_23107);
nand U24060 (N_24060,N_20913,N_23037);
xnor U24061 (N_24061,N_20417,N_23579);
or U24062 (N_24062,N_22530,N_19218);
nand U24063 (N_24063,N_20154,N_18799);
and U24064 (N_24064,N_19080,N_22395);
xor U24065 (N_24065,N_23913,N_22319);
nand U24066 (N_24066,N_20725,N_22653);
xnor U24067 (N_24067,N_19531,N_18917);
nor U24068 (N_24068,N_20586,N_23103);
nand U24069 (N_24069,N_23303,N_22183);
or U24070 (N_24070,N_19579,N_19740);
or U24071 (N_24071,N_19405,N_21346);
nand U24072 (N_24072,N_19322,N_18229);
and U24073 (N_24073,N_20617,N_22808);
nor U24074 (N_24074,N_20868,N_18416);
and U24075 (N_24075,N_22554,N_20910);
and U24076 (N_24076,N_22289,N_19970);
or U24077 (N_24077,N_19827,N_20731);
and U24078 (N_24078,N_22636,N_19109);
or U24079 (N_24079,N_23699,N_23806);
xnor U24080 (N_24080,N_20141,N_18287);
nand U24081 (N_24081,N_21367,N_19380);
and U24082 (N_24082,N_22553,N_18324);
and U24083 (N_24083,N_21172,N_18083);
nand U24084 (N_24084,N_23293,N_20399);
or U24085 (N_24085,N_20445,N_19002);
xor U24086 (N_24086,N_21110,N_23864);
xnor U24087 (N_24087,N_19342,N_23814);
nor U24088 (N_24088,N_23337,N_20718);
or U24089 (N_24089,N_19326,N_23232);
nor U24090 (N_24090,N_19185,N_22830);
and U24091 (N_24091,N_18884,N_23607);
xnor U24092 (N_24092,N_22472,N_23536);
nor U24093 (N_24093,N_22823,N_22220);
xnor U24094 (N_24094,N_18730,N_23901);
nand U24095 (N_24095,N_20357,N_22737);
xor U24096 (N_24096,N_20799,N_22958);
xor U24097 (N_24097,N_22144,N_18621);
nor U24098 (N_24098,N_23763,N_23485);
or U24099 (N_24099,N_19823,N_18212);
nand U24100 (N_24100,N_19099,N_18993);
or U24101 (N_24101,N_19262,N_23267);
and U24102 (N_24102,N_18127,N_19719);
or U24103 (N_24103,N_21271,N_19162);
nand U24104 (N_24104,N_18693,N_22694);
nand U24105 (N_24105,N_20447,N_20474);
or U24106 (N_24106,N_21883,N_23550);
and U24107 (N_24107,N_21259,N_18233);
nor U24108 (N_24108,N_18075,N_22590);
xnor U24109 (N_24109,N_18157,N_21936);
xor U24110 (N_24110,N_19690,N_18132);
nor U24111 (N_24111,N_18204,N_18632);
xor U24112 (N_24112,N_20512,N_19669);
or U24113 (N_24113,N_22264,N_19046);
xnor U24114 (N_24114,N_19814,N_19140);
nor U24115 (N_24115,N_20922,N_22470);
xor U24116 (N_24116,N_20079,N_21908);
or U24117 (N_24117,N_22434,N_22887);
nand U24118 (N_24118,N_22114,N_23934);
and U24119 (N_24119,N_18506,N_22329);
xnor U24120 (N_24120,N_20925,N_19428);
nand U24121 (N_24121,N_19298,N_18986);
nor U24122 (N_24122,N_20233,N_21593);
nor U24123 (N_24123,N_19141,N_23472);
xor U24124 (N_24124,N_18943,N_21143);
nor U24125 (N_24125,N_19734,N_23790);
or U24126 (N_24126,N_21302,N_20096);
and U24127 (N_24127,N_19292,N_21009);
nor U24128 (N_24128,N_21024,N_22520);
nand U24129 (N_24129,N_21974,N_22485);
xor U24130 (N_24130,N_18994,N_23667);
xor U24131 (N_24131,N_20746,N_21348);
or U24132 (N_24132,N_20011,N_23247);
or U24133 (N_24133,N_19453,N_23004);
nand U24134 (N_24134,N_23044,N_19567);
nand U24135 (N_24135,N_19639,N_21867);
xnor U24136 (N_24136,N_23036,N_18758);
or U24137 (N_24137,N_20950,N_22056);
xnor U24138 (N_24138,N_19264,N_23646);
xnor U24139 (N_24139,N_21553,N_20733);
or U24140 (N_24140,N_18946,N_22326);
xor U24141 (N_24141,N_20431,N_23029);
nor U24142 (N_24142,N_21428,N_21649);
nand U24143 (N_24143,N_21653,N_22858);
nand U24144 (N_24144,N_19004,N_20422);
xor U24145 (N_24145,N_22189,N_22774);
and U24146 (N_24146,N_20728,N_18505);
nand U24147 (N_24147,N_21938,N_21356);
nand U24148 (N_24148,N_20498,N_18307);
xnor U24149 (N_24149,N_23923,N_22012);
or U24150 (N_24150,N_20194,N_22250);
xnor U24151 (N_24151,N_23842,N_23961);
nor U24152 (N_24152,N_22904,N_20871);
and U24153 (N_24153,N_23980,N_18332);
or U24154 (N_24154,N_21611,N_18515);
xor U24155 (N_24155,N_20252,N_20712);
nand U24156 (N_24156,N_22061,N_18823);
or U24157 (N_24157,N_19542,N_23697);
nor U24158 (N_24158,N_22037,N_20919);
nand U24159 (N_24159,N_23603,N_23694);
nand U24160 (N_24160,N_22913,N_21158);
or U24161 (N_24161,N_22049,N_22938);
nor U24162 (N_24162,N_19729,N_18190);
nor U24163 (N_24163,N_19954,N_22154);
nor U24164 (N_24164,N_22151,N_20864);
nor U24165 (N_24165,N_22436,N_21038);
xor U24166 (N_24166,N_22489,N_21028);
nor U24167 (N_24167,N_19809,N_20277);
nor U24168 (N_24168,N_21568,N_23296);
nor U24169 (N_24169,N_18074,N_20016);
nand U24170 (N_24170,N_18286,N_21328);
xnor U24171 (N_24171,N_21864,N_20684);
and U24172 (N_24172,N_22131,N_19043);
xor U24173 (N_24173,N_19744,N_21692);
or U24174 (N_24174,N_20259,N_22815);
nor U24175 (N_24175,N_21682,N_18488);
nand U24176 (N_24176,N_20109,N_23454);
nand U24177 (N_24177,N_20494,N_19817);
nor U24178 (N_24178,N_21697,N_23449);
nand U24179 (N_24179,N_21787,N_22098);
nand U24180 (N_24180,N_23555,N_19867);
or U24181 (N_24181,N_23991,N_18375);
xnor U24182 (N_24182,N_21065,N_21156);
and U24183 (N_24183,N_22486,N_22316);
nand U24184 (N_24184,N_22706,N_22716);
nand U24185 (N_24185,N_21552,N_23498);
nor U24186 (N_24186,N_22816,N_22454);
xor U24187 (N_24187,N_20608,N_21098);
and U24188 (N_24188,N_20981,N_18152);
xor U24189 (N_24189,N_23447,N_23756);
nand U24190 (N_24190,N_22674,N_23151);
nand U24191 (N_24191,N_19806,N_22864);
and U24192 (N_24192,N_20467,N_18339);
and U24193 (N_24193,N_21320,N_23895);
nand U24194 (N_24194,N_20317,N_18856);
nor U24195 (N_24195,N_21985,N_22615);
nand U24196 (N_24196,N_18020,N_21144);
and U24197 (N_24197,N_23424,N_23751);
and U24198 (N_24198,N_20645,N_22259);
xor U24199 (N_24199,N_23880,N_20076);
nor U24200 (N_24200,N_18766,N_18807);
nor U24201 (N_24201,N_22310,N_22258);
and U24202 (N_24202,N_22267,N_22241);
and U24203 (N_24203,N_19939,N_18126);
nand U24204 (N_24204,N_18098,N_21270);
and U24205 (N_24205,N_22060,N_19157);
xnor U24206 (N_24206,N_20538,N_18360);
xnor U24207 (N_24207,N_22009,N_23355);
and U24208 (N_24208,N_20290,N_20003);
or U24209 (N_24209,N_22537,N_23334);
nand U24210 (N_24210,N_18689,N_21630);
nor U24211 (N_24211,N_18809,N_23266);
xnor U24212 (N_24212,N_18039,N_19343);
nand U24213 (N_24213,N_23415,N_19120);
or U24214 (N_24214,N_18596,N_18409);
nor U24215 (N_24215,N_18443,N_22602);
nor U24216 (N_24216,N_22668,N_20705);
or U24217 (N_24217,N_19330,N_23503);
nor U24218 (N_24218,N_23617,N_18990);
and U24219 (N_24219,N_22357,N_20900);
and U24220 (N_24220,N_23028,N_21563);
or U24221 (N_24221,N_21388,N_19183);
nor U24222 (N_24222,N_22286,N_21776);
nand U24223 (N_24223,N_20116,N_22788);
xnor U24224 (N_24224,N_20311,N_22599);
xor U24225 (N_24225,N_18805,N_23688);
nor U24226 (N_24226,N_21241,N_23621);
nand U24227 (N_24227,N_18925,N_22327);
and U24228 (N_24228,N_19214,N_21970);
xor U24229 (N_24229,N_20558,N_21121);
or U24230 (N_24230,N_20722,N_20535);
nor U24231 (N_24231,N_19250,N_23304);
nor U24232 (N_24232,N_23145,N_22547);
nor U24233 (N_24233,N_23024,N_22299);
nand U24234 (N_24234,N_19777,N_22153);
or U24235 (N_24235,N_20476,N_20240);
nor U24236 (N_24236,N_18260,N_19435);
and U24237 (N_24237,N_18836,N_18522);
and U24238 (N_24238,N_20126,N_18210);
nand U24239 (N_24239,N_22617,N_22200);
and U24240 (N_24240,N_21853,N_22851);
or U24241 (N_24241,N_20093,N_19008);
nand U24242 (N_24242,N_20069,N_19221);
nand U24243 (N_24243,N_22384,N_22118);
nor U24244 (N_24244,N_21227,N_21193);
nand U24245 (N_24245,N_18037,N_22017);
and U24246 (N_24246,N_20752,N_23322);
nand U24247 (N_24247,N_21554,N_21751);
nand U24248 (N_24248,N_20081,N_20193);
nand U24249 (N_24249,N_22048,N_18289);
nor U24250 (N_24250,N_22024,N_23983);
or U24251 (N_24251,N_23807,N_18697);
xor U24252 (N_24252,N_18338,N_18761);
nand U24253 (N_24253,N_23213,N_22165);
xor U24254 (N_24254,N_23039,N_20807);
and U24255 (N_24255,N_19305,N_22548);
xor U24256 (N_24256,N_22229,N_18391);
and U24257 (N_24257,N_23226,N_23684);
or U24258 (N_24258,N_23246,N_23335);
or U24259 (N_24259,N_22338,N_21459);
nor U24260 (N_24260,N_23050,N_21284);
nor U24261 (N_24261,N_20611,N_23312);
nand U24262 (N_24262,N_23222,N_22457);
and U24263 (N_24263,N_20878,N_19796);
xor U24264 (N_24264,N_20456,N_21131);
and U24265 (N_24265,N_19643,N_22586);
nor U24266 (N_24266,N_21572,N_19735);
xor U24267 (N_24267,N_22452,N_23174);
nand U24268 (N_24268,N_18803,N_20686);
and U24269 (N_24269,N_20411,N_18036);
and U24270 (N_24270,N_18057,N_23288);
xnor U24271 (N_24271,N_22235,N_18924);
nor U24272 (N_24272,N_20734,N_19038);
nand U24273 (N_24273,N_18282,N_22881);
nand U24274 (N_24274,N_22570,N_18553);
and U24275 (N_24275,N_23695,N_23223);
or U24276 (N_24276,N_18585,N_23818);
xor U24277 (N_24277,N_21780,N_19786);
and U24278 (N_24278,N_21642,N_20590);
xnor U24279 (N_24279,N_19582,N_19783);
or U24280 (N_24280,N_19894,N_19064);
and U24281 (N_24281,N_19123,N_19922);
and U24282 (N_24282,N_19266,N_18861);
nor U24283 (N_24283,N_19396,N_19180);
nor U24284 (N_24284,N_22574,N_20205);
or U24285 (N_24285,N_22919,N_18200);
or U24286 (N_24286,N_21551,N_19442);
nor U24287 (N_24287,N_20148,N_18403);
or U24288 (N_24288,N_23346,N_19146);
xor U24289 (N_24289,N_18318,N_18093);
nand U24290 (N_24290,N_19773,N_21993);
or U24291 (N_24291,N_19408,N_22841);
nor U24292 (N_24292,N_22149,N_22960);
and U24293 (N_24293,N_22856,N_23609);
nor U24294 (N_24294,N_22260,N_19682);
and U24295 (N_24295,N_20513,N_22367);
nand U24296 (N_24296,N_21375,N_22193);
nand U24297 (N_24297,N_21033,N_23871);
and U24298 (N_24298,N_19009,N_23351);
nand U24299 (N_24299,N_19495,N_20939);
nand U24300 (N_24300,N_21994,N_19226);
and U24301 (N_24301,N_21170,N_18818);
nand U24302 (N_24302,N_22604,N_21749);
or U24303 (N_24303,N_21929,N_23420);
or U24304 (N_24304,N_23844,N_20469);
and U24305 (N_24305,N_19033,N_23275);
or U24306 (N_24306,N_20741,N_19054);
xor U24307 (N_24307,N_21408,N_19143);
nand U24308 (N_24308,N_22585,N_19358);
nand U24309 (N_24309,N_20443,N_21973);
and U24310 (N_24310,N_23566,N_22109);
xor U24311 (N_24311,N_20363,N_18062);
xnor U24312 (N_24312,N_19699,N_22766);
and U24313 (N_24313,N_23701,N_22022);
xnor U24314 (N_24314,N_22820,N_20649);
and U24315 (N_24315,N_21792,N_23832);
nor U24316 (N_24316,N_23101,N_19134);
nor U24317 (N_24317,N_19793,N_20837);
nor U24318 (N_24318,N_19001,N_20560);
or U24319 (N_24319,N_20313,N_23797);
xnor U24320 (N_24320,N_22639,N_18145);
nor U24321 (N_24321,N_21562,N_19594);
nor U24322 (N_24322,N_20224,N_19612);
xor U24323 (N_24323,N_21747,N_20364);
nor U24324 (N_24324,N_23557,N_19858);
or U24325 (N_24325,N_21855,N_19020);
nand U24326 (N_24326,N_20596,N_23966);
nand U24327 (N_24327,N_21123,N_18970);
xnor U24328 (N_24328,N_21183,N_22971);
xnor U24329 (N_24329,N_19965,N_18405);
nor U24330 (N_24330,N_18273,N_19562);
and U24331 (N_24331,N_23169,N_23388);
and U24332 (N_24332,N_23347,N_21243);
nand U24333 (N_24333,N_22518,N_22630);
or U24334 (N_24334,N_20124,N_23629);
nor U24335 (N_24335,N_23090,N_18812);
nor U24336 (N_24336,N_19834,N_20312);
nor U24337 (N_24337,N_18320,N_23928);
xor U24338 (N_24338,N_21891,N_22651);
nand U24339 (N_24339,N_18568,N_21721);
nand U24340 (N_24340,N_18578,N_20037);
nand U24341 (N_24341,N_22199,N_22622);
and U24342 (N_24342,N_22893,N_20186);
nor U24343 (N_24343,N_18070,N_23625);
nand U24344 (N_24344,N_20263,N_21606);
nand U24345 (N_24345,N_21216,N_22691);
xor U24346 (N_24346,N_18830,N_22923);
or U24347 (N_24347,N_21413,N_22693);
or U24348 (N_24348,N_18552,N_23762);
and U24349 (N_24349,N_21050,N_21924);
nand U24350 (N_24350,N_23839,N_18468);
nor U24351 (N_24351,N_18446,N_21789);
nand U24352 (N_24352,N_22420,N_19362);
and U24353 (N_24353,N_21545,N_23782);
xor U24354 (N_24354,N_22006,N_19245);
xnor U24355 (N_24355,N_18866,N_19136);
and U24356 (N_24356,N_22989,N_21420);
and U24357 (N_24357,N_22112,N_20958);
nor U24358 (N_24358,N_23968,N_19836);
xor U24359 (N_24359,N_22296,N_18016);
nand U24360 (N_24360,N_23545,N_18458);
nand U24361 (N_24361,N_23280,N_20636);
nand U24362 (N_24362,N_23637,N_23785);
nand U24363 (N_24363,N_23808,N_21447);
nor U24364 (N_24364,N_19551,N_22102);
nand U24365 (N_24365,N_18721,N_18312);
nor U24366 (N_24366,N_21174,N_19527);
or U24367 (N_24367,N_22107,N_23058);
nor U24368 (N_24368,N_20726,N_19830);
xnor U24369 (N_24369,N_23330,N_18448);
nand U24370 (N_24370,N_19339,N_23273);
and U24371 (N_24371,N_22792,N_21369);
nand U24372 (N_24372,N_21700,N_18663);
or U24373 (N_24373,N_20867,N_18218);
nor U24374 (N_24374,N_19584,N_20202);
and U24375 (N_24375,N_21213,N_21526);
nand U24376 (N_24376,N_18001,N_20007);
nand U24377 (N_24377,N_19062,N_23329);
xnor U24378 (N_24378,N_23276,N_18412);
xnor U24379 (N_24379,N_19187,N_21229);
xor U24380 (N_24380,N_18288,N_21814);
or U24381 (N_24381,N_18971,N_23064);
and U24382 (N_24382,N_20907,N_23048);
nor U24383 (N_24383,N_23965,N_19170);
xnor U24384 (N_24384,N_23234,N_23540);
xor U24385 (N_24385,N_20437,N_23401);
nand U24386 (N_24386,N_20276,N_21273);
nor U24387 (N_24387,N_19371,N_18460);
nand U24388 (N_24388,N_19952,N_19241);
nand U24389 (N_24389,N_21454,N_20928);
nor U24390 (N_24390,N_21724,N_21533);
nand U24391 (N_24391,N_23628,N_20583);
nand U24392 (N_24392,N_23619,N_21397);
or U24393 (N_24393,N_19249,N_23430);
nor U24394 (N_24394,N_22765,N_20325);
xnor U24395 (N_24395,N_19477,N_23474);
nor U24396 (N_24396,N_18741,N_20406);
xor U24397 (N_24397,N_21952,N_20189);
and U24398 (N_24398,N_23892,N_20176);
nand U24399 (N_24399,N_18017,N_22770);
and U24400 (N_24400,N_20542,N_20239);
xor U24401 (N_24401,N_19701,N_20698);
or U24402 (N_24402,N_23686,N_21569);
and U24403 (N_24403,N_20802,N_22842);
or U24404 (N_24404,N_21659,N_23944);
nand U24405 (N_24405,N_19171,N_23236);
or U24406 (N_24406,N_19720,N_20812);
and U24407 (N_24407,N_20945,N_19596);
and U24408 (N_24408,N_18536,N_21890);
nand U24409 (N_24409,N_22915,N_20553);
and U24410 (N_24410,N_22380,N_19805);
nand U24411 (N_24411,N_20012,N_23171);
xor U24412 (N_24412,N_19387,N_23668);
and U24413 (N_24413,N_20816,N_22576);
xnor U24414 (N_24414,N_22218,N_20314);
nand U24415 (N_24415,N_20316,N_18782);
xnor U24416 (N_24416,N_22888,N_21231);
and U24417 (N_24417,N_18216,N_18878);
nand U24418 (N_24418,N_20876,N_21394);
nand U24419 (N_24419,N_21385,N_20036);
nor U24420 (N_24420,N_23719,N_23176);
xor U24421 (N_24421,N_23217,N_22934);
or U24422 (N_24422,N_21307,N_19932);
nor U24423 (N_24423,N_21169,N_23243);
nand U24424 (N_24424,N_23375,N_18294);
and U24425 (N_24425,N_19654,N_20770);
or U24426 (N_24426,N_20405,N_19439);
xnor U24427 (N_24427,N_18211,N_22275);
nand U24428 (N_24428,N_19570,N_23948);
xor U24429 (N_24429,N_18816,N_21550);
xnor U24430 (N_24430,N_20860,N_21130);
and U24431 (N_24431,N_22983,N_23526);
nand U24432 (N_24432,N_20173,N_23716);
and U24433 (N_24433,N_19552,N_21171);
nand U24434 (N_24434,N_21008,N_22129);
and U24435 (N_24435,N_22391,N_22369);
or U24436 (N_24436,N_21304,N_20488);
or U24437 (N_24437,N_19118,N_18482);
or U24438 (N_24438,N_19706,N_23891);
or U24439 (N_24439,N_22378,N_19090);
nor U24440 (N_24440,N_19961,N_23434);
nand U24441 (N_24441,N_21773,N_23554);
or U24442 (N_24442,N_19422,N_22984);
and U24443 (N_24443,N_19328,N_20279);
nand U24444 (N_24444,N_22158,N_21948);
nand U24445 (N_24445,N_18723,N_21523);
and U24446 (N_24446,N_20099,N_21440);
nand U24447 (N_24447,N_21694,N_23473);
or U24448 (N_24448,N_21333,N_18349);
nand U24449 (N_24449,N_23938,N_22105);
and U24450 (N_24450,N_19991,N_22584);
nand U24451 (N_24451,N_19747,N_18641);
nor U24452 (N_24452,N_23314,N_20057);
and U24453 (N_24453,N_19285,N_20221);
and U24454 (N_24454,N_18315,N_19061);
xor U24455 (N_24455,N_19280,N_18259);
or U24456 (N_24456,N_19843,N_22627);
or U24457 (N_24457,N_21238,N_19731);
and U24458 (N_24458,N_18980,N_20960);
xnor U24459 (N_24459,N_20132,N_23588);
nor U24460 (N_24460,N_19693,N_22127);
or U24461 (N_24461,N_19333,N_21019);
nand U24462 (N_24462,N_19933,N_19896);
and U24463 (N_24463,N_22880,N_18771);
xor U24464 (N_24464,N_22536,N_21456);
and U24465 (N_24465,N_19920,N_18840);
or U24466 (N_24466,N_19897,N_21029);
and U24467 (N_24467,N_23433,N_21357);
nor U24468 (N_24468,N_18793,N_23732);
nand U24469 (N_24469,N_20102,N_19178);
nand U24470 (N_24470,N_23192,N_23874);
or U24471 (N_24471,N_22379,N_20080);
or U24472 (N_24472,N_23417,N_18274);
nor U24473 (N_24473,N_18746,N_22981);
and U24474 (N_24474,N_18120,N_23126);
and U24475 (N_24475,N_23073,N_20211);
nand U24476 (N_24476,N_18196,N_20333);
or U24477 (N_24477,N_23518,N_20874);
and U24478 (N_24478,N_22262,N_21757);
nand U24479 (N_24479,N_18533,N_18804);
nor U24480 (N_24480,N_18507,N_18290);
nor U24481 (N_24481,N_20744,N_20940);
or U24482 (N_24482,N_21232,N_21371);
xor U24483 (N_24483,N_21645,N_18295);
or U24484 (N_24484,N_19378,N_20366);
nand U24485 (N_24485,N_23661,N_23746);
nand U24486 (N_24486,N_23946,N_19801);
and U24487 (N_24487,N_18539,N_22117);
nand U24488 (N_24488,N_19026,N_23918);
nor U24489 (N_24489,N_23670,N_21595);
nor U24490 (N_24490,N_23610,N_21667);
nand U24491 (N_24491,N_18447,N_23469);
nor U24492 (N_24492,N_22874,N_20817);
xor U24493 (N_24493,N_20509,N_19127);
nor U24494 (N_24494,N_20776,N_23104);
nor U24495 (N_24495,N_18995,N_23497);
nor U24496 (N_24496,N_18165,N_20040);
nor U24497 (N_24497,N_21795,N_21124);
nand U24498 (N_24498,N_18267,N_20209);
nand U24499 (N_24499,N_23193,N_23949);
xor U24500 (N_24500,N_19194,N_22705);
or U24501 (N_24501,N_23428,N_18979);
nand U24502 (N_24502,N_19510,N_18313);
and U24503 (N_24503,N_21465,N_19037);
xor U24504 (N_24504,N_23527,N_23572);
nor U24505 (N_24505,N_21961,N_22445);
or U24506 (N_24506,N_20688,N_23200);
nor U24507 (N_24507,N_21374,N_23616);
nand U24508 (N_24508,N_20433,N_22795);
and U24509 (N_24509,N_18658,N_23679);
xor U24510 (N_24510,N_19163,N_23634);
or U24511 (N_24511,N_19637,N_21234);
or U24512 (N_24512,N_18779,N_20604);
nand U24513 (N_24513,N_19168,N_19164);
and U24514 (N_24514,N_21023,N_23602);
and U24515 (N_24515,N_21382,N_21959);
xnor U24516 (N_24516,N_23414,N_23581);
or U24517 (N_24517,N_20091,N_22336);
and U24518 (N_24518,N_19425,N_22213);
nand U24519 (N_24519,N_19846,N_20014);
and U24520 (N_24520,N_22001,N_19269);
xor U24521 (N_24521,N_19018,N_22964);
nand U24522 (N_24522,N_18371,N_21090);
and U24523 (N_24523,N_21186,N_21340);
nor U24524 (N_24524,N_22632,N_20678);
or U24525 (N_24525,N_22206,N_20372);
or U24526 (N_24526,N_22561,N_21717);
and U24527 (N_24527,N_18292,N_20163);
nand U24528 (N_24528,N_18636,N_20888);
or U24529 (N_24529,N_18759,N_20550);
xnor U24530 (N_24530,N_22361,N_19407);
xnor U24531 (N_24531,N_23747,N_22284);
xor U24532 (N_24532,N_21257,N_20555);
xnor U24533 (N_24533,N_18478,N_22195);
xor U24534 (N_24534,N_23191,N_21954);
nand U24535 (N_24535,N_18203,N_19674);
and U24536 (N_24536,N_19723,N_20135);
nand U24537 (N_24537,N_20423,N_22175);
nand U24538 (N_24538,N_20282,N_20631);
xnor U24539 (N_24539,N_20735,N_22473);
and U24540 (N_24540,N_23046,N_18595);
xnor U24541 (N_24541,N_23522,N_23402);
xnor U24542 (N_24542,N_22735,N_21149);
nand U24543 (N_24543,N_19263,N_21969);
nand U24544 (N_24544,N_19537,N_21198);
or U24545 (N_24545,N_22494,N_23467);
xnor U24546 (N_24546,N_18387,N_18579);
or U24547 (N_24547,N_19889,N_18930);
nand U24548 (N_24548,N_23565,N_22052);
or U24549 (N_24549,N_23040,N_23863);
nand U24550 (N_24550,N_20070,N_22468);
xor U24551 (N_24551,N_18453,N_19190);
or U24552 (N_24552,N_18545,N_22318);
and U24553 (N_24553,N_22607,N_22665);
nand U24554 (N_24554,N_18509,N_19198);
and U24555 (N_24555,N_23905,N_22558);
nor U24556 (N_24556,N_21529,N_20319);
nand U24557 (N_24557,N_23410,N_18726);
and U24558 (N_24558,N_19790,N_22970);
xor U24559 (N_24559,N_20997,N_20870);
nor U24560 (N_24560,N_23035,N_18486);
or U24561 (N_24561,N_19707,N_21861);
nand U24562 (N_24562,N_20323,N_19361);
nor U24563 (N_24563,N_19591,N_21949);
nor U24564 (N_24564,N_23031,N_18982);
and U24565 (N_24565,N_20536,N_18845);
nor U24566 (N_24566,N_21242,N_23010);
xnor U24567 (N_24567,N_20480,N_23997);
and U24568 (N_24568,N_20496,N_23173);
or U24569 (N_24569,N_18018,N_22323);
nor U24570 (N_24570,N_18705,N_22311);
nand U24571 (N_24571,N_18650,N_23767);
nand U24572 (N_24572,N_19513,N_19538);
nand U24573 (N_24573,N_18082,N_19875);
nand U24574 (N_24574,N_21574,N_18644);
nand U24575 (N_24575,N_22315,N_21519);
or U24576 (N_24576,N_21881,N_21132);
and U24577 (N_24577,N_20889,N_20425);
xnor U24578 (N_24578,N_18657,N_20961);
and U24579 (N_24579,N_21681,N_19866);
nand U24580 (N_24580,N_19755,N_18813);
xnor U24581 (N_24581,N_20167,N_18306);
and U24582 (N_24582,N_20460,N_19458);
xor U24583 (N_24583,N_22020,N_20212);
and U24584 (N_24584,N_19621,N_21699);
nand U24585 (N_24585,N_23408,N_19975);
nand U24586 (N_24586,N_21104,N_19691);
or U24587 (N_24587,N_23462,N_23437);
and U24588 (N_24588,N_20648,N_20621);
or U24589 (N_24589,N_23974,N_20507);
or U24590 (N_24590,N_22654,N_20395);
nand U24591 (N_24591,N_20121,N_19312);
and U24592 (N_24592,N_18770,N_23198);
xor U24593 (N_24593,N_23284,N_19880);
or U24594 (N_24594,N_23504,N_20006);
and U24595 (N_24595,N_22689,N_21946);
or U24596 (N_24596,N_20344,N_18173);
and U24597 (N_24597,N_21312,N_20017);
and U24598 (N_24598,N_23368,N_21332);
nor U24599 (N_24599,N_23560,N_21311);
or U24600 (N_24600,N_19174,N_23696);
nand U24601 (N_24601,N_20814,N_23812);
nand U24602 (N_24602,N_23843,N_18413);
and U24603 (N_24603,N_20937,N_18379);
or U24604 (N_24604,N_20353,N_23112);
xor U24605 (N_24605,N_22302,N_19093);
or U24606 (N_24606,N_18562,N_19475);
and U24607 (N_24607,N_22279,N_23723);
and U24608 (N_24608,N_22464,N_21042);
xnor U24609 (N_24609,N_20715,N_22976);
xnor U24610 (N_24610,N_20387,N_21522);
or U24611 (N_24611,N_18377,N_19525);
nor U24612 (N_24612,N_20582,N_19186);
and U24613 (N_24613,N_23737,N_20779);
and U24614 (N_24614,N_23867,N_18439);
nand U24615 (N_24615,N_21148,N_21693);
and U24616 (N_24616,N_21249,N_20528);
xnor U24617 (N_24617,N_19329,N_22675);
nor U24618 (N_24618,N_21405,N_18842);
nor U24619 (N_24619,N_20440,N_18541);
or U24620 (N_24620,N_18280,N_23537);
nor U24621 (N_24621,N_23272,N_19990);
xnor U24622 (N_24622,N_19217,N_19718);
nand U24623 (N_24623,N_19753,N_23196);
nand U24624 (N_24624,N_20019,N_19024);
nand U24625 (N_24625,N_21233,N_21000);
and U24626 (N_24626,N_23911,N_20515);
or U24627 (N_24627,N_21915,N_18690);
or U24628 (N_24628,N_19842,N_23549);
nand U24629 (N_24629,N_18665,N_21942);
and U24630 (N_24630,N_21100,N_20162);
nand U24631 (N_24631,N_23998,N_23558);
or U24632 (N_24632,N_21820,N_20673);
nor U24633 (N_24633,N_22638,N_23956);
nor U24634 (N_24634,N_19374,N_21674);
xnor U24635 (N_24635,N_18646,N_22876);
or U24636 (N_24636,N_20767,N_20021);
xor U24637 (N_24637,N_20855,N_18624);
xor U24638 (N_24638,N_19677,N_21543);
or U24639 (N_24639,N_22399,N_20101);
or U24640 (N_24640,N_22094,N_19808);
nand U24641 (N_24641,N_20959,N_18455);
or U24642 (N_24642,N_22211,N_22034);
xor U24643 (N_24643,N_22825,N_23241);
or U24644 (N_24644,N_21457,N_20832);
or U24645 (N_24645,N_21744,N_23106);
nor U24646 (N_24646,N_22358,N_20973);
or U24647 (N_24647,N_22882,N_20839);
nor U24648 (N_24648,N_19045,N_21011);
and U24649 (N_24649,N_19730,N_22669);
xor U24650 (N_24650,N_18590,N_22059);
or U24651 (N_24651,N_20435,N_23741);
or U24652 (N_24652,N_20740,N_18796);
nand U24653 (N_24653,N_20356,N_19775);
and U24654 (N_24654,N_20650,N_21636);
nor U24655 (N_24655,N_20723,N_20674);
nor U24656 (N_24656,N_22917,N_18164);
nor U24657 (N_24657,N_21676,N_19048);
xor U24658 (N_24658,N_23405,N_22031);
nand U24659 (N_24659,N_20294,N_18005);
nor U24660 (N_24660,N_22110,N_19820);
nand U24661 (N_24661,N_23856,N_21943);
nor U24662 (N_24662,N_19427,N_21598);
xor U24663 (N_24663,N_22298,N_20758);
xnor U24664 (N_24664,N_20690,N_18662);
xor U24665 (N_24665,N_19578,N_20084);
xor U24666 (N_24666,N_22488,N_18808);
and U24667 (N_24667,N_22362,N_21180);
and U24668 (N_24668,N_23754,N_21046);
xor U24669 (N_24669,N_20291,N_22297);
or U24670 (N_24670,N_18030,N_20082);
nand U24671 (N_24671,N_20591,N_22562);
nand U24672 (N_24672,N_20699,N_22943);
xnor U24673 (N_24673,N_19664,N_23664);
nor U24674 (N_24674,N_19518,N_21484);
and U24675 (N_24675,N_19191,N_19641);
nor U24676 (N_24676,N_21415,N_22139);
and U24677 (N_24677,N_23097,N_19919);
nand U24678 (N_24678,N_22071,N_18281);
xnor U24679 (N_24679,N_22348,N_19909);
nor U24680 (N_24680,N_18955,N_20043);
and U24681 (N_24681,N_23444,N_21739);
nor U24682 (N_24682,N_20104,N_19656);
nand U24683 (N_24683,N_20697,N_19353);
or U24684 (N_24684,N_18330,N_21264);
nor U24685 (N_24685,N_21609,N_22428);
or U24686 (N_24686,N_21416,N_19113);
xnor U24687 (N_24687,N_22166,N_19569);
nor U24688 (N_24688,N_19994,N_19478);
xnor U24689 (N_24689,N_20257,N_19989);
or U24690 (N_24690,N_23508,N_21878);
xor U24691 (N_24691,N_23300,N_20465);
nand U24692 (N_24692,N_19778,N_20264);
nand U24693 (N_24693,N_23897,N_22040);
nand U24694 (N_24694,N_20100,N_23630);
nand U24695 (N_24695,N_18713,N_21742);
or U24696 (N_24696,N_21474,N_20230);
and U24697 (N_24697,N_19239,N_22821);
nor U24698 (N_24698,N_23725,N_19240);
nand U24699 (N_24699,N_21809,N_20470);
nand U24700 (N_24700,N_22998,N_23826);
nor U24701 (N_24701,N_22740,N_19053);
nor U24702 (N_24702,N_21847,N_21857);
xor U24703 (N_24703,N_22623,N_20050);
nor U24704 (N_24704,N_21047,N_23418);
nand U24705 (N_24705,N_22363,N_20052);
and U24706 (N_24706,N_19474,N_23137);
and U24707 (N_24707,N_22948,N_22784);
nand U24708 (N_24708,N_21401,N_19927);
and U24709 (N_24709,N_22265,N_23505);
nand U24710 (N_24710,N_21955,N_21267);
nand U24711 (N_24711,N_19450,N_18837);
xnor U24712 (N_24712,N_22047,N_20670);
or U24713 (N_24713,N_19826,N_18423);
and U24714 (N_24714,N_22672,N_20373);
or U24715 (N_24715,N_19593,N_18250);
and U24716 (N_24716,N_22763,N_21778);
and U24717 (N_24717,N_20863,N_23307);
xor U24718 (N_24718,N_18495,N_18874);
and U24719 (N_24719,N_20931,N_21843);
and U24720 (N_24720,N_18901,N_21603);
xnor U24721 (N_24721,N_22167,N_18765);
nand U24722 (N_24722,N_21788,N_18944);
nand U24723 (N_24723,N_22019,N_21726);
xnor U24724 (N_24724,N_18527,N_20062);
and U24725 (N_24725,N_21230,N_19644);
and U24726 (N_24726,N_21912,N_19372);
nand U24727 (N_24727,N_23114,N_21471);
xnor U24728 (N_24728,N_19493,N_19349);
and U24729 (N_24729,N_19623,N_20138);
nor U24730 (N_24730,N_21525,N_21866);
nor U24731 (N_24731,N_22238,N_22818);
nor U24732 (N_24732,N_21246,N_19925);
or U24733 (N_24733,N_20564,N_19815);
and U24734 (N_24734,N_19115,N_21783);
nand U24735 (N_24735,N_23344,N_19971);
and U24736 (N_24736,N_22838,N_22417);
nand U24737 (N_24737,N_21081,N_19144);
nand U24738 (N_24738,N_21322,N_19065);
or U24739 (N_24739,N_23940,N_20227);
nor U24740 (N_24740,N_18134,N_18153);
or U24741 (N_24741,N_19583,N_20478);
nor U24742 (N_24742,N_23115,N_21930);
xnor U24743 (N_24743,N_18909,N_18186);
xor U24744 (N_24744,N_19708,N_23478);
and U24745 (N_24745,N_19577,N_18849);
or U24746 (N_24746,N_20552,N_20075);
xor U24747 (N_24747,N_22531,N_23105);
and U24748 (N_24748,N_22878,N_22104);
nand U24749 (N_24749,N_23915,N_22083);
nor U24750 (N_24750,N_21862,N_19461);
xnor U24751 (N_24751,N_23136,N_18627);
or U24752 (N_24752,N_18417,N_19838);
or U24753 (N_24753,N_18939,N_23506);
nor U24754 (N_24754,N_19074,N_22723);
or U24755 (N_24755,N_23510,N_22780);
or U24756 (N_24756,N_19781,N_18348);
nor U24757 (N_24757,N_23739,N_20309);
xor U24758 (N_24758,N_19368,N_22798);
or U24759 (N_24759,N_18019,N_22597);
or U24760 (N_24760,N_21737,N_19175);
xor U24761 (N_24761,N_23623,N_23567);
nor U24762 (N_24762,N_21536,N_22306);
nand U24763 (N_24763,N_22692,N_21195);
nand U24764 (N_24764,N_20527,N_21317);
xor U24765 (N_24765,N_18870,N_18677);
nand U24766 (N_24766,N_19499,N_23008);
and U24767 (N_24767,N_18222,N_19924);
xnor U24768 (N_24768,N_21805,N_23339);
xnor U24769 (N_24769,N_22640,N_21157);
and U24770 (N_24770,N_19317,N_23085);
xnor U24771 (N_24771,N_18341,N_22121);
nand U24772 (N_24772,N_20916,N_21398);
nand U24773 (N_24773,N_19647,N_21845);
nand U24774 (N_24774,N_19308,N_19608);
and U24775 (N_24775,N_20852,N_23034);
nand U24776 (N_24776,N_19558,N_21587);
nor U24777 (N_24777,N_18326,N_20784);
nor U24778 (N_24778,N_19982,N_22791);
and U24779 (N_24779,N_21118,N_23364);
and U24780 (N_24780,N_23465,N_22710);
or U24781 (N_24781,N_23986,N_22756);
and U24782 (N_24782,N_18183,N_18922);
or U24783 (N_24783,N_20970,N_22717);
nand U24784 (N_24784,N_21872,N_19931);
xnor U24785 (N_24785,N_20451,N_20404);
and U24786 (N_24786,N_19492,N_22164);
or U24787 (N_24787,N_19344,N_18668);
nor U24788 (N_24788,N_22475,N_23932);
nand U24789 (N_24789,N_22307,N_23009);
or U24790 (N_24790,N_19948,N_19626);
or U24791 (N_24791,N_19015,N_21673);
or U24792 (N_24792,N_21537,N_18831);
and U24793 (N_24793,N_18054,N_18077);
or U24794 (N_24794,N_19444,N_23310);
nand U24795 (N_24795,N_22626,N_18291);
nand U24796 (N_24796,N_21764,N_19710);
nand U24797 (N_24797,N_21182,N_18526);
or U24798 (N_24798,N_22972,N_20539);
and U24799 (N_24799,N_23298,N_23639);
or U24800 (N_24800,N_22577,N_20068);
xnor U24801 (N_24801,N_21794,N_20629);
xnor U24802 (N_24802,N_22025,N_20196);
nand U24803 (N_24803,N_19417,N_20382);
or U24804 (N_24804,N_18463,N_20915);
nand U24805 (N_24805,N_20053,N_21001);
nor U24806 (N_24806,N_20551,N_19345);
or U24807 (N_24807,N_20502,N_23372);
nor U24808 (N_24808,N_18108,N_23391);
nor U24809 (N_24809,N_23168,N_21651);
nor U24810 (N_24810,N_20436,N_18792);
nand U24811 (N_24811,N_18821,N_19812);
or U24812 (N_24812,N_20668,N_22986);
nand U24813 (N_24813,N_21984,N_22730);
nand U24814 (N_24814,N_22382,N_21512);
xnor U24815 (N_24815,N_22641,N_22010);
nand U24816 (N_24816,N_21196,N_18672);
nand U24817 (N_24817,N_20859,N_21219);
nand U24818 (N_24818,N_19928,N_18886);
and U24819 (N_24819,N_22505,N_21071);
xnor U24820 (N_24820,N_18087,N_20428);
nor U24821 (N_24821,N_21279,N_19955);
and U24822 (N_24822,N_21431,N_20120);
xnor U24823 (N_24823,N_22517,N_20381);
xor U24824 (N_24824,N_22926,N_22546);
nand U24825 (N_24825,N_23930,N_18960);
nand U24826 (N_24826,N_18927,N_20680);
nor U24827 (N_24827,N_21325,N_22985);
xor U24828 (N_24828,N_19382,N_23082);
nand U24829 (N_24829,N_20769,N_20663);
nand U24830 (N_24830,N_18989,N_23299);
nand U24831 (N_24831,N_19411,N_18130);
or U24832 (N_24832,N_20917,N_21579);
nand U24833 (N_24833,N_21003,N_18168);
xnor U24834 (N_24834,N_23979,N_22239);
xnor U24835 (N_24835,N_18667,N_21514);
xor U24836 (N_24836,N_23922,N_21066);
and U24837 (N_24837,N_20996,N_21448);
nand U24838 (N_24838,N_18128,N_20785);
or U24839 (N_24839,N_19275,N_21806);
or U24840 (N_24840,N_18718,N_22198);
or U24841 (N_24841,N_23450,N_18022);
nand U24842 (N_24842,N_18357,N_18739);
nand U24843 (N_24843,N_21838,N_19100);
nor U24844 (N_24844,N_20466,N_20993);
nand U24845 (N_24845,N_20412,N_21093);
and U24846 (N_24846,N_22069,N_20170);
and U24847 (N_24847,N_23142,N_23062);
or U24848 (N_24848,N_21852,N_18176);
nand U24849 (N_24849,N_21534,N_20568);
and U24850 (N_24850,N_23967,N_20038);
and U24851 (N_24851,N_21585,N_18498);
and U24852 (N_24852,N_20906,N_19646);
or U24853 (N_24853,N_23282,N_19105);
or U24854 (N_24854,N_21829,N_19902);
and U24855 (N_24855,N_22435,N_19094);
xnor U24856 (N_24856,N_21573,N_20628);
or U24857 (N_24857,N_21087,N_23801);
nor U24858 (N_24858,N_21406,N_21575);
xor U24859 (N_24859,N_19943,N_19859);
nand U24860 (N_24860,N_22759,N_18048);
nand U24861 (N_24861,N_22847,N_19484);
nor U24862 (N_24862,N_19346,N_20887);
and U24863 (N_24863,N_19697,N_19766);
xor U24864 (N_24864,N_21190,N_22345);
nand U24865 (N_24865,N_23907,N_18563);
or U24866 (N_24866,N_23359,N_20201);
xnor U24867 (N_24867,N_23914,N_21391);
and U24868 (N_24868,N_21640,N_21168);
xor U24869 (N_24869,N_19392,N_20522);
and U24870 (N_24870,N_19243,N_23571);
or U24871 (N_24871,N_18593,N_21826);
xor U24872 (N_24872,N_23179,N_20289);
nor U24873 (N_24873,N_23258,N_19869);
nor U24874 (N_24874,N_19091,N_18835);
or U24875 (N_24875,N_21899,N_20020);
or U24876 (N_24876,N_19271,N_22389);
and U24877 (N_24877,N_23201,N_22634);
or U24878 (N_24878,N_19536,N_23295);
xnor U24879 (N_24879,N_22073,N_21056);
or U24880 (N_24880,N_22087,N_19614);
xor U24881 (N_24881,N_20074,N_23416);
nor U24882 (N_24882,N_23657,N_18159);
xnor U24883 (N_24883,N_18374,N_19160);
and U24884 (N_24884,N_23371,N_18867);
nand U24885 (N_24885,N_19585,N_20105);
nor U24886 (N_24886,N_20484,N_18449);
xor U24887 (N_24887,N_22568,N_22777);
and U24888 (N_24888,N_19853,N_21184);
nand U24889 (N_24889,N_20687,N_23929);
xnor U24890 (N_24890,N_18666,N_22635);
nand U24891 (N_24891,N_22519,N_19212);
nor U24892 (N_24892,N_19223,N_18826);
nand U24893 (N_24893,N_23144,N_23178);
nand U24894 (N_24894,N_23627,N_20532);
nand U24895 (N_24895,N_22512,N_21505);
nor U24896 (N_24896,N_19910,N_19059);
or U24897 (N_24897,N_23601,N_22169);
nand U24898 (N_24898,N_20441,N_20031);
xnor U24899 (N_24899,N_18041,N_20119);
nand U24900 (N_24900,N_21652,N_19572);
or U24901 (N_24901,N_21932,N_21901);
nand U24902 (N_24902,N_19216,N_18628);
xnor U24903 (N_24903,N_21725,N_19166);
xnor U24904 (N_24904,N_18941,N_23706);
nor U24905 (N_24905,N_23455,N_18104);
or U24906 (N_24906,N_21607,N_18797);
nor U24907 (N_24907,N_23205,N_20396);
or U24908 (N_24908,N_22203,N_23135);
or U24909 (N_24909,N_21502,N_22832);
xor U24910 (N_24910,N_22226,N_18327);
and U24911 (N_24911,N_19005,N_22660);
xor U24912 (N_24912,N_18749,N_23859);
nor U24913 (N_24913,N_20426,N_20403);
nand U24914 (N_24914,N_21167,N_18976);
nand U24915 (N_24915,N_18137,N_19604);
and U24916 (N_24916,N_19883,N_20557);
xnor U24917 (N_24917,N_22819,N_18968);
or U24918 (N_24918,N_19724,N_22111);
or U24919 (N_24919,N_21449,N_19535);
nor U24920 (N_24920,N_23265,N_23524);
nand U24921 (N_24921,N_19964,N_19617);
xor U24922 (N_24922,N_21622,N_21349);
nand U24923 (N_24923,N_18471,N_18733);
xor U24924 (N_24924,N_20982,N_23072);
nor U24925 (N_24925,N_18485,N_21647);
or U24926 (N_24926,N_20329,N_22309);
and U24927 (N_24927,N_18181,N_22522);
nand U24928 (N_24928,N_20543,N_18652);
xnor U24929 (N_24929,N_19252,N_18876);
xor U24930 (N_24930,N_22186,N_21476);
and U24931 (N_24931,N_20639,N_23239);
or U24932 (N_24932,N_21746,N_18501);
nand U24933 (N_24933,N_19548,N_18757);
or U24934 (N_24934,N_20385,N_18985);
or U24935 (N_24935,N_23127,N_22567);
xor U24936 (N_24936,N_23614,N_22564);
nand U24937 (N_24937,N_23776,N_20633);
and U24938 (N_24938,N_18484,N_23220);
and U24939 (N_24939,N_19227,N_22438);
nand U24940 (N_24940,N_18296,N_20630);
nand U24941 (N_24941,N_19169,N_19400);
nor U24942 (N_24942,N_22011,N_20929);
xor U24943 (N_24943,N_20810,N_19414);
and U24944 (N_24944,N_21134,N_22405);
xnor U24945 (N_24945,N_19541,N_22659);
or U24946 (N_24946,N_20851,N_20223);
nand U24947 (N_24947,N_21037,N_21577);
and U24948 (N_24948,N_19923,N_23795);
or U24949 (N_24949,N_19335,N_18121);
or U24950 (N_24950,N_18573,N_23352);
or U24951 (N_24951,N_19364,N_19101);
and U24952 (N_24952,N_18908,N_18383);
nand U24953 (N_24953,N_20340,N_22745);
nor U24954 (N_24954,N_20540,N_21831);
xor U24955 (N_24955,N_21439,N_21210);
and U24956 (N_24956,N_19286,N_20025);
xnor U24957 (N_24957,N_23781,N_18915);
and U24958 (N_24958,N_23404,N_22621);
or U24959 (N_24959,N_18311,N_22592);
and U24960 (N_24960,N_20861,N_21034);
and U24961 (N_24961,N_19052,N_19244);
nor U24962 (N_24962,N_21962,N_20094);
nor U24963 (N_24963,N_18843,N_21926);
nor U24964 (N_24964,N_22843,N_23804);
nor U24965 (N_24965,N_23138,N_19553);
nor U24966 (N_24966,N_23678,N_20004);
nand U24967 (N_24967,N_18963,N_22321);
xor U24968 (N_24968,N_22079,N_18352);
nor U24969 (N_24969,N_20903,N_22032);
or U24970 (N_24970,N_20107,N_18609);
or U24971 (N_24971,N_18437,N_21521);
nand U24972 (N_24972,N_19456,N_19615);
or U24973 (N_24973,N_22991,N_20336);
or U24974 (N_24974,N_18271,N_19694);
nor U24975 (N_24975,N_20879,N_20707);
nor U24976 (N_24976,N_20976,N_22426);
or U24977 (N_24977,N_19630,N_21689);
and U24978 (N_24978,N_18325,N_20738);
nor U24979 (N_24979,N_23095,N_21052);
and U24980 (N_24980,N_23154,N_18433);
nand U24981 (N_24981,N_19236,N_21914);
xor U24982 (N_24982,N_18814,N_21141);
nor U24983 (N_24983,N_19446,N_19206);
or U24984 (N_24984,N_18329,N_21663);
nand U24985 (N_24985,N_20840,N_23140);
or U24986 (N_24986,N_19156,N_19732);
xor U24987 (N_24987,N_23409,N_19995);
xnor U24988 (N_24988,N_18472,N_23872);
or U24989 (N_24989,N_20965,N_21882);
or U24990 (N_24990,N_20108,N_23854);
xor U24991 (N_24991,N_19911,N_20041);
or U24992 (N_24992,N_18147,N_20818);
xor U24993 (N_24993,N_22091,N_19261);
nand U24994 (N_24994,N_21661,N_18857);
nand U24995 (N_24995,N_23001,N_19996);
or U24996 (N_24996,N_21069,N_18513);
nand U24997 (N_24997,N_19769,N_23677);
xnor U24998 (N_24998,N_19650,N_20054);
xnor U24999 (N_24999,N_21113,N_19290);
and U25000 (N_25000,N_18366,N_19248);
or U25001 (N_25001,N_19984,N_22133);
xnor U25002 (N_25002,N_18669,N_20491);
and U25003 (N_25003,N_18774,N_19763);
nor U25004 (N_25004,N_22404,N_19976);
nand U25005 (N_25005,N_19071,N_19782);
and U25006 (N_25006,N_18362,N_21140);
nor U25007 (N_25007,N_22873,N_23546);
xor U25008 (N_25008,N_18477,N_18107);
nand U25009 (N_25009,N_21486,N_23523);
nor U25010 (N_25010,N_18569,N_21877);
nand U25011 (N_25011,N_20315,N_22176);
nand U25012 (N_25012,N_20113,N_20503);
nor U25013 (N_25013,N_20368,N_18481);
nand U25014 (N_25014,N_21584,N_18897);
nor U25015 (N_25015,N_21619,N_18892);
or U25016 (N_25016,N_18706,N_18161);
nor U25017 (N_25017,N_23847,N_20432);
and U25018 (N_25018,N_23568,N_19696);
nand U25019 (N_25019,N_23959,N_19947);
nor U25020 (N_25020,N_22231,N_20199);
xnor U25021 (N_25021,N_22775,N_18462);
or U25022 (N_25022,N_21590,N_20307);
nand U25023 (N_25023,N_23204,N_20623);
nor U25024 (N_25024,N_18113,N_18557);
nand U25025 (N_25025,N_21226,N_19818);
nor U25026 (N_25026,N_18333,N_18776);
xor U25027 (N_25027,N_20458,N_20140);
nand U25028 (N_25028,N_20844,N_19470);
nand U25029 (N_25029,N_19926,N_18715);
nand U25030 (N_25030,N_22368,N_19803);
nand U25031 (N_25031,N_21043,N_20523);
nor U25032 (N_25032,N_22190,N_22587);
xnor U25033 (N_25033,N_21272,N_21445);
nand U25034 (N_25034,N_19432,N_23955);
nor U25035 (N_25035,N_23278,N_18442);
and U25036 (N_25036,N_22746,N_22980);
or U25037 (N_25037,N_19337,N_21931);
or U25038 (N_25038,N_21485,N_22403);
nand U25039 (N_25039,N_22987,N_23484);
xor U25040 (N_25040,N_19798,N_23141);
nand U25041 (N_25041,N_20658,N_18174);
nand U25042 (N_25042,N_18844,N_19029);
and U25043 (N_25043,N_19979,N_19309);
and U25044 (N_25044,N_21458,N_22525);
xnor U25045 (N_25045,N_22503,N_21637);
nor U25046 (N_25046,N_21477,N_18977);
or U25047 (N_25047,N_23166,N_21392);
or U25048 (N_25048,N_22439,N_20923);
nand U25049 (N_25049,N_21053,N_20272);
and U25050 (N_25050,N_22778,N_18264);
or U25051 (N_25051,N_21736,N_19340);
xor U25052 (N_25052,N_22804,N_19871);
xnor U25053 (N_25053,N_23384,N_19519);
and U25054 (N_25054,N_22254,N_19751);
and U25055 (N_25055,N_21723,N_23681);
nor U25056 (N_25056,N_20968,N_18304);
and U25057 (N_25057,N_22698,N_23530);
xnor U25058 (N_25058,N_20957,N_22891);
nand U25059 (N_25059,N_20462,N_20866);
nand U25060 (N_25060,N_21335,N_20214);
xor U25061 (N_25061,N_21129,N_20393);
xor U25062 (N_25062,N_21070,N_21509);
xnor U25063 (N_25063,N_18430,N_21832);
or U25064 (N_25064,N_19360,N_18440);
or U25065 (N_25065,N_20822,N_21347);
xnor U25066 (N_25066,N_18368,N_22725);
or U25067 (N_25067,N_22383,N_20566);
xnor U25068 (N_25068,N_21054,N_19070);
or U25069 (N_25069,N_21941,N_23702);
xnor U25070 (N_25070,N_23868,N_18956);
xnor U25071 (N_25071,N_20607,N_20809);
or U25072 (N_25072,N_21326,N_20165);
nand U25073 (N_25073,N_23620,N_23071);
nor U25074 (N_25074,N_21309,N_22666);
nor U25075 (N_25075,N_20614,N_21290);
nand U25076 (N_25076,N_23717,N_23130);
xnor U25077 (N_25077,N_23441,N_18503);
nor U25078 (N_25078,N_19904,N_22510);
and U25079 (N_25079,N_22603,N_18225);
nand U25080 (N_25080,N_19150,N_19077);
nand U25081 (N_25081,N_19665,N_23728);
nor U25082 (N_25082,N_19139,N_19204);
nand U25083 (N_25083,N_23188,N_20585);
or U25084 (N_25084,N_21294,N_19151);
nor U25085 (N_25085,N_18245,N_20398);
nand U25086 (N_25086,N_22524,N_19228);
nand U25087 (N_25087,N_21396,N_22898);
or U25088 (N_25088,N_21112,N_21489);
xnor U25089 (N_25089,N_20792,N_23033);
and U25090 (N_25090,N_21106,N_23651);
or U25091 (N_25091,N_18000,N_18514);
nor U25092 (N_25092,N_23735,N_19049);
nor U25093 (N_25093,N_21343,N_23963);
or U25094 (N_25094,N_23250,N_19205);
and U25095 (N_25095,N_18750,N_18534);
or U25096 (N_25096,N_21321,N_19743);
xnor U25097 (N_25097,N_22365,N_19472);
and U25098 (N_25098,N_21539,N_21686);
or U25099 (N_25099,N_20514,N_20966);
nand U25100 (N_25100,N_20369,N_23221);
and U25101 (N_25101,N_19028,N_22513);
and U25102 (N_25102,N_20226,N_20371);
xor U25103 (N_25103,N_22162,N_21613);
xor U25104 (N_25104,N_19356,N_22526);
nor U25105 (N_25105,N_21253,N_19512);
xor U25106 (N_25106,N_23969,N_23580);
nor U25107 (N_25107,N_19556,N_19403);
or U25108 (N_25108,N_18767,N_23379);
or U25109 (N_25109,N_23014,N_20833);
xnor U25110 (N_25110,N_23363,N_18060);
nor U25111 (N_25111,N_18021,N_20483);
xnor U25112 (N_25112,N_19011,N_19628);
xor U25113 (N_25113,N_18625,N_22767);
and U25114 (N_25114,N_21261,N_18492);
nor U25115 (N_25115,N_18323,N_23333);
or U25116 (N_25116,N_20848,N_22092);
xnor U25117 (N_25117,N_21498,N_21151);
xor U25118 (N_25118,N_19313,N_22201);
and U25119 (N_25119,N_18717,N_20136);
and U25120 (N_25120,N_23962,N_22095);
nand U25121 (N_25121,N_21414,N_23152);
or U25122 (N_25122,N_22776,N_19030);
and U25123 (N_25123,N_19116,N_23939);
nor U25124 (N_25124,N_21732,N_19618);
or U25125 (N_25125,N_21600,N_18725);
or U25126 (N_25126,N_21361,N_22116);
xnor U25127 (N_25127,N_21308,N_23059);
xor U25128 (N_25128,N_23121,N_20865);
and U25129 (N_25129,N_23426,N_18768);
nand U25130 (N_25130,N_23999,N_23412);
and U25131 (N_25131,N_21711,N_20570);
nand U25132 (N_25132,N_23063,N_20287);
and U25133 (N_25133,N_22227,N_19845);
nand U25134 (N_25134,N_19895,N_22802);
nand U25135 (N_25135,N_19321,N_20786);
and U25136 (N_25136,N_19027,N_22232);
nand U25137 (N_25137,N_23225,N_18691);
and U25138 (N_25138,N_22240,N_20664);
and U25139 (N_25139,N_22342,N_19479);
nand U25140 (N_25140,N_22507,N_21990);
xnor U25141 (N_25141,N_23952,N_18911);
xor U25142 (N_25142,N_20924,N_23055);
and U25143 (N_25143,N_21506,N_21417);
or U25144 (N_25144,N_18603,N_22661);
or U25145 (N_25145,N_20455,N_19254);
nor U25146 (N_25146,N_18570,N_18012);
xnor U25147 (N_25147,N_20097,N_20028);
nor U25148 (N_25148,N_20602,N_19316);
nor U25149 (N_25149,N_21380,N_19161);
and U25150 (N_25150,N_18538,N_19487);
nand U25151 (N_25151,N_23598,N_21518);
xor U25152 (N_25152,N_22839,N_23648);
nand U25153 (N_25153,N_22377,N_18367);
nor U25154 (N_25154,N_18825,N_18661);
nor U25155 (N_25155,N_20169,N_19224);
and U25156 (N_25156,N_23252,N_20400);
or U25157 (N_25157,N_21126,N_21770);
nand U25158 (N_25158,N_23829,N_22914);
and U25159 (N_25159,N_20328,N_21215);
and U25160 (N_25160,N_18883,N_20595);
nand U25161 (N_25161,N_18202,N_22386);
and U25162 (N_25162,N_23724,N_20765);
nor U25163 (N_25163,N_21520,N_22192);
xnor U25164 (N_25164,N_18097,N_22850);
nand U25165 (N_25165,N_22813,N_20641);
or U25166 (N_25166,N_20208,N_21235);
and U25167 (N_25167,N_21656,N_18748);
and U25168 (N_25168,N_23652,N_22120);
nor U25169 (N_25169,N_22549,N_20869);
xnor U25170 (N_25170,N_21923,N_18252);
nor U25171 (N_25171,N_22965,N_18586);
or U25172 (N_25172,N_22844,N_20984);
xnor U25173 (N_25173,N_19595,N_19386);
and U25174 (N_25174,N_20572,N_21076);
and U25175 (N_25175,N_22274,N_21411);
nor U25176 (N_25176,N_22664,N_21586);
nand U25177 (N_25177,N_22046,N_19507);
xor U25178 (N_25178,N_21702,N_21496);
nand U25179 (N_25179,N_19597,N_19833);
nand U25180 (N_25180,N_18034,N_20979);
or U25181 (N_25181,N_21482,N_22014);
nor U25182 (N_25182,N_23618,N_20655);
or U25183 (N_25183,N_20295,N_23155);
nand U25184 (N_25184,N_23492,N_22711);
nor U25185 (N_25185,N_19898,N_22555);
xor U25186 (N_25186,N_22566,N_19047);
xor U25187 (N_25187,N_18402,N_19725);
nor U25188 (N_25188,N_23257,N_20626);
xor U25189 (N_25189,N_22479,N_19145);
xor U25190 (N_25190,N_18606,N_18359);
and U25191 (N_25191,N_21538,N_19958);
or U25192 (N_25192,N_19155,N_20745);
or U25193 (N_25193,N_22406,N_22645);
and U25194 (N_25194,N_23270,N_22591);
nor U25195 (N_25195,N_22600,N_23778);
xor U25196 (N_25196,N_19832,N_22908);
and U25197 (N_25197,N_18207,N_21728);
nor U25198 (N_25198,N_19073,N_19985);
nor U25199 (N_25199,N_23559,N_20603);
or U25200 (N_25200,N_18777,N_23666);
xor U25201 (N_25201,N_23824,N_22704);
nand U25202 (N_25202,N_20956,N_23078);
or U25203 (N_25203,N_21022,N_18828);
nand U25204 (N_25204,N_19088,N_20642);
and U25205 (N_25205,N_22332,N_20269);
nand U25206 (N_25206,N_19799,N_20821);
xnor U25207 (N_25207,N_23606,N_20027);
xor U25208 (N_25208,N_18014,N_23139);
xnor U25209 (N_25209,N_18089,N_22885);
and U25210 (N_25210,N_18928,N_22729);
and U25211 (N_25211,N_21753,N_18839);
and U25212 (N_25212,N_18520,N_18112);
and U25213 (N_25213,N_21091,N_21262);
nor U25214 (N_25214,N_19429,N_20593);
nand U25215 (N_25215,N_21933,N_21605);
nand U25216 (N_25216,N_20122,N_23030);
nor U25217 (N_25217,N_20841,N_19232);
or U25218 (N_25218,N_18456,N_19181);
and U25219 (N_25219,N_22631,N_22720);
and U25220 (N_25220,N_22330,N_20991);
and U25221 (N_25221,N_20236,N_22579);
and U25222 (N_25222,N_18376,N_22927);
nand U25223 (N_25223,N_23313,N_21252);
or U25224 (N_25224,N_21909,N_21031);
and U25225 (N_25225,N_19107,N_20288);
nand U25226 (N_25226,N_21368,N_19079);
nand U25227 (N_25227,N_18441,N_21743);
and U25228 (N_25228,N_18105,N_23183);
nand U25229 (N_25229,N_21021,N_19741);
nor U25230 (N_25230,N_22540,N_20938);
xnor U25231 (N_25231,N_20702,N_18124);
nand U25232 (N_25232,N_19999,N_20969);
or U25233 (N_25233,N_23650,N_18162);
nand U25234 (N_25234,N_18129,N_19110);
and U25235 (N_25235,N_22159,N_22906);
or U25236 (N_25236,N_22521,N_18073);
or U25237 (N_25237,N_22809,N_22628);
and U25238 (N_25238,N_18728,N_23227);
and U25239 (N_25239,N_20281,N_18114);
xor U25240 (N_25240,N_21255,N_21461);
or U25241 (N_25241,N_19727,N_20002);
nor U25242 (N_25242,N_19179,N_23705);
or U25243 (N_25243,N_23869,N_23740);
nor U25244 (N_25244,N_22501,N_21650);
xor U25245 (N_25245,N_21925,N_22324);
nand U25246 (N_25246,N_18798,N_19440);
or U25247 (N_25247,N_18064,N_22135);
xor U25248 (N_25248,N_20506,N_21558);
and U25249 (N_25249,N_19874,N_22304);
xor U25250 (N_25250,N_23015,N_23075);
or U25251 (N_25251,N_22437,N_21082);
nand U25252 (N_25252,N_22865,N_19177);
or U25253 (N_25253,N_22271,N_20559);
or U25254 (N_25254,N_18700,N_20324);
xnor U25255 (N_25255,N_22263,N_23710);
nor U25256 (N_25256,N_23438,N_18241);
nand U25257 (N_25257,N_20210,N_19128);
and U25258 (N_25258,N_18929,N_23837);
or U25259 (N_25259,N_19819,N_22335);
xnor U25260 (N_25260,N_20544,N_22170);
and U25261 (N_25261,N_21982,N_22500);
and U25262 (N_25262,N_22173,N_19566);
nand U25263 (N_25263,N_20951,N_22251);
nand U25264 (N_25264,N_18346,N_22237);
nor U25265 (N_25265,N_20574,N_20125);
or U25266 (N_25266,N_21701,N_22090);
and U25267 (N_25267,N_21763,N_22356);
or U25268 (N_25268,N_19267,N_22534);
xor U25269 (N_25269,N_20127,N_20152);
and U25270 (N_25270,N_20766,N_23823);
or U25271 (N_25271,N_23023,N_18811);
or U25272 (N_25272,N_22673,N_23772);
nor U25273 (N_25273,N_21754,N_20298);
nor U25274 (N_25274,N_20795,N_22398);
and U25275 (N_25275,N_20187,N_20921);
xnor U25276 (N_25276,N_20801,N_21014);
and U25277 (N_25277,N_23528,N_18688);
xnor U25278 (N_25278,N_21849,N_19148);
xor U25279 (N_25279,N_21176,N_21733);
xor U25280 (N_25280,N_23553,N_21638);
or U25281 (N_25281,N_23500,N_20256);
xnor U25282 (N_25282,N_23936,N_21508);
or U25283 (N_25283,N_20271,N_18358);
and U25284 (N_25284,N_20384,N_21999);
xor U25285 (N_25285,N_22373,N_19978);
or U25286 (N_25286,N_20719,N_23647);
and U25287 (N_25287,N_22612,N_22975);
nand U25288 (N_25288,N_23342,N_20820);
or U25289 (N_25289,N_21516,N_21841);
or U25290 (N_25290,N_19129,N_18707);
or U25291 (N_25291,N_23264,N_20689);
xor U25292 (N_25292,N_21295,N_18465);
and U25293 (N_25293,N_20700,N_20278);
nor U25294 (N_25294,N_22849,N_19042);
nand U25295 (N_25295,N_22583,N_21310);
and U25296 (N_25296,N_23065,N_22163);
or U25297 (N_25297,N_18916,N_19576);
nand U25298 (N_25298,N_21407,N_22205);
or U25299 (N_25299,N_18871,N_19581);
xnor U25300 (N_25300,N_23689,N_20174);
nand U25301 (N_25301,N_18508,N_23827);
or U25302 (N_25302,N_23177,N_18670);
xnor U25303 (N_25303,N_19138,N_19255);
nand U25304 (N_25304,N_22608,N_21833);
nand U25305 (N_25305,N_22496,N_18354);
nor U25306 (N_25306,N_18736,N_19172);
xor U25307 (N_25307,N_20354,N_21030);
nand U25308 (N_25308,N_22837,N_23656);
xor U25309 (N_25309,N_23297,N_22982);
xnor U25310 (N_25310,N_21395,N_22924);
xnor U25311 (N_25311,N_21655,N_23079);
xor U25312 (N_25312,N_22747,N_22005);
and U25313 (N_25313,N_18013,N_21288);
or U25314 (N_25314,N_19957,N_22230);
xor U25315 (N_25315,N_23068,N_20720);
nand U25316 (N_25316,N_18299,N_19471);
xor U25317 (N_25317,N_19888,N_18559);
or U25318 (N_25318,N_20444,N_22539);
xnor U25319 (N_25319,N_18959,N_21051);
xor U25320 (N_25320,N_18719,N_22016);
nand U25321 (N_25321,N_23865,N_19283);
or U25322 (N_25322,N_19419,N_23249);
xor U25323 (N_25323,N_20516,N_21685);
and U25324 (N_25324,N_19890,N_22471);
nand U25325 (N_25325,N_20238,N_21589);
nor U25326 (N_25326,N_21988,N_22905);
xor U25327 (N_25327,N_20489,N_18953);
xnor U25328 (N_25328,N_22026,N_23552);
or U25329 (N_25329,N_18542,N_23311);
nor U25330 (N_25330,N_21907,N_20739);
or U25331 (N_25331,N_20156,N_21657);
or U25332 (N_25332,N_22614,N_18714);
xor U25333 (N_25333,N_19520,N_18948);
xor U25334 (N_25334,N_21228,N_23957);
nand U25335 (N_25335,N_20706,N_18125);
nand U25336 (N_25336,N_19728,N_18887);
or U25337 (N_25337,N_22322,N_23690);
or U25338 (N_25338,N_19348,N_20836);
xnor U25339 (N_25339,N_21092,N_19207);
xnor U25340 (N_25340,N_18500,N_23229);
nor U25341 (N_25341,N_20421,N_21793);
nor U25342 (N_25342,N_18610,N_19167);
or U25343 (N_25343,N_21706,N_19603);
or U25344 (N_25344,N_18275,N_22483);
nand U25345 (N_25345,N_23902,N_22050);
and U25346 (N_25346,N_18110,N_20033);
nand U25347 (N_25347,N_20691,N_21177);
xor U25348 (N_25348,N_19413,N_22419);
nand U25349 (N_25349,N_22004,N_21425);
nor U25350 (N_25350,N_22899,N_18848);
xnor U25351 (N_25351,N_23047,N_19013);
nor U25352 (N_25352,N_22070,N_21244);
xor U25353 (N_25353,N_19906,N_20157);
and U25354 (N_25354,N_23816,N_18058);
or U25355 (N_25355,N_19192,N_22739);
nand U25356 (N_25356,N_21383,N_20153);
or U25357 (N_25357,N_18256,N_23562);
nand U25358 (N_25358,N_23132,N_18100);
and U25359 (N_25359,N_23516,N_21117);
nor U25360 (N_25360,N_19588,N_18228);
or U25361 (N_25361,N_20696,N_19022);
and U25362 (N_25362,N_19676,N_18011);
nand U25363 (N_25363,N_22188,N_20089);
and U25364 (N_25364,N_18622,N_20464);
and U25365 (N_25365,N_20529,N_20972);
xnor U25366 (N_25366,N_20030,N_19199);
xor U25367 (N_25367,N_23574,N_22764);
nand U25368 (N_25368,N_22606,N_23165);
or U25369 (N_25369,N_23594,N_23883);
xor U25370 (N_25370,N_21748,N_22551);
nor U25371 (N_25371,N_20829,N_18510);
and U25372 (N_25372,N_21804,N_23397);
nand U25373 (N_25373,N_22233,N_23429);
nand U25374 (N_25374,N_21889,N_21327);
and U25375 (N_25375,N_18875,N_18119);
xor U25376 (N_25376,N_22822,N_20106);
nor U25377 (N_25377,N_18664,N_18523);
nor U25378 (N_25378,N_21466,N_20394);
and U25379 (N_25379,N_20775,N_20998);
nand U25380 (N_25380,N_18895,N_23122);
xnor U25381 (N_25381,N_21715,N_19737);
nand U25382 (N_25382,N_18618,N_21316);
xnor U25383 (N_25383,N_18247,N_22317);
nor U25384 (N_25384,N_20268,N_21771);
nand U25385 (N_25385,N_19546,N_21612);
nand U25386 (N_25386,N_18794,N_22872);
nor U25387 (N_25387,N_19683,N_18115);
nand U25388 (N_25388,N_20143,N_23389);
and U25389 (N_25389,N_21777,N_19398);
and U25390 (N_25390,N_19014,N_18094);
and U25391 (N_25391,N_18524,N_21906);
xor U25392 (N_25392,N_23185,N_21615);
or U25393 (N_25393,N_21330,N_19481);
and U25394 (N_25394,N_20397,N_23544);
xnor U25395 (N_25395,N_23261,N_18528);
or U25396 (N_25396,N_22773,N_19165);
nand U25397 (N_25397,N_20948,N_22833);
nand U25398 (N_25398,N_19438,N_19616);
xor U25399 (N_25399,N_18331,N_23916);
and U25400 (N_25400,N_20501,N_18676);
and U25401 (N_25401,N_21902,N_18254);
nor U25402 (N_25402,N_21760,N_22075);
and U25403 (N_25403,N_18293,N_19590);
nand U25404 (N_25404,N_20300,N_18834);
and U25405 (N_25405,N_18163,N_19600);
or U25406 (N_25406,N_22057,N_23791);
xnor U25407 (N_25407,N_22860,N_19885);
xor U25408 (N_25408,N_18898,N_21817);
nand U25409 (N_25409,N_21731,N_21823);
nor U25410 (N_25410,N_20182,N_23294);
xor U25411 (N_25411,N_21927,N_23374);
nand U25412 (N_25412,N_18071,N_22962);
nor U25413 (N_25413,N_21283,N_22366);
or U25414 (N_25414,N_22038,N_19797);
xnor U25415 (N_25415,N_21147,N_18619);
and U25416 (N_25416,N_23440,N_20826);
and U25417 (N_25417,N_23231,N_20580);
nand U25418 (N_25418,N_20219,N_21345);
xor U25419 (N_25419,N_23289,N_21185);
nor U25420 (N_25420,N_19667,N_22613);
xnor U25421 (N_25421,N_22861,N_22803);
nand U25422 (N_25422,N_20768,N_19666);
nor U25423 (N_25423,N_18068,N_23160);
or U25424 (N_25424,N_22359,N_22650);
or U25425 (N_25425,N_19211,N_21646);
or U25426 (N_25426,N_20783,N_22093);
nand U25427 (N_25427,N_22867,N_23783);
or U25428 (N_25428,N_18738,N_22854);
nand U25429 (N_25429,N_22624,N_23638);
nand U25430 (N_25430,N_18480,N_22029);
xor U25431 (N_25431,N_21819,N_22556);
or U25432 (N_25432,N_21540,N_23775);
nand U25433 (N_25433,N_21007,N_23736);
nand U25434 (N_25434,N_23750,N_22544);
nor U25435 (N_25435,N_21390,N_21810);
nor U25436 (N_25436,N_21710,N_23453);
nor U25437 (N_25437,N_23509,N_19771);
and U25438 (N_25438,N_23903,N_20732);
and U25439 (N_25439,N_23501,N_19601);
xnor U25440 (N_25440,N_18967,N_20481);
or U25441 (N_25441,N_18601,N_23715);
nor U25442 (N_25442,N_23143,N_18337);
and U25443 (N_25443,N_21236,N_18276);
or U25444 (N_25444,N_21635,N_18419);
nand U25445 (N_25445,N_22532,N_22499);
and U25446 (N_25446,N_22033,N_18059);
xor U25447 (N_25447,N_22293,N_23387);
or U25448 (N_25448,N_23356,N_20335);
and U25449 (N_25449,N_18716,N_18940);
nand U25450 (N_25450,N_21879,N_19847);
or U25451 (N_25451,N_19761,N_23331);
or U25452 (N_25452,N_19557,N_21240);
and U25453 (N_25453,N_23460,N_19974);
xnor U25454 (N_25454,N_18914,N_21956);
or U25455 (N_25455,N_21083,N_21277);
nand U25456 (N_25456,N_23133,N_20985);
and U25457 (N_25457,N_21105,N_22538);
nand U25458 (N_25458,N_18494,N_23535);
xor U25459 (N_25459,N_21886,N_20085);
nor U25460 (N_25460,N_22007,N_18239);
and U25461 (N_25461,N_19684,N_21581);
nand U25462 (N_25462,N_18236,N_18997);
xnor U25463 (N_25463,N_21830,N_18266);
and U25464 (N_25464,N_21687,N_19350);
or U25465 (N_25465,N_21768,N_20834);
nand U25466 (N_25466,N_18411,N_18195);
nor U25467 (N_25467,N_22786,N_23893);
nor U25468 (N_25468,N_19242,N_21785);
xor U25469 (N_25469,N_23476,N_23576);
or U25470 (N_25470,N_18473,N_21292);
xor U25471 (N_25471,N_22542,N_23216);
nand U25472 (N_25472,N_21120,N_22413);
nand U25473 (N_25473,N_18345,N_22180);
xnor U25474 (N_25474,N_23392,N_23671);
nor U25475 (N_25475,N_18027,N_19960);
or U25476 (N_25476,N_20562,N_23019);
nand U25477 (N_25477,N_20475,N_23182);
nand U25478 (N_25478,N_18556,N_19580);
nand U25479 (N_25479,N_19040,N_22695);
and U25480 (N_25480,N_18384,N_22054);
or U25481 (N_25481,N_20452,N_23110);
xnor U25482 (N_25482,N_19726,N_22143);
xnor U25483 (N_25483,N_21712,N_18978);
and U25484 (N_25484,N_23038,N_18131);
xnor U25485 (N_25485,N_22721,N_23411);
nor U25486 (N_25486,N_18109,N_20653);
and U25487 (N_25487,N_22836,N_19131);
nand U25488 (N_25488,N_21698,N_22868);
xnor U25489 (N_25489,N_20310,N_20083);
nor U25490 (N_25490,N_19220,N_21842);
nand U25491 (N_25491,N_19963,N_23147);
or U25492 (N_25492,N_23027,N_22068);
or U25493 (N_25493,N_22769,N_22074);
or U25494 (N_25494,N_20206,N_21863);
nand U25495 (N_25495,N_19498,N_21971);
and U25496 (N_25496,N_18336,N_20181);
or U25497 (N_25497,N_18158,N_23260);
or U25498 (N_25498,N_18078,N_19483);
and U25499 (N_25499,N_20061,N_22724);
xnor U25500 (N_25500,N_21025,N_20999);
nor U25501 (N_25501,N_18138,N_21282);
or U25502 (N_25502,N_21088,N_22221);
nor U25503 (N_25503,N_20594,N_22308);
nor U25504 (N_25504,N_18461,N_20472);
nand U25505 (N_25505,N_19300,N_18235);
nor U25506 (N_25506,N_23102,N_23032);
xnor U25507 (N_25507,N_21314,N_23987);
nand U25508 (N_25508,N_20815,N_21162);
xnor U25509 (N_25509,N_21296,N_18382);
nand U25510 (N_25510,N_18902,N_19423);
nor U25511 (N_25511,N_18535,N_21384);
nand U25512 (N_25512,N_19828,N_18355);
or U25513 (N_25513,N_19016,N_22580);
and U25514 (N_25514,N_20751,N_21372);
and U25515 (N_25515,N_18984,N_20001);
nor U25516 (N_25516,N_21453,N_19395);
nor U25517 (N_25517,N_18135,N_22429);
nor U25518 (N_25518,N_18398,N_22541);
nor U25519 (N_25519,N_19289,N_23338);
or U25520 (N_25520,N_19912,N_18891);
or U25521 (N_25521,N_19341,N_23644);
and U25522 (N_25522,N_21884,N_21387);
xor U25523 (N_25523,N_21669,N_19373);
and U25524 (N_25524,N_21848,N_18754);
and U25525 (N_25525,N_21207,N_21222);
nand U25526 (N_25526,N_23118,N_18003);
and U25527 (N_25527,N_20774,N_21490);
nor U25528 (N_25528,N_21703,N_18853);
nand U25529 (N_25529,N_19256,N_18404);
xnor U25530 (N_25530,N_22283,N_18406);
xnor U25531 (N_25531,N_18576,N_23507);
and U25532 (N_25532,N_18675,N_18184);
nand U25533 (N_25533,N_18351,N_21965);
nor U25534 (N_25534,N_19000,N_18342);
or U25535 (N_25535,N_20383,N_21658);
nand U25536 (N_25536,N_23268,N_20032);
nand U25537 (N_25537,N_22957,N_23370);
and U25538 (N_25538,N_20573,N_20541);
nand U25539 (N_25539,N_19391,N_20524);
and U25540 (N_25540,N_18597,N_19916);
and U25541 (N_25541,N_20046,N_22748);
nor U25542 (N_25542,N_21324,N_22679);
and U25543 (N_25543,N_21418,N_22089);
or U25544 (N_25544,N_18314,N_20531);
nor U25545 (N_25545,N_18133,N_18209);
nor U25546 (N_25546,N_18992,N_22013);
or U25547 (N_25547,N_22469,N_20962);
and U25548 (N_25548,N_21964,N_22081);
nand U25549 (N_25549,N_20873,N_21339);
xor U25550 (N_25550,N_19768,N_23794);
and U25551 (N_25551,N_22397,N_21075);
xor U25552 (N_25552,N_20644,N_18521);
nand U25553 (N_25553,N_21435,N_19132);
or U25554 (N_25554,N_21412,N_22411);
nand U25555 (N_25555,N_19501,N_22234);
nor U25556 (N_25556,N_19987,N_18243);
and U25557 (N_25557,N_22866,N_19359);
nand U25558 (N_25558,N_19705,N_22462);
nand U25559 (N_25559,N_23228,N_18144);
and U25560 (N_25560,N_18681,N_20533);
nand U25561 (N_25561,N_19872,N_23259);
nor U25562 (N_25562,N_19822,N_23043);
nand U25563 (N_25563,N_19816,N_21089);
and U25564 (N_25564,N_20704,N_23317);
nor U25565 (N_25565,N_21263,N_21745);
or U25566 (N_25566,N_23919,N_23357);
xor U25567 (N_25567,N_21836,N_19057);
nand U25568 (N_25568,N_21727,N_22222);
nor U25569 (N_25569,N_22601,N_21921);
nor U25570 (N_25570,N_23349,N_21621);
and U25571 (N_25571,N_21409,N_21940);
nor U25572 (N_25572,N_19500,N_18009);
and U25573 (N_25573,N_18308,N_22374);
and U25574 (N_25574,N_23933,N_18659);
xnor U25575 (N_25575,N_21341,N_21557);
xnor U25576 (N_25576,N_19521,N_18408);
nor U25577 (N_25577,N_23760,N_18268);
or U25578 (N_25578,N_20609,N_19465);
xnor U25579 (N_25579,N_21163,N_18561);
xor U25580 (N_25580,N_23613,N_21627);
and U25581 (N_25581,N_23436,N_19272);
or U25582 (N_25582,N_21828,N_20321);
or U25583 (N_25583,N_21026,N_18385);
or U25584 (N_25584,N_19854,N_18146);
nor U25585 (N_25585,N_23674,N_23599);
xor U25586 (N_25586,N_22782,N_22039);
nor U25587 (N_25587,N_21825,N_18328);
or U25588 (N_25588,N_18554,N_21654);
nor U25589 (N_25589,N_18483,N_23793);
nand U25590 (N_25590,N_18966,N_23005);
xor U25591 (N_25591,N_19103,N_23134);
nor U25592 (N_25592,N_19482,N_20063);
and U25593 (N_25593,N_22588,N_20166);
and U25594 (N_25594,N_19711,N_19892);
or U25595 (N_25595,N_19767,N_19149);
and U25596 (N_25596,N_22460,N_21576);
and U25597 (N_25597,N_21677,N_20360);
and U25598 (N_25598,N_18491,N_23365);
or U25599 (N_25599,N_20308,N_22108);
nand U25600 (N_25600,N_18199,N_22477);
and U25601 (N_25601,N_21691,N_23362);
and U25602 (N_25602,N_19173,N_19511);
nand U25603 (N_25603,N_20184,N_21664);
nand U25604 (N_25604,N_18820,N_19406);
nand U25605 (N_25605,N_18772,N_19108);
and U25606 (N_25606,N_18270,N_19469);
nand U25607 (N_25607,N_21900,N_22758);
nand U25608 (N_25608,N_23400,N_21101);
nand U25609 (N_25609,N_19802,N_18242);
and U25610 (N_25610,N_20845,N_21429);
nor U25611 (N_25611,N_21741,N_19721);
and U25612 (N_25612,N_19865,N_22333);
or U25613 (N_25613,N_22493,N_23163);
and U25614 (N_25614,N_22053,N_22280);
xnor U25615 (N_25615,N_18734,N_23811);
or U25616 (N_25616,N_21444,N_19491);
or U25617 (N_25617,N_21491,N_23488);
and U25618 (N_25618,N_18445,N_21402);
xor U25619 (N_25619,N_23494,N_18686);
nand U25620 (N_25620,N_23726,N_20828);
nor U25621 (N_25621,N_23532,N_18819);
nor U25622 (N_25622,N_20980,N_20362);
nand U25623 (N_25623,N_20846,N_21208);
and U25624 (N_25624,N_19130,N_23533);
and U25625 (N_25625,N_19393,N_20255);
xor U25626 (N_25626,N_22857,N_20284);
nor U25627 (N_25627,N_20847,N_21799);
and U25628 (N_25628,N_21251,N_22449);
and U25629 (N_25629,N_19006,N_18436);
nand U25630 (N_25630,N_20534,N_20374);
or U25631 (N_25631,N_21128,N_22349);
or U25632 (N_25632,N_20110,N_18056);
nand U25633 (N_25633,N_22202,N_22147);
and U25634 (N_25634,N_22125,N_22216);
nand U25635 (N_25635,N_18025,N_19063);
nand U25636 (N_25636,N_23604,N_19813);
nor U25637 (N_25637,N_19878,N_18602);
nand U25638 (N_25638,N_22939,N_22208);
or U25639 (N_25639,N_22869,N_20015);
nand U25640 (N_25640,N_21813,N_20438);
xor U25641 (N_25641,N_19410,N_20018);
nand U25642 (N_25642,N_18566,N_18103);
xnor U25643 (N_25643,N_18053,N_23093);
nand U25644 (N_25644,N_22506,N_23003);
or U25645 (N_25645,N_22618,N_18046);
nor U25646 (N_25646,N_18361,N_21660);
nor U25647 (N_25647,N_22728,N_21858);
xor U25648 (N_25648,N_19433,N_20409);
or U25649 (N_25649,N_22625,N_23291);
or U25650 (N_25650,N_20056,N_19716);
and U25651 (N_25651,N_22827,N_22722);
xnor U25652 (N_25652,N_20198,N_20448);
nor U25653 (N_25653,N_23149,N_20479);
nor U25654 (N_25654,N_22959,N_19265);
and U25655 (N_25655,N_20525,N_21027);
and U25656 (N_25656,N_22796,N_23421);
or U25657 (N_25657,N_20407,N_22688);
or U25658 (N_25658,N_23306,N_21803);
or U25659 (N_25659,N_21473,N_21109);
nand U25660 (N_25660,N_21895,N_19189);
or U25661 (N_25661,N_21424,N_21765);
or U25662 (N_25662,N_19824,N_21758);
xor U25663 (N_25663,N_22863,N_20554);
nand U25664 (N_25664,N_20710,N_20854);
nor U25665 (N_25665,N_22937,N_18123);
and U25666 (N_25666,N_23167,N_19788);
or U25667 (N_25667,N_23128,N_21386);
xor U25668 (N_25668,N_21913,N_23578);
nand U25669 (N_25669,N_20134,N_21532);
nand U25670 (N_25670,N_18035,N_21137);
nand U25671 (N_25671,N_18050,N_23605);
or U25672 (N_25672,N_20265,N_23153);
nand U25673 (N_25673,N_22119,N_23069);
nand U25674 (N_25674,N_22415,N_19295);
nor U25675 (N_25675,N_20782,N_23543);
and U25676 (N_25676,N_22291,N_19508);
or U25677 (N_25677,N_18872,N_21816);
xor U25678 (N_25678,N_21578,N_23534);
nor U25679 (N_25679,N_18347,N_21306);
or U25680 (N_25680,N_22785,N_21258);
or U25681 (N_25681,N_18444,N_22168);
or U25682 (N_25682,N_22123,N_22670);
nor U25683 (N_25683,N_23238,N_19900);
nand U25684 (N_25684,N_22752,N_23978);
and U25685 (N_25685,N_21822,N_21049);
xor U25686 (N_25686,N_22187,N_23833);
nor U25687 (N_25687,N_19383,N_18099);
and U25688 (N_25688,N_21559,N_22444);
nor U25689 (N_25689,N_20000,N_22408);
nand U25690 (N_25690,N_20662,N_23292);
xnor U25691 (N_25691,N_20164,N_19381);
nand U25692 (N_25692,N_23326,N_21675);
and U25693 (N_25693,N_19657,N_19260);
nor U25694 (N_25694,N_19454,N_20988);
xor U25695 (N_25695,N_18517,N_20857);
nor U25696 (N_25696,N_18945,N_19887);
xnor U25697 (N_25697,N_22099,N_18584);
nand U25698 (N_25698,N_22853,N_19550);
nor U25699 (N_25699,N_20386,N_20571);
and U25700 (N_25700,N_23286,N_19886);
xor U25701 (N_25701,N_22743,N_18277);
nand U25702 (N_25702,N_18855,N_20891);
nor U25703 (N_25703,N_19473,N_23759);
and U25704 (N_25704,N_18906,N_21782);
xor U25705 (N_25705,N_18611,N_23323);
nor U25706 (N_25706,N_19636,N_18642);
nor U25707 (N_25707,N_23720,N_23655);
or U25708 (N_25708,N_20410,N_22442);
and U25709 (N_25709,N_23584,N_19208);
nand U25710 (N_25710,N_18428,N_19627);
xnor U25711 (N_25711,N_23954,N_22314);
or U25712 (N_25712,N_21625,N_23990);
xnor U25713 (N_25713,N_21966,N_22140);
nand U25714 (N_25714,N_21212,N_23624);
or U25715 (N_25715,N_18435,N_21501);
nand U25716 (N_25716,N_23975,N_21085);
nand U25717 (N_25717,N_19095,N_22979);
nor U25718 (N_25718,N_23148,N_21281);
nand U25719 (N_25719,N_21939,N_20656);
or U25720 (N_25720,N_20830,N_20671);
nor U25721 (N_25721,N_23561,N_23499);
or U25722 (N_25722,N_23007,N_23067);
nand U25723 (N_25723,N_21102,N_22410);
nand U25724 (N_25724,N_19680,N_21289);
nand U25725 (N_25725,N_21542,N_19661);
and U25726 (N_25726,N_23491,N_23360);
xor U25727 (N_25727,N_22423,N_20920);
xor U25728 (N_25728,N_18518,N_22487);
and U25729 (N_25729,N_22124,N_22677);
nand U25730 (N_25730,N_23887,N_21073);
nand U25731 (N_25731,N_22196,N_23828);
nand U25732 (N_25732,N_20413,N_20192);
nand U25733 (N_25733,N_19746,N_18838);
nor U25734 (N_25734,N_21381,N_18063);
or U25735 (N_25735,N_23170,N_20241);
nor U25736 (N_25736,N_19085,N_19367);
or U25737 (N_25737,N_18983,N_18660);
xnor U25738 (N_25738,N_20330,N_20078);
xor U25739 (N_25739,N_20912,N_22637);
xnor U25740 (N_25740,N_22990,N_23888);
and U25741 (N_25741,N_22731,N_23608);
and U25742 (N_25742,N_18987,N_23407);
or U25743 (N_25743,N_20565,N_20487);
nor U25744 (N_25744,N_22294,N_21492);
xnor U25745 (N_25745,N_23089,N_18420);
nor U25746 (N_25746,N_18961,N_18787);
xnor U25747 (N_25747,N_18365,N_18305);
nor U25748 (N_25748,N_18858,N_18432);
or U25749 (N_25749,N_19154,N_20365);
xnor U25750 (N_25750,N_23470,N_19903);
or U25751 (N_25751,N_23838,N_18143);
nand U25752 (N_25752,N_21876,N_23641);
or U25753 (N_25753,N_23976,N_19821);
xnor U25754 (N_25754,N_20424,N_21286);
nand U25755 (N_25755,N_21064,N_22550);
nor U25756 (N_25756,N_18426,N_23432);
nand U25757 (N_25757,N_22834,N_21766);
xor U25758 (N_25758,N_20332,N_21220);
xnor U25759 (N_25759,N_18815,N_20504);
nor U25760 (N_25760,N_19044,N_22690);
or U25761 (N_25761,N_21624,N_21188);
nor U25762 (N_25762,N_21287,N_19050);
nor U25763 (N_25763,N_21260,N_19651);
xnor U25764 (N_25764,N_22684,N_18623);
xnor U25765 (N_25765,N_19640,N_19276);
or U25766 (N_25766,N_23727,N_19412);
nand U25767 (N_25767,N_18737,N_19377);
xnor U25768 (N_25768,N_22707,N_23687);
xnor U25769 (N_25769,N_19733,N_19929);
or U25770 (N_25770,N_19879,N_23378);
xor U25771 (N_25771,N_22288,N_20880);
nand U25772 (N_25772,N_18847,N_20377);
nand U25773 (N_25773,N_22051,N_18905);
nor U25774 (N_25774,N_20297,N_18319);
nand U25775 (N_25775,N_19940,N_23972);
or U25776 (N_25776,N_20797,N_20714);
nand U25777 (N_25777,N_22212,N_19385);
or U25778 (N_25778,N_22515,N_23622);
xor U25779 (N_25779,N_22787,N_18248);
nor U25780 (N_25780,N_22446,N_21096);
nor U25781 (N_25781,N_21989,N_18704);
xor U25782 (N_25782,N_21800,N_21403);
and U25783 (N_25783,N_18102,N_18232);
xor U25784 (N_25784,N_21633,N_22456);
or U25785 (N_25785,N_19795,N_23026);
xnor U25786 (N_25786,N_21892,N_21133);
or U25787 (N_25787,N_19332,N_20497);
xor U25788 (N_25788,N_20249,N_22642);
xnor U25789 (N_25789,N_18450,N_23422);
nand U25790 (N_25790,N_23600,N_19311);
nor U25791 (N_25791,N_22273,N_20610);
and U25792 (N_25792,N_23743,N_19284);
or U25793 (N_25793,N_22385,N_22749);
nand U25794 (N_25794,N_21122,N_21135);
xnor U25795 (N_25795,N_19864,N_19196);
and U25796 (N_25796,N_22973,N_20933);
nand U25797 (N_25797,N_21399,N_21479);
nand U25798 (N_25798,N_19457,N_22733);
nand U25799 (N_25799,N_19182,N_22080);
nor U25800 (N_25800,N_18221,N_23845);
nor U25801 (N_25801,N_21204,N_21707);
xnor U25802 (N_25802,N_18957,N_22559);
nand U25803 (N_25803,N_18952,N_23511);
nand U25804 (N_25804,N_23502,N_19488);
nand U25805 (N_25805,N_22015,N_23186);
nand U25806 (N_25806,N_18587,N_23704);
nor U25807 (N_25807,N_20943,N_19757);
or U25808 (N_25808,N_21280,N_20677);
xor U25809 (N_25809,N_18223,N_18516);
and U25810 (N_25810,N_22244,N_19652);
nand U25811 (N_25811,N_21997,N_21455);
or U25812 (N_25812,N_21720,N_18474);
or U25813 (N_25813,N_21761,N_18401);
or U25814 (N_25814,N_19397,N_20884);
and U25815 (N_25815,N_18998,N_19409);
nor U25816 (N_25816,N_21547,N_20587);
nand U25817 (N_25817,N_19717,N_19645);
or U25818 (N_25818,N_21097,N_18684);
and U25819 (N_25819,N_18278,N_18298);
or U25820 (N_25820,N_22961,N_21433);
nand U25821 (N_25821,N_21269,N_22726);
and U25822 (N_25822,N_20178,N_19713);
and U25823 (N_25823,N_23809,N_19997);
nor U25824 (N_25824,N_23452,N_19850);
and U25825 (N_25825,N_21596,N_19188);
xnor U25826 (N_25826,N_22946,N_20716);
xnor U25827 (N_25827,N_21299,N_21684);
or U25828 (N_25828,N_22789,N_21352);
nor U25829 (N_25829,N_18703,N_23443);
nor U25830 (N_25830,N_20911,N_19017);
and U25831 (N_25831,N_21305,N_22044);
and U25832 (N_25832,N_22467,N_18069);
nand U25833 (N_25833,N_22977,N_20659);
or U25834 (N_25834,N_18090,N_21986);
or U25835 (N_25835,N_22371,N_23593);
or U25836 (N_25836,N_23350,N_18564);
or U25837 (N_25837,N_21639,N_19496);
or U25838 (N_25838,N_19238,N_19451);
nand U25839 (N_25839,N_22911,N_22994);
nor U25840 (N_25840,N_20613,N_19076);
or U25841 (N_25841,N_18047,N_18188);
nand U25842 (N_25842,N_22443,N_22242);
and U25843 (N_25843,N_23495,N_19800);
or U25844 (N_25844,N_20989,N_19375);
and U25845 (N_25845,N_23873,N_18392);
xor U25846 (N_25846,N_19455,N_18451);
and U25847 (N_25847,N_20701,N_21599);
or U25848 (N_25848,N_18540,N_20248);
xnor U25849 (N_25849,N_18613,N_22718);
and U25850 (N_25850,N_21099,N_22931);
xor U25851 (N_25851,N_20856,N_23045);
or U25852 (N_25852,N_22582,N_23857);
xor U25853 (N_25853,N_21821,N_23187);
and U25854 (N_25854,N_22902,N_19288);
nor U25855 (N_25855,N_22999,N_21718);
nor U25856 (N_25856,N_20160,N_20118);
or U25857 (N_25857,N_23369,N_23590);
or U25858 (N_25858,N_23635,N_19421);
nand U25859 (N_25859,N_20895,N_18396);
xnor U25860 (N_25860,N_23858,N_19415);
and U25861 (N_25861,N_23796,N_22409);
nor U25862 (N_25862,N_18558,N_23320);
or U25863 (N_25863,N_21442,N_19437);
nand U25864 (N_25864,N_22571,N_18756);
and U25865 (N_25865,N_20579,N_20355);
xor U25866 (N_25866,N_23285,N_18032);
nor U25867 (N_25867,N_18936,N_21197);
xor U25868 (N_25868,N_22396,N_19745);
xor U25869 (N_25869,N_19135,N_18904);
or U25870 (N_25870,N_23769,N_20676);
or U25871 (N_25871,N_19158,N_18214);
or U25872 (N_25872,N_19634,N_23091);
nand U25873 (N_25873,N_20681,N_20651);
xnor U25874 (N_25874,N_19159,N_23993);
and U25875 (N_25875,N_19849,N_19829);
xnor U25876 (N_25876,N_18780,N_22320);
or U25877 (N_25877,N_22828,N_22393);
xor U25878 (N_25878,N_18732,N_22177);
or U25879 (N_25879,N_22269,N_19416);
nor U25880 (N_25880,N_22372,N_18869);
and U25881 (N_25881,N_20139,N_22648);
nor U25882 (N_25882,N_23766,N_19681);
nand U25883 (N_25883,N_22829,N_20620);
and U25884 (N_25884,N_23377,N_18790);
and U25885 (N_25885,N_22589,N_23210);
or U25886 (N_25886,N_23631,N_22400);
nor U25887 (N_25887,N_22141,N_23049);
nor U25888 (N_25888,N_20342,N_23889);
or U25889 (N_25889,N_18246,N_22451);
xor U25890 (N_25890,N_20250,N_21006);
and U25891 (N_25891,N_23947,N_20280);
nand U25892 (N_25892,N_20222,N_20510);
xnor U25893 (N_25893,N_22951,N_22907);
and U25894 (N_25894,N_23066,N_18751);
xnor U25895 (N_25895,N_19653,N_21095);
or U25896 (N_25896,N_18745,N_22002);
nor U25897 (N_25897,N_19736,N_19448);
nand U25898 (N_25898,N_20742,N_23309);
xnor U25899 (N_25899,N_23733,N_20301);
xor U25900 (N_25900,N_21223,N_18954);
nand U25901 (N_25901,N_21979,N_22949);
nor U25902 (N_25902,N_21976,N_21796);
nor U25903 (N_25903,N_21535,N_21276);
and U25904 (N_25904,N_22932,N_20843);
nand U25905 (N_25905,N_20890,N_21730);
xnor U25906 (N_25906,N_18234,N_22146);
or U25907 (N_25907,N_20967,N_19756);
and U25908 (N_25908,N_23240,N_18253);
xnor U25909 (N_25909,N_23281,N_19516);
xnor U25910 (N_25910,N_20299,N_20024);
nor U25911 (N_25911,N_23821,N_22557);
xnor U25912 (N_25912,N_23846,N_19629);
or U25913 (N_25913,N_21154,N_21041);
nand U25914 (N_25914,N_22174,N_23951);
nor U25915 (N_25915,N_19893,N_21548);
and U25916 (N_25916,N_21178,N_19257);
nor U25917 (N_25917,N_18824,N_20254);
nand U25918 (N_25918,N_19060,N_21055);
and U25919 (N_25919,N_21338,N_23924);
nor U25920 (N_25920,N_18167,N_18049);
or U25921 (N_25921,N_20823,N_21708);
nor U25922 (N_25922,N_23672,N_18778);
or U25923 (N_25923,N_20346,N_21665);
xor U25924 (N_25924,N_18801,N_20675);
nor U25925 (N_25925,N_21935,N_19606);
xor U25926 (N_25926,N_19320,N_22331);
or U25927 (N_25927,N_23539,N_20827);
xnor U25928 (N_25928,N_22997,N_22256);
xor U25929 (N_25929,N_21616,N_21293);
nor U25930 (N_25930,N_23904,N_23061);
xnor U25931 (N_25931,N_19573,N_18555);
nand U25932 (N_25932,N_19222,N_19201);
or U25933 (N_25933,N_23953,N_23787);
xnor U25934 (N_25934,N_23855,N_18429);
nor U25935 (N_25935,N_18788,N_21868);
xor U25936 (N_25936,N_18525,N_22713);
and U25937 (N_25937,N_20521,N_23336);
nand U25938 (N_25938,N_21998,N_21812);
nand U25939 (N_25939,N_21560,N_20612);
nor U25940 (N_25940,N_19565,N_23057);
and U25941 (N_25941,N_21150,N_23758);
or U25942 (N_25942,N_18010,N_22402);
and U25943 (N_25943,N_20090,N_22427);
xnor U25944 (N_25944,N_21427,N_21629);
xor U25945 (N_25945,N_23262,N_23109);
xor U25946 (N_25946,N_20345,N_21044);
and U25947 (N_25947,N_23245,N_18002);
and U25948 (N_25948,N_21016,N_23585);
or U25949 (N_25949,N_22862,N_20892);
nor U25950 (N_25950,N_18343,N_21644);
and U25951 (N_25951,N_18708,N_22753);
nand U25952 (N_25952,N_22649,N_19401);
or U25953 (N_25953,N_18262,N_20754);
nor U25954 (N_25954,N_22852,N_21846);
xor U25955 (N_25955,N_19632,N_22353);
xor U25956 (N_25956,N_19844,N_20862);
and U25957 (N_25957,N_18061,N_20682);
nand U25958 (N_25958,N_21566,N_21209);
xor U25959 (N_25959,N_21626,N_18258);
and U25960 (N_25960,N_20974,N_22978);
and U25961 (N_25961,N_21452,N_22078);
xnor U25962 (N_25962,N_22741,N_21503);
and U25963 (N_25963,N_21564,N_23698);
nand U25964 (N_25964,N_23208,N_19055);
nand U25965 (N_25965,N_18575,N_20749);
or U25966 (N_25966,N_21648,N_22703);
or U25967 (N_25967,N_18201,N_22030);
or U25968 (N_25968,N_20216,N_18213);
nor U25969 (N_25969,N_19277,N_22712);
nor U25970 (N_25970,N_20114,N_22433);
nand U25971 (N_25971,N_22021,N_18571);
and U25972 (N_25972,N_18272,N_19084);
nand U25973 (N_25973,N_21953,N_18198);
nand U25974 (N_25974,N_18605,N_19789);
or U25975 (N_25975,N_21944,N_23748);
xor U25976 (N_25976,N_20493,N_21802);
xor U25977 (N_25977,N_18852,N_22347);
and U25978 (N_25978,N_21894,N_20218);
nor U25979 (N_25979,N_18612,N_23124);
and U25980 (N_25980,N_21840,N_19210);
or U25981 (N_25981,N_21419,N_23514);
or U25982 (N_25982,N_18999,N_23830);
nand U25983 (N_25983,N_20526,N_18285);
xor U25984 (N_25984,N_20640,N_23011);
and U25985 (N_25985,N_19021,N_19066);
nor U25986 (N_25986,N_22738,N_18565);
nor U25987 (N_25987,N_23860,N_20794);
xor U25988 (N_25988,N_19738,N_23489);
or U25989 (N_25989,N_18393,N_19649);
or U25990 (N_25990,N_19945,N_18033);
xor U25991 (N_25991,N_18224,N_18934);
nor U25992 (N_25992,N_20990,N_19503);
xnor U25993 (N_25993,N_22643,N_23451);
or U25994 (N_25994,N_19490,N_22875);
and U25995 (N_25995,N_18389,N_20172);
or U25996 (N_25996,N_19698,N_20446);
nor U25997 (N_25997,N_23945,N_18497);
xnor U25998 (N_25998,N_20026,N_23712);
and U25999 (N_25999,N_21032,N_21978);
and U26000 (N_26000,N_20519,N_22126);
and U26001 (N_26001,N_18882,N_20453);
nor U26002 (N_26002,N_23209,N_22295);
nor U26003 (N_26003,N_21679,N_23982);
and U26004 (N_26004,N_18673,N_18964);
nand U26005 (N_26005,N_18372,N_23731);
and U26006 (N_26006,N_18006,N_18923);
and U26007 (N_26007,N_23172,N_21250);
nand U26008 (N_26008,N_20145,N_18187);
nand U26009 (N_26009,N_19592,N_22204);
nand U26010 (N_26010,N_23764,N_23318);
and U26011 (N_26011,N_21873,N_20231);
or U26012 (N_26012,N_22897,N_18452);
xnor U26013 (N_26013,N_20213,N_18710);
or U26014 (N_26014,N_23025,N_22160);
nor U26015 (N_26015,N_21767,N_23056);
nand U26016 (N_26016,N_23382,N_23927);
nor U26017 (N_26017,N_23287,N_20625);
or U26018 (N_26018,N_19258,N_19539);
or U26019 (N_26019,N_19522,N_20825);
nor U26020 (N_26020,N_22812,N_20800);
and U26021 (N_26021,N_23745,N_23879);
and U26022 (N_26022,N_21187,N_21301);
nor U26023 (N_26023,N_20517,N_22303);
and U26024 (N_26024,N_19791,N_23805);
nand U26025 (N_26025,N_18731,N_22128);
nand U26026 (N_26026,N_21164,N_18079);
and U26027 (N_26027,N_22228,N_20242);
xor U26028 (N_26028,N_23427,N_20361);
nand U26029 (N_26029,N_21818,N_18230);
or U26030 (N_26030,N_20619,N_22096);
xor U26031 (N_26031,N_21752,N_19296);
nor U26032 (N_26032,N_18800,N_20077);
nand U26033 (N_26033,N_20204,N_20304);
or U26034 (N_26034,N_22681,N_18850);
and U26035 (N_26035,N_19097,N_22890);
nand U26036 (N_26036,N_20637,N_22390);
xor U26037 (N_26037,N_21175,N_20530);
nand U26038 (N_26038,N_18865,N_22285);
and U26039 (N_26039,N_23950,N_20158);
or U26040 (N_26040,N_18969,N_20897);
xor U26041 (N_26041,N_23685,N_20787);
or U26042 (N_26042,N_19420,N_21199);
nor U26043 (N_26043,N_23973,N_23981);
xor U26044 (N_26044,N_23490,N_22578);
or U26045 (N_26045,N_21342,N_22686);
or U26046 (N_26046,N_22859,N_22797);
nand U26047 (N_26047,N_18369,N_19126);
nand U26048 (N_26048,N_19068,N_22224);
nand U26049 (N_26049,N_20380,N_21815);
and U26050 (N_26050,N_22573,N_19119);
or U26051 (N_26051,N_22940,N_22947);
nand U26052 (N_26052,N_18604,N_22272);
or U26053 (N_26053,N_22266,N_18548);
and U26054 (N_26054,N_19992,N_20592);
nand U26055 (N_26055,N_19502,N_19445);
nor U26056 (N_26056,N_21555,N_18873);
and U26057 (N_26057,N_18817,N_20246);
and U26058 (N_26058,N_21377,N_19200);
xor U26059 (N_26059,N_22762,N_20657);
and U26060 (N_26060,N_21709,N_23642);
nor U26061 (N_26061,N_22925,N_19388);
nor U26062 (N_26062,N_22282,N_19540);
nor U26063 (N_26063,N_20065,N_21239);
nor U26064 (N_26064,N_23592,N_23984);
xnor U26065 (N_26065,N_23041,N_18931);
or U26066 (N_26066,N_18626,N_23052);
nand U26067 (N_26067,N_20262,N_19672);
xor U26068 (N_26068,N_18647,N_23660);
xnor U26069 (N_26069,N_21358,N_23403);
and U26070 (N_26070,N_23875,N_22831);
nand U26071 (N_26071,N_22027,N_18965);
nor U26072 (N_26072,N_20111,N_19142);
nand U26073 (N_26073,N_21353,N_22509);
or U26074 (N_26074,N_18490,N_22680);
nor U26075 (N_26075,N_21360,N_23519);
nand U26076 (N_26076,N_23233,N_22197);
xnor U26077 (N_26077,N_22461,N_23419);
nor U26078 (N_26078,N_22552,N_23020);
nor U26079 (N_26079,N_22794,N_20144);
or U26080 (N_26080,N_23876,N_19554);
nor U26081 (N_26081,N_22903,N_23587);
nor U26082 (N_26082,N_20486,N_18086);
nand U26083 (N_26083,N_20616,N_23425);
nor U26084 (N_26084,N_19089,N_22498);
or U26085 (N_26085,N_22043,N_23992);
nand U26086 (N_26086,N_20622,N_22845);
or U26087 (N_26087,N_18687,N_22956);
xnor U26088 (N_26088,N_20632,N_23738);
or U26089 (N_26089,N_20898,N_21670);
or U26090 (N_26090,N_23813,N_20894);
nand U26091 (N_26091,N_20638,N_22122);
nand U26092 (N_26092,N_18868,N_21344);
nand U26093 (N_26093,N_19121,N_20986);
nand U26094 (N_26094,N_20721,N_18694);
and U26095 (N_26095,N_20806,N_23771);
xnor U26096 (N_26096,N_22171,N_20600);
nand U26097 (N_26097,N_18321,N_22676);
and U26098 (N_26098,N_23931,N_23825);
xnor U26099 (N_26099,N_22683,N_20459);
or U26100 (N_26100,N_21781,N_18421);
or U26101 (N_26101,N_22328,N_23707);
nor U26102 (N_26102,N_19233,N_22066);
nor U26103 (N_26103,N_19969,N_19599);
nand U26104 (N_26104,N_20234,N_18237);
nand U26105 (N_26105,N_18981,N_20660);
and U26106 (N_26106,N_20190,N_21323);
or U26107 (N_26107,N_20904,N_19390);
nor U26108 (N_26108,N_18380,N_21666);
xnor U26109 (N_26109,N_20133,N_19938);
nand U26110 (N_26110,N_22511,N_18024);
nor U26111 (N_26111,N_23542,N_23885);
nor U26112 (N_26112,N_19402,N_22184);
or U26113 (N_26113,N_21462,N_19792);
or U26114 (N_26114,N_19301,N_22950);
nor U26115 (N_26115,N_21977,N_18388);
nor U26116 (N_26116,N_23683,N_23074);
and U26117 (N_26117,N_21960,N_19936);
xnor U26118 (N_26118,N_23682,N_22388);
or U26119 (N_26119,N_22963,N_19784);
and U26120 (N_26120,N_19942,N_19941);
or U26121 (N_26121,N_18775,N_22103);
xor U26122 (N_26122,N_23290,N_19962);
or U26123 (N_26123,N_21963,N_19274);
and U26124 (N_26124,N_23964,N_21880);
nand U26125 (N_26125,N_18942,N_23920);
or U26126 (N_26126,N_19545,N_23653);
nor U26127 (N_26127,N_21714,N_19700);
and U26128 (N_26128,N_23755,N_22394);
nand U26129 (N_26129,N_23475,N_21614);
xnor U26130 (N_26130,N_21354,N_20499);
or U26131 (N_26131,N_20039,N_19908);
nand U26132 (N_26132,N_18643,N_21464);
xor U26133 (N_26133,N_21202,N_22783);
or U26134 (N_26134,N_19860,N_18913);
and U26135 (N_26135,N_21057,N_21274);
or U26136 (N_26136,N_22194,N_18208);
and U26137 (N_26137,N_21421,N_20370);
nand U26138 (N_26138,N_18464,N_18080);
and U26139 (N_26139,N_23002,N_19765);
or U26140 (N_26140,N_19770,N_20748);
nor U26141 (N_26141,N_22392,N_23203);
and U26142 (N_26142,N_23157,N_18679);
nand U26143 (N_26143,N_19825,N_20253);
nand U26144 (N_26144,N_18890,N_20225);
nor U26145 (N_26145,N_21628,N_20713);
xor U26146 (N_26146,N_18040,N_23834);
and U26147 (N_26147,N_18640,N_20188);
and U26148 (N_26148,N_21671,N_19524);
xnor U26149 (N_26149,N_18353,N_23354);
nor U26150 (N_26150,N_21561,N_18155);
or U26151 (N_26151,N_20647,N_22933);
nand U26152 (N_26152,N_23461,N_22003);
and U26153 (N_26153,N_18512,N_18150);
and U26154 (N_26154,N_22732,N_21152);
nor U26155 (N_26155,N_18459,N_20932);
or U26156 (N_26156,N_22088,N_19901);
nand U26157 (N_26157,N_18674,N_19568);
xnor U26158 (N_26158,N_21865,N_20331);
xnor U26159 (N_26159,N_23636,N_23835);
xor U26160 (N_26160,N_23315,N_18085);
nand U26161 (N_26161,N_20022,N_22067);
or U26162 (N_26162,N_20343,N_22646);
and U26163 (N_26163,N_18434,N_20430);
or U26164 (N_26164,N_23305,N_18088);
nor U26165 (N_26165,N_19056,N_20703);
nor U26166 (N_26166,N_23242,N_23691);
nor U26167 (N_26167,N_20390,N_18919);
and U26168 (N_26168,N_22355,N_19497);
or U26169 (N_26169,N_20575,N_23669);
nand U26170 (N_26170,N_20875,N_19441);
and U26171 (N_26171,N_18279,N_20183);
nand U26172 (N_26172,N_22185,N_23486);
and U26173 (N_26173,N_22036,N_22287);
nand U26174 (N_26174,N_23383,N_23471);
and U26175 (N_26175,N_22210,N_18755);
and U26176 (N_26176,N_21173,N_18487);
nand U26177 (N_26177,N_20266,N_23483);
or U26178 (N_26178,N_23100,N_18067);
and U26179 (N_26179,N_21497,N_21138);
xor U26180 (N_26180,N_18390,N_18111);
nor U26181 (N_26181,N_21756,N_23394);
nor U26182 (N_26182,N_18851,N_18549);
or U26183 (N_26183,N_23129,N_19125);
nor U26184 (N_26184,N_18574,N_21035);
or U26185 (N_26185,N_23381,N_22418);
nor U26186 (N_26186,N_23512,N_23316);
and U26187 (N_26187,N_23711,N_19523);
or U26188 (N_26188,N_22652,N_20123);
or U26189 (N_26189,N_20944,N_19633);
nor U26190 (N_26190,N_18783,N_19430);
nor U26191 (N_26191,N_18701,N_22995);
xor U26192 (N_26192,N_19619,N_18550);
or U26193 (N_26193,N_20500,N_20429);
and U26194 (N_26194,N_20599,N_18846);
nand U26195 (N_26195,N_18918,N_19019);
xor U26196 (N_26196,N_21634,N_21827);
nand U26197 (N_26197,N_21662,N_23773);
or U26198 (N_26198,N_21950,N_23017);
nand U26199 (N_26199,N_22790,N_18240);
and U26200 (N_26200,N_19673,N_22253);
nor U26201 (N_26201,N_19111,N_21801);
xnor U26202 (N_26202,N_23730,N_23547);
and U26203 (N_26203,N_19930,N_22191);
or U26204 (N_26204,N_20155,N_22941);
and U26205 (N_26205,N_19452,N_23081);
or U26206 (N_26206,N_22760,N_23321);
nor U26207 (N_26207,N_23693,N_18572);
or U26208 (N_26208,N_20358,N_18711);
or U26209 (N_26209,N_21355,N_21807);
nand U26210 (N_26210,N_20724,N_18303);
xor U26211 (N_26211,N_18764,N_23373);
or U26212 (N_26212,N_22150,N_22840);
xnor U26213 (N_26213,N_19443,N_22594);
nand U26214 (N_26214,N_19831,N_20215);
xor U26215 (N_26215,N_19072,N_19780);
and U26216 (N_26216,N_23556,N_18900);
or U26217 (N_26217,N_19935,N_20045);
nand U26218 (N_26218,N_18156,N_19748);
and U26219 (N_26219,N_20679,N_19460);
or U26220 (N_26220,N_19807,N_23150);
nor U26221 (N_26221,N_18671,N_22252);
or U26222 (N_26222,N_22701,N_20762);
xor U26223 (N_26223,N_23994,N_22236);
nor U26224 (N_26224,N_18182,N_21376);
nand U26225 (N_26225,N_23445,N_22533);
nand U26226 (N_26226,N_19515,N_23774);
or U26227 (N_26227,N_22610,N_19336);
nor U26228 (N_26228,N_19293,N_19384);
or U26229 (N_26229,N_18529,N_18418);
and U26230 (N_26230,N_20578,N_22662);
nand U26231 (N_26231,N_23325,N_21690);
xnor U26232 (N_26232,N_20449,N_23479);
nor U26233 (N_26233,N_20561,N_23626);
or U26234 (N_26234,N_21791,N_19609);
or U26235 (N_26235,N_22560,N_23092);
or U26236 (N_26236,N_21992,N_20261);
nor U26237 (N_26237,N_18373,N_18880);
and U26238 (N_26238,N_21967,N_18140);
or U26239 (N_26239,N_22563,N_22575);
or U26240 (N_26240,N_21808,N_22700);
xor U26241 (N_26241,N_19648,N_23703);
and U26242 (N_26242,N_23870,N_19988);
nor U26243 (N_26243,N_22793,N_20296);
nand U26244 (N_26244,N_18937,N_23271);
or U26245 (N_26245,N_20419,N_22480);
nand U26246 (N_26246,N_21688,N_19758);
or U26247 (N_26247,N_19467,N_18215);
or U26248 (N_26248,N_18475,N_20567);
and U26249 (N_26249,N_19624,N_22008);
nand U26250 (N_26250,N_18802,N_20235);
nor U26251 (N_26251,N_20615,N_19112);
and U26252 (N_26252,N_20416,N_23900);
nor U26253 (N_26253,N_23194,N_18028);
and U26254 (N_26254,N_19891,N_18727);
nor U26255 (N_26255,N_19325,N_20258);
xnor U26256 (N_26256,N_23643,N_19586);
and U26257 (N_26257,N_21443,N_19003);
or U26258 (N_26258,N_23446,N_22215);
nor U26259 (N_26259,N_21874,N_21370);
nand U26260 (N_26260,N_19315,N_19760);
nor U26261 (N_26261,N_20129,N_22339);
nand U26262 (N_26262,N_22042,N_21922);
xor U26263 (N_26263,N_21002,N_22605);
nor U26264 (N_26264,N_22663,N_19899);
xor U26265 (N_26265,N_22528,N_22929);
nand U26266 (N_26266,N_18885,N_21983);
nand U26267 (N_26267,N_20757,N_23366);
xor U26268 (N_26268,N_19695,N_23254);
nor U26269 (N_26269,N_21136,N_23423);
and U26270 (N_26270,N_21839,N_20337);
xnor U26271 (N_26271,N_20646,N_18231);
nand U26272 (N_26272,N_20947,N_23218);
nand U26273 (N_26273,N_23831,N_21010);
or U26274 (N_26274,N_19946,N_18470);
xor U26275 (N_26275,N_18096,N_20508);
nand U26276 (N_26276,N_19610,N_22412);
xnor U26277 (N_26277,N_19486,N_19102);
nand U26278 (N_26278,N_20137,N_21224);
nor U26279 (N_26279,N_20034,N_20537);
xnor U26280 (N_26280,N_18284,N_18084);
nor U26281 (N_26281,N_21040,N_23798);
nand U26282 (N_26282,N_21524,N_21478);
nand U26283 (N_26283,N_19369,N_22901);
nand U26284 (N_26284,N_22817,N_21331);
or U26285 (N_26285,N_18302,N_22421);
nor U26286 (N_26286,N_19704,N_21062);
or U26287 (N_26287,N_19137,N_18920);
xor U26288 (N_26288,N_19785,N_21487);
nand U26289 (N_26289,N_19840,N_18431);
and U26290 (N_26290,N_23515,N_20274);
xnor U26291 (N_26291,N_22620,N_19712);
xnor U26292 (N_26292,N_18189,N_19279);
nor U26293 (N_26293,N_19968,N_20930);
and U26294 (N_26294,N_22719,N_20772);
and U26295 (N_26295,N_18860,N_20935);
xnor U26296 (N_26296,N_21504,N_18151);
and U26297 (N_26297,N_22137,N_23396);
nand U26298 (N_26298,N_20197,N_22581);
nor U26299 (N_26299,N_18171,N_19032);
or U26300 (N_26300,N_20185,N_18795);
and U26301 (N_26301,N_20885,N_23431);
xnor U26302 (N_26302,N_21604,N_23051);
or U26303 (N_26303,N_23230,N_23146);
nand U26304 (N_26304,N_19678,N_19980);
nor U26305 (N_26305,N_22696,N_18729);
nor U26306 (N_26306,N_18172,N_21450);
xor U26307 (N_26307,N_21499,N_23253);
or U26308 (N_26308,N_23390,N_21005);
and U26309 (N_26309,N_23120,N_18206);
or U26310 (N_26310,N_22270,N_20492);
nand U26311 (N_26311,N_18467,N_22894);
nor U26312 (N_26312,N_20635,N_21432);
nor U26313 (N_26313,N_22217,N_20711);
or U26314 (N_26314,N_23324,N_18635);
or U26315 (N_26315,N_20654,N_18101);
and U26316 (N_26316,N_23841,N_23659);
nand U26317 (N_26317,N_19122,N_22341);
or U26318 (N_26318,N_20747,N_23457);
or U26319 (N_26319,N_22425,N_20882);
nor U26320 (N_26320,N_18551,N_22502);
nor U26321 (N_26321,N_21893,N_18386);
xor U26322 (N_26322,N_21620,N_21247);
and U26323 (N_26323,N_23332,N_21074);
nand U26324 (N_26324,N_19877,N_18653);
xnor U26325 (N_26325,N_18544,N_22161);
nor U26326 (N_26326,N_21214,N_20347);
xor U26327 (N_26327,N_18973,N_21201);
nor U26328 (N_26328,N_19574,N_21115);
and U26329 (N_26329,N_21790,N_23395);
and U26330 (N_26330,N_19133,N_20798);
nor U26331 (N_26331,N_21400,N_18177);
xnor U26332 (N_26332,N_21077,N_22207);
and U26333 (N_26333,N_18175,N_21114);
and U26334 (N_26334,N_23881,N_22484);
nor U26335 (N_26335,N_18806,N_23882);
and U26336 (N_26336,N_19431,N_20293);
or U26337 (N_26337,N_18007,N_20661);
xor U26338 (N_26338,N_21483,N_18692);
nand U26339 (N_26339,N_22751,N_21898);
or U26340 (N_26340,N_18031,N_21601);
nor U26341 (N_26341,N_18786,N_23777);
or U26342 (N_26342,N_21937,N_22249);
or U26343 (N_26343,N_23802,N_23084);
and U26344 (N_26344,N_19660,N_19873);
xor U26345 (N_26345,N_19082,N_20352);
and U26346 (N_26346,N_22245,N_20087);
and U26347 (N_26347,N_19559,N_22916);
and U26348 (N_26348,N_22424,N_19528);
or U26349 (N_26349,N_22945,N_18407);
or U26350 (N_26350,N_18547,N_23175);
nor U26351 (N_26351,N_21919,N_18972);
nand U26352 (N_26352,N_20035,N_22492);
nand U26353 (N_26353,N_23770,N_21493);
xnor U26354 (N_26354,N_18092,N_22954);
or U26355 (N_26355,N_18747,N_23076);
nand U26356 (N_26356,N_23675,N_19561);
xnor U26357 (N_26357,N_19575,N_23890);
and U26358 (N_26358,N_22755,N_20482);
or U26359 (N_26359,N_18888,N_21254);
nor U26360 (N_26360,N_19972,N_19856);
nand U26361 (N_26361,N_22023,N_19310);
nand U26362 (N_26362,N_20391,N_20954);
or U26363 (N_26363,N_21947,N_21835);
nor U26364 (N_26364,N_20490,N_20175);
nand U26365 (N_26365,N_18695,N_19981);
nand U26366 (N_26366,N_19235,N_18191);
and U26367 (N_26367,N_22877,N_23662);
nor U26368 (N_26368,N_23935,N_20548);
or U26369 (N_26369,N_20401,N_22376);
nand U26370 (N_26370,N_19993,N_19967);
nand U26371 (N_26371,N_20853,N_23224);
and U26372 (N_26372,N_20067,N_19722);
xnor U26373 (N_26373,N_18709,N_20047);
nor U26374 (N_26374,N_18238,N_20442);
nor U26375 (N_26375,N_18877,N_20624);
nand U26376 (N_26376,N_19714,N_21631);
nor U26377 (N_26377,N_19868,N_20392);
and U26378 (N_26378,N_20305,N_18896);
or U26379 (N_26379,N_21480,N_20872);
or U26380 (N_26380,N_23345,N_21704);
and U26381 (N_26381,N_19034,N_21740);
nor U26382 (N_26382,N_18065,N_20146);
nor U26383 (N_26383,N_20128,N_22157);
xor U26384 (N_26384,N_22113,N_19104);
nand U26385 (N_26385,N_22884,N_22106);
xnor U26386 (N_26386,N_20995,N_18301);
and U26387 (N_26387,N_19631,N_18620);
xnor U26388 (N_26388,N_22855,N_22988);
or U26389 (N_26389,N_21291,N_18316);
or U26390 (N_26390,N_20685,N_21165);
or U26391 (N_26391,N_23996,N_19587);
nor U26392 (N_26392,N_23525,N_19352);
nand U26393 (N_26393,N_20439,N_23803);
nor U26394 (N_26394,N_22930,N_19863);
nand U26395 (N_26395,N_22918,N_22440);
nand U26396 (N_26396,N_21957,N_21200);
nor U26397 (N_26397,N_20072,N_21772);
and U26398 (N_26398,N_23439,N_20955);
nor U26399 (N_26399,N_18117,N_18589);
nand U26400 (N_26400,N_23468,N_18197);
xor U26401 (N_26401,N_21488,N_19464);
nand U26402 (N_26402,N_23477,N_22699);
and U26403 (N_26403,N_19370,N_23757);
nand U26404 (N_26404,N_22261,N_18827);
xnor U26405 (N_26405,N_21004,N_23583);
nor U26406 (N_26406,N_18680,N_20901);
and U26407 (N_26407,N_23538,N_23910);
or U26408 (N_26408,N_20584,N_18577);
and U26409 (N_26409,N_22401,N_20736);
or U26410 (N_26410,N_19811,N_19534);
and U26411 (N_26411,N_23800,N_21438);
nand U26412 (N_26412,N_19688,N_20601);
and U26413 (N_26413,N_18762,N_19620);
and U26414 (N_26414,N_23235,N_21528);
xor U26415 (N_26415,N_23909,N_21769);
and U26416 (N_26416,N_21996,N_23206);
xnor U26417 (N_26417,N_20468,N_23080);
nand U26418 (N_26418,N_23083,N_19069);
or U26419 (N_26419,N_23917,N_19092);
xor U26420 (N_26420,N_23466,N_22761);
or U26421 (N_26421,N_22709,N_21127);
and U26422 (N_26422,N_23925,N_23493);
and U26423 (N_26423,N_18300,N_22352);
nand U26424 (N_26424,N_20669,N_18899);
or U26425 (N_26425,N_20927,N_21672);
nand U26426 (N_26426,N_18226,N_18160);
nor U26427 (N_26427,N_23564,N_21975);
and U26428 (N_26428,N_19281,N_20103);
nand U26429 (N_26429,N_19147,N_19944);
and U26430 (N_26430,N_22702,N_23822);
or U26431 (N_26431,N_20195,N_22912);
nor U26432 (N_26432,N_22545,N_23053);
or U26433 (N_26433,N_20150,N_18227);
nand U26434 (N_26434,N_19622,N_20251);
and U26435 (N_26435,N_19876,N_20023);
nand U26436 (N_26436,N_22246,N_20791);
nor U26437 (N_26437,N_23263,N_23125);
nor U26438 (N_26438,N_22942,N_21570);
and U26439 (N_26439,N_22101,N_23898);
and U26440 (N_26440,N_19598,N_18949);
nor U26441 (N_26441,N_21507,N_21441);
and U26442 (N_26442,N_23958,N_23244);
or U26443 (N_26443,N_20159,N_22155);
or U26444 (N_26444,N_20771,N_23744);
nand U26445 (N_26445,N_18493,N_20992);
xnor U26446 (N_26446,N_21142,N_19884);
nor U26447 (N_26447,N_23054,N_18469);
xnor U26448 (N_26448,N_20149,N_22459);
nand U26449 (N_26449,N_21211,N_18179);
nand U26450 (N_26450,N_23851,N_18863);
nor U26451 (N_26451,N_19197,N_22407);
nand U26452 (N_26452,N_21145,N_19679);
and U26453 (N_26453,N_20773,N_22465);
xnor U26454 (N_26454,N_23094,N_22134);
nand U26455 (N_26455,N_21871,N_19702);
xnor U26456 (N_26456,N_22744,N_18269);
nor U26457 (N_26457,N_18592,N_19426);
or U26458 (N_26458,N_19282,N_20759);
nand U26459 (N_26459,N_21735,N_21153);
xor U26460 (N_26460,N_20576,N_23277);
or U26461 (N_26461,N_18142,N_22077);
xor U26462 (N_26462,N_21641,N_21036);
or U26463 (N_26463,N_23361,N_21928);
nor U26464 (N_26464,N_21217,N_23123);
or U26465 (N_26465,N_22453,N_18008);
and U26466 (N_26466,N_21897,N_18257);
or U26467 (N_26467,N_19555,N_22214);
nor U26468 (N_26468,N_23308,N_23709);
nor U26469 (N_26469,N_23481,N_18744);
and U26470 (N_26470,N_19686,N_23215);
nand U26471 (N_26471,N_18045,N_23480);
or U26472 (N_26472,N_20803,N_22247);
nor U26473 (N_26473,N_22800,N_19468);
or U26474 (N_26474,N_21351,N_23658);
and U26475 (N_26475,N_22928,N_19184);
or U26476 (N_26476,N_23086,N_23906);
xor U26477 (N_26477,N_21981,N_21888);
or U26478 (N_26478,N_23926,N_18340);
nand U26479 (N_26479,N_20781,N_18537);
xnor U26480 (N_26480,N_20339,N_18615);
nor U26481 (N_26481,N_19176,N_20471);
or U26482 (N_26482,N_21722,N_21680);
and U26483 (N_26483,N_19247,N_22974);
xor U26484 (N_26484,N_22644,N_21968);
xor U26485 (N_26485,N_20243,N_19625);
nor U26486 (N_26486,N_18029,N_23016);
xnor U26487 (N_26487,N_21018,N_19759);
or U26488 (N_26488,N_18832,N_22351);
or U26489 (N_26489,N_23563,N_23111);
or U26490 (N_26490,N_21108,N_23721);
xnor U26491 (N_26491,N_19685,N_22447);
nor U26492 (N_26492,N_20934,N_18023);
xnor U26493 (N_26493,N_21987,N_22058);
nor U26494 (N_26494,N_19810,N_22619);
nand U26495 (N_26495,N_19306,N_23482);
and U26496 (N_26496,N_18938,N_23850);
or U26497 (N_26497,N_21268,N_22870);
nor U26498 (N_26498,N_20191,N_23131);
and U26499 (N_26499,N_22656,N_21951);
or U26500 (N_26500,N_22145,N_19219);
and U26501 (N_26501,N_18958,N_18864);
xor U26502 (N_26502,N_19297,N_23768);
nor U26503 (N_26503,N_19035,N_19949);
nor U26504 (N_26504,N_18760,N_20881);
xor U26505 (N_26505,N_23663,N_22900);
or U26506 (N_26506,N_18219,N_19549);
or U26507 (N_26507,N_19779,N_19934);
and U26508 (N_26508,N_23632,N_20941);
or U26509 (N_26509,N_22062,N_20902);
xor U26510 (N_26510,N_23765,N_18394);
xor U26511 (N_26511,N_20229,N_21495);
and U26512 (N_26512,N_19366,N_21389);
and U26513 (N_26513,N_18594,N_18425);
nor U26514 (N_26514,N_20179,N_22742);
nor U26515 (N_26515,N_18399,N_18608);
xor U26516 (N_26516,N_19195,N_19613);
xnor U26517 (N_26517,N_20849,N_19259);
nor U26518 (N_26518,N_19658,N_19703);
or U26519 (N_26519,N_19096,N_21774);
nand U26520 (N_26520,N_19739,N_18637);
and U26521 (N_26521,N_20727,N_21017);
nand U26522 (N_26522,N_18350,N_18217);
nand U26523 (N_26523,N_19804,N_19857);
nor U26524 (N_26524,N_18502,N_18169);
or U26525 (N_26525,N_23937,N_22495);
and U26526 (N_26526,N_22132,N_21610);
or U26527 (N_26527,N_19959,N_21762);
nand U26528 (N_26528,N_21446,N_23708);
and U26529 (N_26529,N_20217,N_23654);
xor U26530 (N_26530,N_21191,N_18560);
nand U26531 (N_26531,N_21079,N_21834);
nor U26532 (N_26532,N_19347,N_20764);
nand U26533 (N_26533,N_19921,N_23582);
and U26534 (N_26534,N_20349,N_21159);
xor U26535 (N_26535,N_21784,N_20060);
nor U26536 (N_26536,N_19379,N_22474);
and U26537 (N_26537,N_18038,N_22441);
nand U26538 (N_26538,N_23788,N_23219);
xor U26539 (N_26539,N_22148,N_20049);
nand U26540 (N_26540,N_19039,N_19237);
nand U26541 (N_26541,N_23713,N_18317);
nor U26542 (N_26542,N_21313,N_21713);
xor U26543 (N_26543,N_19635,N_21591);
xnor U26544 (N_26544,N_18026,N_22491);
nor U26545 (N_26545,N_22734,N_22936);
nand U26546 (N_26546,N_22178,N_20142);
and U26547 (N_26547,N_23458,N_21116);
or U26548 (N_26548,N_19774,N_21824);
and U26549 (N_26549,N_19532,N_22826);
nor U26550 (N_26550,N_23853,N_20778);
nor U26551 (N_26551,N_22799,N_18042);
nand U26552 (N_26552,N_19655,N_23207);
nor U26553 (N_26553,N_21160,N_22633);
or U26554 (N_26554,N_22768,N_22889);
xor U26555 (N_26555,N_21225,N_19354);
nand U26556 (N_26556,N_19334,N_20695);
and U26557 (N_26557,N_20348,N_23327);
or U26558 (N_26558,N_22305,N_20378);
xor U26559 (N_26559,N_20808,N_22257);
or U26560 (N_26560,N_21580,N_23734);
xor U26561 (N_26561,N_20546,N_23463);
and U26562 (N_26562,N_21632,N_20761);
nand U26563 (N_26563,N_18651,N_23098);
or U26564 (N_26564,N_22028,N_23849);
or U26565 (N_26565,N_21475,N_19881);
nand U26566 (N_26566,N_18438,N_20066);
nand U26567 (N_26567,N_21729,N_20819);
nor U26568 (N_26568,N_18988,N_23006);
or U26569 (N_26569,N_19058,N_21334);
and U26570 (N_26570,N_18912,N_23274);
nor U26571 (N_26571,N_22172,N_22781);
or U26572 (N_26572,N_19287,N_19659);
nand U26573 (N_26573,N_20750,N_23161);
xor U26574 (N_26574,N_22225,N_23367);
xor U26575 (N_26575,N_19447,N_19506);
and U26576 (N_26576,N_18580,N_22312);
nand U26577 (N_26577,N_21869,N_23248);
nor U26578 (N_26578,N_23908,N_23676);
and U26579 (N_26579,N_20095,N_23799);
or U26580 (N_26580,N_23862,N_20220);
nand U26581 (N_26581,N_18178,N_23836);
xor U26582 (N_26582,N_23988,N_19363);
and U26583 (N_26583,N_19689,N_22886);
or U26584 (N_26584,N_22156,N_23319);
nor U26585 (N_26585,N_20790,N_23729);
xnor U26586 (N_26586,N_20098,N_23341);
and U26587 (N_26587,N_19794,N_19117);
and U26588 (N_26588,N_22879,N_20267);
xnor U26589 (N_26589,N_22343,N_20858);
xor U26590 (N_26590,N_20286,N_20117);
nand U26591 (N_26591,N_23752,N_18122);
and U26592 (N_26592,N_18634,N_19504);
xor U26593 (N_26593,N_18769,N_18052);
nor U26594 (N_26594,N_23886,N_20180);
or U26595 (N_26595,N_20569,N_21980);
nor U26596 (N_26596,N_22543,N_20367);
xnor U26597 (N_26597,N_22346,N_23521);
or U26598 (N_26598,N_21695,N_20717);
nor U26599 (N_26599,N_18543,N_21107);
and U26600 (N_26600,N_23977,N_21205);
xnor U26601 (N_26601,N_19462,N_18091);
nor U26602 (N_26602,N_22514,N_22772);
and U26603 (N_26603,N_23251,N_20926);
xnor U26604 (N_26604,N_19215,N_18532);
nor U26605 (N_26605,N_18702,N_19671);
nand U26606 (N_26606,N_21278,N_18712);
nand U26607 (N_26607,N_21221,N_20351);
xnor U26608 (N_26608,N_22516,N_20350);
and U26609 (N_26609,N_23496,N_22209);
and U26610 (N_26610,N_20953,N_20563);
nand U26611 (N_26611,N_20334,N_19662);
nand U26612 (N_26612,N_23301,N_22450);
or U26613 (N_26613,N_18344,N_18926);
nor U26614 (N_26614,N_22136,N_19543);
or U26615 (N_26615,N_18194,N_20831);
or U26616 (N_26616,N_22281,N_18699);
nor U26617 (N_26617,N_19278,N_19839);
nand U26618 (N_26618,N_21072,N_18297);
nor U26619 (N_26619,N_18685,N_19404);
and U26620 (N_26620,N_21719,N_20463);
nor U26621 (N_26621,N_20667,N_20359);
nand U26622 (N_26622,N_18720,N_19687);
xor U26623 (N_26623,N_23548,N_21844);
nor U26624 (N_26624,N_18907,N_20598);
xnor U26625 (N_26625,N_20896,N_20058);
nor U26626 (N_26626,N_23789,N_22523);
and U26627 (N_26627,N_21080,N_20275);
or U26628 (N_26628,N_18893,N_19086);
nand U26629 (N_26629,N_23995,N_20683);
nand U26630 (N_26630,N_19213,N_21111);
and U26631 (N_26631,N_22921,N_23612);
and U26632 (N_26632,N_20693,N_22714);
or U26633 (N_26633,N_18582,N_22504);
nor U26634 (N_26634,N_19977,N_21298);
and U26635 (N_26635,N_22708,N_21275);
nor U26636 (N_26636,N_22430,N_21265);
nor U26637 (N_26637,N_18364,N_21716);
xor U26638 (N_26638,N_19514,N_20905);
nor U26639 (N_26639,N_22896,N_18220);
xor U26640 (N_26640,N_20285,N_23753);
and U26641 (N_26641,N_22835,N_20813);
nand U26642 (N_26642,N_21588,N_18854);
nand U26643 (N_26643,N_18476,N_21469);
xnor U26644 (N_26644,N_23640,N_18519);
nor U26645 (N_26645,N_21155,N_22072);
xor U26646 (N_26646,N_21119,N_19841);
nand U26647 (N_26647,N_23866,N_21039);
or U26648 (N_26648,N_22647,N_23448);
or U26649 (N_26649,N_18051,N_22414);
or U26650 (N_26650,N_19862,N_20292);
nand U26651 (N_26651,N_18356,N_23848);
nand U26652 (N_26652,N_19365,N_19251);
nand U26653 (N_26653,N_21683,N_22278);
or U26654 (N_26654,N_22910,N_21859);
nand U26655 (N_26655,N_23328,N_20511);
nand U26656 (N_26656,N_19078,N_23792);
or U26657 (N_26657,N_21426,N_18309);
nor U26658 (N_26658,N_21181,N_20051);
nor U26659 (N_26659,N_23077,N_21206);
and U26660 (N_26660,N_20589,N_21918);
or U26661 (N_26661,N_19294,N_23575);
or U26662 (N_26662,N_19338,N_22810);
or U26663 (N_26663,N_22476,N_18081);
nand U26664 (N_26664,N_22966,N_21582);
nand U26665 (N_26665,N_20168,N_21995);
nand U26666 (N_26666,N_22508,N_18881);
nor U26667 (N_26667,N_21608,N_22968);
or U26668 (N_26668,N_20893,N_21549);
nand U26669 (N_26669,N_23070,N_21103);
nor U26670 (N_26670,N_22301,N_22996);
nand U26671 (N_26671,N_19772,N_19953);
nand U26672 (N_26672,N_19787,N_19067);
or U26673 (N_26673,N_21379,N_20652);
or U26674 (N_26674,N_19449,N_19152);
xnor U26675 (N_26675,N_21410,N_20450);
and U26676 (N_26676,N_20303,N_23164);
nand U26677 (N_26677,N_21887,N_21067);
nand U26678 (N_26678,N_21494,N_20977);
or U26679 (N_26679,N_21048,N_19436);
and U26680 (N_26680,N_18933,N_22000);
nand U26681 (N_26681,N_21059,N_20088);
nand U26682 (N_26682,N_22381,N_19852);
nor U26683 (N_26683,N_22824,N_23551);
xnor U26684 (N_26684,N_20457,N_21434);
xor U26685 (N_26685,N_20556,N_21013);
xor U26686 (N_26686,N_21192,N_22655);
nand U26687 (N_26687,N_23673,N_18170);
xor U26688 (N_26688,N_22130,N_19675);
nor U26689 (N_26689,N_18591,N_23156);
nand U26690 (N_26690,N_20477,N_22248);
or U26691 (N_26691,N_21463,N_18335);
nor U26692 (N_26692,N_18454,N_19776);
or U26693 (N_26693,N_19424,N_22458);
and U26694 (N_26694,N_19355,N_20388);
nor U26695 (N_26695,N_21300,N_19973);
or U26696 (N_26696,N_21297,N_20971);
or U26697 (N_26697,N_21567,N_20454);
nor U26698 (N_26698,N_21530,N_18696);
nand U26699 (N_26699,N_19950,N_20245);
and U26700 (N_26700,N_20618,N_18588);
and U26701 (N_26701,N_23591,N_22895);
xor U26702 (N_26702,N_21934,N_19327);
nor U26703 (N_26703,N_19010,N_22455);
and U26704 (N_26704,N_20260,N_20952);
nand U26705 (N_26705,N_18466,N_22993);
nand U26706 (N_26706,N_19762,N_22337);
xor U26707 (N_26707,N_20200,N_18614);
and U26708 (N_26708,N_18479,N_22085);
and U26709 (N_26709,N_22370,N_23569);
nand U26710 (N_26710,N_18616,N_19114);
xor U26711 (N_26711,N_21189,N_21958);
nor U26712 (N_26712,N_18581,N_21125);
or U26713 (N_26713,N_23722,N_22685);
nor U26714 (N_26714,N_23202,N_19526);
xnor U26715 (N_26715,N_21363,N_22616);
nor U26716 (N_26716,N_23212,N_23096);
and U26717 (N_26717,N_18631,N_20520);
or U26718 (N_26718,N_23214,N_23541);
xor U26719 (N_26719,N_22595,N_18261);
or U26720 (N_26720,N_20009,N_21359);
and U26721 (N_26721,N_18424,N_23761);
xnor U26722 (N_26722,N_23013,N_20071);
nand U26723 (N_26723,N_20461,N_21058);
nor U26724 (N_26724,N_23393,N_21437);
xnor U26725 (N_26725,N_20666,N_21468);
or U26726 (N_26726,N_19023,N_23116);
nand U26727 (N_26727,N_20883,N_21472);
nand U26728 (N_26728,N_19480,N_20665);
xnor U26729 (N_26729,N_18363,N_22490);
nor U26730 (N_26730,N_20547,N_19389);
or U26731 (N_26731,N_23633,N_22344);
nor U26732 (N_26732,N_21696,N_20306);
nor U26733 (N_26733,N_20273,N_19202);
nor U26734 (N_26734,N_21511,N_18724);
nand U26735 (N_26735,N_23852,N_21451);
xnor U26736 (N_26736,N_18400,N_19025);
nand U26737 (N_26737,N_22527,N_18742);
and U26738 (N_26738,N_21366,N_18378);
nor U26739 (N_26739,N_23343,N_18743);
nor U26740 (N_26740,N_19153,N_19966);
nand U26741 (N_26741,N_22482,N_21467);
or U26742 (N_26742,N_23353,N_18531);
nor U26743 (N_26743,N_21541,N_23878);
nor U26744 (N_26744,N_19642,N_22657);
nor U26745 (N_26745,N_18598,N_23820);
nor U26746 (N_26746,N_23817,N_18106);
nor U26747 (N_26747,N_19331,N_22814);
and U26748 (N_26748,N_21556,N_20415);
nand U26749 (N_26749,N_20605,N_22955);
and U26750 (N_26750,N_18118,N_20375);
nand U26751 (N_26751,N_22375,N_19517);
xnor U26752 (N_26752,N_20942,N_22807);
nor U26753 (N_26753,N_20909,N_20597);
xnor U26754 (N_26754,N_20824,N_20414);
nor U26755 (N_26755,N_19668,N_23692);
nand U26756 (N_26756,N_22354,N_22598);
nand U26757 (N_26757,N_18141,N_18283);
and U26758 (N_26758,N_20147,N_23380);
nor U26759 (N_26759,N_21393,N_20694);
nor U26760 (N_26760,N_23442,N_21705);
nand U26761 (N_26761,N_21364,N_20760);
or U26762 (N_26762,N_18004,N_19914);
and U26763 (N_26763,N_22671,N_22179);
and U26764 (N_26764,N_19913,N_19209);
or U26765 (N_26765,N_20796,N_21991);
or U26766 (N_26766,N_18410,N_20485);
or U26767 (N_26767,N_18192,N_18066);
nand U26768 (N_26768,N_20672,N_20042);
nor U26769 (N_26769,N_20842,N_18763);
nor U26770 (N_26770,N_18599,N_21860);
nor U26771 (N_26771,N_20577,N_19087);
or U26772 (N_26772,N_20048,N_20131);
nand U26773 (N_26773,N_20420,N_19083);
nand U26774 (N_26774,N_18044,N_19742);
and U26775 (N_26775,N_22593,N_21245);
and U26776 (N_26776,N_22018,N_21285);
xnor U26777 (N_26777,N_22757,N_22431);
xor U26778 (N_26778,N_21798,N_19611);
nor U26779 (N_26779,N_18148,N_18903);
xnor U26780 (N_26780,N_19861,N_20151);
and U26781 (N_26781,N_21337,N_22340);
and U26782 (N_26782,N_21755,N_20013);
and U26783 (N_26783,N_19268,N_20755);
xor U26784 (N_26784,N_18740,N_19607);
and U26785 (N_26785,N_18630,N_23435);
nand U26786 (N_26786,N_23012,N_22678);
xnor U26787 (N_26787,N_19314,N_21759);
and U26788 (N_26788,N_18656,N_19291);
nand U26789 (N_26789,N_21623,N_23586);
nor U26790 (N_26790,N_22182,N_23749);
nand U26791 (N_26791,N_20495,N_19905);
nand U26792 (N_26792,N_18255,N_20322);
and U26793 (N_26793,N_19530,N_19692);
xnor U26794 (N_26794,N_18781,N_20341);
xor U26795 (N_26795,N_21851,N_20338);
and U26796 (N_26796,N_23283,N_21500);
and U26797 (N_26797,N_21602,N_21423);
and U26798 (N_26798,N_19715,N_20763);
nor U26799 (N_26799,N_18648,N_20402);
nand U26800 (N_26800,N_21373,N_23021);
xor U26801 (N_26801,N_23896,N_23714);
and U26802 (N_26802,N_20899,N_18655);
nand U26803 (N_26803,N_23531,N_21515);
and U26804 (N_26804,N_22629,N_18722);
and U26805 (N_26805,N_22138,N_22416);
xnor U26806 (N_26806,N_21430,N_18822);
or U26807 (N_26807,N_23718,N_20987);
nor U26808 (N_26808,N_22422,N_18116);
nor U26809 (N_26809,N_19463,N_21903);
xnor U26810 (N_26810,N_22715,N_21571);
xnor U26811 (N_26811,N_19051,N_19837);
xnor U26812 (N_26812,N_19007,N_22255);
and U26813 (N_26813,N_18567,N_21146);
and U26814 (N_26814,N_20978,N_22811);
nand U26815 (N_26815,N_20244,N_20207);
or U26816 (N_26816,N_20161,N_23985);
nor U26817 (N_26817,N_20753,N_22806);
nor U26818 (N_26818,N_20434,N_18784);
nor U26819 (N_26819,N_20908,N_21510);
nor U26820 (N_26820,N_19882,N_22697);
xor U26821 (N_26821,N_21068,N_18810);
or U26822 (N_26822,N_22667,N_20789);
xor U26823 (N_26823,N_21139,N_22727);
nor U26824 (N_26824,N_20318,N_20029);
xnor U26825 (N_26825,N_23513,N_22055);
and U26826 (N_26826,N_22565,N_21910);
and U26827 (N_26827,N_19848,N_21513);
or U26828 (N_26828,N_21837,N_19376);
nand U26829 (N_26829,N_20983,N_18947);
or U26830 (N_26830,N_20811,N_21045);
nand U26831 (N_26831,N_18205,N_20918);
or U26832 (N_26832,N_19986,N_18859);
nand U26833 (N_26833,N_19602,N_23894);
xor U26834 (N_26834,N_18789,N_20302);
or U26835 (N_26835,N_21315,N_22529);
xor U26836 (N_26836,N_19231,N_18136);
nand U26837 (N_26837,N_19749,N_22892);
and U26838 (N_26838,N_19466,N_23256);
nor U26839 (N_26839,N_22736,N_23810);
and U26840 (N_26840,N_18166,N_19302);
nor U26841 (N_26841,N_23899,N_23158);
nor U26842 (N_26842,N_20518,N_20064);
nand U26843 (N_26843,N_22922,N_23700);
and U26844 (N_26844,N_21256,N_22313);
nand U26845 (N_26845,N_23589,N_23018);
or U26846 (N_26846,N_23255,N_21203);
or U26847 (N_26847,N_19434,N_22497);
nand U26848 (N_26848,N_22805,N_19754);
or U26849 (N_26849,N_19229,N_18962);
and U26850 (N_26850,N_21565,N_21594);
xor U26851 (N_26851,N_20737,N_23088);
xnor U26852 (N_26852,N_18263,N_19225);
xnor U26853 (N_26853,N_22076,N_23680);
nand U26854 (N_26854,N_21870,N_21797);
xor U26855 (N_26855,N_19750,N_21020);
or U26856 (N_26856,N_21266,N_21365);
nor U26857 (N_26857,N_19547,N_19193);
xnor U26858 (N_26858,N_19318,N_23971);
or U26859 (N_26859,N_19835,N_22682);
xor U26860 (N_26860,N_22065,N_18889);
or U26861 (N_26861,N_21885,N_23596);
nor U26862 (N_26862,N_18511,N_18645);
and U26863 (N_26863,N_22969,N_20805);
nand U26864 (N_26864,N_19571,N_23459);
nand U26865 (N_26865,N_21350,N_19418);
xnor U26866 (N_26866,N_18991,N_21905);
or U26867 (N_26867,N_21856,N_19907);
and U26868 (N_26868,N_23197,N_22300);
and U26869 (N_26869,N_23195,N_19589);
nor U26870 (N_26870,N_23840,N_21544);
xnor U26871 (N_26871,N_22754,N_19663);
xor U26872 (N_26872,N_18629,N_23615);
and U26873 (N_26873,N_21422,N_19304);
and U26874 (N_26874,N_20005,N_18600);
and U26875 (N_26875,N_18154,N_20283);
nor U26876 (N_26876,N_20780,N_20964);
nand U26877 (N_26877,N_22115,N_22466);
or U26878 (N_26878,N_23119,N_22572);
or U26879 (N_26879,N_19529,N_22935);
nand U26880 (N_26880,N_20073,N_18607);
and U26881 (N_26881,N_23665,N_18785);
and U26882 (N_26882,N_18076,N_23742);
nor U26883 (N_26883,N_23517,N_23162);
and U26884 (N_26884,N_18095,N_23099);
and U26885 (N_26885,N_19307,N_19036);
nor U26886 (N_26886,N_23022,N_22569);
xnor U26887 (N_26887,N_22463,N_18639);
and U26888 (N_26888,N_20326,N_20756);
nand U26889 (N_26889,N_19560,N_19476);
and U26890 (N_26890,N_23520,N_18244);
or U26891 (N_26891,N_20327,N_23042);
or U26892 (N_26892,N_22350,N_22883);
nand U26893 (N_26893,N_21920,N_23960);
or U26894 (N_26894,N_19203,N_23819);
and U26895 (N_26895,N_21086,N_18496);
or U26896 (N_26896,N_19533,N_22609);
nand U26897 (N_26897,N_23861,N_20709);
or U26898 (N_26898,N_19351,N_21303);
nor U26899 (N_26899,N_23921,N_23487);
nor U26900 (N_26900,N_21775,N_18841);
nor U26901 (N_26901,N_23398,N_18698);
nand U26902 (N_26902,N_23645,N_19357);
nor U26903 (N_26903,N_20946,N_22223);
nor U26904 (N_26904,N_22909,N_22920);
or U26905 (N_26905,N_20963,N_19459);
and U26906 (N_26906,N_19764,N_18894);
xnor U26907 (N_26907,N_21597,N_23877);
nand U26908 (N_26908,N_21850,N_23181);
and U26909 (N_26909,N_20643,N_20044);
nand U26910 (N_26910,N_20112,N_22658);
nand U26911 (N_26911,N_23464,N_21583);
nand U26912 (N_26912,N_18427,N_20389);
nand U26913 (N_26913,N_20708,N_22045);
nor U26914 (N_26914,N_23456,N_22276);
nor U26915 (N_26915,N_20473,N_18683);
xor U26916 (N_26916,N_18149,N_18072);
xor U26917 (N_26917,N_22953,N_22084);
or U26918 (N_26918,N_21481,N_22064);
and U26919 (N_26919,N_21896,N_19752);
or U26920 (N_26920,N_22771,N_21194);
or U26921 (N_26921,N_20171,N_20379);
nand U26922 (N_26922,N_21904,N_22277);
nand U26923 (N_26923,N_23780,N_22871);
xor U26924 (N_26924,N_18055,N_22750);
xor U26925 (N_26925,N_22082,N_18678);
and U26926 (N_26926,N_23302,N_18633);
and U26927 (N_26927,N_23786,N_23000);
nand U26928 (N_26928,N_22152,N_21875);
nand U26929 (N_26929,N_20877,N_19670);
or U26930 (N_26930,N_21617,N_20408);
nor U26931 (N_26931,N_22360,N_18310);
nor U26932 (N_26932,N_20130,N_21063);
xnor U26933 (N_26933,N_20788,N_18015);
xnor U26934 (N_26934,N_21318,N_20994);
or U26935 (N_26935,N_18415,N_18334);
nand U26936 (N_26936,N_18975,N_19299);
or U26937 (N_26937,N_19709,N_18381);
nand U26938 (N_26938,N_19494,N_21618);
xor U26939 (N_26939,N_18921,N_18583);
or U26940 (N_26940,N_21179,N_19323);
or U26941 (N_26941,N_20549,N_21972);
or U26942 (N_26942,N_20729,N_18489);
xor U26943 (N_26943,N_21811,N_20270);
or U26944 (N_26944,N_19394,N_23358);
nor U26945 (N_26945,N_20055,N_18546);
nor U26946 (N_26946,N_18322,N_23577);
nor U26947 (N_26947,N_21362,N_21738);
and U26948 (N_26948,N_23784,N_22448);
nor U26949 (N_26949,N_22290,N_23108);
or U26950 (N_26950,N_18265,N_23597);
nand U26951 (N_26951,N_21084,N_18504);
nand U26952 (N_26952,N_20232,N_21248);
xnor U26953 (N_26953,N_19489,N_22334);
xnor U26954 (N_26954,N_18682,N_22952);
and U26955 (N_26955,N_23269,N_20237);
or U26956 (N_26956,N_19998,N_20850);
and U26957 (N_26957,N_20743,N_20588);
nor U26958 (N_26958,N_22097,N_21060);
xnor U26959 (N_26959,N_23117,N_22063);
nor U26960 (N_26960,N_21078,N_19563);
xnor U26961 (N_26961,N_23573,N_20914);
xnor U26962 (N_26962,N_20247,N_18996);
or U26963 (N_26963,N_22478,N_21750);
and U26964 (N_26964,N_23199,N_18649);
or U26965 (N_26965,N_21404,N_20059);
or U26966 (N_26966,N_18752,N_22848);
nand U26967 (N_26967,N_19951,N_21917);
or U26968 (N_26968,N_20777,N_21319);
nor U26969 (N_26969,N_21734,N_18753);
or U26970 (N_26970,N_22086,N_19273);
nand U26971 (N_26971,N_21470,N_19234);
xor U26972 (N_26972,N_21061,N_19399);
or U26973 (N_26973,N_22535,N_19081);
and U26974 (N_26974,N_20793,N_21643);
or U26975 (N_26975,N_22219,N_19106);
nor U26976 (N_26976,N_18829,N_22846);
and U26977 (N_26977,N_23348,N_18638);
and U26978 (N_26978,N_23406,N_21460);
nor U26979 (N_26979,N_18879,N_22801);
and U26980 (N_26980,N_19324,N_18185);
nand U26981 (N_26981,N_22944,N_22687);
and U26982 (N_26982,N_19505,N_18833);
xor U26983 (N_26983,N_18932,N_23943);
xor U26984 (N_26984,N_18139,N_21779);
or U26985 (N_26985,N_18249,N_21592);
nor U26986 (N_26986,N_21161,N_19319);
nor U26987 (N_26987,N_19012,N_21436);
nand U26988 (N_26988,N_19098,N_18370);
and U26989 (N_26989,N_22181,N_22243);
and U26990 (N_26990,N_19253,N_23386);
xnor U26991 (N_26991,N_23189,N_20092);
or U26992 (N_26992,N_20949,N_22611);
nand U26993 (N_26993,N_20975,N_20838);
xnor U26994 (N_26994,N_21527,N_18862);
or U26995 (N_26995,N_20010,N_20730);
or U26996 (N_26996,N_20581,N_23385);
xnor U26997 (N_26997,N_23159,N_19983);
and U26998 (N_26998,N_23942,N_22596);
and U26999 (N_26999,N_19246,N_20086);
nand U27000 (N_27000,N_19323,N_20935);
xnor U27001 (N_27001,N_23559,N_18443);
nor U27002 (N_27002,N_21202,N_22569);
nand U27003 (N_27003,N_18607,N_22301);
and U27004 (N_27004,N_22961,N_20017);
xnor U27005 (N_27005,N_19695,N_23285);
and U27006 (N_27006,N_19836,N_21367);
and U27007 (N_27007,N_21769,N_19875);
or U27008 (N_27008,N_19591,N_22391);
xnor U27009 (N_27009,N_23205,N_19063);
or U27010 (N_27010,N_20717,N_23059);
and U27011 (N_27011,N_22426,N_20104);
nand U27012 (N_27012,N_21652,N_23981);
or U27013 (N_27013,N_23446,N_23489);
nand U27014 (N_27014,N_21873,N_20738);
nor U27015 (N_27015,N_21885,N_18545);
nor U27016 (N_27016,N_19309,N_19303);
or U27017 (N_27017,N_22968,N_21344);
and U27018 (N_27018,N_21548,N_22764);
nor U27019 (N_27019,N_21365,N_22671);
nand U27020 (N_27020,N_18042,N_23814);
xor U27021 (N_27021,N_22276,N_22987);
and U27022 (N_27022,N_22191,N_21279);
nor U27023 (N_27023,N_19432,N_19028);
and U27024 (N_27024,N_22342,N_19559);
xnor U27025 (N_27025,N_21878,N_23659);
xnor U27026 (N_27026,N_19209,N_19554);
or U27027 (N_27027,N_22261,N_22463);
nand U27028 (N_27028,N_23521,N_22253);
xnor U27029 (N_27029,N_20256,N_20189);
xor U27030 (N_27030,N_19712,N_19968);
and U27031 (N_27031,N_20572,N_18943);
xor U27032 (N_27032,N_22449,N_23735);
and U27033 (N_27033,N_22452,N_22636);
nor U27034 (N_27034,N_18808,N_18656);
or U27035 (N_27035,N_20763,N_21038);
or U27036 (N_27036,N_18568,N_22061);
nor U27037 (N_27037,N_20795,N_22902);
nor U27038 (N_27038,N_23650,N_18471);
nor U27039 (N_27039,N_20338,N_19678);
or U27040 (N_27040,N_22814,N_22741);
or U27041 (N_27041,N_20333,N_19547);
xnor U27042 (N_27042,N_19998,N_19553);
nand U27043 (N_27043,N_21076,N_19185);
or U27044 (N_27044,N_22968,N_22120);
or U27045 (N_27045,N_21748,N_21105);
nand U27046 (N_27046,N_18649,N_18185);
or U27047 (N_27047,N_18890,N_22162);
xor U27048 (N_27048,N_19436,N_21930);
nor U27049 (N_27049,N_20637,N_21754);
and U27050 (N_27050,N_21547,N_22794);
xnor U27051 (N_27051,N_19847,N_22732);
xor U27052 (N_27052,N_22893,N_18332);
and U27053 (N_27053,N_23196,N_21774);
or U27054 (N_27054,N_19274,N_18225);
nor U27055 (N_27055,N_18273,N_22195);
nor U27056 (N_27056,N_23709,N_23539);
nand U27057 (N_27057,N_21757,N_23470);
nand U27058 (N_27058,N_23921,N_20462);
xnor U27059 (N_27059,N_23477,N_20812);
or U27060 (N_27060,N_22667,N_21122);
nor U27061 (N_27061,N_19900,N_23939);
nand U27062 (N_27062,N_23260,N_23562);
and U27063 (N_27063,N_23913,N_20403);
nand U27064 (N_27064,N_22284,N_21607);
or U27065 (N_27065,N_20435,N_18590);
nor U27066 (N_27066,N_23493,N_22419);
nor U27067 (N_27067,N_19419,N_18627);
nand U27068 (N_27068,N_20221,N_21659);
nor U27069 (N_27069,N_23410,N_18820);
and U27070 (N_27070,N_22993,N_21060);
nor U27071 (N_27071,N_19756,N_23987);
xor U27072 (N_27072,N_20668,N_23479);
nor U27073 (N_27073,N_23131,N_18636);
xnor U27074 (N_27074,N_22507,N_22580);
and U27075 (N_27075,N_23979,N_21271);
or U27076 (N_27076,N_22234,N_18816);
xor U27077 (N_27077,N_22946,N_19151);
and U27078 (N_27078,N_23137,N_20359);
or U27079 (N_27079,N_19551,N_18634);
and U27080 (N_27080,N_18147,N_20663);
nand U27081 (N_27081,N_23062,N_23733);
xor U27082 (N_27082,N_21707,N_19095);
nand U27083 (N_27083,N_21253,N_19820);
xor U27084 (N_27084,N_18560,N_22294);
nor U27085 (N_27085,N_19354,N_20467);
and U27086 (N_27086,N_20572,N_20331);
xnor U27087 (N_27087,N_22391,N_18545);
nor U27088 (N_27088,N_21354,N_18958);
and U27089 (N_27089,N_20046,N_22127);
and U27090 (N_27090,N_21045,N_22823);
and U27091 (N_27091,N_21625,N_21478);
or U27092 (N_27092,N_21234,N_22598);
xor U27093 (N_27093,N_23710,N_23686);
nor U27094 (N_27094,N_23393,N_21867);
or U27095 (N_27095,N_18882,N_23504);
nand U27096 (N_27096,N_19102,N_22718);
or U27097 (N_27097,N_18619,N_18767);
or U27098 (N_27098,N_20571,N_23047);
or U27099 (N_27099,N_20821,N_23365);
nor U27100 (N_27100,N_22474,N_21691);
nand U27101 (N_27101,N_23250,N_18497);
xnor U27102 (N_27102,N_19279,N_20897);
nor U27103 (N_27103,N_21752,N_23804);
nor U27104 (N_27104,N_18414,N_18372);
or U27105 (N_27105,N_18794,N_19368);
and U27106 (N_27106,N_23443,N_21984);
and U27107 (N_27107,N_22104,N_21219);
or U27108 (N_27108,N_18389,N_21279);
and U27109 (N_27109,N_21579,N_18840);
nor U27110 (N_27110,N_22711,N_23120);
or U27111 (N_27111,N_18435,N_18669);
and U27112 (N_27112,N_18053,N_19722);
nand U27113 (N_27113,N_23161,N_18284);
nand U27114 (N_27114,N_19547,N_21459);
nor U27115 (N_27115,N_21930,N_19068);
xor U27116 (N_27116,N_20394,N_22818);
or U27117 (N_27117,N_19375,N_23041);
or U27118 (N_27118,N_20712,N_21918);
nor U27119 (N_27119,N_22709,N_20160);
and U27120 (N_27120,N_20550,N_21769);
xnor U27121 (N_27121,N_21333,N_20158);
xnor U27122 (N_27122,N_18604,N_22795);
xor U27123 (N_27123,N_23345,N_19397);
xnor U27124 (N_27124,N_22716,N_23277);
nor U27125 (N_27125,N_20887,N_22397);
nand U27126 (N_27126,N_21065,N_20644);
nor U27127 (N_27127,N_20070,N_19252);
xor U27128 (N_27128,N_21742,N_22197);
nand U27129 (N_27129,N_20179,N_20026);
nand U27130 (N_27130,N_21861,N_20669);
and U27131 (N_27131,N_18351,N_21106);
nand U27132 (N_27132,N_18950,N_19963);
xnor U27133 (N_27133,N_23224,N_18638);
or U27134 (N_27134,N_23828,N_21339);
and U27135 (N_27135,N_22446,N_21525);
or U27136 (N_27136,N_20588,N_21124);
or U27137 (N_27137,N_19771,N_23412);
or U27138 (N_27138,N_21466,N_23316);
xor U27139 (N_27139,N_23693,N_18550);
xnor U27140 (N_27140,N_18241,N_21560);
or U27141 (N_27141,N_19692,N_23663);
xor U27142 (N_27142,N_21025,N_19640);
xnor U27143 (N_27143,N_21779,N_23501);
xor U27144 (N_27144,N_23259,N_20648);
and U27145 (N_27145,N_21447,N_20209);
or U27146 (N_27146,N_19243,N_19789);
nor U27147 (N_27147,N_22527,N_22956);
nand U27148 (N_27148,N_19166,N_20876);
xor U27149 (N_27149,N_22732,N_19579);
nand U27150 (N_27150,N_22064,N_20159);
xnor U27151 (N_27151,N_23479,N_22369);
nor U27152 (N_27152,N_23200,N_23842);
nor U27153 (N_27153,N_22761,N_22604);
or U27154 (N_27154,N_20619,N_19719);
xnor U27155 (N_27155,N_21749,N_19456);
and U27156 (N_27156,N_20157,N_18553);
nor U27157 (N_27157,N_20202,N_22162);
or U27158 (N_27158,N_21941,N_20096);
or U27159 (N_27159,N_20988,N_19422);
nand U27160 (N_27160,N_18847,N_23202);
xor U27161 (N_27161,N_23885,N_21753);
or U27162 (N_27162,N_18791,N_21120);
and U27163 (N_27163,N_22326,N_22251);
and U27164 (N_27164,N_23939,N_20402);
and U27165 (N_27165,N_22079,N_18219);
xnor U27166 (N_27166,N_21382,N_23479);
nand U27167 (N_27167,N_18539,N_23474);
and U27168 (N_27168,N_22328,N_19475);
or U27169 (N_27169,N_20605,N_23053);
nor U27170 (N_27170,N_21252,N_21311);
nor U27171 (N_27171,N_23630,N_18624);
nand U27172 (N_27172,N_23552,N_23336);
xor U27173 (N_27173,N_20506,N_19134);
or U27174 (N_27174,N_18985,N_18990);
nand U27175 (N_27175,N_21669,N_23161);
and U27176 (N_27176,N_20101,N_18626);
and U27177 (N_27177,N_19873,N_21345);
or U27178 (N_27178,N_21191,N_19969);
xor U27179 (N_27179,N_20011,N_18368);
xnor U27180 (N_27180,N_23368,N_21745);
xnor U27181 (N_27181,N_18184,N_22713);
or U27182 (N_27182,N_21414,N_22489);
or U27183 (N_27183,N_21799,N_19519);
nor U27184 (N_27184,N_19470,N_20753);
or U27185 (N_27185,N_23957,N_21927);
nand U27186 (N_27186,N_22739,N_22814);
and U27187 (N_27187,N_22555,N_19606);
and U27188 (N_27188,N_23084,N_21736);
nor U27189 (N_27189,N_18659,N_18688);
or U27190 (N_27190,N_20138,N_21128);
nor U27191 (N_27191,N_23484,N_21467);
nand U27192 (N_27192,N_18751,N_20380);
and U27193 (N_27193,N_21982,N_21033);
nand U27194 (N_27194,N_19742,N_23612);
and U27195 (N_27195,N_23029,N_18265);
and U27196 (N_27196,N_23911,N_21129);
xnor U27197 (N_27197,N_19308,N_21800);
or U27198 (N_27198,N_23503,N_23751);
nor U27199 (N_27199,N_23921,N_19072);
nor U27200 (N_27200,N_23063,N_20248);
or U27201 (N_27201,N_22528,N_23948);
nor U27202 (N_27202,N_19442,N_21616);
nor U27203 (N_27203,N_19345,N_23528);
and U27204 (N_27204,N_23553,N_22483);
or U27205 (N_27205,N_21325,N_19975);
and U27206 (N_27206,N_20577,N_18908);
and U27207 (N_27207,N_20442,N_19300);
xor U27208 (N_27208,N_18484,N_19334);
xor U27209 (N_27209,N_21241,N_23258);
nand U27210 (N_27210,N_18522,N_18528);
xor U27211 (N_27211,N_20848,N_23998);
or U27212 (N_27212,N_19909,N_23274);
nand U27213 (N_27213,N_23881,N_21706);
nor U27214 (N_27214,N_22342,N_22092);
and U27215 (N_27215,N_20698,N_21873);
nand U27216 (N_27216,N_18022,N_23134);
nor U27217 (N_27217,N_18941,N_20437);
xnor U27218 (N_27218,N_22950,N_23978);
or U27219 (N_27219,N_21116,N_21233);
and U27220 (N_27220,N_18838,N_18124);
nor U27221 (N_27221,N_23353,N_20738);
nand U27222 (N_27222,N_19802,N_22154);
and U27223 (N_27223,N_23440,N_21675);
xnor U27224 (N_27224,N_19351,N_18406);
or U27225 (N_27225,N_18951,N_20720);
nand U27226 (N_27226,N_21551,N_18174);
nor U27227 (N_27227,N_20505,N_19858);
nor U27228 (N_27228,N_19200,N_18056);
nor U27229 (N_27229,N_22960,N_18899);
or U27230 (N_27230,N_18100,N_20818);
xor U27231 (N_27231,N_22101,N_19324);
nand U27232 (N_27232,N_21181,N_19356);
nor U27233 (N_27233,N_23637,N_22036);
and U27234 (N_27234,N_21109,N_18951);
nor U27235 (N_27235,N_20365,N_18490);
and U27236 (N_27236,N_18731,N_22018);
nor U27237 (N_27237,N_18420,N_19473);
nor U27238 (N_27238,N_18810,N_22550);
nand U27239 (N_27239,N_19439,N_22689);
nor U27240 (N_27240,N_22683,N_22545);
or U27241 (N_27241,N_18501,N_18624);
or U27242 (N_27242,N_22350,N_19786);
nor U27243 (N_27243,N_19765,N_21615);
or U27244 (N_27244,N_20624,N_18762);
and U27245 (N_27245,N_19060,N_23752);
and U27246 (N_27246,N_21421,N_20587);
nand U27247 (N_27247,N_22199,N_21705);
nor U27248 (N_27248,N_18534,N_18582);
nor U27249 (N_27249,N_23526,N_18979);
nor U27250 (N_27250,N_23152,N_23981);
and U27251 (N_27251,N_23205,N_22399);
nand U27252 (N_27252,N_18837,N_23399);
xor U27253 (N_27253,N_22446,N_21637);
xor U27254 (N_27254,N_22654,N_23923);
nor U27255 (N_27255,N_19975,N_20649);
and U27256 (N_27256,N_22542,N_18608);
or U27257 (N_27257,N_20114,N_19209);
nand U27258 (N_27258,N_18787,N_22587);
nor U27259 (N_27259,N_22146,N_23896);
or U27260 (N_27260,N_19558,N_20541);
and U27261 (N_27261,N_22332,N_18206);
nand U27262 (N_27262,N_20002,N_23379);
nor U27263 (N_27263,N_18680,N_22421);
xor U27264 (N_27264,N_21120,N_21247);
xor U27265 (N_27265,N_21924,N_20978);
or U27266 (N_27266,N_20782,N_23639);
nor U27267 (N_27267,N_18100,N_18283);
nor U27268 (N_27268,N_21236,N_18841);
and U27269 (N_27269,N_23717,N_20150);
and U27270 (N_27270,N_20565,N_18830);
xor U27271 (N_27271,N_21749,N_19603);
nand U27272 (N_27272,N_21453,N_20556);
nor U27273 (N_27273,N_20728,N_18826);
xor U27274 (N_27274,N_21930,N_18492);
and U27275 (N_27275,N_20494,N_20521);
or U27276 (N_27276,N_21637,N_20471);
nand U27277 (N_27277,N_23256,N_22822);
and U27278 (N_27278,N_19539,N_22789);
or U27279 (N_27279,N_23239,N_18338);
or U27280 (N_27280,N_22963,N_19405);
nor U27281 (N_27281,N_23680,N_22231);
nor U27282 (N_27282,N_21442,N_18556);
xor U27283 (N_27283,N_22088,N_20522);
xnor U27284 (N_27284,N_22552,N_20228);
or U27285 (N_27285,N_20959,N_21137);
nand U27286 (N_27286,N_20532,N_23800);
nand U27287 (N_27287,N_18952,N_18141);
or U27288 (N_27288,N_21350,N_22410);
or U27289 (N_27289,N_19895,N_23746);
nor U27290 (N_27290,N_19377,N_19889);
xnor U27291 (N_27291,N_20790,N_21691);
nand U27292 (N_27292,N_22361,N_22904);
xor U27293 (N_27293,N_18858,N_23562);
xor U27294 (N_27294,N_19275,N_19967);
nor U27295 (N_27295,N_18302,N_18632);
xnor U27296 (N_27296,N_21415,N_21492);
nand U27297 (N_27297,N_23080,N_18102);
xnor U27298 (N_27298,N_21929,N_20660);
or U27299 (N_27299,N_19670,N_19466);
nand U27300 (N_27300,N_23546,N_22136);
nand U27301 (N_27301,N_23488,N_22973);
nand U27302 (N_27302,N_20204,N_22357);
xnor U27303 (N_27303,N_19052,N_19814);
or U27304 (N_27304,N_23781,N_18064);
or U27305 (N_27305,N_21957,N_19997);
nand U27306 (N_27306,N_18610,N_23014);
nand U27307 (N_27307,N_20493,N_19057);
and U27308 (N_27308,N_19676,N_18142);
and U27309 (N_27309,N_21366,N_19962);
nand U27310 (N_27310,N_22626,N_21909);
nand U27311 (N_27311,N_23317,N_18098);
nand U27312 (N_27312,N_19174,N_18248);
and U27313 (N_27313,N_18640,N_19126);
nor U27314 (N_27314,N_21162,N_20840);
nand U27315 (N_27315,N_22249,N_19339);
and U27316 (N_27316,N_21959,N_18220);
or U27317 (N_27317,N_22261,N_21042);
and U27318 (N_27318,N_19185,N_19078);
nor U27319 (N_27319,N_23064,N_23394);
xnor U27320 (N_27320,N_18987,N_19166);
or U27321 (N_27321,N_18551,N_21684);
and U27322 (N_27322,N_18183,N_19571);
xnor U27323 (N_27323,N_21336,N_18006);
xor U27324 (N_27324,N_23627,N_21969);
xor U27325 (N_27325,N_19098,N_23326);
or U27326 (N_27326,N_23077,N_21551);
xor U27327 (N_27327,N_21929,N_19928);
nor U27328 (N_27328,N_23473,N_23798);
and U27329 (N_27329,N_21396,N_18738);
nand U27330 (N_27330,N_22678,N_19441);
nand U27331 (N_27331,N_21328,N_20236);
nand U27332 (N_27332,N_23647,N_20462);
and U27333 (N_27333,N_21210,N_19442);
and U27334 (N_27334,N_23862,N_19677);
xor U27335 (N_27335,N_19228,N_19137);
nor U27336 (N_27336,N_22617,N_18308);
xor U27337 (N_27337,N_21326,N_23439);
nor U27338 (N_27338,N_22306,N_21822);
xnor U27339 (N_27339,N_20605,N_20538);
xor U27340 (N_27340,N_19715,N_22925);
xnor U27341 (N_27341,N_23447,N_20768);
and U27342 (N_27342,N_23010,N_22637);
and U27343 (N_27343,N_18695,N_18060);
nand U27344 (N_27344,N_20323,N_22801);
or U27345 (N_27345,N_19529,N_23226);
xor U27346 (N_27346,N_20707,N_21752);
or U27347 (N_27347,N_23067,N_22506);
or U27348 (N_27348,N_23156,N_20351);
xnor U27349 (N_27349,N_23861,N_22173);
and U27350 (N_27350,N_20607,N_19755);
nor U27351 (N_27351,N_21300,N_19000);
nor U27352 (N_27352,N_23518,N_18439);
xor U27353 (N_27353,N_22652,N_18255);
nand U27354 (N_27354,N_21537,N_18839);
nor U27355 (N_27355,N_23916,N_18743);
and U27356 (N_27356,N_23948,N_19006);
nor U27357 (N_27357,N_22863,N_21954);
xor U27358 (N_27358,N_19473,N_19356);
xor U27359 (N_27359,N_19460,N_19172);
and U27360 (N_27360,N_23008,N_21630);
xnor U27361 (N_27361,N_19516,N_23381);
and U27362 (N_27362,N_21231,N_19250);
nand U27363 (N_27363,N_20968,N_19916);
and U27364 (N_27364,N_22835,N_21123);
or U27365 (N_27365,N_22542,N_19819);
xnor U27366 (N_27366,N_18846,N_23237);
or U27367 (N_27367,N_20397,N_21424);
or U27368 (N_27368,N_21893,N_19648);
xnor U27369 (N_27369,N_20195,N_22346);
xnor U27370 (N_27370,N_22572,N_21925);
or U27371 (N_27371,N_18504,N_20327);
nor U27372 (N_27372,N_20779,N_21891);
xnor U27373 (N_27373,N_22805,N_18671);
xor U27374 (N_27374,N_22573,N_21476);
and U27375 (N_27375,N_23609,N_20281);
nand U27376 (N_27376,N_19178,N_21180);
or U27377 (N_27377,N_23845,N_23038);
or U27378 (N_27378,N_23632,N_18020);
xor U27379 (N_27379,N_19889,N_23607);
nand U27380 (N_27380,N_18961,N_18351);
xnor U27381 (N_27381,N_18298,N_22090);
nand U27382 (N_27382,N_21093,N_18301);
nand U27383 (N_27383,N_22188,N_20466);
or U27384 (N_27384,N_20663,N_19720);
xor U27385 (N_27385,N_18024,N_21247);
nor U27386 (N_27386,N_23684,N_18791);
nor U27387 (N_27387,N_18471,N_20668);
nand U27388 (N_27388,N_21915,N_20273);
nor U27389 (N_27389,N_21151,N_18926);
xnor U27390 (N_27390,N_19081,N_18127);
and U27391 (N_27391,N_19630,N_18610);
xor U27392 (N_27392,N_21766,N_22600);
xor U27393 (N_27393,N_18710,N_21673);
or U27394 (N_27394,N_22119,N_23597);
and U27395 (N_27395,N_20502,N_20613);
nor U27396 (N_27396,N_21672,N_22677);
xnor U27397 (N_27397,N_18688,N_20283);
xor U27398 (N_27398,N_22362,N_19078);
and U27399 (N_27399,N_20701,N_20552);
nor U27400 (N_27400,N_19099,N_19710);
nor U27401 (N_27401,N_23888,N_23282);
and U27402 (N_27402,N_18278,N_19467);
and U27403 (N_27403,N_19840,N_23608);
xnor U27404 (N_27404,N_20426,N_18896);
or U27405 (N_27405,N_22119,N_18985);
or U27406 (N_27406,N_18990,N_22486);
and U27407 (N_27407,N_23197,N_20180);
or U27408 (N_27408,N_23026,N_23132);
nand U27409 (N_27409,N_21398,N_21250);
and U27410 (N_27410,N_20667,N_23816);
and U27411 (N_27411,N_22272,N_23450);
xor U27412 (N_27412,N_18749,N_22727);
xor U27413 (N_27413,N_20476,N_22337);
nor U27414 (N_27414,N_19827,N_22773);
or U27415 (N_27415,N_23566,N_23784);
or U27416 (N_27416,N_19223,N_18772);
or U27417 (N_27417,N_20823,N_18184);
nor U27418 (N_27418,N_22250,N_22761);
nand U27419 (N_27419,N_21801,N_21982);
xnor U27420 (N_27420,N_21359,N_20462);
xnor U27421 (N_27421,N_20602,N_21537);
nor U27422 (N_27422,N_19683,N_22065);
and U27423 (N_27423,N_21977,N_22274);
nand U27424 (N_27424,N_19037,N_19159);
or U27425 (N_27425,N_23384,N_19191);
xor U27426 (N_27426,N_21711,N_18582);
nand U27427 (N_27427,N_19165,N_21769);
or U27428 (N_27428,N_22930,N_18228);
nor U27429 (N_27429,N_23846,N_22400);
xor U27430 (N_27430,N_21185,N_19007);
xnor U27431 (N_27431,N_20973,N_23028);
nand U27432 (N_27432,N_21454,N_20679);
or U27433 (N_27433,N_18897,N_20413);
and U27434 (N_27434,N_20812,N_21025);
xor U27435 (N_27435,N_23499,N_23352);
or U27436 (N_27436,N_19327,N_22442);
xnor U27437 (N_27437,N_19781,N_19066);
and U27438 (N_27438,N_19186,N_23998);
and U27439 (N_27439,N_20447,N_18386);
nor U27440 (N_27440,N_20598,N_19240);
nand U27441 (N_27441,N_20844,N_22457);
and U27442 (N_27442,N_20313,N_21217);
nand U27443 (N_27443,N_19511,N_23136);
nor U27444 (N_27444,N_19968,N_18612);
and U27445 (N_27445,N_23274,N_19444);
nand U27446 (N_27446,N_20183,N_19389);
nand U27447 (N_27447,N_18169,N_21195);
and U27448 (N_27448,N_19814,N_21847);
xor U27449 (N_27449,N_20838,N_18312);
or U27450 (N_27450,N_21035,N_18191);
xnor U27451 (N_27451,N_18494,N_18656);
xnor U27452 (N_27452,N_19873,N_20711);
and U27453 (N_27453,N_18638,N_23376);
nor U27454 (N_27454,N_18998,N_21748);
nand U27455 (N_27455,N_20253,N_21700);
nor U27456 (N_27456,N_21086,N_21063);
and U27457 (N_27457,N_21150,N_23740);
xnor U27458 (N_27458,N_21009,N_22491);
nor U27459 (N_27459,N_21737,N_21478);
or U27460 (N_27460,N_23440,N_20969);
xor U27461 (N_27461,N_19705,N_18486);
xor U27462 (N_27462,N_19952,N_18096);
nor U27463 (N_27463,N_22393,N_22285);
nand U27464 (N_27464,N_18931,N_22528);
or U27465 (N_27465,N_19305,N_22911);
nor U27466 (N_27466,N_19237,N_20803);
or U27467 (N_27467,N_18992,N_19518);
or U27468 (N_27468,N_18400,N_19677);
or U27469 (N_27469,N_22085,N_22884);
nand U27470 (N_27470,N_22702,N_21444);
xnor U27471 (N_27471,N_18769,N_18881);
or U27472 (N_27472,N_18087,N_23166);
nor U27473 (N_27473,N_18263,N_23167);
and U27474 (N_27474,N_23341,N_21946);
xor U27475 (N_27475,N_23170,N_21218);
nand U27476 (N_27476,N_18944,N_20267);
or U27477 (N_27477,N_20700,N_19022);
xnor U27478 (N_27478,N_19014,N_22045);
and U27479 (N_27479,N_18901,N_23895);
nand U27480 (N_27480,N_23866,N_20490);
or U27481 (N_27481,N_18346,N_21817);
or U27482 (N_27482,N_18446,N_22466);
and U27483 (N_27483,N_21405,N_19543);
or U27484 (N_27484,N_23702,N_22722);
nand U27485 (N_27485,N_19746,N_18197);
and U27486 (N_27486,N_19992,N_18662);
or U27487 (N_27487,N_22406,N_18315);
and U27488 (N_27488,N_22534,N_20646);
xor U27489 (N_27489,N_22426,N_21866);
xor U27490 (N_27490,N_20459,N_19918);
nand U27491 (N_27491,N_20442,N_18611);
and U27492 (N_27492,N_20319,N_18250);
or U27493 (N_27493,N_18259,N_21138);
nor U27494 (N_27494,N_23286,N_23258);
and U27495 (N_27495,N_19225,N_22335);
nand U27496 (N_27496,N_18003,N_19933);
nor U27497 (N_27497,N_20199,N_19216);
and U27498 (N_27498,N_19784,N_21865);
or U27499 (N_27499,N_22528,N_19862);
xor U27500 (N_27500,N_18159,N_18635);
nand U27501 (N_27501,N_18489,N_18867);
nor U27502 (N_27502,N_18935,N_22026);
and U27503 (N_27503,N_21659,N_18888);
nor U27504 (N_27504,N_19811,N_21037);
nor U27505 (N_27505,N_21067,N_21787);
or U27506 (N_27506,N_20231,N_18135);
or U27507 (N_27507,N_22803,N_23088);
or U27508 (N_27508,N_23401,N_19417);
nor U27509 (N_27509,N_23076,N_19041);
nand U27510 (N_27510,N_20398,N_19728);
nor U27511 (N_27511,N_19611,N_20506);
nor U27512 (N_27512,N_23752,N_22200);
and U27513 (N_27513,N_23499,N_22618);
nand U27514 (N_27514,N_20094,N_20642);
or U27515 (N_27515,N_22239,N_21201);
or U27516 (N_27516,N_22502,N_18222);
and U27517 (N_27517,N_19715,N_19962);
nor U27518 (N_27518,N_18771,N_23055);
and U27519 (N_27519,N_22196,N_20638);
or U27520 (N_27520,N_19475,N_21034);
or U27521 (N_27521,N_21178,N_23786);
xor U27522 (N_27522,N_19043,N_20181);
xnor U27523 (N_27523,N_21997,N_23081);
or U27524 (N_27524,N_22119,N_19563);
and U27525 (N_27525,N_21899,N_23962);
or U27526 (N_27526,N_19441,N_22686);
nand U27527 (N_27527,N_22231,N_22648);
xor U27528 (N_27528,N_22414,N_18040);
or U27529 (N_27529,N_22475,N_20882);
xor U27530 (N_27530,N_19276,N_22205);
nor U27531 (N_27531,N_23248,N_21321);
xor U27532 (N_27532,N_20875,N_19511);
xnor U27533 (N_27533,N_22036,N_22105);
or U27534 (N_27534,N_20116,N_18867);
nand U27535 (N_27535,N_22610,N_22292);
nor U27536 (N_27536,N_21124,N_21516);
or U27537 (N_27537,N_21614,N_22056);
nand U27538 (N_27538,N_21036,N_20647);
xnor U27539 (N_27539,N_18912,N_23140);
and U27540 (N_27540,N_18116,N_20038);
and U27541 (N_27541,N_19813,N_20876);
nor U27542 (N_27542,N_20298,N_22490);
xnor U27543 (N_27543,N_18070,N_18927);
nor U27544 (N_27544,N_23506,N_22103);
or U27545 (N_27545,N_20125,N_18967);
nor U27546 (N_27546,N_20415,N_19114);
nor U27547 (N_27547,N_22234,N_18388);
xnor U27548 (N_27548,N_21953,N_19160);
xnor U27549 (N_27549,N_21050,N_23838);
or U27550 (N_27550,N_23136,N_22784);
xor U27551 (N_27551,N_20538,N_21514);
nand U27552 (N_27552,N_21232,N_23780);
nand U27553 (N_27553,N_23844,N_23876);
and U27554 (N_27554,N_19140,N_23117);
nand U27555 (N_27555,N_18755,N_22931);
xor U27556 (N_27556,N_19570,N_21104);
xor U27557 (N_27557,N_20529,N_20675);
and U27558 (N_27558,N_18606,N_19925);
nor U27559 (N_27559,N_18653,N_20916);
xor U27560 (N_27560,N_19143,N_21186);
and U27561 (N_27561,N_22610,N_19863);
nor U27562 (N_27562,N_20393,N_18338);
xor U27563 (N_27563,N_22235,N_23017);
xnor U27564 (N_27564,N_22534,N_19250);
and U27565 (N_27565,N_22523,N_20248);
and U27566 (N_27566,N_21686,N_22286);
and U27567 (N_27567,N_21771,N_21989);
and U27568 (N_27568,N_22493,N_22061);
nor U27569 (N_27569,N_20441,N_20262);
or U27570 (N_27570,N_18732,N_19334);
and U27571 (N_27571,N_23330,N_22702);
nand U27572 (N_27572,N_23392,N_22393);
nor U27573 (N_27573,N_20671,N_21192);
nor U27574 (N_27574,N_19459,N_20494);
nor U27575 (N_27575,N_18707,N_21299);
nor U27576 (N_27576,N_18729,N_21955);
nand U27577 (N_27577,N_23454,N_18235);
nand U27578 (N_27578,N_19336,N_18366);
xnor U27579 (N_27579,N_19087,N_19170);
xnor U27580 (N_27580,N_23195,N_19805);
xnor U27581 (N_27581,N_20744,N_23651);
nor U27582 (N_27582,N_18693,N_21699);
nand U27583 (N_27583,N_19929,N_22704);
and U27584 (N_27584,N_18993,N_19711);
or U27585 (N_27585,N_19383,N_23250);
or U27586 (N_27586,N_19496,N_22920);
or U27587 (N_27587,N_18099,N_23596);
and U27588 (N_27588,N_20834,N_23154);
nand U27589 (N_27589,N_21507,N_18859);
and U27590 (N_27590,N_23979,N_19217);
nor U27591 (N_27591,N_18470,N_20214);
nor U27592 (N_27592,N_18569,N_18688);
and U27593 (N_27593,N_21694,N_21716);
and U27594 (N_27594,N_22769,N_18014);
nand U27595 (N_27595,N_22301,N_19747);
and U27596 (N_27596,N_22443,N_18382);
or U27597 (N_27597,N_18374,N_22336);
xor U27598 (N_27598,N_18300,N_23311);
xnor U27599 (N_27599,N_19042,N_18970);
xor U27600 (N_27600,N_18676,N_18664);
nor U27601 (N_27601,N_21492,N_22629);
or U27602 (N_27602,N_20146,N_23245);
nand U27603 (N_27603,N_21813,N_23751);
xor U27604 (N_27604,N_21732,N_20566);
xnor U27605 (N_27605,N_21867,N_18084);
xor U27606 (N_27606,N_19690,N_22160);
or U27607 (N_27607,N_21024,N_21047);
nor U27608 (N_27608,N_22563,N_22117);
nor U27609 (N_27609,N_19729,N_22824);
nand U27610 (N_27610,N_18814,N_18816);
and U27611 (N_27611,N_22927,N_22476);
nand U27612 (N_27612,N_21628,N_20083);
or U27613 (N_27613,N_22737,N_18892);
nand U27614 (N_27614,N_20959,N_22777);
or U27615 (N_27615,N_19827,N_23930);
xnor U27616 (N_27616,N_18716,N_19684);
or U27617 (N_27617,N_21667,N_21024);
and U27618 (N_27618,N_20707,N_19307);
nor U27619 (N_27619,N_19944,N_22899);
and U27620 (N_27620,N_20423,N_23734);
nor U27621 (N_27621,N_20014,N_20501);
nor U27622 (N_27622,N_19744,N_22043);
xor U27623 (N_27623,N_19878,N_22631);
xor U27624 (N_27624,N_20609,N_19827);
nor U27625 (N_27625,N_20052,N_22627);
and U27626 (N_27626,N_23551,N_23642);
nand U27627 (N_27627,N_19677,N_18802);
xnor U27628 (N_27628,N_22528,N_22485);
nor U27629 (N_27629,N_19158,N_21145);
or U27630 (N_27630,N_19244,N_18482);
nand U27631 (N_27631,N_21493,N_19515);
or U27632 (N_27632,N_22852,N_23330);
or U27633 (N_27633,N_18205,N_22783);
nor U27634 (N_27634,N_23011,N_23937);
nor U27635 (N_27635,N_19794,N_21850);
nand U27636 (N_27636,N_19409,N_22513);
xor U27637 (N_27637,N_23112,N_23913);
and U27638 (N_27638,N_20459,N_20331);
nand U27639 (N_27639,N_22750,N_20490);
xnor U27640 (N_27640,N_19962,N_18956);
nor U27641 (N_27641,N_22231,N_23205);
or U27642 (N_27642,N_22394,N_18171);
nor U27643 (N_27643,N_20256,N_18297);
or U27644 (N_27644,N_19839,N_19943);
and U27645 (N_27645,N_20763,N_23270);
xor U27646 (N_27646,N_21573,N_18764);
and U27647 (N_27647,N_22921,N_18681);
xnor U27648 (N_27648,N_23816,N_21779);
nand U27649 (N_27649,N_23069,N_21242);
and U27650 (N_27650,N_23694,N_22506);
or U27651 (N_27651,N_21012,N_21347);
or U27652 (N_27652,N_18241,N_18703);
xnor U27653 (N_27653,N_22794,N_23459);
and U27654 (N_27654,N_19268,N_20041);
nor U27655 (N_27655,N_22879,N_21736);
xor U27656 (N_27656,N_18318,N_21232);
nor U27657 (N_27657,N_20766,N_21479);
and U27658 (N_27658,N_22597,N_21534);
and U27659 (N_27659,N_23446,N_22458);
and U27660 (N_27660,N_21181,N_19442);
xor U27661 (N_27661,N_21607,N_20910);
nor U27662 (N_27662,N_21235,N_22516);
xor U27663 (N_27663,N_23629,N_19384);
or U27664 (N_27664,N_22419,N_18580);
or U27665 (N_27665,N_21832,N_18971);
and U27666 (N_27666,N_20988,N_18435);
nand U27667 (N_27667,N_21695,N_19809);
and U27668 (N_27668,N_23266,N_21728);
nand U27669 (N_27669,N_20506,N_20020);
and U27670 (N_27670,N_19969,N_18073);
or U27671 (N_27671,N_19589,N_20615);
nor U27672 (N_27672,N_21438,N_19197);
and U27673 (N_27673,N_23024,N_22680);
or U27674 (N_27674,N_20593,N_21904);
nor U27675 (N_27675,N_20543,N_23865);
or U27676 (N_27676,N_23038,N_19315);
nand U27677 (N_27677,N_23859,N_18490);
or U27678 (N_27678,N_21723,N_22668);
and U27679 (N_27679,N_20468,N_20714);
xnor U27680 (N_27680,N_20354,N_21105);
nor U27681 (N_27681,N_21637,N_21998);
nand U27682 (N_27682,N_22855,N_20559);
xnor U27683 (N_27683,N_18278,N_21853);
xor U27684 (N_27684,N_23790,N_19713);
or U27685 (N_27685,N_19930,N_23733);
nor U27686 (N_27686,N_20520,N_23725);
nand U27687 (N_27687,N_22774,N_21682);
and U27688 (N_27688,N_19250,N_19300);
nor U27689 (N_27689,N_23132,N_20757);
xor U27690 (N_27690,N_22842,N_23525);
or U27691 (N_27691,N_23454,N_19140);
nor U27692 (N_27692,N_22156,N_18964);
nor U27693 (N_27693,N_21003,N_18104);
or U27694 (N_27694,N_22427,N_22936);
xnor U27695 (N_27695,N_18398,N_23695);
xor U27696 (N_27696,N_21228,N_23151);
or U27697 (N_27697,N_18088,N_23219);
nand U27698 (N_27698,N_22252,N_22587);
and U27699 (N_27699,N_21657,N_22079);
xnor U27700 (N_27700,N_19157,N_23596);
xor U27701 (N_27701,N_19202,N_22492);
nand U27702 (N_27702,N_21855,N_19908);
nor U27703 (N_27703,N_20361,N_18156);
nor U27704 (N_27704,N_20551,N_22925);
nand U27705 (N_27705,N_18470,N_19524);
nand U27706 (N_27706,N_18986,N_18980);
nor U27707 (N_27707,N_22484,N_18207);
or U27708 (N_27708,N_19465,N_23384);
nand U27709 (N_27709,N_20960,N_21081);
nor U27710 (N_27710,N_19848,N_19537);
xnor U27711 (N_27711,N_23271,N_22188);
or U27712 (N_27712,N_19043,N_18190);
nor U27713 (N_27713,N_22144,N_20555);
nand U27714 (N_27714,N_23968,N_20506);
or U27715 (N_27715,N_19973,N_19902);
nand U27716 (N_27716,N_20509,N_21782);
nor U27717 (N_27717,N_22011,N_23452);
and U27718 (N_27718,N_23051,N_19536);
nand U27719 (N_27719,N_18479,N_23189);
and U27720 (N_27720,N_23547,N_22925);
nand U27721 (N_27721,N_19047,N_23964);
nor U27722 (N_27722,N_22899,N_20199);
nand U27723 (N_27723,N_20851,N_23545);
nand U27724 (N_27724,N_18899,N_18877);
or U27725 (N_27725,N_21291,N_18085);
xnor U27726 (N_27726,N_19010,N_21833);
or U27727 (N_27727,N_19000,N_19128);
and U27728 (N_27728,N_22840,N_19755);
or U27729 (N_27729,N_20044,N_21726);
xnor U27730 (N_27730,N_19259,N_19918);
and U27731 (N_27731,N_22693,N_21274);
xnor U27732 (N_27732,N_23653,N_22469);
xor U27733 (N_27733,N_23033,N_23161);
xor U27734 (N_27734,N_23399,N_22257);
or U27735 (N_27735,N_21913,N_19923);
nand U27736 (N_27736,N_22230,N_22988);
nor U27737 (N_27737,N_20064,N_23521);
and U27738 (N_27738,N_22675,N_21675);
xnor U27739 (N_27739,N_21062,N_18788);
nor U27740 (N_27740,N_23018,N_22666);
and U27741 (N_27741,N_20706,N_21014);
nand U27742 (N_27742,N_22620,N_18129);
nand U27743 (N_27743,N_20261,N_21938);
nand U27744 (N_27744,N_18427,N_23065);
xnor U27745 (N_27745,N_21464,N_19701);
nor U27746 (N_27746,N_19515,N_21628);
or U27747 (N_27747,N_18320,N_18540);
or U27748 (N_27748,N_20690,N_18196);
or U27749 (N_27749,N_19417,N_20544);
nand U27750 (N_27750,N_20111,N_21327);
xnor U27751 (N_27751,N_21177,N_20628);
nor U27752 (N_27752,N_21968,N_23393);
or U27753 (N_27753,N_21112,N_19920);
xor U27754 (N_27754,N_18170,N_23350);
and U27755 (N_27755,N_19006,N_18520);
nand U27756 (N_27756,N_20926,N_23656);
nor U27757 (N_27757,N_21612,N_18236);
nor U27758 (N_27758,N_21742,N_21853);
and U27759 (N_27759,N_23953,N_20937);
xnor U27760 (N_27760,N_18156,N_20690);
nand U27761 (N_27761,N_23228,N_22511);
nand U27762 (N_27762,N_19341,N_22941);
nor U27763 (N_27763,N_19509,N_20755);
or U27764 (N_27764,N_18322,N_18307);
nand U27765 (N_27765,N_21860,N_18057);
and U27766 (N_27766,N_20020,N_18857);
nand U27767 (N_27767,N_23502,N_20153);
and U27768 (N_27768,N_21476,N_21092);
and U27769 (N_27769,N_20687,N_22701);
or U27770 (N_27770,N_22420,N_18294);
xor U27771 (N_27771,N_22294,N_19467);
nor U27772 (N_27772,N_22246,N_21083);
xor U27773 (N_27773,N_20731,N_18232);
xor U27774 (N_27774,N_21758,N_18038);
nand U27775 (N_27775,N_20712,N_20329);
and U27776 (N_27776,N_18369,N_23410);
xor U27777 (N_27777,N_20023,N_19183);
or U27778 (N_27778,N_23418,N_19290);
or U27779 (N_27779,N_20658,N_20920);
nor U27780 (N_27780,N_21811,N_19414);
nand U27781 (N_27781,N_23383,N_23356);
and U27782 (N_27782,N_23426,N_19429);
and U27783 (N_27783,N_21750,N_21100);
xnor U27784 (N_27784,N_18634,N_22509);
or U27785 (N_27785,N_23088,N_22372);
nand U27786 (N_27786,N_18027,N_22383);
or U27787 (N_27787,N_20709,N_19951);
xor U27788 (N_27788,N_22154,N_23375);
and U27789 (N_27789,N_19431,N_19640);
nor U27790 (N_27790,N_22755,N_19059);
nand U27791 (N_27791,N_18225,N_20784);
nor U27792 (N_27792,N_19588,N_19809);
nand U27793 (N_27793,N_18041,N_20110);
or U27794 (N_27794,N_22095,N_18902);
or U27795 (N_27795,N_20760,N_20239);
nor U27796 (N_27796,N_21027,N_21886);
or U27797 (N_27797,N_23624,N_23740);
or U27798 (N_27798,N_18644,N_21545);
and U27799 (N_27799,N_20919,N_19179);
and U27800 (N_27800,N_21979,N_19114);
nand U27801 (N_27801,N_21287,N_18127);
xnor U27802 (N_27802,N_22331,N_22032);
or U27803 (N_27803,N_22780,N_18635);
xnor U27804 (N_27804,N_23958,N_23922);
nand U27805 (N_27805,N_19405,N_18640);
xnor U27806 (N_27806,N_21974,N_21678);
xor U27807 (N_27807,N_18379,N_18982);
xnor U27808 (N_27808,N_23823,N_18250);
xnor U27809 (N_27809,N_21425,N_19999);
nor U27810 (N_27810,N_23028,N_19443);
nor U27811 (N_27811,N_19424,N_22086);
xor U27812 (N_27812,N_22906,N_19448);
nor U27813 (N_27813,N_19649,N_21456);
or U27814 (N_27814,N_19263,N_19387);
nor U27815 (N_27815,N_20806,N_23823);
or U27816 (N_27816,N_18058,N_19260);
xor U27817 (N_27817,N_23147,N_21441);
xor U27818 (N_27818,N_18646,N_22301);
nor U27819 (N_27819,N_23963,N_21769);
nor U27820 (N_27820,N_18625,N_22107);
and U27821 (N_27821,N_20997,N_18830);
and U27822 (N_27822,N_19496,N_22287);
xnor U27823 (N_27823,N_21505,N_19174);
xor U27824 (N_27824,N_20663,N_20919);
nor U27825 (N_27825,N_18039,N_21875);
nor U27826 (N_27826,N_21664,N_19003);
and U27827 (N_27827,N_22979,N_21683);
or U27828 (N_27828,N_19905,N_23302);
nor U27829 (N_27829,N_18467,N_18163);
xor U27830 (N_27830,N_19862,N_23153);
nor U27831 (N_27831,N_18759,N_20194);
xnor U27832 (N_27832,N_20419,N_19516);
and U27833 (N_27833,N_18886,N_21770);
xnor U27834 (N_27834,N_18429,N_18775);
or U27835 (N_27835,N_18620,N_22531);
or U27836 (N_27836,N_21796,N_20562);
nand U27837 (N_27837,N_21630,N_23420);
xnor U27838 (N_27838,N_18008,N_19690);
nor U27839 (N_27839,N_21457,N_20556);
and U27840 (N_27840,N_19074,N_19362);
xnor U27841 (N_27841,N_19353,N_20878);
and U27842 (N_27842,N_18091,N_21643);
nor U27843 (N_27843,N_19729,N_22237);
or U27844 (N_27844,N_19688,N_19142);
or U27845 (N_27845,N_21344,N_23455);
and U27846 (N_27846,N_21893,N_20332);
xnor U27847 (N_27847,N_23419,N_19514);
nand U27848 (N_27848,N_20765,N_22179);
or U27849 (N_27849,N_21777,N_23775);
and U27850 (N_27850,N_20231,N_19479);
or U27851 (N_27851,N_18408,N_19196);
nand U27852 (N_27852,N_22653,N_21908);
and U27853 (N_27853,N_20261,N_21643);
nor U27854 (N_27854,N_23868,N_21444);
and U27855 (N_27855,N_22420,N_19052);
nor U27856 (N_27856,N_18424,N_18293);
xnor U27857 (N_27857,N_19372,N_21258);
and U27858 (N_27858,N_22724,N_20961);
or U27859 (N_27859,N_18248,N_19994);
or U27860 (N_27860,N_19424,N_21727);
and U27861 (N_27861,N_20834,N_20976);
and U27862 (N_27862,N_20925,N_23140);
or U27863 (N_27863,N_20249,N_23034);
nor U27864 (N_27864,N_22784,N_18026);
nor U27865 (N_27865,N_20422,N_19395);
or U27866 (N_27866,N_20046,N_19551);
or U27867 (N_27867,N_22743,N_22044);
and U27868 (N_27868,N_20052,N_21744);
xor U27869 (N_27869,N_23643,N_22881);
xor U27870 (N_27870,N_20447,N_21753);
and U27871 (N_27871,N_21240,N_19517);
nand U27872 (N_27872,N_19488,N_23566);
nand U27873 (N_27873,N_21408,N_20388);
nand U27874 (N_27874,N_20630,N_19502);
or U27875 (N_27875,N_23267,N_18413);
nand U27876 (N_27876,N_18073,N_19438);
nor U27877 (N_27877,N_23360,N_19735);
nand U27878 (N_27878,N_19014,N_20128);
xnor U27879 (N_27879,N_18788,N_20193);
nor U27880 (N_27880,N_20022,N_21684);
nand U27881 (N_27881,N_23635,N_19232);
nor U27882 (N_27882,N_22517,N_22105);
nor U27883 (N_27883,N_21225,N_20031);
nor U27884 (N_27884,N_18447,N_19995);
xor U27885 (N_27885,N_18727,N_22448);
nand U27886 (N_27886,N_23770,N_19379);
nand U27887 (N_27887,N_23726,N_20227);
xor U27888 (N_27888,N_20490,N_22298);
nor U27889 (N_27889,N_21635,N_20557);
and U27890 (N_27890,N_19319,N_21307);
nand U27891 (N_27891,N_22034,N_19690);
nor U27892 (N_27892,N_22726,N_22311);
and U27893 (N_27893,N_18125,N_22852);
or U27894 (N_27894,N_19449,N_23832);
nand U27895 (N_27895,N_21299,N_22468);
and U27896 (N_27896,N_22529,N_19715);
nand U27897 (N_27897,N_23889,N_21473);
xor U27898 (N_27898,N_21637,N_20687);
or U27899 (N_27899,N_22622,N_22564);
xor U27900 (N_27900,N_23812,N_18849);
and U27901 (N_27901,N_21819,N_19889);
nand U27902 (N_27902,N_21269,N_20070);
nor U27903 (N_27903,N_23790,N_23938);
and U27904 (N_27904,N_21848,N_18784);
xor U27905 (N_27905,N_23423,N_20990);
or U27906 (N_27906,N_19493,N_21269);
nand U27907 (N_27907,N_19558,N_18655);
xor U27908 (N_27908,N_22965,N_20976);
nand U27909 (N_27909,N_23036,N_20474);
nor U27910 (N_27910,N_18708,N_21706);
and U27911 (N_27911,N_19468,N_22476);
or U27912 (N_27912,N_22521,N_23141);
nand U27913 (N_27913,N_22731,N_23705);
nand U27914 (N_27914,N_18597,N_22783);
or U27915 (N_27915,N_19542,N_20370);
nor U27916 (N_27916,N_23586,N_21447);
nand U27917 (N_27917,N_19907,N_21351);
or U27918 (N_27918,N_22672,N_22264);
and U27919 (N_27919,N_18707,N_19370);
and U27920 (N_27920,N_22751,N_20067);
xor U27921 (N_27921,N_18007,N_21581);
or U27922 (N_27922,N_19696,N_21882);
xnor U27923 (N_27923,N_23572,N_19809);
nor U27924 (N_27924,N_18466,N_23900);
nand U27925 (N_27925,N_20470,N_20897);
nand U27926 (N_27926,N_21973,N_23434);
nor U27927 (N_27927,N_22246,N_20439);
nand U27928 (N_27928,N_21525,N_18883);
or U27929 (N_27929,N_19382,N_19253);
and U27930 (N_27930,N_21258,N_19154);
nand U27931 (N_27931,N_20444,N_21861);
nor U27932 (N_27932,N_21978,N_18800);
nand U27933 (N_27933,N_21011,N_18538);
xnor U27934 (N_27934,N_21578,N_22809);
and U27935 (N_27935,N_22373,N_18479);
xor U27936 (N_27936,N_22179,N_23053);
or U27937 (N_27937,N_22793,N_22250);
xor U27938 (N_27938,N_18241,N_19247);
xnor U27939 (N_27939,N_21909,N_23972);
or U27940 (N_27940,N_21115,N_22538);
and U27941 (N_27941,N_23839,N_19964);
and U27942 (N_27942,N_22575,N_18741);
xor U27943 (N_27943,N_19034,N_20240);
nor U27944 (N_27944,N_19474,N_23007);
xnor U27945 (N_27945,N_22029,N_23941);
and U27946 (N_27946,N_22998,N_23941);
nand U27947 (N_27947,N_20905,N_23311);
nand U27948 (N_27948,N_18403,N_23745);
xnor U27949 (N_27949,N_21608,N_20582);
and U27950 (N_27950,N_19305,N_22236);
xor U27951 (N_27951,N_23935,N_21788);
or U27952 (N_27952,N_21493,N_19633);
nand U27953 (N_27953,N_18670,N_20598);
nor U27954 (N_27954,N_20650,N_22946);
or U27955 (N_27955,N_21150,N_22461);
xor U27956 (N_27956,N_22714,N_20394);
nor U27957 (N_27957,N_23086,N_19735);
nor U27958 (N_27958,N_20608,N_18683);
xor U27959 (N_27959,N_21566,N_21328);
and U27960 (N_27960,N_23528,N_21868);
nand U27961 (N_27961,N_22622,N_20871);
and U27962 (N_27962,N_19480,N_18588);
xnor U27963 (N_27963,N_21212,N_18179);
xor U27964 (N_27964,N_20377,N_18922);
nor U27965 (N_27965,N_18586,N_19042);
nor U27966 (N_27966,N_23734,N_19098);
nor U27967 (N_27967,N_23853,N_20213);
and U27968 (N_27968,N_21534,N_22144);
or U27969 (N_27969,N_19188,N_20230);
nor U27970 (N_27970,N_20260,N_22929);
xnor U27971 (N_27971,N_18498,N_22980);
or U27972 (N_27972,N_23334,N_21629);
and U27973 (N_27973,N_21127,N_22677);
xor U27974 (N_27974,N_18287,N_22059);
nand U27975 (N_27975,N_22362,N_23947);
and U27976 (N_27976,N_21502,N_21792);
xor U27977 (N_27977,N_21819,N_18375);
xnor U27978 (N_27978,N_19728,N_21550);
nor U27979 (N_27979,N_20587,N_21230);
xor U27980 (N_27980,N_22442,N_22243);
nor U27981 (N_27981,N_23736,N_18245);
and U27982 (N_27982,N_23482,N_20710);
and U27983 (N_27983,N_23142,N_23656);
nor U27984 (N_27984,N_23619,N_21005);
nor U27985 (N_27985,N_19656,N_19959);
nand U27986 (N_27986,N_23463,N_22687);
nor U27987 (N_27987,N_23493,N_19650);
nor U27988 (N_27988,N_21876,N_19656);
nor U27989 (N_27989,N_20533,N_19804);
nand U27990 (N_27990,N_19364,N_18442);
nor U27991 (N_27991,N_23087,N_22356);
xnor U27992 (N_27992,N_22736,N_19001);
nor U27993 (N_27993,N_22205,N_22329);
and U27994 (N_27994,N_18677,N_20432);
or U27995 (N_27995,N_20039,N_19689);
and U27996 (N_27996,N_23222,N_21865);
nand U27997 (N_27997,N_18378,N_21935);
nor U27998 (N_27998,N_18991,N_19306);
and U27999 (N_27999,N_18124,N_22771);
or U28000 (N_28000,N_22237,N_21710);
and U28001 (N_28001,N_19454,N_20842);
and U28002 (N_28002,N_18287,N_18078);
nor U28003 (N_28003,N_23992,N_23899);
and U28004 (N_28004,N_23865,N_23097);
and U28005 (N_28005,N_19884,N_23588);
xnor U28006 (N_28006,N_19319,N_20077);
nor U28007 (N_28007,N_20203,N_23970);
nand U28008 (N_28008,N_19951,N_22165);
and U28009 (N_28009,N_19852,N_18500);
nor U28010 (N_28010,N_20281,N_22327);
xnor U28011 (N_28011,N_19496,N_21907);
xor U28012 (N_28012,N_21610,N_21756);
nor U28013 (N_28013,N_20643,N_19594);
xnor U28014 (N_28014,N_21180,N_19083);
xor U28015 (N_28015,N_22365,N_20394);
or U28016 (N_28016,N_23943,N_18596);
xnor U28017 (N_28017,N_21252,N_18511);
nor U28018 (N_28018,N_22931,N_21972);
nand U28019 (N_28019,N_18641,N_19694);
nand U28020 (N_28020,N_20705,N_21576);
or U28021 (N_28021,N_21844,N_19014);
and U28022 (N_28022,N_20690,N_23203);
or U28023 (N_28023,N_18970,N_23598);
nor U28024 (N_28024,N_19546,N_22570);
and U28025 (N_28025,N_21075,N_21965);
xor U28026 (N_28026,N_19232,N_19622);
or U28027 (N_28027,N_20052,N_18130);
nand U28028 (N_28028,N_18060,N_21694);
or U28029 (N_28029,N_21985,N_23093);
or U28030 (N_28030,N_19460,N_23005);
and U28031 (N_28031,N_21356,N_23004);
nand U28032 (N_28032,N_23619,N_21011);
nand U28033 (N_28033,N_18060,N_23591);
xnor U28034 (N_28034,N_23228,N_18521);
or U28035 (N_28035,N_22664,N_23814);
or U28036 (N_28036,N_20343,N_21261);
nand U28037 (N_28037,N_23312,N_23569);
nor U28038 (N_28038,N_18244,N_21023);
nand U28039 (N_28039,N_21206,N_21031);
nor U28040 (N_28040,N_21233,N_21026);
or U28041 (N_28041,N_19310,N_23395);
or U28042 (N_28042,N_23608,N_19240);
nand U28043 (N_28043,N_19066,N_20931);
and U28044 (N_28044,N_23862,N_18540);
and U28045 (N_28045,N_18819,N_21949);
nor U28046 (N_28046,N_21180,N_19889);
or U28047 (N_28047,N_21078,N_23439);
nor U28048 (N_28048,N_20242,N_22615);
xnor U28049 (N_28049,N_21425,N_20935);
or U28050 (N_28050,N_21448,N_20756);
or U28051 (N_28051,N_18105,N_23408);
or U28052 (N_28052,N_22401,N_23080);
nand U28053 (N_28053,N_23400,N_18640);
xor U28054 (N_28054,N_21097,N_20187);
and U28055 (N_28055,N_21413,N_20840);
nand U28056 (N_28056,N_21134,N_19387);
xor U28057 (N_28057,N_18342,N_23408);
nor U28058 (N_28058,N_22115,N_18266);
or U28059 (N_28059,N_20686,N_21514);
or U28060 (N_28060,N_18859,N_19595);
or U28061 (N_28061,N_21445,N_19122);
nor U28062 (N_28062,N_19113,N_22835);
and U28063 (N_28063,N_22836,N_23204);
nand U28064 (N_28064,N_20550,N_19284);
xnor U28065 (N_28065,N_18874,N_20586);
nor U28066 (N_28066,N_23716,N_19069);
and U28067 (N_28067,N_21325,N_21646);
nor U28068 (N_28068,N_22592,N_22896);
and U28069 (N_28069,N_20321,N_23508);
and U28070 (N_28070,N_18121,N_21233);
or U28071 (N_28071,N_20826,N_19345);
nand U28072 (N_28072,N_18670,N_18975);
xnor U28073 (N_28073,N_18829,N_18749);
or U28074 (N_28074,N_20822,N_19543);
xnor U28075 (N_28075,N_18253,N_18630);
nand U28076 (N_28076,N_23332,N_18415);
nand U28077 (N_28077,N_23698,N_21395);
or U28078 (N_28078,N_22781,N_21684);
nand U28079 (N_28079,N_22309,N_21759);
nand U28080 (N_28080,N_19834,N_21182);
nor U28081 (N_28081,N_23503,N_18192);
nor U28082 (N_28082,N_23485,N_21062);
nand U28083 (N_28083,N_19355,N_23810);
nor U28084 (N_28084,N_18057,N_21335);
nand U28085 (N_28085,N_19143,N_22422);
or U28086 (N_28086,N_19605,N_18601);
xor U28087 (N_28087,N_22335,N_23473);
and U28088 (N_28088,N_22891,N_20539);
or U28089 (N_28089,N_22802,N_21701);
or U28090 (N_28090,N_22499,N_23829);
nand U28091 (N_28091,N_23125,N_18545);
xor U28092 (N_28092,N_18925,N_23792);
and U28093 (N_28093,N_23437,N_20387);
and U28094 (N_28094,N_20615,N_22578);
or U28095 (N_28095,N_21399,N_22755);
nor U28096 (N_28096,N_20919,N_18436);
xor U28097 (N_28097,N_22937,N_19423);
or U28098 (N_28098,N_22231,N_23528);
nor U28099 (N_28099,N_21057,N_20125);
and U28100 (N_28100,N_20253,N_18233);
nor U28101 (N_28101,N_19274,N_18902);
nor U28102 (N_28102,N_18148,N_22490);
xnor U28103 (N_28103,N_20113,N_20271);
xor U28104 (N_28104,N_23216,N_20801);
nand U28105 (N_28105,N_18701,N_19624);
nor U28106 (N_28106,N_20670,N_23987);
nor U28107 (N_28107,N_19390,N_23487);
or U28108 (N_28108,N_21907,N_21761);
or U28109 (N_28109,N_18326,N_20840);
nor U28110 (N_28110,N_22172,N_18471);
nor U28111 (N_28111,N_22113,N_18130);
and U28112 (N_28112,N_19721,N_22107);
or U28113 (N_28113,N_22283,N_18197);
xor U28114 (N_28114,N_18587,N_21593);
and U28115 (N_28115,N_23257,N_19532);
or U28116 (N_28116,N_23013,N_20131);
and U28117 (N_28117,N_21682,N_22364);
or U28118 (N_28118,N_19462,N_19661);
xor U28119 (N_28119,N_19894,N_23033);
xnor U28120 (N_28120,N_21323,N_20509);
and U28121 (N_28121,N_23010,N_23963);
nor U28122 (N_28122,N_23736,N_21536);
nand U28123 (N_28123,N_22863,N_19784);
xor U28124 (N_28124,N_22240,N_22323);
and U28125 (N_28125,N_18119,N_23113);
or U28126 (N_28126,N_20602,N_22451);
or U28127 (N_28127,N_21355,N_22951);
xnor U28128 (N_28128,N_21851,N_21063);
xor U28129 (N_28129,N_21366,N_19512);
nor U28130 (N_28130,N_23744,N_21853);
xnor U28131 (N_28131,N_19568,N_21117);
nor U28132 (N_28132,N_20159,N_22315);
or U28133 (N_28133,N_21259,N_19729);
nand U28134 (N_28134,N_18535,N_18209);
nand U28135 (N_28135,N_22503,N_22212);
nand U28136 (N_28136,N_21928,N_21130);
nor U28137 (N_28137,N_20592,N_21438);
or U28138 (N_28138,N_18349,N_20041);
and U28139 (N_28139,N_18712,N_19485);
xor U28140 (N_28140,N_20908,N_21703);
and U28141 (N_28141,N_22565,N_21781);
nand U28142 (N_28142,N_18112,N_20690);
nand U28143 (N_28143,N_18765,N_22001);
nand U28144 (N_28144,N_19745,N_18116);
nand U28145 (N_28145,N_22507,N_22548);
or U28146 (N_28146,N_20497,N_18653);
and U28147 (N_28147,N_21945,N_18592);
nand U28148 (N_28148,N_23531,N_19934);
xor U28149 (N_28149,N_21615,N_20244);
xnor U28150 (N_28150,N_18723,N_19706);
or U28151 (N_28151,N_23442,N_21086);
nand U28152 (N_28152,N_21462,N_21760);
xor U28153 (N_28153,N_21179,N_22635);
or U28154 (N_28154,N_23998,N_19821);
or U28155 (N_28155,N_19800,N_23029);
or U28156 (N_28156,N_20575,N_22287);
nand U28157 (N_28157,N_18388,N_19420);
xnor U28158 (N_28158,N_21655,N_23696);
or U28159 (N_28159,N_23978,N_19936);
nand U28160 (N_28160,N_19499,N_23758);
nor U28161 (N_28161,N_23942,N_21875);
or U28162 (N_28162,N_18284,N_21074);
or U28163 (N_28163,N_18499,N_18506);
nand U28164 (N_28164,N_19340,N_18281);
xor U28165 (N_28165,N_20222,N_21873);
and U28166 (N_28166,N_20540,N_22430);
nand U28167 (N_28167,N_22262,N_18740);
and U28168 (N_28168,N_23179,N_21270);
nand U28169 (N_28169,N_19708,N_20930);
nand U28170 (N_28170,N_19570,N_21942);
or U28171 (N_28171,N_18074,N_22031);
nor U28172 (N_28172,N_23869,N_20036);
nor U28173 (N_28173,N_23373,N_23587);
and U28174 (N_28174,N_22398,N_20518);
and U28175 (N_28175,N_18470,N_20864);
and U28176 (N_28176,N_18682,N_19579);
or U28177 (N_28177,N_22537,N_22562);
xor U28178 (N_28178,N_19306,N_20843);
or U28179 (N_28179,N_23926,N_19685);
nor U28180 (N_28180,N_23912,N_23472);
xor U28181 (N_28181,N_21984,N_21248);
or U28182 (N_28182,N_23172,N_21420);
nand U28183 (N_28183,N_18915,N_22546);
and U28184 (N_28184,N_22613,N_21537);
nor U28185 (N_28185,N_23069,N_21125);
xnor U28186 (N_28186,N_21938,N_20851);
or U28187 (N_28187,N_18356,N_22690);
nand U28188 (N_28188,N_22933,N_21956);
and U28189 (N_28189,N_19436,N_22034);
xnor U28190 (N_28190,N_21066,N_21418);
or U28191 (N_28191,N_22738,N_23401);
or U28192 (N_28192,N_19000,N_20497);
and U28193 (N_28193,N_20132,N_21584);
and U28194 (N_28194,N_19543,N_19100);
nor U28195 (N_28195,N_19184,N_19614);
nand U28196 (N_28196,N_20743,N_18573);
or U28197 (N_28197,N_21627,N_19952);
nand U28198 (N_28198,N_19521,N_20520);
nor U28199 (N_28199,N_22116,N_21395);
or U28200 (N_28200,N_23449,N_20852);
nand U28201 (N_28201,N_23740,N_22745);
and U28202 (N_28202,N_19682,N_19169);
xor U28203 (N_28203,N_18761,N_23432);
xnor U28204 (N_28204,N_20833,N_18219);
xor U28205 (N_28205,N_21593,N_23245);
nor U28206 (N_28206,N_21707,N_18509);
and U28207 (N_28207,N_21761,N_19431);
or U28208 (N_28208,N_18934,N_21941);
xnor U28209 (N_28209,N_20330,N_18126);
nand U28210 (N_28210,N_21537,N_20286);
nand U28211 (N_28211,N_23436,N_23699);
nor U28212 (N_28212,N_23515,N_22344);
and U28213 (N_28213,N_19255,N_23881);
or U28214 (N_28214,N_22783,N_23633);
or U28215 (N_28215,N_21157,N_21396);
or U28216 (N_28216,N_22342,N_18593);
nand U28217 (N_28217,N_21025,N_20276);
nor U28218 (N_28218,N_18309,N_23566);
nand U28219 (N_28219,N_18883,N_20630);
or U28220 (N_28220,N_18183,N_20676);
or U28221 (N_28221,N_18159,N_21072);
and U28222 (N_28222,N_18739,N_20359);
nor U28223 (N_28223,N_22789,N_19848);
nand U28224 (N_28224,N_22262,N_20035);
and U28225 (N_28225,N_20336,N_20766);
nor U28226 (N_28226,N_19601,N_18327);
xor U28227 (N_28227,N_22755,N_22212);
and U28228 (N_28228,N_18230,N_19842);
nor U28229 (N_28229,N_21351,N_22706);
nor U28230 (N_28230,N_19836,N_19856);
or U28231 (N_28231,N_22275,N_22583);
xnor U28232 (N_28232,N_20231,N_21177);
and U28233 (N_28233,N_21557,N_20499);
or U28234 (N_28234,N_23729,N_22064);
xor U28235 (N_28235,N_20545,N_19916);
or U28236 (N_28236,N_19502,N_21051);
or U28237 (N_28237,N_21824,N_21308);
nor U28238 (N_28238,N_22628,N_21749);
and U28239 (N_28239,N_20639,N_23711);
and U28240 (N_28240,N_18613,N_21903);
xor U28241 (N_28241,N_20755,N_21601);
or U28242 (N_28242,N_18708,N_18933);
nor U28243 (N_28243,N_19586,N_21582);
xnor U28244 (N_28244,N_21237,N_18301);
or U28245 (N_28245,N_23117,N_20621);
nand U28246 (N_28246,N_23212,N_18071);
nor U28247 (N_28247,N_20029,N_21218);
nand U28248 (N_28248,N_23525,N_21105);
xor U28249 (N_28249,N_18587,N_22018);
nor U28250 (N_28250,N_18767,N_22564);
nand U28251 (N_28251,N_22547,N_22271);
nand U28252 (N_28252,N_21913,N_23152);
nand U28253 (N_28253,N_19917,N_21697);
xnor U28254 (N_28254,N_22432,N_22775);
xor U28255 (N_28255,N_21493,N_21563);
xnor U28256 (N_28256,N_18776,N_23197);
nor U28257 (N_28257,N_19082,N_22917);
and U28258 (N_28258,N_22857,N_20762);
nor U28259 (N_28259,N_19171,N_21428);
nand U28260 (N_28260,N_18127,N_22520);
nor U28261 (N_28261,N_20347,N_21695);
nor U28262 (N_28262,N_21031,N_23908);
and U28263 (N_28263,N_23660,N_18240);
nand U28264 (N_28264,N_19623,N_21631);
nand U28265 (N_28265,N_19603,N_18120);
nor U28266 (N_28266,N_18452,N_23004);
nand U28267 (N_28267,N_23138,N_22390);
nand U28268 (N_28268,N_18936,N_22177);
and U28269 (N_28269,N_22994,N_21776);
nand U28270 (N_28270,N_21151,N_21169);
nand U28271 (N_28271,N_21319,N_22903);
nand U28272 (N_28272,N_18108,N_22317);
nand U28273 (N_28273,N_19215,N_23570);
nand U28274 (N_28274,N_21625,N_19708);
or U28275 (N_28275,N_18877,N_21897);
nor U28276 (N_28276,N_22462,N_23682);
or U28277 (N_28277,N_22932,N_18662);
or U28278 (N_28278,N_18575,N_22005);
nor U28279 (N_28279,N_21076,N_22651);
xnor U28280 (N_28280,N_19612,N_20054);
or U28281 (N_28281,N_22851,N_20927);
or U28282 (N_28282,N_22732,N_19465);
nor U28283 (N_28283,N_22991,N_22653);
and U28284 (N_28284,N_23426,N_20204);
nor U28285 (N_28285,N_22593,N_20951);
nand U28286 (N_28286,N_22491,N_19557);
nand U28287 (N_28287,N_22013,N_18225);
or U28288 (N_28288,N_18792,N_19362);
nor U28289 (N_28289,N_23465,N_22115);
and U28290 (N_28290,N_23136,N_20652);
nand U28291 (N_28291,N_21546,N_18684);
or U28292 (N_28292,N_21656,N_18730);
or U28293 (N_28293,N_22664,N_22734);
xor U28294 (N_28294,N_21609,N_21820);
nor U28295 (N_28295,N_22442,N_23920);
and U28296 (N_28296,N_19135,N_23656);
nor U28297 (N_28297,N_21127,N_19809);
and U28298 (N_28298,N_20072,N_21919);
nand U28299 (N_28299,N_21636,N_19951);
or U28300 (N_28300,N_23550,N_23750);
nand U28301 (N_28301,N_20151,N_21361);
xnor U28302 (N_28302,N_22359,N_22150);
xor U28303 (N_28303,N_22358,N_18235);
nand U28304 (N_28304,N_22658,N_18064);
nand U28305 (N_28305,N_18327,N_19466);
and U28306 (N_28306,N_23978,N_19369);
nor U28307 (N_28307,N_19854,N_23936);
and U28308 (N_28308,N_22274,N_20119);
nand U28309 (N_28309,N_18903,N_22351);
xnor U28310 (N_28310,N_18131,N_20200);
and U28311 (N_28311,N_20234,N_22608);
xnor U28312 (N_28312,N_18133,N_20024);
and U28313 (N_28313,N_23569,N_18899);
nand U28314 (N_28314,N_22181,N_20809);
and U28315 (N_28315,N_20556,N_22793);
nand U28316 (N_28316,N_20524,N_21936);
or U28317 (N_28317,N_18211,N_21617);
nand U28318 (N_28318,N_23520,N_23305);
nand U28319 (N_28319,N_23453,N_20069);
xor U28320 (N_28320,N_20582,N_18462);
xnor U28321 (N_28321,N_23586,N_18129);
nor U28322 (N_28322,N_21073,N_19945);
nor U28323 (N_28323,N_19111,N_18599);
and U28324 (N_28324,N_19127,N_19391);
nand U28325 (N_28325,N_23491,N_20519);
and U28326 (N_28326,N_23700,N_20237);
and U28327 (N_28327,N_18004,N_21738);
nand U28328 (N_28328,N_21580,N_19849);
and U28329 (N_28329,N_19807,N_23601);
nor U28330 (N_28330,N_18700,N_21872);
nand U28331 (N_28331,N_19950,N_19691);
xnor U28332 (N_28332,N_21015,N_19013);
nand U28333 (N_28333,N_19385,N_18576);
nor U28334 (N_28334,N_22977,N_20192);
and U28335 (N_28335,N_20745,N_20033);
or U28336 (N_28336,N_19646,N_20347);
or U28337 (N_28337,N_22445,N_21235);
xnor U28338 (N_28338,N_23444,N_19894);
xnor U28339 (N_28339,N_22322,N_20266);
nor U28340 (N_28340,N_19379,N_23969);
xnor U28341 (N_28341,N_19504,N_22586);
nand U28342 (N_28342,N_19261,N_20403);
nand U28343 (N_28343,N_20995,N_18864);
nand U28344 (N_28344,N_18144,N_20677);
xnor U28345 (N_28345,N_23913,N_18750);
or U28346 (N_28346,N_19474,N_19045);
nor U28347 (N_28347,N_20560,N_18194);
and U28348 (N_28348,N_19909,N_19141);
nor U28349 (N_28349,N_18598,N_23546);
xor U28350 (N_28350,N_20889,N_21307);
nand U28351 (N_28351,N_22138,N_20192);
and U28352 (N_28352,N_22822,N_19066);
xnor U28353 (N_28353,N_21700,N_23845);
nor U28354 (N_28354,N_20700,N_19262);
xor U28355 (N_28355,N_18227,N_20119);
and U28356 (N_28356,N_18252,N_21590);
nor U28357 (N_28357,N_19014,N_21615);
nand U28358 (N_28358,N_19042,N_23223);
and U28359 (N_28359,N_19023,N_22262);
nor U28360 (N_28360,N_22570,N_22230);
and U28361 (N_28361,N_21644,N_20563);
nor U28362 (N_28362,N_23136,N_19883);
nor U28363 (N_28363,N_22909,N_20355);
nor U28364 (N_28364,N_23116,N_21307);
nor U28365 (N_28365,N_23865,N_19494);
nand U28366 (N_28366,N_22541,N_18897);
xnor U28367 (N_28367,N_18574,N_21795);
xor U28368 (N_28368,N_21149,N_21674);
xor U28369 (N_28369,N_23178,N_23895);
or U28370 (N_28370,N_23582,N_20515);
and U28371 (N_28371,N_21843,N_22578);
nand U28372 (N_28372,N_22576,N_18040);
and U28373 (N_28373,N_21357,N_18689);
and U28374 (N_28374,N_20242,N_19709);
nand U28375 (N_28375,N_18649,N_21309);
or U28376 (N_28376,N_20638,N_18878);
nand U28377 (N_28377,N_20306,N_18566);
nand U28378 (N_28378,N_19029,N_21998);
nand U28379 (N_28379,N_23512,N_19242);
nor U28380 (N_28380,N_23013,N_23064);
or U28381 (N_28381,N_18128,N_19953);
nand U28382 (N_28382,N_21560,N_21103);
xor U28383 (N_28383,N_22802,N_20977);
nor U28384 (N_28384,N_18213,N_21836);
nor U28385 (N_28385,N_20845,N_19416);
or U28386 (N_28386,N_22199,N_23375);
nand U28387 (N_28387,N_21116,N_22363);
xor U28388 (N_28388,N_18772,N_22710);
xnor U28389 (N_28389,N_20772,N_23372);
nand U28390 (N_28390,N_18157,N_19698);
nand U28391 (N_28391,N_22902,N_20169);
xor U28392 (N_28392,N_18941,N_21893);
or U28393 (N_28393,N_19395,N_22189);
or U28394 (N_28394,N_21995,N_21231);
nor U28395 (N_28395,N_22493,N_20768);
and U28396 (N_28396,N_22409,N_21306);
or U28397 (N_28397,N_20821,N_22924);
and U28398 (N_28398,N_19230,N_22515);
xor U28399 (N_28399,N_22670,N_19573);
nor U28400 (N_28400,N_18230,N_22865);
nor U28401 (N_28401,N_19008,N_18383);
nand U28402 (N_28402,N_22516,N_22072);
nor U28403 (N_28403,N_21983,N_20952);
xnor U28404 (N_28404,N_21346,N_19040);
nor U28405 (N_28405,N_19930,N_18106);
or U28406 (N_28406,N_20065,N_22745);
xor U28407 (N_28407,N_22771,N_23849);
and U28408 (N_28408,N_19109,N_20971);
or U28409 (N_28409,N_22914,N_18497);
nand U28410 (N_28410,N_22024,N_21717);
or U28411 (N_28411,N_18323,N_20830);
and U28412 (N_28412,N_19188,N_20460);
xor U28413 (N_28413,N_23482,N_20777);
or U28414 (N_28414,N_22512,N_23927);
nand U28415 (N_28415,N_22650,N_23476);
nand U28416 (N_28416,N_19024,N_19478);
or U28417 (N_28417,N_21143,N_18789);
or U28418 (N_28418,N_23688,N_19321);
nand U28419 (N_28419,N_19823,N_18427);
nor U28420 (N_28420,N_21800,N_18426);
and U28421 (N_28421,N_21954,N_19016);
xnor U28422 (N_28422,N_18096,N_22528);
nor U28423 (N_28423,N_19182,N_20116);
xor U28424 (N_28424,N_19664,N_21517);
xor U28425 (N_28425,N_22318,N_20593);
xnor U28426 (N_28426,N_19270,N_20582);
xor U28427 (N_28427,N_22112,N_21036);
nand U28428 (N_28428,N_18878,N_23528);
nand U28429 (N_28429,N_20562,N_18169);
or U28430 (N_28430,N_18675,N_19133);
or U28431 (N_28431,N_22211,N_18805);
xnor U28432 (N_28432,N_23453,N_22860);
nor U28433 (N_28433,N_18401,N_23585);
and U28434 (N_28434,N_22182,N_18838);
or U28435 (N_28435,N_20990,N_23176);
xnor U28436 (N_28436,N_22407,N_18660);
or U28437 (N_28437,N_21271,N_23402);
xor U28438 (N_28438,N_19873,N_18755);
xnor U28439 (N_28439,N_19795,N_23452);
and U28440 (N_28440,N_19653,N_23587);
nor U28441 (N_28441,N_18825,N_19186);
nand U28442 (N_28442,N_21746,N_22207);
or U28443 (N_28443,N_21936,N_21120);
or U28444 (N_28444,N_21256,N_23200);
nand U28445 (N_28445,N_18930,N_23702);
or U28446 (N_28446,N_19358,N_23725);
and U28447 (N_28447,N_21370,N_21967);
nor U28448 (N_28448,N_21320,N_18007);
nand U28449 (N_28449,N_23614,N_21605);
or U28450 (N_28450,N_19943,N_19722);
xor U28451 (N_28451,N_19034,N_18923);
nand U28452 (N_28452,N_19244,N_18085);
nor U28453 (N_28453,N_22384,N_20294);
or U28454 (N_28454,N_18367,N_21158);
and U28455 (N_28455,N_20262,N_22205);
and U28456 (N_28456,N_18534,N_20524);
or U28457 (N_28457,N_20588,N_23517);
or U28458 (N_28458,N_18133,N_23764);
and U28459 (N_28459,N_20079,N_18410);
or U28460 (N_28460,N_21195,N_20881);
or U28461 (N_28461,N_21625,N_22897);
xor U28462 (N_28462,N_20816,N_19097);
and U28463 (N_28463,N_22806,N_19043);
nand U28464 (N_28464,N_22971,N_19354);
nor U28465 (N_28465,N_22944,N_23284);
nor U28466 (N_28466,N_19809,N_21129);
nand U28467 (N_28467,N_23192,N_18504);
xor U28468 (N_28468,N_18324,N_19243);
or U28469 (N_28469,N_18442,N_21635);
nand U28470 (N_28470,N_19447,N_22803);
and U28471 (N_28471,N_22305,N_21187);
or U28472 (N_28472,N_18627,N_18691);
and U28473 (N_28473,N_18115,N_18772);
or U28474 (N_28474,N_20124,N_23136);
xnor U28475 (N_28475,N_18487,N_23277);
or U28476 (N_28476,N_18269,N_21256);
or U28477 (N_28477,N_19298,N_21920);
xor U28478 (N_28478,N_22458,N_18980);
nor U28479 (N_28479,N_19561,N_21740);
nand U28480 (N_28480,N_21938,N_23585);
nand U28481 (N_28481,N_18498,N_19007);
and U28482 (N_28482,N_20341,N_21728);
nor U28483 (N_28483,N_20899,N_19545);
nor U28484 (N_28484,N_19914,N_23485);
nor U28485 (N_28485,N_22222,N_22756);
and U28486 (N_28486,N_23963,N_22226);
or U28487 (N_28487,N_23864,N_19481);
or U28488 (N_28488,N_18460,N_22730);
xnor U28489 (N_28489,N_21452,N_19467);
nor U28490 (N_28490,N_19742,N_18604);
or U28491 (N_28491,N_19288,N_22518);
and U28492 (N_28492,N_23329,N_22843);
nand U28493 (N_28493,N_22748,N_18239);
or U28494 (N_28494,N_22709,N_20382);
nand U28495 (N_28495,N_19322,N_22138);
nor U28496 (N_28496,N_23987,N_18409);
xnor U28497 (N_28497,N_20326,N_20446);
nor U28498 (N_28498,N_21165,N_22474);
xor U28499 (N_28499,N_20859,N_23672);
or U28500 (N_28500,N_19924,N_22137);
or U28501 (N_28501,N_21524,N_23582);
nor U28502 (N_28502,N_23453,N_23589);
nand U28503 (N_28503,N_20147,N_23758);
or U28504 (N_28504,N_21326,N_19893);
xor U28505 (N_28505,N_23283,N_18392);
or U28506 (N_28506,N_21082,N_22766);
nor U28507 (N_28507,N_18408,N_22418);
or U28508 (N_28508,N_18125,N_21227);
xnor U28509 (N_28509,N_22944,N_23390);
or U28510 (N_28510,N_21796,N_22058);
and U28511 (N_28511,N_20302,N_23847);
and U28512 (N_28512,N_21165,N_23422);
xnor U28513 (N_28513,N_20487,N_21981);
and U28514 (N_28514,N_23558,N_21770);
or U28515 (N_28515,N_19950,N_21457);
and U28516 (N_28516,N_18862,N_21218);
and U28517 (N_28517,N_21382,N_23676);
xnor U28518 (N_28518,N_20765,N_23082);
or U28519 (N_28519,N_18625,N_22692);
nand U28520 (N_28520,N_19656,N_18125);
and U28521 (N_28521,N_18315,N_21675);
and U28522 (N_28522,N_18731,N_21617);
and U28523 (N_28523,N_20975,N_19119);
nand U28524 (N_28524,N_19438,N_23557);
nor U28525 (N_28525,N_21657,N_22820);
and U28526 (N_28526,N_21217,N_22203);
and U28527 (N_28527,N_18724,N_18424);
or U28528 (N_28528,N_21792,N_19907);
nand U28529 (N_28529,N_23379,N_18723);
or U28530 (N_28530,N_21601,N_20220);
xnor U28531 (N_28531,N_18877,N_22654);
xor U28532 (N_28532,N_18995,N_19811);
xor U28533 (N_28533,N_20703,N_18098);
xor U28534 (N_28534,N_18504,N_18091);
nor U28535 (N_28535,N_20666,N_23939);
or U28536 (N_28536,N_19444,N_18085);
xnor U28537 (N_28537,N_23803,N_20489);
xnor U28538 (N_28538,N_20848,N_21822);
and U28539 (N_28539,N_23060,N_20507);
xor U28540 (N_28540,N_23473,N_19665);
nor U28541 (N_28541,N_18085,N_19108);
xnor U28542 (N_28542,N_19743,N_18352);
and U28543 (N_28543,N_22061,N_22023);
nor U28544 (N_28544,N_19061,N_20905);
xor U28545 (N_28545,N_21266,N_19638);
or U28546 (N_28546,N_22861,N_19041);
xor U28547 (N_28547,N_22773,N_20711);
or U28548 (N_28548,N_21222,N_21673);
and U28549 (N_28549,N_18351,N_21326);
nand U28550 (N_28550,N_20622,N_20078);
and U28551 (N_28551,N_20636,N_20831);
or U28552 (N_28552,N_19060,N_23343);
nand U28553 (N_28553,N_19353,N_21108);
or U28554 (N_28554,N_21478,N_22138);
or U28555 (N_28555,N_20990,N_22626);
xor U28556 (N_28556,N_21000,N_23053);
nand U28557 (N_28557,N_20173,N_21120);
nor U28558 (N_28558,N_21904,N_20182);
nor U28559 (N_28559,N_21336,N_22711);
nor U28560 (N_28560,N_23152,N_18586);
xor U28561 (N_28561,N_19006,N_19875);
nor U28562 (N_28562,N_20282,N_18279);
xor U28563 (N_28563,N_18205,N_23275);
and U28564 (N_28564,N_23924,N_23221);
and U28565 (N_28565,N_23749,N_21801);
nand U28566 (N_28566,N_20399,N_18144);
and U28567 (N_28567,N_23057,N_18239);
nor U28568 (N_28568,N_23022,N_20686);
nor U28569 (N_28569,N_18849,N_23566);
and U28570 (N_28570,N_18947,N_21569);
nand U28571 (N_28571,N_19005,N_20226);
or U28572 (N_28572,N_20390,N_20535);
xnor U28573 (N_28573,N_20722,N_21339);
nor U28574 (N_28574,N_19914,N_22360);
and U28575 (N_28575,N_21386,N_19183);
and U28576 (N_28576,N_18099,N_19793);
and U28577 (N_28577,N_18651,N_21552);
or U28578 (N_28578,N_22841,N_19577);
nor U28579 (N_28579,N_22027,N_20630);
nor U28580 (N_28580,N_20572,N_18724);
nor U28581 (N_28581,N_19053,N_23870);
xor U28582 (N_28582,N_21850,N_21890);
xor U28583 (N_28583,N_18793,N_19028);
nand U28584 (N_28584,N_20868,N_18376);
xnor U28585 (N_28585,N_20250,N_23493);
or U28586 (N_28586,N_23999,N_18298);
and U28587 (N_28587,N_22853,N_22543);
nor U28588 (N_28588,N_22370,N_22198);
nand U28589 (N_28589,N_21351,N_23252);
xnor U28590 (N_28590,N_20949,N_23418);
nand U28591 (N_28591,N_19833,N_19136);
or U28592 (N_28592,N_22446,N_18730);
nand U28593 (N_28593,N_18697,N_22240);
and U28594 (N_28594,N_20926,N_18777);
xnor U28595 (N_28595,N_21977,N_22526);
xor U28596 (N_28596,N_23326,N_21242);
or U28597 (N_28597,N_23063,N_18697);
nand U28598 (N_28598,N_19340,N_20578);
and U28599 (N_28599,N_18040,N_20186);
xnor U28600 (N_28600,N_21247,N_22721);
or U28601 (N_28601,N_21633,N_18082);
nor U28602 (N_28602,N_23446,N_23996);
or U28603 (N_28603,N_22143,N_21722);
xor U28604 (N_28604,N_18527,N_18895);
or U28605 (N_28605,N_20327,N_23395);
xnor U28606 (N_28606,N_19559,N_18178);
nand U28607 (N_28607,N_19294,N_19108);
nand U28608 (N_28608,N_18887,N_22403);
nor U28609 (N_28609,N_20716,N_19420);
or U28610 (N_28610,N_18891,N_22534);
nor U28611 (N_28611,N_19914,N_20598);
nand U28612 (N_28612,N_19405,N_20202);
or U28613 (N_28613,N_22624,N_19935);
nand U28614 (N_28614,N_20767,N_19770);
nand U28615 (N_28615,N_23104,N_19510);
xor U28616 (N_28616,N_20884,N_20963);
nor U28617 (N_28617,N_21754,N_20350);
or U28618 (N_28618,N_18110,N_22781);
and U28619 (N_28619,N_18182,N_22368);
or U28620 (N_28620,N_20806,N_23774);
and U28621 (N_28621,N_21678,N_23017);
and U28622 (N_28622,N_21859,N_23966);
nor U28623 (N_28623,N_22232,N_19607);
and U28624 (N_28624,N_19697,N_22570);
nor U28625 (N_28625,N_19372,N_21180);
and U28626 (N_28626,N_21156,N_18331);
nor U28627 (N_28627,N_19806,N_21783);
and U28628 (N_28628,N_18665,N_22726);
and U28629 (N_28629,N_18150,N_18648);
nor U28630 (N_28630,N_20517,N_21683);
xnor U28631 (N_28631,N_21559,N_19993);
or U28632 (N_28632,N_19692,N_18170);
nor U28633 (N_28633,N_21638,N_22885);
and U28634 (N_28634,N_18415,N_20320);
nand U28635 (N_28635,N_18564,N_22675);
or U28636 (N_28636,N_18151,N_22533);
and U28637 (N_28637,N_20108,N_20185);
nand U28638 (N_28638,N_19010,N_21071);
and U28639 (N_28639,N_23563,N_20049);
or U28640 (N_28640,N_19640,N_19982);
nand U28641 (N_28641,N_20961,N_20257);
xnor U28642 (N_28642,N_22872,N_22083);
nor U28643 (N_28643,N_21820,N_20095);
nand U28644 (N_28644,N_18506,N_22936);
or U28645 (N_28645,N_21618,N_18061);
nor U28646 (N_28646,N_23638,N_21511);
xor U28647 (N_28647,N_18702,N_19275);
or U28648 (N_28648,N_23576,N_21235);
or U28649 (N_28649,N_19901,N_21185);
xor U28650 (N_28650,N_18413,N_20966);
xor U28651 (N_28651,N_23364,N_19053);
and U28652 (N_28652,N_22621,N_19260);
or U28653 (N_28653,N_20204,N_23725);
nand U28654 (N_28654,N_23768,N_22900);
or U28655 (N_28655,N_22742,N_23203);
nand U28656 (N_28656,N_19027,N_23521);
xor U28657 (N_28657,N_23932,N_22097);
and U28658 (N_28658,N_18700,N_20785);
and U28659 (N_28659,N_19865,N_20257);
nand U28660 (N_28660,N_22769,N_21757);
nand U28661 (N_28661,N_23158,N_21418);
nand U28662 (N_28662,N_20281,N_22830);
nor U28663 (N_28663,N_19847,N_22883);
nand U28664 (N_28664,N_21643,N_19130);
nand U28665 (N_28665,N_20291,N_18214);
nand U28666 (N_28666,N_23801,N_18774);
nor U28667 (N_28667,N_21903,N_23282);
and U28668 (N_28668,N_19675,N_22247);
xnor U28669 (N_28669,N_23181,N_19171);
nand U28670 (N_28670,N_19613,N_23884);
xnor U28671 (N_28671,N_18677,N_19855);
or U28672 (N_28672,N_23164,N_22954);
or U28673 (N_28673,N_22271,N_22367);
nor U28674 (N_28674,N_22936,N_21723);
xnor U28675 (N_28675,N_23363,N_21680);
or U28676 (N_28676,N_20830,N_22163);
nand U28677 (N_28677,N_19992,N_23729);
xnor U28678 (N_28678,N_21455,N_22097);
or U28679 (N_28679,N_20235,N_19504);
xor U28680 (N_28680,N_20070,N_21135);
xor U28681 (N_28681,N_23336,N_18016);
or U28682 (N_28682,N_23760,N_22901);
and U28683 (N_28683,N_22530,N_22247);
xor U28684 (N_28684,N_23046,N_21095);
xnor U28685 (N_28685,N_18430,N_20607);
xor U28686 (N_28686,N_20944,N_22442);
xor U28687 (N_28687,N_23881,N_18785);
xnor U28688 (N_28688,N_22284,N_19079);
nand U28689 (N_28689,N_20811,N_19294);
xnor U28690 (N_28690,N_21632,N_18070);
or U28691 (N_28691,N_22803,N_21672);
xor U28692 (N_28692,N_23266,N_22281);
nor U28693 (N_28693,N_21417,N_18625);
nand U28694 (N_28694,N_23255,N_23653);
nand U28695 (N_28695,N_18532,N_20718);
nor U28696 (N_28696,N_20878,N_22526);
nor U28697 (N_28697,N_20920,N_20002);
nor U28698 (N_28698,N_18692,N_19001);
nor U28699 (N_28699,N_23439,N_18202);
or U28700 (N_28700,N_21369,N_21521);
nand U28701 (N_28701,N_23906,N_20816);
or U28702 (N_28702,N_23858,N_18027);
and U28703 (N_28703,N_20341,N_21104);
nand U28704 (N_28704,N_20770,N_23020);
nor U28705 (N_28705,N_23950,N_22485);
and U28706 (N_28706,N_20261,N_18126);
xnor U28707 (N_28707,N_18044,N_22709);
nor U28708 (N_28708,N_22974,N_23410);
nor U28709 (N_28709,N_20058,N_21066);
nor U28710 (N_28710,N_19385,N_19288);
and U28711 (N_28711,N_20156,N_23449);
nor U28712 (N_28712,N_20473,N_19966);
nor U28713 (N_28713,N_20986,N_22236);
nand U28714 (N_28714,N_23152,N_22943);
and U28715 (N_28715,N_22288,N_23497);
nand U28716 (N_28716,N_23322,N_23326);
xnor U28717 (N_28717,N_20397,N_18136);
and U28718 (N_28718,N_20645,N_22060);
and U28719 (N_28719,N_22844,N_22288);
or U28720 (N_28720,N_18646,N_18872);
xnor U28721 (N_28721,N_21293,N_23361);
nand U28722 (N_28722,N_22627,N_21064);
or U28723 (N_28723,N_19170,N_21719);
xor U28724 (N_28724,N_20533,N_19378);
or U28725 (N_28725,N_21432,N_21539);
nand U28726 (N_28726,N_21446,N_20606);
and U28727 (N_28727,N_20152,N_21582);
and U28728 (N_28728,N_20220,N_18538);
xnor U28729 (N_28729,N_19799,N_21630);
nand U28730 (N_28730,N_22891,N_22243);
nand U28731 (N_28731,N_19304,N_23663);
and U28732 (N_28732,N_21381,N_20292);
nor U28733 (N_28733,N_22576,N_18602);
nand U28734 (N_28734,N_18396,N_18692);
xnor U28735 (N_28735,N_20186,N_20803);
nor U28736 (N_28736,N_19861,N_22679);
nand U28737 (N_28737,N_23338,N_21390);
nand U28738 (N_28738,N_23297,N_19524);
and U28739 (N_28739,N_19320,N_23355);
xor U28740 (N_28740,N_19487,N_19451);
nand U28741 (N_28741,N_23285,N_23437);
and U28742 (N_28742,N_18271,N_20000);
and U28743 (N_28743,N_20640,N_18327);
or U28744 (N_28744,N_19873,N_20081);
nor U28745 (N_28745,N_20440,N_20447);
xor U28746 (N_28746,N_20003,N_21037);
and U28747 (N_28747,N_21459,N_18100);
xnor U28748 (N_28748,N_19842,N_22715);
xor U28749 (N_28749,N_21483,N_18878);
xnor U28750 (N_28750,N_21179,N_20068);
nand U28751 (N_28751,N_22507,N_18128);
xor U28752 (N_28752,N_22136,N_20774);
nor U28753 (N_28753,N_22274,N_18023);
nand U28754 (N_28754,N_18216,N_19577);
nand U28755 (N_28755,N_18875,N_21485);
xor U28756 (N_28756,N_23802,N_20020);
or U28757 (N_28757,N_23855,N_23434);
or U28758 (N_28758,N_19779,N_21561);
nand U28759 (N_28759,N_23650,N_19688);
nand U28760 (N_28760,N_23730,N_18063);
and U28761 (N_28761,N_20586,N_20470);
or U28762 (N_28762,N_19840,N_23993);
xor U28763 (N_28763,N_18639,N_19817);
xnor U28764 (N_28764,N_18807,N_19671);
nand U28765 (N_28765,N_18163,N_23075);
or U28766 (N_28766,N_22139,N_23837);
or U28767 (N_28767,N_21340,N_23273);
and U28768 (N_28768,N_20173,N_23204);
or U28769 (N_28769,N_19021,N_19089);
nand U28770 (N_28770,N_22029,N_21620);
or U28771 (N_28771,N_22739,N_20189);
and U28772 (N_28772,N_20335,N_18564);
and U28773 (N_28773,N_19247,N_20395);
nor U28774 (N_28774,N_20082,N_21720);
nor U28775 (N_28775,N_19934,N_22339);
nand U28776 (N_28776,N_20552,N_20726);
or U28777 (N_28777,N_21282,N_23634);
xor U28778 (N_28778,N_20074,N_23027);
nor U28779 (N_28779,N_21255,N_19591);
and U28780 (N_28780,N_20613,N_18192);
and U28781 (N_28781,N_19416,N_19245);
nand U28782 (N_28782,N_20871,N_19537);
and U28783 (N_28783,N_19203,N_20805);
and U28784 (N_28784,N_18078,N_22459);
nand U28785 (N_28785,N_19853,N_20501);
and U28786 (N_28786,N_20187,N_23390);
nand U28787 (N_28787,N_21553,N_20970);
xnor U28788 (N_28788,N_18141,N_18315);
xor U28789 (N_28789,N_23019,N_22237);
or U28790 (N_28790,N_19669,N_23539);
xor U28791 (N_28791,N_21898,N_23083);
and U28792 (N_28792,N_23428,N_18406);
xnor U28793 (N_28793,N_22235,N_23623);
nand U28794 (N_28794,N_23345,N_20663);
or U28795 (N_28795,N_23904,N_18428);
xnor U28796 (N_28796,N_21572,N_22201);
or U28797 (N_28797,N_23311,N_23342);
nor U28798 (N_28798,N_22931,N_22340);
nand U28799 (N_28799,N_20312,N_21982);
nor U28800 (N_28800,N_23353,N_22128);
xnor U28801 (N_28801,N_21807,N_19128);
nor U28802 (N_28802,N_21257,N_22141);
and U28803 (N_28803,N_22136,N_22610);
xor U28804 (N_28804,N_20298,N_18347);
and U28805 (N_28805,N_23673,N_19316);
and U28806 (N_28806,N_22873,N_18678);
xor U28807 (N_28807,N_23504,N_20742);
nor U28808 (N_28808,N_21299,N_19234);
nor U28809 (N_28809,N_23688,N_23773);
or U28810 (N_28810,N_23186,N_20895);
nor U28811 (N_28811,N_18433,N_18804);
and U28812 (N_28812,N_18367,N_23190);
nor U28813 (N_28813,N_19212,N_22353);
or U28814 (N_28814,N_19169,N_23547);
nand U28815 (N_28815,N_20735,N_23699);
or U28816 (N_28816,N_21614,N_19705);
nand U28817 (N_28817,N_20822,N_23674);
xor U28818 (N_28818,N_18305,N_22843);
nor U28819 (N_28819,N_19878,N_23610);
xnor U28820 (N_28820,N_23253,N_18410);
xor U28821 (N_28821,N_18867,N_19630);
or U28822 (N_28822,N_18259,N_23585);
nor U28823 (N_28823,N_20597,N_21974);
and U28824 (N_28824,N_22250,N_19149);
nor U28825 (N_28825,N_21095,N_19690);
nand U28826 (N_28826,N_23441,N_22829);
xor U28827 (N_28827,N_22309,N_19886);
nor U28828 (N_28828,N_22124,N_20098);
nand U28829 (N_28829,N_19089,N_21924);
nand U28830 (N_28830,N_20196,N_18198);
or U28831 (N_28831,N_22838,N_23525);
nand U28832 (N_28832,N_18909,N_19952);
nand U28833 (N_28833,N_22598,N_23350);
nand U28834 (N_28834,N_19087,N_20823);
or U28835 (N_28835,N_22159,N_21251);
and U28836 (N_28836,N_19915,N_22318);
nand U28837 (N_28837,N_19633,N_20158);
nor U28838 (N_28838,N_22416,N_19181);
xor U28839 (N_28839,N_22107,N_19571);
nor U28840 (N_28840,N_21983,N_23771);
and U28841 (N_28841,N_23025,N_18939);
xnor U28842 (N_28842,N_18761,N_18963);
nor U28843 (N_28843,N_18892,N_19344);
nand U28844 (N_28844,N_19661,N_23659);
nor U28845 (N_28845,N_20631,N_22510);
and U28846 (N_28846,N_20756,N_19749);
nand U28847 (N_28847,N_19382,N_18338);
and U28848 (N_28848,N_23319,N_22596);
nor U28849 (N_28849,N_19153,N_23457);
xor U28850 (N_28850,N_22575,N_18905);
and U28851 (N_28851,N_19799,N_19631);
and U28852 (N_28852,N_20574,N_18570);
and U28853 (N_28853,N_18032,N_23846);
xor U28854 (N_28854,N_23587,N_20776);
nor U28855 (N_28855,N_21780,N_20561);
xnor U28856 (N_28856,N_22091,N_20054);
or U28857 (N_28857,N_23440,N_23770);
xor U28858 (N_28858,N_18794,N_18546);
and U28859 (N_28859,N_19774,N_18943);
nor U28860 (N_28860,N_23413,N_20245);
nor U28861 (N_28861,N_20716,N_21655);
nand U28862 (N_28862,N_19145,N_23599);
and U28863 (N_28863,N_22786,N_20812);
nand U28864 (N_28864,N_21051,N_20489);
or U28865 (N_28865,N_22988,N_19191);
nor U28866 (N_28866,N_23697,N_20593);
and U28867 (N_28867,N_19933,N_22710);
and U28868 (N_28868,N_21943,N_19235);
or U28869 (N_28869,N_18183,N_19711);
and U28870 (N_28870,N_23629,N_18504);
xor U28871 (N_28871,N_23262,N_22298);
or U28872 (N_28872,N_19391,N_22557);
nand U28873 (N_28873,N_23874,N_23939);
nand U28874 (N_28874,N_19651,N_22269);
xnor U28875 (N_28875,N_19047,N_23624);
nor U28876 (N_28876,N_22564,N_18522);
xnor U28877 (N_28877,N_19149,N_23397);
and U28878 (N_28878,N_22960,N_21214);
xnor U28879 (N_28879,N_23940,N_19815);
and U28880 (N_28880,N_20200,N_19957);
nand U28881 (N_28881,N_19971,N_23345);
nand U28882 (N_28882,N_20683,N_20012);
nand U28883 (N_28883,N_19434,N_22190);
nor U28884 (N_28884,N_22430,N_20310);
nor U28885 (N_28885,N_23555,N_19248);
nand U28886 (N_28886,N_22255,N_19835);
xor U28887 (N_28887,N_23405,N_18498);
or U28888 (N_28888,N_18947,N_18888);
or U28889 (N_28889,N_22147,N_21028);
or U28890 (N_28890,N_18262,N_22274);
and U28891 (N_28891,N_20139,N_18094);
nor U28892 (N_28892,N_23748,N_23090);
nand U28893 (N_28893,N_21107,N_22431);
and U28894 (N_28894,N_20831,N_18528);
xnor U28895 (N_28895,N_18005,N_22095);
and U28896 (N_28896,N_22253,N_18135);
or U28897 (N_28897,N_21835,N_22222);
nor U28898 (N_28898,N_19096,N_21599);
nand U28899 (N_28899,N_23911,N_23086);
xnor U28900 (N_28900,N_22731,N_23552);
xor U28901 (N_28901,N_22868,N_23670);
nor U28902 (N_28902,N_19439,N_19618);
xnor U28903 (N_28903,N_21433,N_21053);
or U28904 (N_28904,N_19092,N_18854);
nor U28905 (N_28905,N_22783,N_22387);
and U28906 (N_28906,N_18091,N_19161);
nand U28907 (N_28907,N_22066,N_20723);
nor U28908 (N_28908,N_18227,N_22752);
nand U28909 (N_28909,N_22112,N_23568);
xnor U28910 (N_28910,N_21796,N_21641);
nand U28911 (N_28911,N_18567,N_23940);
nor U28912 (N_28912,N_21091,N_22576);
xnor U28913 (N_28913,N_23915,N_18066);
xor U28914 (N_28914,N_18442,N_19233);
nand U28915 (N_28915,N_21945,N_20742);
or U28916 (N_28916,N_22793,N_22338);
xnor U28917 (N_28917,N_19765,N_21431);
nor U28918 (N_28918,N_18833,N_18940);
nand U28919 (N_28919,N_21524,N_22045);
and U28920 (N_28920,N_21001,N_19961);
nor U28921 (N_28921,N_19996,N_23527);
or U28922 (N_28922,N_23621,N_19514);
and U28923 (N_28923,N_20051,N_20297);
xor U28924 (N_28924,N_23948,N_23227);
nand U28925 (N_28925,N_21438,N_20728);
nand U28926 (N_28926,N_23666,N_19135);
and U28927 (N_28927,N_21408,N_18526);
nor U28928 (N_28928,N_19231,N_23164);
xnor U28929 (N_28929,N_19351,N_20483);
xnor U28930 (N_28930,N_23133,N_22772);
and U28931 (N_28931,N_19971,N_19051);
and U28932 (N_28932,N_21559,N_21602);
nor U28933 (N_28933,N_22294,N_18211);
nor U28934 (N_28934,N_18601,N_23569);
and U28935 (N_28935,N_19905,N_18266);
or U28936 (N_28936,N_23200,N_23929);
nor U28937 (N_28937,N_22307,N_21442);
xnor U28938 (N_28938,N_23481,N_22290);
and U28939 (N_28939,N_21214,N_20272);
or U28940 (N_28940,N_19894,N_20220);
xor U28941 (N_28941,N_20272,N_19197);
and U28942 (N_28942,N_18131,N_22065);
nor U28943 (N_28943,N_21153,N_22426);
nor U28944 (N_28944,N_19446,N_23922);
and U28945 (N_28945,N_21358,N_19124);
nor U28946 (N_28946,N_18063,N_21514);
or U28947 (N_28947,N_19365,N_23081);
and U28948 (N_28948,N_23409,N_20245);
xnor U28949 (N_28949,N_23248,N_22015);
and U28950 (N_28950,N_20874,N_20294);
nor U28951 (N_28951,N_23601,N_23605);
and U28952 (N_28952,N_18158,N_22510);
and U28953 (N_28953,N_19305,N_22776);
nand U28954 (N_28954,N_19352,N_22637);
and U28955 (N_28955,N_18675,N_18686);
or U28956 (N_28956,N_20268,N_18408);
xnor U28957 (N_28957,N_20649,N_20506);
nand U28958 (N_28958,N_22675,N_18667);
xnor U28959 (N_28959,N_21105,N_22364);
and U28960 (N_28960,N_23390,N_23516);
nand U28961 (N_28961,N_18409,N_23528);
and U28962 (N_28962,N_21376,N_22137);
and U28963 (N_28963,N_20966,N_21721);
and U28964 (N_28964,N_19457,N_22752);
xnor U28965 (N_28965,N_20254,N_21492);
nand U28966 (N_28966,N_22373,N_20713);
and U28967 (N_28967,N_23394,N_22835);
nor U28968 (N_28968,N_20400,N_23622);
and U28969 (N_28969,N_18924,N_19434);
nor U28970 (N_28970,N_20750,N_23355);
and U28971 (N_28971,N_22948,N_19983);
nor U28972 (N_28972,N_18568,N_18050);
and U28973 (N_28973,N_18205,N_21647);
nor U28974 (N_28974,N_22107,N_20861);
or U28975 (N_28975,N_21389,N_18469);
xnor U28976 (N_28976,N_22585,N_21811);
nand U28977 (N_28977,N_18892,N_21765);
nand U28978 (N_28978,N_18055,N_21915);
xor U28979 (N_28979,N_22048,N_23251);
and U28980 (N_28980,N_18195,N_21630);
and U28981 (N_28981,N_22114,N_23484);
and U28982 (N_28982,N_18179,N_23667);
and U28983 (N_28983,N_21776,N_23776);
xnor U28984 (N_28984,N_19644,N_18010);
xor U28985 (N_28985,N_18558,N_23587);
xor U28986 (N_28986,N_18085,N_22606);
nand U28987 (N_28987,N_18482,N_20280);
nor U28988 (N_28988,N_18186,N_23807);
or U28989 (N_28989,N_22279,N_23740);
and U28990 (N_28990,N_18114,N_19169);
nor U28991 (N_28991,N_23422,N_23963);
or U28992 (N_28992,N_18801,N_23659);
xnor U28993 (N_28993,N_18280,N_19320);
nor U28994 (N_28994,N_22506,N_22048);
and U28995 (N_28995,N_23338,N_18448);
nand U28996 (N_28996,N_19776,N_23586);
nor U28997 (N_28997,N_22531,N_23445);
nor U28998 (N_28998,N_22217,N_22875);
nor U28999 (N_28999,N_21517,N_21594);
or U29000 (N_29000,N_19966,N_21483);
nor U29001 (N_29001,N_18089,N_19643);
and U29002 (N_29002,N_19512,N_21013);
nand U29003 (N_29003,N_23971,N_19295);
or U29004 (N_29004,N_23803,N_18837);
and U29005 (N_29005,N_18632,N_23506);
xor U29006 (N_29006,N_18793,N_20195);
nand U29007 (N_29007,N_19889,N_18440);
and U29008 (N_29008,N_20404,N_21140);
xor U29009 (N_29009,N_19675,N_18937);
xor U29010 (N_29010,N_20236,N_23998);
nor U29011 (N_29011,N_21719,N_21202);
and U29012 (N_29012,N_19363,N_19002);
nor U29013 (N_29013,N_20937,N_22736);
nor U29014 (N_29014,N_22486,N_23145);
or U29015 (N_29015,N_20869,N_21705);
nor U29016 (N_29016,N_18762,N_20238);
and U29017 (N_29017,N_23597,N_23478);
or U29018 (N_29018,N_19319,N_20810);
or U29019 (N_29019,N_18474,N_18582);
xnor U29020 (N_29020,N_20933,N_20665);
nor U29021 (N_29021,N_20791,N_19921);
nor U29022 (N_29022,N_20707,N_23317);
xor U29023 (N_29023,N_19432,N_19116);
and U29024 (N_29024,N_20416,N_23133);
nor U29025 (N_29025,N_22912,N_18449);
or U29026 (N_29026,N_23835,N_19039);
xnor U29027 (N_29027,N_22614,N_20640);
xnor U29028 (N_29028,N_23608,N_22621);
nand U29029 (N_29029,N_19884,N_19281);
nand U29030 (N_29030,N_21435,N_21207);
or U29031 (N_29031,N_21869,N_22018);
and U29032 (N_29032,N_21866,N_22533);
nand U29033 (N_29033,N_18577,N_22111);
xnor U29034 (N_29034,N_19296,N_20896);
and U29035 (N_29035,N_19382,N_21887);
or U29036 (N_29036,N_23394,N_21007);
or U29037 (N_29037,N_18216,N_22886);
or U29038 (N_29038,N_22664,N_22997);
and U29039 (N_29039,N_20391,N_22370);
nand U29040 (N_29040,N_23113,N_22887);
xnor U29041 (N_29041,N_19686,N_23285);
or U29042 (N_29042,N_21417,N_22213);
and U29043 (N_29043,N_21681,N_23034);
nor U29044 (N_29044,N_22795,N_18981);
nand U29045 (N_29045,N_19080,N_21504);
nor U29046 (N_29046,N_22269,N_19677);
xnor U29047 (N_29047,N_23957,N_19908);
nand U29048 (N_29048,N_23819,N_22538);
nand U29049 (N_29049,N_20981,N_20378);
or U29050 (N_29050,N_20260,N_18718);
nand U29051 (N_29051,N_20047,N_23924);
nor U29052 (N_29052,N_19924,N_18947);
nor U29053 (N_29053,N_22905,N_22316);
or U29054 (N_29054,N_22367,N_23855);
nand U29055 (N_29055,N_19116,N_20038);
or U29056 (N_29056,N_21809,N_21556);
nand U29057 (N_29057,N_23407,N_23964);
nor U29058 (N_29058,N_19227,N_21547);
xor U29059 (N_29059,N_18231,N_18252);
nand U29060 (N_29060,N_21120,N_20663);
nor U29061 (N_29061,N_22515,N_21103);
or U29062 (N_29062,N_21096,N_20955);
nor U29063 (N_29063,N_22355,N_18335);
nor U29064 (N_29064,N_21669,N_21231);
nand U29065 (N_29065,N_20950,N_22107);
or U29066 (N_29066,N_19956,N_23088);
nand U29067 (N_29067,N_20711,N_19162);
nand U29068 (N_29068,N_18987,N_19959);
nor U29069 (N_29069,N_22876,N_18097);
xnor U29070 (N_29070,N_19031,N_20617);
xor U29071 (N_29071,N_20899,N_19498);
or U29072 (N_29072,N_23405,N_20698);
nand U29073 (N_29073,N_20853,N_23608);
xor U29074 (N_29074,N_20147,N_18583);
nand U29075 (N_29075,N_23730,N_20649);
xnor U29076 (N_29076,N_23733,N_19438);
and U29077 (N_29077,N_22256,N_23439);
nand U29078 (N_29078,N_23025,N_22476);
or U29079 (N_29079,N_22047,N_21260);
or U29080 (N_29080,N_21519,N_18698);
xor U29081 (N_29081,N_23979,N_22573);
nor U29082 (N_29082,N_22102,N_19626);
nor U29083 (N_29083,N_22259,N_20929);
or U29084 (N_29084,N_23687,N_22063);
xor U29085 (N_29085,N_21683,N_19887);
nand U29086 (N_29086,N_20116,N_22640);
or U29087 (N_29087,N_21866,N_20528);
nor U29088 (N_29088,N_21479,N_18920);
or U29089 (N_29089,N_21308,N_21114);
or U29090 (N_29090,N_20392,N_19180);
nor U29091 (N_29091,N_22829,N_23169);
xnor U29092 (N_29092,N_18525,N_21217);
nor U29093 (N_29093,N_19024,N_18965);
or U29094 (N_29094,N_21107,N_19204);
xnor U29095 (N_29095,N_18218,N_22533);
nor U29096 (N_29096,N_23176,N_18500);
and U29097 (N_29097,N_23698,N_21531);
nand U29098 (N_29098,N_21152,N_20680);
and U29099 (N_29099,N_18428,N_23480);
nand U29100 (N_29100,N_22506,N_21217);
xnor U29101 (N_29101,N_20992,N_21479);
nand U29102 (N_29102,N_21857,N_20542);
nand U29103 (N_29103,N_19178,N_19230);
nand U29104 (N_29104,N_20423,N_19604);
and U29105 (N_29105,N_22465,N_19329);
nand U29106 (N_29106,N_21230,N_22666);
or U29107 (N_29107,N_21525,N_19936);
and U29108 (N_29108,N_20049,N_23349);
and U29109 (N_29109,N_20134,N_19088);
xor U29110 (N_29110,N_22348,N_20143);
and U29111 (N_29111,N_23788,N_19619);
and U29112 (N_29112,N_19988,N_23612);
nand U29113 (N_29113,N_18447,N_20155);
xor U29114 (N_29114,N_21236,N_18236);
nor U29115 (N_29115,N_19952,N_23221);
and U29116 (N_29116,N_21258,N_18688);
and U29117 (N_29117,N_23522,N_23503);
and U29118 (N_29118,N_19516,N_21781);
or U29119 (N_29119,N_23708,N_21474);
and U29120 (N_29120,N_18995,N_23973);
nand U29121 (N_29121,N_20419,N_20569);
nand U29122 (N_29122,N_20272,N_21567);
or U29123 (N_29123,N_20600,N_21048);
and U29124 (N_29124,N_23608,N_23343);
and U29125 (N_29125,N_19015,N_23304);
nor U29126 (N_29126,N_19115,N_22041);
and U29127 (N_29127,N_20227,N_19473);
nand U29128 (N_29128,N_21914,N_21449);
xor U29129 (N_29129,N_19442,N_18215);
and U29130 (N_29130,N_20855,N_20008);
nand U29131 (N_29131,N_18452,N_22937);
xor U29132 (N_29132,N_21024,N_18541);
and U29133 (N_29133,N_20905,N_23863);
and U29134 (N_29134,N_19010,N_19716);
and U29135 (N_29135,N_19426,N_19040);
xnor U29136 (N_29136,N_23438,N_20441);
nor U29137 (N_29137,N_19410,N_23603);
nand U29138 (N_29138,N_18936,N_21932);
nand U29139 (N_29139,N_23144,N_22801);
nand U29140 (N_29140,N_21033,N_22468);
xnor U29141 (N_29141,N_20437,N_21127);
nand U29142 (N_29142,N_18450,N_20919);
nor U29143 (N_29143,N_21346,N_20733);
nand U29144 (N_29144,N_22048,N_19229);
nand U29145 (N_29145,N_20770,N_20624);
nand U29146 (N_29146,N_18561,N_22030);
or U29147 (N_29147,N_22079,N_23582);
nand U29148 (N_29148,N_21488,N_20439);
or U29149 (N_29149,N_18553,N_23960);
and U29150 (N_29150,N_22914,N_21348);
nor U29151 (N_29151,N_18534,N_21712);
xor U29152 (N_29152,N_18492,N_19506);
or U29153 (N_29153,N_19404,N_18078);
or U29154 (N_29154,N_18421,N_18675);
nand U29155 (N_29155,N_20331,N_21723);
nor U29156 (N_29156,N_18169,N_23639);
nand U29157 (N_29157,N_18246,N_18933);
or U29158 (N_29158,N_22463,N_23245);
and U29159 (N_29159,N_20389,N_21720);
and U29160 (N_29160,N_21075,N_21865);
xor U29161 (N_29161,N_22986,N_20328);
nor U29162 (N_29162,N_19828,N_19629);
and U29163 (N_29163,N_19362,N_23893);
nor U29164 (N_29164,N_22339,N_23002);
xor U29165 (N_29165,N_19425,N_21705);
or U29166 (N_29166,N_22941,N_19197);
or U29167 (N_29167,N_20460,N_23354);
and U29168 (N_29168,N_22878,N_19798);
or U29169 (N_29169,N_21924,N_20214);
xor U29170 (N_29170,N_22997,N_22280);
nand U29171 (N_29171,N_22426,N_22781);
nand U29172 (N_29172,N_22404,N_22554);
or U29173 (N_29173,N_22776,N_22611);
xnor U29174 (N_29174,N_18328,N_19676);
nor U29175 (N_29175,N_18700,N_19784);
xnor U29176 (N_29176,N_19758,N_23318);
nor U29177 (N_29177,N_23274,N_21419);
nand U29178 (N_29178,N_18201,N_20797);
and U29179 (N_29179,N_23890,N_19685);
or U29180 (N_29180,N_20816,N_20434);
nor U29181 (N_29181,N_18317,N_18702);
and U29182 (N_29182,N_21984,N_21814);
xnor U29183 (N_29183,N_20421,N_18283);
nor U29184 (N_29184,N_19265,N_20933);
and U29185 (N_29185,N_20900,N_18417);
and U29186 (N_29186,N_19200,N_23129);
and U29187 (N_29187,N_18315,N_23408);
nor U29188 (N_29188,N_21633,N_23093);
or U29189 (N_29189,N_18703,N_20292);
nand U29190 (N_29190,N_23124,N_18513);
and U29191 (N_29191,N_21560,N_23088);
xnor U29192 (N_29192,N_18783,N_19164);
and U29193 (N_29193,N_21590,N_19494);
and U29194 (N_29194,N_23476,N_21794);
nand U29195 (N_29195,N_21658,N_18945);
nand U29196 (N_29196,N_18142,N_23755);
or U29197 (N_29197,N_21453,N_22316);
xnor U29198 (N_29198,N_18326,N_20347);
nand U29199 (N_29199,N_20460,N_19038);
or U29200 (N_29200,N_19623,N_23353);
or U29201 (N_29201,N_21859,N_23877);
xnor U29202 (N_29202,N_20254,N_22303);
nand U29203 (N_29203,N_22590,N_20202);
xnor U29204 (N_29204,N_21290,N_22518);
and U29205 (N_29205,N_22942,N_19935);
nor U29206 (N_29206,N_19660,N_20048);
xnor U29207 (N_29207,N_22706,N_23249);
xor U29208 (N_29208,N_22574,N_19023);
and U29209 (N_29209,N_18279,N_19599);
xnor U29210 (N_29210,N_19229,N_20191);
nand U29211 (N_29211,N_21026,N_18011);
nand U29212 (N_29212,N_20339,N_19626);
or U29213 (N_29213,N_18703,N_21119);
nand U29214 (N_29214,N_18886,N_18566);
and U29215 (N_29215,N_20860,N_23699);
nor U29216 (N_29216,N_23651,N_19638);
or U29217 (N_29217,N_19858,N_19146);
nand U29218 (N_29218,N_18536,N_20347);
nand U29219 (N_29219,N_18633,N_20761);
nor U29220 (N_29220,N_18971,N_23788);
nor U29221 (N_29221,N_21784,N_18707);
xor U29222 (N_29222,N_19607,N_23178);
and U29223 (N_29223,N_20798,N_23098);
and U29224 (N_29224,N_18304,N_23885);
nor U29225 (N_29225,N_18552,N_19244);
or U29226 (N_29226,N_23610,N_19485);
and U29227 (N_29227,N_23340,N_21948);
or U29228 (N_29228,N_21595,N_23941);
or U29229 (N_29229,N_19244,N_20170);
nand U29230 (N_29230,N_22656,N_19773);
and U29231 (N_29231,N_20482,N_20337);
xnor U29232 (N_29232,N_23310,N_19743);
xor U29233 (N_29233,N_23678,N_20455);
and U29234 (N_29234,N_18935,N_21125);
or U29235 (N_29235,N_21873,N_20719);
nor U29236 (N_29236,N_19422,N_22935);
xnor U29237 (N_29237,N_19347,N_20181);
nand U29238 (N_29238,N_23358,N_22221);
xor U29239 (N_29239,N_18927,N_21940);
xnor U29240 (N_29240,N_18952,N_19284);
nand U29241 (N_29241,N_22762,N_21729);
nor U29242 (N_29242,N_23490,N_21898);
or U29243 (N_29243,N_20185,N_21643);
xor U29244 (N_29244,N_23848,N_19448);
and U29245 (N_29245,N_20338,N_23615);
nand U29246 (N_29246,N_19731,N_22021);
xor U29247 (N_29247,N_18388,N_18041);
or U29248 (N_29248,N_19028,N_19142);
nand U29249 (N_29249,N_23151,N_22535);
nand U29250 (N_29250,N_21114,N_20748);
nand U29251 (N_29251,N_22700,N_23808);
and U29252 (N_29252,N_20001,N_23599);
nor U29253 (N_29253,N_22690,N_19975);
and U29254 (N_29254,N_22363,N_21069);
xnor U29255 (N_29255,N_18344,N_18590);
nor U29256 (N_29256,N_20989,N_19581);
xnor U29257 (N_29257,N_20168,N_21759);
and U29258 (N_29258,N_21529,N_20414);
and U29259 (N_29259,N_18978,N_21821);
and U29260 (N_29260,N_21568,N_23620);
xnor U29261 (N_29261,N_22928,N_23890);
nand U29262 (N_29262,N_20062,N_18477);
nor U29263 (N_29263,N_22011,N_22222);
and U29264 (N_29264,N_23424,N_19427);
or U29265 (N_29265,N_19245,N_23874);
or U29266 (N_29266,N_18211,N_18292);
xnor U29267 (N_29267,N_23621,N_19817);
nand U29268 (N_29268,N_19178,N_20916);
or U29269 (N_29269,N_22408,N_18077);
nor U29270 (N_29270,N_18777,N_19552);
nor U29271 (N_29271,N_19086,N_21338);
or U29272 (N_29272,N_19364,N_21622);
or U29273 (N_29273,N_19275,N_23138);
or U29274 (N_29274,N_20709,N_19443);
or U29275 (N_29275,N_22148,N_20376);
nor U29276 (N_29276,N_22753,N_19390);
xor U29277 (N_29277,N_18117,N_21887);
or U29278 (N_29278,N_18068,N_19609);
or U29279 (N_29279,N_18489,N_18922);
and U29280 (N_29280,N_18209,N_21741);
xor U29281 (N_29281,N_21936,N_19473);
or U29282 (N_29282,N_22196,N_23452);
or U29283 (N_29283,N_23325,N_21924);
xnor U29284 (N_29284,N_23085,N_22222);
xor U29285 (N_29285,N_18817,N_23656);
and U29286 (N_29286,N_18382,N_18423);
and U29287 (N_29287,N_20680,N_22022);
xnor U29288 (N_29288,N_22579,N_23401);
or U29289 (N_29289,N_19049,N_19317);
xnor U29290 (N_29290,N_21288,N_19668);
or U29291 (N_29291,N_21930,N_23095);
xor U29292 (N_29292,N_20910,N_18523);
nor U29293 (N_29293,N_23008,N_21696);
xor U29294 (N_29294,N_18955,N_18848);
nand U29295 (N_29295,N_23764,N_18907);
and U29296 (N_29296,N_23889,N_21270);
xnor U29297 (N_29297,N_19691,N_22892);
xnor U29298 (N_29298,N_21904,N_23080);
nor U29299 (N_29299,N_18143,N_23880);
or U29300 (N_29300,N_22122,N_23446);
or U29301 (N_29301,N_21627,N_19859);
xnor U29302 (N_29302,N_20236,N_21011);
nor U29303 (N_29303,N_18288,N_18164);
and U29304 (N_29304,N_20343,N_23402);
and U29305 (N_29305,N_20552,N_23882);
nor U29306 (N_29306,N_21092,N_20147);
nor U29307 (N_29307,N_21031,N_19277);
xnor U29308 (N_29308,N_19654,N_18655);
nand U29309 (N_29309,N_19267,N_22569);
or U29310 (N_29310,N_18154,N_21683);
nor U29311 (N_29311,N_23411,N_19788);
or U29312 (N_29312,N_21843,N_22969);
nor U29313 (N_29313,N_23704,N_18113);
xnor U29314 (N_29314,N_22161,N_22140);
or U29315 (N_29315,N_22164,N_18986);
or U29316 (N_29316,N_18063,N_21632);
and U29317 (N_29317,N_18059,N_20665);
xnor U29318 (N_29318,N_20427,N_22515);
nor U29319 (N_29319,N_23946,N_22219);
nand U29320 (N_29320,N_19099,N_20049);
or U29321 (N_29321,N_23103,N_21433);
or U29322 (N_29322,N_22247,N_22112);
and U29323 (N_29323,N_18768,N_18987);
nor U29324 (N_29324,N_21327,N_19488);
nor U29325 (N_29325,N_18026,N_20388);
or U29326 (N_29326,N_19096,N_22034);
and U29327 (N_29327,N_21265,N_19313);
xnor U29328 (N_29328,N_23168,N_23663);
nor U29329 (N_29329,N_20148,N_20075);
or U29330 (N_29330,N_20504,N_19378);
nand U29331 (N_29331,N_21969,N_22457);
nor U29332 (N_29332,N_21585,N_18914);
nand U29333 (N_29333,N_22355,N_21347);
xnor U29334 (N_29334,N_19383,N_22292);
and U29335 (N_29335,N_22521,N_23025);
xor U29336 (N_29336,N_21258,N_19639);
or U29337 (N_29337,N_18008,N_22990);
or U29338 (N_29338,N_20060,N_20031);
nor U29339 (N_29339,N_18253,N_23061);
nand U29340 (N_29340,N_21936,N_18467);
xor U29341 (N_29341,N_22730,N_20418);
nor U29342 (N_29342,N_20779,N_22434);
or U29343 (N_29343,N_22941,N_20235);
xor U29344 (N_29344,N_22712,N_21590);
or U29345 (N_29345,N_23584,N_20261);
and U29346 (N_29346,N_22475,N_21859);
or U29347 (N_29347,N_23177,N_19126);
nor U29348 (N_29348,N_23565,N_19257);
nand U29349 (N_29349,N_22411,N_19336);
nor U29350 (N_29350,N_22336,N_23666);
nand U29351 (N_29351,N_22181,N_18414);
xnor U29352 (N_29352,N_23731,N_18586);
or U29353 (N_29353,N_22482,N_21011);
nand U29354 (N_29354,N_18455,N_22146);
nor U29355 (N_29355,N_21794,N_18071);
nand U29356 (N_29356,N_22004,N_22984);
or U29357 (N_29357,N_21786,N_21465);
nand U29358 (N_29358,N_23941,N_21443);
nand U29359 (N_29359,N_21161,N_21074);
xor U29360 (N_29360,N_23075,N_18638);
xor U29361 (N_29361,N_20061,N_20436);
nand U29362 (N_29362,N_21299,N_21144);
xnor U29363 (N_29363,N_22391,N_20872);
nand U29364 (N_29364,N_23388,N_20062);
or U29365 (N_29365,N_22485,N_19832);
or U29366 (N_29366,N_20344,N_18566);
nor U29367 (N_29367,N_19444,N_19996);
and U29368 (N_29368,N_19192,N_20250);
or U29369 (N_29369,N_18581,N_20374);
nand U29370 (N_29370,N_23332,N_21450);
nand U29371 (N_29371,N_20708,N_20243);
xor U29372 (N_29372,N_20109,N_21423);
xor U29373 (N_29373,N_23823,N_21550);
and U29374 (N_29374,N_22411,N_22581);
or U29375 (N_29375,N_23475,N_18604);
and U29376 (N_29376,N_19875,N_20101);
xnor U29377 (N_29377,N_23780,N_18567);
nor U29378 (N_29378,N_23754,N_18102);
xnor U29379 (N_29379,N_22706,N_22153);
xnor U29380 (N_29380,N_20716,N_22886);
or U29381 (N_29381,N_22976,N_18599);
xnor U29382 (N_29382,N_21393,N_23006);
xor U29383 (N_29383,N_19242,N_23791);
nor U29384 (N_29384,N_20914,N_22966);
nor U29385 (N_29385,N_20645,N_22895);
xnor U29386 (N_29386,N_20291,N_18432);
nand U29387 (N_29387,N_20999,N_18849);
nand U29388 (N_29388,N_18556,N_18820);
nor U29389 (N_29389,N_18380,N_22345);
or U29390 (N_29390,N_23760,N_21737);
and U29391 (N_29391,N_19551,N_23828);
or U29392 (N_29392,N_18800,N_19285);
nand U29393 (N_29393,N_20141,N_21816);
nor U29394 (N_29394,N_21327,N_20273);
or U29395 (N_29395,N_18683,N_23711);
xor U29396 (N_29396,N_20050,N_22927);
nand U29397 (N_29397,N_20564,N_19229);
nand U29398 (N_29398,N_20035,N_22029);
or U29399 (N_29399,N_23201,N_20312);
xnor U29400 (N_29400,N_23938,N_20972);
nor U29401 (N_29401,N_18937,N_19135);
nand U29402 (N_29402,N_19148,N_23695);
nand U29403 (N_29403,N_19301,N_18096);
nor U29404 (N_29404,N_21035,N_21159);
nor U29405 (N_29405,N_20418,N_23772);
or U29406 (N_29406,N_23880,N_18583);
nor U29407 (N_29407,N_21371,N_19030);
or U29408 (N_29408,N_23746,N_19787);
xnor U29409 (N_29409,N_23417,N_21729);
nor U29410 (N_29410,N_19877,N_22619);
nor U29411 (N_29411,N_21303,N_21638);
nand U29412 (N_29412,N_22105,N_19739);
xnor U29413 (N_29413,N_23582,N_21345);
or U29414 (N_29414,N_22107,N_22347);
or U29415 (N_29415,N_20626,N_18013);
xnor U29416 (N_29416,N_18058,N_21700);
and U29417 (N_29417,N_18847,N_18394);
nand U29418 (N_29418,N_19428,N_23939);
xor U29419 (N_29419,N_23430,N_20311);
nand U29420 (N_29420,N_22582,N_19709);
xnor U29421 (N_29421,N_18602,N_21528);
and U29422 (N_29422,N_20217,N_18311);
nor U29423 (N_29423,N_18041,N_20735);
nor U29424 (N_29424,N_18686,N_23036);
xnor U29425 (N_29425,N_18911,N_22758);
or U29426 (N_29426,N_18481,N_23642);
or U29427 (N_29427,N_20220,N_20503);
nor U29428 (N_29428,N_19199,N_19874);
and U29429 (N_29429,N_22110,N_19832);
nand U29430 (N_29430,N_22797,N_22456);
and U29431 (N_29431,N_21411,N_19110);
or U29432 (N_29432,N_23927,N_20573);
or U29433 (N_29433,N_20088,N_20615);
nor U29434 (N_29434,N_23016,N_20848);
and U29435 (N_29435,N_20574,N_21344);
or U29436 (N_29436,N_19040,N_22564);
or U29437 (N_29437,N_23667,N_19326);
xnor U29438 (N_29438,N_22586,N_19837);
or U29439 (N_29439,N_18321,N_22148);
or U29440 (N_29440,N_19183,N_23980);
nor U29441 (N_29441,N_20071,N_20441);
nor U29442 (N_29442,N_18688,N_19099);
nor U29443 (N_29443,N_22917,N_23614);
nand U29444 (N_29444,N_22210,N_19964);
nor U29445 (N_29445,N_19248,N_20006);
nor U29446 (N_29446,N_21165,N_19637);
nand U29447 (N_29447,N_19327,N_20925);
or U29448 (N_29448,N_18290,N_21718);
nand U29449 (N_29449,N_18739,N_23813);
nand U29450 (N_29450,N_18706,N_21219);
xor U29451 (N_29451,N_18007,N_19605);
or U29452 (N_29452,N_18327,N_18782);
xnor U29453 (N_29453,N_19804,N_22203);
nand U29454 (N_29454,N_23637,N_20183);
nor U29455 (N_29455,N_23339,N_22724);
nand U29456 (N_29456,N_19424,N_19348);
or U29457 (N_29457,N_20208,N_23449);
nand U29458 (N_29458,N_22542,N_21386);
and U29459 (N_29459,N_19585,N_21664);
xnor U29460 (N_29460,N_22372,N_18269);
and U29461 (N_29461,N_21767,N_18599);
xnor U29462 (N_29462,N_20161,N_19149);
nand U29463 (N_29463,N_21130,N_20460);
nand U29464 (N_29464,N_20454,N_22103);
nand U29465 (N_29465,N_22950,N_20305);
nand U29466 (N_29466,N_19238,N_20677);
nand U29467 (N_29467,N_20771,N_22564);
and U29468 (N_29468,N_20204,N_18763);
or U29469 (N_29469,N_18413,N_20578);
or U29470 (N_29470,N_19748,N_20723);
or U29471 (N_29471,N_21951,N_18682);
nand U29472 (N_29472,N_20507,N_21753);
or U29473 (N_29473,N_19449,N_19694);
nor U29474 (N_29474,N_23613,N_23194);
or U29475 (N_29475,N_19532,N_21920);
xnor U29476 (N_29476,N_21564,N_20633);
and U29477 (N_29477,N_22292,N_20575);
or U29478 (N_29478,N_23359,N_20792);
nand U29479 (N_29479,N_21477,N_21206);
nor U29480 (N_29480,N_23328,N_21843);
xnor U29481 (N_29481,N_19367,N_21518);
xor U29482 (N_29482,N_22907,N_23987);
or U29483 (N_29483,N_20244,N_22290);
or U29484 (N_29484,N_19271,N_19026);
xnor U29485 (N_29485,N_22603,N_20344);
nand U29486 (N_29486,N_21292,N_21545);
or U29487 (N_29487,N_19404,N_21499);
xnor U29488 (N_29488,N_22290,N_23765);
xor U29489 (N_29489,N_20034,N_18656);
or U29490 (N_29490,N_18843,N_20212);
nor U29491 (N_29491,N_20273,N_22577);
nand U29492 (N_29492,N_21569,N_20702);
xnor U29493 (N_29493,N_21309,N_23166);
xnor U29494 (N_29494,N_22759,N_18652);
nor U29495 (N_29495,N_22907,N_21726);
and U29496 (N_29496,N_18369,N_22984);
xor U29497 (N_29497,N_22256,N_22963);
or U29498 (N_29498,N_20503,N_22100);
xnor U29499 (N_29499,N_20662,N_21638);
nand U29500 (N_29500,N_23394,N_18044);
xnor U29501 (N_29501,N_21945,N_23991);
and U29502 (N_29502,N_23591,N_19157);
xnor U29503 (N_29503,N_20669,N_19208);
nor U29504 (N_29504,N_18016,N_19875);
or U29505 (N_29505,N_23731,N_20420);
nand U29506 (N_29506,N_19518,N_20995);
or U29507 (N_29507,N_21986,N_18050);
nor U29508 (N_29508,N_21355,N_22977);
and U29509 (N_29509,N_20711,N_23421);
xnor U29510 (N_29510,N_22100,N_18561);
nor U29511 (N_29511,N_18234,N_21580);
nor U29512 (N_29512,N_23569,N_20797);
nand U29513 (N_29513,N_20933,N_23241);
nand U29514 (N_29514,N_22856,N_20174);
xnor U29515 (N_29515,N_23058,N_21010);
nor U29516 (N_29516,N_18421,N_19098);
xnor U29517 (N_29517,N_18490,N_21988);
nand U29518 (N_29518,N_21886,N_20621);
xnor U29519 (N_29519,N_23161,N_19226);
xor U29520 (N_29520,N_22183,N_21163);
or U29521 (N_29521,N_23696,N_20074);
and U29522 (N_29522,N_21893,N_18193);
or U29523 (N_29523,N_23069,N_20780);
xor U29524 (N_29524,N_18615,N_19588);
nor U29525 (N_29525,N_20057,N_19118);
and U29526 (N_29526,N_18578,N_22729);
and U29527 (N_29527,N_19757,N_21127);
and U29528 (N_29528,N_18805,N_22124);
or U29529 (N_29529,N_21183,N_20686);
xnor U29530 (N_29530,N_18812,N_20848);
and U29531 (N_29531,N_19496,N_23452);
and U29532 (N_29532,N_21637,N_22010);
nor U29533 (N_29533,N_18418,N_20377);
xnor U29534 (N_29534,N_18865,N_18324);
xnor U29535 (N_29535,N_20927,N_21213);
nor U29536 (N_29536,N_23598,N_23979);
or U29537 (N_29537,N_18422,N_23987);
or U29538 (N_29538,N_20667,N_21750);
nor U29539 (N_29539,N_19083,N_20473);
nor U29540 (N_29540,N_19494,N_19543);
and U29541 (N_29541,N_20401,N_21545);
nand U29542 (N_29542,N_20462,N_21106);
xnor U29543 (N_29543,N_19738,N_20327);
and U29544 (N_29544,N_19118,N_22633);
nor U29545 (N_29545,N_19030,N_18439);
or U29546 (N_29546,N_22062,N_19486);
nand U29547 (N_29547,N_23719,N_20948);
nor U29548 (N_29548,N_19993,N_21571);
nor U29549 (N_29549,N_23644,N_20721);
or U29550 (N_29550,N_20116,N_22460);
xnor U29551 (N_29551,N_21909,N_21579);
or U29552 (N_29552,N_22089,N_18329);
nor U29553 (N_29553,N_22316,N_23711);
or U29554 (N_29554,N_23480,N_23209);
xor U29555 (N_29555,N_23025,N_23115);
and U29556 (N_29556,N_23355,N_20607);
or U29557 (N_29557,N_18827,N_18545);
and U29558 (N_29558,N_19951,N_19961);
or U29559 (N_29559,N_21800,N_23900);
xor U29560 (N_29560,N_20904,N_22662);
nor U29561 (N_29561,N_23008,N_21412);
or U29562 (N_29562,N_18623,N_21933);
nand U29563 (N_29563,N_20338,N_22793);
xor U29564 (N_29564,N_18175,N_20247);
and U29565 (N_29565,N_20691,N_18856);
and U29566 (N_29566,N_18484,N_20115);
nor U29567 (N_29567,N_23322,N_19860);
xnor U29568 (N_29568,N_22692,N_22288);
xnor U29569 (N_29569,N_23708,N_21203);
nor U29570 (N_29570,N_18735,N_23323);
and U29571 (N_29571,N_20521,N_21388);
or U29572 (N_29572,N_23353,N_18420);
xnor U29573 (N_29573,N_22597,N_23320);
and U29574 (N_29574,N_23515,N_18827);
nor U29575 (N_29575,N_19752,N_21367);
xnor U29576 (N_29576,N_18002,N_22984);
xor U29577 (N_29577,N_23290,N_19774);
nand U29578 (N_29578,N_19928,N_19715);
and U29579 (N_29579,N_21244,N_23592);
nand U29580 (N_29580,N_23054,N_18519);
and U29581 (N_29581,N_21703,N_19161);
and U29582 (N_29582,N_21807,N_23647);
or U29583 (N_29583,N_22693,N_22877);
nor U29584 (N_29584,N_22255,N_22752);
xnor U29585 (N_29585,N_21363,N_23534);
nor U29586 (N_29586,N_23878,N_23183);
nor U29587 (N_29587,N_22161,N_20544);
and U29588 (N_29588,N_20470,N_18607);
nor U29589 (N_29589,N_20427,N_19514);
or U29590 (N_29590,N_19719,N_23242);
or U29591 (N_29591,N_20923,N_21951);
nor U29592 (N_29592,N_19387,N_21073);
nand U29593 (N_29593,N_22888,N_20093);
nand U29594 (N_29594,N_21751,N_18397);
or U29595 (N_29595,N_18961,N_20370);
and U29596 (N_29596,N_22849,N_20940);
or U29597 (N_29597,N_21113,N_21148);
and U29598 (N_29598,N_21668,N_20349);
nand U29599 (N_29599,N_19681,N_21021);
and U29600 (N_29600,N_23470,N_21098);
or U29601 (N_29601,N_21802,N_18826);
or U29602 (N_29602,N_19713,N_22921);
xor U29603 (N_29603,N_21595,N_21864);
xor U29604 (N_29604,N_20794,N_21518);
xor U29605 (N_29605,N_19819,N_23634);
and U29606 (N_29606,N_23519,N_22674);
xor U29607 (N_29607,N_21481,N_23377);
or U29608 (N_29608,N_21995,N_22132);
and U29609 (N_29609,N_21317,N_22019);
or U29610 (N_29610,N_21680,N_19797);
and U29611 (N_29611,N_21226,N_20164);
and U29612 (N_29612,N_18549,N_19610);
nand U29613 (N_29613,N_19511,N_22359);
and U29614 (N_29614,N_23722,N_21003);
and U29615 (N_29615,N_23784,N_19442);
or U29616 (N_29616,N_19300,N_21357);
nand U29617 (N_29617,N_19285,N_22618);
or U29618 (N_29618,N_20155,N_23344);
xor U29619 (N_29619,N_19273,N_19450);
nor U29620 (N_29620,N_20044,N_18418);
and U29621 (N_29621,N_19815,N_19383);
and U29622 (N_29622,N_20436,N_21533);
xor U29623 (N_29623,N_20475,N_23482);
xor U29624 (N_29624,N_19445,N_21938);
or U29625 (N_29625,N_22450,N_20917);
nand U29626 (N_29626,N_22571,N_23283);
nand U29627 (N_29627,N_22721,N_18527);
nand U29628 (N_29628,N_20020,N_20076);
and U29629 (N_29629,N_23855,N_22072);
or U29630 (N_29630,N_20672,N_23836);
nor U29631 (N_29631,N_21313,N_21773);
and U29632 (N_29632,N_20742,N_21705);
xnor U29633 (N_29633,N_20447,N_21472);
xor U29634 (N_29634,N_19942,N_18633);
xnor U29635 (N_29635,N_22140,N_22636);
or U29636 (N_29636,N_22801,N_22300);
nand U29637 (N_29637,N_19912,N_18847);
and U29638 (N_29638,N_22069,N_19701);
or U29639 (N_29639,N_20207,N_22971);
and U29640 (N_29640,N_22068,N_21140);
xnor U29641 (N_29641,N_21216,N_22910);
or U29642 (N_29642,N_19012,N_21088);
nand U29643 (N_29643,N_19001,N_22677);
and U29644 (N_29644,N_22166,N_21278);
or U29645 (N_29645,N_19837,N_19450);
nand U29646 (N_29646,N_18059,N_23431);
nor U29647 (N_29647,N_20739,N_19643);
nand U29648 (N_29648,N_18280,N_20909);
nand U29649 (N_29649,N_20373,N_19044);
and U29650 (N_29650,N_21547,N_23195);
nor U29651 (N_29651,N_20737,N_20586);
nor U29652 (N_29652,N_18120,N_21121);
xnor U29653 (N_29653,N_23125,N_21441);
nor U29654 (N_29654,N_18774,N_22563);
nor U29655 (N_29655,N_18986,N_23685);
or U29656 (N_29656,N_23672,N_18677);
xnor U29657 (N_29657,N_20817,N_22592);
xor U29658 (N_29658,N_20696,N_22142);
xnor U29659 (N_29659,N_21905,N_23017);
nand U29660 (N_29660,N_20733,N_22055);
nor U29661 (N_29661,N_21832,N_22186);
and U29662 (N_29662,N_19266,N_21579);
and U29663 (N_29663,N_19092,N_21848);
and U29664 (N_29664,N_19277,N_20988);
xnor U29665 (N_29665,N_21329,N_19217);
and U29666 (N_29666,N_23648,N_22922);
xor U29667 (N_29667,N_18826,N_20165);
xor U29668 (N_29668,N_23386,N_20688);
or U29669 (N_29669,N_22592,N_20871);
nor U29670 (N_29670,N_19713,N_19201);
or U29671 (N_29671,N_18750,N_21669);
xor U29672 (N_29672,N_19734,N_21572);
and U29673 (N_29673,N_21809,N_21485);
xor U29674 (N_29674,N_18583,N_21510);
nand U29675 (N_29675,N_22529,N_18178);
nor U29676 (N_29676,N_21941,N_21606);
nand U29677 (N_29677,N_22156,N_19623);
xor U29678 (N_29678,N_18898,N_20815);
nand U29679 (N_29679,N_20111,N_23229);
and U29680 (N_29680,N_21714,N_23263);
xor U29681 (N_29681,N_18004,N_21940);
nand U29682 (N_29682,N_21217,N_23754);
or U29683 (N_29683,N_20899,N_18399);
nand U29684 (N_29684,N_19196,N_22546);
and U29685 (N_29685,N_22912,N_19429);
or U29686 (N_29686,N_20990,N_19061);
xnor U29687 (N_29687,N_19822,N_21835);
and U29688 (N_29688,N_18816,N_22440);
and U29689 (N_29689,N_20141,N_18977);
and U29690 (N_29690,N_22062,N_18125);
or U29691 (N_29691,N_22333,N_19138);
nor U29692 (N_29692,N_21968,N_19657);
and U29693 (N_29693,N_19233,N_19878);
nand U29694 (N_29694,N_18257,N_21783);
nor U29695 (N_29695,N_18163,N_20681);
nor U29696 (N_29696,N_23526,N_18365);
nor U29697 (N_29697,N_22224,N_19518);
nand U29698 (N_29698,N_19504,N_21438);
nor U29699 (N_29699,N_23789,N_23352);
nor U29700 (N_29700,N_19466,N_22439);
xor U29701 (N_29701,N_18823,N_21120);
nor U29702 (N_29702,N_23458,N_19968);
and U29703 (N_29703,N_21692,N_22206);
xor U29704 (N_29704,N_18226,N_23321);
xor U29705 (N_29705,N_22997,N_18629);
and U29706 (N_29706,N_22863,N_23589);
nand U29707 (N_29707,N_20419,N_18449);
nand U29708 (N_29708,N_21294,N_23007);
or U29709 (N_29709,N_21010,N_20101);
or U29710 (N_29710,N_20398,N_18206);
or U29711 (N_29711,N_19748,N_19782);
and U29712 (N_29712,N_22559,N_18760);
and U29713 (N_29713,N_20431,N_18475);
nor U29714 (N_29714,N_20052,N_22238);
or U29715 (N_29715,N_23387,N_22411);
and U29716 (N_29716,N_22119,N_21209);
xnor U29717 (N_29717,N_18191,N_20807);
or U29718 (N_29718,N_21912,N_20367);
xnor U29719 (N_29719,N_18228,N_18150);
or U29720 (N_29720,N_20526,N_19072);
and U29721 (N_29721,N_19826,N_22809);
nand U29722 (N_29722,N_23371,N_23843);
and U29723 (N_29723,N_18515,N_18666);
nor U29724 (N_29724,N_22153,N_23486);
nor U29725 (N_29725,N_21280,N_22137);
nand U29726 (N_29726,N_20934,N_18849);
and U29727 (N_29727,N_18260,N_21548);
xnor U29728 (N_29728,N_19126,N_18306);
nor U29729 (N_29729,N_19835,N_19417);
nand U29730 (N_29730,N_20399,N_22170);
and U29731 (N_29731,N_20175,N_18513);
nor U29732 (N_29732,N_22358,N_19017);
nand U29733 (N_29733,N_23591,N_19657);
xnor U29734 (N_29734,N_22740,N_21989);
and U29735 (N_29735,N_21833,N_18975);
nor U29736 (N_29736,N_22407,N_23375);
or U29737 (N_29737,N_20330,N_19607);
nand U29738 (N_29738,N_21385,N_21274);
nand U29739 (N_29739,N_18569,N_23154);
or U29740 (N_29740,N_21658,N_21063);
and U29741 (N_29741,N_21932,N_18081);
or U29742 (N_29742,N_22174,N_20766);
or U29743 (N_29743,N_18372,N_23635);
xnor U29744 (N_29744,N_20114,N_20806);
nand U29745 (N_29745,N_22681,N_19530);
or U29746 (N_29746,N_22315,N_21074);
nor U29747 (N_29747,N_22038,N_19587);
or U29748 (N_29748,N_22008,N_22042);
or U29749 (N_29749,N_22713,N_20733);
nor U29750 (N_29750,N_18764,N_21526);
nand U29751 (N_29751,N_21386,N_20622);
or U29752 (N_29752,N_21650,N_20534);
nand U29753 (N_29753,N_21003,N_19500);
nand U29754 (N_29754,N_21575,N_18968);
nor U29755 (N_29755,N_18299,N_19240);
nand U29756 (N_29756,N_21051,N_22750);
and U29757 (N_29757,N_19535,N_19195);
nand U29758 (N_29758,N_18553,N_20957);
nor U29759 (N_29759,N_19994,N_19382);
xnor U29760 (N_29760,N_23980,N_23115);
or U29761 (N_29761,N_21096,N_21868);
nor U29762 (N_29762,N_21228,N_22169);
or U29763 (N_29763,N_21847,N_18007);
nand U29764 (N_29764,N_20794,N_19957);
nand U29765 (N_29765,N_20598,N_23023);
or U29766 (N_29766,N_23146,N_19708);
and U29767 (N_29767,N_21807,N_18336);
or U29768 (N_29768,N_23603,N_20196);
and U29769 (N_29769,N_21846,N_18351);
and U29770 (N_29770,N_21741,N_21044);
and U29771 (N_29771,N_20212,N_23162);
or U29772 (N_29772,N_18209,N_22393);
nor U29773 (N_29773,N_22153,N_21309);
and U29774 (N_29774,N_18179,N_20394);
or U29775 (N_29775,N_21880,N_23254);
nor U29776 (N_29776,N_21011,N_20314);
and U29777 (N_29777,N_22158,N_19135);
or U29778 (N_29778,N_21358,N_20720);
or U29779 (N_29779,N_21577,N_18635);
or U29780 (N_29780,N_20575,N_22155);
nand U29781 (N_29781,N_21582,N_23919);
and U29782 (N_29782,N_18722,N_22277);
or U29783 (N_29783,N_21601,N_19175);
xnor U29784 (N_29784,N_19595,N_23925);
or U29785 (N_29785,N_20267,N_20911);
xnor U29786 (N_29786,N_20134,N_18172);
xor U29787 (N_29787,N_21306,N_20842);
xor U29788 (N_29788,N_19918,N_22117);
and U29789 (N_29789,N_20890,N_18389);
or U29790 (N_29790,N_21900,N_20427);
nand U29791 (N_29791,N_22695,N_23047);
xnor U29792 (N_29792,N_20141,N_19276);
nand U29793 (N_29793,N_21165,N_23021);
xor U29794 (N_29794,N_23993,N_23862);
and U29795 (N_29795,N_19039,N_20073);
or U29796 (N_29796,N_23241,N_22478);
xor U29797 (N_29797,N_18715,N_18404);
nor U29798 (N_29798,N_19900,N_23701);
nand U29799 (N_29799,N_23470,N_19267);
nor U29800 (N_29800,N_22630,N_23843);
nor U29801 (N_29801,N_21647,N_21274);
and U29802 (N_29802,N_23214,N_20111);
nor U29803 (N_29803,N_19227,N_21844);
nand U29804 (N_29804,N_21516,N_21801);
xor U29805 (N_29805,N_22388,N_19403);
nand U29806 (N_29806,N_18016,N_23069);
and U29807 (N_29807,N_23273,N_19234);
xor U29808 (N_29808,N_23163,N_20678);
nand U29809 (N_29809,N_22068,N_23465);
xor U29810 (N_29810,N_18807,N_19435);
nor U29811 (N_29811,N_20849,N_18587);
and U29812 (N_29812,N_20605,N_20770);
xor U29813 (N_29813,N_23742,N_19563);
nand U29814 (N_29814,N_22826,N_23602);
and U29815 (N_29815,N_19433,N_23071);
xnor U29816 (N_29816,N_18275,N_19995);
nand U29817 (N_29817,N_19512,N_20393);
xor U29818 (N_29818,N_19075,N_23928);
xnor U29819 (N_29819,N_23091,N_18205);
nand U29820 (N_29820,N_20391,N_23820);
nor U29821 (N_29821,N_18063,N_22751);
nand U29822 (N_29822,N_22293,N_23992);
nor U29823 (N_29823,N_21931,N_20013);
xnor U29824 (N_29824,N_21995,N_19075);
nand U29825 (N_29825,N_23344,N_19839);
and U29826 (N_29826,N_22265,N_23560);
or U29827 (N_29827,N_18930,N_23631);
and U29828 (N_29828,N_22461,N_18828);
nor U29829 (N_29829,N_19274,N_22356);
or U29830 (N_29830,N_23180,N_20723);
or U29831 (N_29831,N_21482,N_22916);
or U29832 (N_29832,N_23761,N_23442);
nand U29833 (N_29833,N_21091,N_19712);
nor U29834 (N_29834,N_19168,N_21359);
or U29835 (N_29835,N_19956,N_23817);
and U29836 (N_29836,N_20038,N_22475);
and U29837 (N_29837,N_20808,N_19791);
and U29838 (N_29838,N_18594,N_18513);
or U29839 (N_29839,N_18074,N_22110);
xnor U29840 (N_29840,N_19228,N_19803);
nor U29841 (N_29841,N_22120,N_21187);
nand U29842 (N_29842,N_21076,N_20990);
nand U29843 (N_29843,N_23316,N_21886);
nand U29844 (N_29844,N_22788,N_20429);
or U29845 (N_29845,N_22560,N_19291);
or U29846 (N_29846,N_20328,N_23947);
and U29847 (N_29847,N_19964,N_18111);
xnor U29848 (N_29848,N_18671,N_21330);
nor U29849 (N_29849,N_20137,N_19668);
nor U29850 (N_29850,N_19722,N_20134);
or U29851 (N_29851,N_19155,N_20647);
xor U29852 (N_29852,N_20431,N_19286);
xnor U29853 (N_29853,N_23396,N_18790);
and U29854 (N_29854,N_20005,N_20169);
xor U29855 (N_29855,N_20625,N_23601);
nand U29856 (N_29856,N_19803,N_19862);
nand U29857 (N_29857,N_21054,N_18677);
nor U29858 (N_29858,N_18889,N_23365);
nor U29859 (N_29859,N_23610,N_18512);
nor U29860 (N_29860,N_19993,N_19971);
and U29861 (N_29861,N_22410,N_20520);
and U29862 (N_29862,N_18978,N_21142);
nand U29863 (N_29863,N_22491,N_18522);
nand U29864 (N_29864,N_20455,N_21919);
xor U29865 (N_29865,N_19133,N_20952);
xor U29866 (N_29866,N_19982,N_19946);
nor U29867 (N_29867,N_18722,N_21138);
nor U29868 (N_29868,N_23134,N_22995);
nand U29869 (N_29869,N_21620,N_23513);
or U29870 (N_29870,N_23321,N_19920);
or U29871 (N_29871,N_21801,N_23852);
xor U29872 (N_29872,N_21920,N_18273);
and U29873 (N_29873,N_23432,N_21157);
or U29874 (N_29874,N_19420,N_22916);
xor U29875 (N_29875,N_23832,N_22790);
nor U29876 (N_29876,N_19139,N_23755);
and U29877 (N_29877,N_18374,N_18518);
or U29878 (N_29878,N_19620,N_20658);
xor U29879 (N_29879,N_23569,N_21111);
nor U29880 (N_29880,N_22426,N_22024);
nand U29881 (N_29881,N_19962,N_21204);
and U29882 (N_29882,N_20560,N_20421);
xor U29883 (N_29883,N_19735,N_18362);
or U29884 (N_29884,N_18044,N_22652);
and U29885 (N_29885,N_22018,N_21281);
nor U29886 (N_29886,N_22016,N_19625);
or U29887 (N_29887,N_18319,N_18673);
or U29888 (N_29888,N_22056,N_19091);
nand U29889 (N_29889,N_20831,N_19465);
xnor U29890 (N_29890,N_23211,N_19160);
and U29891 (N_29891,N_22858,N_18956);
xor U29892 (N_29892,N_20856,N_22584);
xnor U29893 (N_29893,N_20254,N_23743);
nand U29894 (N_29894,N_23777,N_19335);
or U29895 (N_29895,N_21465,N_21689);
nor U29896 (N_29896,N_19329,N_21786);
nor U29897 (N_29897,N_20673,N_21076);
nor U29898 (N_29898,N_21178,N_22413);
and U29899 (N_29899,N_21870,N_19404);
nor U29900 (N_29900,N_22774,N_22551);
nor U29901 (N_29901,N_18382,N_21618);
nor U29902 (N_29902,N_21973,N_18020);
nand U29903 (N_29903,N_23050,N_22956);
and U29904 (N_29904,N_23119,N_19493);
nor U29905 (N_29905,N_18393,N_19838);
and U29906 (N_29906,N_22735,N_20208);
or U29907 (N_29907,N_18938,N_22804);
nor U29908 (N_29908,N_20286,N_18519);
nand U29909 (N_29909,N_18463,N_20263);
nor U29910 (N_29910,N_18369,N_20112);
and U29911 (N_29911,N_23914,N_21437);
or U29912 (N_29912,N_22034,N_18088);
nor U29913 (N_29913,N_18079,N_21018);
nor U29914 (N_29914,N_21608,N_18699);
nor U29915 (N_29915,N_18930,N_21819);
and U29916 (N_29916,N_19830,N_20687);
xnor U29917 (N_29917,N_22513,N_18736);
xor U29918 (N_29918,N_21439,N_23936);
nor U29919 (N_29919,N_22645,N_18241);
xnor U29920 (N_29920,N_21686,N_19443);
and U29921 (N_29921,N_18456,N_18254);
or U29922 (N_29922,N_23955,N_22417);
nor U29923 (N_29923,N_21988,N_18273);
xor U29924 (N_29924,N_20756,N_21029);
or U29925 (N_29925,N_21092,N_19689);
xnor U29926 (N_29926,N_19226,N_20645);
or U29927 (N_29927,N_19736,N_19316);
xnor U29928 (N_29928,N_22240,N_23081);
and U29929 (N_29929,N_21403,N_18488);
nor U29930 (N_29930,N_19513,N_18802);
xnor U29931 (N_29931,N_20137,N_23552);
and U29932 (N_29932,N_19594,N_21552);
nand U29933 (N_29933,N_23701,N_18456);
nor U29934 (N_29934,N_18510,N_18640);
or U29935 (N_29935,N_19120,N_21205);
xor U29936 (N_29936,N_22450,N_21579);
or U29937 (N_29937,N_20328,N_22341);
nand U29938 (N_29938,N_19104,N_18428);
and U29939 (N_29939,N_21960,N_19490);
or U29940 (N_29940,N_23238,N_20049);
xnor U29941 (N_29941,N_23639,N_22144);
and U29942 (N_29942,N_18437,N_23319);
nor U29943 (N_29943,N_22144,N_21402);
or U29944 (N_29944,N_19203,N_18242);
nor U29945 (N_29945,N_20403,N_22317);
and U29946 (N_29946,N_19986,N_21305);
nor U29947 (N_29947,N_19881,N_19150);
or U29948 (N_29948,N_19787,N_23003);
nor U29949 (N_29949,N_21804,N_22399);
and U29950 (N_29950,N_23424,N_23723);
and U29951 (N_29951,N_21627,N_18226);
and U29952 (N_29952,N_22890,N_19679);
or U29953 (N_29953,N_21671,N_23466);
or U29954 (N_29954,N_18036,N_18977);
xor U29955 (N_29955,N_19206,N_21661);
nor U29956 (N_29956,N_20576,N_20360);
and U29957 (N_29957,N_23650,N_22412);
nand U29958 (N_29958,N_21113,N_22103);
xnor U29959 (N_29959,N_19816,N_21810);
and U29960 (N_29960,N_21760,N_18059);
and U29961 (N_29961,N_20342,N_19471);
and U29962 (N_29962,N_19541,N_20499);
xnor U29963 (N_29963,N_19534,N_19503);
and U29964 (N_29964,N_23762,N_19500);
nor U29965 (N_29965,N_20263,N_18217);
and U29966 (N_29966,N_23483,N_21596);
nand U29967 (N_29967,N_22283,N_18879);
and U29968 (N_29968,N_18121,N_23040);
nand U29969 (N_29969,N_20525,N_23355);
nor U29970 (N_29970,N_18678,N_19998);
and U29971 (N_29971,N_21854,N_23888);
nand U29972 (N_29972,N_19316,N_20004);
xnor U29973 (N_29973,N_21690,N_20738);
and U29974 (N_29974,N_22209,N_23974);
and U29975 (N_29975,N_22251,N_22127);
or U29976 (N_29976,N_18392,N_21011);
nor U29977 (N_29977,N_19840,N_23279);
nand U29978 (N_29978,N_20397,N_21759);
and U29979 (N_29979,N_19751,N_18545);
or U29980 (N_29980,N_23587,N_18466);
nand U29981 (N_29981,N_19262,N_23537);
nand U29982 (N_29982,N_21648,N_20971);
nor U29983 (N_29983,N_18876,N_20794);
nand U29984 (N_29984,N_18442,N_23859);
nor U29985 (N_29985,N_18716,N_22606);
and U29986 (N_29986,N_22758,N_21894);
xor U29987 (N_29987,N_20812,N_22215);
or U29988 (N_29988,N_18195,N_21825);
and U29989 (N_29989,N_21029,N_23924);
or U29990 (N_29990,N_22118,N_20651);
nand U29991 (N_29991,N_21148,N_21658);
or U29992 (N_29992,N_18095,N_22442);
nand U29993 (N_29993,N_21208,N_20265);
and U29994 (N_29994,N_23104,N_22406);
and U29995 (N_29995,N_18519,N_21687);
nor U29996 (N_29996,N_19258,N_22964);
xnor U29997 (N_29997,N_23956,N_19604);
nand U29998 (N_29998,N_19960,N_20966);
xnor U29999 (N_29999,N_20161,N_18690);
xnor UO_0 (O_0,N_29343,N_25997);
or UO_1 (O_1,N_25990,N_29661);
and UO_2 (O_2,N_25415,N_25405);
nor UO_3 (O_3,N_29034,N_27381);
or UO_4 (O_4,N_26064,N_24273);
xnor UO_5 (O_5,N_29308,N_29589);
and UO_6 (O_6,N_29928,N_27139);
nor UO_7 (O_7,N_28374,N_28091);
nand UO_8 (O_8,N_24331,N_26929);
nor UO_9 (O_9,N_24295,N_27127);
nor UO_10 (O_10,N_27816,N_24172);
nor UO_11 (O_11,N_24050,N_25046);
nor UO_12 (O_12,N_29756,N_27164);
nand UO_13 (O_13,N_26624,N_29057);
nand UO_14 (O_14,N_26922,N_29749);
nor UO_15 (O_15,N_24061,N_26164);
nor UO_16 (O_16,N_29606,N_27762);
or UO_17 (O_17,N_26298,N_24938);
or UO_18 (O_18,N_25139,N_25572);
and UO_19 (O_19,N_24461,N_28717);
or UO_20 (O_20,N_26748,N_29154);
nor UO_21 (O_21,N_27203,N_28659);
nor UO_22 (O_22,N_25772,N_26021);
xor UO_23 (O_23,N_28350,N_24256);
xor UO_24 (O_24,N_24152,N_25000);
xor UO_25 (O_25,N_27346,N_25477);
and UO_26 (O_26,N_28042,N_25544);
or UO_27 (O_27,N_27558,N_24864);
nor UO_28 (O_28,N_27174,N_29335);
and UO_29 (O_29,N_26848,N_29344);
nor UO_30 (O_30,N_26172,N_27040);
nand UO_31 (O_31,N_25939,N_29189);
xnor UO_32 (O_32,N_24131,N_27342);
nor UO_33 (O_33,N_26450,N_27949);
nor UO_34 (O_34,N_24786,N_28459);
nand UO_35 (O_35,N_24490,N_28199);
xnor UO_36 (O_36,N_27058,N_28803);
and UO_37 (O_37,N_26525,N_25362);
nor UO_38 (O_38,N_27639,N_26803);
or UO_39 (O_39,N_24194,N_27124);
and UO_40 (O_40,N_28325,N_27288);
xnor UO_41 (O_41,N_29161,N_29988);
or UO_42 (O_42,N_29056,N_25336);
nand UO_43 (O_43,N_24663,N_27348);
and UO_44 (O_44,N_24740,N_28444);
nor UO_45 (O_45,N_26263,N_27480);
nand UO_46 (O_46,N_24922,N_25966);
nor UO_47 (O_47,N_26116,N_24683);
nand UO_48 (O_48,N_29851,N_27322);
and UO_49 (O_49,N_27080,N_28848);
nand UO_50 (O_50,N_28814,N_29775);
and UO_51 (O_51,N_27141,N_28297);
and UO_52 (O_52,N_29257,N_25947);
xnor UO_53 (O_53,N_28642,N_28117);
and UO_54 (O_54,N_24121,N_29115);
and UO_55 (O_55,N_24517,N_27024);
or UO_56 (O_56,N_26109,N_26860);
or UO_57 (O_57,N_27207,N_26451);
nand UO_58 (O_58,N_28635,N_24913);
nand UO_59 (O_59,N_29726,N_24896);
nor UO_60 (O_60,N_25443,N_25660);
nand UO_61 (O_61,N_25271,N_29625);
nor UO_62 (O_62,N_24316,N_24629);
and UO_63 (O_63,N_25112,N_29081);
nand UO_64 (O_64,N_27531,N_24435);
nor UO_65 (O_65,N_28303,N_27289);
nand UO_66 (O_66,N_24905,N_28389);
and UO_67 (O_67,N_25324,N_24552);
and UO_68 (O_68,N_24682,N_25060);
xnor UO_69 (O_69,N_24619,N_25227);
nand UO_70 (O_70,N_26968,N_28694);
nand UO_71 (O_71,N_25177,N_25432);
and UO_72 (O_72,N_25172,N_29963);
nand UO_73 (O_73,N_29750,N_29285);
nand UO_74 (O_74,N_27858,N_25108);
or UO_75 (O_75,N_27105,N_26679);
nor UO_76 (O_76,N_28442,N_27025);
xnor UO_77 (O_77,N_28646,N_25246);
xnor UO_78 (O_78,N_24892,N_28971);
or UO_79 (O_79,N_28720,N_28311);
or UO_80 (O_80,N_27197,N_25728);
or UO_81 (O_81,N_24322,N_24506);
xor UO_82 (O_82,N_24776,N_25492);
xor UO_83 (O_83,N_25674,N_24471);
nor UO_84 (O_84,N_29401,N_25501);
nand UO_85 (O_85,N_27967,N_24719);
or UO_86 (O_86,N_24804,N_28552);
or UO_87 (O_87,N_24747,N_29117);
nor UO_88 (O_88,N_24981,N_29437);
nand UO_89 (O_89,N_25483,N_28281);
nor UO_90 (O_90,N_27552,N_27400);
xor UO_91 (O_91,N_25089,N_29703);
xor UO_92 (O_92,N_29181,N_24606);
or UO_93 (O_93,N_26360,N_29708);
nand UO_94 (O_94,N_28929,N_26325);
or UO_95 (O_95,N_28804,N_25926);
nand UO_96 (O_96,N_29230,N_27768);
and UO_97 (O_97,N_27975,N_27672);
nor UO_98 (O_98,N_29441,N_26401);
xor UO_99 (O_99,N_27880,N_28284);
xor UO_100 (O_100,N_25645,N_25955);
and UO_101 (O_101,N_27498,N_27045);
and UO_102 (O_102,N_28559,N_24123);
nand UO_103 (O_103,N_25449,N_25963);
and UO_104 (O_104,N_24563,N_25727);
or UO_105 (O_105,N_29325,N_27849);
nand UO_106 (O_106,N_27625,N_24242);
nand UO_107 (O_107,N_26448,N_27367);
nand UO_108 (O_108,N_28165,N_29168);
nand UO_109 (O_109,N_28242,N_27947);
and UO_110 (O_110,N_27415,N_28737);
and UO_111 (O_111,N_28033,N_24154);
or UO_112 (O_112,N_25949,N_25145);
xor UO_113 (O_113,N_24234,N_26566);
nor UO_114 (O_114,N_29779,N_24560);
nor UO_115 (O_115,N_25014,N_24781);
nand UO_116 (O_116,N_29911,N_26965);
nor UO_117 (O_117,N_26125,N_26546);
nor UO_118 (O_118,N_26913,N_27553);
or UO_119 (O_119,N_25066,N_25684);
and UO_120 (O_120,N_24026,N_29753);
and UO_121 (O_121,N_28329,N_27933);
xor UO_122 (O_122,N_29826,N_24440);
nand UO_123 (O_123,N_24543,N_27336);
nor UO_124 (O_124,N_27930,N_24879);
nand UO_125 (O_125,N_25261,N_26117);
or UO_126 (O_126,N_24674,N_28081);
and UO_127 (O_127,N_24483,N_27153);
or UO_128 (O_128,N_27393,N_26949);
and UO_129 (O_129,N_24333,N_26771);
xnor UO_130 (O_130,N_27526,N_28621);
xnor UO_131 (O_131,N_26186,N_29083);
and UO_132 (O_132,N_25021,N_24173);
nor UO_133 (O_133,N_29504,N_27529);
nand UO_134 (O_134,N_26911,N_26408);
nor UO_135 (O_135,N_24760,N_28691);
nand UO_136 (O_136,N_28792,N_24263);
or UO_137 (O_137,N_26647,N_25111);
xnor UO_138 (O_138,N_27783,N_29188);
or UO_139 (O_139,N_28488,N_24924);
xor UO_140 (O_140,N_27865,N_28775);
nor UO_141 (O_141,N_24571,N_24268);
nand UO_142 (O_142,N_29946,N_24699);
nand UO_143 (O_143,N_25871,N_24193);
and UO_144 (O_144,N_28100,N_29784);
nand UO_145 (O_145,N_29719,N_26698);
or UO_146 (O_146,N_24287,N_25157);
and UO_147 (O_147,N_28530,N_25159);
and UO_148 (O_148,N_27927,N_28658);
nor UO_149 (O_149,N_26188,N_29608);
xnor UO_150 (O_150,N_28221,N_28783);
xnor UO_151 (O_151,N_27056,N_28336);
nand UO_152 (O_152,N_29355,N_25864);
or UO_153 (O_153,N_29588,N_26684);
nor UO_154 (O_154,N_28246,N_27456);
and UO_155 (O_155,N_25913,N_28678);
or UO_156 (O_156,N_29214,N_28158);
nand UO_157 (O_157,N_29242,N_26670);
and UO_158 (O_158,N_24254,N_28432);
nand UO_159 (O_159,N_27165,N_27380);
or UO_160 (O_160,N_29402,N_28386);
nand UO_161 (O_161,N_26407,N_25798);
or UO_162 (O_162,N_27107,N_25444);
nor UO_163 (O_163,N_26359,N_29924);
nor UO_164 (O_164,N_26043,N_24056);
and UO_165 (O_165,N_26403,N_28813);
xnor UO_166 (O_166,N_25075,N_25081);
nor UO_167 (O_167,N_24579,N_27991);
and UO_168 (O_168,N_27414,N_29627);
and UO_169 (O_169,N_24431,N_28131);
xor UO_170 (O_170,N_26919,N_26356);
nor UO_171 (O_171,N_27626,N_27210);
nand UO_172 (O_172,N_26273,N_25440);
and UO_173 (O_173,N_27151,N_25267);
xor UO_174 (O_174,N_28353,N_29116);
nor UO_175 (O_175,N_27546,N_27999);
or UO_176 (O_176,N_29194,N_24145);
nor UO_177 (O_177,N_29793,N_27824);
or UO_178 (O_178,N_24837,N_29629);
or UO_179 (O_179,N_28791,N_27795);
and UO_180 (O_180,N_28431,N_27700);
and UO_181 (O_181,N_28087,N_26813);
xor UO_182 (O_182,N_24842,N_24303);
and UO_183 (O_183,N_28112,N_28435);
and UO_184 (O_184,N_28639,N_26974);
and UO_185 (O_185,N_29112,N_26784);
xnor UO_186 (O_186,N_27302,N_28761);
or UO_187 (O_187,N_29463,N_25920);
nor UO_188 (O_188,N_29326,N_28312);
nor UO_189 (O_189,N_27473,N_24603);
or UO_190 (O_190,N_27185,N_25635);
xnor UO_191 (O_191,N_26462,N_27066);
xnor UO_192 (O_192,N_27859,N_25846);
nor UO_193 (O_193,N_25346,N_28757);
xnor UO_194 (O_194,N_29878,N_27216);
or UO_195 (O_195,N_29091,N_29718);
and UO_196 (O_196,N_29987,N_28317);
nand UO_197 (O_197,N_26822,N_24686);
xnor UO_198 (O_198,N_24601,N_27032);
nand UO_199 (O_199,N_24023,N_26823);
and UO_200 (O_200,N_29646,N_27397);
nor UO_201 (O_201,N_28664,N_26687);
xor UO_202 (O_202,N_24714,N_29050);
nand UO_203 (O_203,N_26983,N_29426);
xor UO_204 (O_204,N_26899,N_28385);
nor UO_205 (O_205,N_24111,N_29932);
or UO_206 (O_206,N_27007,N_29918);
nor UO_207 (O_207,N_24280,N_26237);
xnor UO_208 (O_208,N_25950,N_28995);
or UO_209 (O_209,N_24100,N_27838);
nor UO_210 (O_210,N_24209,N_29813);
nand UO_211 (O_211,N_27026,N_25115);
nor UO_212 (O_212,N_29481,N_27786);
xor UO_213 (O_213,N_24124,N_24417);
or UO_214 (O_214,N_25166,N_24546);
nor UO_215 (O_215,N_26418,N_24385);
nor UO_216 (O_216,N_26554,N_28676);
xor UO_217 (O_217,N_24350,N_24646);
nand UO_218 (O_218,N_29432,N_29533);
or UO_219 (O_219,N_24752,N_29954);
nor UO_220 (O_220,N_25377,N_24328);
and UO_221 (O_221,N_27855,N_27134);
or UO_222 (O_222,N_26124,N_27049);
nand UO_223 (O_223,N_25775,N_27466);
nor UO_224 (O_224,N_24665,N_25489);
nor UO_225 (O_225,N_27372,N_25892);
xor UO_226 (O_226,N_25753,N_25826);
or UO_227 (O_227,N_28301,N_28521);
and UO_228 (O_228,N_24176,N_29591);
and UO_229 (O_229,N_26209,N_29002);
or UO_230 (O_230,N_27976,N_24232);
and UO_231 (O_231,N_24470,N_25817);
nor UO_232 (O_232,N_27198,N_28476);
nor UO_233 (O_233,N_25317,N_27262);
or UO_234 (O_234,N_27805,N_29716);
or UO_235 (O_235,N_27726,N_26674);
and UO_236 (O_236,N_24219,N_29974);
or UO_237 (O_237,N_27407,N_27461);
nor UO_238 (O_238,N_26299,N_26948);
and UO_239 (O_239,N_26023,N_29534);
nor UO_240 (O_240,N_29539,N_24927);
xnor UO_241 (O_241,N_25142,N_24153);
nor UO_242 (O_242,N_25124,N_24183);
nor UO_243 (O_243,N_24736,N_24778);
nand UO_244 (O_244,N_28942,N_28710);
or UO_245 (O_245,N_28322,N_27962);
nor UO_246 (O_246,N_28926,N_28376);
or UO_247 (O_247,N_26222,N_28426);
nand UO_248 (O_248,N_24359,N_27484);
nand UO_249 (O_249,N_26597,N_28893);
and UO_250 (O_250,N_26709,N_27359);
nand UO_251 (O_251,N_29675,N_27054);
xor UO_252 (O_252,N_26874,N_27736);
and UO_253 (O_253,N_29183,N_25685);
nand UO_254 (O_254,N_26495,N_28508);
xor UO_255 (O_255,N_26569,N_27735);
or UO_256 (O_256,N_27450,N_25325);
and UO_257 (O_257,N_24910,N_29372);
nor UO_258 (O_258,N_29455,N_24832);
nand UO_259 (O_259,N_29762,N_25872);
xnor UO_260 (O_260,N_28863,N_28203);
or UO_261 (O_261,N_26639,N_25549);
nor UO_262 (O_262,N_29386,N_27964);
nor UO_263 (O_263,N_24511,N_26484);
xnor UO_264 (O_264,N_27811,N_26643);
and UO_265 (O_265,N_29579,N_27455);
xor UO_266 (O_266,N_26686,N_29648);
or UO_267 (O_267,N_28269,N_24956);
and UO_268 (O_268,N_26627,N_26447);
and UO_269 (O_269,N_25977,N_27368);
and UO_270 (O_270,N_28927,N_24749);
nand UO_271 (O_271,N_24725,N_24524);
nor UO_272 (O_272,N_27852,N_29819);
or UO_273 (O_273,N_26248,N_27196);
or UO_274 (O_274,N_29713,N_28633);
xnor UO_275 (O_275,N_26699,N_25245);
nand UO_276 (O_276,N_24166,N_27744);
xor UO_277 (O_277,N_28064,N_28118);
and UO_278 (O_278,N_29542,N_27649);
and UO_279 (O_279,N_24772,N_26726);
xor UO_280 (O_280,N_26957,N_28941);
or UO_281 (O_281,N_27901,N_24383);
nor UO_282 (O_282,N_26873,N_26570);
xor UO_283 (O_283,N_27512,N_24092);
and UO_284 (O_284,N_26166,N_24836);
nand UO_285 (O_285,N_27409,N_24319);
and UO_286 (O_286,N_25792,N_29806);
nor UO_287 (O_287,N_25153,N_27004);
and UO_288 (O_288,N_25958,N_25236);
xor UO_289 (O_289,N_28984,N_29883);
xor UO_290 (O_290,N_29487,N_28826);
or UO_291 (O_291,N_27750,N_27360);
nor UO_292 (O_292,N_24365,N_28596);
nand UO_293 (O_293,N_29131,N_24707);
and UO_294 (O_294,N_24667,N_24679);
nand UO_295 (O_295,N_24867,N_24831);
nand UO_296 (O_296,N_27278,N_25965);
or UO_297 (O_297,N_26144,N_26892);
xnor UO_298 (O_298,N_29106,N_24897);
or UO_299 (O_299,N_27717,N_28765);
or UO_300 (O_300,N_27001,N_29674);
or UO_301 (O_301,N_25269,N_25927);
and UO_302 (O_302,N_24535,N_26039);
nor UO_303 (O_303,N_24126,N_27503);
nor UO_304 (O_304,N_25059,N_27585);
nor UO_305 (O_305,N_28089,N_26029);
xnor UO_306 (O_306,N_27022,N_25366);
xor UO_307 (O_307,N_29262,N_24069);
or UO_308 (O_308,N_27477,N_28668);
nor UO_309 (O_309,N_25044,N_28975);
and UO_310 (O_310,N_28843,N_24114);
nand UO_311 (O_311,N_24642,N_27312);
xor UO_312 (O_312,N_24053,N_27023);
nor UO_313 (O_313,N_28293,N_25090);
nor UO_314 (O_314,N_26497,N_25680);
nand UO_315 (O_315,N_24190,N_24341);
or UO_316 (O_316,N_29382,N_27813);
nor UO_317 (O_317,N_28039,N_28485);
or UO_318 (O_318,N_29073,N_28913);
nand UO_319 (O_319,N_28475,N_29584);
nand UO_320 (O_320,N_24159,N_25825);
nand UO_321 (O_321,N_28471,N_25322);
and UO_322 (O_322,N_29869,N_25526);
or UO_323 (O_323,N_29628,N_24810);
or UO_324 (O_324,N_26307,N_25559);
or UO_325 (O_325,N_25176,N_28196);
xor UO_326 (O_326,N_26837,N_24139);
or UO_327 (O_327,N_25371,N_28250);
nor UO_328 (O_328,N_27604,N_26781);
and UO_329 (O_329,N_24748,N_26632);
nor UO_330 (O_330,N_27634,N_27041);
nand UO_331 (O_331,N_24021,N_26113);
or UO_332 (O_332,N_27948,N_26316);
or UO_333 (O_333,N_27707,N_27223);
xor UO_334 (O_334,N_27969,N_25815);
nor UO_335 (O_335,N_25074,N_29316);
nor UO_336 (O_336,N_28541,N_28959);
xor UO_337 (O_337,N_27444,N_29936);
nand UO_338 (O_338,N_26474,N_26322);
and UO_339 (O_339,N_26390,N_27090);
and UO_340 (O_340,N_29933,N_28839);
or UO_341 (O_341,N_25612,N_24978);
nor UO_342 (O_342,N_24272,N_24589);
nand UO_343 (O_343,N_24570,N_29324);
xor UO_344 (O_344,N_29972,N_25458);
and UO_345 (O_345,N_28265,N_27423);
and UO_346 (O_346,N_26045,N_29417);
xnor UO_347 (O_347,N_24645,N_27067);
or UO_348 (O_348,N_24208,N_27660);
and UO_349 (O_349,N_28790,N_25585);
or UO_350 (O_350,N_24951,N_28636);
and UO_351 (O_351,N_26989,N_29536);
xnor UO_352 (O_352,N_26309,N_28032);
xor UO_353 (O_353,N_28360,N_27109);
nor UO_354 (O_354,N_27984,N_25714);
nand UO_355 (O_355,N_28438,N_29097);
nand UO_356 (O_356,N_24243,N_25859);
and UO_357 (O_357,N_29418,N_27803);
nor UO_358 (O_358,N_25352,N_27365);
nor UO_359 (O_359,N_26522,N_24871);
or UO_360 (O_360,N_24632,N_28028);
or UO_361 (O_361,N_26003,N_27428);
nand UO_362 (O_362,N_24575,N_24376);
xnor UO_363 (O_363,N_27490,N_28592);
nand UO_364 (O_364,N_25387,N_27084);
xor UO_365 (O_365,N_27872,N_27468);
and UO_366 (O_366,N_28056,N_29714);
or UO_367 (O_367,N_28878,N_25796);
xnor UO_368 (O_368,N_28419,N_27081);
xor UO_369 (O_369,N_24636,N_26438);
nor UO_370 (O_370,N_25654,N_29634);
and UO_371 (O_371,N_25156,N_25408);
or UO_372 (O_372,N_29951,N_27422);
and UO_373 (O_373,N_24529,N_24149);
nor UO_374 (O_374,N_24132,N_28615);
xnor UO_375 (O_375,N_25876,N_24787);
nand UO_376 (O_376,N_26455,N_26320);
xor UO_377 (O_377,N_25785,N_29103);
nor UO_378 (O_378,N_29420,N_27663);
or UO_379 (O_379,N_29647,N_24761);
nand UO_380 (O_380,N_26996,N_28579);
nand UO_381 (O_381,N_26910,N_25276);
nor UO_382 (O_382,N_27167,N_29226);
nor UO_383 (O_383,N_24485,N_29952);
nand UO_384 (O_384,N_29198,N_29768);
and UO_385 (O_385,N_28557,N_29577);
and UO_386 (O_386,N_24403,N_28218);
nand UO_387 (O_387,N_26787,N_29614);
and UO_388 (O_388,N_27188,N_24205);
xor UO_389 (O_389,N_27183,N_26135);
and UO_390 (O_390,N_24229,N_26206);
xor UO_391 (O_391,N_28163,N_28292);
xor UO_392 (O_392,N_29502,N_26564);
or UO_393 (O_393,N_29009,N_28168);
and UO_394 (O_394,N_28420,N_29252);
nand UO_395 (O_395,N_28811,N_28865);
nor UO_396 (O_396,N_26828,N_25803);
or UO_397 (O_397,N_26622,N_28680);
nor UO_398 (O_398,N_27199,N_29472);
nand UO_399 (O_399,N_27374,N_27541);
or UO_400 (O_400,N_25481,N_25895);
or UO_401 (O_401,N_28111,N_25962);
nand UO_402 (O_402,N_29535,N_26347);
nor UO_403 (O_403,N_25369,N_26312);
or UO_404 (O_404,N_26470,N_26844);
nand UO_405 (O_405,N_25183,N_26654);
nor UO_406 (O_406,N_27285,N_26226);
nor UO_407 (O_407,N_25472,N_27297);
nand UO_408 (O_408,N_28750,N_29669);
nor UO_409 (O_409,N_24408,N_28068);
and UO_410 (O_410,N_25766,N_27763);
nor UO_411 (O_411,N_29339,N_24542);
xor UO_412 (O_412,N_26001,N_27913);
nor UO_413 (O_413,N_26349,N_28686);
nand UO_414 (O_414,N_25531,N_29158);
or UO_415 (O_415,N_29844,N_29421);
nand UO_416 (O_416,N_29126,N_25085);
nand UO_417 (O_417,N_24313,N_29644);
and UO_418 (O_418,N_25850,N_25017);
nand UO_419 (O_419,N_24849,N_27110);
and UO_420 (O_420,N_24826,N_28457);
and UO_421 (O_421,N_27130,N_29528);
nor UO_422 (O_422,N_25563,N_26238);
nand UO_423 (O_423,N_24024,N_25231);
and UO_424 (O_424,N_25218,N_25462);
and UO_425 (O_425,N_28285,N_24577);
xor UO_426 (O_426,N_28358,N_29052);
nor UO_427 (O_427,N_25622,N_29261);
and UO_428 (O_428,N_26946,N_27097);
and UO_429 (O_429,N_28059,N_25149);
xnor UO_430 (O_430,N_25786,N_28335);
and UO_431 (O_431,N_28237,N_24655);
nor UO_432 (O_432,N_26834,N_25535);
xnor UO_433 (O_433,N_27800,N_28260);
or UO_434 (O_434,N_25981,N_26052);
or UO_435 (O_435,N_29738,N_24693);
xnor UO_436 (O_436,N_26225,N_24215);
or UO_437 (O_437,N_29476,N_27405);
nor UO_438 (O_438,N_26344,N_29953);
nor UO_439 (O_439,N_26078,N_25437);
and UO_440 (O_440,N_24358,N_29479);
nor UO_441 (O_441,N_29686,N_28201);
xnor UO_442 (O_442,N_26330,N_26138);
or UO_443 (O_443,N_28090,N_25426);
or UO_444 (O_444,N_28525,N_26293);
xor UO_445 (O_445,N_25607,N_29916);
nand UO_446 (O_446,N_28076,N_29555);
and UO_447 (O_447,N_27996,N_28896);
nand UO_448 (O_448,N_28810,N_27510);
and UO_449 (O_449,N_29248,N_27968);
or UO_450 (O_450,N_28327,N_26097);
or UO_451 (O_451,N_24116,N_25133);
nor UO_452 (O_452,N_24433,N_28660);
or UO_453 (O_453,N_25606,N_24954);
xnor UO_454 (O_454,N_28828,N_28645);
nand UO_455 (O_455,N_28429,N_29379);
nor UO_456 (O_456,N_26881,N_29939);
or UO_457 (O_457,N_26680,N_26667);
nand UO_458 (O_458,N_25239,N_26400);
nor UO_459 (O_459,N_28663,N_28688);
or UO_460 (O_460,N_29245,N_26866);
and UO_461 (O_461,N_29396,N_26548);
or UO_462 (O_462,N_24594,N_28495);
nand UO_463 (O_463,N_26435,N_26292);
xor UO_464 (O_464,N_29216,N_24661);
nor UO_465 (O_465,N_27464,N_25941);
and UO_466 (O_466,N_27245,N_28960);
or UO_467 (O_467,N_26137,N_25084);
and UO_468 (O_468,N_29664,N_27832);
nor UO_469 (O_469,N_29438,N_28911);
nor UO_470 (O_470,N_27010,N_26749);
and UO_471 (O_471,N_26926,N_26806);
xnor UO_472 (O_472,N_26835,N_29556);
or UO_473 (O_473,N_29825,N_29696);
or UO_474 (O_474,N_28051,N_26423);
nor UO_475 (O_475,N_24507,N_27094);
and UO_476 (O_476,N_25533,N_25129);
xor UO_477 (O_477,N_29681,N_29607);
and UO_478 (O_478,N_24275,N_25180);
and UO_479 (O_479,N_27350,N_27892);
xor UO_480 (O_480,N_25736,N_27449);
xnor UO_481 (O_481,N_26783,N_24844);
xor UO_482 (O_482,N_26121,N_25809);
xnor UO_483 (O_483,N_25457,N_24068);
or UO_484 (O_484,N_29691,N_26473);
nand UO_485 (O_485,N_24734,N_24712);
nand UO_486 (O_486,N_27059,N_26846);
xnor UO_487 (O_487,N_28366,N_24448);
nor UO_488 (O_488,N_26762,N_24684);
or UO_489 (O_489,N_29159,N_26802);
xor UO_490 (O_490,N_26034,N_26310);
nor UO_491 (O_491,N_25099,N_29766);
xor UO_492 (O_492,N_26703,N_29038);
or UO_493 (O_493,N_27317,N_25182);
xor UO_494 (O_494,N_27688,N_29662);
and UO_495 (O_495,N_29613,N_27021);
nand UO_496 (O_496,N_29095,N_28964);
or UO_497 (O_497,N_25070,N_29548);
nand UO_498 (O_498,N_28490,N_27711);
nor UO_499 (O_499,N_24953,N_28700);
or UO_500 (O_500,N_28454,N_28591);
or UO_501 (O_501,N_29410,N_24708);
and UO_502 (O_502,N_26227,N_27519);
or UO_503 (O_503,N_26442,N_25800);
xor UO_504 (O_504,N_24251,N_25206);
and UO_505 (O_505,N_28978,N_26270);
xnor UO_506 (O_506,N_25422,N_28271);
nand UO_507 (O_507,N_27703,N_26601);
and UO_508 (O_508,N_26046,N_28267);
xor UO_509 (O_509,N_29239,N_24059);
xnor UO_510 (O_510,N_28945,N_25793);
nor UO_511 (O_511,N_28186,N_29640);
and UO_512 (O_512,N_24763,N_25486);
nor UO_513 (O_513,N_25822,N_25668);
or UO_514 (O_514,N_25633,N_25720);
nand UO_515 (O_515,N_25820,N_25940);
xor UO_516 (O_516,N_28604,N_25024);
or UO_517 (O_517,N_29167,N_26069);
nand UO_518 (O_518,N_24673,N_28561);
nand UO_519 (O_519,N_28902,N_24067);
xor UO_520 (O_520,N_29047,N_24266);
xnor UO_521 (O_521,N_25745,N_27857);
and UO_522 (O_522,N_29576,N_28263);
and UO_523 (O_523,N_24586,N_28598);
nor UO_524 (O_524,N_25233,N_27944);
nand UO_525 (O_525,N_25274,N_26884);
nor UO_526 (O_526,N_28189,N_28497);
or UO_527 (O_527,N_25163,N_25242);
and UO_528 (O_528,N_28095,N_28565);
xnor UO_529 (O_529,N_25171,N_27038);
nor UO_530 (O_530,N_28818,N_27100);
or UO_531 (O_531,N_25810,N_29152);
nor UO_532 (O_532,N_24312,N_29135);
or UO_533 (O_533,N_24746,N_29010);
or UO_534 (O_534,N_24741,N_25162);
xor UO_535 (O_535,N_28812,N_29059);
xnor UO_536 (O_536,N_26986,N_28370);
or UO_537 (O_537,N_29484,N_27836);
xor UO_538 (O_538,N_28328,N_27891);
xnor UO_539 (O_539,N_24422,N_28015);
xor UO_540 (O_540,N_25228,N_27404);
nor UO_541 (O_541,N_26128,N_26945);
nor UO_542 (O_542,N_24115,N_28504);
nor UO_543 (O_543,N_25524,N_26770);
nand UO_544 (O_544,N_27299,N_28088);
xnor UO_545 (O_545,N_29929,N_25514);
xnor UO_546 (O_546,N_27387,N_25378);
or UO_547 (O_547,N_27113,N_26065);
xnor UO_548 (O_548,N_29153,N_25316);
xnor UO_549 (O_549,N_29349,N_25191);
nand UO_550 (O_550,N_27345,N_28379);
and UO_551 (O_551,N_29294,N_24814);
nand UO_552 (O_552,N_27738,N_25360);
nor UO_553 (O_553,N_28616,N_27119);
or UO_554 (O_554,N_29016,N_25647);
xor UO_555 (O_555,N_28417,N_26074);
nor UO_556 (O_556,N_29751,N_24289);
and UO_557 (O_557,N_29133,N_24841);
or UO_558 (O_558,N_29390,N_25368);
nand UO_559 (O_559,N_25064,N_26004);
nand UO_560 (O_560,N_26236,N_28305);
nor UO_561 (O_561,N_25048,N_27798);
and UO_562 (O_562,N_25557,N_29573);
and UO_563 (O_563,N_27622,N_28256);
nand UO_564 (O_564,N_25088,N_29968);
xnor UO_565 (O_565,N_25903,N_24903);
and UO_566 (O_566,N_27758,N_25758);
and UO_567 (O_567,N_26811,N_27971);
nor UO_568 (O_568,N_28355,N_24827);
nand UO_569 (O_569,N_28522,N_25746);
nand UO_570 (O_570,N_29850,N_26852);
or UO_571 (O_571,N_25038,N_26799);
nor UO_572 (O_572,N_24730,N_24668);
nor UO_573 (O_573,N_26305,N_26824);
xor UO_574 (O_574,N_29715,N_29653);
xnor UO_575 (O_575,N_28083,N_28982);
and UO_576 (O_576,N_26702,N_28513);
and UO_577 (O_577,N_25788,N_28278);
nand UO_578 (O_578,N_29785,N_28409);
or UO_579 (O_579,N_26200,N_26545);
and UO_580 (O_580,N_27772,N_26296);
xor UO_581 (O_581,N_26315,N_24766);
nor UO_582 (O_582,N_28208,N_28005);
nor UO_583 (O_583,N_27687,N_29488);
xnor UO_584 (O_584,N_28215,N_26142);
and UO_585 (O_585,N_25923,N_28772);
and UO_586 (O_586,N_27528,N_27135);
nor UO_587 (O_587,N_28021,N_28424);
and UO_588 (O_588,N_24882,N_28570);
nor UO_589 (O_589,N_28733,N_27161);
nor UO_590 (O_590,N_24047,N_25126);
nand UO_591 (O_591,N_24624,N_29179);
or UO_592 (O_592,N_27851,N_28973);
and UO_593 (O_593,N_25445,N_29847);
nand UO_594 (O_594,N_24614,N_24675);
and UO_595 (O_595,N_25385,N_27386);
and UO_596 (O_596,N_28983,N_26977);
or UO_597 (O_597,N_24883,N_29346);
nand UO_598 (O_598,N_28503,N_28096);
and UO_599 (O_599,N_27416,N_26997);
nand UO_600 (O_600,N_25396,N_28306);
nand UO_601 (O_601,N_26535,N_24382);
nor UO_602 (O_602,N_27764,N_29880);
xnor UO_603 (O_603,N_29272,N_28859);
or UO_604 (O_604,N_24522,N_26460);
or UO_605 (O_605,N_26656,N_26809);
nor UO_606 (O_606,N_25468,N_29098);
xor UO_607 (O_607,N_26434,N_27193);
or UO_608 (O_608,N_25224,N_25033);
nor UO_609 (O_609,N_27447,N_24930);
xnor UO_610 (O_610,N_25620,N_24569);
and UO_611 (O_611,N_25118,N_27268);
nand UO_612 (O_612,N_29821,N_27754);
or UO_613 (O_613,N_27052,N_28837);
nor UO_614 (O_614,N_27908,N_26614);
nor UO_615 (O_615,N_24874,N_29811);
and UO_616 (O_616,N_28673,N_24010);
or UO_617 (O_617,N_29456,N_24660);
and UO_618 (O_618,N_29594,N_28721);
nand UO_619 (O_619,N_24137,N_25345);
nand UO_620 (O_620,N_29110,N_28849);
xnor UO_621 (O_621,N_24474,N_24491);
xor UO_622 (O_622,N_26741,N_29392);
and UO_623 (O_623,N_25953,N_24476);
and UO_624 (O_624,N_25320,N_26585);
nor UO_625 (O_625,N_24727,N_28310);
and UO_626 (O_626,N_29531,N_29986);
and UO_627 (O_627,N_28887,N_29466);
or UO_628 (O_628,N_27395,N_26220);
nor UO_629 (O_629,N_25330,N_26355);
nor UO_630 (O_630,N_26943,N_24110);
nor UO_631 (O_631,N_26251,N_28756);
nor UO_632 (O_632,N_29615,N_28852);
xor UO_633 (O_633,N_28544,N_26671);
xnor UO_634 (O_634,N_26284,N_25179);
or UO_635 (O_635,N_26410,N_24245);
and UO_636 (O_636,N_27215,N_28648);
nand UO_637 (O_637,N_25057,N_27596);
xor UO_638 (O_638,N_27518,N_25291);
and UO_639 (O_639,N_28725,N_25706);
and UO_640 (O_640,N_28780,N_28656);
or UO_641 (O_641,N_28494,N_27580);
and UO_642 (O_642,N_27509,N_25930);
nor UO_643 (O_643,N_25248,N_25100);
and UO_644 (O_644,N_27411,N_25030);
xnor UO_645 (O_645,N_28233,N_24227);
nor UO_646 (O_646,N_28077,N_26514);
nor UO_647 (O_647,N_25529,N_28798);
nor UO_648 (O_648,N_24654,N_29692);
and UO_649 (O_649,N_27614,N_27425);
xor UO_650 (O_650,N_29416,N_24834);
nor UO_651 (O_651,N_27378,N_29446);
nand UO_652 (O_652,N_25890,N_24715);
xnor UO_653 (O_653,N_27746,N_25539);
or UO_654 (O_654,N_26914,N_27611);
nand UO_655 (O_655,N_26020,N_25453);
xor UO_656 (O_656,N_28864,N_28895);
nor UO_657 (O_657,N_28901,N_25726);
or UO_658 (O_658,N_25418,N_25303);
xnor UO_659 (O_659,N_24169,N_26280);
or UO_660 (O_660,N_28043,N_27590);
nand UO_661 (O_661,N_25818,N_27489);
and UO_662 (O_662,N_29684,N_26103);
nand UO_663 (O_663,N_29166,N_28754);
or UO_664 (O_664,N_27740,N_28411);
nand UO_665 (O_665,N_27437,N_28789);
xnor UO_666 (O_666,N_27474,N_29760);
or UO_667 (O_667,N_26731,N_24413);
nand UO_668 (O_668,N_28086,N_26129);
and UO_669 (O_669,N_26623,N_29225);
and UO_670 (O_670,N_28589,N_24743);
and UO_671 (O_671,N_29199,N_26105);
xnor UO_672 (O_672,N_26147,N_28994);
nor UO_673 (O_673,N_29792,N_29228);
xnor UO_674 (O_674,N_28768,N_25174);
nor UO_675 (O_675,N_25912,N_26817);
and UO_676 (O_676,N_24912,N_25282);
nand UO_677 (O_677,N_24424,N_24898);
and UO_678 (O_678,N_24944,N_28177);
nor UO_679 (O_679,N_25400,N_27938);
nand UO_680 (O_680,N_26482,N_26258);
nor UO_681 (O_681,N_25484,N_24397);
or UO_682 (O_682,N_26879,N_26553);
nand UO_683 (O_683,N_27894,N_25877);
or UO_684 (O_684,N_25860,N_27575);
xor UO_685 (O_685,N_29741,N_24616);
and UO_686 (O_686,N_24943,N_28125);
xnor UO_687 (O_687,N_28324,N_27793);
or UO_688 (O_688,N_26810,N_25446);
or UO_689 (O_689,N_26468,N_24789);
or UO_690 (O_690,N_25701,N_25834);
or UO_691 (O_691,N_27051,N_28928);
xor UO_692 (O_692,N_27269,N_24627);
nor UO_693 (O_693,N_29210,N_25067);
nor UO_694 (O_694,N_26286,N_26501);
and UO_695 (O_695,N_29011,N_28249);
xor UO_696 (O_696,N_26976,N_29497);
nor UO_697 (O_697,N_26414,N_25510);
nor UO_698 (O_698,N_28408,N_29585);
xor UO_699 (O_699,N_27767,N_29840);
nor UO_700 (O_700,N_28715,N_29494);
nor UO_701 (O_701,N_24862,N_25284);
or UO_702 (O_702,N_27612,N_29287);
xor UO_703 (O_703,N_27307,N_26114);
nor UO_704 (O_704,N_28564,N_25596);
nand UO_705 (O_705,N_27465,N_28013);
and UO_706 (O_706,N_26711,N_25733);
and UO_707 (O_707,N_28551,N_29884);
xor UO_708 (O_708,N_24239,N_27055);
xor UO_709 (O_709,N_25634,N_28602);
nand UO_710 (O_710,N_28628,N_26077);
or UO_711 (O_711,N_24744,N_28456);
nor UO_712 (O_712,N_25214,N_27621);
xnor UO_713 (O_713,N_27778,N_28643);
nand UO_714 (O_714,N_29480,N_29413);
nand UO_715 (O_715,N_24677,N_27255);
and UO_716 (O_716,N_24925,N_24425);
and UO_717 (O_717,N_25315,N_24909);
xnor UO_718 (O_718,N_28996,N_28622);
nand UO_719 (O_719,N_28239,N_27027);
nor UO_720 (O_720,N_25076,N_25215);
xnor UO_721 (O_721,N_28012,N_28704);
nor UO_722 (O_722,N_26644,N_26014);
xnor UO_723 (O_723,N_25374,N_28923);
or UO_724 (O_724,N_25729,N_29398);
or UO_725 (O_725,N_26141,N_27815);
or UO_726 (O_726,N_26615,N_27655);
xor UO_727 (O_727,N_27881,N_29604);
xor UO_728 (O_728,N_29582,N_25160);
nand UO_729 (O_729,N_26661,N_25528);
xnor UO_730 (O_730,N_24723,N_24449);
or UO_731 (O_731,N_28610,N_24108);
nor UO_732 (O_732,N_24462,N_29254);
and UO_733 (O_733,N_29781,N_28613);
xnor UO_734 (O_734,N_24052,N_25709);
xnor UO_735 (O_735,N_24515,N_26233);
xnor UO_736 (O_736,N_24755,N_26005);
and UO_737 (O_737,N_27823,N_26889);
nand UO_738 (O_738,N_25299,N_28903);
nand UO_739 (O_739,N_25970,N_24302);
xor UO_740 (O_740,N_24751,N_26695);
and UO_741 (O_741,N_26738,N_24246);
xor UO_742 (O_742,N_28245,N_24688);
nor UO_743 (O_743,N_26556,N_29314);
xnor UO_744 (O_744,N_24373,N_26982);
and UO_745 (O_745,N_25558,N_28275);
and UO_746 (O_746,N_25795,N_29962);
nor UO_747 (O_747,N_24003,N_27327);
nand UO_748 (O_748,N_28823,N_27844);
nor UO_749 (O_749,N_29204,N_26967);
or UO_750 (O_750,N_24720,N_29834);
nand UO_751 (O_751,N_24527,N_25661);
nor UO_752 (O_752,N_27033,N_26197);
or UO_753 (O_753,N_24285,N_25716);
and UO_754 (O_754,N_27682,N_29599);
nor UO_755 (O_755,N_25188,N_28638);
and UO_756 (O_756,N_25192,N_25007);
xor UO_757 (O_757,N_26354,N_29310);
nor UO_758 (O_758,N_29682,N_29976);
and UO_759 (O_759,N_26933,N_24444);
nor UO_760 (O_760,N_28985,N_24923);
nor UO_761 (O_761,N_28634,N_26406);
nor UO_762 (O_762,N_24429,N_24652);
nand UO_763 (O_763,N_27961,N_27633);
and UO_764 (O_764,N_29055,N_27029);
or UO_765 (O_765,N_25146,N_25605);
xor UO_766 (O_766,N_29340,N_27115);
xor UO_767 (O_767,N_27847,N_28805);
or UO_768 (O_768,N_28749,N_27577);
nor UO_769 (O_769,N_25835,N_26637);
and UO_770 (O_770,N_27701,N_27862);
xor UO_771 (O_771,N_28573,N_26715);
nor UO_772 (O_772,N_25498,N_29283);
nand UO_773 (O_773,N_26063,N_26366);
xnor UO_774 (O_774,N_25523,N_24931);
nand UO_775 (O_775,N_24034,N_26002);
xor UO_776 (O_776,N_27311,N_24066);
nor UO_777 (O_777,N_27666,N_26373);
xnor UO_778 (O_778,N_25403,N_24420);
nor UO_779 (O_779,N_25015,N_26737);
or UO_780 (O_780,N_28375,N_26500);
xor UO_781 (O_781,N_29601,N_25771);
nand UO_782 (O_782,N_27417,N_28906);
nor UO_783 (O_783,N_24811,N_25723);
or UO_784 (O_784,N_29270,N_29523);
nand UO_785 (O_785,N_24676,N_24113);
nand UO_786 (O_786,N_24984,N_28252);
nand UO_787 (O_787,N_26477,N_27722);
and UO_788 (O_788,N_28236,N_26174);
xor UO_789 (O_789,N_27559,N_27571);
and UO_790 (O_790,N_26246,N_24179);
xor UO_791 (O_791,N_24573,N_29383);
nor UO_792 (O_792,N_27544,N_29912);
nand UO_793 (O_793,N_27452,N_27313);
nor UO_794 (O_794,N_28987,N_26786);
nand UO_795 (O_795,N_24493,N_26862);
nand UO_796 (O_796,N_25849,N_26740);
xnor UO_797 (O_797,N_25065,N_25513);
or UO_798 (O_798,N_28211,N_28827);
or UO_799 (O_799,N_24843,N_28461);
and UO_800 (O_800,N_28412,N_29746);
or UO_801 (O_801,N_29336,N_24077);
and UO_802 (O_802,N_25814,N_29218);
and UO_803 (O_803,N_24937,N_29776);
and UO_804 (O_804,N_25574,N_27479);
xnor UO_805 (O_805,N_28917,N_27820);
and UO_806 (O_806,N_29171,N_29688);
nor UO_807 (O_807,N_26465,N_27266);
and UO_808 (O_808,N_28883,N_24148);
or UO_809 (O_809,N_25508,N_25399);
and UO_810 (O_810,N_27946,N_24850);
xor UO_811 (O_811,N_26212,N_25730);
and UO_812 (O_812,N_26191,N_25616);
nor UO_813 (O_813,N_27492,N_27117);
nand UO_814 (O_814,N_25705,N_29967);
nand UO_815 (O_815,N_24342,N_27533);
and UO_816 (O_816,N_25543,N_28891);
nor UO_817 (O_817,N_29318,N_29575);
and UO_818 (O_818,N_28529,N_28788);
nand UO_819 (O_819,N_29593,N_28300);
and UO_820 (O_820,N_27344,N_24398);
or UO_821 (O_821,N_29101,N_25783);
nor UO_822 (O_822,N_28993,N_27974);
and UO_823 (O_823,N_27310,N_26058);
nor UO_824 (O_824,N_24320,N_27941);
or UO_825 (O_825,N_29724,N_25569);
xnor UO_826 (O_826,N_24489,N_28763);
nand UO_827 (O_827,N_25054,N_29665);
nand UO_828 (O_828,N_29385,N_28404);
nor UO_829 (O_829,N_24830,N_29232);
and UO_830 (O_830,N_27662,N_27235);
nand UO_831 (O_831,N_24099,N_29023);
xnor UO_832 (O_832,N_29454,N_28861);
nand UO_833 (O_833,N_28354,N_27839);
nor UO_834 (O_834,N_27669,N_24394);
nand UO_835 (O_835,N_25551,N_25628);
nand UO_836 (O_836,N_29364,N_29434);
nor UO_837 (O_837,N_28004,N_24664);
nor UO_838 (O_838,N_25151,N_28160);
nor UO_839 (O_839,N_29375,N_28670);
nor UO_840 (O_840,N_29583,N_28922);
nor UO_841 (O_841,N_27292,N_26145);
xor UO_842 (O_842,N_25938,N_29264);
or UO_843 (O_843,N_26185,N_28871);
nor UO_844 (O_844,N_27030,N_26677);
nand UO_845 (O_845,N_24704,N_24102);
or UO_846 (O_846,N_24775,N_24557);
nand UO_847 (O_847,N_28787,N_28195);
or UO_848 (O_848,N_28466,N_27061);
xnor UO_849 (O_849,N_26042,N_28705);
or UO_850 (O_850,N_26693,N_27208);
or UO_851 (O_851,N_28176,N_27549);
and UO_852 (O_852,N_25732,N_26839);
nand UO_853 (O_853,N_24803,N_28362);
or UO_854 (O_854,N_28629,N_27042);
nor UO_855 (O_855,N_27790,N_29499);
nand UO_856 (O_856,N_29041,N_24164);
and UO_857 (O_857,N_25991,N_25954);
and UO_858 (O_858,N_25478,N_24191);
xor UO_859 (O_859,N_28905,N_29468);
nor UO_860 (O_860,N_24770,N_24013);
and UO_861 (O_861,N_24959,N_26939);
xnor UO_862 (O_862,N_28025,N_26928);
nor UO_863 (O_863,N_25383,N_25681);
xnor UO_864 (O_864,N_29842,N_29229);
xnor UO_865 (O_865,N_28000,N_25114);
or UO_866 (O_866,N_28808,N_29906);
nor UO_867 (O_867,N_27501,N_28145);
xnor UO_868 (O_868,N_25801,N_25541);
nor UO_869 (O_869,N_25980,N_29271);
or UO_870 (O_870,N_27643,N_26239);
and UO_871 (O_871,N_26198,N_29876);
and UO_872 (O_872,N_28637,N_29391);
and UO_873 (O_873,N_27619,N_24961);
or UO_874 (O_874,N_28755,N_29247);
and UO_875 (O_875,N_24167,N_24177);
nor UO_876 (O_876,N_27817,N_29863);
nor UO_877 (O_877,N_28707,N_25420);
nor UO_878 (O_878,N_27883,N_25208);
and UO_879 (O_879,N_24564,N_24224);
or UO_880 (O_880,N_24784,N_26342);
xnor UO_881 (O_881,N_25636,N_27384);
and UO_882 (O_882,N_26952,N_28644);
xnor UO_883 (O_883,N_24255,N_24678);
nor UO_884 (O_884,N_28026,N_26894);
or UO_885 (O_885,N_26529,N_29170);
and UO_886 (O_886,N_29567,N_24651);
nand UO_887 (O_887,N_26404,N_29459);
nor UO_888 (O_888,N_27305,N_27481);
and UO_889 (O_889,N_27543,N_27222);
or UO_890 (O_890,N_26167,N_28065);
or UO_891 (O_891,N_24314,N_28820);
and UO_892 (O_892,N_25041,N_29250);
and UO_893 (O_893,N_29723,N_24378);
or UO_894 (O_894,N_27671,N_27093);
nor UO_895 (O_895,N_27551,N_24630);
nand UO_896 (O_896,N_24372,N_28464);
xor UO_897 (O_897,N_26944,N_28674);
nor UO_898 (O_898,N_24692,N_29816);
nor UO_899 (O_899,N_26100,N_28712);
and UO_900 (O_900,N_26951,N_27168);
nor UO_901 (O_901,N_26066,N_26530);
nand UO_902 (O_902,N_29959,N_24928);
or UO_903 (O_903,N_26089,N_26688);
or UO_904 (O_904,N_29174,N_29305);
or UO_905 (O_905,N_25833,N_24202);
xor UO_906 (O_906,N_29678,N_26662);
nor UO_907 (O_907,N_25646,N_24214);
or UO_908 (O_908,N_27043,N_25210);
xor UO_909 (O_909,N_27147,N_26027);
and UO_910 (O_910,N_27083,N_25068);
xor UO_911 (O_911,N_29854,N_26436);
or UO_912 (O_912,N_29100,N_25439);
and UO_913 (O_913,N_27047,N_24503);
nand UO_914 (O_914,N_28532,N_29276);
and UO_915 (O_915,N_25580,N_26441);
nor UO_916 (O_916,N_27209,N_27899);
and UO_917 (O_917,N_24381,N_29200);
xnor UO_918 (O_918,N_29865,N_28174);
nor UO_919 (O_919,N_28834,N_28153);
and UO_920 (O_920,N_25625,N_27650);
nand UO_921 (O_921,N_25197,N_26712);
and UO_922 (O_922,N_26631,N_29529);
or UO_923 (O_923,N_28558,N_26000);
or UO_924 (O_924,N_27240,N_26334);
and UO_925 (O_925,N_27472,N_25592);
or UO_926 (O_926,N_27352,N_27169);
xnor UO_927 (O_927,N_26311,N_27155);
and UO_928 (O_928,N_28977,N_29736);
or UO_929 (O_929,N_29347,N_26490);
or UO_930 (O_930,N_27394,N_25244);
nand UO_931 (O_931,N_24181,N_29622);
and UO_932 (O_932,N_28107,N_25995);
and UO_933 (O_933,N_24888,N_26621);
nand UO_934 (O_934,N_27572,N_26980);
or UO_935 (O_935,N_26766,N_24213);
nand UO_936 (O_936,N_27273,N_27789);
or UO_937 (O_937,N_25424,N_25614);
nand UO_938 (O_938,N_27458,N_29005);
nand UO_939 (O_939,N_29747,N_26289);
xor UO_940 (O_940,N_25518,N_29836);
nand UO_941 (O_941,N_27656,N_25993);
and UO_942 (O_942,N_24415,N_28469);
and UO_943 (O_943,N_24298,N_27089);
and UO_944 (O_944,N_24895,N_25451);
nor UO_945 (O_945,N_24286,N_24983);
nand UO_946 (O_946,N_24808,N_29699);
nor UO_947 (O_947,N_24374,N_27692);
or UO_948 (O_948,N_28223,N_25748);
or UO_949 (O_949,N_29118,N_26018);
nand UO_950 (O_950,N_29898,N_29845);
or UO_951 (O_951,N_28094,N_28862);
and UO_952 (O_952,N_29321,N_29307);
xor UO_953 (O_953,N_26717,N_24576);
nand UO_954 (O_954,N_27829,N_25767);
nor UO_955 (O_955,N_28302,N_28907);
and UO_956 (O_956,N_26028,N_27439);
nor UO_957 (O_957,N_24583,N_26800);
nor UO_958 (O_958,N_28690,N_28164);
nor UO_959 (O_959,N_26264,N_25207);
xor UO_960 (O_960,N_26499,N_28082);
nor UO_961 (O_961,N_29367,N_28206);
and UO_962 (O_962,N_28198,N_25086);
xnor UO_963 (O_963,N_24364,N_26692);
xnor UO_964 (O_964,N_26157,N_24412);
nand UO_965 (O_965,N_29368,N_24094);
nor UO_966 (O_966,N_28954,N_29820);
nor UO_967 (O_967,N_25964,N_25318);
nor UO_968 (O_968,N_29062,N_24315);
and UO_969 (O_969,N_25967,N_27676);
and UO_970 (O_970,N_27907,N_26890);
xnor UO_971 (O_971,N_26562,N_26019);
xnor UO_972 (O_972,N_28046,N_25482);
nor UO_973 (O_973,N_25534,N_27578);
and UO_974 (O_974,N_27217,N_25092);
nor UO_975 (O_975,N_25069,N_28990);
and UO_976 (O_976,N_28548,N_29043);
xor UO_977 (O_977,N_24467,N_24146);
or UO_978 (O_978,N_27914,N_29807);
nor UO_979 (O_979,N_27835,N_26123);
nor UO_980 (O_980,N_26750,N_25648);
xnor UO_981 (O_981,N_27190,N_29143);
or UO_982 (O_982,N_24446,N_26927);
or UO_983 (O_983,N_24450,N_26533);
or UO_984 (O_984,N_27985,N_28873);
xor UO_985 (O_985,N_24464,N_28607);
or UO_986 (O_986,N_28567,N_29190);
nand UO_987 (O_987,N_27358,N_29134);
or UO_988 (O_988,N_29471,N_28238);
xor UO_989 (O_989,N_29830,N_29492);
xnor UO_990 (O_990,N_28338,N_24439);
nand UO_991 (O_991,N_25917,N_28609);
nor UO_992 (O_992,N_27020,N_27705);
xor UO_993 (O_993,N_27355,N_24758);
xor UO_994 (O_994,N_26478,N_26641);
xnor UO_995 (O_995,N_29652,N_25921);
and UO_996 (O_996,N_28693,N_24293);
nor UO_997 (O_997,N_26867,N_26869);
nor UO_998 (O_998,N_26836,N_27048);
nor UO_999 (O_999,N_24797,N_28703);
or UO_1000 (O_1000,N_27095,N_26788);
xnor UO_1001 (O_1001,N_28270,N_25141);
or UO_1002 (O_1002,N_28677,N_28888);
or UO_1003 (O_1003,N_25982,N_25556);
and UO_1004 (O_1004,N_28556,N_28752);
or UO_1005 (O_1005,N_26568,N_25717);
nor UO_1006 (O_1006,N_24957,N_26070);
and UO_1007 (O_1007,N_24549,N_26214);
xor UO_1008 (O_1008,N_27819,N_26326);
nand UO_1009 (O_1009,N_26483,N_29087);
xnor UO_1010 (O_1010,N_28620,N_27873);
nand UO_1011 (O_1011,N_27451,N_28334);
xor UO_1012 (O_1012,N_29113,N_25079);
xor UO_1013 (O_1013,N_24296,N_24008);
and UO_1014 (O_1014,N_26331,N_27111);
xor UO_1015 (O_1015,N_27653,N_25466);
nand UO_1016 (O_1016,N_29474,N_26827);
nor UO_1017 (O_1017,N_27483,N_27267);
or UO_1018 (O_1018,N_27377,N_24201);
nand UO_1019 (O_1019,N_26527,N_25755);
nor UO_1020 (O_1020,N_28289,N_29483);
or UO_1021 (O_1021,N_24348,N_24902);
nand UO_1022 (O_1022,N_29667,N_24097);
nand UO_1023 (O_1023,N_25259,N_28699);
and UO_1024 (O_1024,N_29342,N_25883);
and UO_1025 (O_1025,N_28736,N_29808);
nand UO_1026 (O_1026,N_29302,N_24936);
xnor UO_1027 (O_1027,N_28807,N_28393);
or UO_1028 (O_1028,N_26668,N_25682);
or UO_1029 (O_1029,N_24233,N_27545);
xor UO_1030 (O_1030,N_28352,N_24346);
xnor UO_1031 (O_1031,N_29334,N_28356);
nor UO_1032 (O_1032,N_24160,N_29223);
nor UO_1033 (O_1033,N_27356,N_27608);
nor UO_1034 (O_1034,N_26901,N_28169);
nor UO_1035 (O_1035,N_25071,N_24595);
xor UO_1036 (O_1036,N_26900,N_29937);
and UO_1037 (O_1037,N_29780,N_28516);
nor UO_1038 (O_1038,N_29296,N_29824);
nand UO_1039 (O_1039,N_25116,N_27710);
and UO_1040 (O_1040,N_29656,N_25342);
nand UO_1041 (O_1041,N_28912,N_25213);
or UO_1042 (O_1042,N_24788,N_27517);
nor UO_1043 (O_1043,N_27331,N_28748);
nand UO_1044 (O_1044,N_29561,N_25517);
nor UO_1045 (O_1045,N_26856,N_27632);
or UO_1046 (O_1046,N_26332,N_28899);
and UO_1047 (O_1047,N_26082,N_27864);
nor UO_1048 (O_1048,N_26591,N_28368);
xor UO_1049 (O_1049,N_25147,N_28782);
or UO_1050 (O_1050,N_28601,N_24040);
xor UO_1051 (O_1051,N_27103,N_26371);
and UO_1052 (O_1052,N_25827,N_28625);
nand UO_1053 (O_1053,N_25667,N_24647);
nor UO_1054 (O_1054,N_29444,N_27069);
or UO_1055 (O_1055,N_26084,N_25697);
and UO_1056 (O_1056,N_25293,N_27733);
nand UO_1057 (O_1057,N_28121,N_25465);
nor UO_1058 (O_1058,N_24029,N_27371);
and UO_1059 (O_1059,N_24290,N_24617);
nand UO_1060 (O_1060,N_27910,N_27694);
and UO_1061 (O_1061,N_29358,N_27459);
xnor UO_1062 (O_1062,N_27804,N_25791);
nand UO_1063 (O_1063,N_26333,N_27469);
nor UO_1064 (O_1064,N_26247,N_25136);
nor UO_1065 (O_1065,N_26243,N_25300);
or UO_1066 (O_1066,N_24274,N_29517);
and UO_1067 (O_1067,N_24633,N_25043);
nor UO_1068 (O_1068,N_26339,N_29679);
or UO_1069 (O_1069,N_28320,N_25824);
nor UO_1070 (O_1070,N_24057,N_28771);
nand UO_1071 (O_1071,N_27780,N_28377);
nor UO_1072 (O_1072,N_28740,N_25382);
nand UO_1073 (O_1073,N_29450,N_24473);
nor UO_1074 (O_1074,N_29352,N_29597);
or UO_1075 (O_1075,N_24825,N_28586);
or UO_1076 (O_1076,N_24582,N_27659);
nor UO_1077 (O_1077,N_27429,N_28735);
nor UO_1078 (O_1078,N_29881,N_29566);
nand UO_1079 (O_1079,N_28480,N_27791);
or UO_1080 (O_1080,N_24987,N_25747);
or UO_1081 (O_1081,N_28433,N_26524);
nand UO_1082 (O_1082,N_28967,N_27176);
nor UO_1083 (O_1083,N_26966,N_25427);
or UO_1084 (O_1084,N_27424,N_28222);
nand UO_1085 (O_1085,N_24599,N_27229);
and UO_1086 (O_1086,N_25120,N_29196);
nor UO_1087 (O_1087,N_26594,N_28924);
xor UO_1088 (O_1088,N_29151,N_25673);
and UO_1089 (O_1089,N_24357,N_28257);
xnor UO_1090 (O_1090,N_26118,N_24291);
xnor UO_1091 (O_1091,N_29862,N_28739);
and UO_1092 (O_1092,N_24119,N_27570);
or UO_1093 (O_1093,N_29886,N_24504);
nand UO_1094 (O_1094,N_29026,N_24203);
nor UO_1095 (O_1095,N_24631,N_27869);
and UO_1096 (O_1096,N_27712,N_24657);
xor UO_1097 (O_1097,N_24084,N_25658);
nor UO_1098 (O_1098,N_25537,N_26673);
nand UO_1099 (O_1099,N_24133,N_29509);
nand UO_1100 (O_1100,N_29657,N_24241);
nor UO_1101 (O_1101,N_27934,N_25039);
or UO_1102 (O_1102,N_28309,N_24891);
or UO_1103 (O_1103,N_26255,N_24942);
nor UO_1104 (O_1104,N_29136,N_26504);
xor UO_1105 (O_1105,N_26778,N_28367);
and UO_1106 (O_1106,N_29764,N_28569);
or UO_1107 (O_1107,N_25838,N_27332);
nand UO_1108 (O_1108,N_26120,N_26010);
nor UO_1109 (O_1109,N_25567,N_25899);
or UO_1110 (O_1110,N_26733,N_27156);
xnor UO_1111 (O_1111,N_27399,N_29791);
or UO_1112 (O_1112,N_27620,N_28535);
nor UO_1113 (O_1113,N_28014,N_29322);
xor UO_1114 (O_1114,N_28357,N_24391);
or UO_1115 (O_1115,N_27243,N_26031);
nand UO_1116 (O_1116,N_24217,N_24220);
nor UO_1117 (O_1117,N_28235,N_24301);
nand UO_1118 (O_1118,N_25496,N_29580);
and UO_1119 (O_1119,N_25929,N_27995);
nor UO_1120 (O_1120,N_26650,N_24801);
nand UO_1121 (O_1121,N_24399,N_29680);
nand UO_1122 (O_1122,N_24618,N_29033);
nand UO_1123 (O_1123,N_24074,N_27540);
and UO_1124 (O_1124,N_28732,N_25525);
or UO_1125 (O_1125,N_28661,N_24265);
nand UO_1126 (O_1126,N_27039,N_26742);
nand UO_1127 (O_1127,N_25055,N_25220);
and UO_1128 (O_1128,N_27125,N_26374);
or UO_1129 (O_1129,N_24621,N_28428);
nor UO_1130 (O_1130,N_25878,N_29077);
and UO_1131 (O_1131,N_27993,N_25735);
xnor UO_1132 (O_1132,N_24389,N_27002);
xor UO_1133 (O_1133,N_24640,N_29004);
or UO_1134 (O_1134,N_25639,N_25961);
or UO_1135 (O_1135,N_26805,N_25487);
nor UO_1136 (O_1136,N_28781,N_24806);
nand UO_1137 (O_1137,N_29537,N_28134);
nand UO_1138 (O_1138,N_24807,N_24338);
or UO_1139 (O_1139,N_25773,N_27936);
xnor UO_1140 (O_1140,N_27150,N_28742);
nand UO_1141 (O_1141,N_29740,N_27583);
and UO_1142 (O_1142,N_28069,N_29278);
nand UO_1143 (O_1143,N_28969,N_25107);
nor UO_1144 (O_1144,N_25770,N_25461);
xnor UO_1145 (O_1145,N_26794,N_26567);
xnor UO_1146 (O_1146,N_26958,N_26324);
nor UO_1147 (O_1147,N_25488,N_27737);
nor UO_1148 (O_1148,N_25262,N_28774);
and UO_1149 (O_1149,N_25061,N_29042);
or UO_1150 (O_1150,N_28441,N_26552);
and UO_1151 (O_1151,N_24049,N_26792);
and UO_1152 (O_1152,N_24016,N_26526);
xor UO_1153 (O_1153,N_27295,N_24165);
or UO_1154 (O_1154,N_29111,N_26300);
nor UO_1155 (O_1155,N_26541,N_29645);
and UO_1156 (O_1156,N_29274,N_24681);
nor UO_1157 (O_1157,N_25006,N_26102);
or UO_1158 (O_1158,N_25474,N_27149);
and UO_1159 (O_1159,N_25279,N_24284);
xor UO_1160 (O_1160,N_24401,N_26492);
or UO_1161 (O_1161,N_25865,N_25234);
and UO_1162 (O_1162,N_28483,N_24421);
xnor UO_1163 (O_1163,N_25608,N_25561);
nand UO_1164 (O_1164,N_26037,N_26090);
nor UO_1165 (O_1165,N_28138,N_24500);
or UO_1166 (O_1166,N_25704,N_28255);
xnor UO_1167 (O_1167,N_25338,N_26657);
and UO_1168 (O_1168,N_28786,N_25522);
nor UO_1169 (O_1169,N_28583,N_29841);
nand UO_1170 (O_1170,N_28226,N_25229);
or UO_1171 (O_1171,N_26377,N_25721);
or UO_1172 (O_1172,N_26419,N_24584);
and UO_1173 (O_1173,N_27260,N_29306);
nor UO_1174 (O_1174,N_28016,N_27945);
nor UO_1175 (O_1175,N_24419,N_28944);
and UO_1176 (O_1176,N_24932,N_24592);
and UO_1177 (O_1177,N_29148,N_27986);
nand UO_1178 (O_1178,N_26190,N_27298);
and UO_1179 (O_1179,N_26855,N_29160);
and UO_1180 (O_1180,N_26704,N_29176);
nor UO_1181 (O_1181,N_24762,N_29586);
xnor UO_1182 (O_1182,N_25189,N_25910);
and UO_1183 (O_1183,N_26456,N_26736);
and UO_1184 (O_1184,N_29506,N_24310);
nor UO_1185 (O_1185,N_25725,N_24607);
and UO_1186 (O_1186,N_29871,N_27727);
xnor UO_1187 (O_1187,N_26880,N_26672);
xnor UO_1188 (O_1188,N_24337,N_24992);
or UO_1189 (O_1189,N_25185,N_24064);
nand UO_1190 (O_1190,N_29551,N_27628);
nor UO_1191 (O_1191,N_24520,N_24031);
or UO_1192 (O_1192,N_29044,N_29802);
nor UO_1193 (O_1193,N_29722,N_27652);
xnor UO_1194 (O_1194,N_25699,N_26369);
and UO_1195 (O_1195,N_25918,N_29018);
or UO_1196 (O_1196,N_29730,N_24379);
xnor UO_1197 (O_1197,N_26664,N_26421);
or UO_1198 (O_1198,N_29619,N_29609);
and UO_1199 (O_1199,N_28566,N_25094);
xor UO_1200 (O_1200,N_28886,N_27686);
and UO_1201 (O_1201,N_26184,N_29412);
or UO_1202 (O_1202,N_27937,N_29088);
nand UO_1203 (O_1203,N_25626,N_29810);
nand UO_1204 (O_1204,N_29258,N_26480);
xor UO_1205 (O_1205,N_26905,N_29545);
or UO_1206 (O_1206,N_27884,N_27500);
or UO_1207 (O_1207,N_26610,N_24637);
xor UO_1208 (O_1208,N_28365,N_29767);
nand UO_1209 (O_1209,N_24717,N_24045);
and UO_1210 (O_1210,N_26026,N_28845);
and UO_1211 (O_1211,N_26970,N_29086);
or UO_1212 (O_1212,N_29293,N_28728);
or UO_1213 (O_1213,N_26761,N_24096);
and UO_1214 (O_1214,N_27616,N_28833);
nand UO_1215 (O_1215,N_26151,N_27658);
xor UO_1216 (O_1216,N_25581,N_26363);
xnor UO_1217 (O_1217,N_26361,N_26267);
and UO_1218 (O_1218,N_26651,N_24876);
nand UO_1219 (O_1219,N_26751,N_27597);
nand UO_1220 (O_1220,N_26199,N_26753);
and UO_1221 (O_1221,N_28194,N_26579);
or UO_1222 (O_1222,N_28797,N_25867);
xnor UO_1223 (O_1223,N_24705,N_26394);
xnor UO_1224 (O_1224,N_27759,N_25752);
and UO_1225 (O_1225,N_28770,N_27252);
and UO_1226 (O_1226,N_27431,N_24198);
or UO_1227 (O_1227,N_29612,N_26994);
or UO_1228 (O_1228,N_26973,N_28904);
nand UO_1229 (O_1229,N_25623,N_24171);
xnor UO_1230 (O_1230,N_27441,N_28608);
and UO_1231 (O_1231,N_24168,N_28045);
nor UO_1232 (O_1232,N_26259,N_27635);
xnor UO_1233 (O_1233,N_25689,N_25604);
and UO_1234 (O_1234,N_24639,N_28425);
nor UO_1235 (O_1235,N_24994,N_29449);
or UO_1236 (O_1236,N_29093,N_24105);
xnor UO_1237 (O_1237,N_24178,N_26277);
nand UO_1238 (O_1238,N_27960,N_24901);
xnor UO_1239 (O_1239,N_26665,N_27261);
nand UO_1240 (O_1240,N_24822,N_25436);
nand UO_1241 (O_1241,N_27286,N_27535);
or UO_1242 (O_1242,N_24812,N_26219);
xnor UO_1243 (O_1243,N_27878,N_27118);
and UO_1244 (O_1244,N_24764,N_29956);
xor UO_1245 (O_1245,N_28261,N_26397);
xnor UO_1246 (O_1246,N_25916,N_26271);
nor UO_1247 (O_1247,N_25335,N_28465);
nor UO_1248 (O_1248,N_27734,N_28140);
or UO_1249 (O_1249,N_25562,N_24147);
nand UO_1250 (O_1250,N_25077,N_27166);
xor UO_1251 (O_1251,N_26288,N_29763);
nand UO_1252 (O_1252,N_25564,N_24437);
or UO_1253 (O_1253,N_24777,N_28214);
or UO_1254 (O_1254,N_24349,N_25540);
nor UO_1255 (O_1255,N_28909,N_29925);
xnor UO_1256 (O_1256,N_29049,N_26068);
nand UO_1257 (O_1257,N_29827,N_28509);
nand UO_1258 (O_1258,N_24277,N_24966);
and UO_1259 (O_1259,N_26708,N_27776);
and UO_1260 (O_1260,N_29435,N_25848);
and UO_1261 (O_1261,N_25621,N_29332);
nand UO_1262 (O_1262,N_26513,N_27390);
nand UO_1263 (O_1263,N_26013,N_28120);
or UO_1264 (O_1264,N_25695,N_24626);
xnor UO_1265 (O_1265,N_28342,N_26532);
and UO_1266 (O_1266,N_28279,N_25600);
and UO_1267 (O_1267,N_26171,N_25641);
and UO_1268 (O_1268,N_29797,N_29978);
nor UO_1269 (O_1269,N_24083,N_24561);
xor UO_1270 (O_1270,N_27555,N_28136);
xor UO_1271 (O_1271,N_25713,N_26177);
nor UO_1272 (O_1272,N_26350,N_28146);
nor UO_1273 (O_1273,N_26789,N_27195);
nand UO_1274 (O_1274,N_24793,N_27351);
nor UO_1275 (O_1275,N_26217,N_28036);
nor UO_1276 (O_1276,N_24305,N_29071);
nor UO_1277 (O_1277,N_29950,N_25520);
xnor UO_1278 (O_1278,N_27797,N_27112);
or UO_1279 (O_1279,N_29475,N_24531);
nand UO_1280 (O_1280,N_25010,N_27708);
or UO_1281 (O_1281,N_24979,N_27184);
xor UO_1282 (O_1282,N_26015,N_29096);
nand UO_1283 (O_1283,N_28148,N_26882);
xor UO_1284 (O_1284,N_28829,N_28619);
or UO_1285 (O_1285,N_28143,N_29064);
nand UO_1286 (O_1286,N_25979,N_29201);
nor UO_1287 (O_1287,N_26721,N_27956);
or UO_1288 (O_1288,N_27104,N_25694);
or UO_1289 (O_1289,N_26816,N_28070);
or UO_1290 (O_1290,N_28618,N_28836);
or UO_1291 (O_1291,N_25677,N_26798);
nand UO_1292 (O_1292,N_29141,N_24608);
nand UO_1293 (O_1293,N_24565,N_29809);
nor UO_1294 (O_1294,N_26007,N_29019);
nand UO_1295 (O_1295,N_27265,N_26775);
and UO_1296 (O_1296,N_26683,N_27357);
nand UO_1297 (O_1297,N_24222,N_25546);
nand UO_1298 (O_1298,N_27693,N_25178);
and UO_1299 (O_1299,N_25598,N_26959);
xnor UO_1300 (O_1300,N_29422,N_29380);
nor UO_1301 (O_1301,N_28137,N_26426);
nand UO_1302 (O_1302,N_27063,N_28505);
and UO_1303 (O_1303,N_26777,N_27376);
nand UO_1304 (O_1304,N_27709,N_28401);
or UO_1305 (O_1305,N_27341,N_24447);
xor UO_1306 (O_1306,N_27966,N_28858);
nor UO_1307 (O_1307,N_28337,N_25802);
xor UO_1308 (O_1308,N_25696,N_29164);
nand UO_1309 (O_1309,N_25683,N_29979);
nand UO_1310 (O_1310,N_25034,N_26719);
nor UO_1311 (O_1311,N_28514,N_27812);
xnor UO_1312 (O_1312,N_25049,N_24325);
nand UO_1313 (O_1313,N_25571,N_28947);
nor UO_1314 (O_1314,N_28190,N_27191);
xnor UO_1315 (O_1315,N_26887,N_24819);
and UO_1316 (O_1316,N_26904,N_28119);
nor UO_1317 (O_1317,N_25022,N_28458);
or UO_1318 (O_1318,N_27977,N_28506);
nand UO_1319 (O_1319,N_28966,N_25969);
nand UO_1320 (O_1320,N_24479,N_27248);
nor UO_1321 (O_1321,N_28695,N_24140);
or UO_1322 (O_1322,N_26228,N_25105);
and UO_1323 (O_1323,N_27582,N_26780);
xor UO_1324 (O_1324,N_28776,N_28767);
nor UO_1325 (O_1325,N_29361,N_25194);
xor UO_1326 (O_1326,N_26608,N_24893);
nand UO_1327 (O_1327,N_24351,N_26274);
and UO_1328 (O_1328,N_25603,N_25425);
and UO_1329 (O_1329,N_28470,N_28547);
nor UO_1330 (O_1330,N_24900,N_29207);
xnor UO_1331 (O_1331,N_26183,N_29995);
nor UO_1332 (O_1332,N_26250,N_24030);
or UO_1333 (O_1333,N_27771,N_24615);
xor UO_1334 (O_1334,N_24886,N_24880);
or UO_1335 (O_1335,N_27826,N_26075);
nor UO_1336 (O_1336,N_28440,N_28679);
nand UO_1337 (O_1337,N_25722,N_29045);
and UO_1338 (O_1338,N_25512,N_26449);
nand UO_1339 (O_1339,N_28054,N_25886);
or UO_1340 (O_1340,N_27462,N_25578);
or UO_1341 (O_1341,N_26232,N_28098);
nor UO_1342 (O_1342,N_26306,N_26829);
and UO_1343 (O_1343,N_26842,N_27537);
and UO_1344 (O_1344,N_29514,N_27391);
or UO_1345 (O_1345,N_28479,N_27654);
xnor UO_1346 (O_1346,N_28632,N_28655);
and UO_1347 (O_1347,N_29373,N_24134);
nand UO_1348 (O_1348,N_26223,N_24721);
and UO_1349 (O_1349,N_29992,N_28155);
nor UO_1350 (O_1350,N_26093,N_26755);
and UO_1351 (O_1351,N_27599,N_26155);
xnor UO_1352 (O_1352,N_25253,N_27647);
or UO_1353 (O_1353,N_28876,N_28816);
xor UO_1354 (O_1354,N_24109,N_24866);
or UO_1355 (O_1355,N_25805,N_26774);
and UO_1356 (O_1356,N_24700,N_24868);
xor UO_1357 (O_1357,N_26583,N_28217);
xnor UO_1358 (O_1358,N_28759,N_25286);
nand UO_1359 (O_1359,N_29938,N_24051);
and UO_1360 (O_1360,N_27343,N_26576);
nor UO_1361 (O_1361,N_25361,N_28856);
xnor UO_1362 (O_1362,N_24042,N_24353);
and UO_1363 (O_1363,N_29119,N_28115);
and UO_1364 (O_1364,N_27315,N_28427);
and UO_1365 (O_1365,N_24009,N_27595);
xor UO_1366 (O_1366,N_29737,N_29079);
nand UO_1367 (O_1367,N_26059,N_27392);
xor UO_1368 (O_1368,N_24709,N_28288);
nor UO_1369 (O_1369,N_26134,N_29654);
nor UO_1370 (O_1370,N_28017,N_27679);
nand UO_1371 (O_1371,N_29904,N_29260);
and UO_1372 (O_1372,N_29672,N_29231);
xor UO_1373 (O_1373,N_26503,N_29224);
xnor UO_1374 (O_1374,N_28333,N_29949);
and UO_1375 (O_1375,N_26847,N_29903);
nand UO_1376 (O_1376,N_29720,N_27471);
nand UO_1377 (O_1377,N_26776,N_25289);
or UO_1378 (O_1378,N_24184,N_25309);
nand UO_1379 (O_1379,N_24430,N_29084);
or UO_1380 (O_1380,N_29769,N_26620);
or UO_1381 (O_1381,N_25832,N_25868);
xnor UO_1382 (O_1382,N_27194,N_29982);
or UO_1383 (O_1383,N_26463,N_29235);
nand UO_1384 (O_1384,N_27713,N_26295);
and UO_1385 (O_1385,N_25842,N_28953);
nor UO_1386 (O_1386,N_27442,N_25700);
nor UO_1387 (O_1387,N_26960,N_28681);
xor UO_1388 (O_1388,N_25390,N_27831);
nand UO_1389 (O_1389,N_29022,N_24835);
xnor UO_1390 (O_1390,N_25130,N_25797);
or UO_1391 (O_1391,N_29900,N_25230);
nor UO_1392 (O_1392,N_26883,N_26471);
and UO_1393 (O_1393,N_25630,N_27728);
xnor UO_1394 (O_1394,N_25582,N_28061);
or UO_1395 (O_1395,N_27853,N_26808);
nand UO_1396 (O_1396,N_28099,N_25216);
xor UO_1397 (O_1397,N_26156,N_27953);
and UO_1398 (O_1398,N_25710,N_26110);
xnor UO_1399 (O_1399,N_26872,N_27550);
nand UO_1400 (O_1400,N_29486,N_29739);
nand UO_1401 (O_1401,N_27770,N_27755);
or UO_1402 (O_1402,N_29794,N_29683);
nor UO_1403 (O_1403,N_29457,N_27955);
or UO_1404 (O_1404,N_26765,N_26636);
nor UO_1405 (O_1405,N_27856,N_29544);
xnor UO_1406 (O_1406,N_28122,N_27645);
nor UO_1407 (O_1407,N_28243,N_26396);
and UO_1408 (O_1408,N_28234,N_24347);
and UO_1409 (O_1409,N_25137,N_28210);
xnor UO_1410 (O_1410,N_27082,N_24820);
nor UO_1411 (O_1411,N_25698,N_27979);
xnor UO_1412 (O_1412,N_24691,N_28835);
and UO_1413 (O_1413,N_27098,N_27062);
and UO_1414 (O_1414,N_27638,N_28697);
nor UO_1415 (O_1415,N_25757,N_28937);
nor UO_1416 (O_1416,N_28486,N_27256);
or UO_1417 (O_1417,N_29031,N_26660);
xor UO_1418 (O_1418,N_29165,N_29859);
xor UO_1419 (O_1419,N_25241,N_24666);
xnor UO_1420 (O_1420,N_25779,N_26550);
nand UO_1421 (O_1421,N_29721,N_26757);
xor UO_1422 (O_1422,N_29558,N_25703);
nand UO_1423 (O_1423,N_26057,N_28702);
or UO_1424 (O_1424,N_29805,N_27952);
xor UO_1425 (O_1425,N_28443,N_26574);
xnor UO_1426 (O_1426,N_27364,N_29516);
or UO_1427 (O_1427,N_26025,N_25398);
nand UO_1428 (O_1428,N_26234,N_26073);
or UO_1429 (O_1429,N_26895,N_24093);
or UO_1430 (O_1430,N_26412,N_28200);
and UO_1431 (O_1431,N_28395,N_25650);
and UO_1432 (O_1432,N_28545,N_28869);
nand UO_1433 (O_1433,N_27321,N_25226);
or UO_1434 (O_1434,N_26431,N_25536);
xnor UO_1435 (O_1435,N_27773,N_26317);
or UO_1436 (O_1436,N_28123,N_29905);
xnor UO_1437 (O_1437,N_26773,N_24625);
xnor UO_1438 (O_1438,N_27745,N_24915);
nand UO_1439 (O_1439,N_24237,N_25337);
xnor UO_1440 (O_1440,N_27730,N_27435);
or UO_1441 (O_1441,N_26962,N_29734);
xnor UO_1442 (O_1442,N_25434,N_29089);
and UO_1443 (O_1443,N_27131,N_26937);
nor UO_1444 (O_1444,N_24143,N_24230);
nand UO_1445 (O_1445,N_25494,N_29660);
or UO_1446 (O_1446,N_25365,N_28919);
nor UO_1447 (O_1447,N_27796,N_28970);
xor UO_1448 (O_1448,N_24759,N_25764);
xor UO_1449 (O_1449,N_26875,N_24007);
and UO_1450 (O_1450,N_26510,N_27006);
nand UO_1451 (O_1451,N_25430,N_27732);
xor UO_1452 (O_1452,N_28961,N_26101);
xnor UO_1453 (O_1453,N_28477,N_27340);
nand UO_1454 (O_1454,N_26241,N_24311);
and UO_1455 (O_1455,N_29114,N_24604);
nor UO_1456 (O_1456,N_26942,N_25251);
nor UO_1457 (O_1457,N_28533,N_26690);
and UO_1458 (O_1458,N_24071,N_29489);
or UO_1459 (O_1459,N_27232,N_24670);
and UO_1460 (O_1460,N_25354,N_28669);
or UO_1461 (O_1461,N_27602,N_24344);
xnor UO_1462 (O_1462,N_24189,N_26056);
or UO_1463 (O_1463,N_25591,N_24380);
nand UO_1464 (O_1464,N_27623,N_24918);
or UO_1465 (O_1465,N_24253,N_24162);
nand UO_1466 (O_1466,N_28580,N_25778);
nor UO_1467 (O_1467,N_28957,N_26584);
xor UO_1468 (O_1468,N_29298,N_28925);
nor UO_1469 (O_1469,N_28867,N_24710);
and UO_1470 (O_1470,N_27426,N_25491);
or UO_1471 (O_1471,N_26607,N_29393);
nor UO_1472 (O_1472,N_27760,N_28220);
or UO_1473 (O_1473,N_28764,N_26464);
and UO_1474 (O_1474,N_25978,N_25219);
xor UO_1475 (O_1475,N_28147,N_27467);
nor UO_1476 (O_1476,N_26375,N_24512);
nor UO_1477 (O_1477,N_29142,N_29337);
nand UO_1478 (O_1478,N_26179,N_27180);
and UO_1479 (O_1479,N_29193,N_25350);
and UO_1480 (O_1480,N_28709,N_28943);
xor UO_1481 (O_1481,N_29443,N_26011);
or UO_1482 (O_1482,N_26729,N_24044);
xnor UO_1483 (O_1483,N_25080,N_29812);
and UO_1484 (O_1484,N_29186,N_29795);
xor UO_1485 (O_1485,N_28724,N_28229);
or UO_1486 (O_1486,N_26491,N_24494);
or UO_1487 (O_1487,N_24041,N_25288);
and UO_1488 (O_1488,N_28821,N_27609);
or UO_1489 (O_1489,N_28104,N_29503);
nand UO_1490 (O_1490,N_29376,N_26252);
or UO_1491 (O_1491,N_26617,N_28369);
and UO_1492 (O_1492,N_25036,N_24033);
nand UO_1493 (O_1493,N_24459,N_28900);
nor UO_1494 (O_1494,N_27724,N_24530);
nor UO_1495 (O_1495,N_24488,N_29040);
nor UO_1496 (O_1496,N_29890,N_24107);
xor UO_1497 (O_1497,N_25222,N_28142);
nor UO_1498 (O_1498,N_28630,N_29758);
nand UO_1499 (O_1499,N_25837,N_24297);
xor UO_1500 (O_1500,N_26984,N_27511);
nor UO_1501 (O_1501,N_29798,N_26368);
xnor UO_1502 (O_1502,N_29397,N_28330);
nor UO_1503 (O_1503,N_26563,N_24355);
xnor UO_1504 (O_1504,N_28006,N_27725);
xnor UO_1505 (O_1505,N_27765,N_29945);
nand UO_1506 (O_1506,N_28588,N_26700);
nand UO_1507 (O_1507,N_26335,N_29846);
or UO_1508 (O_1508,N_24247,N_25258);
nor UO_1509 (O_1509,N_24309,N_29092);
and UO_1510 (O_1510,N_27173,N_27806);
xnor UO_1511 (O_1511,N_25394,N_26508);
nor UO_1512 (O_1512,N_25902,N_24921);
nor UO_1513 (O_1513,N_28492,N_29108);
nand UO_1514 (O_1514,N_26076,N_25782);
nor UO_1515 (O_1515,N_24231,N_25083);
nor UO_1516 (O_1516,N_28092,N_29540);
and UO_1517 (O_1517,N_29990,N_29215);
and UO_1518 (O_1518,N_25602,N_25306);
or UO_1519 (O_1519,N_29671,N_29777);
or UO_1520 (O_1520,N_27146,N_28009);
nand UO_1521 (O_1521,N_26493,N_27337);
nor UO_1522 (O_1522,N_27072,N_25542);
nor UO_1523 (O_1523,N_26588,N_24481);
nand UO_1524 (O_1524,N_27280,N_25333);
nor UO_1525 (O_1525,N_26859,N_28824);
nor UO_1526 (O_1526,N_29920,N_24070);
xnor UO_1527 (O_1527,N_29975,N_26626);
nand UO_1528 (O_1528,N_29837,N_25750);
or UO_1529 (O_1529,N_25138,N_25273);
and UO_1530 (O_1530,N_24482,N_29304);
xor UO_1531 (O_1531,N_27157,N_25738);
or UO_1532 (O_1532,N_29560,N_26746);
xnor UO_1533 (O_1533,N_28746,N_29461);
or UO_1534 (O_1534,N_24974,N_25799);
nand UO_1535 (O_1535,N_28894,N_27314);
or UO_1536 (O_1536,N_28538,N_25861);
or UO_1537 (O_1537,N_25905,N_25052);
or UO_1538 (O_1538,N_28184,N_28084);
nor UO_1539 (O_1539,N_27868,N_27716);
and UO_1540 (O_1540,N_27323,N_29605);
nor UO_1541 (O_1541,N_24022,N_25853);
or UO_1542 (O_1542,N_26694,N_28549);
or UO_1543 (O_1543,N_28390,N_27075);
xnor UO_1544 (O_1544,N_29553,N_27277);
or UO_1545 (O_1545,N_24952,N_27601);
or UO_1546 (O_1546,N_27943,N_26592);
nand UO_1547 (O_1547,N_24728,N_25063);
nor UO_1548 (O_1548,N_29015,N_27326);
nand UO_1549 (O_1549,N_27508,N_25460);
nand UO_1550 (O_1550,N_24038,N_24695);
xnor UO_1551 (O_1551,N_28936,N_26853);
xnor UO_1552 (O_1552,N_28207,N_26505);
nor UO_1553 (O_1553,N_27911,N_26739);
nand UO_1554 (O_1554,N_29981,N_24104);
or UO_1555 (O_1555,N_27003,N_28914);
nand UO_1556 (O_1556,N_26338,N_27446);
or UO_1557 (O_1557,N_26260,N_28626);
nor UO_1558 (O_1558,N_29238,N_28109);
nor UO_1559 (O_1559,N_27743,N_26472);
xor UO_1560 (O_1560,N_29351,N_27814);
xor UO_1561 (O_1561,N_29887,N_25509);
xnor UO_1562 (O_1562,N_27140,N_24656);
nand UO_1563 (O_1563,N_29549,N_27579);
nand UO_1564 (O_1564,N_26897,N_29572);
or UO_1565 (O_1565,N_24559,N_29027);
or UO_1566 (O_1566,N_24505,N_28020);
nand UO_1567 (O_1567,N_27427,N_25597);
nor UO_1568 (O_1568,N_29458,N_24085);
nand UO_1569 (O_1569,N_25401,N_27186);
nor UO_1570 (O_1570,N_27101,N_25254);
xnor UO_1571 (O_1571,N_24195,N_26388);
nor UO_1572 (O_1572,N_25297,N_28930);
xor UO_1573 (O_1573,N_26428,N_25816);
xor UO_1574 (O_1574,N_27497,N_29901);
and UO_1575 (O_1575,N_26558,N_29685);
xor UO_1576 (O_1576,N_26038,N_24887);
xor UO_1577 (O_1577,N_27070,N_25102);
nand UO_1578 (O_1578,N_25760,N_25946);
nand UO_1579 (O_1579,N_27438,N_29997);
or UO_1580 (O_1580,N_24278,N_26262);
nor UO_1581 (O_1581,N_26104,N_26148);
nor UO_1582 (O_1582,N_29032,N_24369);
nor UO_1583 (O_1583,N_24141,N_25450);
or UO_1584 (O_1584,N_24908,N_26544);
xnor UO_1585 (O_1585,N_25935,N_26150);
nand UO_1586 (O_1586,N_25168,N_28391);
and UO_1587 (O_1587,N_25012,N_27721);
nor UO_1588 (O_1588,N_28499,N_26924);
nor UO_1589 (O_1589,N_26821,N_29522);
xnor UO_1590 (O_1590,N_25255,N_29137);
nor UO_1591 (O_1591,N_26054,N_25610);
or UO_1592 (O_1592,N_29482,N_25851);
xnor UO_1593 (O_1593,N_29156,N_29991);
nand UO_1594 (O_1594,N_29658,N_27879);
nor UO_1595 (O_1595,N_26376,N_25891);
xnor UO_1596 (O_1596,N_24135,N_27981);
nand UO_1597 (O_1597,N_27719,N_24737);
or UO_1598 (O_1598,N_25907,N_27253);
xor UO_1599 (O_1599,N_24782,N_24940);
and UO_1600 (O_1600,N_25657,N_27249);
and UO_1601 (O_1601,N_27521,N_29694);
and UO_1602 (O_1602,N_27413,N_25857);
or UO_1603 (O_1603,N_28445,N_25305);
nor UO_1604 (O_1604,N_27889,N_27751);
or UO_1605 (O_1605,N_29697,N_27603);
nand UO_1606 (O_1606,N_25268,N_29275);
and UO_1607 (O_1607,N_26517,N_26204);
nand UO_1608 (O_1608,N_24914,N_29365);
xor UO_1609 (O_1609,N_25087,N_29596);
nand UO_1610 (O_1610,N_25391,N_26415);
or UO_1611 (O_1611,N_27485,N_28170);
xor UO_1612 (O_1612,N_27828,N_25232);
nor UO_1613 (O_1613,N_26175,N_29491);
xor UO_1614 (O_1614,N_29046,N_27715);
nor UO_1615 (O_1615,N_28939,N_24885);
and UO_1616 (O_1616,N_27172,N_29894);
or UO_1617 (O_1617,N_25678,N_26130);
nand UO_1618 (O_1618,N_27171,N_27206);
nand UO_1619 (O_1619,N_29357,N_28723);
xnor UO_1620 (O_1620,N_28313,N_24544);
nor UO_1621 (O_1621,N_25994,N_24000);
xor UO_1622 (O_1622,N_26523,N_25127);
and UO_1623 (O_1623,N_28178,N_27328);
nand UO_1624 (O_1624,N_28349,N_28652);
nor UO_1625 (O_1625,N_26565,N_29569);
or UO_1626 (O_1626,N_24899,N_26950);
nor UO_1627 (O_1627,N_25311,N_28842);
xor UO_1628 (O_1628,N_29090,N_26646);
or UO_1629 (O_1629,N_29374,N_28314);
and UO_1630 (O_1630,N_29208,N_27667);
nor UO_1631 (O_1631,N_26319,N_28130);
nand UO_1632 (O_1632,N_24452,N_24813);
and UO_1633 (O_1633,N_29789,N_25125);
xnor UO_1634 (O_1634,N_27284,N_29639);
and UO_1635 (O_1635,N_27843,N_25256);
or UO_1636 (O_1636,N_28192,N_24122);
nor UO_1637 (O_1637,N_24977,N_28072);
and UO_1638 (O_1638,N_26165,N_29632);
nand UO_1639 (O_1639,N_26453,N_29742);
or UO_1640 (O_1640,N_24144,N_25642);
nand UO_1641 (O_1641,N_29140,N_27050);
nor UO_1642 (O_1642,N_27617,N_27842);
and UO_1643 (O_1643,N_27699,N_29877);
nand UO_1644 (O_1644,N_26291,N_27270);
or UO_1645 (O_1645,N_27846,N_26091);
xor UO_1646 (O_1646,N_28361,N_29445);
xor UO_1647 (O_1647,N_25340,N_24990);
and UO_1648 (O_1648,N_25702,N_29068);
nand UO_1649 (O_1649,N_24020,N_26902);
nor UO_1650 (O_1650,N_26111,N_26304);
nor UO_1651 (O_1651,N_26094,N_25976);
nor UO_1652 (O_1652,N_26012,N_28381);
and UO_1653 (O_1653,N_26210,N_29191);
or UO_1654 (O_1654,N_27959,N_28976);
nor UO_1655 (O_1655,N_26893,N_29896);
or UO_1656 (O_1656,N_24566,N_28468);
nand UO_1657 (O_1657,N_27918,N_26903);
nand UO_1658 (O_1658,N_27132,N_24821);
xor UO_1659 (O_1659,N_24919,N_29848);
nand UO_1660 (O_1660,N_28227,N_28326);
nor UO_1661 (O_1661,N_29727,N_29559);
nand UO_1662 (O_1662,N_27935,N_28364);
and UO_1663 (O_1663,N_27224,N_25821);
nor UO_1664 (O_1664,N_25813,N_25370);
and UO_1665 (O_1665,N_26099,N_25323);
xnor UO_1666 (O_1666,N_29399,N_25521);
xnor UO_1667 (O_1667,N_29518,N_26730);
nand UO_1668 (O_1668,N_24792,N_26281);
nor UO_1669 (O_1669,N_28931,N_28378);
nand UO_1670 (O_1670,N_29132,N_29348);
nor UO_1671 (O_1671,N_24845,N_26327);
nor UO_1672 (O_1672,N_24125,N_26159);
xnor UO_1673 (O_1673,N_28347,N_29121);
or UO_1674 (O_1674,N_25983,N_26936);
and UO_1675 (O_1675,N_27028,N_24904);
xor UO_1676 (O_1676,N_27263,N_26634);
nand UO_1677 (O_1677,N_24151,N_28259);
and UO_1678 (O_1678,N_25652,N_27214);
and UO_1679 (O_1679,N_27919,N_26713);
and UO_1680 (O_1680,N_26743,N_26938);
xor UO_1681 (O_1681,N_25856,N_25123);
and UO_1682 (O_1682,N_28809,N_29524);
or UO_1683 (O_1683,N_24180,N_26297);
and UO_1684 (O_1684,N_26710,N_29428);
xor UO_1685 (O_1685,N_26318,N_29550);
or UO_1686 (O_1686,N_26287,N_27741);
xnor UO_1687 (O_1687,N_27636,N_28224);
and UO_1688 (O_1688,N_27860,N_26722);
xnor UO_1689 (O_1689,N_29984,N_24393);
and UO_1690 (O_1690,N_26763,N_24690);
and UO_1691 (O_1691,N_29094,N_28241);
and UO_1692 (O_1692,N_26119,N_28482);
xor UO_1693 (O_1693,N_27983,N_25278);
nor UO_1694 (O_1694,N_24264,N_25367);
nand UO_1695 (O_1695,N_27402,N_27774);
nor UO_1696 (O_1696,N_24120,N_27009);
xor UO_1697 (O_1697,N_29219,N_27306);
nand UO_1698 (O_1698,N_24175,N_25554);
and UO_1699 (O_1699,N_24672,N_29206);
nor UO_1700 (O_1700,N_24468,N_25155);
nor UO_1701 (O_1701,N_24001,N_28584);
or UO_1702 (O_1702,N_25040,N_24073);
xnor UO_1703 (O_1703,N_25669,N_29618);
nand UO_1704 (O_1704,N_25583,N_29039);
or UO_1705 (O_1705,N_28448,N_29241);
or UO_1706 (O_1706,N_27053,N_28571);
and UO_1707 (O_1707,N_27182,N_26494);
nand UO_1708 (O_1708,N_29263,N_27272);
xnor UO_1709 (O_1709,N_25355,N_25298);
xor UO_1710 (O_1710,N_26458,N_28416);
and UO_1711 (O_1711,N_26194,N_28402);
nand UO_1712 (O_1712,N_29701,N_29389);
nand UO_1713 (O_1713,N_27834,N_24423);
xor UO_1714 (O_1714,N_24794,N_29745);
nor UO_1715 (O_1715,N_29501,N_27293);
nand UO_1716 (O_1716,N_24738,N_26230);
nand UO_1717 (O_1717,N_29874,N_28777);
xnor UO_1718 (O_1718,N_24240,N_27921);
nor UO_1719 (O_1719,N_25527,N_28543);
nor UO_1720 (O_1720,N_24851,N_28030);
nor UO_1721 (O_1721,N_27057,N_29330);
nand UO_1722 (O_1722,N_25686,N_24414);
or UO_1723 (O_1723,N_27681,N_29870);
nor UO_1724 (O_1724,N_24174,N_25743);
nor UO_1725 (O_1725,N_26764,N_27036);
nor UO_1726 (O_1726,N_28972,N_27460);
xor UO_1727 (O_1727,N_29301,N_26840);
or UO_1728 (O_1728,N_24926,N_29773);
nand UO_1729 (O_1729,N_25711,N_26854);
or UO_1730 (O_1730,N_27871,N_28380);
nor UO_1731 (O_1731,N_29104,N_28520);
nor UO_1732 (O_1732,N_25280,N_27178);
or UO_1733 (O_1733,N_28946,N_26467);
nand UO_1734 (O_1734,N_28450,N_25593);
xnor UO_1735 (O_1735,N_25794,N_26127);
and UO_1736 (O_1736,N_27099,N_26329);
and UO_1737 (O_1737,N_24859,N_27532);
and UO_1738 (O_1738,N_27646,N_24982);
nand UO_1739 (O_1739,N_29127,N_28474);
and UO_1740 (O_1740,N_28304,N_25435);
xor UO_1741 (O_1741,N_28889,N_28870);
xor UO_1742 (O_1742,N_27642,N_26178);
xnor UO_1743 (O_1743,N_26387,N_27940);
nand UO_1744 (O_1744,N_27593,N_26040);
nand UO_1745 (O_1745,N_25308,N_24718);
xor UO_1746 (O_1746,N_28318,N_27192);
xnor UO_1747 (O_1747,N_28264,N_29495);
or UO_1748 (O_1748,N_25679,N_26629);
nor UO_1749 (O_1749,N_25986,N_26947);
nand UO_1750 (O_1750,N_26678,N_27904);
xor UO_1751 (O_1751,N_28581,N_25334);
and UO_1752 (O_1752,N_25763,N_25719);
or UO_1753 (O_1753,N_24791,N_25845);
or UO_1754 (O_1754,N_24103,N_25113);
and UO_1755 (O_1755,N_24510,N_27520);
xor UO_1756 (O_1756,N_29130,N_28162);
nor UO_1757 (O_1757,N_29782,N_24689);
nor UO_1758 (O_1758,N_26832,N_27507);
nand UO_1759 (O_1759,N_24739,N_24079);
or UO_1760 (O_1760,N_25911,N_25588);
and UO_1761 (O_1761,N_27723,N_24685);
nand UO_1762 (O_1762,N_27213,N_29249);
nor UO_1763 (O_1763,N_26328,N_27560);
or UO_1764 (O_1764,N_28258,N_28067);
nand UO_1765 (O_1765,N_26507,N_29526);
and UO_1766 (O_1766,N_24076,N_26909);
nand UO_1767 (O_1767,N_26560,N_27792);
nor UO_1768 (O_1768,N_26603,N_26669);
or UO_1769 (O_1769,N_24307,N_28180);
and UO_1770 (O_1770,N_25863,N_26409);
nor UO_1771 (O_1771,N_28213,N_24698);
and UO_1772 (O_1772,N_29907,N_24118);
xnor UO_1773 (O_1773,N_25343,N_27756);
nand UO_1774 (O_1774,N_28734,N_26240);
nand UO_1775 (O_1775,N_26528,N_24207);
or UO_1776 (O_1776,N_28692,N_27294);
xnor UO_1777 (O_1777,N_28055,N_29610);
nor UO_1778 (O_1778,N_27274,N_29001);
nor UO_1779 (O_1779,N_26279,N_28392);
or UO_1780 (O_1780,N_25392,N_25042);
or UO_1781 (O_1781,N_24955,N_28097);
or UO_1782 (O_1782,N_24745,N_26152);
or UO_1783 (O_1783,N_25431,N_25384);
nor UO_1784 (O_1784,N_25359,N_26205);
xor UO_1785 (O_1785,N_25960,N_27665);
nor UO_1786 (O_1786,N_24973,N_25053);
xnor UO_1787 (O_1787,N_26457,N_28527);
nor UO_1788 (O_1788,N_29470,N_28132);
xor UO_1789 (O_1789,N_27128,N_27282);
xnor UO_1790 (O_1790,N_26891,N_28546);
nand UO_1791 (O_1791,N_25252,N_28745);
nand UO_1792 (O_1792,N_24260,N_24613);
nor UO_1793 (O_1793,N_27160,N_26619);
nand UO_1794 (O_1794,N_24249,N_26389);
nand UO_1795 (O_1795,N_24939,N_29300);
nor UO_1796 (O_1796,N_27592,N_24248);
nor UO_1797 (O_1797,N_24294,N_24802);
nand UO_1798 (O_1798,N_24156,N_26160);
nand UO_1799 (O_1799,N_24257,N_28363);
xor UO_1800 (O_1800,N_24828,N_27769);
nand UO_1801 (O_1801,N_29563,N_24659);
nand UO_1802 (O_1802,N_25553,N_28262);
nor UO_1803 (O_1803,N_29616,N_25609);
nor UO_1804 (O_1804,N_25001,N_26981);
and UO_1805 (O_1805,N_28003,N_29733);
and UO_1806 (O_1806,N_28968,N_27591);
xor UO_1807 (O_1807,N_28762,N_24985);
and UO_1808 (O_1808,N_27896,N_29512);
nor UO_1809 (O_1809,N_26868,N_29460);
or UO_1810 (O_1810,N_29833,N_28662);
xnor UO_1811 (O_1811,N_26978,N_25776);
nor UO_1812 (O_1812,N_26044,N_29864);
or UO_1813 (O_1813,N_25026,N_28103);
and UO_1814 (O_1814,N_25852,N_29282);
and UO_1815 (O_1815,N_24487,N_29327);
xnor UO_1816 (O_1816,N_29493,N_28418);
xor UO_1817 (O_1817,N_26294,N_24964);
nor UO_1818 (O_1818,N_25277,N_26454);
and UO_1819 (O_1819,N_29532,N_26132);
nand UO_1820 (O_1820,N_26752,N_28151);
and UO_1821 (O_1821,N_29013,N_28382);
and UO_1822 (O_1822,N_29147,N_27388);
and UO_1823 (O_1823,N_29860,N_25885);
nand UO_1824 (O_1824,N_25158,N_24703);
xnor UO_1825 (O_1825,N_25957,N_24336);
nand UO_1826 (O_1826,N_24492,N_25331);
nor UO_1827 (O_1827,N_25037,N_27627);
or UO_1828 (O_1828,N_29149,N_28449);
and UO_1829 (O_1829,N_24847,N_24441);
or UO_1830 (O_1830,N_29125,N_28185);
nor UO_1831 (O_1831,N_24002,N_29704);
and UO_1832 (O_1832,N_28193,N_29787);
xnor UO_1833 (O_1833,N_24724,N_28071);
nand UO_1834 (O_1834,N_29635,N_26990);
xnor UO_1835 (O_1835,N_28135,N_25595);
nor UO_1836 (O_1836,N_25473,N_26108);
or UO_1837 (O_1837,N_28593,N_25250);
and UO_1838 (O_1838,N_25109,N_26476);
nand UO_1839 (O_1839,N_28578,N_27398);
and UO_1840 (O_1840,N_27909,N_26244);
nand UO_1841 (O_1841,N_27419,N_27779);
nand UO_1842 (O_1842,N_27091,N_26067);
nor UO_1843 (O_1843,N_29277,N_28965);
or UO_1844 (O_1844,N_29525,N_25173);
nand UO_1845 (O_1845,N_29676,N_28191);
nand UO_1846 (O_1846,N_24972,N_25319);
nand UO_1847 (O_1847,N_25898,N_24611);
nand UO_1848 (O_1848,N_26168,N_26437);
and UO_1849 (O_1849,N_27640,N_25356);
and UO_1850 (O_1850,N_29790,N_24556);
nand UO_1851 (O_1851,N_25599,N_26420);
xor UO_1852 (O_1852,N_24941,N_24226);
nand UO_1853 (O_1853,N_26486,N_25217);
or UO_1854 (O_1854,N_26573,N_28916);
nor UO_1855 (O_1855,N_27493,N_25106);
or UO_1856 (O_1856,N_26963,N_28247);
nand UO_1857 (O_1857,N_29590,N_24262);
and UO_1858 (O_1858,N_26956,N_29403);
nand UO_1859 (O_1859,N_24711,N_28410);
or UO_1860 (O_1860,N_28542,N_26906);
xor UO_1861 (O_1861,N_26348,N_26444);
xor UO_1862 (O_1862,N_28063,N_26341);
xnor UO_1863 (O_1863,N_29209,N_28002);
or UO_1864 (O_1864,N_28272,N_25589);
nand UO_1865 (O_1865,N_24976,N_25404);
nand UO_1866 (O_1866,N_25296,N_24395);
xnor UO_1867 (O_1867,N_29172,N_24553);
or UO_1868 (O_1868,N_24075,N_25169);
xor UO_1869 (O_1869,N_24218,N_24161);
nor UO_1870 (O_1870,N_28539,N_28815);
nand UO_1871 (O_1871,N_29320,N_24039);
or UO_1872 (O_1872,N_26367,N_24779);
nand UO_1873 (O_1873,N_29910,N_27373);
or UO_1874 (O_1874,N_27251,N_26728);
and UO_1875 (O_1875,N_26659,N_28649);
xnor UO_1876 (O_1876,N_27598,N_29943);
xor UO_1877 (O_1877,N_27231,N_24729);
or UO_1878 (O_1878,N_24438,N_27929);
nor UO_1879 (O_1879,N_27753,N_26675);
nor UO_1880 (O_1880,N_25932,N_26440);
or UO_1881 (O_1881,N_28531,N_29541);
or UO_1882 (O_1882,N_24687,N_24798);
nor UO_1883 (O_1883,N_24445,N_25854);
or UO_1884 (O_1884,N_24186,N_26511);
nand UO_1885 (O_1885,N_25687,N_28597);
xnor UO_1886 (O_1886,N_28719,N_26735);
xnor UO_1887 (O_1887,N_25417,N_27085);
or UO_1888 (O_1888,N_29868,N_25238);
or UO_1889 (O_1889,N_25756,N_29279);
and UO_1890 (O_1890,N_26321,N_25480);
nand UO_1891 (O_1891,N_27684,N_29251);
nor UO_1892 (O_1892,N_24623,N_28665);
or UO_1893 (O_1893,N_27011,N_28452);
nand UO_1894 (O_1894,N_28882,N_25045);
and UO_1895 (O_1895,N_28627,N_24018);
nand UO_1896 (O_1896,N_24858,N_29557);
or UO_1897 (O_1897,N_29360,N_28344);
nand UO_1898 (O_1898,N_25666,N_29964);
and UO_1899 (O_1899,N_25928,N_29411);
nor UO_1900 (O_1900,N_29439,N_25152);
or UO_1901 (O_1901,N_28018,N_28802);
or UO_1902 (O_1902,N_28512,N_24006);
and UO_1903 (O_1903,N_27443,N_28819);
xnor UO_1904 (O_1904,N_28348,N_29955);
or UO_1905 (O_1905,N_29702,N_24396);
xor UO_1906 (O_1906,N_29317,N_27845);
xor UO_1907 (O_1907,N_25888,N_27016);
xnor UO_1908 (O_1908,N_24182,N_25548);
nand UO_1909 (O_1909,N_27275,N_24054);
or UO_1910 (O_1910,N_28280,N_25204);
nor UO_1911 (O_1911,N_25879,N_28299);
nor UO_1912 (O_1912,N_29857,N_29259);
or UO_1913 (O_1913,N_24733,N_26572);
nor UO_1914 (O_1914,N_29195,N_28769);
and UO_1915 (O_1915,N_29122,N_28511);
or UO_1916 (O_1916,N_29292,N_27144);
xnor UO_1917 (O_1917,N_24532,N_25047);
and UO_1918 (O_1918,N_26534,N_28758);
xor UO_1919 (O_1919,N_26697,N_28657);
and UO_1920 (O_1920,N_29578,N_25314);
nand UO_1921 (O_1921,N_28997,N_25339);
nand UO_1922 (O_1922,N_25781,N_24578);
nor UO_1923 (O_1923,N_24330,N_29350);
xnor UO_1924 (O_1924,N_29602,N_28437);
and UO_1925 (O_1925,N_28139,N_27353);
and UO_1926 (O_1926,N_27951,N_29728);
nand UO_1927 (O_1927,N_27863,N_27086);
nor UO_1928 (O_1928,N_25304,N_25464);
nand UO_1929 (O_1929,N_29829,N_29521);
and UO_1930 (O_1930,N_24300,N_26876);
xnor UO_1931 (O_1931,N_29451,N_25198);
and UO_1932 (O_1932,N_29407,N_29922);
and UO_1933 (O_1933,N_25584,N_29973);
or UO_1934 (O_1934,N_26732,N_26580);
and UO_1935 (O_1935,N_24388,N_25502);
nor UO_1936 (O_1936,N_27664,N_27912);
nor UO_1937 (O_1937,N_26381,N_26024);
xnor UO_1938 (O_1938,N_24757,N_29237);
and UO_1939 (O_1939,N_26642,N_27702);
or UO_1940 (O_1940,N_29288,N_24999);
nor UO_1941 (O_1941,N_25909,N_24223);
nor UO_1942 (O_1942,N_27175,N_29003);
and UO_1943 (O_1943,N_25874,N_26971);
nand UO_1944 (O_1944,N_29146,N_29236);
nor UO_1945 (O_1945,N_28603,N_28078);
or UO_1946 (O_1946,N_25373,N_25110);
or UO_1947 (O_1947,N_29965,N_29291);
xor UO_1948 (O_1948,N_29424,N_24432);
nor UO_1949 (O_1949,N_27670,N_24555);
nand UO_1950 (O_1950,N_28048,N_26353);
xnor UO_1951 (O_1951,N_26352,N_28910);
and UO_1952 (O_1952,N_29801,N_29709);
xor UO_1953 (O_1953,N_26920,N_29020);
and UO_1954 (O_1954,N_26115,N_24332);
nor UO_1955 (O_1955,N_24460,N_25754);
nand UO_1956 (O_1956,N_26378,N_29295);
nand UO_1957 (O_1957,N_25187,N_25448);
nand UO_1958 (O_1958,N_27225,N_27366);
nand UO_1959 (O_1959,N_26575,N_27678);
nand UO_1960 (O_1960,N_24989,N_29786);
xor UO_1961 (O_1961,N_26870,N_28274);
and UO_1962 (O_1962,N_25959,N_24484);
or UO_1963 (O_1963,N_26122,N_27802);
nand UO_1964 (O_1964,N_27610,N_29867);
and UO_1965 (O_1965,N_28980,N_28838);
or UO_1966 (O_1966,N_25505,N_27060);
nand UO_1967 (O_1967,N_27005,N_25103);
nand UO_1968 (O_1968,N_25263,N_27212);
or UO_1969 (O_1969,N_28102,N_25397);
xor UO_1970 (O_1970,N_29289,N_27389);
nor UO_1971 (O_1971,N_27237,N_29329);
nor UO_1972 (O_1972,N_26112,N_29072);
xor UO_1973 (O_1973,N_24799,N_24356);
xnor UO_1974 (O_1974,N_27478,N_24513);
nand UO_1975 (O_1975,N_27014,N_24387);
and UO_1976 (O_1976,N_26358,N_26083);
nor UO_1977 (O_1977,N_27808,N_25774);
nand UO_1978 (O_1978,N_24101,N_29202);
nor UO_1979 (O_1979,N_25759,N_26831);
nor UO_1980 (O_1980,N_26479,N_29931);
or UO_1981 (O_1981,N_27126,N_25631);
nand UO_1982 (O_1982,N_27078,N_28523);
xor UO_1983 (O_1983,N_26691,N_26163);
or UO_1984 (O_1984,N_29240,N_25161);
or UO_1985 (O_1985,N_28040,N_27903);
and UO_1986 (O_1986,N_29966,N_27615);
nor UO_1987 (O_1987,N_26187,N_28576);
xnor UO_1988 (O_1988,N_29362,N_25573);
nand UO_1989 (O_1989,N_27637,N_29804);
xor UO_1990 (O_1990,N_24129,N_25023);
nand UO_1991 (O_1991,N_29069,N_29570);
nor UO_1992 (O_1992,N_27624,N_24334);
or UO_1993 (O_1993,N_29313,N_25406);
and UO_1994 (O_1994,N_28687,N_27504);
or UO_1995 (O_1995,N_27495,N_29173);
nor UO_1996 (O_1996,N_26398,N_25516);
and UO_1997 (O_1997,N_25395,N_28741);
and UO_1998 (O_1998,N_27031,N_25221);
xor UO_1999 (O_1999,N_29400,N_26797);
or UO_2000 (O_2000,N_26932,N_29832);
nand UO_2001 (O_2001,N_25914,N_27574);
nand UO_2002 (O_2002,N_28726,N_26758);
xor UO_2003 (O_2003,N_25485,N_26992);
nor UO_2004 (O_2004,N_28563,N_29695);
xor UO_2005 (O_2005,N_24644,N_28890);
xor UO_2006 (O_2006,N_24170,N_28491);
xnor UO_2007 (O_2007,N_27361,N_25101);
and UO_2008 (O_2008,N_24463,N_24554);
nor UO_2009 (O_2009,N_28585,N_29333);
or UO_2010 (O_2010,N_29620,N_27470);
xor UO_2011 (O_2011,N_26850,N_24269);
xor UO_2012 (O_2012,N_29915,N_25862);
or UO_2013 (O_2013,N_27129,N_28340);
and UO_2014 (O_2014,N_29520,N_28066);
xor UO_2015 (O_2015,N_25847,N_27420);
nor UO_2016 (O_2016,N_29831,N_26549);
nand UO_2017 (O_2017,N_27211,N_26481);
nor UO_2018 (O_2018,N_24541,N_26830);
nand UO_2019 (O_2019,N_25121,N_25164);
and UO_2020 (O_2020,N_28572,N_26961);
or UO_2021 (O_2021,N_27329,N_28624);
nand UO_2022 (O_2022,N_29711,N_27233);
nand UO_2023 (O_2023,N_26502,N_27821);
xnor UO_2024 (O_2024,N_25275,N_26268);
and UO_2025 (O_2025,N_25357,N_24400);
or UO_2026 (O_2026,N_27900,N_27965);
nand UO_2027 (O_2027,N_29838,N_27958);
or UO_2028 (O_2028,N_28057,N_24537);
xor UO_2029 (O_2029,N_28487,N_29630);
and UO_2030 (O_2030,N_29280,N_28453);
xnor UO_2031 (O_2031,N_24098,N_25429);
nand UO_2032 (O_2032,N_27588,N_25975);
or UO_2033 (O_2033,N_25438,N_24005);
xnor UO_2034 (O_2034,N_27850,N_24742);
and UO_2035 (O_2035,N_29543,N_29012);
xnor UO_2036 (O_2036,N_26496,N_26935);
nor UO_2037 (O_2037,N_27565,N_26701);
nand UO_2038 (O_2038,N_25312,N_25618);
nand UO_2039 (O_2039,N_28493,N_24805);
nand UO_2040 (O_2040,N_24407,N_26430);
nor UO_2041 (O_2041,N_25579,N_26955);
and UO_2042 (O_2042,N_25313,N_26030);
or UO_2043 (O_2043,N_24386,N_27202);
and UO_2044 (O_2044,N_25326,N_24035);
or UO_2045 (O_2045,N_25447,N_29712);
or UO_2046 (O_2046,N_24335,N_27290);
or UO_2047 (O_2047,N_24765,N_24548);
xnor UO_2048 (O_2048,N_28553,N_25828);
nand UO_2049 (O_2049,N_29710,N_24477);
and UO_2050 (O_2050,N_25577,N_25104);
xnor UO_2051 (O_2051,N_29985,N_24078);
nor UO_2052 (O_2052,N_27319,N_24980);
nand UO_2053 (O_2053,N_26488,N_28590);
nand UO_2054 (O_2054,N_29405,N_26249);
and UO_2055 (O_2055,N_25119,N_29668);
or UO_2056 (O_2056,N_29107,N_26439);
nand UO_2057 (O_2057,N_24590,N_24323);
and UO_2058 (O_2058,N_25659,N_26176);
or UO_2059 (O_2059,N_27034,N_28423);
nand UO_2060 (O_2060,N_24649,N_28126);
nand UO_2061 (O_2061,N_27690,N_27177);
and UO_2062 (O_2062,N_26598,N_26282);
or UO_2063 (O_2063,N_29852,N_25344);
and UO_2064 (O_2064,N_29562,N_27542);
nand UO_2065 (O_2065,N_25421,N_29338);
or UO_2066 (O_2066,N_26618,N_28282);
nor UO_2067 (O_2067,N_25942,N_26769);
nand UO_2068 (O_2068,N_24970,N_26635);
or UO_2069 (O_2069,N_25349,N_29028);
and UO_2070 (O_2070,N_25247,N_24643);
or UO_2071 (O_2071,N_25664,N_29743);
nor UO_2072 (O_2072,N_29858,N_29075);
nor UO_2073 (O_2073,N_26727,N_25148);
nor UO_2074 (O_2074,N_25003,N_28388);
xnor UO_2075 (O_2075,N_24920,N_26628);
or UO_2076 (O_2076,N_25839,N_27406);
or UO_2077 (O_2077,N_28024,N_28956);
or UO_2078 (O_2078,N_28600,N_24427);
nand UO_2079 (O_2079,N_24036,N_25538);
and UO_2080 (O_2080,N_28955,N_26061);
and UO_2081 (O_2081,N_28577,N_25281);
nor UO_2082 (O_2082,N_25671,N_27445);
nor UO_2083 (O_2083,N_25919,N_28860);
nand UO_2084 (O_2084,N_29621,N_28447);
or UO_2085 (O_2085,N_26581,N_26393);
or UO_2086 (O_2086,N_25575,N_29892);
and UO_2087 (O_2087,N_29856,N_25731);
nand UO_2088 (O_2088,N_27012,N_29913);
and UO_2089 (O_2089,N_26593,N_28879);
and UO_2090 (O_2090,N_25018,N_28073);
nor UO_2091 (O_2091,N_28999,N_25934);
or UO_2092 (O_2092,N_24935,N_29266);
and UO_2093 (O_2093,N_24697,N_27587);
xnor UO_2094 (O_2094,N_25441,N_29331);
nand UO_2095 (O_2095,N_25290,N_25992);
nor UO_2096 (O_2096,N_27200,N_25134);
nand UO_2097 (O_2097,N_26313,N_26793);
nor UO_2098 (O_2098,N_28152,N_27606);
nor UO_2099 (O_2099,N_24612,N_29866);
xor UO_2100 (O_2100,N_24127,N_28747);
nor UO_2101 (O_2101,N_25294,N_28171);
xor UO_2102 (O_2102,N_28031,N_27704);
nand UO_2103 (O_2103,N_27494,N_25264);
and UO_2104 (O_2104,N_27145,N_29574);
nor UO_2105 (O_2105,N_25790,N_28766);
xnor UO_2106 (O_2106,N_27675,N_27837);
or UO_2107 (O_2107,N_24426,N_29519);
nand UO_2108 (O_2108,N_29914,N_24377);
and UO_2109 (O_2109,N_28472,N_25050);
nor UO_2110 (O_2110,N_28248,N_28478);
and UO_2111 (O_2111,N_27015,N_27383);
xnor UO_2112 (O_2112,N_26051,N_27657);
xor UO_2113 (O_2113,N_29234,N_29465);
nor UO_2114 (O_2114,N_29067,N_25376);
xor UO_2115 (O_2115,N_24894,N_28830);
xor UO_2116 (O_2116,N_26658,N_29772);
or UO_2117 (O_2117,N_26995,N_29600);
and UO_2118 (O_2118,N_29637,N_29253);
and UO_2119 (O_2119,N_27957,N_26009);
xnor UO_2120 (O_2120,N_24037,N_29187);
nand UO_2121 (O_2121,N_28727,N_29989);
nand UO_2122 (O_2122,N_29893,N_28880);
and UO_2123 (O_2123,N_26133,N_29394);
and UO_2124 (O_2124,N_24326,N_28113);
xnor UO_2125 (O_2125,N_24650,N_26991);
xnor UO_2126 (O_2126,N_24934,N_25032);
or UO_2127 (O_2127,N_26916,N_25078);
nand UO_2128 (O_2128,N_24572,N_28540);
nand UO_2129 (O_2129,N_24958,N_24443);
xnor UO_2130 (O_2130,N_28575,N_28167);
xnor UO_2131 (O_2131,N_29442,N_24968);
nand UO_2132 (O_2132,N_29899,N_25656);
or UO_2133 (O_2133,N_27523,N_28696);
xnor UO_2134 (O_2134,N_27887,N_27631);
nor UO_2135 (O_2135,N_28266,N_28672);
nand UO_2136 (O_2136,N_28932,N_24363);
xor UO_2137 (O_2137,N_29377,N_25499);
nand UO_2138 (O_2138,N_29598,N_29464);
nand UO_2139 (O_2139,N_28181,N_28689);
or UO_2140 (O_2140,N_29649,N_25375);
nor UO_2141 (O_2141,N_24750,N_24568);
nor UO_2142 (O_2142,N_29129,N_26445);
nor UO_2143 (O_2143,N_29048,N_28316);
and UO_2144 (O_2144,N_24597,N_26725);
nand UO_2145 (O_2145,N_28446,N_24773);
or UO_2146 (O_2146,N_25287,N_28029);
xnor UO_2147 (O_2147,N_28850,N_28892);
and UO_2148 (O_2148,N_26605,N_25613);
xor UO_2149 (O_2149,N_24235,N_28654);
nand UO_2150 (O_2150,N_26917,N_25019);
and UO_2151 (O_2151,N_28034,N_28187);
and UO_2152 (O_2152,N_26877,N_27742);
xor UO_2153 (O_2153,N_28554,N_27729);
nor UO_2154 (O_2154,N_28582,N_28058);
or UO_2155 (O_2155,N_25235,N_28528);
xnor UO_2156 (O_2156,N_25454,N_29105);
nand UO_2157 (O_2157,N_28182,N_25203);
nand UO_2158 (O_2158,N_29007,N_28920);
nand UO_2159 (O_2159,N_24308,N_28708);
nand UO_2160 (O_2160,N_28202,N_28935);
or UO_2161 (O_2161,N_24829,N_28106);
nor UO_2162 (O_2162,N_26796,N_26953);
xnor UO_2163 (O_2163,N_28044,N_25167);
nand UO_2164 (O_2164,N_27706,N_29642);
and UO_2165 (O_2165,N_28866,N_29303);
and UO_2166 (O_2166,N_29626,N_26384);
xor UO_2167 (O_2167,N_25691,N_29957);
nand UO_2168 (O_2168,N_29568,N_28785);
and UO_2169 (O_2169,N_24138,N_26429);
xnor UO_2170 (O_2170,N_25807,N_24574);
xor UO_2171 (O_2171,N_29759,N_29006);
nand UO_2172 (O_2172,N_29595,N_26380);
or UO_2173 (O_2173,N_27220,N_28800);
nand UO_2174 (O_2174,N_27121,N_25651);
nand UO_2175 (O_2175,N_25830,N_29035);
or UO_2176 (O_2176,N_29025,N_27354);
xor UO_2177 (O_2177,N_29942,N_27291);
xor UO_2178 (O_2178,N_26433,N_26716);
nand UO_2179 (O_2179,N_29085,N_24210);
nor UO_2180 (O_2180,N_25186,N_27801);
xor UO_2181 (O_2181,N_27077,N_27304);
xor UO_2182 (O_2182,N_24547,N_25506);
nand UO_2183 (O_2183,N_28254,N_26088);
or UO_2184 (O_2184,N_24027,N_25900);
and UO_2185 (O_2185,N_27576,N_27963);
nand UO_2186 (O_2186,N_24796,N_29221);
and UO_2187 (O_2187,N_27848,N_25768);
or UO_2188 (O_2188,N_28875,N_27142);
nand UO_2189 (O_2189,N_25936,N_26092);
or UO_2190 (O_2190,N_27219,N_29872);
or UO_2191 (O_2191,N_26106,N_27162);
and UO_2192 (O_2192,N_27123,N_25617);
nor UO_2193 (O_2193,N_26930,N_28933);
nor UO_2194 (O_2194,N_28216,N_29700);
nor UO_2195 (O_2195,N_26714,N_29014);
nor UO_2196 (O_2196,N_24884,N_28518);
or UO_2197 (O_2197,N_28105,N_27303);
xor UO_2198 (O_2198,N_25560,N_26616);
nand UO_2199 (O_2199,N_29879,N_29944);
nor UO_2200 (O_2200,N_28413,N_28631);
and UO_2201 (O_2201,N_28286,N_27584);
xor UO_2202 (O_2202,N_29823,N_24019);
xor UO_2203 (O_2203,N_27874,N_29233);
nor UO_2204 (O_2204,N_26107,N_24324);
xnor UO_2205 (O_2205,N_25184,N_27087);
nand UO_2206 (O_2206,N_29419,N_24598);
nor UO_2207 (O_2207,N_26724,N_26745);
and UO_2208 (O_2208,N_25128,N_25351);
nand UO_2209 (O_2209,N_24716,N_26551);
and UO_2210 (O_2210,N_28986,N_27300);
or UO_2211 (O_2211,N_25190,N_28295);
and UO_2212 (O_2212,N_28144,N_28481);
nand UO_2213 (O_2213,N_29971,N_24562);
xor UO_2214 (O_2214,N_29717,N_28451);
xor UO_2215 (O_2215,N_26432,N_24155);
and UO_2216 (O_2216,N_28682,N_27116);
or UO_2217 (O_2217,N_24163,N_27454);
nor UO_2218 (O_2218,N_28594,N_29770);
nand UO_2219 (O_2219,N_28421,N_25409);
nor UO_2220 (O_2220,N_29265,N_27102);
nand UO_2221 (O_2221,N_27539,N_24306);
nand UO_2222 (O_2222,N_26016,N_28560);
nand UO_2223 (O_2223,N_26666,N_27505);
and UO_2224 (O_2224,N_27696,N_26062);
nand UO_2225 (O_2225,N_25547,N_24090);
or UO_2226 (O_2226,N_29473,N_28730);
and UO_2227 (O_2227,N_28430,N_27538);
nor UO_2228 (O_2228,N_29960,N_26362);
and UO_2229 (O_2229,N_25433,N_26265);
xor UO_2230 (O_2230,N_28341,N_29592);
and UO_2231 (O_2231,N_26934,N_26988);
nor UO_2232 (O_2232,N_28240,N_26395);
nand UO_2233 (O_2233,N_26571,N_29169);
nand UO_2234 (O_2234,N_26383,N_26925);
nor UO_2235 (O_2235,N_24442,N_26795);
and UO_2236 (O_2236,N_29817,N_27330);
nand UO_2237 (O_2237,N_27296,N_29477);
xor UO_2238 (O_2238,N_29430,N_29017);
xnor UO_2239 (O_2239,N_27564,N_28339);
nor UO_2240 (O_2240,N_26173,N_24368);
or UO_2241 (O_2241,N_26050,N_25943);
nor UO_2242 (O_2242,N_24861,N_29180);
or UO_2243 (O_2243,N_29917,N_24824);
nor UO_2244 (O_2244,N_29923,N_24453);
and UO_2245 (O_2245,N_25237,N_25988);
nand UO_2246 (O_2246,N_28287,N_26898);
nor UO_2247 (O_2247,N_27258,N_27714);
xor UO_2248 (O_2248,N_25624,N_29623);
and UO_2249 (O_2249,N_27890,N_29527);
and UO_2250 (O_2250,N_24833,N_29689);
nand UO_2251 (O_2251,N_24187,N_24095);
and UO_2252 (O_2252,N_28156,N_25925);
xor UO_2253 (O_2253,N_28093,N_28711);
and UO_2254 (O_2254,N_26609,N_26416);
nand UO_2255 (O_2255,N_28296,N_27897);
or UO_2256 (O_2256,N_29843,N_27246);
nor UO_2257 (O_2257,N_29996,N_25407);
nand UO_2258 (O_2258,N_28047,N_26275);
nand UO_2259 (O_2259,N_24469,N_28881);
and UO_2260 (O_2260,N_28537,N_28885);
nor UO_2261 (O_2261,N_24480,N_25285);
and UO_2262 (O_2262,N_28718,N_27496);
xnor UO_2263 (O_2263,N_25413,N_25823);
nand UO_2264 (O_2264,N_29849,N_28041);
nor UO_2265 (O_2265,N_25532,N_26302);
nand UO_2266 (O_2266,N_24609,N_26600);
nor UO_2267 (O_2267,N_28166,N_28253);
and UO_2268 (O_2268,N_29000,N_27163);
or UO_2269 (O_2269,N_26080,N_29853);
or UO_2270 (O_2270,N_24854,N_25762);
nand UO_2271 (O_2271,N_29184,N_25175);
nand UO_2272 (O_2272,N_29839,N_26561);
and UO_2273 (O_2273,N_26337,N_25051);
and UO_2274 (O_2274,N_26095,N_24907);
xor UO_2275 (O_2275,N_26707,N_27453);
or UO_2276 (O_2276,N_27088,N_26218);
or UO_2277 (O_2277,N_29835,N_29882);
nor UO_2278 (O_2278,N_25199,N_24997);
and UO_2279 (O_2279,N_24200,N_28948);
nand UO_2280 (O_2280,N_29409,N_26633);
or UO_2281 (O_2281,N_29729,N_27514);
or UO_2282 (O_2282,N_26964,N_25380);
xnor UO_2283 (O_2283,N_28114,N_26211);
xor UO_2284 (O_2284,N_24671,N_28197);
xnor UO_2285 (O_2285,N_24384,N_25008);
or UO_2286 (O_2286,N_28731,N_28019);
or UO_2287 (O_2287,N_29082,N_27567);
and UO_2288 (O_2288,N_26599,N_29217);
or UO_2289 (O_2289,N_28273,N_28562);
nor UO_2290 (O_2290,N_24949,N_28857);
or UO_2291 (O_2291,N_28840,N_24648);
nor UO_2292 (O_2292,N_24800,N_24869);
or UO_2293 (O_2293,N_24783,N_26718);
nand UO_2294 (O_2294,N_27987,N_29211);
nand UO_2295 (O_2295,N_24434,N_29885);
or UO_2296 (O_2296,N_29395,N_29099);
nor UO_2297 (O_2297,N_28958,N_26254);
or UO_2298 (O_2298,N_25996,N_24890);
and UO_2299 (O_2299,N_25973,N_25201);
and UO_2300 (O_2300,N_28276,N_27825);
nand UO_2301 (O_2301,N_27316,N_27830);
and UO_2302 (O_2302,N_28507,N_29496);
and UO_2303 (O_2303,N_24411,N_27475);
xnor UO_2304 (O_2304,N_26085,N_26857);
xnor UO_2305 (O_2305,N_26578,N_27044);
nand UO_2306 (O_2306,N_26734,N_28079);
nor UO_2307 (O_2307,N_25715,N_29175);
xnor UO_2308 (O_2308,N_25670,N_28641);
nand UO_2309 (O_2309,N_25550,N_26767);
or UO_2310 (O_2310,N_28855,N_28574);
nand UO_2311 (O_2311,N_26060,N_28623);
xnor UO_2312 (O_2312,N_26385,N_29469);
and UO_2313 (O_2313,N_28729,N_26224);
nor UO_2314 (O_2314,N_28701,N_24087);
or UO_2315 (O_2315,N_26515,N_29053);
or UO_2316 (O_2316,N_25402,N_25611);
xor UO_2317 (O_2317,N_27680,N_26756);
xnor UO_2318 (O_2318,N_28397,N_24962);
and UO_2319 (O_2319,N_26538,N_25410);
nor UO_2320 (O_2320,N_24192,N_25135);
and UO_2321 (O_2321,N_25922,N_26604);
xnor UO_2322 (O_2322,N_24436,N_26759);
or UO_2323 (O_2323,N_25707,N_26888);
nand UO_2324 (O_2324,N_24270,N_25836);
nand UO_2325 (O_2325,N_25507,N_28463);
nor UO_2326 (O_2326,N_24428,N_26652);
nor UO_2327 (O_2327,N_25353,N_29323);
xnor UO_2328 (O_2328,N_26979,N_25093);
xnor UO_2329 (O_2329,N_27761,N_26972);
xor UO_2330 (O_2330,N_24988,N_27487);
nor UO_2331 (O_2331,N_28744,N_27629);
nand UO_2332 (O_2332,N_25844,N_28268);
nor UO_2333 (O_2333,N_24585,N_24769);
and UO_2334 (O_2334,N_26587,N_26098);
or UO_2335 (O_2335,N_27403,N_26411);
nor UO_2336 (O_2336,N_24696,N_28612);
nor UO_2337 (O_2337,N_27915,N_29873);
xor UO_2338 (O_2338,N_29144,N_29940);
nor UO_2339 (O_2339,N_29008,N_29732);
xor UO_2340 (O_2340,N_26645,N_27972);
nor UO_2341 (O_2341,N_27752,N_25841);
or UO_2342 (O_2342,N_25013,N_27515);
nand UO_2343 (O_2343,N_25150,N_28291);
or UO_2344 (O_2344,N_27718,N_26405);
nor UO_2345 (O_2345,N_25098,N_27784);
or UO_2346 (O_2346,N_28998,N_27841);
xnor UO_2347 (O_2347,N_25787,N_25974);
nand UO_2348 (O_2348,N_24840,N_27013);
xnor UO_2349 (O_2349,N_25875,N_24713);
nor UO_2350 (O_2350,N_24267,N_28988);
nor UO_2351 (O_2351,N_27661,N_28149);
xnor UO_2352 (O_2352,N_26531,N_26475);
or UO_2353 (O_2353,N_26516,N_27534);
or UO_2354 (O_2354,N_26993,N_25831);
and UO_2355 (O_2355,N_25676,N_27788);
and UO_2356 (O_2356,N_28595,N_24753);
and UO_2357 (O_2357,N_28979,N_26582);
nor UO_2358 (O_2358,N_26681,N_24004);
xnor UO_2359 (O_2359,N_27939,N_29467);
or UO_2360 (O_2360,N_27440,N_28779);
nand UO_2361 (O_2361,N_26851,N_26340);
and UO_2362 (O_2362,N_28384,N_29934);
or UO_2363 (O_2363,N_25887,N_28455);
nor UO_2364 (O_2364,N_24662,N_27159);
and UO_2365 (O_2365,N_26180,N_24502);
xnor UO_2366 (O_2366,N_24197,N_29815);
xnor UO_2367 (O_2367,N_28396,N_26364);
nand UO_2368 (O_2368,N_29299,N_27349);
xnor UO_2369 (O_2369,N_26192,N_25082);
nand UO_2370 (O_2370,N_24418,N_25649);
nand UO_2371 (O_2371,N_26301,N_29633);
or UO_2372 (O_2372,N_24790,N_24283);
or UO_2373 (O_2373,N_27557,N_27506);
nand UO_2374 (O_2374,N_25515,N_27143);
and UO_2375 (O_2375,N_27401,N_24211);
and UO_2376 (O_2376,N_27179,N_27568);
or UO_2377 (O_2377,N_28080,N_25347);
nor UO_2378 (O_2378,N_25503,N_24641);
or UO_2379 (O_2379,N_26612,N_25688);
nor UO_2380 (O_2380,N_25565,N_26466);
nand UO_2381 (O_2381,N_24466,N_29462);
or UO_2382 (O_2382,N_26143,N_25944);
nor UO_2383 (O_2383,N_29369,N_27499);
nor UO_2384 (O_2384,N_24580,N_28501);
nor UO_2385 (O_2385,N_25740,N_29312);
or UO_2386 (O_2386,N_28035,N_28023);
and UO_2387 (O_2387,N_28387,N_28992);
xor UO_2388 (O_2388,N_29948,N_27605);
nand UO_2389 (O_2389,N_27563,N_27379);
nor UO_2390 (O_2390,N_24339,N_27882);
or UO_2391 (O_2391,N_27782,N_25718);
or UO_2392 (O_2392,N_24870,N_26841);
nand UO_2393 (O_2393,N_27895,N_27924);
or UO_2394 (O_2394,N_25777,N_28173);
or UO_2395 (O_2395,N_27370,N_24680);
and UO_2396 (O_2396,N_28359,N_28496);
or UO_2397 (O_2397,N_25091,N_24055);
nand UO_2398 (O_2398,N_27276,N_25672);
or UO_2399 (O_2399,N_26285,N_26229);
and UO_2400 (O_2400,N_27228,N_25475);
or UO_2401 (O_2401,N_24221,N_28183);
or UO_2402 (O_2402,N_26201,N_25894);
or UO_2403 (O_2403,N_24771,N_25880);
or UO_2404 (O_2404,N_27065,N_26998);
nor UO_2405 (O_2405,N_29197,N_25665);
nand UO_2406 (O_2406,N_29145,N_27071);
nor UO_2407 (O_2407,N_29185,N_25594);
nor UO_2408 (O_2408,N_26804,N_29311);
or UO_2409 (O_2409,N_28372,N_29511);
nand UO_2410 (O_2410,N_27281,N_27932);
and UO_2411 (O_2411,N_26586,N_28473);
nor UO_2412 (O_2412,N_24591,N_24508);
nor UO_2413 (O_2413,N_28877,N_27482);
nand UO_2414 (O_2414,N_24622,N_26266);
and UO_2415 (O_2415,N_27547,N_28962);
nor UO_2416 (O_2416,N_25302,N_24658);
and UO_2417 (O_2417,N_25056,N_29155);
xnor UO_2418 (O_2418,N_27513,N_25004);
or UO_2419 (O_2419,N_26589,N_25972);
and UO_2420 (O_2420,N_29505,N_28407);
or UO_2421 (O_2421,N_26878,N_25744);
or UO_2422 (O_2422,N_24965,N_26807);
and UO_2423 (O_2423,N_26858,N_24863);
and UO_2424 (O_2424,N_27347,N_26815);
or UO_2425 (O_2425,N_29256,N_28251);
nor UO_2426 (O_2426,N_26469,N_26314);
and UO_2427 (O_2427,N_28743,N_27152);
or UO_2428 (O_2428,N_26539,N_29744);
or UO_2429 (O_2429,N_24390,N_24228);
or UO_2430 (O_2430,N_27613,N_26235);
or UO_2431 (O_2431,N_29587,N_24933);
nor UO_2432 (O_2432,N_24299,N_28489);
nor UO_2433 (O_2433,N_26213,N_27064);
nor UO_2434 (O_2434,N_29666,N_29783);
xnor UO_2435 (O_2435,N_26685,N_28001);
nand UO_2436 (O_2436,N_29102,N_25870);
xnor UO_2437 (O_2437,N_24457,N_28343);
and UO_2438 (O_2438,N_29926,N_27870);
nor UO_2439 (O_2439,N_29076,N_26825);
or UO_2440 (O_2440,N_28209,N_24028);
and UO_2441 (O_2441,N_28383,N_24967);
nor UO_2442 (O_2442,N_28161,N_27648);
or UO_2443 (O_2443,N_29366,N_27573);
or UO_2444 (O_2444,N_26303,N_26392);
xor UO_2445 (O_2445,N_25780,N_25884);
nand UO_2446 (O_2446,N_24853,N_28753);
or UO_2447 (O_2447,N_29800,N_24911);
nor UO_2448 (O_2448,N_27502,N_27230);
xor UO_2449 (O_2449,N_28011,N_25893);
nor UO_2450 (O_2450,N_27242,N_27046);
nand UO_2451 (O_2451,N_28108,N_27204);
and UO_2452 (O_2452,N_29643,N_24276);
xnor UO_2453 (O_2453,N_29659,N_25576);
or UO_2454 (O_2454,N_26915,N_27698);
xor UO_2455 (O_2455,N_26577,N_25393);
nand UO_2456 (O_2456,N_26372,N_29999);
nand UO_2457 (O_2457,N_29788,N_28085);
xnor UO_2458 (O_2458,N_27382,N_26487);
xnor UO_2459 (O_2459,N_24818,N_26602);
nand UO_2460 (O_2460,N_29363,N_26785);
xnor UO_2461 (O_2461,N_26649,N_24735);
xor UO_2462 (O_2462,N_25765,N_29384);
nor UO_2463 (O_2463,N_24112,N_26169);
nand UO_2464 (O_2464,N_28498,N_24993);
nand UO_2465 (O_2465,N_24354,N_26032);
and UO_2466 (O_2466,N_28846,N_29408);
nor UO_2467 (O_2467,N_26351,N_24567);
nand UO_2468 (O_2468,N_25869,N_29998);
or UO_2469 (O_2469,N_27017,N_28398);
and UO_2470 (O_2470,N_25881,N_29803);
or UO_2471 (O_2471,N_28898,N_27674);
or UO_2472 (O_2472,N_24212,N_28599);
and UO_2473 (O_2473,N_24948,N_29508);
nor UO_2474 (O_2474,N_27651,N_29670);
nand UO_2475 (O_2475,N_29755,N_26819);
and UO_2476 (O_2476,N_26519,N_26871);
nand UO_2477 (O_2477,N_24454,N_25897);
xor UO_2478 (O_2478,N_25952,N_28225);
nand UO_2479 (O_2479,N_27749,N_24856);
and UO_2480 (O_2480,N_25640,N_29855);
and UO_2481 (O_2481,N_26779,N_24947);
nor UO_2482 (O_2482,N_29061,N_24839);
xnor UO_2483 (O_2483,N_26506,N_28536);
or UO_2484 (O_2484,N_29530,N_28874);
and UO_2485 (O_2485,N_26999,N_24244);
nor UO_2486 (O_2486,N_28277,N_24072);
and UO_2487 (O_2487,N_24258,N_25985);
xor UO_2488 (O_2488,N_26193,N_24998);
and UO_2489 (O_2489,N_25712,N_29581);
nand UO_2490 (O_2490,N_26071,N_27236);
and UO_2491 (O_2491,N_26941,N_27886);
xor UO_2492 (O_2492,N_28519,N_24343);
nand UO_2493 (O_2493,N_26782,N_25479);
nand UO_2494 (O_2494,N_28307,N_29690);
nor UO_2495 (O_2495,N_25901,N_26126);
nor UO_2496 (O_2496,N_25073,N_27247);
nand UO_2497 (O_2497,N_27488,N_29888);
nor UO_2498 (O_2498,N_27250,N_27218);
nand UO_2499 (O_2499,N_25332,N_26754);
nand UO_2500 (O_2500,N_26863,N_28751);
or UO_2501 (O_2501,N_29447,N_26975);
nand UO_2502 (O_2502,N_24048,N_28794);
xor UO_2503 (O_2503,N_27524,N_25655);
nor UO_2504 (O_2504,N_27920,N_25459);
xor UO_2505 (O_2505,N_28205,N_25971);
xnor UO_2506 (O_2506,N_29080,N_25619);
nand UO_2507 (O_2507,N_25906,N_27898);
or UO_2508 (O_2508,N_28793,N_24917);
nand UO_2509 (O_2509,N_29919,N_28204);
nand UO_2510 (O_2510,N_28950,N_27408);
nor UO_2511 (O_2511,N_26425,N_26606);
or UO_2512 (O_2512,N_25310,N_28854);
xnor UO_2513 (O_2513,N_26203,N_25493);
xor UO_2514 (O_2514,N_27430,N_28331);
or UO_2515 (O_2515,N_28371,N_24865);
nand UO_2516 (O_2516,N_25956,N_24392);
nand UO_2517 (O_2517,N_24731,N_26290);
nor UO_2518 (O_2518,N_27928,N_28784);
and UO_2519 (O_2519,N_26812,N_26540);
or UO_2520 (O_2520,N_26261,N_26918);
xnor UO_2521 (O_2521,N_24465,N_25265);
and UO_2522 (O_2522,N_28294,N_25260);
and UO_2523 (O_2523,N_28116,N_26543);
nand UO_2524 (O_2524,N_25411,N_29078);
nor UO_2525 (O_2525,N_24089,N_28831);
xor UO_2526 (O_2526,N_28921,N_25341);
and UO_2527 (O_2527,N_27685,N_29024);
or UO_2528 (O_2528,N_25568,N_28129);
or UO_2529 (O_2529,N_29754,N_28323);
nand UO_2530 (O_2530,N_27731,N_27925);
nand UO_2531 (O_2531,N_26838,N_27154);
xnor UO_2532 (O_2532,N_28738,N_24157);
xor UO_2533 (O_2533,N_26648,N_24082);
and UO_2534 (O_2534,N_27226,N_27412);
nand UO_2535 (O_2535,N_25662,N_27259);
or UO_2536 (O_2536,N_26443,N_29510);
nor UO_2537 (O_2537,N_24352,N_25989);
nand UO_2538 (O_2538,N_27068,N_27822);
nor UO_2539 (O_2539,N_24620,N_24971);
xnor UO_2540 (O_2540,N_27369,N_26146);
and UO_2541 (O_2541,N_28698,N_25035);
nor UO_2542 (O_2542,N_24288,N_27257);
and UO_2543 (O_2543,N_29774,N_29030);
nand UO_2544 (O_2544,N_25829,N_24199);
and UO_2545 (O_2545,N_24706,N_25348);
and UO_2546 (O_2546,N_25530,N_25812);
xor UO_2547 (O_2547,N_28008,N_26760);
and UO_2548 (O_2548,N_27138,N_24345);
nor UO_2549 (O_2549,N_24472,N_28713);
or UO_2550 (O_2550,N_29063,N_24857);
nor UO_2551 (O_2551,N_26640,N_29507);
and UO_2552 (O_2552,N_29902,N_28414);
nor UO_2553 (O_2553,N_24406,N_28230);
nand UO_2554 (O_2554,N_27695,N_27923);
xnor UO_2555 (O_2555,N_27008,N_28436);
and UO_2556 (O_2556,N_27781,N_26596);
nand UO_2557 (O_2557,N_28399,N_25724);
or UO_2558 (O_2558,N_24588,N_28647);
xor UO_2559 (O_2559,N_29212,N_24823);
xnor UO_2560 (O_2560,N_28684,N_26379);
and UO_2561 (O_2561,N_26521,N_28685);
nor UO_2562 (O_2562,N_25789,N_24329);
nor UO_2563 (O_2563,N_24063,N_29328);
nor UO_2564 (O_2564,N_24478,N_29281);
and UO_2565 (O_2565,N_25002,N_24106);
nor UO_2566 (O_2566,N_29315,N_27244);
or UO_2567 (O_2567,N_27324,N_26087);
nor UO_2568 (O_2568,N_25193,N_25455);
nor UO_2569 (O_2569,N_25243,N_24785);
and UO_2570 (O_2570,N_28940,N_26278);
or UO_2571 (O_2571,N_25257,N_26954);
xor UO_2572 (O_2572,N_25742,N_29564);
xnor UO_2573 (O_2573,N_24304,N_29120);
nand UO_2574 (O_2574,N_27922,N_29222);
nand UO_2575 (O_2575,N_25587,N_27287);
xor UO_2576 (O_2576,N_27739,N_24975);
nand UO_2577 (O_2577,N_25632,N_25131);
xor UO_2578 (O_2578,N_24025,N_25627);
xor UO_2579 (O_2579,N_26245,N_27586);
or UO_2580 (O_2580,N_24702,N_29378);
xnor UO_2581 (O_2581,N_24877,N_29138);
or UO_2582 (O_2582,N_26136,N_29286);
nor UO_2583 (O_2583,N_29693,N_24261);
or UO_2584 (O_2584,N_24292,N_24960);
or UO_2585 (O_2585,N_25031,N_29983);
nor UO_2586 (O_2586,N_26022,N_25200);
nor UO_2587 (O_2587,N_24185,N_28550);
xnor UO_2588 (O_2588,N_26402,N_25948);
or UO_2589 (O_2589,N_26536,N_29150);
nor UO_2590 (O_2590,N_27748,N_29246);
xor UO_2591 (O_2591,N_25692,N_26907);
nand UO_2592 (O_2592,N_28510,N_29070);
xor UO_2593 (O_2593,N_27114,N_29638);
xnor UO_2594 (O_2594,N_27641,N_26706);
nor UO_2595 (O_2595,N_26908,N_27120);
and UO_2596 (O_2596,N_25283,N_26625);
nand UO_2597 (O_2597,N_24046,N_29554);
xor UO_2598 (O_2598,N_27926,N_26461);
nor UO_2599 (O_2599,N_27076,N_26655);
nor UO_2600 (O_2600,N_25629,N_27385);
nand UO_2601 (O_2601,N_24366,N_24816);
nand UO_2602 (O_2602,N_24533,N_24371);
nand UO_2603 (O_2603,N_28568,N_28817);
and UO_2604 (O_2604,N_28007,N_26923);
nand UO_2605 (O_2605,N_28150,N_28027);
xnor UO_2606 (O_2606,N_26427,N_29436);
nand UO_2607 (O_2607,N_28022,N_29309);
and UO_2608 (O_2608,N_24370,N_28405);
nand UO_2609 (O_2609,N_29796,N_24986);
nor UO_2610 (O_2610,N_24525,N_28133);
nand UO_2611 (O_2611,N_24086,N_27362);
and UO_2612 (O_2612,N_29799,N_28760);
or UO_2613 (O_2613,N_26931,N_29255);
xnor UO_2614 (O_2614,N_25240,N_29994);
or UO_2615 (O_2615,N_27241,N_28534);
nor UO_2616 (O_2616,N_24732,N_26079);
or UO_2617 (O_2617,N_29603,N_28908);
xnor UO_2618 (O_2618,N_29060,N_29178);
nor UO_2619 (O_2619,N_26365,N_25945);
nor UO_2620 (O_2620,N_26557,N_25029);
nor UO_2621 (O_2621,N_24060,N_25266);
nand UO_2622 (O_2622,N_27122,N_27092);
nor UO_2623 (O_2623,N_25414,N_25586);
nand UO_2624 (O_2624,N_26801,N_28010);
nand UO_2625 (O_2625,N_24875,N_25143);
and UO_2626 (O_2626,N_24496,N_26196);
or UO_2627 (O_2627,N_28799,N_27556);
xnor UO_2628 (O_2628,N_27035,N_24518);
nor UO_2629 (O_2629,N_29074,N_28897);
or UO_2630 (O_2630,N_26216,N_26814);
nor UO_2631 (O_2631,N_29284,N_27073);
nand UO_2632 (O_2632,N_24969,N_27989);
nor UO_2633 (O_2633,N_25419,N_26272);
or UO_2634 (O_2634,N_25908,N_24995);
nor UO_2635 (O_2635,N_27333,N_26489);
and UO_2636 (O_2636,N_27221,N_25025);
or UO_2637 (O_2637,N_28517,N_29552);
xnor UO_2638 (O_2638,N_25855,N_25097);
xor UO_2639 (O_2639,N_25784,N_27906);
xnor UO_2640 (O_2640,N_24252,N_28651);
and UO_2641 (O_2641,N_29404,N_28074);
nand UO_2642 (O_2642,N_28938,N_29725);
or UO_2643 (O_2643,N_29698,N_27950);
xnor UO_2644 (O_2644,N_29319,N_24017);
or UO_2645 (O_2645,N_26131,N_29356);
or UO_2646 (O_2646,N_29895,N_27554);
and UO_2647 (O_2647,N_27618,N_24963);
and UO_2648 (O_2648,N_29687,N_26720);
and UO_2649 (O_2649,N_28617,N_29182);
xnor UO_2650 (O_2650,N_25469,N_25205);
nand UO_2651 (O_2651,N_27079,N_28484);
xor UO_2652 (O_2652,N_26768,N_26096);
xnor UO_2653 (O_2653,N_25072,N_26638);
nand UO_2654 (O_2654,N_29203,N_26790);
xnor UO_2655 (O_2655,N_25555,N_29891);
nor UO_2656 (O_2656,N_27916,N_25212);
nand UO_2657 (O_2657,N_26864,N_24945);
or UO_2658 (O_2658,N_25321,N_28060);
and UO_2659 (O_2659,N_29706,N_24361);
xnor UO_2660 (O_2660,N_27432,N_26055);
nor UO_2661 (O_2661,N_28400,N_29617);
nand UO_2662 (O_2662,N_29611,N_29058);
nand UO_2663 (O_2663,N_26153,N_27827);
xnor UO_2664 (O_2664,N_27338,N_28050);
or UO_2665 (O_2665,N_25858,N_26861);
and UO_2666 (O_2666,N_29297,N_26547);
xor UO_2667 (O_2667,N_28212,N_26845);
nor UO_2668 (O_2668,N_24236,N_24653);
and UO_2669 (O_2669,N_29269,N_25096);
or UO_2670 (O_2670,N_26520,N_27818);
nor UO_2671 (O_2671,N_27205,N_25122);
and UO_2672 (O_2672,N_25456,N_28232);
xor UO_2673 (O_2673,N_28154,N_24362);
and UO_2674 (O_2674,N_26049,N_25806);
and UO_2675 (O_2675,N_26162,N_28462);
nand UO_2676 (O_2676,N_27982,N_24282);
or UO_2677 (O_2677,N_27876,N_25062);
nor UO_2678 (O_2678,N_24602,N_28722);
nand UO_2679 (O_2679,N_24521,N_26723);
or UO_2680 (O_2680,N_24499,N_25295);
nor UO_2681 (O_2681,N_24996,N_25301);
nor UO_2682 (O_2682,N_24416,N_25663);
nor UO_2683 (O_2683,N_27861,N_25209);
and UO_2684 (O_2684,N_27607,N_27840);
nor UO_2685 (O_2685,N_27600,N_24780);
xnor UO_2686 (O_2686,N_28952,N_26242);
xnor UO_2687 (O_2687,N_27630,N_27363);
and UO_2688 (O_2688,N_25769,N_26559);
nand UO_2689 (O_2689,N_25519,N_29875);
or UO_2690 (O_2690,N_24634,N_26417);
and UO_2691 (O_2691,N_24501,N_28844);
nor UO_2692 (O_2692,N_26865,N_26072);
and UO_2693 (O_2693,N_25027,N_29970);
and UO_2694 (O_2694,N_24404,N_26422);
xor UO_2695 (O_2695,N_28062,N_24409);
nor UO_2696 (O_2696,N_26689,N_27589);
or UO_2697 (O_2697,N_27668,N_29243);
or UO_2698 (O_2698,N_29213,N_24150);
nor UO_2699 (O_2699,N_26791,N_28872);
or UO_2700 (O_2700,N_24536,N_25497);
nor UO_2701 (O_2701,N_29822,N_24204);
and UO_2702 (O_2702,N_28124,N_27581);
nor UO_2703 (O_2703,N_24701,N_27018);
xnor UO_2704 (O_2704,N_28179,N_24015);
xnor UO_2705 (O_2705,N_25968,N_24486);
xor UO_2706 (O_2706,N_24669,N_29220);
or UO_2707 (O_2707,N_28822,N_27019);
nor UO_2708 (O_2708,N_25328,N_25442);
nor UO_2709 (O_2709,N_25734,N_28650);
nor UO_2710 (O_2710,N_27396,N_24726);
and UO_2711 (O_2711,N_27990,N_29547);
and UO_2712 (O_2712,N_29705,N_28110);
or UO_2713 (O_2713,N_27998,N_28934);
or UO_2714 (O_2714,N_26139,N_28706);
xnor UO_2715 (O_2715,N_29192,N_29958);
nand UO_2716 (O_2716,N_27561,N_28714);
or UO_2717 (O_2717,N_29771,N_25452);
and UO_2718 (O_2718,N_28460,N_25693);
nand UO_2719 (O_2719,N_29651,N_28290);
xor UO_2720 (O_2720,N_25643,N_29123);
and UO_2721 (O_2721,N_26253,N_25270);
or UO_2722 (O_2722,N_24929,N_24317);
xnor UO_2723 (O_2723,N_29655,N_27548);
and UO_2724 (O_2724,N_27807,N_24600);
nand UO_2725 (O_2725,N_25272,N_29433);
and UO_2726 (O_2726,N_28049,N_28434);
xor UO_2727 (O_2727,N_29423,N_25931);
xnor UO_2728 (O_2728,N_26940,N_27463);
or UO_2729 (O_2729,N_28526,N_27954);
nand UO_2730 (O_2730,N_27530,N_29429);
and UO_2731 (O_2731,N_29818,N_27875);
or UO_2732 (O_2732,N_24032,N_29778);
nor UO_2733 (O_2733,N_25873,N_29761);
nor UO_2734 (O_2734,N_29139,N_25933);
or UO_2735 (O_2735,N_26921,N_25028);
or UO_2736 (O_2736,N_28773,N_24458);
nor UO_2737 (O_2737,N_29636,N_25987);
nand UO_2738 (O_2738,N_24065,N_25545);
nand UO_2739 (O_2739,N_26345,N_26843);
nor UO_2740 (O_2740,N_26969,N_27133);
nand UO_2741 (O_2741,N_26772,N_29908);
and UO_2742 (O_2742,N_29054,N_24991);
and UO_2743 (O_2743,N_27525,N_27189);
nand UO_2744 (O_2744,N_27785,N_28555);
nand UO_2745 (O_2745,N_24596,N_29021);
nor UO_2746 (O_2746,N_24225,N_27522);
or UO_2747 (O_2747,N_24271,N_28052);
nor UO_2748 (O_2748,N_26189,N_25511);
nand UO_2749 (O_2749,N_27148,N_26509);
xor UO_2750 (O_2750,N_28502,N_24340);
or UO_2751 (O_2751,N_29752,N_28683);
or UO_2752 (O_2752,N_24128,N_27683);
and UO_2753 (O_2753,N_24011,N_25951);
xor UO_2754 (O_2754,N_28345,N_24528);
nor UO_2755 (O_2755,N_28439,N_28394);
or UO_2756 (O_2756,N_28796,N_25889);
nor UO_2757 (O_2757,N_26705,N_25225);
and UO_2758 (O_2758,N_28159,N_29631);
xor UO_2759 (O_2759,N_28037,N_27747);
and UO_2760 (O_2760,N_24509,N_27516);
and UO_2761 (O_2761,N_28671,N_25999);
xor UO_2762 (O_2762,N_24694,N_24581);
nand UO_2763 (O_2763,N_27794,N_24872);
nor UO_2764 (O_2764,N_24117,N_25327);
nor UO_2765 (O_2765,N_25638,N_27893);
nand UO_2766 (O_2766,N_24534,N_29128);
nor UO_2767 (O_2767,N_24281,N_28853);
and UO_2768 (O_2768,N_24916,N_25416);
or UO_2769 (O_2769,N_24593,N_29227);
or UO_2770 (O_2770,N_28500,N_25749);
and UO_2771 (O_2771,N_27594,N_26202);
and UO_2772 (O_2772,N_25467,N_27994);
or UO_2773 (O_2773,N_25364,N_29066);
xnor UO_2774 (O_2774,N_29036,N_29897);
or UO_2775 (O_2775,N_27491,N_28832);
nor UO_2776 (O_2776,N_24846,N_28219);
or UO_2777 (O_2777,N_25570,N_25937);
and UO_2778 (O_2778,N_24906,N_28319);
and UO_2779 (O_2779,N_25741,N_27264);
or UO_2780 (O_2780,N_29414,N_25690);
xor UO_2781 (O_2781,N_26158,N_29498);
nor UO_2782 (O_2782,N_27234,N_29448);
and UO_2783 (O_2783,N_24848,N_26399);
nand UO_2784 (O_2784,N_25737,N_25675);
and UO_2785 (O_2785,N_27866,N_28605);
xnor UO_2786 (O_2786,N_24774,N_29157);
or UO_2787 (O_2787,N_24279,N_26542);
or UO_2788 (O_2788,N_27992,N_27809);
nor UO_2789 (O_2789,N_25495,N_24768);
and UO_2790 (O_2790,N_25249,N_24881);
and UO_2791 (O_2791,N_27905,N_26413);
or UO_2792 (O_2792,N_27988,N_24405);
nor UO_2793 (O_2793,N_29889,N_25095);
nor UO_2794 (O_2794,N_27334,N_25211);
and UO_2795 (O_2795,N_29748,N_24142);
or UO_2796 (O_2796,N_28640,N_29930);
nor UO_2797 (O_2797,N_29757,N_27421);
or UO_2798 (O_2798,N_27181,N_24475);
or UO_2799 (O_2799,N_25292,N_24375);
nor UO_2800 (O_2800,N_27037,N_25653);
xnor UO_2801 (O_2801,N_27227,N_26207);
nand UO_2802 (O_2802,N_27436,N_27476);
xnor UO_2803 (O_2803,N_24815,N_28244);
nor UO_2804 (O_2804,N_24456,N_24545);
or UO_2805 (O_2805,N_26256,N_24817);
nor UO_2806 (O_2806,N_24610,N_24495);
nand UO_2807 (O_2807,N_25924,N_29921);
nor UO_2808 (O_2808,N_27187,N_24526);
nor UO_2809 (O_2809,N_29861,N_28231);
xnor UO_2810 (O_2810,N_26308,N_29515);
and UO_2811 (O_2811,N_26140,N_27757);
or UO_2812 (O_2812,N_25708,N_27170);
or UO_2813 (O_2813,N_28981,N_27301);
xnor UO_2814 (O_2814,N_26215,N_25470);
or UO_2815 (O_2815,N_25998,N_29037);
or UO_2816 (O_2816,N_24538,N_28403);
and UO_2817 (O_2817,N_25223,N_26041);
or UO_2818 (O_2818,N_29431,N_25615);
or UO_2819 (O_2819,N_28611,N_29065);
xnor UO_2820 (O_2820,N_26149,N_26985);
xnor UO_2821 (O_2821,N_27238,N_27279);
xnor UO_2822 (O_2822,N_26221,N_28915);
nor UO_2823 (O_2823,N_29677,N_26512);
and UO_2824 (O_2824,N_24250,N_26276);
nor UO_2825 (O_2825,N_29538,N_25644);
and UO_2826 (O_2826,N_29267,N_29353);
or UO_2827 (O_2827,N_26663,N_28406);
and UO_2828 (O_2828,N_29650,N_27787);
nand UO_2829 (O_2829,N_25412,N_26017);
nand UO_2830 (O_2830,N_28675,N_24873);
xnor UO_2831 (O_2831,N_29354,N_24410);
and UO_2832 (O_2832,N_24058,N_29624);
nand UO_2833 (O_2833,N_25915,N_24158);
nor UO_2834 (O_2834,N_26555,N_24238);
xor UO_2835 (O_2835,N_26452,N_26896);
xnor UO_2836 (O_2836,N_29565,N_25423);
nand UO_2837 (O_2837,N_29765,N_28283);
or UO_2838 (O_2838,N_28587,N_29969);
nor UO_2839 (O_2839,N_25196,N_27375);
nand UO_2840 (O_2840,N_26181,N_28989);
xnor UO_2841 (O_2841,N_24519,N_28415);
xor UO_2842 (O_2842,N_27074,N_24498);
xor UO_2843 (O_2843,N_27433,N_29500);
nor UO_2844 (O_2844,N_27973,N_28795);
and UO_2845 (O_2845,N_26485,N_24514);
xor UO_2846 (O_2846,N_25463,N_26820);
or UO_2847 (O_2847,N_24014,N_25154);
nand UO_2848 (O_2848,N_27566,N_26195);
nor UO_2849 (O_2849,N_29707,N_24946);
xor UO_2850 (O_2850,N_24043,N_26886);
or UO_2851 (O_2851,N_29571,N_28963);
and UO_2852 (O_2852,N_25381,N_27283);
xor UO_2853 (O_2853,N_29387,N_26036);
xnor UO_2854 (O_2854,N_27562,N_28991);
xor UO_2855 (O_2855,N_27833,N_27766);
or UO_2856 (O_2856,N_25011,N_27434);
or UO_2857 (O_2857,N_26161,N_27410);
nand UO_2858 (O_2858,N_25379,N_27970);
or UO_2859 (O_2859,N_28868,N_29205);
or UO_2860 (O_2860,N_27106,N_29513);
and UO_2861 (O_2861,N_26048,N_27201);
and UO_2862 (O_2862,N_24080,N_25428);
or UO_2863 (O_2863,N_24188,N_29359);
xnor UO_2864 (O_2864,N_25601,N_28422);
and UO_2865 (O_2865,N_29163,N_26537);
and UO_2866 (O_2866,N_25566,N_25358);
or UO_2867 (O_2867,N_29935,N_28666);
nand UO_2868 (O_2868,N_29927,N_26885);
xor UO_2869 (O_2869,N_24081,N_25811);
nor UO_2870 (O_2870,N_25386,N_27137);
or UO_2871 (O_2871,N_29961,N_27777);
xnor UO_2872 (O_2872,N_29485,N_28949);
xnor UO_2873 (O_2873,N_26269,N_26170);
and UO_2874 (O_2874,N_29051,N_25819);
nand UO_2875 (O_2875,N_28346,N_28128);
xor UO_2876 (O_2876,N_29273,N_24360);
nor UO_2877 (O_2877,N_25307,N_29427);
or UO_2878 (O_2878,N_26498,N_27339);
nand UO_2879 (O_2879,N_26590,N_29440);
xor UO_2880 (O_2880,N_28351,N_24852);
or UO_2881 (O_2881,N_25866,N_29029);
nand UO_2882 (O_2882,N_24497,N_24540);
or UO_2883 (O_2883,N_25140,N_29947);
and UO_2884 (O_2884,N_28974,N_26696);
nand UO_2885 (O_2885,N_26047,N_27448);
xnor UO_2886 (O_2886,N_29415,N_27720);
nor UO_2887 (O_2887,N_25500,N_29453);
nand UO_2888 (O_2888,N_24206,N_28801);
nand UO_2889 (O_2889,N_28228,N_25195);
or UO_2890 (O_2890,N_26611,N_29244);
nor UO_2891 (O_2891,N_26747,N_27536);
and UO_2892 (O_2892,N_28172,N_29268);
nand UO_2893 (O_2893,N_25372,N_28315);
or UO_2894 (O_2894,N_24259,N_24635);
nand UO_2895 (O_2895,N_28825,N_24860);
nand UO_2896 (O_2896,N_25389,N_24558);
nand UO_2897 (O_2897,N_27697,N_28884);
or UO_2898 (O_2898,N_26682,N_26459);
nor UO_2899 (O_2899,N_25165,N_29828);
or UO_2900 (O_2900,N_27335,N_25590);
or UO_2901 (O_2901,N_24012,N_26231);
nor UO_2902 (O_2902,N_25016,N_27810);
and UO_2903 (O_2903,N_26035,N_29371);
or UO_2904 (O_2904,N_24754,N_25058);
or UO_2905 (O_2905,N_26257,N_25471);
or UO_2906 (O_2906,N_24091,N_28308);
nor UO_2907 (O_2907,N_27096,N_28157);
xor UO_2908 (O_2908,N_25904,N_26653);
xor UO_2909 (O_2909,N_24367,N_26518);
or UO_2910 (O_2910,N_29663,N_29381);
nor UO_2911 (O_2911,N_24516,N_24327);
or UO_2912 (O_2912,N_28806,N_29388);
nand UO_2913 (O_2913,N_27980,N_24638);
and UO_2914 (O_2914,N_26008,N_24062);
nor UO_2915 (O_2915,N_29162,N_27309);
nor UO_2916 (O_2916,N_28918,N_24889);
nand UO_2917 (O_2917,N_27254,N_24136);
nor UO_2918 (O_2918,N_26357,N_26382);
nand UO_2919 (O_2919,N_26182,N_28101);
xnor UO_2920 (O_2920,N_27486,N_29124);
and UO_2921 (O_2921,N_27877,N_29425);
and UO_2922 (O_2922,N_27136,N_26744);
nor UO_2923 (O_2923,N_25761,N_24402);
or UO_2924 (O_2924,N_28851,N_25552);
xor UO_2925 (O_2925,N_25363,N_29941);
nor UO_2926 (O_2926,N_24088,N_25490);
xor UO_2927 (O_2927,N_27318,N_29909);
nand UO_2928 (O_2928,N_26424,N_28841);
and UO_2929 (O_2929,N_28373,N_24722);
xnor UO_2930 (O_2930,N_27978,N_24587);
or UO_2931 (O_2931,N_26208,N_25144);
xnor UO_2932 (O_2932,N_25882,N_27457);
nand UO_2933 (O_2933,N_25020,N_25637);
nor UO_2934 (O_2934,N_28332,N_25808);
nand UO_2935 (O_2935,N_27271,N_27239);
nor UO_2936 (O_2936,N_27569,N_28716);
or UO_2937 (O_2937,N_28653,N_26818);
nor UO_2938 (O_2938,N_24216,N_29177);
and UO_2939 (O_2939,N_27691,N_24767);
or UO_2940 (O_2940,N_29673,N_25739);
or UO_2941 (O_2941,N_28515,N_29977);
nor UO_2942 (O_2942,N_24795,N_29109);
nor UO_2943 (O_2943,N_27108,N_26613);
or UO_2944 (O_2944,N_26336,N_28606);
nor UO_2945 (O_2945,N_28778,N_29452);
xnor UO_2946 (O_2946,N_29341,N_25009);
or UO_2947 (O_2947,N_28127,N_25843);
nor UO_2948 (O_2948,N_24878,N_28467);
and UO_2949 (O_2949,N_24756,N_29814);
nand UO_2950 (O_2950,N_25476,N_28175);
xor UO_2951 (O_2951,N_25329,N_25804);
or UO_2952 (O_2952,N_25005,N_25751);
xnor UO_2953 (O_2953,N_28667,N_26386);
and UO_2954 (O_2954,N_28053,N_27158);
nor UO_2955 (O_2955,N_25117,N_24950);
nand UO_2956 (O_2956,N_27325,N_25132);
or UO_2957 (O_2957,N_26154,N_28188);
nor UO_2958 (O_2958,N_27917,N_24551);
xor UO_2959 (O_2959,N_26343,N_26833);
nand UO_2960 (O_2960,N_28298,N_24628);
xor UO_2961 (O_2961,N_24605,N_26346);
nor UO_2962 (O_2962,N_28847,N_24523);
and UO_2963 (O_2963,N_27997,N_26086);
or UO_2964 (O_2964,N_28614,N_26676);
and UO_2965 (O_2965,N_27000,N_24321);
and UO_2966 (O_2966,N_25202,N_26446);
xor UO_2967 (O_2967,N_27418,N_26323);
and UO_2968 (O_2968,N_26849,N_25896);
and UO_2969 (O_2969,N_29546,N_28075);
nand UO_2970 (O_2970,N_28141,N_27673);
xnor UO_2971 (O_2971,N_28524,N_26391);
nor UO_2972 (O_2972,N_26033,N_28321);
or UO_2973 (O_2973,N_24318,N_25840);
and UO_2974 (O_2974,N_24550,N_26081);
nand UO_2975 (O_2975,N_27799,N_29290);
nand UO_2976 (O_2976,N_29735,N_27320);
or UO_2977 (O_2977,N_29406,N_24838);
and UO_2978 (O_2978,N_27885,N_25181);
xnor UO_2979 (O_2979,N_27931,N_24855);
nand UO_2980 (O_2980,N_27854,N_27888);
nor UO_2981 (O_2981,N_25504,N_28038);
or UO_2982 (O_2982,N_25170,N_25388);
nand UO_2983 (O_2983,N_26630,N_27867);
or UO_2984 (O_2984,N_26595,N_29641);
xor UO_2985 (O_2985,N_26006,N_24451);
nor UO_2986 (O_2986,N_29478,N_27308);
nand UO_2987 (O_2987,N_24130,N_26826);
or UO_2988 (O_2988,N_26912,N_27689);
xor UO_2989 (O_2989,N_27677,N_24455);
nor UO_2990 (O_2990,N_26370,N_26283);
nor UO_2991 (O_2991,N_25984,N_27942);
nor UO_2992 (O_2992,N_27902,N_29370);
nor UO_2993 (O_2993,N_24809,N_24196);
nand UO_2994 (O_2994,N_29490,N_24539);
nor UO_2995 (O_2995,N_27527,N_27644);
nor UO_2996 (O_2996,N_26053,N_28951);
and UO_2997 (O_2997,N_29345,N_29980);
or UO_2998 (O_2998,N_27775,N_29731);
or UO_2999 (O_2999,N_29993,N_26987);
xnor UO_3000 (O_3000,N_28692,N_25245);
and UO_3001 (O_3001,N_26146,N_26782);
nand UO_3002 (O_3002,N_28341,N_26580);
or UO_3003 (O_3003,N_24480,N_27227);
and UO_3004 (O_3004,N_24034,N_24488);
nand UO_3005 (O_3005,N_27942,N_28327);
xor UO_3006 (O_3006,N_26350,N_29190);
nand UO_3007 (O_3007,N_26412,N_29605);
or UO_3008 (O_3008,N_25352,N_24363);
xor UO_3009 (O_3009,N_28981,N_28123);
xnor UO_3010 (O_3010,N_28107,N_25864);
nand UO_3011 (O_3011,N_27453,N_27006);
or UO_3012 (O_3012,N_26831,N_25729);
and UO_3013 (O_3013,N_24063,N_25863);
nand UO_3014 (O_3014,N_24890,N_28927);
nand UO_3015 (O_3015,N_27297,N_28056);
nor UO_3016 (O_3016,N_26335,N_26482);
nand UO_3017 (O_3017,N_29863,N_24226);
xnor UO_3018 (O_3018,N_24293,N_26852);
nor UO_3019 (O_3019,N_24702,N_26211);
xnor UO_3020 (O_3020,N_24523,N_28926);
or UO_3021 (O_3021,N_28130,N_27244);
nor UO_3022 (O_3022,N_28238,N_26384);
or UO_3023 (O_3023,N_27854,N_28106);
or UO_3024 (O_3024,N_24047,N_24035);
and UO_3025 (O_3025,N_24584,N_29047);
and UO_3026 (O_3026,N_26172,N_27900);
xnor UO_3027 (O_3027,N_26880,N_28450);
nor UO_3028 (O_3028,N_27671,N_26307);
xnor UO_3029 (O_3029,N_25223,N_27699);
and UO_3030 (O_3030,N_26185,N_26803);
xnor UO_3031 (O_3031,N_27675,N_26325);
nand UO_3032 (O_3032,N_27573,N_28628);
nor UO_3033 (O_3033,N_26082,N_28212);
xnor UO_3034 (O_3034,N_29098,N_27675);
nand UO_3035 (O_3035,N_25276,N_29239);
nand UO_3036 (O_3036,N_27260,N_28691);
nand UO_3037 (O_3037,N_28583,N_25976);
or UO_3038 (O_3038,N_25733,N_29387);
xnor UO_3039 (O_3039,N_27250,N_28446);
nand UO_3040 (O_3040,N_28780,N_25477);
nand UO_3041 (O_3041,N_27869,N_29840);
nand UO_3042 (O_3042,N_28599,N_24964);
xor UO_3043 (O_3043,N_28324,N_26823);
and UO_3044 (O_3044,N_25448,N_26619);
nor UO_3045 (O_3045,N_25778,N_27155);
nand UO_3046 (O_3046,N_28269,N_29817);
xor UO_3047 (O_3047,N_25514,N_28088);
nand UO_3048 (O_3048,N_29608,N_29110);
or UO_3049 (O_3049,N_26084,N_27418);
nor UO_3050 (O_3050,N_28268,N_27884);
xor UO_3051 (O_3051,N_24353,N_27717);
nand UO_3052 (O_3052,N_26207,N_27645);
or UO_3053 (O_3053,N_27440,N_25788);
or UO_3054 (O_3054,N_29668,N_27934);
nand UO_3055 (O_3055,N_25780,N_24003);
xor UO_3056 (O_3056,N_25573,N_26372);
nor UO_3057 (O_3057,N_27252,N_27525);
nor UO_3058 (O_3058,N_24301,N_27699);
or UO_3059 (O_3059,N_27655,N_24621);
and UO_3060 (O_3060,N_28921,N_27671);
or UO_3061 (O_3061,N_29186,N_25223);
or UO_3062 (O_3062,N_25353,N_28637);
or UO_3063 (O_3063,N_27514,N_26444);
xnor UO_3064 (O_3064,N_25940,N_24191);
xnor UO_3065 (O_3065,N_25661,N_28068);
and UO_3066 (O_3066,N_28333,N_24926);
and UO_3067 (O_3067,N_26060,N_26930);
nor UO_3068 (O_3068,N_25683,N_29845);
nand UO_3069 (O_3069,N_26276,N_27555);
nand UO_3070 (O_3070,N_26708,N_25202);
nand UO_3071 (O_3071,N_26952,N_28641);
xnor UO_3072 (O_3072,N_27197,N_28063);
and UO_3073 (O_3073,N_27815,N_25471);
or UO_3074 (O_3074,N_24701,N_26147);
xor UO_3075 (O_3075,N_25619,N_26313);
xnor UO_3076 (O_3076,N_26926,N_29393);
nor UO_3077 (O_3077,N_27305,N_26444);
nor UO_3078 (O_3078,N_28030,N_29048);
xnor UO_3079 (O_3079,N_24139,N_27206);
xnor UO_3080 (O_3080,N_29188,N_25732);
nor UO_3081 (O_3081,N_25449,N_26315);
nand UO_3082 (O_3082,N_28749,N_29049);
nor UO_3083 (O_3083,N_29882,N_25024);
or UO_3084 (O_3084,N_24052,N_27752);
or UO_3085 (O_3085,N_24656,N_26375);
and UO_3086 (O_3086,N_26305,N_27759);
and UO_3087 (O_3087,N_28945,N_29739);
and UO_3088 (O_3088,N_26210,N_27392);
nor UO_3089 (O_3089,N_29023,N_28013);
nor UO_3090 (O_3090,N_28959,N_28629);
and UO_3091 (O_3091,N_29775,N_26972);
nand UO_3092 (O_3092,N_25246,N_28985);
nor UO_3093 (O_3093,N_25594,N_26375);
nand UO_3094 (O_3094,N_29603,N_25084);
xor UO_3095 (O_3095,N_27554,N_27201);
nor UO_3096 (O_3096,N_27091,N_24687);
and UO_3097 (O_3097,N_28460,N_24068);
nor UO_3098 (O_3098,N_27263,N_28563);
nand UO_3099 (O_3099,N_24071,N_29509);
xnor UO_3100 (O_3100,N_24888,N_25025);
and UO_3101 (O_3101,N_24935,N_25058);
xor UO_3102 (O_3102,N_27315,N_26109);
nor UO_3103 (O_3103,N_24474,N_29780);
nor UO_3104 (O_3104,N_28142,N_29746);
xor UO_3105 (O_3105,N_27700,N_24734);
nand UO_3106 (O_3106,N_29392,N_24149);
xor UO_3107 (O_3107,N_27894,N_27113);
and UO_3108 (O_3108,N_29044,N_29829);
nand UO_3109 (O_3109,N_28801,N_28211);
or UO_3110 (O_3110,N_26296,N_24563);
nand UO_3111 (O_3111,N_26397,N_27686);
nand UO_3112 (O_3112,N_26435,N_25602);
nand UO_3113 (O_3113,N_28034,N_29456);
and UO_3114 (O_3114,N_25871,N_26619);
nand UO_3115 (O_3115,N_27034,N_29662);
nand UO_3116 (O_3116,N_25351,N_29741);
or UO_3117 (O_3117,N_25010,N_29620);
and UO_3118 (O_3118,N_24689,N_26646);
nor UO_3119 (O_3119,N_27436,N_29828);
xor UO_3120 (O_3120,N_26511,N_26645);
nor UO_3121 (O_3121,N_25041,N_24642);
nor UO_3122 (O_3122,N_25223,N_26834);
nor UO_3123 (O_3123,N_25609,N_28399);
xor UO_3124 (O_3124,N_27200,N_25743);
xnor UO_3125 (O_3125,N_27198,N_27243);
nor UO_3126 (O_3126,N_24021,N_26293);
nor UO_3127 (O_3127,N_25012,N_29897);
nor UO_3128 (O_3128,N_29060,N_28126);
nor UO_3129 (O_3129,N_25307,N_24746);
xor UO_3130 (O_3130,N_26636,N_24589);
xnor UO_3131 (O_3131,N_27181,N_26061);
and UO_3132 (O_3132,N_27463,N_24123);
xnor UO_3133 (O_3133,N_25787,N_28208);
or UO_3134 (O_3134,N_25734,N_27265);
or UO_3135 (O_3135,N_29983,N_25969);
and UO_3136 (O_3136,N_28815,N_24823);
and UO_3137 (O_3137,N_26769,N_28955);
and UO_3138 (O_3138,N_27994,N_28490);
xnor UO_3139 (O_3139,N_29945,N_29899);
and UO_3140 (O_3140,N_24574,N_25518);
nand UO_3141 (O_3141,N_27088,N_28496);
xnor UO_3142 (O_3142,N_24324,N_26399);
and UO_3143 (O_3143,N_25845,N_29962);
xor UO_3144 (O_3144,N_26782,N_25580);
nand UO_3145 (O_3145,N_25354,N_24023);
and UO_3146 (O_3146,N_29681,N_26159);
xor UO_3147 (O_3147,N_27121,N_27833);
nor UO_3148 (O_3148,N_26325,N_28467);
or UO_3149 (O_3149,N_25551,N_28595);
nor UO_3150 (O_3150,N_24960,N_25464);
nor UO_3151 (O_3151,N_24222,N_25387);
and UO_3152 (O_3152,N_27158,N_25510);
nor UO_3153 (O_3153,N_27975,N_25967);
and UO_3154 (O_3154,N_27789,N_27343);
nand UO_3155 (O_3155,N_27180,N_27300);
nand UO_3156 (O_3156,N_29806,N_27094);
or UO_3157 (O_3157,N_24668,N_27879);
or UO_3158 (O_3158,N_29721,N_27243);
nand UO_3159 (O_3159,N_28332,N_29662);
xnor UO_3160 (O_3160,N_28376,N_29531);
xor UO_3161 (O_3161,N_26730,N_29362);
nor UO_3162 (O_3162,N_27147,N_26417);
or UO_3163 (O_3163,N_24564,N_27372);
nor UO_3164 (O_3164,N_25723,N_28179);
nor UO_3165 (O_3165,N_29257,N_24402);
nand UO_3166 (O_3166,N_24712,N_24352);
nor UO_3167 (O_3167,N_27933,N_25595);
and UO_3168 (O_3168,N_28532,N_28129);
and UO_3169 (O_3169,N_26485,N_29235);
nor UO_3170 (O_3170,N_27836,N_24022);
and UO_3171 (O_3171,N_26919,N_26083);
and UO_3172 (O_3172,N_24906,N_29677);
or UO_3173 (O_3173,N_24511,N_28273);
or UO_3174 (O_3174,N_28002,N_27676);
or UO_3175 (O_3175,N_27694,N_26905);
or UO_3176 (O_3176,N_25523,N_26514);
nor UO_3177 (O_3177,N_24006,N_29954);
xor UO_3178 (O_3178,N_28523,N_25293);
and UO_3179 (O_3179,N_26065,N_24276);
nand UO_3180 (O_3180,N_27099,N_29927);
xor UO_3181 (O_3181,N_28454,N_25411);
or UO_3182 (O_3182,N_29794,N_24064);
nand UO_3183 (O_3183,N_25690,N_25873);
nor UO_3184 (O_3184,N_29687,N_29337);
nor UO_3185 (O_3185,N_27656,N_27534);
and UO_3186 (O_3186,N_28303,N_28513);
nor UO_3187 (O_3187,N_28963,N_29389);
xor UO_3188 (O_3188,N_25267,N_29939);
xnor UO_3189 (O_3189,N_29266,N_28302);
xor UO_3190 (O_3190,N_28284,N_26109);
nand UO_3191 (O_3191,N_27967,N_29952);
nor UO_3192 (O_3192,N_26832,N_27494);
nor UO_3193 (O_3193,N_26931,N_24339);
or UO_3194 (O_3194,N_28165,N_24537);
and UO_3195 (O_3195,N_29091,N_28984);
and UO_3196 (O_3196,N_25964,N_24079);
and UO_3197 (O_3197,N_24852,N_26835);
nor UO_3198 (O_3198,N_27668,N_25314);
and UO_3199 (O_3199,N_26792,N_26384);
or UO_3200 (O_3200,N_27822,N_25340);
nand UO_3201 (O_3201,N_27961,N_29023);
and UO_3202 (O_3202,N_24820,N_27853);
nand UO_3203 (O_3203,N_29939,N_25447);
nand UO_3204 (O_3204,N_26594,N_24405);
nand UO_3205 (O_3205,N_25419,N_24197);
nand UO_3206 (O_3206,N_26145,N_27481);
or UO_3207 (O_3207,N_28116,N_26788);
nor UO_3208 (O_3208,N_25553,N_27060);
and UO_3209 (O_3209,N_27053,N_25263);
nor UO_3210 (O_3210,N_26411,N_26908);
or UO_3211 (O_3211,N_24278,N_25407);
or UO_3212 (O_3212,N_26377,N_24987);
nor UO_3213 (O_3213,N_28424,N_25802);
nor UO_3214 (O_3214,N_26967,N_24841);
xor UO_3215 (O_3215,N_27710,N_28888);
or UO_3216 (O_3216,N_28947,N_24126);
nor UO_3217 (O_3217,N_29103,N_25377);
or UO_3218 (O_3218,N_27775,N_29923);
xnor UO_3219 (O_3219,N_26769,N_29605);
nand UO_3220 (O_3220,N_25913,N_24728);
or UO_3221 (O_3221,N_28254,N_28386);
nor UO_3222 (O_3222,N_25437,N_25850);
xnor UO_3223 (O_3223,N_24012,N_27759);
nand UO_3224 (O_3224,N_24090,N_26410);
xnor UO_3225 (O_3225,N_29230,N_29899);
nor UO_3226 (O_3226,N_24599,N_28044);
nand UO_3227 (O_3227,N_29091,N_29985);
xor UO_3228 (O_3228,N_29410,N_25098);
nand UO_3229 (O_3229,N_24053,N_26713);
and UO_3230 (O_3230,N_28174,N_26859);
nor UO_3231 (O_3231,N_26884,N_26679);
and UO_3232 (O_3232,N_27820,N_24912);
xor UO_3233 (O_3233,N_26038,N_25042);
nor UO_3234 (O_3234,N_25323,N_25427);
and UO_3235 (O_3235,N_27254,N_25713);
nor UO_3236 (O_3236,N_28272,N_29101);
xor UO_3237 (O_3237,N_28964,N_26894);
xor UO_3238 (O_3238,N_26306,N_25068);
nand UO_3239 (O_3239,N_28912,N_24480);
nor UO_3240 (O_3240,N_24650,N_28918);
xor UO_3241 (O_3241,N_26881,N_24513);
nand UO_3242 (O_3242,N_29711,N_28962);
nand UO_3243 (O_3243,N_29054,N_27560);
or UO_3244 (O_3244,N_26214,N_25179);
and UO_3245 (O_3245,N_27281,N_26786);
nor UO_3246 (O_3246,N_24010,N_24305);
nand UO_3247 (O_3247,N_27488,N_26705);
nor UO_3248 (O_3248,N_24393,N_26977);
and UO_3249 (O_3249,N_27617,N_24314);
nand UO_3250 (O_3250,N_25265,N_28022);
nand UO_3251 (O_3251,N_25703,N_26857);
xnor UO_3252 (O_3252,N_24228,N_26560);
xnor UO_3253 (O_3253,N_27620,N_25033);
nor UO_3254 (O_3254,N_29486,N_29391);
nor UO_3255 (O_3255,N_27032,N_25199);
xnor UO_3256 (O_3256,N_28090,N_29209);
and UO_3257 (O_3257,N_28092,N_26105);
xnor UO_3258 (O_3258,N_29856,N_29860);
nand UO_3259 (O_3259,N_27695,N_25868);
and UO_3260 (O_3260,N_26454,N_26378);
xnor UO_3261 (O_3261,N_25381,N_24139);
or UO_3262 (O_3262,N_29801,N_26849);
and UO_3263 (O_3263,N_27307,N_27953);
or UO_3264 (O_3264,N_29270,N_29698);
and UO_3265 (O_3265,N_26949,N_25982);
nor UO_3266 (O_3266,N_26589,N_24723);
or UO_3267 (O_3267,N_28745,N_26824);
nor UO_3268 (O_3268,N_26756,N_28795);
and UO_3269 (O_3269,N_27427,N_24326);
nor UO_3270 (O_3270,N_26876,N_29512);
xnor UO_3271 (O_3271,N_29147,N_24670);
nand UO_3272 (O_3272,N_28043,N_26125);
or UO_3273 (O_3273,N_28081,N_25468);
and UO_3274 (O_3274,N_27241,N_27160);
or UO_3275 (O_3275,N_26990,N_24471);
nand UO_3276 (O_3276,N_26400,N_26387);
or UO_3277 (O_3277,N_27285,N_27741);
or UO_3278 (O_3278,N_29576,N_27621);
or UO_3279 (O_3279,N_28824,N_29916);
or UO_3280 (O_3280,N_29232,N_29219);
and UO_3281 (O_3281,N_27288,N_28855);
nor UO_3282 (O_3282,N_28008,N_24810);
nor UO_3283 (O_3283,N_27585,N_24483);
xnor UO_3284 (O_3284,N_28951,N_29066);
and UO_3285 (O_3285,N_25055,N_26813);
nand UO_3286 (O_3286,N_29110,N_26174);
nand UO_3287 (O_3287,N_25460,N_27201);
nor UO_3288 (O_3288,N_26979,N_29041);
nand UO_3289 (O_3289,N_24423,N_24178);
nand UO_3290 (O_3290,N_25945,N_24896);
nand UO_3291 (O_3291,N_25232,N_25632);
nand UO_3292 (O_3292,N_29732,N_28852);
nand UO_3293 (O_3293,N_29736,N_28107);
xor UO_3294 (O_3294,N_29961,N_26433);
or UO_3295 (O_3295,N_28270,N_27367);
or UO_3296 (O_3296,N_29669,N_24798);
or UO_3297 (O_3297,N_29058,N_24036);
xor UO_3298 (O_3298,N_26302,N_28766);
nor UO_3299 (O_3299,N_26474,N_24908);
nor UO_3300 (O_3300,N_26841,N_26621);
or UO_3301 (O_3301,N_26308,N_25884);
or UO_3302 (O_3302,N_25827,N_24095);
and UO_3303 (O_3303,N_27318,N_27291);
and UO_3304 (O_3304,N_24190,N_25668);
xnor UO_3305 (O_3305,N_28670,N_25160);
nand UO_3306 (O_3306,N_27941,N_25255);
and UO_3307 (O_3307,N_24599,N_25080);
nand UO_3308 (O_3308,N_26169,N_27419);
nand UO_3309 (O_3309,N_24056,N_24578);
and UO_3310 (O_3310,N_25106,N_26390);
xor UO_3311 (O_3311,N_29603,N_24857);
nand UO_3312 (O_3312,N_29226,N_29639);
nor UO_3313 (O_3313,N_24410,N_27745);
nor UO_3314 (O_3314,N_28548,N_28708);
xor UO_3315 (O_3315,N_24145,N_29174);
nor UO_3316 (O_3316,N_27762,N_26115);
and UO_3317 (O_3317,N_28093,N_25234);
nor UO_3318 (O_3318,N_28143,N_28664);
and UO_3319 (O_3319,N_26498,N_27962);
nand UO_3320 (O_3320,N_24597,N_25434);
nor UO_3321 (O_3321,N_29798,N_28261);
nor UO_3322 (O_3322,N_29857,N_27714);
and UO_3323 (O_3323,N_29268,N_24370);
or UO_3324 (O_3324,N_24513,N_28118);
or UO_3325 (O_3325,N_26319,N_25806);
and UO_3326 (O_3326,N_27654,N_28180);
or UO_3327 (O_3327,N_25538,N_25407);
xor UO_3328 (O_3328,N_26438,N_28831);
and UO_3329 (O_3329,N_29006,N_26942);
xor UO_3330 (O_3330,N_27048,N_24824);
or UO_3331 (O_3331,N_26821,N_24784);
nor UO_3332 (O_3332,N_25745,N_28781);
nand UO_3333 (O_3333,N_24549,N_28375);
nor UO_3334 (O_3334,N_25715,N_26915);
and UO_3335 (O_3335,N_25954,N_25103);
nor UO_3336 (O_3336,N_26714,N_27876);
or UO_3337 (O_3337,N_27707,N_29825);
and UO_3338 (O_3338,N_26740,N_26277);
nor UO_3339 (O_3339,N_29470,N_28512);
xor UO_3340 (O_3340,N_29496,N_27055);
xor UO_3341 (O_3341,N_26663,N_28132);
and UO_3342 (O_3342,N_28090,N_24277);
or UO_3343 (O_3343,N_28694,N_24211);
nand UO_3344 (O_3344,N_24055,N_29051);
nand UO_3345 (O_3345,N_25771,N_29660);
nor UO_3346 (O_3346,N_28476,N_24737);
and UO_3347 (O_3347,N_24858,N_24617);
or UO_3348 (O_3348,N_26803,N_24036);
or UO_3349 (O_3349,N_24280,N_26881);
xnor UO_3350 (O_3350,N_27504,N_25078);
nand UO_3351 (O_3351,N_28895,N_27788);
nand UO_3352 (O_3352,N_28038,N_26279);
nand UO_3353 (O_3353,N_29254,N_26605);
xnor UO_3354 (O_3354,N_27522,N_28610);
xnor UO_3355 (O_3355,N_25267,N_25706);
and UO_3356 (O_3356,N_27643,N_24682);
xnor UO_3357 (O_3357,N_27855,N_27070);
nor UO_3358 (O_3358,N_24001,N_28256);
or UO_3359 (O_3359,N_27683,N_24746);
nor UO_3360 (O_3360,N_26254,N_26930);
or UO_3361 (O_3361,N_24377,N_29569);
nor UO_3362 (O_3362,N_26048,N_26457);
nand UO_3363 (O_3363,N_27016,N_24423);
or UO_3364 (O_3364,N_24923,N_26057);
and UO_3365 (O_3365,N_25086,N_25581);
xnor UO_3366 (O_3366,N_25744,N_25533);
nand UO_3367 (O_3367,N_24975,N_29481);
nand UO_3368 (O_3368,N_26241,N_26743);
nand UO_3369 (O_3369,N_25901,N_24258);
and UO_3370 (O_3370,N_24875,N_27184);
and UO_3371 (O_3371,N_27221,N_24861);
xnor UO_3372 (O_3372,N_27143,N_24795);
nor UO_3373 (O_3373,N_25921,N_28391);
nor UO_3374 (O_3374,N_24627,N_28346);
or UO_3375 (O_3375,N_28387,N_29075);
nand UO_3376 (O_3376,N_26571,N_27117);
nand UO_3377 (O_3377,N_26827,N_25703);
xor UO_3378 (O_3378,N_27598,N_27070);
and UO_3379 (O_3379,N_27868,N_25370);
xnor UO_3380 (O_3380,N_28831,N_24101);
and UO_3381 (O_3381,N_26023,N_28370);
xor UO_3382 (O_3382,N_25363,N_25506);
xor UO_3383 (O_3383,N_26866,N_29893);
xnor UO_3384 (O_3384,N_27022,N_28924);
nand UO_3385 (O_3385,N_24997,N_28010);
xnor UO_3386 (O_3386,N_26283,N_29012);
nand UO_3387 (O_3387,N_25175,N_29222);
or UO_3388 (O_3388,N_24542,N_24698);
nor UO_3389 (O_3389,N_27346,N_27367);
xor UO_3390 (O_3390,N_28251,N_29176);
nand UO_3391 (O_3391,N_27471,N_26942);
and UO_3392 (O_3392,N_29195,N_28968);
and UO_3393 (O_3393,N_25976,N_27622);
nor UO_3394 (O_3394,N_24631,N_24484);
xnor UO_3395 (O_3395,N_25310,N_28206);
nand UO_3396 (O_3396,N_29714,N_29327);
nor UO_3397 (O_3397,N_25115,N_29666);
nor UO_3398 (O_3398,N_24271,N_24066);
nand UO_3399 (O_3399,N_26716,N_28546);
xor UO_3400 (O_3400,N_25017,N_25863);
or UO_3401 (O_3401,N_29008,N_27898);
xor UO_3402 (O_3402,N_28554,N_27596);
nor UO_3403 (O_3403,N_28463,N_25930);
or UO_3404 (O_3404,N_27766,N_25494);
and UO_3405 (O_3405,N_29658,N_24647);
nand UO_3406 (O_3406,N_24647,N_26927);
and UO_3407 (O_3407,N_24824,N_24862);
and UO_3408 (O_3408,N_28792,N_26380);
and UO_3409 (O_3409,N_26447,N_28329);
nand UO_3410 (O_3410,N_27813,N_25988);
or UO_3411 (O_3411,N_24041,N_24412);
xor UO_3412 (O_3412,N_29563,N_27022);
or UO_3413 (O_3413,N_29409,N_28242);
nand UO_3414 (O_3414,N_26882,N_29855);
and UO_3415 (O_3415,N_28790,N_27234);
nand UO_3416 (O_3416,N_28753,N_28178);
xor UO_3417 (O_3417,N_28667,N_26687);
and UO_3418 (O_3418,N_27724,N_26029);
nand UO_3419 (O_3419,N_26522,N_27022);
nor UO_3420 (O_3420,N_24376,N_27189);
and UO_3421 (O_3421,N_25211,N_29065);
nor UO_3422 (O_3422,N_29831,N_29633);
or UO_3423 (O_3423,N_26178,N_24798);
nand UO_3424 (O_3424,N_26788,N_25102);
and UO_3425 (O_3425,N_26388,N_24953);
and UO_3426 (O_3426,N_25297,N_29423);
nand UO_3427 (O_3427,N_29670,N_26206);
and UO_3428 (O_3428,N_26093,N_25107);
xor UO_3429 (O_3429,N_27696,N_24048);
and UO_3430 (O_3430,N_27969,N_24751);
nand UO_3431 (O_3431,N_27697,N_28194);
and UO_3432 (O_3432,N_26295,N_26559);
nor UO_3433 (O_3433,N_24596,N_24704);
or UO_3434 (O_3434,N_25494,N_28355);
xnor UO_3435 (O_3435,N_25195,N_25958);
nand UO_3436 (O_3436,N_28420,N_24551);
xnor UO_3437 (O_3437,N_24555,N_29353);
xnor UO_3438 (O_3438,N_24040,N_27102);
or UO_3439 (O_3439,N_26467,N_28883);
or UO_3440 (O_3440,N_25086,N_26025);
xor UO_3441 (O_3441,N_25336,N_25943);
and UO_3442 (O_3442,N_24898,N_25116);
and UO_3443 (O_3443,N_28418,N_26017);
nor UO_3444 (O_3444,N_29708,N_24096);
and UO_3445 (O_3445,N_26105,N_28446);
nand UO_3446 (O_3446,N_26534,N_26589);
nand UO_3447 (O_3447,N_25345,N_27698);
or UO_3448 (O_3448,N_24463,N_28338);
xnor UO_3449 (O_3449,N_24357,N_26358);
and UO_3450 (O_3450,N_27223,N_27828);
nand UO_3451 (O_3451,N_28529,N_25361);
nor UO_3452 (O_3452,N_25381,N_29805);
xnor UO_3453 (O_3453,N_26189,N_27188);
nand UO_3454 (O_3454,N_28929,N_24720);
and UO_3455 (O_3455,N_25871,N_24431);
or UO_3456 (O_3456,N_29297,N_25234);
nand UO_3457 (O_3457,N_26950,N_27792);
nor UO_3458 (O_3458,N_29416,N_26271);
nor UO_3459 (O_3459,N_24751,N_25640);
nor UO_3460 (O_3460,N_25587,N_28460);
nor UO_3461 (O_3461,N_28951,N_24475);
nor UO_3462 (O_3462,N_27060,N_25056);
or UO_3463 (O_3463,N_29868,N_29397);
xnor UO_3464 (O_3464,N_25513,N_28557);
nor UO_3465 (O_3465,N_26778,N_24912);
nor UO_3466 (O_3466,N_25762,N_25509);
xnor UO_3467 (O_3467,N_28439,N_26535);
or UO_3468 (O_3468,N_27275,N_29921);
or UO_3469 (O_3469,N_28427,N_24424);
xnor UO_3470 (O_3470,N_24593,N_27300);
nor UO_3471 (O_3471,N_25976,N_28958);
nor UO_3472 (O_3472,N_29757,N_24111);
nor UO_3473 (O_3473,N_25195,N_26136);
nor UO_3474 (O_3474,N_25211,N_28029);
nand UO_3475 (O_3475,N_29654,N_26660);
or UO_3476 (O_3476,N_25892,N_24428);
nand UO_3477 (O_3477,N_27438,N_29471);
and UO_3478 (O_3478,N_29879,N_27134);
and UO_3479 (O_3479,N_29305,N_27046);
xnor UO_3480 (O_3480,N_26831,N_25427);
nand UO_3481 (O_3481,N_27222,N_27315);
nor UO_3482 (O_3482,N_26967,N_25961);
xnor UO_3483 (O_3483,N_24417,N_26164);
xor UO_3484 (O_3484,N_24718,N_24382);
and UO_3485 (O_3485,N_28132,N_25476);
nand UO_3486 (O_3486,N_28880,N_27622);
nand UO_3487 (O_3487,N_27458,N_27970);
nor UO_3488 (O_3488,N_27096,N_24591);
and UO_3489 (O_3489,N_24032,N_28018);
nand UO_3490 (O_3490,N_25095,N_24405);
or UO_3491 (O_3491,N_24678,N_28628);
and UO_3492 (O_3492,N_29410,N_28796);
nor UO_3493 (O_3493,N_25203,N_26462);
nor UO_3494 (O_3494,N_28953,N_27178);
or UO_3495 (O_3495,N_24800,N_29905);
xor UO_3496 (O_3496,N_27795,N_29463);
or UO_3497 (O_3497,N_28106,N_24644);
xor UO_3498 (O_3498,N_25744,N_27359);
nor UO_3499 (O_3499,N_26380,N_24092);
endmodule