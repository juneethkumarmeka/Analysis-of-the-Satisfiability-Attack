module basic_2000_20000_2500_10_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_175,In_1606);
or U1 (N_1,In_460,In_554);
nand U2 (N_2,In_867,In_1856);
nand U3 (N_3,In_1912,In_1181);
or U4 (N_4,In_1789,In_663);
or U5 (N_5,In_1418,In_794);
or U6 (N_6,In_1233,In_1027);
and U7 (N_7,In_1374,In_1538);
or U8 (N_8,In_917,In_1978);
nand U9 (N_9,In_1093,In_110);
nor U10 (N_10,In_1268,In_1331);
nand U11 (N_11,In_306,In_1623);
xor U12 (N_12,In_1929,In_774);
and U13 (N_13,In_1705,In_1953);
or U14 (N_14,In_499,In_401);
nor U15 (N_15,In_90,In_419);
or U16 (N_16,In_829,In_1216);
nor U17 (N_17,In_980,In_1753);
or U18 (N_18,In_479,In_1097);
nand U19 (N_19,In_1373,In_935);
xnor U20 (N_20,In_1486,In_1434);
and U21 (N_21,In_28,In_645);
and U22 (N_22,In_1478,In_654);
or U23 (N_23,In_797,In_924);
and U24 (N_24,In_1143,In_83);
nor U25 (N_25,In_1370,In_439);
nand U26 (N_26,In_108,In_1344);
nand U27 (N_27,In_1513,In_810);
or U28 (N_28,In_846,In_1082);
or U29 (N_29,In_74,In_805);
nand U30 (N_30,In_235,In_928);
and U31 (N_31,In_18,In_1278);
and U32 (N_32,In_435,In_1274);
and U33 (N_33,In_1426,In_82);
and U34 (N_34,In_1157,In_327);
and U35 (N_35,In_1456,In_1096);
xor U36 (N_36,In_1488,In_1160);
and U37 (N_37,In_377,In_1709);
nand U38 (N_38,In_1225,In_723);
xnor U39 (N_39,In_936,In_1925);
or U40 (N_40,In_1724,In_1182);
or U41 (N_41,In_800,In_397);
and U42 (N_42,In_107,In_537);
nor U43 (N_43,In_815,In_530);
nor U44 (N_44,In_940,In_325);
and U45 (N_45,In_691,In_265);
nand U46 (N_46,In_411,In_313);
and U47 (N_47,In_1603,In_1845);
xor U48 (N_48,In_332,In_448);
and U49 (N_49,In_553,In_260);
or U50 (N_50,In_261,In_453);
nand U51 (N_51,In_741,In_1654);
nor U52 (N_52,In_1868,In_1118);
and U53 (N_53,In_1894,In_1955);
and U54 (N_54,In_1698,In_727);
nor U55 (N_55,In_292,In_1435);
and U56 (N_56,In_1039,In_1008);
or U57 (N_57,In_34,In_1341);
or U58 (N_58,In_1794,In_358);
or U59 (N_59,In_444,In_476);
nor U60 (N_60,In_1253,In_1446);
xor U61 (N_61,In_1037,In_489);
nand U62 (N_62,In_1134,In_272);
and U63 (N_63,In_264,In_1360);
or U64 (N_64,In_1240,In_1916);
nand U65 (N_65,In_964,In_66);
and U66 (N_66,In_161,In_944);
nor U67 (N_67,In_467,In_801);
or U68 (N_68,In_369,In_1392);
or U69 (N_69,In_1757,In_1590);
or U70 (N_70,In_1232,In_355);
and U71 (N_71,In_290,In_667);
or U72 (N_72,In_1734,In_1895);
and U73 (N_73,In_985,In_1920);
xor U74 (N_74,In_1166,In_966);
xor U75 (N_75,In_360,In_1677);
nor U76 (N_76,In_1057,In_63);
nor U77 (N_77,In_1617,In_975);
nand U78 (N_78,In_1884,In_1474);
and U79 (N_79,In_1537,In_1439);
nor U80 (N_80,In_947,In_1797);
or U81 (N_81,In_482,In_968);
nand U82 (N_82,In_30,In_149);
nor U83 (N_83,In_621,In_1948);
nor U84 (N_84,In_67,In_1294);
or U85 (N_85,In_109,In_819);
and U86 (N_86,In_1365,In_481);
or U87 (N_87,In_714,In_211);
xor U88 (N_88,In_299,In_735);
nor U89 (N_89,In_638,In_248);
nand U90 (N_90,In_1583,In_27);
nor U91 (N_91,In_338,In_697);
nor U92 (N_92,In_1672,In_1577);
nand U93 (N_93,In_521,In_1259);
and U94 (N_94,In_147,In_1621);
nor U95 (N_95,In_1864,In_748);
or U96 (N_96,In_1979,In_1077);
or U97 (N_97,In_1988,In_1578);
nand U98 (N_98,In_1207,In_843);
and U99 (N_99,In_1256,In_642);
and U100 (N_100,In_1247,In_1930);
and U101 (N_101,In_1174,In_1443);
nand U102 (N_102,In_1178,In_600);
nor U103 (N_103,In_88,In_830);
nor U104 (N_104,In_738,In_71);
and U105 (N_105,In_523,In_1170);
and U106 (N_106,In_341,In_1980);
and U107 (N_107,In_1737,In_1349);
and U108 (N_108,In_1714,In_339);
nand U109 (N_109,In_808,In_171);
xor U110 (N_110,In_999,In_623);
xor U111 (N_111,In_422,In_212);
nor U112 (N_112,In_1249,In_1084);
or U113 (N_113,In_69,In_677);
or U114 (N_114,In_181,In_792);
nand U115 (N_115,In_1071,In_506);
or U116 (N_116,In_121,In_1716);
or U117 (N_117,In_1248,In_1465);
nor U118 (N_118,In_1112,In_170);
nand U119 (N_119,In_1176,In_1999);
and U120 (N_120,In_1356,In_1368);
or U121 (N_121,In_1956,In_758);
or U122 (N_122,In_43,In_1751);
nor U123 (N_123,In_685,In_312);
nor U124 (N_124,In_1552,In_73);
or U125 (N_125,In_694,In_647);
nand U126 (N_126,In_1943,In_1770);
and U127 (N_127,In_952,In_1154);
and U128 (N_128,In_1842,In_434);
xnor U129 (N_129,In_798,In_1711);
or U130 (N_130,In_122,In_719);
or U131 (N_131,In_1006,In_698);
or U132 (N_132,In_1932,In_1505);
or U133 (N_133,In_400,In_364);
nand U134 (N_134,In_681,In_726);
or U135 (N_135,In_1874,In_1620);
or U136 (N_136,In_957,In_1320);
or U137 (N_137,In_1908,In_737);
or U138 (N_138,In_441,In_1324);
xor U139 (N_139,In_1415,In_1347);
or U140 (N_140,In_456,In_713);
and U141 (N_141,In_1931,In_1832);
nand U142 (N_142,In_1109,In_1732);
nor U143 (N_143,In_383,In_1198);
nand U144 (N_144,In_670,In_240);
nor U145 (N_145,In_988,In_1735);
nor U146 (N_146,In_901,In_20);
and U147 (N_147,In_1188,In_1025);
nor U148 (N_148,In_1726,In_1860);
nand U149 (N_149,In_1602,In_1872);
and U150 (N_150,In_1830,In_1394);
or U151 (N_151,In_1179,In_138);
and U152 (N_152,In_615,In_1404);
and U153 (N_153,In_593,In_1481);
and U154 (N_154,In_430,In_1237);
nor U155 (N_155,In_1444,In_1030);
and U156 (N_156,In_836,In_1263);
xnor U157 (N_157,In_1959,In_569);
and U158 (N_158,In_49,In_330);
or U159 (N_159,In_1464,In_1799);
and U160 (N_160,In_446,In_1150);
nand U161 (N_161,In_1473,In_1622);
xnor U162 (N_162,In_1660,In_1846);
xnor U163 (N_163,In_180,In_958);
nor U164 (N_164,In_1448,In_1740);
nand U165 (N_165,In_1026,In_1075);
xor U166 (N_166,In_1345,In_854);
nor U167 (N_167,In_1954,In_1431);
nand U168 (N_168,In_1339,In_1055);
nor U169 (N_169,In_1241,In_372);
nand U170 (N_170,In_1318,In_1524);
xor U171 (N_171,In_1888,In_436);
and U172 (N_172,In_1200,In_1838);
and U173 (N_173,In_1681,In_596);
nor U174 (N_174,In_907,In_1739);
nand U175 (N_175,In_1982,In_911);
nand U176 (N_176,In_608,In_889);
and U177 (N_177,In_1246,In_1857);
and U178 (N_178,In_1610,In_268);
nand U179 (N_179,In_60,In_15);
nand U180 (N_180,In_1822,In_1397);
xor U181 (N_181,In_1784,In_918);
nand U182 (N_182,In_1229,In_1715);
or U183 (N_183,In_44,In_1796);
nand U184 (N_184,In_1546,In_1922);
or U185 (N_185,In_1967,In_906);
nand U186 (N_186,In_1924,In_1403);
nand U187 (N_187,In_1629,In_349);
xor U188 (N_188,In_320,In_862);
xor U189 (N_189,In_183,In_524);
and U190 (N_190,In_463,In_1183);
xor U191 (N_191,In_768,In_1512);
nor U192 (N_192,In_1708,In_1293);
nand U193 (N_193,In_1015,In_733);
nand U194 (N_194,In_731,In_547);
nor U195 (N_195,In_133,In_1094);
or U196 (N_196,In_579,In_827);
nor U197 (N_197,In_1767,In_494);
xor U198 (N_198,In_1467,In_1201);
or U199 (N_199,In_223,In_237);
nor U200 (N_200,In_1707,In_575);
nand U201 (N_201,In_1353,In_452);
nand U202 (N_202,In_1522,In_1171);
and U203 (N_203,In_1421,In_106);
or U204 (N_204,In_462,In_1139);
or U205 (N_205,In_5,In_413);
xor U206 (N_206,In_510,In_1079);
nor U207 (N_207,In_1539,In_722);
nand U208 (N_208,In_1848,In_578);
xor U209 (N_209,In_1001,In_1658);
xor U210 (N_210,In_514,In_1054);
or U211 (N_211,In_1102,In_1640);
or U212 (N_212,In_1744,In_1202);
and U213 (N_213,In_931,In_1591);
or U214 (N_214,In_747,In_669);
nand U215 (N_215,In_1409,In_1161);
nor U216 (N_216,In_1477,In_409);
and U217 (N_217,In_939,In_821);
xor U218 (N_218,In_915,In_1580);
and U219 (N_219,In_1485,In_594);
nor U220 (N_220,In_314,In_197);
nand U221 (N_221,In_130,In_495);
nor U222 (N_222,In_150,In_566);
xor U223 (N_223,In_89,In_1779);
and U224 (N_224,In_899,In_1438);
nand U225 (N_225,In_1910,In_883);
and U226 (N_226,In_0,In_62);
nand U227 (N_227,In_631,In_475);
nand U228 (N_228,In_459,In_1400);
and U229 (N_229,In_449,In_930);
nand U230 (N_230,In_1264,In_291);
and U231 (N_231,In_201,In_619);
and U232 (N_232,In_1503,In_1164);
or U233 (N_233,In_1490,In_913);
nand U234 (N_234,In_824,In_1386);
nand U235 (N_235,In_425,In_266);
nor U236 (N_236,In_1604,In_1046);
nand U237 (N_237,In_336,In_1049);
or U238 (N_238,In_131,In_371);
nand U239 (N_239,In_111,In_1065);
xor U240 (N_240,In_280,In_1628);
and U241 (N_241,In_1657,In_94);
and U242 (N_242,In_259,In_1103);
xor U243 (N_243,In_1540,In_156);
nor U244 (N_244,In_263,In_421);
nor U245 (N_245,In_246,In_1803);
and U246 (N_246,In_873,In_618);
or U247 (N_247,In_1892,In_159);
and U248 (N_248,In_923,In_763);
nor U249 (N_249,In_14,In_736);
or U250 (N_250,In_644,In_662);
nand U251 (N_251,In_1091,In_1131);
nand U252 (N_252,In_1398,In_381);
nor U253 (N_253,In_1428,In_390);
xor U254 (N_254,In_994,In_1371);
nor U255 (N_255,In_1226,In_388);
nor U256 (N_256,In_806,In_26);
nand U257 (N_257,In_1303,In_1376);
nand U258 (N_258,In_978,In_1720);
or U259 (N_259,In_269,In_176);
and U260 (N_260,In_1661,In_309);
and U261 (N_261,In_675,In_695);
xnor U262 (N_262,In_294,In_610);
and U263 (N_263,In_1937,In_1936);
nor U264 (N_264,In_983,In_1375);
nand U265 (N_265,In_611,In_565);
nand U266 (N_266,In_428,In_1491);
nor U267 (N_267,In_205,In_1136);
nor U268 (N_268,In_1587,In_1034);
and U269 (N_269,In_1257,In_1977);
and U270 (N_270,In_1024,In_404);
and U271 (N_271,In_218,In_210);
nand U272 (N_272,In_1985,In_1909);
or U273 (N_273,In_650,In_859);
nand U274 (N_274,In_16,In_828);
or U275 (N_275,In_1964,In_1701);
nand U276 (N_276,In_1120,In_1033);
or U277 (N_277,In_1457,In_1719);
nand U278 (N_278,In_787,In_1752);
nor U279 (N_279,In_188,In_1607);
xor U280 (N_280,In_1142,In_1975);
and U281 (N_281,In_1489,In_1108);
nor U282 (N_282,In_1949,In_981);
nor U283 (N_283,In_1668,In_822);
or U284 (N_284,In_1795,In_105);
nor U285 (N_285,In_1815,In_1514);
and U286 (N_286,In_541,In_771);
or U287 (N_287,In_1544,In_454);
or U288 (N_288,In_973,In_1563);
and U289 (N_289,In_139,In_1642);
nand U290 (N_290,In_1588,In_832);
and U291 (N_291,In_574,In_21);
nor U292 (N_292,In_729,In_960);
or U293 (N_293,In_394,In_535);
nand U294 (N_294,In_1307,In_443);
or U295 (N_295,In_1871,In_203);
and U296 (N_296,In_13,In_245);
or U297 (N_297,In_279,In_674);
and U298 (N_298,In_696,In_1593);
and U299 (N_299,In_1921,In_1687);
nand U300 (N_300,In_37,In_1335);
or U301 (N_301,In_1825,In_607);
and U302 (N_302,In_1463,In_693);
nand U303 (N_303,In_1683,In_79);
and U304 (N_304,In_1191,In_1265);
nor U305 (N_305,In_816,In_890);
and U306 (N_306,In_934,In_469);
and U307 (N_307,In_1840,In_1942);
xor U308 (N_308,In_289,In_1205);
and U309 (N_309,In_1568,In_359);
nor U310 (N_310,In_564,In_581);
and U311 (N_311,In_1211,In_704);
xor U312 (N_312,In_234,In_52);
nor U313 (N_313,In_1765,In_1381);
nand U314 (N_314,In_1405,In_1482);
nor U315 (N_315,In_293,In_335);
nor U316 (N_316,In_204,In_1940);
and U317 (N_317,In_1786,In_1685);
and U318 (N_318,In_1454,In_1697);
or U319 (N_319,In_1935,In_1252);
xor U320 (N_320,In_864,In_126);
nand U321 (N_321,In_1238,In_1251);
nand U322 (N_322,In_1035,In_301);
or U323 (N_323,In_1863,In_1385);
nand U324 (N_324,In_1957,In_1882);
and U325 (N_325,In_368,In_1509);
nand U326 (N_326,In_785,In_1560);
nor U327 (N_327,In_1245,In_119);
or U328 (N_328,In_707,In_1173);
nor U329 (N_329,In_55,In_1816);
and U330 (N_330,In_438,In_949);
nand U331 (N_331,In_884,In_331);
or U332 (N_332,In_1083,In_365);
nor U333 (N_333,In_1993,In_324);
xor U334 (N_334,In_1343,In_746);
xnor U335 (N_335,In_273,In_516);
nand U336 (N_336,In_875,In_1749);
and U337 (N_337,In_124,In_1432);
and U338 (N_338,In_376,In_847);
xor U339 (N_339,In_429,In_1287);
and U340 (N_340,In_625,In_1138);
and U341 (N_341,In_1571,In_1380);
nor U342 (N_342,In_128,In_1011);
and U343 (N_343,In_190,In_597);
or U344 (N_344,In_1938,In_1776);
xnor U345 (N_345,In_970,In_1674);
nor U346 (N_346,In_1301,In_1228);
and U347 (N_347,In_1833,In_252);
xnor U348 (N_348,In_1986,In_1133);
nor U349 (N_349,In_1748,In_1213);
or U350 (N_350,In_366,In_213);
nand U351 (N_351,In_1123,In_1762);
nor U352 (N_352,In_1831,In_297);
nor U353 (N_353,In_542,In_1926);
or U354 (N_354,In_1204,In_1122);
xnor U355 (N_355,In_195,In_1219);
nor U356 (N_356,In_328,In_657);
and U357 (N_357,In_174,In_592);
and U358 (N_358,In_851,In_503);
nand U359 (N_359,In_989,In_1731);
nand U360 (N_360,In_752,In_1021);
or U361 (N_361,In_1364,In_959);
and U362 (N_362,In_315,In_809);
and U363 (N_363,In_57,In_1016);
and U364 (N_364,In_790,In_560);
xor U365 (N_365,In_703,In_1627);
or U366 (N_366,In_215,In_648);
nand U367 (N_367,In_1558,In_1260);
nor U368 (N_368,In_1041,In_1718);
nand U369 (N_369,In_1665,In_567);
nor U370 (N_370,In_393,In_896);
or U371 (N_371,In_765,In_634);
nor U372 (N_372,In_730,In_1377);
or U373 (N_373,In_1609,In_874);
nor U374 (N_374,In_23,In_1745);
nor U375 (N_375,In_1086,In_281);
xnor U376 (N_376,In_1197,In_87);
or U377 (N_377,In_151,In_1644);
and U378 (N_378,In_761,In_326);
xor U379 (N_379,In_1323,In_1236);
xnor U380 (N_380,In_1650,In_700);
and U381 (N_381,In_220,In_185);
or U382 (N_382,In_1144,In_1453);
nor U383 (N_383,In_347,In_1458);
or U384 (N_384,In_38,In_137);
and U385 (N_385,In_876,In_1515);
and U386 (N_386,In_711,In_440);
or U387 (N_387,In_323,In_114);
or U388 (N_388,In_1111,In_750);
nor U389 (N_389,In_1327,In_1827);
nor U390 (N_390,In_559,In_1747);
xnor U391 (N_391,In_1866,In_1530);
or U392 (N_392,In_1313,In_627);
nor U393 (N_393,In_1682,In_891);
nor U394 (N_394,In_1028,In_298);
and U395 (N_395,In_416,In_1305);
or U396 (N_396,In_937,In_1430);
nor U397 (N_397,In_382,In_1785);
nor U398 (N_398,In_497,In_1449);
nand U399 (N_399,In_392,In_872);
nand U400 (N_400,In_1413,In_1774);
nand U401 (N_401,In_1483,In_1793);
and U402 (N_402,In_1152,In_1061);
and U403 (N_403,In_1511,In_1963);
and U404 (N_404,In_656,In_835);
or U405 (N_405,In_1877,In_1382);
nand U406 (N_406,In_739,In_403);
nor U407 (N_407,In_905,In_1276);
nand U408 (N_408,In_51,In_417);
nand U409 (N_409,In_540,In_660);
nand U410 (N_410,In_189,In_1780);
or U411 (N_411,In_1212,In_941);
nand U412 (N_412,In_1390,In_48);
xnor U413 (N_413,In_1754,In_1129);
and U414 (N_414,In_1873,In_1332);
or U415 (N_415,In_1728,In_1067);
nand U416 (N_416,In_491,In_1532);
or U417 (N_417,In_665,In_141);
or U418 (N_418,In_433,In_904);
nor U419 (N_419,In_1997,In_97);
nor U420 (N_420,In_643,In_337);
and U421 (N_421,In_1834,In_1192);
nand U422 (N_422,In_3,In_1471);
xnor U423 (N_423,In_39,In_142);
nor U424 (N_424,In_892,In_536);
nor U425 (N_425,In_1040,In_840);
nand U426 (N_426,In_1973,In_1630);
xnor U427 (N_427,In_591,In_1239);
xor U428 (N_428,In_1529,In_839);
and U429 (N_429,In_1535,In_64);
nand U430 (N_430,In_184,In_1378);
xor U431 (N_431,In_1414,In_29);
and U432 (N_432,In_1808,In_85);
nand U433 (N_433,In_1566,In_1080);
and U434 (N_434,In_384,In_1525);
nand U435 (N_435,In_1574,In_1594);
or U436 (N_436,In_1941,In_351);
and U437 (N_437,In_148,In_375);
and U438 (N_438,In_1905,In_65);
and U439 (N_439,In_274,In_35);
and U440 (N_440,In_480,In_96);
nor U441 (N_441,In_858,In_1423);
nor U442 (N_442,In_1777,In_1536);
nand U443 (N_443,In_12,In_818);
nor U444 (N_444,In_115,In_1099);
nor U445 (N_445,In_1311,In_1440);
xnor U446 (N_446,In_120,In_533);
xnor U447 (N_447,In_1140,In_997);
and U448 (N_448,In_676,In_1792);
nor U449 (N_449,In_455,In_308);
xnor U450 (N_450,In_1688,In_244);
nand U451 (N_451,In_1673,In_1304);
nor U452 (N_452,In_426,In_1826);
xnor U453 (N_453,In_1852,In_528);
nand U454 (N_454,In_943,In_1266);
and U455 (N_455,In_1402,In_740);
or U456 (N_456,In_1694,In_606);
or U457 (N_457,In_1424,In_814);
nor U458 (N_458,In_1723,In_1292);
or U459 (N_459,In_1007,In_1078);
nor U460 (N_460,In_1710,In_912);
nand U461 (N_461,In_902,In_1670);
nand U462 (N_462,In_1406,In_143);
or U463 (N_463,In_92,In_1072);
nor U464 (N_464,In_666,In_1820);
and U465 (N_465,In_307,In_1717);
or U466 (N_466,In_515,In_962);
nand U467 (N_467,In_1998,In_932);
and U468 (N_468,In_486,In_1053);
nor U469 (N_469,In_998,In_701);
nor U470 (N_470,In_1124,In_1811);
nand U471 (N_471,In_910,In_1234);
or U472 (N_472,In_492,In_938);
or U473 (N_473,In_98,In_751);
or U474 (N_474,In_471,In_1556);
xnor U475 (N_475,In_9,In_1523);
nand U476 (N_476,In_1756,In_1651);
nor U477 (N_477,In_196,In_76);
nand U478 (N_478,In_1554,In_1060);
or U479 (N_479,In_193,In_1755);
nand U480 (N_480,In_1655,In_1639);
xor U481 (N_481,In_1175,In_1965);
nand U482 (N_482,In_1854,In_1653);
or U483 (N_483,In_40,In_1961);
or U484 (N_484,In_101,In_47);
xnor U485 (N_485,In_451,In_1012);
nand U486 (N_486,In_352,In_1638);
and U487 (N_487,In_198,In_1357);
nand U488 (N_488,In_1498,In_1847);
xor U489 (N_489,In_1151,In_1417);
nand U490 (N_490,In_343,In_1476);
or U491 (N_491,In_278,In_179);
nor U492 (N_492,In_1081,In_688);
or U493 (N_493,In_1441,In_1379);
nand U494 (N_494,In_483,In_760);
and U495 (N_495,In_1363,In_1584);
nor U496 (N_496,In_861,In_1667);
nand U497 (N_497,In_1972,In_764);
or U498 (N_498,In_852,In_1288);
nor U499 (N_499,In_1231,In_288);
nor U500 (N_500,In_230,In_1813);
and U501 (N_501,In_56,In_1906);
nor U502 (N_502,In_1581,In_1611);
and U503 (N_503,In_206,In_1194);
or U504 (N_504,In_317,In_795);
or U505 (N_505,In_191,In_632);
nand U506 (N_506,In_1547,In_420);
xnor U507 (N_507,In_1104,In_734);
or U508 (N_508,In_464,In_1887);
nor U509 (N_509,In_1009,In_692);
or U510 (N_510,In_1098,In_186);
nor U511 (N_511,In_1684,In_1277);
nor U512 (N_512,In_802,In_1678);
or U513 (N_513,In_1952,In_945);
nand U514 (N_514,In_1968,In_1891);
and U515 (N_515,In_437,In_1597);
xor U516 (N_516,In_1399,In_1898);
nor U517 (N_517,In_921,In_466);
nand U518 (N_518,In_661,In_283);
nor U519 (N_519,In_1676,In_605);
and U520 (N_520,In_755,In_834);
and U521 (N_521,In_984,In_672);
or U522 (N_522,In_548,In_791);
nor U523 (N_523,In_1896,In_991);
or U524 (N_524,In_1828,In_72);
or U525 (N_525,In_226,In_427);
nor U526 (N_526,In_1562,In_617);
nor U527 (N_527,In_342,In_1470);
xor U528 (N_528,In_1422,In_1976);
nor U529 (N_529,In_742,In_1989);
nand U530 (N_530,In_1823,In_951);
nor U531 (N_531,In_744,In_146);
nor U532 (N_532,In_1817,In_219);
nand U533 (N_533,In_1244,In_1411);
nand U534 (N_534,In_1121,In_1169);
nand U535 (N_535,In_1088,In_1059);
nand U536 (N_536,In_70,In_982);
nand U537 (N_537,In_1325,In_1495);
nand U538 (N_538,In_1911,In_46);
or U539 (N_539,In_1763,In_511);
nand U540 (N_540,In_1531,In_1996);
and U541 (N_541,In_671,In_1613);
or U542 (N_542,In_1032,In_690);
and U543 (N_543,In_473,In_1902);
xor U544 (N_544,In_1814,In_1172);
nand U545 (N_545,In_262,In_652);
nor U546 (N_546,In_908,In_1336);
and U547 (N_547,In_1328,In_284);
and U548 (N_548,In_1506,In_950);
nand U549 (N_549,In_702,In_1275);
or U550 (N_550,In_517,In_898);
and U551 (N_551,In_1865,In_1487);
nor U552 (N_552,In_1396,In_1113);
or U553 (N_553,In_1044,In_418);
and U554 (N_554,In_682,In_100);
nor U555 (N_555,In_1507,In_1878);
nor U556 (N_556,In_1358,In_6);
nand U557 (N_557,In_588,In_1600);
or U558 (N_558,In_465,In_1217);
and U559 (N_559,In_842,In_504);
nand U560 (N_560,In_231,In_1383);
nor U561 (N_561,In_318,In_534);
nand U562 (N_562,In_1451,In_362);
nand U563 (N_563,In_25,In_1419);
or U564 (N_564,In_1798,In_1915);
and U565 (N_565,In_1608,In_487);
or U566 (N_566,In_833,In_1196);
nor U567 (N_567,In_214,In_136);
and U568 (N_568,In_1105,In_1612);
or U569 (N_569,In_1647,In_974);
nand U570 (N_570,In_1971,In_1599);
nand U571 (N_571,In_551,In_1527);
and U572 (N_572,In_1659,In_803);
or U573 (N_573,In_963,In_1369);
nor U574 (N_574,In_1761,In_1810);
xor U575 (N_575,In_820,In_1372);
nor U576 (N_576,In_779,In_493);
nor U577 (N_577,In_1010,In_1759);
and U578 (N_578,In_961,In_500);
nor U579 (N_579,In_1555,In_470);
nand U580 (N_580,In_340,In_972);
xor U581 (N_581,In_601,In_68);
or U582 (N_582,In_54,In_1062);
and U583 (N_583,In_775,In_1455);
nor U584 (N_584,In_778,In_2);
nor U585 (N_585,In_572,In_93);
or U586 (N_586,In_258,In_1992);
and U587 (N_587,In_1666,In_1867);
nor U588 (N_588,In_1843,In_42);
and U589 (N_589,In_965,In_1427);
and U590 (N_590,In_659,In_1412);
xnor U591 (N_591,In_1893,In_1788);
or U592 (N_592,In_956,In_1291);
nor U593 (N_593,In_885,In_1821);
nand U594 (N_594,In_33,In_1582);
nor U595 (N_595,In_562,In_257);
nor U596 (N_596,In_1945,In_424);
nor U597 (N_597,In_50,In_539);
nand U598 (N_598,In_1177,In_796);
or U599 (N_599,In_887,In_41);
or U600 (N_600,In_776,In_316);
and U601 (N_601,In_1675,In_1573);
and U602 (N_602,In_1760,In_152);
and U603 (N_603,In_1004,In_1351);
or U604 (N_604,In_1819,In_1746);
nor U605 (N_605,In_1452,In_1900);
and U606 (N_606,In_894,In_633);
nand U607 (N_607,In_720,In_10);
or U608 (N_608,In_1156,In_837);
nand U609 (N_609,In_302,In_485);
nand U610 (N_610,In_850,In_1758);
nand U611 (N_611,In_1733,In_1983);
xor U612 (N_612,In_254,In_450);
and U613 (N_613,In_1849,In_1624);
or U614 (N_614,In_386,In_583);
or U615 (N_615,In_160,In_7);
xor U616 (N_616,In_1570,In_1002);
and U617 (N_617,In_224,In_116);
and U618 (N_618,In_1844,In_8);
nand U619 (N_619,In_300,In_844);
or U620 (N_620,In_285,In_1258);
nor U621 (N_621,In_1870,In_955);
nor U622 (N_622,In_389,In_484);
nand U623 (N_623,In_1618,In_754);
and U624 (N_624,In_1729,In_1914);
nand U625 (N_625,In_1074,In_1869);
and U626 (N_626,In_1185,In_1391);
nor U627 (N_627,In_1020,In_172);
nor U628 (N_628,In_1790,In_1579);
nand U629 (N_629,In_1876,In_367);
nand U630 (N_630,In_1768,In_415);
or U631 (N_631,In_1807,In_769);
or U632 (N_632,In_1663,In_1850);
and U633 (N_633,In_895,In_927);
nand U634 (N_634,In_1189,In_721);
nand U635 (N_635,In_1520,In_1981);
nor U636 (N_636,In_1596,In_103);
xnor U637 (N_637,In_1899,In_577);
nand U638 (N_638,In_1279,In_1484);
or U639 (N_639,In_361,In_882);
or U640 (N_640,In_766,In_1730);
nor U641 (N_641,In_1771,In_102);
and U642 (N_642,In_571,In_710);
nand U643 (N_643,In_871,In_333);
xor U644 (N_644,In_334,In_613);
nand U645 (N_645,In_1713,In_1367);
nand U646 (N_646,In_1585,In_877);
nand U647 (N_647,In_900,In_1861);
and U648 (N_648,In_1282,In_641);
xor U649 (N_649,In_1296,In_1115);
xnor U650 (N_650,In_112,In_979);
or U651 (N_651,In_513,In_1003);
and U652 (N_652,In_78,In_1393);
and U653 (N_653,In_986,In_757);
xnor U654 (N_654,In_1146,In_310);
or U655 (N_655,In_1128,In_612);
nand U656 (N_656,In_1502,In_1806);
nor U657 (N_657,In_1669,In_992);
nor U658 (N_658,In_236,In_1526);
nand U659 (N_659,In_77,In_1076);
nand U660 (N_660,In_354,In_1564);
nor U661 (N_661,In_158,In_200);
nor U662 (N_662,In_1395,In_1114);
and U663 (N_663,In_75,In_1939);
and U664 (N_664,In_295,In_749);
nand U665 (N_665,In_544,In_1167);
and U666 (N_666,In_1286,In_45);
xor U667 (N_667,In_1800,In_1933);
and U668 (N_668,In_182,In_127);
nor U669 (N_669,In_1671,In_1703);
nand U670 (N_670,In_1772,In_501);
nor U671 (N_671,In_1553,In_831);
nand U672 (N_672,In_1429,In_1261);
nand U673 (N_673,In_36,In_391);
nor U674 (N_674,In_651,In_270);
xnor U675 (N_675,In_395,In_1220);
xor U676 (N_676,In_305,In_789);
or U677 (N_677,In_1496,In_1309);
nand U678 (N_678,In_845,In_1342);
xnor U679 (N_679,In_946,In_1326);
nor U680 (N_680,In_1333,In_1447);
nor U681 (N_681,In_773,In_276);
nor U682 (N_682,In_1664,In_538);
xnor U683 (N_683,In_468,In_1500);
nor U684 (N_684,In_1637,In_1433);
or U685 (N_685,In_1782,In_1903);
nor U686 (N_686,In_1619,In_95);
and U687 (N_687,In_1662,In_1149);
nand U688 (N_688,In_1727,In_217);
nor U689 (N_689,In_919,In_1235);
nand U690 (N_690,In_1545,In_1107);
or U691 (N_691,In_399,In_732);
nand U692 (N_692,In_255,In_1712);
or U693 (N_693,In_1387,In_568);
and U694 (N_694,In_1883,In_251);
nand U695 (N_695,In_849,In_1300);
nor U696 (N_696,In_1519,In_256);
nand U697 (N_697,In_1425,In_1853);
and U698 (N_698,In_953,In_1919);
and U699 (N_699,In_1,In_1802);
nor U700 (N_700,In_640,In_683);
or U701 (N_701,In_1410,In_474);
and U702 (N_702,In_1885,In_817);
xnor U703 (N_703,In_712,In_780);
or U704 (N_704,In_512,In_777);
xnor U705 (N_705,In_1738,In_1330);
nor U706 (N_706,In_228,In_1601);
or U707 (N_707,In_609,In_545);
nand U708 (N_708,In_1289,In_1295);
or U709 (N_709,In_1889,In_679);
or U710 (N_710,In_582,In_135);
and U711 (N_711,In_772,In_799);
nand U712 (N_712,In_1442,In_782);
nor U713 (N_713,In_848,In_1090);
and U714 (N_714,In_1262,In_1270);
and U715 (N_715,In_1841,In_1126);
or U716 (N_716,In_668,In_1479);
or U717 (N_717,In_445,In_1407);
or U718 (N_718,In_216,In_942);
nand U719 (N_719,In_1565,In_167);
and U720 (N_720,In_922,In_811);
nand U721 (N_721,In_550,In_1047);
and U722 (N_722,In_520,In_527);
and U723 (N_723,In_1700,In_1466);
and U724 (N_724,In_1722,In_125);
or U725 (N_725,In_346,In_1472);
nand U726 (N_726,In_1984,In_1310);
or U727 (N_727,In_706,In_353);
nand U728 (N_728,In_1605,In_1018);
and U729 (N_729,In_1636,In_1742);
and U730 (N_730,In_1280,In_1631);
nand U731 (N_731,In_250,In_1064);
xor U732 (N_732,In_178,In_1812);
and U733 (N_733,In_1764,In_1492);
nor U734 (N_734,In_1595,In_595);
nor U735 (N_735,In_118,In_1706);
xnor U736 (N_736,In_1508,In_1316);
nand U737 (N_737,In_1306,In_1193);
nor U738 (N_738,In_1679,In_177);
nand U739 (N_739,In_164,In_457);
nor U740 (N_740,In_1050,In_865);
xor U741 (N_741,In_1743,In_1804);
or U742 (N_742,In_1218,In_868);
nor U743 (N_743,In_1721,In_1469);
nor U744 (N_744,In_1119,In_916);
nor U745 (N_745,In_1214,In_1652);
xor U746 (N_746,In_199,In_909);
nor U747 (N_747,In_653,In_1561);
and U748 (N_748,In_1881,In_432);
nand U749 (N_749,In_1960,In_1056);
nor U750 (N_750,In_914,In_1901);
and U751 (N_751,In_1934,In_678);
nor U752 (N_752,In_1135,In_1958);
and U753 (N_753,In_61,In_396);
nand U754 (N_754,In_1572,In_1184);
nand U755 (N_755,In_573,In_717);
nand U756 (N_756,In_1928,In_1215);
nand U757 (N_757,In_823,In_209);
nand U758 (N_758,In_684,In_969);
and U759 (N_759,In_1648,In_556);
nor U760 (N_760,In_1633,In_507);
nor U761 (N_761,In_113,In_267);
xor U762 (N_762,In_329,In_1209);
nor U763 (N_763,In_350,In_207);
nor U764 (N_764,In_1051,In_1907);
nor U765 (N_765,In_1987,In_59);
nand U766 (N_766,In_933,In_1990);
nand U767 (N_767,In_555,In_977);
or U768 (N_768,In_546,In_812);
nor U769 (N_769,In_1693,In_1829);
xor U770 (N_770,In_458,In_275);
or U771 (N_771,In_1408,In_153);
xor U772 (N_772,In_1087,In_1147);
nor U773 (N_773,In_380,In_402);
or U774 (N_774,In_1242,In_53);
nor U775 (N_775,In_410,In_866);
and U776 (N_776,In_461,In_664);
or U777 (N_777,In_1361,In_1089);
nor U778 (N_778,In_1950,In_344);
xor U779 (N_779,In_373,In_1634);
nand U780 (N_780,In_1329,In_166);
nand U781 (N_781,In_1317,In_756);
or U782 (N_782,In_1890,In_549);
nor U783 (N_783,In_271,In_1125);
and U784 (N_784,In_637,In_165);
nor U785 (N_785,In_442,In_1013);
nor U786 (N_786,In_519,In_1947);
xor U787 (N_787,In_1528,In_1116);
nor U788 (N_788,In_1766,In_1995);
nor U789 (N_789,In_1148,In_287);
nor U790 (N_790,In_1879,In_17);
or U791 (N_791,In_781,In_759);
xor U792 (N_792,In_604,In_1913);
nand U793 (N_793,In_971,In_117);
nor U794 (N_794,In_1516,In_1346);
or U795 (N_795,In_1168,In_526);
nor U796 (N_796,In_1643,In_1559);
or U797 (N_797,In_241,In_995);
nor U798 (N_798,In_192,In_926);
xor U799 (N_799,In_1255,In_238);
and U800 (N_800,In_1736,In_522);
or U801 (N_801,In_86,In_705);
xnor U802 (N_802,In_1388,In_163);
or U803 (N_803,In_1557,In_84);
nand U804 (N_804,In_242,In_232);
nand U805 (N_805,In_239,In_247);
and U806 (N_806,In_1224,In_1206);
or U807 (N_807,In_1696,In_1319);
nor U808 (N_808,In_1321,In_976);
and U809 (N_809,In_1510,In_762);
or U810 (N_810,In_1969,In_624);
or U811 (N_811,In_1946,In_628);
nor U812 (N_812,In_1966,In_1615);
nor U813 (N_813,In_169,In_363);
nand U814 (N_814,In_880,In_414);
or U815 (N_815,In_1645,In_406);
nor U816 (N_816,In_658,In_1073);
or U817 (N_817,In_1101,In_1117);
nor U818 (N_818,In_715,In_1692);
and U819 (N_819,In_1686,In_897);
nand U820 (N_820,In_1058,In_1534);
and U821 (N_821,In_1835,In_888);
nor U822 (N_822,In_1680,In_1155);
nand U823 (N_823,In_1775,In_743);
or U824 (N_824,In_303,In_1501);
and U825 (N_825,In_1302,In_1781);
nor U826 (N_826,In_243,In_387);
nand U827 (N_827,In_636,In_655);
and U828 (N_828,In_1384,In_1927);
or U829 (N_829,In_1420,In_1180);
xor U830 (N_830,In_1106,In_531);
and U831 (N_831,In_1052,In_1163);
or U832 (N_832,In_1699,In_1145);
and U833 (N_833,In_570,In_1267);
or U834 (N_834,In_886,In_1352);
and U835 (N_835,In_1141,In_1043);
nor U836 (N_836,In_286,In_1023);
or U837 (N_837,In_1656,In_753);
or U838 (N_838,In_1250,In_1066);
and U839 (N_839,In_145,In_1285);
or U840 (N_840,In_929,In_561);
nand U841 (N_841,In_857,In_1308);
and U842 (N_842,In_1576,In_584);
xnor U843 (N_843,In_826,In_1551);
and U844 (N_844,In_32,In_1019);
nor U845 (N_845,In_1991,In_1695);
or U846 (N_846,In_379,In_580);
or U847 (N_847,In_304,In_1271);
and U848 (N_848,In_1354,In_1962);
nand U849 (N_849,In_140,In_1063);
nor U850 (N_850,In_155,In_1322);
or U851 (N_851,In_1070,In_793);
nor U852 (N_852,In_954,In_680);
nor U853 (N_853,In_408,In_173);
nor U854 (N_854,In_1416,In_1085);
or U855 (N_855,In_1031,In_1017);
and U856 (N_856,In_639,In_1635);
xnor U857 (N_857,In_249,In_144);
xor U858 (N_858,In_1436,In_370);
or U859 (N_859,In_1014,In_687);
nand U860 (N_860,In_1923,In_948);
nand U861 (N_861,In_187,In_1475);
xnor U862 (N_862,In_1000,In_488);
nand U863 (N_863,In_590,In_1626);
or U864 (N_864,In_319,In_19);
nand U865 (N_865,In_99,In_1350);
and U866 (N_866,In_1362,In_813);
nand U867 (N_867,In_1459,In_1095);
and U868 (N_868,In_1859,In_233);
or U869 (N_869,In_345,In_993);
xnor U870 (N_870,In_532,In_508);
nand U871 (N_871,In_855,In_1851);
nand U872 (N_872,In_81,In_282);
and U873 (N_873,In_1646,In_1970);
nand U874 (N_874,In_552,In_1159);
and U875 (N_875,In_838,In_1068);
nor U876 (N_876,In_1195,In_208);
nor U877 (N_877,In_1297,In_1208);
nor U878 (N_878,In_587,In_770);
nand U879 (N_879,In_356,In_1809);
or U880 (N_880,In_1517,In_784);
or U881 (N_881,In_502,In_586);
and U882 (N_882,In_509,In_1389);
or U883 (N_883,In_841,In_1480);
nand U884 (N_884,In_1494,In_1127);
or U885 (N_885,In_1359,In_1269);
or U886 (N_886,In_525,In_1917);
xnor U887 (N_887,In_1616,In_1548);
xor U888 (N_888,In_1130,In_202);
xnor U889 (N_889,In_1691,In_616);
nor U890 (N_890,In_825,In_589);
nand U891 (N_891,In_893,In_1299);
nand U892 (N_892,In_1132,In_1460);
or U893 (N_893,In_576,In_1787);
nand U894 (N_894,In_154,In_162);
or U895 (N_895,In_1190,In_967);
nand U896 (N_896,In_716,In_804);
nand U897 (N_897,In_699,In_767);
and U898 (N_898,In_563,In_620);
and U899 (N_899,In_1165,In_1186);
and U900 (N_900,In_1312,In_708);
nand U901 (N_901,In_881,In_1272);
nor U902 (N_902,In_431,In_1689);
and U903 (N_903,In_786,In_1690);
or U904 (N_904,In_1586,In_194);
xor U905 (N_905,In_602,In_412);
nand U906 (N_906,In_357,In_996);
and U907 (N_907,In_478,In_856);
xnor U908 (N_908,In_221,In_1533);
nand U909 (N_909,In_505,In_1855);
and U910 (N_910,In_649,In_1045);
or U911 (N_911,In_718,In_1918);
and U912 (N_912,In_920,In_253);
or U913 (N_913,In_277,In_1223);
and U914 (N_914,In_614,In_1199);
xnor U915 (N_915,In_222,In_1994);
and U916 (N_916,In_529,In_1337);
or U917 (N_917,In_788,In_1243);
nand U918 (N_918,In_1210,In_322);
and U919 (N_919,In_1069,In_22);
and U920 (N_920,In_1137,In_689);
xor U921 (N_921,In_1801,In_132);
nand U922 (N_922,In_626,In_1298);
nand U923 (N_923,In_987,In_1493);
and U924 (N_924,In_1450,In_225);
nand U925 (N_925,In_1543,In_1158);
and U926 (N_926,In_472,In_1542);
and U927 (N_927,In_229,In_745);
or U928 (N_928,In_1773,In_1769);
nand U929 (N_929,In_311,In_1598);
and U930 (N_930,In_490,In_673);
xor U931 (N_931,In_1462,In_407);
nor U932 (N_932,In_1589,In_1641);
xnor U933 (N_933,In_1461,In_1836);
and U934 (N_934,In_1338,In_477);
nor U935 (N_935,In_1355,In_1518);
or U936 (N_936,In_878,In_1702);
and U937 (N_937,In_725,In_1783);
or U938 (N_938,In_1366,In_585);
nor U939 (N_939,In_1340,In_1649);
and U940 (N_940,In_635,In_1818);
nand U941 (N_941,In_990,In_1401);
nand U942 (N_942,In_4,In_157);
nand U943 (N_943,In_543,In_1875);
xor U944 (N_944,In_1725,In_58);
or U945 (N_945,In_863,In_599);
or U946 (N_946,In_853,In_1858);
and U947 (N_947,In_31,In_1944);
nor U948 (N_948,In_1541,In_296);
or U949 (N_949,In_398,In_1741);
nand U950 (N_950,In_1521,In_1048);
and U951 (N_951,In_496,In_1592);
nor U952 (N_952,In_646,In_1187);
xnor U953 (N_953,In_1468,In_860);
or U954 (N_954,In_1886,In_227);
nor U955 (N_955,In_1497,In_1791);
nor U956 (N_956,In_1038,In_1445);
nand U957 (N_957,In_374,In_1273);
nand U958 (N_958,In_1092,In_518);
nand U959 (N_959,In_709,In_168);
or U960 (N_960,In_1281,In_1549);
nor U961 (N_961,In_1504,In_603);
nor U962 (N_962,In_1162,In_385);
nand U963 (N_963,In_1437,In_1897);
xnor U964 (N_964,In_1283,In_728);
or U965 (N_965,In_1284,In_1221);
xnor U966 (N_966,In_1704,In_1036);
nor U967 (N_967,In_630,In_686);
or U968 (N_968,In_1904,In_423);
nand U969 (N_969,In_903,In_1222);
nor U970 (N_970,In_348,In_1974);
or U971 (N_971,In_1778,In_1839);
nand U972 (N_972,In_557,In_321);
nor U973 (N_973,In_104,In_378);
nand U974 (N_974,In_1290,In_1880);
xnor U975 (N_975,In_129,In_1005);
or U976 (N_976,In_91,In_1110);
nand U977 (N_977,In_724,In_405);
nand U978 (N_978,In_1567,In_807);
or U979 (N_979,In_1153,In_134);
or U980 (N_980,In_783,In_1348);
nor U981 (N_981,In_1805,In_1334);
nor U982 (N_982,In_1042,In_24);
nand U983 (N_983,In_1100,In_1632);
nor U984 (N_984,In_123,In_879);
and U985 (N_985,In_1550,In_1499);
nand U986 (N_986,In_1314,In_1254);
nand U987 (N_987,In_11,In_598);
or U988 (N_988,In_1022,In_1029);
and U989 (N_989,In_1750,In_870);
nor U990 (N_990,In_622,In_1824);
nand U991 (N_991,In_447,In_1575);
and U992 (N_992,In_925,In_1951);
nand U993 (N_993,In_498,In_1837);
nand U994 (N_994,In_1203,In_1315);
nor U995 (N_995,In_1625,In_1230);
nand U996 (N_996,In_1227,In_629);
or U997 (N_997,In_1862,In_869);
nor U998 (N_998,In_558,In_80);
nand U999 (N_999,In_1614,In_1569);
nand U1000 (N_1000,In_612,In_510);
nor U1001 (N_1001,In_636,In_1668);
and U1002 (N_1002,In_746,In_367);
or U1003 (N_1003,In_570,In_681);
nand U1004 (N_1004,In_679,In_1521);
xor U1005 (N_1005,In_1109,In_41);
xnor U1006 (N_1006,In_1808,In_1077);
nor U1007 (N_1007,In_1944,In_283);
or U1008 (N_1008,In_1714,In_993);
and U1009 (N_1009,In_1565,In_967);
or U1010 (N_1010,In_1383,In_488);
nand U1011 (N_1011,In_1826,In_568);
nor U1012 (N_1012,In_1844,In_703);
nor U1013 (N_1013,In_120,In_460);
and U1014 (N_1014,In_84,In_1722);
and U1015 (N_1015,In_971,In_602);
nand U1016 (N_1016,In_392,In_1146);
nor U1017 (N_1017,In_539,In_951);
nand U1018 (N_1018,In_1756,In_347);
nand U1019 (N_1019,In_1655,In_120);
and U1020 (N_1020,In_1308,In_750);
xor U1021 (N_1021,In_576,In_873);
nand U1022 (N_1022,In_161,In_1031);
nor U1023 (N_1023,In_1805,In_1832);
nor U1024 (N_1024,In_1483,In_1974);
nor U1025 (N_1025,In_1859,In_1039);
and U1026 (N_1026,In_681,In_1884);
or U1027 (N_1027,In_1226,In_995);
nor U1028 (N_1028,In_710,In_1656);
nand U1029 (N_1029,In_309,In_230);
nor U1030 (N_1030,In_1316,In_162);
nand U1031 (N_1031,In_447,In_923);
nor U1032 (N_1032,In_997,In_1078);
and U1033 (N_1033,In_1197,In_1757);
nor U1034 (N_1034,In_1683,In_1497);
and U1035 (N_1035,In_1633,In_601);
and U1036 (N_1036,In_765,In_425);
xnor U1037 (N_1037,In_1015,In_1491);
or U1038 (N_1038,In_229,In_1195);
nor U1039 (N_1039,In_1155,In_454);
and U1040 (N_1040,In_809,In_1210);
nand U1041 (N_1041,In_1226,In_22);
and U1042 (N_1042,In_916,In_1345);
nand U1043 (N_1043,In_1793,In_1720);
or U1044 (N_1044,In_1464,In_1259);
or U1045 (N_1045,In_1853,In_144);
and U1046 (N_1046,In_1355,In_1521);
nor U1047 (N_1047,In_349,In_1054);
or U1048 (N_1048,In_50,In_72);
nor U1049 (N_1049,In_1467,In_416);
nand U1050 (N_1050,In_1457,In_171);
xor U1051 (N_1051,In_836,In_628);
nand U1052 (N_1052,In_671,In_1603);
and U1053 (N_1053,In_1938,In_807);
nor U1054 (N_1054,In_1883,In_424);
nand U1055 (N_1055,In_1470,In_1917);
xor U1056 (N_1056,In_840,In_80);
and U1057 (N_1057,In_583,In_1821);
or U1058 (N_1058,In_1603,In_1778);
nand U1059 (N_1059,In_1518,In_1796);
and U1060 (N_1060,In_1223,In_1679);
nor U1061 (N_1061,In_391,In_230);
or U1062 (N_1062,In_1040,In_666);
nand U1063 (N_1063,In_1427,In_449);
or U1064 (N_1064,In_948,In_1015);
nor U1065 (N_1065,In_1364,In_1908);
and U1066 (N_1066,In_1991,In_90);
nor U1067 (N_1067,In_1334,In_1541);
or U1068 (N_1068,In_1258,In_486);
nand U1069 (N_1069,In_631,In_202);
or U1070 (N_1070,In_1591,In_168);
or U1071 (N_1071,In_115,In_1007);
or U1072 (N_1072,In_846,In_1677);
or U1073 (N_1073,In_1869,In_206);
or U1074 (N_1074,In_1412,In_899);
and U1075 (N_1075,In_1590,In_653);
or U1076 (N_1076,In_1515,In_1273);
or U1077 (N_1077,In_1330,In_1482);
xnor U1078 (N_1078,In_1493,In_24);
nand U1079 (N_1079,In_1109,In_976);
nor U1080 (N_1080,In_738,In_1186);
xor U1081 (N_1081,In_1737,In_769);
nor U1082 (N_1082,In_789,In_1644);
nor U1083 (N_1083,In_1317,In_903);
or U1084 (N_1084,In_1321,In_1817);
nand U1085 (N_1085,In_1629,In_1265);
xnor U1086 (N_1086,In_32,In_1056);
or U1087 (N_1087,In_811,In_132);
or U1088 (N_1088,In_108,In_807);
nand U1089 (N_1089,In_1680,In_1310);
and U1090 (N_1090,In_482,In_1187);
nor U1091 (N_1091,In_939,In_706);
nor U1092 (N_1092,In_1148,In_1885);
and U1093 (N_1093,In_1707,In_350);
and U1094 (N_1094,In_339,In_192);
or U1095 (N_1095,In_1742,In_1820);
xnor U1096 (N_1096,In_1879,In_843);
nand U1097 (N_1097,In_1901,In_996);
nor U1098 (N_1098,In_753,In_875);
nand U1099 (N_1099,In_287,In_1177);
nand U1100 (N_1100,In_152,In_1383);
nor U1101 (N_1101,In_348,In_1902);
nand U1102 (N_1102,In_930,In_1625);
and U1103 (N_1103,In_1562,In_1344);
and U1104 (N_1104,In_1770,In_596);
nand U1105 (N_1105,In_105,In_1168);
nand U1106 (N_1106,In_540,In_1122);
or U1107 (N_1107,In_1442,In_66);
and U1108 (N_1108,In_1428,In_489);
and U1109 (N_1109,In_1947,In_1191);
or U1110 (N_1110,In_1654,In_867);
nor U1111 (N_1111,In_700,In_323);
xor U1112 (N_1112,In_1393,In_1575);
nor U1113 (N_1113,In_1221,In_698);
or U1114 (N_1114,In_428,In_1238);
or U1115 (N_1115,In_1890,In_1288);
and U1116 (N_1116,In_962,In_1030);
and U1117 (N_1117,In_1888,In_1833);
or U1118 (N_1118,In_1949,In_752);
or U1119 (N_1119,In_2,In_1154);
xnor U1120 (N_1120,In_467,In_1990);
nor U1121 (N_1121,In_43,In_704);
nor U1122 (N_1122,In_344,In_1206);
nand U1123 (N_1123,In_613,In_650);
xnor U1124 (N_1124,In_32,In_721);
or U1125 (N_1125,In_1076,In_929);
or U1126 (N_1126,In_546,In_1810);
or U1127 (N_1127,In_1185,In_243);
xor U1128 (N_1128,In_1484,In_1780);
xnor U1129 (N_1129,In_1126,In_50);
nand U1130 (N_1130,In_587,In_190);
and U1131 (N_1131,In_173,In_1479);
nand U1132 (N_1132,In_1389,In_1406);
nor U1133 (N_1133,In_1513,In_589);
xor U1134 (N_1134,In_258,In_1598);
and U1135 (N_1135,In_300,In_1144);
or U1136 (N_1136,In_1709,In_1883);
xor U1137 (N_1137,In_1538,In_762);
nor U1138 (N_1138,In_1289,In_11);
nor U1139 (N_1139,In_276,In_1434);
nand U1140 (N_1140,In_1929,In_1453);
and U1141 (N_1141,In_1198,In_1327);
or U1142 (N_1142,In_1932,In_1535);
nor U1143 (N_1143,In_1830,In_125);
or U1144 (N_1144,In_763,In_1266);
nor U1145 (N_1145,In_700,In_1809);
nand U1146 (N_1146,In_1613,In_1276);
nand U1147 (N_1147,In_1352,In_1373);
nand U1148 (N_1148,In_504,In_1428);
nand U1149 (N_1149,In_410,In_288);
xor U1150 (N_1150,In_1145,In_406);
nor U1151 (N_1151,In_140,In_843);
xor U1152 (N_1152,In_142,In_653);
nand U1153 (N_1153,In_1648,In_365);
nor U1154 (N_1154,In_200,In_339);
nand U1155 (N_1155,In_1462,In_1010);
or U1156 (N_1156,In_591,In_1743);
nor U1157 (N_1157,In_585,In_820);
nor U1158 (N_1158,In_932,In_771);
nand U1159 (N_1159,In_461,In_206);
or U1160 (N_1160,In_664,In_729);
or U1161 (N_1161,In_1831,In_976);
or U1162 (N_1162,In_166,In_1216);
nor U1163 (N_1163,In_1815,In_924);
nand U1164 (N_1164,In_736,In_301);
nand U1165 (N_1165,In_735,In_25);
nor U1166 (N_1166,In_240,In_878);
and U1167 (N_1167,In_476,In_985);
nand U1168 (N_1168,In_605,In_1648);
nor U1169 (N_1169,In_337,In_1808);
and U1170 (N_1170,In_158,In_724);
and U1171 (N_1171,In_806,In_652);
nor U1172 (N_1172,In_1543,In_1161);
nor U1173 (N_1173,In_692,In_1297);
nor U1174 (N_1174,In_1238,In_1099);
and U1175 (N_1175,In_1631,In_66);
or U1176 (N_1176,In_1594,In_1698);
nor U1177 (N_1177,In_871,In_153);
or U1178 (N_1178,In_148,In_1880);
nand U1179 (N_1179,In_1216,In_924);
and U1180 (N_1180,In_38,In_1541);
nor U1181 (N_1181,In_466,In_751);
nand U1182 (N_1182,In_1605,In_333);
nor U1183 (N_1183,In_1398,In_1071);
nor U1184 (N_1184,In_1769,In_1368);
or U1185 (N_1185,In_430,In_1048);
and U1186 (N_1186,In_1327,In_825);
nand U1187 (N_1187,In_1115,In_1901);
nand U1188 (N_1188,In_1634,In_1609);
nor U1189 (N_1189,In_1527,In_1125);
nor U1190 (N_1190,In_907,In_1897);
and U1191 (N_1191,In_1499,In_1636);
nor U1192 (N_1192,In_1745,In_1656);
or U1193 (N_1193,In_1590,In_813);
nand U1194 (N_1194,In_1992,In_188);
or U1195 (N_1195,In_1955,In_1112);
nor U1196 (N_1196,In_282,In_1329);
nand U1197 (N_1197,In_137,In_283);
nand U1198 (N_1198,In_1242,In_219);
or U1199 (N_1199,In_809,In_1285);
nand U1200 (N_1200,In_1998,In_1602);
xor U1201 (N_1201,In_120,In_843);
nor U1202 (N_1202,In_1166,In_428);
and U1203 (N_1203,In_1140,In_227);
nand U1204 (N_1204,In_1966,In_647);
and U1205 (N_1205,In_40,In_266);
nand U1206 (N_1206,In_588,In_238);
and U1207 (N_1207,In_897,In_1177);
and U1208 (N_1208,In_740,In_603);
nand U1209 (N_1209,In_570,In_1482);
nor U1210 (N_1210,In_1750,In_1624);
and U1211 (N_1211,In_505,In_1470);
or U1212 (N_1212,In_1873,In_197);
xnor U1213 (N_1213,In_1163,In_1059);
and U1214 (N_1214,In_565,In_908);
and U1215 (N_1215,In_1103,In_1325);
xor U1216 (N_1216,In_229,In_1778);
and U1217 (N_1217,In_1858,In_1639);
or U1218 (N_1218,In_1242,In_682);
nand U1219 (N_1219,In_638,In_236);
or U1220 (N_1220,In_400,In_1051);
and U1221 (N_1221,In_1366,In_1476);
xor U1222 (N_1222,In_1290,In_495);
nand U1223 (N_1223,In_50,In_1534);
nor U1224 (N_1224,In_277,In_1029);
nand U1225 (N_1225,In_1045,In_790);
nor U1226 (N_1226,In_892,In_1493);
xnor U1227 (N_1227,In_1780,In_643);
nor U1228 (N_1228,In_1716,In_1183);
nand U1229 (N_1229,In_1558,In_371);
or U1230 (N_1230,In_626,In_1183);
nand U1231 (N_1231,In_134,In_807);
nor U1232 (N_1232,In_1598,In_177);
nor U1233 (N_1233,In_1039,In_1551);
nor U1234 (N_1234,In_1399,In_167);
nor U1235 (N_1235,In_1373,In_526);
xnor U1236 (N_1236,In_651,In_1334);
or U1237 (N_1237,In_1239,In_513);
nor U1238 (N_1238,In_1422,In_846);
and U1239 (N_1239,In_1022,In_1582);
nor U1240 (N_1240,In_828,In_1325);
and U1241 (N_1241,In_327,In_1154);
and U1242 (N_1242,In_1169,In_1580);
nor U1243 (N_1243,In_1624,In_70);
nor U1244 (N_1244,In_93,In_757);
nor U1245 (N_1245,In_1360,In_1874);
nor U1246 (N_1246,In_183,In_1570);
and U1247 (N_1247,In_325,In_1381);
nand U1248 (N_1248,In_736,In_1020);
nand U1249 (N_1249,In_1267,In_1251);
nand U1250 (N_1250,In_1759,In_421);
and U1251 (N_1251,In_1173,In_576);
nor U1252 (N_1252,In_1813,In_870);
and U1253 (N_1253,In_220,In_1887);
or U1254 (N_1254,In_1134,In_336);
and U1255 (N_1255,In_255,In_1612);
nor U1256 (N_1256,In_1378,In_1719);
xor U1257 (N_1257,In_286,In_1375);
nand U1258 (N_1258,In_312,In_888);
nand U1259 (N_1259,In_690,In_693);
xor U1260 (N_1260,In_1602,In_1272);
or U1261 (N_1261,In_1366,In_1381);
and U1262 (N_1262,In_832,In_609);
and U1263 (N_1263,In_507,In_77);
nand U1264 (N_1264,In_1313,In_1883);
and U1265 (N_1265,In_97,In_409);
nand U1266 (N_1266,In_826,In_955);
nor U1267 (N_1267,In_1424,In_64);
nand U1268 (N_1268,In_1037,In_47);
nand U1269 (N_1269,In_607,In_136);
and U1270 (N_1270,In_1771,In_1484);
nand U1271 (N_1271,In_159,In_806);
or U1272 (N_1272,In_1657,In_208);
nor U1273 (N_1273,In_1627,In_1841);
and U1274 (N_1274,In_888,In_1552);
nand U1275 (N_1275,In_391,In_1888);
nor U1276 (N_1276,In_734,In_672);
and U1277 (N_1277,In_1421,In_1629);
nand U1278 (N_1278,In_1076,In_1168);
nand U1279 (N_1279,In_1187,In_271);
nand U1280 (N_1280,In_822,In_1434);
nor U1281 (N_1281,In_179,In_906);
nor U1282 (N_1282,In_827,In_777);
nor U1283 (N_1283,In_1426,In_1060);
or U1284 (N_1284,In_283,In_1536);
or U1285 (N_1285,In_804,In_1250);
or U1286 (N_1286,In_683,In_1708);
nand U1287 (N_1287,In_1767,In_393);
or U1288 (N_1288,In_501,In_1908);
xnor U1289 (N_1289,In_1053,In_1498);
or U1290 (N_1290,In_202,In_1148);
nand U1291 (N_1291,In_63,In_113);
nor U1292 (N_1292,In_1245,In_940);
or U1293 (N_1293,In_619,In_76);
nor U1294 (N_1294,In_1645,In_539);
nand U1295 (N_1295,In_574,In_354);
or U1296 (N_1296,In_1366,In_144);
nor U1297 (N_1297,In_272,In_793);
or U1298 (N_1298,In_911,In_286);
nand U1299 (N_1299,In_1439,In_1622);
nor U1300 (N_1300,In_134,In_864);
nand U1301 (N_1301,In_1665,In_1234);
nand U1302 (N_1302,In_87,In_479);
and U1303 (N_1303,In_1471,In_1351);
xnor U1304 (N_1304,In_695,In_497);
and U1305 (N_1305,In_1138,In_1651);
nor U1306 (N_1306,In_297,In_1629);
and U1307 (N_1307,In_1540,In_1508);
nand U1308 (N_1308,In_717,In_666);
nor U1309 (N_1309,In_1399,In_534);
and U1310 (N_1310,In_1483,In_1618);
or U1311 (N_1311,In_1392,In_268);
or U1312 (N_1312,In_742,In_902);
xnor U1313 (N_1313,In_524,In_1569);
nor U1314 (N_1314,In_1843,In_1993);
or U1315 (N_1315,In_828,In_1);
or U1316 (N_1316,In_124,In_1628);
nor U1317 (N_1317,In_881,In_1540);
or U1318 (N_1318,In_558,In_794);
and U1319 (N_1319,In_827,In_1142);
nand U1320 (N_1320,In_1708,In_1236);
nor U1321 (N_1321,In_697,In_412);
nor U1322 (N_1322,In_1533,In_849);
xnor U1323 (N_1323,In_907,In_639);
nand U1324 (N_1324,In_1809,In_1067);
xnor U1325 (N_1325,In_854,In_558);
nor U1326 (N_1326,In_1483,In_1851);
or U1327 (N_1327,In_121,In_939);
and U1328 (N_1328,In_1185,In_131);
nor U1329 (N_1329,In_1971,In_97);
nand U1330 (N_1330,In_1594,In_1780);
and U1331 (N_1331,In_1673,In_1868);
nand U1332 (N_1332,In_592,In_774);
or U1333 (N_1333,In_1598,In_646);
nand U1334 (N_1334,In_619,In_1620);
and U1335 (N_1335,In_852,In_1947);
nand U1336 (N_1336,In_1030,In_319);
nor U1337 (N_1337,In_986,In_1589);
or U1338 (N_1338,In_1125,In_864);
nand U1339 (N_1339,In_102,In_1787);
nor U1340 (N_1340,In_226,In_1453);
or U1341 (N_1341,In_1399,In_1682);
or U1342 (N_1342,In_1804,In_32);
and U1343 (N_1343,In_29,In_590);
or U1344 (N_1344,In_796,In_1582);
nand U1345 (N_1345,In_1767,In_1876);
nand U1346 (N_1346,In_896,In_1989);
nand U1347 (N_1347,In_1366,In_551);
xor U1348 (N_1348,In_1326,In_704);
nand U1349 (N_1349,In_1803,In_746);
nand U1350 (N_1350,In_575,In_835);
or U1351 (N_1351,In_1720,In_1869);
nor U1352 (N_1352,In_1131,In_1005);
xnor U1353 (N_1353,In_1343,In_8);
xnor U1354 (N_1354,In_1763,In_129);
or U1355 (N_1355,In_1363,In_1545);
and U1356 (N_1356,In_1324,In_1966);
nor U1357 (N_1357,In_1328,In_382);
nand U1358 (N_1358,In_1820,In_624);
xnor U1359 (N_1359,In_1487,In_381);
and U1360 (N_1360,In_1351,In_284);
or U1361 (N_1361,In_634,In_719);
nand U1362 (N_1362,In_1073,In_1384);
nor U1363 (N_1363,In_155,In_627);
nand U1364 (N_1364,In_1585,In_487);
and U1365 (N_1365,In_1179,In_391);
nor U1366 (N_1366,In_1319,In_363);
nor U1367 (N_1367,In_857,In_323);
nor U1368 (N_1368,In_864,In_1007);
nor U1369 (N_1369,In_1978,In_1633);
and U1370 (N_1370,In_933,In_1164);
and U1371 (N_1371,In_185,In_1164);
nand U1372 (N_1372,In_574,In_1854);
xnor U1373 (N_1373,In_1305,In_1785);
or U1374 (N_1374,In_1251,In_1381);
xnor U1375 (N_1375,In_1564,In_771);
xor U1376 (N_1376,In_587,In_684);
nor U1377 (N_1377,In_1098,In_171);
nor U1378 (N_1378,In_17,In_127);
nor U1379 (N_1379,In_1868,In_397);
or U1380 (N_1380,In_647,In_864);
or U1381 (N_1381,In_1907,In_1318);
nand U1382 (N_1382,In_59,In_1019);
xnor U1383 (N_1383,In_1042,In_1503);
nor U1384 (N_1384,In_1043,In_1537);
nor U1385 (N_1385,In_1143,In_1681);
xnor U1386 (N_1386,In_136,In_896);
nor U1387 (N_1387,In_960,In_1205);
or U1388 (N_1388,In_820,In_1991);
and U1389 (N_1389,In_71,In_581);
nor U1390 (N_1390,In_1635,In_228);
or U1391 (N_1391,In_1406,In_1190);
xnor U1392 (N_1392,In_33,In_1497);
or U1393 (N_1393,In_39,In_1828);
or U1394 (N_1394,In_221,In_870);
or U1395 (N_1395,In_911,In_1068);
nor U1396 (N_1396,In_402,In_1303);
nor U1397 (N_1397,In_763,In_1427);
nor U1398 (N_1398,In_850,In_1965);
or U1399 (N_1399,In_1887,In_906);
nand U1400 (N_1400,In_520,In_913);
nor U1401 (N_1401,In_1834,In_967);
nand U1402 (N_1402,In_580,In_1120);
or U1403 (N_1403,In_1905,In_1404);
or U1404 (N_1404,In_1829,In_1244);
and U1405 (N_1405,In_1678,In_1612);
and U1406 (N_1406,In_405,In_447);
nor U1407 (N_1407,In_1282,In_1394);
or U1408 (N_1408,In_221,In_296);
nor U1409 (N_1409,In_1223,In_899);
or U1410 (N_1410,In_1445,In_960);
nor U1411 (N_1411,In_1623,In_1676);
nor U1412 (N_1412,In_1495,In_770);
nor U1413 (N_1413,In_581,In_1203);
or U1414 (N_1414,In_530,In_286);
nor U1415 (N_1415,In_309,In_1991);
and U1416 (N_1416,In_1999,In_408);
nand U1417 (N_1417,In_1425,In_860);
nor U1418 (N_1418,In_596,In_502);
and U1419 (N_1419,In_1113,In_823);
nand U1420 (N_1420,In_1707,In_191);
nor U1421 (N_1421,In_609,In_1079);
nand U1422 (N_1422,In_971,In_1098);
and U1423 (N_1423,In_1527,In_1189);
and U1424 (N_1424,In_1527,In_1765);
nand U1425 (N_1425,In_202,In_983);
nor U1426 (N_1426,In_949,In_188);
nand U1427 (N_1427,In_1810,In_1727);
nor U1428 (N_1428,In_1942,In_641);
and U1429 (N_1429,In_542,In_968);
xor U1430 (N_1430,In_426,In_1048);
nor U1431 (N_1431,In_934,In_557);
or U1432 (N_1432,In_904,In_1772);
and U1433 (N_1433,In_1716,In_76);
nor U1434 (N_1434,In_509,In_1350);
nand U1435 (N_1435,In_1707,In_1291);
nor U1436 (N_1436,In_224,In_1854);
or U1437 (N_1437,In_793,In_1764);
nor U1438 (N_1438,In_760,In_1866);
xnor U1439 (N_1439,In_1437,In_1388);
nor U1440 (N_1440,In_452,In_1656);
nor U1441 (N_1441,In_1921,In_1702);
and U1442 (N_1442,In_1748,In_1379);
xnor U1443 (N_1443,In_976,In_980);
or U1444 (N_1444,In_751,In_1213);
and U1445 (N_1445,In_1123,In_1318);
nand U1446 (N_1446,In_821,In_1549);
and U1447 (N_1447,In_642,In_597);
xor U1448 (N_1448,In_368,In_1212);
or U1449 (N_1449,In_1651,In_73);
or U1450 (N_1450,In_1304,In_1590);
and U1451 (N_1451,In_886,In_225);
or U1452 (N_1452,In_1975,In_467);
nand U1453 (N_1453,In_200,In_1818);
nand U1454 (N_1454,In_1673,In_480);
or U1455 (N_1455,In_1704,In_43);
and U1456 (N_1456,In_1869,In_130);
nor U1457 (N_1457,In_1163,In_1242);
nand U1458 (N_1458,In_1,In_444);
nor U1459 (N_1459,In_1428,In_377);
or U1460 (N_1460,In_727,In_1837);
or U1461 (N_1461,In_567,In_148);
or U1462 (N_1462,In_865,In_368);
nor U1463 (N_1463,In_1057,In_449);
nor U1464 (N_1464,In_1101,In_1727);
nand U1465 (N_1465,In_1441,In_1272);
nor U1466 (N_1466,In_1305,In_1848);
or U1467 (N_1467,In_1952,In_283);
and U1468 (N_1468,In_1105,In_95);
nand U1469 (N_1469,In_1661,In_477);
or U1470 (N_1470,In_112,In_885);
or U1471 (N_1471,In_104,In_112);
nand U1472 (N_1472,In_320,In_921);
nand U1473 (N_1473,In_683,In_727);
nor U1474 (N_1474,In_141,In_1222);
and U1475 (N_1475,In_1164,In_912);
and U1476 (N_1476,In_47,In_969);
or U1477 (N_1477,In_764,In_974);
or U1478 (N_1478,In_1894,In_1736);
and U1479 (N_1479,In_1611,In_508);
nand U1480 (N_1480,In_77,In_1101);
nand U1481 (N_1481,In_823,In_1112);
and U1482 (N_1482,In_1337,In_1257);
nor U1483 (N_1483,In_186,In_1722);
and U1484 (N_1484,In_1666,In_1689);
xnor U1485 (N_1485,In_1792,In_1957);
and U1486 (N_1486,In_511,In_1379);
xor U1487 (N_1487,In_112,In_1450);
and U1488 (N_1488,In_915,In_421);
nor U1489 (N_1489,In_886,In_1978);
nor U1490 (N_1490,In_1599,In_551);
or U1491 (N_1491,In_437,In_239);
and U1492 (N_1492,In_1574,In_26);
nand U1493 (N_1493,In_340,In_160);
and U1494 (N_1494,In_1323,In_698);
nand U1495 (N_1495,In_486,In_741);
nand U1496 (N_1496,In_1708,In_716);
and U1497 (N_1497,In_791,In_163);
and U1498 (N_1498,In_1484,In_521);
nand U1499 (N_1499,In_1088,In_393);
and U1500 (N_1500,In_1080,In_1457);
nor U1501 (N_1501,In_1305,In_1047);
nor U1502 (N_1502,In_335,In_733);
or U1503 (N_1503,In_685,In_85);
nand U1504 (N_1504,In_1731,In_1369);
nor U1505 (N_1505,In_1047,In_269);
and U1506 (N_1506,In_102,In_553);
and U1507 (N_1507,In_1834,In_1722);
nor U1508 (N_1508,In_1095,In_1308);
or U1509 (N_1509,In_585,In_1031);
or U1510 (N_1510,In_1843,In_279);
and U1511 (N_1511,In_902,In_654);
and U1512 (N_1512,In_1055,In_253);
nand U1513 (N_1513,In_1131,In_840);
or U1514 (N_1514,In_589,In_1067);
nor U1515 (N_1515,In_404,In_577);
nand U1516 (N_1516,In_985,In_1937);
or U1517 (N_1517,In_1558,In_1177);
nand U1518 (N_1518,In_1683,In_1572);
and U1519 (N_1519,In_1264,In_194);
nor U1520 (N_1520,In_819,In_1738);
nand U1521 (N_1521,In_1520,In_1287);
nor U1522 (N_1522,In_1733,In_991);
nor U1523 (N_1523,In_1284,In_1018);
and U1524 (N_1524,In_1342,In_160);
or U1525 (N_1525,In_1736,In_1668);
and U1526 (N_1526,In_1203,In_1880);
and U1527 (N_1527,In_418,In_816);
nor U1528 (N_1528,In_1239,In_968);
nand U1529 (N_1529,In_1282,In_1972);
or U1530 (N_1530,In_1545,In_1661);
nor U1531 (N_1531,In_1023,In_1885);
and U1532 (N_1532,In_275,In_389);
xor U1533 (N_1533,In_1168,In_215);
nand U1534 (N_1534,In_15,In_1168);
nor U1535 (N_1535,In_596,In_746);
nor U1536 (N_1536,In_589,In_391);
and U1537 (N_1537,In_1497,In_427);
or U1538 (N_1538,In_884,In_1124);
nor U1539 (N_1539,In_1092,In_1020);
nand U1540 (N_1540,In_1407,In_966);
or U1541 (N_1541,In_708,In_133);
nand U1542 (N_1542,In_415,In_1989);
nand U1543 (N_1543,In_770,In_1019);
and U1544 (N_1544,In_931,In_81);
or U1545 (N_1545,In_1917,In_1980);
or U1546 (N_1546,In_1582,In_147);
nor U1547 (N_1547,In_1102,In_283);
nor U1548 (N_1548,In_1249,In_578);
nand U1549 (N_1549,In_1677,In_1536);
nand U1550 (N_1550,In_1719,In_1122);
and U1551 (N_1551,In_1847,In_675);
and U1552 (N_1552,In_1916,In_402);
or U1553 (N_1553,In_1297,In_68);
or U1554 (N_1554,In_1466,In_1845);
xnor U1555 (N_1555,In_571,In_698);
nand U1556 (N_1556,In_70,In_239);
xor U1557 (N_1557,In_660,In_1022);
nand U1558 (N_1558,In_229,In_1020);
or U1559 (N_1559,In_1841,In_474);
and U1560 (N_1560,In_1435,In_590);
nand U1561 (N_1561,In_126,In_985);
or U1562 (N_1562,In_1241,In_1534);
and U1563 (N_1563,In_935,In_706);
nor U1564 (N_1564,In_1289,In_669);
nand U1565 (N_1565,In_1464,In_586);
nor U1566 (N_1566,In_1438,In_1445);
and U1567 (N_1567,In_1640,In_1772);
nand U1568 (N_1568,In_1338,In_1829);
and U1569 (N_1569,In_369,In_591);
nand U1570 (N_1570,In_426,In_1936);
xnor U1571 (N_1571,In_1153,In_87);
and U1572 (N_1572,In_400,In_1621);
and U1573 (N_1573,In_1602,In_1509);
nand U1574 (N_1574,In_1868,In_479);
and U1575 (N_1575,In_1510,In_435);
nand U1576 (N_1576,In_565,In_1788);
nor U1577 (N_1577,In_594,In_1541);
nand U1578 (N_1578,In_937,In_1806);
xnor U1579 (N_1579,In_987,In_494);
and U1580 (N_1580,In_1014,In_1415);
and U1581 (N_1581,In_434,In_1445);
or U1582 (N_1582,In_1347,In_330);
nand U1583 (N_1583,In_1738,In_1407);
nor U1584 (N_1584,In_564,In_1872);
nand U1585 (N_1585,In_265,In_1761);
nand U1586 (N_1586,In_1236,In_1377);
nor U1587 (N_1587,In_968,In_760);
and U1588 (N_1588,In_1986,In_538);
nand U1589 (N_1589,In_174,In_1805);
nand U1590 (N_1590,In_125,In_1377);
or U1591 (N_1591,In_190,In_1718);
nor U1592 (N_1592,In_177,In_1480);
and U1593 (N_1593,In_75,In_1950);
and U1594 (N_1594,In_1197,In_601);
and U1595 (N_1595,In_1769,In_795);
nand U1596 (N_1596,In_1079,In_1600);
nor U1597 (N_1597,In_131,In_1585);
nor U1598 (N_1598,In_1970,In_590);
or U1599 (N_1599,In_1242,In_236);
nor U1600 (N_1600,In_1121,In_1301);
nor U1601 (N_1601,In_1032,In_406);
nor U1602 (N_1602,In_779,In_664);
or U1603 (N_1603,In_609,In_1331);
or U1604 (N_1604,In_1818,In_1569);
or U1605 (N_1605,In_1608,In_1087);
and U1606 (N_1606,In_98,In_752);
nand U1607 (N_1607,In_978,In_2);
and U1608 (N_1608,In_1329,In_617);
or U1609 (N_1609,In_1159,In_476);
nor U1610 (N_1610,In_1242,In_963);
nor U1611 (N_1611,In_1465,In_1507);
nor U1612 (N_1612,In_1049,In_244);
or U1613 (N_1613,In_558,In_990);
or U1614 (N_1614,In_1480,In_1841);
nor U1615 (N_1615,In_1624,In_274);
or U1616 (N_1616,In_28,In_415);
nor U1617 (N_1617,In_1871,In_1930);
nand U1618 (N_1618,In_1464,In_277);
nand U1619 (N_1619,In_1345,In_890);
and U1620 (N_1620,In_232,In_306);
or U1621 (N_1621,In_41,In_766);
nand U1622 (N_1622,In_702,In_175);
nand U1623 (N_1623,In_198,In_785);
nand U1624 (N_1624,In_1466,In_1685);
nand U1625 (N_1625,In_1185,In_1307);
nor U1626 (N_1626,In_1061,In_389);
or U1627 (N_1627,In_1455,In_511);
nor U1628 (N_1628,In_153,In_1071);
nor U1629 (N_1629,In_1934,In_399);
and U1630 (N_1630,In_37,In_1786);
nor U1631 (N_1631,In_1462,In_94);
nand U1632 (N_1632,In_1877,In_940);
and U1633 (N_1633,In_486,In_898);
nor U1634 (N_1634,In_1355,In_1372);
and U1635 (N_1635,In_1919,In_1697);
xor U1636 (N_1636,In_1073,In_1667);
nand U1637 (N_1637,In_1739,In_1901);
nand U1638 (N_1638,In_921,In_1461);
xnor U1639 (N_1639,In_1772,In_365);
nor U1640 (N_1640,In_1285,In_437);
or U1641 (N_1641,In_740,In_326);
nand U1642 (N_1642,In_939,In_1724);
or U1643 (N_1643,In_618,In_329);
or U1644 (N_1644,In_268,In_1712);
xor U1645 (N_1645,In_877,In_1908);
or U1646 (N_1646,In_625,In_1729);
or U1647 (N_1647,In_829,In_1019);
and U1648 (N_1648,In_734,In_1614);
nor U1649 (N_1649,In_420,In_1956);
nor U1650 (N_1650,In_1993,In_226);
nor U1651 (N_1651,In_59,In_1553);
xor U1652 (N_1652,In_222,In_1567);
nand U1653 (N_1653,In_1667,In_663);
nor U1654 (N_1654,In_238,In_503);
and U1655 (N_1655,In_1274,In_16);
nand U1656 (N_1656,In_1819,In_1345);
nand U1657 (N_1657,In_1637,In_502);
xor U1658 (N_1658,In_1007,In_969);
nand U1659 (N_1659,In_85,In_568);
or U1660 (N_1660,In_34,In_805);
nand U1661 (N_1661,In_658,In_1800);
nor U1662 (N_1662,In_1967,In_330);
and U1663 (N_1663,In_778,In_1412);
nor U1664 (N_1664,In_224,In_646);
or U1665 (N_1665,In_1333,In_1187);
and U1666 (N_1666,In_1191,In_1117);
or U1667 (N_1667,In_738,In_1978);
or U1668 (N_1668,In_1517,In_345);
or U1669 (N_1669,In_1842,In_1830);
xnor U1670 (N_1670,In_1138,In_766);
nor U1671 (N_1671,In_1196,In_1111);
nor U1672 (N_1672,In_1237,In_453);
and U1673 (N_1673,In_1618,In_1513);
nor U1674 (N_1674,In_1176,In_343);
xor U1675 (N_1675,In_207,In_101);
and U1676 (N_1676,In_500,In_1319);
or U1677 (N_1677,In_1663,In_1896);
nand U1678 (N_1678,In_1196,In_1662);
or U1679 (N_1679,In_542,In_159);
nand U1680 (N_1680,In_1154,In_1290);
or U1681 (N_1681,In_283,In_1975);
or U1682 (N_1682,In_307,In_280);
or U1683 (N_1683,In_7,In_1854);
and U1684 (N_1684,In_1478,In_404);
nor U1685 (N_1685,In_768,In_413);
nor U1686 (N_1686,In_55,In_1722);
nor U1687 (N_1687,In_1151,In_1902);
nand U1688 (N_1688,In_1987,In_540);
nor U1689 (N_1689,In_118,In_1539);
or U1690 (N_1690,In_545,In_386);
and U1691 (N_1691,In_654,In_307);
or U1692 (N_1692,In_329,In_230);
nand U1693 (N_1693,In_1224,In_1470);
nand U1694 (N_1694,In_656,In_515);
xor U1695 (N_1695,In_529,In_204);
nor U1696 (N_1696,In_770,In_1591);
and U1697 (N_1697,In_38,In_1225);
or U1698 (N_1698,In_1297,In_503);
or U1699 (N_1699,In_701,In_817);
nor U1700 (N_1700,In_364,In_250);
or U1701 (N_1701,In_124,In_1534);
nor U1702 (N_1702,In_883,In_1864);
nor U1703 (N_1703,In_1684,In_619);
and U1704 (N_1704,In_380,In_330);
and U1705 (N_1705,In_1349,In_683);
xnor U1706 (N_1706,In_673,In_1942);
nor U1707 (N_1707,In_1246,In_611);
and U1708 (N_1708,In_1560,In_1502);
nor U1709 (N_1709,In_336,In_352);
nand U1710 (N_1710,In_1932,In_624);
or U1711 (N_1711,In_865,In_904);
or U1712 (N_1712,In_1405,In_8);
or U1713 (N_1713,In_633,In_1445);
nor U1714 (N_1714,In_1810,In_322);
or U1715 (N_1715,In_1773,In_1095);
nor U1716 (N_1716,In_656,In_1923);
or U1717 (N_1717,In_518,In_1675);
or U1718 (N_1718,In_1603,In_916);
nand U1719 (N_1719,In_230,In_1782);
nand U1720 (N_1720,In_962,In_499);
and U1721 (N_1721,In_1833,In_392);
or U1722 (N_1722,In_598,In_1267);
or U1723 (N_1723,In_1541,In_1077);
or U1724 (N_1724,In_1945,In_987);
or U1725 (N_1725,In_1974,In_1415);
xnor U1726 (N_1726,In_584,In_832);
xor U1727 (N_1727,In_1412,In_1485);
nor U1728 (N_1728,In_1044,In_1033);
nor U1729 (N_1729,In_922,In_1374);
nor U1730 (N_1730,In_55,In_623);
and U1731 (N_1731,In_1614,In_834);
nand U1732 (N_1732,In_1168,In_884);
nor U1733 (N_1733,In_1121,In_297);
and U1734 (N_1734,In_649,In_1781);
and U1735 (N_1735,In_975,In_1077);
nand U1736 (N_1736,In_1588,In_184);
xnor U1737 (N_1737,In_934,In_232);
or U1738 (N_1738,In_999,In_484);
nand U1739 (N_1739,In_128,In_403);
nor U1740 (N_1740,In_1103,In_1171);
nor U1741 (N_1741,In_797,In_488);
nor U1742 (N_1742,In_772,In_1323);
or U1743 (N_1743,In_1107,In_1299);
nand U1744 (N_1744,In_388,In_1450);
and U1745 (N_1745,In_1732,In_1033);
and U1746 (N_1746,In_1401,In_59);
or U1747 (N_1747,In_552,In_394);
nand U1748 (N_1748,In_1356,In_1228);
nand U1749 (N_1749,In_564,In_283);
xor U1750 (N_1750,In_1878,In_300);
nor U1751 (N_1751,In_1613,In_1536);
nor U1752 (N_1752,In_87,In_284);
nand U1753 (N_1753,In_1280,In_1618);
nand U1754 (N_1754,In_1887,In_557);
nand U1755 (N_1755,In_571,In_729);
xor U1756 (N_1756,In_905,In_198);
or U1757 (N_1757,In_1592,In_425);
nand U1758 (N_1758,In_1293,In_1969);
and U1759 (N_1759,In_1003,In_1057);
nor U1760 (N_1760,In_885,In_1852);
or U1761 (N_1761,In_1793,In_1619);
nand U1762 (N_1762,In_1318,In_609);
nor U1763 (N_1763,In_937,In_763);
xor U1764 (N_1764,In_1200,In_1496);
and U1765 (N_1765,In_643,In_1540);
xor U1766 (N_1766,In_128,In_123);
nor U1767 (N_1767,In_1626,In_221);
and U1768 (N_1768,In_1095,In_1251);
xor U1769 (N_1769,In_357,In_1611);
nand U1770 (N_1770,In_609,In_1697);
and U1771 (N_1771,In_1058,In_219);
nor U1772 (N_1772,In_425,In_719);
xor U1773 (N_1773,In_1134,In_1560);
nand U1774 (N_1774,In_1633,In_1969);
nand U1775 (N_1775,In_1778,In_1355);
nand U1776 (N_1776,In_1157,In_1485);
or U1777 (N_1777,In_801,In_1996);
and U1778 (N_1778,In_56,In_1090);
nor U1779 (N_1779,In_643,In_1335);
nand U1780 (N_1780,In_1787,In_1619);
and U1781 (N_1781,In_1055,In_578);
xnor U1782 (N_1782,In_484,In_895);
and U1783 (N_1783,In_1222,In_1874);
and U1784 (N_1784,In_962,In_792);
nand U1785 (N_1785,In_1370,In_1128);
xnor U1786 (N_1786,In_1671,In_1590);
xor U1787 (N_1787,In_1455,In_1925);
nor U1788 (N_1788,In_1777,In_463);
nand U1789 (N_1789,In_145,In_1996);
xor U1790 (N_1790,In_1809,In_1116);
nor U1791 (N_1791,In_744,In_225);
and U1792 (N_1792,In_819,In_1161);
nand U1793 (N_1793,In_1513,In_695);
or U1794 (N_1794,In_1100,In_470);
nor U1795 (N_1795,In_1909,In_926);
and U1796 (N_1796,In_1959,In_1821);
xor U1797 (N_1797,In_892,In_463);
nor U1798 (N_1798,In_1698,In_193);
nand U1799 (N_1799,In_355,In_421);
or U1800 (N_1800,In_591,In_434);
or U1801 (N_1801,In_69,In_710);
or U1802 (N_1802,In_57,In_771);
nor U1803 (N_1803,In_825,In_1096);
or U1804 (N_1804,In_277,In_463);
nand U1805 (N_1805,In_440,In_3);
and U1806 (N_1806,In_329,In_413);
nor U1807 (N_1807,In_1961,In_680);
xnor U1808 (N_1808,In_826,In_1950);
nor U1809 (N_1809,In_482,In_1665);
nand U1810 (N_1810,In_853,In_146);
nor U1811 (N_1811,In_526,In_1809);
nor U1812 (N_1812,In_1222,In_1350);
nand U1813 (N_1813,In_843,In_659);
or U1814 (N_1814,In_208,In_28);
or U1815 (N_1815,In_685,In_22);
nand U1816 (N_1816,In_1447,In_1758);
or U1817 (N_1817,In_755,In_822);
xnor U1818 (N_1818,In_20,In_22);
and U1819 (N_1819,In_110,In_1327);
or U1820 (N_1820,In_1202,In_1694);
nor U1821 (N_1821,In_1071,In_1373);
or U1822 (N_1822,In_1483,In_958);
or U1823 (N_1823,In_1996,In_260);
or U1824 (N_1824,In_928,In_1913);
and U1825 (N_1825,In_1582,In_56);
nor U1826 (N_1826,In_1379,In_1208);
or U1827 (N_1827,In_44,In_296);
or U1828 (N_1828,In_1444,In_100);
or U1829 (N_1829,In_578,In_1622);
and U1830 (N_1830,In_1415,In_862);
nor U1831 (N_1831,In_1066,In_1378);
nor U1832 (N_1832,In_310,In_1643);
nor U1833 (N_1833,In_1860,In_1094);
and U1834 (N_1834,In_1587,In_1608);
and U1835 (N_1835,In_188,In_104);
nand U1836 (N_1836,In_1168,In_1749);
and U1837 (N_1837,In_1026,In_202);
and U1838 (N_1838,In_663,In_1984);
or U1839 (N_1839,In_1857,In_33);
or U1840 (N_1840,In_308,In_817);
nand U1841 (N_1841,In_7,In_1766);
nand U1842 (N_1842,In_100,In_899);
nor U1843 (N_1843,In_1052,In_1140);
nor U1844 (N_1844,In_870,In_99);
and U1845 (N_1845,In_1510,In_366);
and U1846 (N_1846,In_1594,In_349);
nand U1847 (N_1847,In_1135,In_1545);
nor U1848 (N_1848,In_1922,In_1849);
or U1849 (N_1849,In_142,In_156);
and U1850 (N_1850,In_1378,In_781);
nor U1851 (N_1851,In_812,In_1253);
and U1852 (N_1852,In_1019,In_1319);
nand U1853 (N_1853,In_1655,In_184);
or U1854 (N_1854,In_1047,In_277);
nor U1855 (N_1855,In_1452,In_1968);
nand U1856 (N_1856,In_990,In_1505);
nor U1857 (N_1857,In_1642,In_617);
or U1858 (N_1858,In_787,In_455);
nor U1859 (N_1859,In_759,In_386);
xor U1860 (N_1860,In_1560,In_20);
nand U1861 (N_1861,In_934,In_61);
and U1862 (N_1862,In_433,In_1409);
nand U1863 (N_1863,In_1243,In_100);
and U1864 (N_1864,In_878,In_467);
nand U1865 (N_1865,In_1622,In_991);
and U1866 (N_1866,In_653,In_708);
nor U1867 (N_1867,In_911,In_311);
nor U1868 (N_1868,In_536,In_288);
nor U1869 (N_1869,In_1277,In_1898);
nand U1870 (N_1870,In_328,In_1158);
and U1871 (N_1871,In_1559,In_761);
and U1872 (N_1872,In_781,In_808);
and U1873 (N_1873,In_1287,In_1258);
or U1874 (N_1874,In_742,In_1215);
nor U1875 (N_1875,In_753,In_578);
xnor U1876 (N_1876,In_755,In_1648);
and U1877 (N_1877,In_753,In_1693);
nor U1878 (N_1878,In_1194,In_1474);
and U1879 (N_1879,In_1251,In_1541);
and U1880 (N_1880,In_987,In_614);
nand U1881 (N_1881,In_404,In_180);
and U1882 (N_1882,In_1542,In_852);
and U1883 (N_1883,In_1720,In_510);
nand U1884 (N_1884,In_1051,In_1147);
nor U1885 (N_1885,In_179,In_326);
nand U1886 (N_1886,In_1192,In_1664);
nand U1887 (N_1887,In_1414,In_1346);
and U1888 (N_1888,In_412,In_17);
nand U1889 (N_1889,In_1883,In_1170);
nand U1890 (N_1890,In_961,In_1006);
and U1891 (N_1891,In_1966,In_1341);
nor U1892 (N_1892,In_348,In_617);
nor U1893 (N_1893,In_1004,In_1860);
nor U1894 (N_1894,In_1812,In_247);
or U1895 (N_1895,In_137,In_1751);
or U1896 (N_1896,In_469,In_129);
or U1897 (N_1897,In_1724,In_733);
nor U1898 (N_1898,In_1983,In_1101);
nor U1899 (N_1899,In_889,In_1782);
nor U1900 (N_1900,In_1900,In_1600);
or U1901 (N_1901,In_266,In_269);
nand U1902 (N_1902,In_670,In_1908);
or U1903 (N_1903,In_1232,In_260);
and U1904 (N_1904,In_1068,In_485);
nand U1905 (N_1905,In_1951,In_757);
nand U1906 (N_1906,In_1812,In_1455);
nand U1907 (N_1907,In_1053,In_246);
nor U1908 (N_1908,In_174,In_1901);
xor U1909 (N_1909,In_569,In_751);
xor U1910 (N_1910,In_1862,In_1280);
and U1911 (N_1911,In_961,In_301);
or U1912 (N_1912,In_403,In_873);
and U1913 (N_1913,In_1399,In_808);
nand U1914 (N_1914,In_158,In_226);
and U1915 (N_1915,In_204,In_1075);
and U1916 (N_1916,In_1299,In_843);
nand U1917 (N_1917,In_1664,In_430);
nand U1918 (N_1918,In_1518,In_416);
nor U1919 (N_1919,In_1455,In_952);
or U1920 (N_1920,In_1034,In_732);
or U1921 (N_1921,In_1858,In_1860);
and U1922 (N_1922,In_1114,In_271);
or U1923 (N_1923,In_1556,In_817);
xnor U1924 (N_1924,In_1121,In_475);
and U1925 (N_1925,In_1473,In_1613);
nor U1926 (N_1926,In_266,In_880);
or U1927 (N_1927,In_598,In_1575);
nand U1928 (N_1928,In_1922,In_1136);
xnor U1929 (N_1929,In_855,In_886);
nor U1930 (N_1930,In_43,In_465);
nand U1931 (N_1931,In_1103,In_440);
xnor U1932 (N_1932,In_350,In_953);
or U1933 (N_1933,In_1282,In_617);
xnor U1934 (N_1934,In_1379,In_1210);
xnor U1935 (N_1935,In_1513,In_1638);
xor U1936 (N_1936,In_201,In_1808);
and U1937 (N_1937,In_126,In_550);
or U1938 (N_1938,In_567,In_875);
nand U1939 (N_1939,In_1968,In_1026);
nor U1940 (N_1940,In_871,In_1700);
or U1941 (N_1941,In_1924,In_1251);
nand U1942 (N_1942,In_1720,In_1245);
or U1943 (N_1943,In_1307,In_1437);
and U1944 (N_1944,In_1879,In_174);
and U1945 (N_1945,In_1637,In_1122);
nor U1946 (N_1946,In_1211,In_1428);
nor U1947 (N_1947,In_1683,In_630);
or U1948 (N_1948,In_1402,In_1985);
nand U1949 (N_1949,In_379,In_1206);
nand U1950 (N_1950,In_571,In_1515);
and U1951 (N_1951,In_1401,In_1793);
or U1952 (N_1952,In_572,In_371);
and U1953 (N_1953,In_866,In_1302);
or U1954 (N_1954,In_826,In_574);
and U1955 (N_1955,In_1580,In_1831);
and U1956 (N_1956,In_270,In_605);
nor U1957 (N_1957,In_1469,In_158);
nor U1958 (N_1958,In_59,In_120);
or U1959 (N_1959,In_851,In_1814);
xor U1960 (N_1960,In_1190,In_588);
nor U1961 (N_1961,In_1151,In_122);
nand U1962 (N_1962,In_1321,In_300);
nor U1963 (N_1963,In_1051,In_1392);
nor U1964 (N_1964,In_1108,In_530);
or U1965 (N_1965,In_1062,In_630);
nor U1966 (N_1966,In_947,In_1614);
and U1967 (N_1967,In_623,In_497);
xnor U1968 (N_1968,In_116,In_1179);
or U1969 (N_1969,In_1747,In_685);
xor U1970 (N_1970,In_1013,In_1479);
nor U1971 (N_1971,In_1009,In_51);
nor U1972 (N_1972,In_1127,In_865);
nand U1973 (N_1973,In_577,In_1771);
or U1974 (N_1974,In_1272,In_401);
or U1975 (N_1975,In_505,In_548);
and U1976 (N_1976,In_1346,In_1936);
and U1977 (N_1977,In_406,In_429);
nor U1978 (N_1978,In_1487,In_1900);
or U1979 (N_1979,In_1603,In_508);
nor U1980 (N_1980,In_16,In_1844);
and U1981 (N_1981,In_1927,In_704);
xor U1982 (N_1982,In_1858,In_1722);
and U1983 (N_1983,In_1385,In_540);
and U1984 (N_1984,In_1257,In_480);
nand U1985 (N_1985,In_85,In_678);
or U1986 (N_1986,In_689,In_1995);
xnor U1987 (N_1987,In_1106,In_758);
or U1988 (N_1988,In_991,In_1544);
nand U1989 (N_1989,In_1347,In_1123);
and U1990 (N_1990,In_47,In_1627);
xnor U1991 (N_1991,In_1101,In_1329);
xnor U1992 (N_1992,In_1168,In_34);
or U1993 (N_1993,In_654,In_1724);
and U1994 (N_1994,In_479,In_1792);
nand U1995 (N_1995,In_1169,In_1684);
nor U1996 (N_1996,In_1242,In_1603);
nand U1997 (N_1997,In_1048,In_1243);
or U1998 (N_1998,In_292,In_1496);
and U1999 (N_1999,In_769,In_1976);
and U2000 (N_2000,N_1065,N_1846);
nand U2001 (N_2001,N_536,N_54);
nand U2002 (N_2002,N_1014,N_1140);
nor U2003 (N_2003,N_1521,N_79);
nor U2004 (N_2004,N_481,N_1571);
and U2005 (N_2005,N_1904,N_707);
nor U2006 (N_2006,N_459,N_1713);
xnor U2007 (N_2007,N_1733,N_268);
xor U2008 (N_2008,N_880,N_1730);
nor U2009 (N_2009,N_87,N_408);
nor U2010 (N_2010,N_1778,N_1418);
nor U2011 (N_2011,N_620,N_557);
xnor U2012 (N_2012,N_1731,N_1216);
and U2013 (N_2013,N_1799,N_1832);
nand U2014 (N_2014,N_864,N_1231);
xor U2015 (N_2015,N_1596,N_1035);
nand U2016 (N_2016,N_492,N_1732);
and U2017 (N_2017,N_920,N_611);
xor U2018 (N_2018,N_68,N_1136);
xnor U2019 (N_2019,N_43,N_285);
or U2020 (N_2020,N_1541,N_117);
nor U2021 (N_2021,N_271,N_1610);
nor U2022 (N_2022,N_593,N_961);
and U2023 (N_2023,N_1645,N_606);
nand U2024 (N_2024,N_99,N_899);
nand U2025 (N_2025,N_755,N_1743);
and U2026 (N_2026,N_155,N_433);
nand U2027 (N_2027,N_739,N_1700);
or U2028 (N_2028,N_1539,N_1289);
nor U2029 (N_2029,N_1634,N_113);
and U2030 (N_2030,N_512,N_1847);
or U2031 (N_2031,N_1725,N_1311);
or U2032 (N_2032,N_551,N_941);
and U2033 (N_2033,N_1083,N_347);
nand U2034 (N_2034,N_1457,N_998);
nand U2035 (N_2035,N_766,N_1511);
nor U2036 (N_2036,N_1456,N_1918);
and U2037 (N_2037,N_1785,N_1451);
nor U2038 (N_2038,N_817,N_1840);
and U2039 (N_2039,N_369,N_663);
nand U2040 (N_2040,N_1431,N_1007);
nor U2041 (N_2041,N_575,N_891);
nand U2042 (N_2042,N_748,N_49);
and U2043 (N_2043,N_44,N_1705);
nor U2044 (N_2044,N_795,N_80);
nand U2045 (N_2045,N_538,N_919);
xor U2046 (N_2046,N_737,N_178);
and U2047 (N_2047,N_1244,N_1678);
xnor U2048 (N_2048,N_576,N_1550);
nor U2049 (N_2049,N_1950,N_1404);
nand U2050 (N_2050,N_953,N_639);
nor U2051 (N_2051,N_1503,N_53);
and U2052 (N_2052,N_545,N_1393);
nor U2053 (N_2053,N_1240,N_283);
xnor U2054 (N_2054,N_1992,N_1218);
and U2055 (N_2055,N_570,N_1622);
nor U2056 (N_2056,N_406,N_958);
or U2057 (N_2057,N_236,N_111);
nor U2058 (N_2058,N_1419,N_1722);
nor U2059 (N_2059,N_1538,N_509);
nor U2060 (N_2060,N_995,N_1093);
nand U2061 (N_2061,N_1841,N_1894);
xor U2062 (N_2062,N_86,N_645);
nor U2063 (N_2063,N_1797,N_1814);
or U2064 (N_2064,N_287,N_1059);
nand U2065 (N_2065,N_222,N_1766);
or U2066 (N_2066,N_352,N_847);
nand U2067 (N_2067,N_187,N_373);
or U2068 (N_2068,N_1892,N_1500);
or U2069 (N_2069,N_371,N_1224);
and U2070 (N_2070,N_1761,N_1777);
nor U2071 (N_2071,N_705,N_982);
nor U2072 (N_2072,N_1756,N_384);
or U2073 (N_2073,N_344,N_1440);
nor U2074 (N_2074,N_1661,N_46);
nand U2075 (N_2075,N_1825,N_1251);
nand U2076 (N_2076,N_1718,N_4);
or U2077 (N_2077,N_813,N_1055);
and U2078 (N_2078,N_1721,N_1727);
or U2079 (N_2079,N_1046,N_587);
nand U2080 (N_2080,N_1577,N_490);
nand U2081 (N_2081,N_1480,N_1956);
and U2082 (N_2082,N_1837,N_225);
nor U2083 (N_2083,N_797,N_360);
or U2084 (N_2084,N_1542,N_330);
nor U2085 (N_2085,N_1303,N_1292);
nor U2086 (N_2086,N_853,N_1029);
and U2087 (N_2087,N_789,N_23);
nor U2088 (N_2088,N_984,N_463);
or U2089 (N_2089,N_1890,N_977);
nand U2090 (N_2090,N_269,N_124);
and U2091 (N_2091,N_1019,N_220);
and U2092 (N_2092,N_1986,N_1908);
nand U2093 (N_2093,N_134,N_1828);
and U2094 (N_2094,N_1822,N_912);
xor U2095 (N_2095,N_596,N_1675);
or U2096 (N_2096,N_807,N_1606);
nand U2097 (N_2097,N_708,N_359);
and U2098 (N_2098,N_260,N_416);
or U2099 (N_2099,N_729,N_978);
nand U2100 (N_2100,N_231,N_337);
nor U2101 (N_2101,N_1633,N_1482);
or U2102 (N_2102,N_962,N_427);
xor U2103 (N_2103,N_295,N_1214);
and U2104 (N_2104,N_1913,N_956);
or U2105 (N_2105,N_1448,N_1692);
nor U2106 (N_2106,N_1769,N_1242);
xor U2107 (N_2107,N_464,N_905);
or U2108 (N_2108,N_527,N_135);
and U2109 (N_2109,N_294,N_1217);
nand U2110 (N_2110,N_764,N_868);
nor U2111 (N_2111,N_1391,N_1219);
nor U2112 (N_2112,N_567,N_622);
nor U2113 (N_2113,N_598,N_379);
and U2114 (N_2114,N_1344,N_1208);
and U2115 (N_2115,N_1164,N_787);
nor U2116 (N_2116,N_1807,N_1209);
xnor U2117 (N_2117,N_417,N_655);
and U2118 (N_2118,N_153,N_1910);
nor U2119 (N_2119,N_722,N_1588);
nor U2120 (N_2120,N_1945,N_158);
nand U2121 (N_2121,N_1514,N_665);
or U2122 (N_2122,N_1599,N_1808);
xor U2123 (N_2123,N_1173,N_1408);
or U2124 (N_2124,N_1411,N_1656);
xor U2125 (N_2125,N_937,N_1651);
nor U2126 (N_2126,N_168,N_232);
nor U2127 (N_2127,N_1420,N_1210);
and U2128 (N_2128,N_1490,N_458);
and U2129 (N_2129,N_1954,N_215);
xnor U2130 (N_2130,N_1034,N_1868);
and U2131 (N_2131,N_1342,N_1259);
nor U2132 (N_2132,N_1008,N_848);
nor U2133 (N_2133,N_75,N_834);
xor U2134 (N_2134,N_89,N_1073);
xor U2135 (N_2135,N_671,N_1655);
or U2136 (N_2136,N_1470,N_1308);
nand U2137 (N_2137,N_1512,N_1698);
nor U2138 (N_2138,N_197,N_1994);
nand U2139 (N_2139,N_1466,N_1865);
or U2140 (N_2140,N_444,N_1637);
nand U2141 (N_2141,N_45,N_1193);
nand U2142 (N_2142,N_1189,N_323);
nand U2143 (N_2143,N_1158,N_858);
and U2144 (N_2144,N_873,N_116);
or U2145 (N_2145,N_1145,N_1340);
xnor U2146 (N_2146,N_181,N_1051);
nor U2147 (N_2147,N_480,N_1337);
or U2148 (N_2148,N_405,N_875);
or U2149 (N_2149,N_1669,N_1012);
nor U2150 (N_2150,N_1629,N_216);
nand U2151 (N_2151,N_1299,N_1575);
nand U2152 (N_2152,N_1003,N_223);
nand U2153 (N_2153,N_1013,N_1458);
and U2154 (N_2154,N_1206,N_1001);
or U2155 (N_2155,N_689,N_1737);
and U2156 (N_2156,N_1131,N_97);
nor U2157 (N_2157,N_1381,N_1476);
and U2158 (N_2158,N_652,N_282);
nor U2159 (N_2159,N_595,N_1567);
and U2160 (N_2160,N_940,N_241);
nand U2161 (N_2161,N_1703,N_142);
nor U2162 (N_2162,N_493,N_244);
or U2163 (N_2163,N_1177,N_1502);
nand U2164 (N_2164,N_456,N_469);
nand U2165 (N_2165,N_1943,N_846);
nor U2166 (N_2166,N_1818,N_291);
xor U2167 (N_2167,N_202,N_1366);
or U2168 (N_2168,N_1468,N_183);
and U2169 (N_2169,N_1343,N_1555);
nor U2170 (N_2170,N_1734,N_863);
nand U2171 (N_2171,N_1706,N_683);
and U2172 (N_2172,N_1615,N_1963);
nor U2173 (N_2173,N_255,N_788);
xor U2174 (N_2174,N_1863,N_447);
nand U2175 (N_2175,N_420,N_1617);
or U2176 (N_2176,N_1677,N_192);
nand U2177 (N_2177,N_1556,N_636);
and U2178 (N_2178,N_1642,N_1682);
or U2179 (N_2179,N_145,N_591);
or U2180 (N_2180,N_615,N_981);
or U2181 (N_2181,N_1009,N_1644);
nand U2182 (N_2182,N_1384,N_449);
and U2183 (N_2183,N_95,N_1017);
or U2184 (N_2184,N_1496,N_1223);
or U2185 (N_2185,N_630,N_1653);
nor U2186 (N_2186,N_270,N_1202);
xor U2187 (N_2187,N_165,N_637);
nand U2188 (N_2188,N_1222,N_1916);
or U2189 (N_2189,N_1478,N_1434);
xnor U2190 (N_2190,N_1043,N_1447);
or U2191 (N_2191,N_971,N_1228);
nand U2192 (N_2192,N_1198,N_1015);
nand U2193 (N_2193,N_1063,N_36);
and U2194 (N_2194,N_968,N_1400);
nand U2195 (N_2195,N_1834,N_346);
nor U2196 (N_2196,N_475,N_1033);
xor U2197 (N_2197,N_226,N_1562);
and U2198 (N_2198,N_1282,N_1365);
and U2199 (N_2199,N_980,N_1532);
nand U2200 (N_2200,N_586,N_1039);
or U2201 (N_2201,N_1300,N_108);
nor U2202 (N_2202,N_1385,N_1127);
nor U2203 (N_2203,N_1869,N_879);
nand U2204 (N_2204,N_1409,N_573);
and U2205 (N_2205,N_1776,N_874);
and U2206 (N_2206,N_992,N_1813);
and U2207 (N_2207,N_15,N_1711);
and U2208 (N_2208,N_1955,N_814);
xnor U2209 (N_2209,N_623,N_1752);
and U2210 (N_2210,N_1499,N_1979);
nand U2211 (N_2211,N_804,N_736);
or U2212 (N_2212,N_1339,N_628);
or U2213 (N_2213,N_468,N_1068);
xor U2214 (N_2214,N_1861,N_180);
nor U2215 (N_2215,N_778,N_72);
and U2216 (N_2216,N_1650,N_946);
and U2217 (N_2217,N_686,N_66);
nor U2218 (N_2218,N_421,N_1618);
nor U2219 (N_2219,N_1075,N_1267);
and U2220 (N_2220,N_1744,N_1041);
or U2221 (N_2221,N_1463,N_103);
and U2222 (N_2222,N_1229,N_1489);
nand U2223 (N_2223,N_299,N_203);
or U2224 (N_2224,N_1780,N_1114);
nand U2225 (N_2225,N_1423,N_1566);
nor U2226 (N_2226,N_343,N_391);
or U2227 (N_2227,N_1553,N_310);
xor U2228 (N_2228,N_718,N_965);
nand U2229 (N_2229,N_944,N_1460);
or U2230 (N_2230,N_74,N_1338);
or U2231 (N_2231,N_1554,N_1373);
nand U2232 (N_2232,N_775,N_699);
or U2233 (N_2233,N_1249,N_259);
and U2234 (N_2234,N_157,N_37);
and U2235 (N_2235,N_59,N_1739);
nand U2236 (N_2236,N_979,N_609);
nor U2237 (N_2237,N_497,N_543);
or U2238 (N_2238,N_1163,N_862);
or U2239 (N_2239,N_280,N_1623);
xnor U2240 (N_2240,N_466,N_311);
or U2241 (N_2241,N_1740,N_1302);
and U2242 (N_2242,N_1197,N_230);
and U2243 (N_2243,N_928,N_1268);
or U2244 (N_2244,N_467,N_1741);
nor U2245 (N_2245,N_1835,N_1475);
nand U2246 (N_2246,N_1849,N_1699);
and U2247 (N_2247,N_1269,N_1595);
nand U2248 (N_2248,N_1176,N_1380);
nand U2249 (N_2249,N_460,N_1875);
xor U2250 (N_2250,N_436,N_1695);
nand U2251 (N_2251,N_473,N_1167);
or U2252 (N_2252,N_913,N_893);
xnor U2253 (N_2253,N_1382,N_1704);
nand U2254 (N_2254,N_195,N_462);
or U2255 (N_2255,N_784,N_1611);
and U2256 (N_2256,N_1774,N_229);
or U2257 (N_2257,N_1827,N_289);
and U2258 (N_2258,N_1886,N_1931);
and U2259 (N_2259,N_9,N_1245);
and U2260 (N_2260,N_1836,N_1951);
nor U2261 (N_2261,N_350,N_1565);
or U2262 (N_2262,N_303,N_1446);
or U2263 (N_2263,N_762,N_824);
and U2264 (N_2264,N_1261,N_1771);
nor U2265 (N_2265,N_1791,N_1838);
or U2266 (N_2266,N_1234,N_1996);
or U2267 (N_2267,N_1345,N_18);
or U2268 (N_2268,N_1350,N_1966);
or U2269 (N_2269,N_592,N_1506);
nor U2270 (N_2270,N_810,N_1199);
and U2271 (N_2271,N_380,N_312);
nand U2272 (N_2272,N_274,N_1260);
or U2273 (N_2273,N_354,N_1831);
and U2274 (N_2274,N_1830,N_679);
and U2275 (N_2275,N_771,N_605);
and U2276 (N_2276,N_1759,N_809);
or U2277 (N_2277,N_94,N_1902);
or U2278 (N_2278,N_1125,N_743);
xnor U2279 (N_2279,N_1960,N_1281);
or U2280 (N_2280,N_934,N_518);
nor U2281 (N_2281,N_1270,N_1991);
xnor U2282 (N_2282,N_1369,N_1054);
and U2283 (N_2283,N_451,N_1154);
xnor U2284 (N_2284,N_329,N_1363);
xor U2285 (N_2285,N_658,N_1534);
nand U2286 (N_2286,N_1048,N_844);
nor U2287 (N_2287,N_1889,N_1414);
or U2288 (N_2288,N_1433,N_1246);
or U2289 (N_2289,N_1909,N_1082);
xor U2290 (N_2290,N_1984,N_1062);
nor U2291 (N_2291,N_1768,N_340);
or U2292 (N_2292,N_821,N_1250);
xnor U2293 (N_2293,N_148,N_811);
or U2294 (N_2294,N_991,N_1291);
nand U2295 (N_2295,N_477,N_1469);
nand U2296 (N_2296,N_1087,N_1148);
nand U2297 (N_2297,N_1885,N_594);
or U2298 (N_2298,N_1146,N_887);
or U2299 (N_2299,N_276,N_163);
nor U2300 (N_2300,N_878,N_564);
nor U2301 (N_2301,N_435,N_1124);
nand U2302 (N_2302,N_681,N_684);
nor U2303 (N_2303,N_796,N_935);
nor U2304 (N_2304,N_939,N_510);
nor U2305 (N_2305,N_1150,N_301);
nor U2306 (N_2306,N_262,N_479);
nor U2307 (N_2307,N_438,N_1795);
nand U2308 (N_2308,N_439,N_1265);
or U2309 (N_2309,N_1248,N_666);
nand U2310 (N_2310,N_1099,N_1848);
or U2311 (N_2311,N_989,N_1184);
xnor U2312 (N_2312,N_321,N_1974);
nand U2313 (N_2313,N_372,N_395);
nand U2314 (N_2314,N_305,N_732);
and U2315 (N_2315,N_1652,N_224);
and U2316 (N_2316,N_1067,N_1215);
and U2317 (N_2317,N_375,N_1279);
and U2318 (N_2318,N_948,N_106);
nand U2319 (N_2319,N_1137,N_1399);
nand U2320 (N_2320,N_572,N_1175);
and U2321 (N_2321,N_1111,N_254);
and U2322 (N_2322,N_1569,N_754);
and U2323 (N_2323,N_88,N_1115);
or U2324 (N_2324,N_40,N_1346);
or U2325 (N_2325,N_1295,N_1551);
and U2326 (N_2326,N_768,N_1044);
or U2327 (N_2327,N_643,N_1877);
xor U2328 (N_2328,N_67,N_151);
nor U2329 (N_2329,N_1120,N_1801);
nor U2330 (N_2330,N_1578,N_177);
and U2331 (N_2331,N_924,N_820);
nand U2332 (N_2332,N_1942,N_1389);
and U2333 (N_2333,N_1374,N_247);
and U2334 (N_2334,N_993,N_396);
and U2335 (N_2335,N_1870,N_1372);
nor U2336 (N_2336,N_1547,N_0);
nand U2337 (N_2337,N_136,N_98);
nand U2338 (N_2338,N_1335,N_942);
nand U2339 (N_2339,N_179,N_1570);
nand U2340 (N_2340,N_1712,N_1893);
nor U2341 (N_2341,N_1188,N_1856);
nor U2342 (N_2342,N_1917,N_901);
nor U2343 (N_2343,N_1050,N_1349);
nor U2344 (N_2344,N_1585,N_1221);
and U2345 (N_2345,N_752,N_676);
or U2346 (N_2346,N_1772,N_1928);
nand U2347 (N_2347,N_772,N_1680);
and U2348 (N_2348,N_922,N_550);
nor U2349 (N_2349,N_1762,N_1604);
and U2350 (N_2350,N_1442,N_1920);
nand U2351 (N_2351,N_1192,N_751);
or U2352 (N_2352,N_50,N_32);
or U2353 (N_2353,N_526,N_668);
and U2354 (N_2354,N_1804,N_761);
nor U2355 (N_2355,N_240,N_1921);
nor U2356 (N_2356,N_955,N_246);
or U2357 (N_2357,N_414,N_1058);
and U2358 (N_2358,N_348,N_1781);
or U2359 (N_2359,N_399,N_1313);
and U2360 (N_2360,N_530,N_1388);
nor U2361 (N_2361,N_1540,N_1959);
nand U2362 (N_2362,N_185,N_1488);
nor U2363 (N_2363,N_1763,N_1283);
xnor U2364 (N_2364,N_1590,N_234);
and U2365 (N_2365,N_281,N_670);
nor U2366 (N_2366,N_1481,N_1395);
and U2367 (N_2367,N_1648,N_1226);
nor U2368 (N_2368,N_520,N_769);
or U2369 (N_2369,N_1392,N_217);
or U2370 (N_2370,N_507,N_1810);
or U2371 (N_2371,N_799,N_963);
xor U2372 (N_2372,N_132,N_140);
nand U2373 (N_2373,N_1907,N_1182);
nand U2374 (N_2374,N_1211,N_917);
and U2375 (N_2375,N_1662,N_1980);
or U2376 (N_2376,N_970,N_618);
xor U2377 (N_2377,N_1888,N_489);
xnor U2378 (N_2378,N_10,N_1508);
and U2379 (N_2379,N_191,N_383);
nor U2380 (N_2380,N_1205,N_1518);
or U2381 (N_2381,N_904,N_1694);
nand U2382 (N_2382,N_82,N_1627);
nor U2383 (N_2383,N_1647,N_1845);
xor U2384 (N_2384,N_1510,N_1826);
xor U2385 (N_2385,N_1563,N_1201);
or U2386 (N_2386,N_851,N_1715);
or U2387 (N_2387,N_983,N_688);
and U2388 (N_2388,N_313,N_1608);
nor U2389 (N_2389,N_73,N_1074);
nand U2390 (N_2390,N_1903,N_629);
nor U2391 (N_2391,N_890,N_1495);
nand U2392 (N_2392,N_1753,N_1084);
nand U2393 (N_2393,N_1095,N_1361);
xor U2394 (N_2394,N_1152,N_55);
nand U2395 (N_2395,N_63,N_500);
and U2396 (N_2396,N_713,N_818);
and U2397 (N_2397,N_58,N_1272);
nand U2398 (N_2398,N_1168,N_1277);
xnor U2399 (N_2399,N_672,N_1964);
nor U2400 (N_2400,N_675,N_1174);
nor U2401 (N_2401,N_13,N_125);
nor U2402 (N_2402,N_728,N_339);
or U2403 (N_2403,N_1842,N_62);
nor U2404 (N_2404,N_607,N_1276);
or U2405 (N_2405,N_1169,N_541);
nor U2406 (N_2406,N_1096,N_1533);
nor U2407 (N_2407,N_1207,N_910);
nand U2408 (N_2408,N_5,N_1794);
and U2409 (N_2409,N_1576,N_166);
nor U2410 (N_2410,N_1334,N_1066);
nand U2411 (N_2411,N_1351,N_1589);
xor U2412 (N_2412,N_1284,N_776);
or U2413 (N_2413,N_57,N_1898);
or U2414 (N_2414,N_701,N_1516);
nand U2415 (N_2415,N_1425,N_1657);
or U2416 (N_2416,N_1355,N_1787);
or U2417 (N_2417,N_1612,N_1760);
nor U2418 (N_2418,N_726,N_1674);
or U2419 (N_2419,N_1236,N_1410);
xnor U2420 (N_2420,N_506,N_382);
nand U2421 (N_2421,N_253,N_1757);
nor U2422 (N_2422,N_1993,N_1078);
nand U2423 (N_2423,N_1505,N_204);
or U2424 (N_2424,N_1587,N_1422);
nor U2425 (N_2425,N_1742,N_1758);
nor U2426 (N_2426,N_164,N_1052);
or U2427 (N_2427,N_733,N_700);
or U2428 (N_2428,N_388,N_763);
nor U2429 (N_2429,N_870,N_194);
and U2430 (N_2430,N_302,N_1056);
nand U2431 (N_2431,N_505,N_455);
nand U2432 (N_2432,N_1684,N_1574);
nand U2433 (N_2433,N_1190,N_214);
nand U2434 (N_2434,N_931,N_1047);
or U2435 (N_2435,N_1579,N_1110);
or U2436 (N_2436,N_1040,N_964);
or U2437 (N_2437,N_511,N_1415);
or U2438 (N_2438,N_249,N_119);
or U2439 (N_2439,N_1428,N_300);
or U2440 (N_2440,N_602,N_735);
and U2441 (N_2441,N_1926,N_1919);
and U2442 (N_2442,N_601,N_1278);
nor U2443 (N_2443,N_656,N_121);
nand U2444 (N_2444,N_780,N_865);
or U2445 (N_2445,N_267,N_1728);
nand U2446 (N_2446,N_365,N_740);
and U2447 (N_2447,N_883,N_1568);
nand U2448 (N_2448,N_84,N_1998);
nor U2449 (N_2449,N_419,N_20);
xnor U2450 (N_2450,N_1053,N_803);
or U2451 (N_2451,N_1360,N_1531);
nand U2452 (N_2452,N_1775,N_869);
and U2453 (N_2453,N_1784,N_1104);
nand U2454 (N_2454,N_1851,N_1736);
or U2455 (N_2455,N_1767,N_1027);
and U2456 (N_2456,N_886,N_207);
and U2457 (N_2457,N_1630,N_1997);
or U2458 (N_2458,N_1583,N_721);
xnor U2459 (N_2459,N_1329,N_734);
and U2460 (N_2460,N_1091,N_76);
nor U2461 (N_2461,N_146,N_614);
xnor U2462 (N_2462,N_988,N_664);
or U2463 (N_2463,N_1187,N_1620);
or U2464 (N_2464,N_1421,N_1517);
nand U2465 (N_2465,N_1564,N_1367);
nand U2466 (N_2466,N_1022,N_1726);
nor U2467 (N_2467,N_687,N_51);
or U2468 (N_2468,N_1319,N_680);
or U2469 (N_2469,N_1635,N_1679);
and U2470 (N_2470,N_1935,N_1132);
nand U2471 (N_2471,N_1988,N_517);
nand U2472 (N_2472,N_533,N_1643);
xor U2473 (N_2473,N_115,N_422);
and U2474 (N_2474,N_1179,N_402);
nor U2475 (N_2475,N_193,N_425);
or U2476 (N_2476,N_1196,N_1624);
nand U2477 (N_2477,N_266,N_428);
nor U2478 (N_2478,N_364,N_513);
and U2479 (N_2479,N_159,N_29);
or U2480 (N_2480,N_83,N_716);
and U2481 (N_2481,N_25,N_1107);
nor U2482 (N_2482,N_1445,N_105);
and U2483 (N_2483,N_1754,N_173);
nor U2484 (N_2484,N_653,N_1376);
or U2485 (N_2485,N_897,N_1631);
and U2486 (N_2486,N_1371,N_565);
xnor U2487 (N_2487,N_1560,N_1549);
xnor U2488 (N_2488,N_635,N_172);
nor U2489 (N_2489,N_141,N_1280);
or U2490 (N_2490,N_725,N_1341);
xnor U2491 (N_2491,N_322,N_829);
or U2492 (N_2492,N_1454,N_800);
or U2493 (N_2493,N_997,N_902);
xor U2494 (N_2494,N_1764,N_1332);
xnor U2495 (N_2495,N_104,N_1304);
or U2496 (N_2496,N_1850,N_109);
or U2497 (N_2497,N_1707,N_275);
xnor U2498 (N_2498,N_860,N_288);
and U2499 (N_2499,N_196,N_650);
nand U2500 (N_2500,N_1326,N_26);
and U2501 (N_2501,N_338,N_1815);
xnor U2502 (N_2502,N_1929,N_1852);
nand U2503 (N_2503,N_529,N_1320);
and U2504 (N_2504,N_608,N_660);
nand U2505 (N_2505,N_324,N_201);
and U2506 (N_2506,N_825,N_554);
and U2507 (N_2507,N_1939,N_1086);
nor U2508 (N_2508,N_1896,N_413);
nand U2509 (N_2509,N_437,N_1225);
nor U2510 (N_2510,N_358,N_1688);
and U2511 (N_2511,N_616,N_1501);
and U2512 (N_2512,N_1153,N_855);
xnor U2513 (N_2513,N_745,N_1681);
and U2514 (N_2514,N_926,N_1444);
nor U2515 (N_2515,N_1143,N_1824);
and U2516 (N_2516,N_1709,N_711);
nand U2517 (N_2517,N_638,N_461);
or U2518 (N_2518,N_1593,N_1429);
nor U2519 (N_2519,N_345,N_519);
and U2520 (N_2520,N_61,N_1812);
and U2521 (N_2521,N_952,N_457);
or U2522 (N_2522,N_1880,N_1435);
or U2523 (N_2523,N_1006,N_1605);
and U2524 (N_2524,N_1439,N_1786);
nor U2525 (N_2525,N_1081,N_1621);
or U2526 (N_2526,N_1362,N_452);
nor U2527 (N_2527,N_669,N_133);
and U2528 (N_2528,N_1461,N_1537);
and U2529 (N_2529,N_1368,N_1230);
and U2530 (N_2530,N_138,N_1665);
and U2531 (N_2531,N_884,N_1394);
nor U2532 (N_2532,N_1853,N_1079);
nor U2533 (N_2533,N_574,N_1978);
or U2534 (N_2534,N_102,N_1755);
nand U2535 (N_2535,N_333,N_484);
or U2536 (N_2536,N_1,N_758);
nor U2537 (N_2537,N_1626,N_1181);
nand U2538 (N_2538,N_1171,N_1708);
nor U2539 (N_2539,N_1949,N_631);
and U2540 (N_2540,N_835,N_1690);
nand U2541 (N_2541,N_693,N_150);
and U2542 (N_2542,N_453,N_691);
nand U2543 (N_2543,N_1200,N_1985);
or U2544 (N_2544,N_1806,N_704);
xnor U2545 (N_2545,N_1862,N_1867);
nand U2546 (N_2546,N_128,N_827);
nor U2547 (N_2547,N_781,N_1166);
and U2548 (N_2548,N_198,N_22);
or U2549 (N_2549,N_186,N_805);
or U2550 (N_2550,N_1305,N_1887);
nor U2551 (N_2551,N_1103,N_328);
or U2552 (N_2552,N_233,N_41);
xnor U2553 (N_2553,N_767,N_843);
and U2554 (N_2554,N_1271,N_309);
or U2555 (N_2555,N_243,N_1162);
and U2556 (N_2556,N_1310,N_1948);
and U2557 (N_2557,N_1640,N_1462);
or U2558 (N_2558,N_659,N_1811);
nand U2559 (N_2559,N_1664,N_1745);
and U2560 (N_2560,N_315,N_514);
or U2561 (N_2561,N_1958,N_16);
and U2562 (N_2562,N_1738,N_112);
and U2563 (N_2563,N_1097,N_1356);
and U2564 (N_2564,N_378,N_1659);
nor U2565 (N_2565,N_1773,N_1407);
nor U2566 (N_2566,N_1529,N_833);
or U2567 (N_2567,N_251,N_1318);
nor U2568 (N_2568,N_1118,N_219);
nor U2569 (N_2569,N_1323,N_1873);
and U2570 (N_2570,N_1252,N_1010);
nand U2571 (N_2571,N_139,N_410);
nand U2572 (N_2572,N_1060,N_932);
and U2573 (N_2573,N_1976,N_1572);
and U2574 (N_2574,N_1881,N_1452);
and U2575 (N_2575,N_1693,N_757);
nand U2576 (N_2576,N_85,N_1089);
nor U2577 (N_2577,N_1287,N_566);
or U2578 (N_2578,N_694,N_892);
or U2579 (N_2579,N_731,N_296);
nand U2580 (N_2580,N_1536,N_1802);
and U2581 (N_2581,N_1879,N_1293);
nor U2582 (N_2582,N_1241,N_885);
or U2583 (N_2583,N_1546,N_152);
and U2584 (N_2584,N_888,N_1874);
nand U2585 (N_2585,N_1038,N_866);
nand U2586 (N_2586,N_1649,N_1748);
or U2587 (N_2587,N_261,N_1616);
or U2588 (N_2588,N_1735,N_258);
or U2589 (N_2589,N_1030,N_92);
or U2590 (N_2590,N_1878,N_1983);
nor U2591 (N_2591,N_1872,N_1491);
nor U2592 (N_2592,N_1525,N_854);
and U2593 (N_2593,N_923,N_1936);
nor U2594 (N_2594,N_747,N_28);
and U2595 (N_2595,N_1782,N_548);
or U2596 (N_2596,N_1037,N_353);
or U2597 (N_2597,N_1559,N_1906);
nand U2598 (N_2598,N_1403,N_882);
xor U2599 (N_2599,N_1307,N_411);
or U2600 (N_2600,N_823,N_320);
or U2601 (N_2601,N_130,N_1203);
xor U2602 (N_2602,N_1405,N_1032);
nor U2603 (N_2603,N_1558,N_856);
xor U2604 (N_2604,N_644,N_727);
nand U2605 (N_2605,N_1891,N_278);
nor U2606 (N_2606,N_1069,N_1584);
and U2607 (N_2607,N_496,N_1416);
nor U2608 (N_2608,N_326,N_107);
or U2609 (N_2609,N_528,N_429);
or U2610 (N_2610,N_619,N_1306);
nand U2611 (N_2611,N_966,N_969);
or U2612 (N_2612,N_1328,N_17);
nor U2613 (N_2613,N_936,N_70);
or U2614 (N_2614,N_1884,N_426);
nand U2615 (N_2615,N_756,N_387);
nand U2616 (N_2616,N_206,N_389);
nand U2617 (N_2617,N_1600,N_710);
and U2618 (N_2618,N_1005,N_617);
nand U2619 (N_2619,N_1938,N_1258);
or U2620 (N_2620,N_624,N_100);
or U2621 (N_2621,N_960,N_1800);
and U2622 (N_2622,N_730,N_1232);
nor U2623 (N_2623,N_625,N_508);
nand U2624 (N_2624,N_621,N_1934);
nor U2625 (N_2625,N_1513,N_1535);
nor U2626 (N_2626,N_849,N_1297);
nand U2627 (N_2627,N_290,N_286);
nand U2628 (N_2628,N_1264,N_200);
nand U2629 (N_2629,N_719,N_175);
nand U2630 (N_2630,N_33,N_317);
or U2631 (N_2631,N_1121,N_1417);
or U2632 (N_2632,N_1031,N_1286);
and U2633 (N_2633,N_1602,N_357);
or U2634 (N_2634,N_1126,N_832);
nor U2635 (N_2635,N_678,N_392);
and U2636 (N_2636,N_1788,N_867);
or U2637 (N_2637,N_1018,N_65);
and U2638 (N_2638,N_184,N_600);
nor U2639 (N_2639,N_171,N_1975);
nor U2640 (N_2640,N_1161,N_1170);
nor U2641 (N_2641,N_627,N_1178);
nand U2642 (N_2642,N_1628,N_842);
nor U2643 (N_2643,N_819,N_483);
nor U2644 (N_2644,N_199,N_1839);
or U2645 (N_2645,N_1235,N_1493);
or U2646 (N_2646,N_48,N_443);
nor U2647 (N_2647,N_950,N_1843);
nand U2648 (N_2648,N_1426,N_356);
nor U2649 (N_2649,N_503,N_442);
xnor U2650 (N_2650,N_987,N_1509);
nand U2651 (N_2651,N_1352,N_1357);
or U2652 (N_2652,N_1274,N_1940);
nor U2653 (N_2653,N_539,N_850);
and U2654 (N_2654,N_999,N_1315);
or U2655 (N_2655,N_404,N_838);
and U2656 (N_2656,N_1070,N_1450);
or U2657 (N_2657,N_703,N_1147);
and U2658 (N_2658,N_1749,N_12);
nor U2659 (N_2659,N_1061,N_96);
or U2660 (N_2660,N_515,N_502);
or U2661 (N_2661,N_1504,N_568);
nor U2662 (N_2662,N_717,N_21);
nor U2663 (N_2663,N_1922,N_1437);
nand U2664 (N_2664,N_1961,N_555);
or U2665 (N_2665,N_114,N_450);
nand U2666 (N_2666,N_1798,N_532);
or U2667 (N_2667,N_1901,N_898);
and U2668 (N_2668,N_1676,N_957);
and U2669 (N_2669,N_1683,N_1607);
and U2670 (N_2670,N_238,N_504);
nor U2671 (N_2671,N_34,N_1347);
nand U2672 (N_2672,N_1750,N_368);
and U2673 (N_2673,N_279,N_1438);
or U2674 (N_2674,N_1666,N_1882);
or U2675 (N_2675,N_633,N_1947);
xnor U2676 (N_2676,N_1322,N_1112);
and U2677 (N_2677,N_1497,N_552);
nand U2678 (N_2678,N_1545,N_1479);
or U2679 (N_2679,N_1858,N_610);
or U2680 (N_2680,N_1965,N_1185);
nand U2681 (N_2681,N_908,N_1582);
and U2682 (N_2682,N_1144,N_110);
and U2683 (N_2683,N_1101,N_1494);
and U2684 (N_2684,N_38,N_448);
nand U2685 (N_2685,N_1524,N_894);
and U2686 (N_2686,N_690,N_39);
nor U2687 (N_2687,N_839,N_553);
or U2688 (N_2688,N_582,N_648);
nand U2689 (N_2689,N_256,N_1336);
or U2690 (N_2690,N_1139,N_91);
xnor U2691 (N_2691,N_1573,N_1905);
and U2692 (N_2692,N_1317,N_581);
nor U2693 (N_2693,N_974,N_1989);
nor U2694 (N_2694,N_972,N_162);
and U2695 (N_2695,N_218,N_1911);
or U2696 (N_2696,N_273,N_167);
and U2697 (N_2697,N_1660,N_959);
xor U2698 (N_2698,N_42,N_488);
nand U2699 (N_2699,N_1156,N_129);
nor U2700 (N_2700,N_264,N_1119);
nor U2701 (N_2701,N_1932,N_1990);
nand U2702 (N_2702,N_685,N_1724);
or U2703 (N_2703,N_182,N_1386);
nand U2704 (N_2704,N_316,N_8);
nor U2705 (N_2705,N_590,N_741);
or U2706 (N_2706,N_1673,N_1544);
nor U2707 (N_2707,N_516,N_188);
or U2708 (N_2708,N_304,N_871);
or U2709 (N_2709,N_714,N_1263);
or U2710 (N_2710,N_1135,N_90);
xor U2711 (N_2711,N_1614,N_996);
or U2712 (N_2712,N_24,N_682);
or U2713 (N_2713,N_81,N_1011);
nand U2714 (N_2714,N_1117,N_1746);
or U2715 (N_2715,N_753,N_945);
or U2716 (N_2716,N_1519,N_1301);
or U2717 (N_2717,N_1995,N_603);
and U2718 (N_2718,N_1876,N_1819);
and U2719 (N_2719,N_69,N_535);
nor U2720 (N_2720,N_1233,N_546);
nor U2721 (N_2721,N_634,N_361);
and U2722 (N_2722,N_1378,N_1256);
nand U2723 (N_2723,N_1719,N_1520);
or U2724 (N_2724,N_1255,N_852);
or U2725 (N_2725,N_524,N_1100);
nor U2726 (N_2726,N_808,N_1923);
nand U2727 (N_2727,N_990,N_930);
nor U2728 (N_2728,N_826,N_744);
and U2729 (N_2729,N_1023,N_1330);
or U2730 (N_2730,N_1561,N_1254);
or U2731 (N_2731,N_1441,N_292);
and U2732 (N_2732,N_889,N_1930);
nor U2733 (N_2733,N_1654,N_1102);
nand U2734 (N_2734,N_1639,N_6);
nand U2735 (N_2735,N_1390,N_1625);
and U2736 (N_2736,N_470,N_1160);
nor U2737 (N_2737,N_1820,N_558);
and U2738 (N_2738,N_706,N_872);
or U2739 (N_2739,N_1036,N_1129);
or U2740 (N_2740,N_1977,N_1092);
or U2741 (N_2741,N_78,N_1432);
and U2742 (N_2742,N_351,N_1116);
nor U2743 (N_2743,N_1142,N_632);
nand U2744 (N_2744,N_1090,N_1973);
and U2745 (N_2745,N_308,N_792);
nand U2746 (N_2746,N_363,N_738);
nand U2747 (N_2747,N_985,N_1899);
or U2748 (N_2748,N_1485,N_877);
or U2749 (N_2749,N_580,N_1298);
or U2750 (N_2750,N_1672,N_245);
nand U2751 (N_2751,N_859,N_544);
nand U2752 (N_2752,N_393,N_697);
or U2753 (N_2753,N_715,N_1696);
nand U2754 (N_2754,N_161,N_355);
nand U2755 (N_2755,N_212,N_349);
and U2756 (N_2756,N_126,N_1646);
nand U2757 (N_2757,N_1702,N_794);
or U2758 (N_2758,N_1912,N_646);
nand U2759 (N_2759,N_1717,N_802);
or U2760 (N_2760,N_336,N_1883);
nor U2761 (N_2761,N_1866,N_390);
xor U2762 (N_2762,N_816,N_56);
nor U2763 (N_2763,N_709,N_1609);
nand U2764 (N_2764,N_465,N_954);
or U2765 (N_2765,N_975,N_1829);
and U2766 (N_2766,N_332,N_583);
nand U2767 (N_2767,N_1854,N_418);
or U2768 (N_2768,N_973,N_1296);
nor U2769 (N_2769,N_642,N_1915);
or U2770 (N_2770,N_837,N_487);
and U2771 (N_2771,N_1453,N_1379);
nor U2772 (N_2772,N_933,N_209);
and U2773 (N_2773,N_250,N_1805);
or U2774 (N_2774,N_1714,N_876);
nor U2775 (N_2775,N_495,N_1191);
or U2776 (N_2776,N_1598,N_647);
nand U2777 (N_2777,N_169,N_64);
xnor U2778 (N_2778,N_1860,N_446);
nor U2779 (N_2779,N_1237,N_1071);
and U2780 (N_2780,N_1028,N_377);
nor U2781 (N_2781,N_1937,N_2);
nor U2782 (N_2782,N_588,N_770);
and U2783 (N_2783,N_160,N_131);
or U2784 (N_2784,N_1982,N_1527);
or U2785 (N_2785,N_1424,N_1333);
and U2786 (N_2786,N_423,N_298);
nor U2787 (N_2787,N_1927,N_190);
or U2788 (N_2788,N_1253,N_812);
or U2789 (N_2789,N_7,N_1671);
and U2790 (N_2790,N_248,N_815);
nor U2791 (N_2791,N_916,N_1944);
and U2792 (N_2792,N_1094,N_476);
and U2793 (N_2793,N_774,N_1720);
nand U2794 (N_2794,N_841,N_749);
nor U2795 (N_2795,N_549,N_1855);
nor U2796 (N_2796,N_571,N_651);
nor U2797 (N_2797,N_921,N_1472);
nand U2798 (N_2798,N_314,N_696);
nor U2799 (N_2799,N_1823,N_35);
nor U2800 (N_2800,N_398,N_1464);
nand U2801 (N_2801,N_1523,N_1412);
and U2802 (N_2802,N_1859,N_242);
nor U2803 (N_2803,N_1632,N_1548);
xor U2804 (N_2804,N_857,N_1186);
nor U2805 (N_2805,N_1377,N_1970);
and U2806 (N_2806,N_906,N_929);
or U2807 (N_2807,N_1498,N_1406);
and U2808 (N_2808,N_1275,N_1227);
and U2809 (N_2809,N_208,N_1796);
nor U2810 (N_2810,N_491,N_677);
and U2811 (N_2811,N_143,N_793);
xnor U2812 (N_2812,N_522,N_1603);
nand U2813 (N_2813,N_1021,N_407);
and U2814 (N_2814,N_1592,N_370);
or U2815 (N_2815,N_1436,N_235);
or U2816 (N_2816,N_1586,N_445);
or U2817 (N_2817,N_559,N_1941);
nand U2818 (N_2818,N_221,N_1109);
or U2819 (N_2819,N_1358,N_1077);
or U2820 (N_2820,N_19,N_1157);
or U2821 (N_2821,N_434,N_1401);
or U2822 (N_2822,N_93,N_1792);
nand U2823 (N_2823,N_1601,N_1864);
or U2824 (N_2824,N_77,N_123);
and U2825 (N_2825,N_692,N_1397);
nand U2826 (N_2826,N_903,N_252);
nor U2827 (N_2827,N_938,N_474);
and U2828 (N_2828,N_1266,N_263);
nand U2829 (N_2829,N_1141,N_144);
nor U2830 (N_2830,N_569,N_1262);
xnor U2831 (N_2831,N_1402,N_1816);
and U2832 (N_2832,N_765,N_1971);
and U2833 (N_2833,N_213,N_472);
and U2834 (N_2834,N_1024,N_1933);
or U2835 (N_2835,N_1486,N_1465);
nor U2836 (N_2836,N_649,N_584);
nor U2837 (N_2837,N_562,N_1528);
and U2838 (N_2838,N_547,N_1165);
and U2839 (N_2839,N_60,N_1353);
nand U2840 (N_2840,N_537,N_374);
and U2841 (N_2841,N_911,N_1900);
nor U2842 (N_2842,N_1833,N_1790);
and U2843 (N_2843,N_1686,N_1076);
nor U2844 (N_2844,N_498,N_1515);
or U2845 (N_2845,N_1999,N_454);
nand U2846 (N_2846,N_318,N_1449);
and U2847 (N_2847,N_1106,N_915);
or U2848 (N_2848,N_1467,N_1314);
or U2849 (N_2849,N_1133,N_1149);
or U2850 (N_2850,N_1594,N_394);
or U2851 (N_2851,N_556,N_1016);
and U2852 (N_2852,N_401,N_1619);
xor U2853 (N_2853,N_1312,N_385);
nor U2854 (N_2854,N_147,N_440);
and U2855 (N_2855,N_798,N_1370);
or U2856 (N_2856,N_1691,N_1924);
and U2857 (N_2857,N_1507,N_599);
nor U2858 (N_2858,N_712,N_1247);
nand U2859 (N_2859,N_1020,N_896);
and U2860 (N_2860,N_1552,N_667);
or U2861 (N_2861,N_1324,N_779);
nor U2862 (N_2862,N_1105,N_521);
nor U2863 (N_2863,N_1747,N_585);
and U2864 (N_2864,N_1526,N_1953);
and U2865 (N_2865,N_1471,N_327);
nor U2866 (N_2866,N_156,N_1897);
or U2867 (N_2867,N_783,N_1793);
nor U2868 (N_2868,N_1969,N_881);
nand U2869 (N_2869,N_412,N_1484);
or U2870 (N_2870,N_331,N_1723);
nand U2871 (N_2871,N_1238,N_265);
xor U2872 (N_2872,N_1383,N_1914);
nor U2873 (N_2873,N_746,N_1770);
nand U2874 (N_2874,N_1159,N_482);
nor U2875 (N_2875,N_612,N_1779);
nand U2876 (N_2876,N_52,N_1668);
or U2877 (N_2877,N_205,N_1670);
nor U2878 (N_2878,N_1857,N_210);
nor U2879 (N_2879,N_773,N_947);
nand U2880 (N_2880,N_801,N_1080);
nand U2881 (N_2881,N_1088,N_1729);
nor U2882 (N_2882,N_319,N_1844);
nor U2883 (N_2883,N_367,N_579);
or U2884 (N_2884,N_1821,N_1473);
nor U2885 (N_2885,N_1113,N_560);
or U2886 (N_2886,N_626,N_1387);
or U2887 (N_2887,N_1398,N_272);
nand U2888 (N_2888,N_1492,N_228);
nor U2889 (N_2889,N_1331,N_1273);
or U2890 (N_2890,N_831,N_1183);
or U2891 (N_2891,N_907,N_1477);
nand U2892 (N_2892,N_1687,N_189);
nand U2893 (N_2893,N_409,N_499);
and U2894 (N_2894,N_1765,N_1128);
nand U2895 (N_2895,N_1957,N_1213);
xnor U2896 (N_2896,N_830,N_1239);
xnor U2897 (N_2897,N_1689,N_1925);
and U2898 (N_2898,N_967,N_828);
nor U2899 (N_2899,N_1180,N_1288);
and U2900 (N_2900,N_1557,N_657);
or U2901 (N_2901,N_673,N_257);
nand U2902 (N_2902,N_1026,N_1613);
or U2903 (N_2903,N_531,N_297);
xor U2904 (N_2904,N_698,N_1172);
or U2905 (N_2905,N_1597,N_1697);
or U2906 (N_2906,N_1783,N_1327);
nand U2907 (N_2907,N_1981,N_1895);
nor U2908 (N_2908,N_471,N_1000);
nor U2909 (N_2909,N_478,N_293);
nor U2910 (N_2910,N_641,N_661);
and U2911 (N_2911,N_170,N_1580);
nand U2912 (N_2912,N_1045,N_307);
xnor U2913 (N_2913,N_1427,N_840);
nand U2914 (N_2914,N_1430,N_122);
xnor U2915 (N_2915,N_561,N_1359);
or U2916 (N_2916,N_1123,N_334);
nor U2917 (N_2917,N_895,N_1321);
and U2918 (N_2918,N_1658,N_1004);
nand U2919 (N_2919,N_1751,N_1522);
or U2920 (N_2920,N_1946,N_604);
nor U2921 (N_2921,N_1290,N_27);
nand U2922 (N_2922,N_30,N_534);
and U2923 (N_2923,N_441,N_430);
and U2924 (N_2924,N_1638,N_1716);
and U2925 (N_2925,N_542,N_578);
nor U2926 (N_2926,N_501,N_494);
and U2927 (N_2927,N_14,N_341);
nor U2928 (N_2928,N_1325,N_1871);
nand U2929 (N_2929,N_325,N_986);
or U2930 (N_2930,N_211,N_154);
or U2931 (N_2931,N_1049,N_662);
or U2932 (N_2932,N_759,N_1396);
nand U2933 (N_2933,N_47,N_1002);
or U2934 (N_2934,N_1701,N_1967);
nor U2935 (N_2935,N_486,N_1212);
xnor U2936 (N_2936,N_523,N_927);
and U2937 (N_2937,N_1220,N_1122);
nand U2938 (N_2938,N_1487,N_11);
and U2939 (N_2939,N_577,N_1243);
nand U2940 (N_2940,N_376,N_1025);
and U2941 (N_2941,N_400,N_640);
nand U2942 (N_2942,N_1064,N_836);
nand U2943 (N_2943,N_951,N_174);
and U2944 (N_2944,N_1530,N_1130);
or U2945 (N_2945,N_239,N_176);
and U2946 (N_2946,N_1072,N_540);
nand U2947 (N_2947,N_597,N_403);
or U2948 (N_2948,N_1348,N_1042);
and U2949 (N_2949,N_3,N_1098);
and U2950 (N_2950,N_563,N_1667);
nor U2951 (N_2951,N_806,N_120);
nor U2952 (N_2952,N_397,N_485);
nor U2953 (N_2953,N_777,N_1483);
nand U2954 (N_2954,N_1294,N_284);
or U2955 (N_2955,N_720,N_674);
or U2956 (N_2956,N_1155,N_1809);
and U2957 (N_2957,N_1636,N_1285);
nand U2958 (N_2958,N_386,N_750);
and U2959 (N_2959,N_976,N_1459);
or U2960 (N_2960,N_760,N_1968);
nor U2961 (N_2961,N_1663,N_1455);
nand U2962 (N_2962,N_1591,N_277);
nor U2963 (N_2963,N_1194,N_362);
nor U2964 (N_2964,N_342,N_1710);
nand U2965 (N_2965,N_127,N_1443);
nand U2966 (N_2966,N_1195,N_742);
xor U2967 (N_2967,N_1474,N_782);
nand U2968 (N_2968,N_31,N_1134);
nand U2969 (N_2969,N_791,N_702);
nor U2970 (N_2970,N_1108,N_137);
nand U2971 (N_2971,N_943,N_1543);
nor U2972 (N_2972,N_1354,N_589);
nand U2973 (N_2973,N_1257,N_525);
nand U2974 (N_2974,N_1204,N_1685);
nand U2975 (N_2975,N_1972,N_1803);
and U2976 (N_2976,N_431,N_306);
xor U2977 (N_2977,N_918,N_822);
or U2978 (N_2978,N_1375,N_994);
and U2979 (N_2979,N_1581,N_1817);
nand U2980 (N_2980,N_335,N_1085);
and U2981 (N_2981,N_366,N_724);
or U2982 (N_2982,N_1138,N_1413);
or U2983 (N_2983,N_1151,N_237);
nor U2984 (N_2984,N_415,N_1952);
nor U2985 (N_2985,N_71,N_227);
or U2986 (N_2986,N_925,N_900);
and U2987 (N_2987,N_101,N_845);
nor U2988 (N_2988,N_1364,N_914);
xnor U2989 (N_2989,N_786,N_909);
nor U2990 (N_2990,N_1309,N_432);
and U2991 (N_2991,N_1962,N_785);
and U2992 (N_2992,N_381,N_118);
nand U2993 (N_2993,N_1316,N_790);
nor U2994 (N_2994,N_654,N_1789);
nand U2995 (N_2995,N_1641,N_949);
nand U2996 (N_2996,N_695,N_861);
or U2997 (N_2997,N_149,N_1987);
and U2998 (N_2998,N_424,N_613);
and U2999 (N_2999,N_723,N_1057);
nand U3000 (N_3000,N_1687,N_982);
nor U3001 (N_3001,N_742,N_1017);
or U3002 (N_3002,N_688,N_1306);
and U3003 (N_3003,N_1278,N_1064);
and U3004 (N_3004,N_1211,N_1095);
or U3005 (N_3005,N_1883,N_66);
and U3006 (N_3006,N_212,N_1828);
nand U3007 (N_3007,N_1163,N_1867);
and U3008 (N_3008,N_1395,N_1890);
and U3009 (N_3009,N_1997,N_618);
and U3010 (N_3010,N_961,N_1131);
and U3011 (N_3011,N_562,N_1030);
nor U3012 (N_3012,N_201,N_390);
and U3013 (N_3013,N_107,N_824);
nor U3014 (N_3014,N_252,N_206);
nor U3015 (N_3015,N_824,N_1112);
or U3016 (N_3016,N_178,N_170);
and U3017 (N_3017,N_103,N_429);
nor U3018 (N_3018,N_1257,N_1034);
nor U3019 (N_3019,N_934,N_1236);
and U3020 (N_3020,N_1539,N_354);
nor U3021 (N_3021,N_1485,N_620);
nor U3022 (N_3022,N_1306,N_772);
or U3023 (N_3023,N_1204,N_598);
xor U3024 (N_3024,N_1481,N_1695);
xor U3025 (N_3025,N_192,N_438);
nor U3026 (N_3026,N_743,N_1897);
nand U3027 (N_3027,N_1452,N_898);
and U3028 (N_3028,N_407,N_260);
or U3029 (N_3029,N_1957,N_1472);
or U3030 (N_3030,N_469,N_561);
and U3031 (N_3031,N_1802,N_548);
nand U3032 (N_3032,N_364,N_1426);
nand U3033 (N_3033,N_1629,N_1836);
and U3034 (N_3034,N_1473,N_1158);
xor U3035 (N_3035,N_2,N_1926);
and U3036 (N_3036,N_377,N_809);
nand U3037 (N_3037,N_1004,N_969);
and U3038 (N_3038,N_451,N_120);
and U3039 (N_3039,N_1159,N_1635);
nor U3040 (N_3040,N_59,N_1795);
nand U3041 (N_3041,N_1392,N_1396);
nor U3042 (N_3042,N_1527,N_1517);
or U3043 (N_3043,N_554,N_584);
and U3044 (N_3044,N_1372,N_164);
nand U3045 (N_3045,N_1476,N_924);
nor U3046 (N_3046,N_1185,N_1861);
nand U3047 (N_3047,N_1050,N_320);
nand U3048 (N_3048,N_1698,N_1212);
or U3049 (N_3049,N_841,N_1177);
and U3050 (N_3050,N_1578,N_738);
xnor U3051 (N_3051,N_1109,N_415);
and U3052 (N_3052,N_99,N_339);
nor U3053 (N_3053,N_1606,N_1676);
and U3054 (N_3054,N_1371,N_1504);
and U3055 (N_3055,N_979,N_1985);
nor U3056 (N_3056,N_752,N_969);
nor U3057 (N_3057,N_1869,N_937);
nor U3058 (N_3058,N_1789,N_1521);
nor U3059 (N_3059,N_877,N_684);
xor U3060 (N_3060,N_998,N_1264);
and U3061 (N_3061,N_1692,N_1521);
nor U3062 (N_3062,N_349,N_435);
nor U3063 (N_3063,N_1493,N_288);
and U3064 (N_3064,N_745,N_1460);
nand U3065 (N_3065,N_1678,N_560);
nor U3066 (N_3066,N_1140,N_1055);
or U3067 (N_3067,N_1468,N_1595);
or U3068 (N_3068,N_845,N_991);
or U3069 (N_3069,N_765,N_798);
nor U3070 (N_3070,N_383,N_404);
and U3071 (N_3071,N_859,N_993);
nor U3072 (N_3072,N_537,N_1856);
nor U3073 (N_3073,N_1644,N_429);
nor U3074 (N_3074,N_681,N_384);
nand U3075 (N_3075,N_895,N_926);
or U3076 (N_3076,N_1262,N_1504);
nor U3077 (N_3077,N_120,N_98);
nand U3078 (N_3078,N_771,N_942);
xor U3079 (N_3079,N_1181,N_257);
nor U3080 (N_3080,N_1708,N_190);
and U3081 (N_3081,N_1111,N_1435);
nand U3082 (N_3082,N_265,N_191);
and U3083 (N_3083,N_909,N_775);
nand U3084 (N_3084,N_1118,N_76);
nor U3085 (N_3085,N_320,N_1299);
nand U3086 (N_3086,N_908,N_1091);
and U3087 (N_3087,N_1503,N_1418);
and U3088 (N_3088,N_891,N_1091);
or U3089 (N_3089,N_697,N_1040);
xor U3090 (N_3090,N_38,N_479);
nand U3091 (N_3091,N_91,N_1717);
or U3092 (N_3092,N_1626,N_344);
xor U3093 (N_3093,N_1804,N_227);
nand U3094 (N_3094,N_1643,N_1965);
xnor U3095 (N_3095,N_783,N_126);
xnor U3096 (N_3096,N_784,N_733);
xor U3097 (N_3097,N_1135,N_1217);
nand U3098 (N_3098,N_1583,N_1531);
or U3099 (N_3099,N_1486,N_655);
and U3100 (N_3100,N_1666,N_500);
and U3101 (N_3101,N_1364,N_957);
nand U3102 (N_3102,N_1147,N_286);
nor U3103 (N_3103,N_1503,N_1723);
nand U3104 (N_3104,N_1955,N_853);
nand U3105 (N_3105,N_128,N_583);
xnor U3106 (N_3106,N_167,N_1874);
or U3107 (N_3107,N_445,N_396);
or U3108 (N_3108,N_713,N_721);
nand U3109 (N_3109,N_815,N_301);
xnor U3110 (N_3110,N_1896,N_647);
and U3111 (N_3111,N_1557,N_1733);
or U3112 (N_3112,N_889,N_409);
xnor U3113 (N_3113,N_1828,N_1922);
nor U3114 (N_3114,N_234,N_227);
or U3115 (N_3115,N_644,N_1379);
nand U3116 (N_3116,N_892,N_540);
nor U3117 (N_3117,N_22,N_177);
nand U3118 (N_3118,N_226,N_292);
nor U3119 (N_3119,N_1620,N_1980);
and U3120 (N_3120,N_1586,N_864);
and U3121 (N_3121,N_1862,N_996);
nand U3122 (N_3122,N_799,N_1056);
or U3123 (N_3123,N_1928,N_744);
or U3124 (N_3124,N_283,N_1821);
nor U3125 (N_3125,N_204,N_1408);
xor U3126 (N_3126,N_563,N_1784);
and U3127 (N_3127,N_1899,N_1818);
nor U3128 (N_3128,N_1908,N_409);
or U3129 (N_3129,N_1546,N_1707);
nand U3130 (N_3130,N_792,N_1675);
nor U3131 (N_3131,N_988,N_476);
or U3132 (N_3132,N_696,N_961);
or U3133 (N_3133,N_824,N_1478);
nand U3134 (N_3134,N_399,N_996);
nor U3135 (N_3135,N_1418,N_1915);
nand U3136 (N_3136,N_794,N_1175);
nor U3137 (N_3137,N_903,N_1504);
xor U3138 (N_3138,N_325,N_681);
nor U3139 (N_3139,N_1608,N_808);
or U3140 (N_3140,N_1417,N_890);
and U3141 (N_3141,N_1857,N_1371);
nand U3142 (N_3142,N_1270,N_1696);
nand U3143 (N_3143,N_1477,N_1593);
nor U3144 (N_3144,N_421,N_1441);
and U3145 (N_3145,N_691,N_450);
and U3146 (N_3146,N_1586,N_1439);
xnor U3147 (N_3147,N_561,N_1938);
or U3148 (N_3148,N_1104,N_869);
and U3149 (N_3149,N_521,N_727);
or U3150 (N_3150,N_1987,N_590);
xor U3151 (N_3151,N_1071,N_830);
nor U3152 (N_3152,N_169,N_1140);
nand U3153 (N_3153,N_1209,N_6);
nand U3154 (N_3154,N_497,N_1302);
or U3155 (N_3155,N_1124,N_1000);
nor U3156 (N_3156,N_356,N_533);
and U3157 (N_3157,N_729,N_202);
or U3158 (N_3158,N_664,N_882);
nor U3159 (N_3159,N_685,N_640);
and U3160 (N_3160,N_1720,N_1727);
nor U3161 (N_3161,N_1732,N_940);
or U3162 (N_3162,N_1525,N_1918);
nor U3163 (N_3163,N_883,N_669);
xor U3164 (N_3164,N_306,N_397);
nand U3165 (N_3165,N_413,N_1665);
nor U3166 (N_3166,N_918,N_810);
nand U3167 (N_3167,N_1195,N_1577);
or U3168 (N_3168,N_820,N_880);
and U3169 (N_3169,N_939,N_1633);
and U3170 (N_3170,N_1772,N_285);
and U3171 (N_3171,N_372,N_1427);
or U3172 (N_3172,N_317,N_204);
and U3173 (N_3173,N_505,N_946);
nand U3174 (N_3174,N_1964,N_1217);
nand U3175 (N_3175,N_1982,N_954);
and U3176 (N_3176,N_390,N_1803);
nand U3177 (N_3177,N_1731,N_1526);
nor U3178 (N_3178,N_1000,N_1089);
or U3179 (N_3179,N_1974,N_1475);
or U3180 (N_3180,N_1633,N_1617);
nor U3181 (N_3181,N_417,N_1358);
or U3182 (N_3182,N_486,N_360);
nor U3183 (N_3183,N_138,N_1197);
nor U3184 (N_3184,N_1539,N_1900);
nor U3185 (N_3185,N_1530,N_1730);
xnor U3186 (N_3186,N_887,N_1658);
nor U3187 (N_3187,N_1749,N_769);
or U3188 (N_3188,N_1082,N_1409);
nand U3189 (N_3189,N_922,N_1197);
or U3190 (N_3190,N_1874,N_1621);
nor U3191 (N_3191,N_713,N_1493);
and U3192 (N_3192,N_1797,N_814);
nor U3193 (N_3193,N_1681,N_1543);
and U3194 (N_3194,N_472,N_1323);
nand U3195 (N_3195,N_1612,N_1988);
nor U3196 (N_3196,N_1030,N_1768);
and U3197 (N_3197,N_953,N_1860);
and U3198 (N_3198,N_108,N_617);
nand U3199 (N_3199,N_760,N_1062);
and U3200 (N_3200,N_1692,N_1999);
and U3201 (N_3201,N_617,N_13);
nand U3202 (N_3202,N_870,N_484);
nor U3203 (N_3203,N_1707,N_1394);
nor U3204 (N_3204,N_214,N_447);
nand U3205 (N_3205,N_1583,N_1294);
nand U3206 (N_3206,N_137,N_1485);
or U3207 (N_3207,N_591,N_1663);
and U3208 (N_3208,N_1,N_522);
nand U3209 (N_3209,N_222,N_808);
nor U3210 (N_3210,N_831,N_1376);
nor U3211 (N_3211,N_1235,N_1590);
and U3212 (N_3212,N_1041,N_1676);
or U3213 (N_3213,N_738,N_1165);
nor U3214 (N_3214,N_1102,N_1425);
nand U3215 (N_3215,N_1349,N_1768);
and U3216 (N_3216,N_23,N_423);
nand U3217 (N_3217,N_792,N_623);
or U3218 (N_3218,N_1758,N_1577);
nand U3219 (N_3219,N_539,N_234);
nor U3220 (N_3220,N_1530,N_1297);
or U3221 (N_3221,N_553,N_1170);
nand U3222 (N_3222,N_846,N_1494);
nor U3223 (N_3223,N_1171,N_1854);
and U3224 (N_3224,N_1848,N_372);
nand U3225 (N_3225,N_612,N_829);
and U3226 (N_3226,N_870,N_499);
nand U3227 (N_3227,N_247,N_1172);
nand U3228 (N_3228,N_1904,N_394);
and U3229 (N_3229,N_892,N_1495);
nor U3230 (N_3230,N_738,N_53);
xnor U3231 (N_3231,N_378,N_1122);
or U3232 (N_3232,N_628,N_23);
xor U3233 (N_3233,N_1009,N_117);
or U3234 (N_3234,N_852,N_599);
nor U3235 (N_3235,N_392,N_1039);
nor U3236 (N_3236,N_1831,N_1767);
nor U3237 (N_3237,N_1953,N_1909);
nor U3238 (N_3238,N_386,N_1124);
or U3239 (N_3239,N_161,N_113);
nor U3240 (N_3240,N_542,N_888);
nand U3241 (N_3241,N_1054,N_1530);
xor U3242 (N_3242,N_1099,N_1501);
nor U3243 (N_3243,N_1525,N_567);
and U3244 (N_3244,N_73,N_858);
nand U3245 (N_3245,N_1498,N_195);
nand U3246 (N_3246,N_1855,N_195);
xor U3247 (N_3247,N_1444,N_737);
nor U3248 (N_3248,N_1624,N_1802);
and U3249 (N_3249,N_1393,N_1323);
or U3250 (N_3250,N_730,N_1888);
nand U3251 (N_3251,N_809,N_1214);
nand U3252 (N_3252,N_151,N_612);
and U3253 (N_3253,N_183,N_1810);
xnor U3254 (N_3254,N_411,N_1966);
nor U3255 (N_3255,N_350,N_1322);
nor U3256 (N_3256,N_619,N_1915);
xnor U3257 (N_3257,N_1894,N_802);
or U3258 (N_3258,N_1914,N_952);
nand U3259 (N_3259,N_795,N_132);
nor U3260 (N_3260,N_1108,N_444);
nor U3261 (N_3261,N_1109,N_505);
nor U3262 (N_3262,N_105,N_1389);
nor U3263 (N_3263,N_591,N_1341);
or U3264 (N_3264,N_1384,N_521);
nor U3265 (N_3265,N_731,N_1586);
or U3266 (N_3266,N_793,N_542);
or U3267 (N_3267,N_1931,N_500);
or U3268 (N_3268,N_1258,N_1965);
nand U3269 (N_3269,N_1229,N_331);
nor U3270 (N_3270,N_1040,N_1495);
nor U3271 (N_3271,N_1141,N_889);
and U3272 (N_3272,N_29,N_43);
and U3273 (N_3273,N_1879,N_1193);
nor U3274 (N_3274,N_235,N_1080);
nand U3275 (N_3275,N_545,N_1181);
nand U3276 (N_3276,N_997,N_226);
nand U3277 (N_3277,N_1260,N_15);
nand U3278 (N_3278,N_1282,N_1251);
xor U3279 (N_3279,N_55,N_1948);
and U3280 (N_3280,N_1465,N_1188);
nor U3281 (N_3281,N_1032,N_700);
and U3282 (N_3282,N_303,N_1238);
nand U3283 (N_3283,N_909,N_540);
and U3284 (N_3284,N_1444,N_742);
and U3285 (N_3285,N_95,N_249);
or U3286 (N_3286,N_1586,N_1696);
or U3287 (N_3287,N_1035,N_1224);
and U3288 (N_3288,N_550,N_879);
xnor U3289 (N_3289,N_957,N_1783);
xor U3290 (N_3290,N_770,N_1429);
nor U3291 (N_3291,N_1210,N_1455);
xnor U3292 (N_3292,N_1425,N_1945);
nand U3293 (N_3293,N_30,N_1534);
and U3294 (N_3294,N_469,N_351);
or U3295 (N_3295,N_1902,N_1192);
or U3296 (N_3296,N_756,N_329);
or U3297 (N_3297,N_1733,N_1275);
nand U3298 (N_3298,N_1385,N_6);
nor U3299 (N_3299,N_765,N_1578);
nand U3300 (N_3300,N_414,N_1632);
and U3301 (N_3301,N_878,N_1801);
nand U3302 (N_3302,N_327,N_1935);
and U3303 (N_3303,N_135,N_430);
nor U3304 (N_3304,N_331,N_450);
or U3305 (N_3305,N_1597,N_438);
or U3306 (N_3306,N_93,N_769);
and U3307 (N_3307,N_1138,N_1585);
and U3308 (N_3308,N_890,N_333);
and U3309 (N_3309,N_1649,N_1852);
nor U3310 (N_3310,N_1851,N_1758);
xnor U3311 (N_3311,N_55,N_740);
or U3312 (N_3312,N_1777,N_443);
and U3313 (N_3313,N_433,N_580);
nor U3314 (N_3314,N_325,N_1304);
xnor U3315 (N_3315,N_51,N_744);
or U3316 (N_3316,N_39,N_1236);
nor U3317 (N_3317,N_626,N_1862);
or U3318 (N_3318,N_189,N_1006);
and U3319 (N_3319,N_83,N_1115);
and U3320 (N_3320,N_806,N_1391);
nand U3321 (N_3321,N_1452,N_192);
and U3322 (N_3322,N_1913,N_1120);
or U3323 (N_3323,N_660,N_897);
or U3324 (N_3324,N_479,N_164);
nand U3325 (N_3325,N_1927,N_442);
and U3326 (N_3326,N_1946,N_73);
or U3327 (N_3327,N_1639,N_1156);
nor U3328 (N_3328,N_667,N_1961);
nor U3329 (N_3329,N_1332,N_565);
or U3330 (N_3330,N_60,N_1102);
nor U3331 (N_3331,N_1017,N_434);
or U3332 (N_3332,N_1408,N_267);
or U3333 (N_3333,N_34,N_1770);
nor U3334 (N_3334,N_1253,N_1844);
nand U3335 (N_3335,N_677,N_270);
nor U3336 (N_3336,N_1419,N_285);
nand U3337 (N_3337,N_222,N_215);
nand U3338 (N_3338,N_846,N_85);
or U3339 (N_3339,N_1636,N_1278);
and U3340 (N_3340,N_638,N_37);
and U3341 (N_3341,N_1351,N_1970);
or U3342 (N_3342,N_237,N_457);
and U3343 (N_3343,N_890,N_553);
nor U3344 (N_3344,N_1175,N_184);
and U3345 (N_3345,N_647,N_1635);
or U3346 (N_3346,N_1122,N_1841);
or U3347 (N_3347,N_1214,N_1898);
and U3348 (N_3348,N_419,N_1904);
nor U3349 (N_3349,N_234,N_631);
xor U3350 (N_3350,N_177,N_1821);
xor U3351 (N_3351,N_1744,N_1040);
xnor U3352 (N_3352,N_329,N_64);
nor U3353 (N_3353,N_1319,N_1179);
nor U3354 (N_3354,N_699,N_1704);
nor U3355 (N_3355,N_1809,N_712);
nor U3356 (N_3356,N_1587,N_46);
or U3357 (N_3357,N_1588,N_603);
nor U3358 (N_3358,N_1283,N_546);
or U3359 (N_3359,N_1791,N_1378);
nor U3360 (N_3360,N_1743,N_1555);
or U3361 (N_3361,N_226,N_520);
nand U3362 (N_3362,N_8,N_1756);
xor U3363 (N_3363,N_145,N_852);
xor U3364 (N_3364,N_1475,N_941);
and U3365 (N_3365,N_401,N_1190);
nand U3366 (N_3366,N_1633,N_902);
xnor U3367 (N_3367,N_338,N_69);
and U3368 (N_3368,N_60,N_608);
nand U3369 (N_3369,N_431,N_1150);
nand U3370 (N_3370,N_454,N_809);
nor U3371 (N_3371,N_451,N_670);
and U3372 (N_3372,N_1742,N_1152);
or U3373 (N_3373,N_908,N_385);
nor U3374 (N_3374,N_1370,N_1252);
nand U3375 (N_3375,N_1183,N_1171);
nor U3376 (N_3376,N_892,N_880);
nor U3377 (N_3377,N_234,N_932);
nand U3378 (N_3378,N_165,N_1200);
nand U3379 (N_3379,N_1562,N_1134);
and U3380 (N_3380,N_789,N_166);
and U3381 (N_3381,N_1999,N_1063);
nor U3382 (N_3382,N_1243,N_1068);
xnor U3383 (N_3383,N_105,N_877);
nor U3384 (N_3384,N_756,N_1387);
xor U3385 (N_3385,N_172,N_681);
nand U3386 (N_3386,N_299,N_1811);
and U3387 (N_3387,N_1727,N_1970);
nand U3388 (N_3388,N_782,N_94);
nor U3389 (N_3389,N_1934,N_361);
or U3390 (N_3390,N_332,N_1996);
nand U3391 (N_3391,N_1370,N_1077);
nor U3392 (N_3392,N_1057,N_860);
and U3393 (N_3393,N_1041,N_1663);
nor U3394 (N_3394,N_1731,N_1838);
or U3395 (N_3395,N_1051,N_133);
or U3396 (N_3396,N_27,N_1596);
and U3397 (N_3397,N_1267,N_1506);
nor U3398 (N_3398,N_1429,N_1055);
or U3399 (N_3399,N_135,N_1174);
nand U3400 (N_3400,N_1573,N_574);
and U3401 (N_3401,N_1019,N_1694);
nor U3402 (N_3402,N_568,N_148);
nand U3403 (N_3403,N_1987,N_1414);
nor U3404 (N_3404,N_1453,N_1851);
or U3405 (N_3405,N_1377,N_497);
and U3406 (N_3406,N_1145,N_1397);
nand U3407 (N_3407,N_1482,N_1893);
xnor U3408 (N_3408,N_709,N_152);
xor U3409 (N_3409,N_605,N_232);
or U3410 (N_3410,N_1695,N_318);
or U3411 (N_3411,N_1432,N_89);
nor U3412 (N_3412,N_310,N_353);
nor U3413 (N_3413,N_821,N_557);
nor U3414 (N_3414,N_146,N_1228);
and U3415 (N_3415,N_562,N_1128);
nand U3416 (N_3416,N_1923,N_1779);
nor U3417 (N_3417,N_458,N_572);
xor U3418 (N_3418,N_975,N_1612);
or U3419 (N_3419,N_1131,N_591);
nor U3420 (N_3420,N_427,N_1829);
nor U3421 (N_3421,N_1910,N_988);
and U3422 (N_3422,N_793,N_1363);
nand U3423 (N_3423,N_1033,N_900);
or U3424 (N_3424,N_107,N_435);
and U3425 (N_3425,N_1229,N_1903);
nor U3426 (N_3426,N_60,N_15);
or U3427 (N_3427,N_305,N_241);
xor U3428 (N_3428,N_700,N_327);
nand U3429 (N_3429,N_1486,N_199);
nand U3430 (N_3430,N_1020,N_414);
and U3431 (N_3431,N_914,N_874);
nor U3432 (N_3432,N_1863,N_593);
or U3433 (N_3433,N_38,N_373);
nor U3434 (N_3434,N_1058,N_1525);
nor U3435 (N_3435,N_1267,N_1918);
and U3436 (N_3436,N_1108,N_843);
nor U3437 (N_3437,N_1313,N_1031);
and U3438 (N_3438,N_140,N_1546);
or U3439 (N_3439,N_279,N_491);
and U3440 (N_3440,N_185,N_1506);
nand U3441 (N_3441,N_469,N_674);
nand U3442 (N_3442,N_1875,N_1233);
nor U3443 (N_3443,N_433,N_1312);
and U3444 (N_3444,N_30,N_991);
nand U3445 (N_3445,N_1773,N_823);
nor U3446 (N_3446,N_392,N_1978);
xor U3447 (N_3447,N_846,N_713);
xnor U3448 (N_3448,N_1550,N_110);
and U3449 (N_3449,N_726,N_891);
xnor U3450 (N_3450,N_1753,N_1769);
and U3451 (N_3451,N_1277,N_1802);
nand U3452 (N_3452,N_1294,N_1186);
xnor U3453 (N_3453,N_833,N_525);
nor U3454 (N_3454,N_1435,N_197);
and U3455 (N_3455,N_1327,N_1413);
xor U3456 (N_3456,N_1879,N_1140);
nor U3457 (N_3457,N_1375,N_1590);
nand U3458 (N_3458,N_1373,N_1982);
nor U3459 (N_3459,N_1931,N_551);
nand U3460 (N_3460,N_196,N_698);
xor U3461 (N_3461,N_915,N_1963);
and U3462 (N_3462,N_363,N_622);
xor U3463 (N_3463,N_61,N_75);
nor U3464 (N_3464,N_1986,N_688);
or U3465 (N_3465,N_1886,N_658);
or U3466 (N_3466,N_1031,N_810);
nor U3467 (N_3467,N_532,N_822);
or U3468 (N_3468,N_236,N_647);
or U3469 (N_3469,N_827,N_1793);
or U3470 (N_3470,N_743,N_420);
nor U3471 (N_3471,N_1731,N_1065);
and U3472 (N_3472,N_674,N_466);
and U3473 (N_3473,N_819,N_1379);
nor U3474 (N_3474,N_1054,N_1253);
nor U3475 (N_3475,N_1342,N_18);
or U3476 (N_3476,N_854,N_459);
and U3477 (N_3477,N_218,N_1103);
nand U3478 (N_3478,N_546,N_928);
and U3479 (N_3479,N_1964,N_1946);
xnor U3480 (N_3480,N_955,N_883);
or U3481 (N_3481,N_1811,N_537);
nor U3482 (N_3482,N_269,N_1516);
and U3483 (N_3483,N_1103,N_1203);
and U3484 (N_3484,N_768,N_579);
xnor U3485 (N_3485,N_1370,N_651);
nand U3486 (N_3486,N_1860,N_333);
xnor U3487 (N_3487,N_920,N_421);
nand U3488 (N_3488,N_870,N_1963);
and U3489 (N_3489,N_414,N_133);
nand U3490 (N_3490,N_807,N_210);
or U3491 (N_3491,N_767,N_887);
nor U3492 (N_3492,N_1291,N_478);
nor U3493 (N_3493,N_1526,N_825);
or U3494 (N_3494,N_361,N_831);
nand U3495 (N_3495,N_1604,N_1825);
nand U3496 (N_3496,N_1858,N_1319);
and U3497 (N_3497,N_1246,N_115);
nor U3498 (N_3498,N_565,N_1217);
or U3499 (N_3499,N_1435,N_1169);
nor U3500 (N_3500,N_137,N_519);
and U3501 (N_3501,N_1769,N_670);
nand U3502 (N_3502,N_1429,N_1765);
nor U3503 (N_3503,N_989,N_1660);
nor U3504 (N_3504,N_1434,N_109);
nand U3505 (N_3505,N_441,N_1664);
nand U3506 (N_3506,N_1138,N_1050);
xnor U3507 (N_3507,N_1345,N_1134);
and U3508 (N_3508,N_1135,N_1316);
nand U3509 (N_3509,N_1115,N_1558);
nor U3510 (N_3510,N_439,N_1836);
nor U3511 (N_3511,N_1414,N_1562);
and U3512 (N_3512,N_1264,N_1768);
or U3513 (N_3513,N_1219,N_552);
nand U3514 (N_3514,N_294,N_558);
nor U3515 (N_3515,N_1568,N_1414);
nor U3516 (N_3516,N_473,N_1673);
xnor U3517 (N_3517,N_860,N_380);
or U3518 (N_3518,N_257,N_1481);
or U3519 (N_3519,N_1444,N_1820);
nand U3520 (N_3520,N_529,N_1645);
nor U3521 (N_3521,N_1857,N_81);
or U3522 (N_3522,N_1577,N_332);
and U3523 (N_3523,N_548,N_668);
nand U3524 (N_3524,N_1041,N_1100);
or U3525 (N_3525,N_1638,N_1472);
or U3526 (N_3526,N_329,N_1434);
nor U3527 (N_3527,N_1205,N_519);
nand U3528 (N_3528,N_292,N_23);
nand U3529 (N_3529,N_504,N_148);
and U3530 (N_3530,N_1501,N_1709);
xor U3531 (N_3531,N_1209,N_545);
nor U3532 (N_3532,N_275,N_1324);
and U3533 (N_3533,N_1779,N_620);
and U3534 (N_3534,N_472,N_689);
nand U3535 (N_3535,N_1678,N_1395);
and U3536 (N_3536,N_1845,N_1513);
nand U3537 (N_3537,N_1184,N_1304);
xor U3538 (N_3538,N_1504,N_960);
and U3539 (N_3539,N_625,N_1797);
nand U3540 (N_3540,N_772,N_1875);
nor U3541 (N_3541,N_709,N_744);
nand U3542 (N_3542,N_1688,N_799);
nand U3543 (N_3543,N_1609,N_1612);
or U3544 (N_3544,N_1857,N_142);
or U3545 (N_3545,N_175,N_24);
and U3546 (N_3546,N_281,N_1108);
nor U3547 (N_3547,N_476,N_1912);
xor U3548 (N_3548,N_1701,N_1177);
nor U3549 (N_3549,N_1553,N_936);
nand U3550 (N_3550,N_1012,N_1578);
or U3551 (N_3551,N_887,N_1853);
nor U3552 (N_3552,N_1325,N_1496);
or U3553 (N_3553,N_1617,N_736);
and U3554 (N_3554,N_1742,N_707);
and U3555 (N_3555,N_1324,N_1358);
or U3556 (N_3556,N_7,N_1598);
nand U3557 (N_3557,N_448,N_34);
or U3558 (N_3558,N_1391,N_1271);
and U3559 (N_3559,N_1973,N_587);
xnor U3560 (N_3560,N_281,N_1409);
and U3561 (N_3561,N_1287,N_1818);
and U3562 (N_3562,N_1489,N_245);
nor U3563 (N_3563,N_509,N_689);
and U3564 (N_3564,N_1054,N_386);
nand U3565 (N_3565,N_1863,N_1450);
nand U3566 (N_3566,N_695,N_1767);
nand U3567 (N_3567,N_1408,N_1296);
xor U3568 (N_3568,N_924,N_1324);
or U3569 (N_3569,N_1317,N_1653);
or U3570 (N_3570,N_1008,N_426);
and U3571 (N_3571,N_1004,N_851);
or U3572 (N_3572,N_1449,N_1434);
nand U3573 (N_3573,N_1410,N_1276);
nor U3574 (N_3574,N_843,N_940);
nor U3575 (N_3575,N_358,N_1964);
nor U3576 (N_3576,N_1145,N_1788);
nor U3577 (N_3577,N_1498,N_1564);
and U3578 (N_3578,N_1608,N_1986);
and U3579 (N_3579,N_241,N_381);
nand U3580 (N_3580,N_375,N_293);
and U3581 (N_3581,N_814,N_631);
nor U3582 (N_3582,N_427,N_696);
and U3583 (N_3583,N_917,N_8);
nand U3584 (N_3584,N_98,N_980);
nor U3585 (N_3585,N_1221,N_1484);
and U3586 (N_3586,N_438,N_234);
and U3587 (N_3587,N_0,N_1871);
xor U3588 (N_3588,N_582,N_641);
and U3589 (N_3589,N_314,N_184);
and U3590 (N_3590,N_1817,N_1019);
xnor U3591 (N_3591,N_1008,N_1354);
or U3592 (N_3592,N_1843,N_1524);
nor U3593 (N_3593,N_1441,N_111);
nand U3594 (N_3594,N_1373,N_568);
nand U3595 (N_3595,N_445,N_397);
or U3596 (N_3596,N_1731,N_1782);
nor U3597 (N_3597,N_598,N_1546);
xor U3598 (N_3598,N_383,N_1081);
or U3599 (N_3599,N_1722,N_1219);
or U3600 (N_3600,N_645,N_18);
nand U3601 (N_3601,N_1235,N_1835);
nor U3602 (N_3602,N_1027,N_1897);
and U3603 (N_3603,N_613,N_8);
nor U3604 (N_3604,N_1183,N_703);
nand U3605 (N_3605,N_723,N_374);
or U3606 (N_3606,N_1313,N_1514);
xnor U3607 (N_3607,N_162,N_970);
xor U3608 (N_3608,N_1728,N_1413);
or U3609 (N_3609,N_668,N_991);
nand U3610 (N_3610,N_1818,N_1260);
nand U3611 (N_3611,N_5,N_1069);
nand U3612 (N_3612,N_755,N_1738);
xnor U3613 (N_3613,N_92,N_1299);
nor U3614 (N_3614,N_1636,N_758);
or U3615 (N_3615,N_91,N_611);
xor U3616 (N_3616,N_1804,N_1603);
nor U3617 (N_3617,N_117,N_65);
nor U3618 (N_3618,N_396,N_339);
or U3619 (N_3619,N_83,N_1445);
nor U3620 (N_3620,N_836,N_1354);
or U3621 (N_3621,N_450,N_1689);
and U3622 (N_3622,N_1959,N_1024);
or U3623 (N_3623,N_1596,N_484);
nand U3624 (N_3624,N_1624,N_945);
or U3625 (N_3625,N_1482,N_1357);
and U3626 (N_3626,N_595,N_572);
nand U3627 (N_3627,N_1307,N_777);
nor U3628 (N_3628,N_596,N_1621);
and U3629 (N_3629,N_307,N_1424);
and U3630 (N_3630,N_1686,N_907);
nor U3631 (N_3631,N_1490,N_592);
or U3632 (N_3632,N_1220,N_427);
nand U3633 (N_3633,N_40,N_1289);
or U3634 (N_3634,N_1858,N_1925);
and U3635 (N_3635,N_689,N_612);
and U3636 (N_3636,N_1523,N_1785);
nor U3637 (N_3637,N_365,N_775);
nand U3638 (N_3638,N_659,N_82);
and U3639 (N_3639,N_1119,N_1834);
xnor U3640 (N_3640,N_398,N_1518);
and U3641 (N_3641,N_1295,N_58);
and U3642 (N_3642,N_1767,N_999);
nor U3643 (N_3643,N_112,N_930);
nand U3644 (N_3644,N_434,N_232);
nand U3645 (N_3645,N_1494,N_893);
or U3646 (N_3646,N_1689,N_1572);
or U3647 (N_3647,N_1333,N_1827);
and U3648 (N_3648,N_1806,N_1952);
and U3649 (N_3649,N_1338,N_1837);
nor U3650 (N_3650,N_644,N_851);
and U3651 (N_3651,N_612,N_1619);
nand U3652 (N_3652,N_318,N_1408);
nor U3653 (N_3653,N_302,N_1340);
xnor U3654 (N_3654,N_1439,N_1630);
nor U3655 (N_3655,N_220,N_84);
or U3656 (N_3656,N_1453,N_718);
and U3657 (N_3657,N_244,N_593);
and U3658 (N_3658,N_1333,N_26);
nand U3659 (N_3659,N_836,N_1991);
nand U3660 (N_3660,N_1819,N_1738);
xnor U3661 (N_3661,N_702,N_720);
nand U3662 (N_3662,N_860,N_125);
nand U3663 (N_3663,N_1086,N_1744);
and U3664 (N_3664,N_154,N_27);
xor U3665 (N_3665,N_1433,N_1161);
and U3666 (N_3666,N_346,N_1548);
and U3667 (N_3667,N_1359,N_1912);
or U3668 (N_3668,N_618,N_922);
nand U3669 (N_3669,N_1355,N_110);
and U3670 (N_3670,N_600,N_456);
nor U3671 (N_3671,N_1041,N_1948);
and U3672 (N_3672,N_1471,N_753);
nor U3673 (N_3673,N_1505,N_1917);
nor U3674 (N_3674,N_778,N_738);
nand U3675 (N_3675,N_1178,N_717);
or U3676 (N_3676,N_1144,N_480);
nand U3677 (N_3677,N_1078,N_128);
nor U3678 (N_3678,N_1086,N_943);
nand U3679 (N_3679,N_1532,N_1727);
nand U3680 (N_3680,N_1323,N_521);
nor U3681 (N_3681,N_156,N_275);
nor U3682 (N_3682,N_340,N_1294);
xor U3683 (N_3683,N_1321,N_492);
or U3684 (N_3684,N_296,N_928);
nand U3685 (N_3685,N_713,N_425);
nor U3686 (N_3686,N_218,N_1412);
and U3687 (N_3687,N_1405,N_246);
and U3688 (N_3688,N_1573,N_1627);
and U3689 (N_3689,N_1812,N_1669);
or U3690 (N_3690,N_174,N_966);
nand U3691 (N_3691,N_708,N_1357);
and U3692 (N_3692,N_346,N_839);
and U3693 (N_3693,N_354,N_1468);
xor U3694 (N_3694,N_903,N_998);
and U3695 (N_3695,N_1254,N_751);
nand U3696 (N_3696,N_717,N_1837);
or U3697 (N_3697,N_564,N_23);
and U3698 (N_3698,N_528,N_581);
nand U3699 (N_3699,N_1005,N_78);
or U3700 (N_3700,N_521,N_1852);
and U3701 (N_3701,N_624,N_583);
and U3702 (N_3702,N_450,N_655);
and U3703 (N_3703,N_457,N_1329);
nand U3704 (N_3704,N_999,N_1051);
or U3705 (N_3705,N_977,N_96);
or U3706 (N_3706,N_508,N_491);
nor U3707 (N_3707,N_260,N_1732);
or U3708 (N_3708,N_181,N_59);
nand U3709 (N_3709,N_945,N_1153);
and U3710 (N_3710,N_1540,N_797);
or U3711 (N_3711,N_78,N_1203);
nor U3712 (N_3712,N_505,N_1078);
nand U3713 (N_3713,N_170,N_1447);
nor U3714 (N_3714,N_1245,N_835);
xnor U3715 (N_3715,N_1164,N_293);
nand U3716 (N_3716,N_1344,N_1464);
xor U3717 (N_3717,N_1562,N_158);
xor U3718 (N_3718,N_574,N_59);
xor U3719 (N_3719,N_1908,N_381);
xor U3720 (N_3720,N_1392,N_579);
and U3721 (N_3721,N_771,N_1105);
and U3722 (N_3722,N_726,N_1221);
nand U3723 (N_3723,N_1120,N_273);
xor U3724 (N_3724,N_835,N_1734);
and U3725 (N_3725,N_169,N_1694);
and U3726 (N_3726,N_760,N_1755);
nor U3727 (N_3727,N_1023,N_1451);
and U3728 (N_3728,N_1270,N_584);
or U3729 (N_3729,N_1981,N_752);
nor U3730 (N_3730,N_1752,N_1999);
nand U3731 (N_3731,N_1246,N_1434);
nand U3732 (N_3732,N_293,N_1941);
nand U3733 (N_3733,N_29,N_262);
nand U3734 (N_3734,N_1301,N_134);
nand U3735 (N_3735,N_617,N_760);
nor U3736 (N_3736,N_1757,N_622);
nand U3737 (N_3737,N_1492,N_1748);
nor U3738 (N_3738,N_1140,N_1193);
nand U3739 (N_3739,N_1048,N_247);
nand U3740 (N_3740,N_1581,N_516);
or U3741 (N_3741,N_600,N_1181);
or U3742 (N_3742,N_908,N_617);
nand U3743 (N_3743,N_61,N_980);
and U3744 (N_3744,N_422,N_535);
nand U3745 (N_3745,N_1843,N_822);
or U3746 (N_3746,N_1787,N_1862);
or U3747 (N_3747,N_960,N_329);
and U3748 (N_3748,N_595,N_1575);
or U3749 (N_3749,N_1841,N_292);
or U3750 (N_3750,N_164,N_289);
or U3751 (N_3751,N_1791,N_341);
or U3752 (N_3752,N_363,N_830);
and U3753 (N_3753,N_988,N_179);
nor U3754 (N_3754,N_707,N_1427);
nand U3755 (N_3755,N_537,N_1717);
and U3756 (N_3756,N_1236,N_1076);
and U3757 (N_3757,N_820,N_1727);
nor U3758 (N_3758,N_1336,N_543);
and U3759 (N_3759,N_1708,N_1713);
nand U3760 (N_3760,N_345,N_1069);
and U3761 (N_3761,N_1309,N_1529);
or U3762 (N_3762,N_576,N_1322);
nand U3763 (N_3763,N_877,N_1847);
nor U3764 (N_3764,N_61,N_1557);
or U3765 (N_3765,N_28,N_1417);
nand U3766 (N_3766,N_1067,N_55);
and U3767 (N_3767,N_1452,N_1237);
nand U3768 (N_3768,N_1347,N_1330);
xor U3769 (N_3769,N_1575,N_1026);
nor U3770 (N_3770,N_760,N_942);
or U3771 (N_3771,N_1857,N_525);
and U3772 (N_3772,N_1594,N_1690);
or U3773 (N_3773,N_102,N_1851);
and U3774 (N_3774,N_129,N_1930);
xor U3775 (N_3775,N_490,N_275);
nand U3776 (N_3776,N_1068,N_775);
or U3777 (N_3777,N_1692,N_1218);
nand U3778 (N_3778,N_635,N_1986);
nor U3779 (N_3779,N_1203,N_181);
and U3780 (N_3780,N_1612,N_1192);
nand U3781 (N_3781,N_1704,N_1207);
or U3782 (N_3782,N_1799,N_186);
and U3783 (N_3783,N_1937,N_545);
nor U3784 (N_3784,N_897,N_1600);
or U3785 (N_3785,N_874,N_186);
nor U3786 (N_3786,N_222,N_910);
nor U3787 (N_3787,N_1406,N_420);
xor U3788 (N_3788,N_1369,N_1753);
and U3789 (N_3789,N_627,N_825);
nor U3790 (N_3790,N_184,N_1266);
and U3791 (N_3791,N_1839,N_940);
or U3792 (N_3792,N_1029,N_1740);
and U3793 (N_3793,N_670,N_1321);
and U3794 (N_3794,N_1969,N_1036);
or U3795 (N_3795,N_1289,N_68);
and U3796 (N_3796,N_860,N_1307);
or U3797 (N_3797,N_343,N_1257);
nand U3798 (N_3798,N_269,N_1084);
and U3799 (N_3799,N_134,N_753);
and U3800 (N_3800,N_1700,N_1784);
and U3801 (N_3801,N_1178,N_798);
or U3802 (N_3802,N_14,N_1491);
xnor U3803 (N_3803,N_1050,N_526);
nand U3804 (N_3804,N_1890,N_1374);
nand U3805 (N_3805,N_326,N_723);
xor U3806 (N_3806,N_736,N_1638);
and U3807 (N_3807,N_1483,N_336);
and U3808 (N_3808,N_360,N_1005);
and U3809 (N_3809,N_103,N_1883);
nor U3810 (N_3810,N_1502,N_1506);
and U3811 (N_3811,N_1357,N_1233);
or U3812 (N_3812,N_1866,N_1947);
nand U3813 (N_3813,N_1576,N_1973);
nor U3814 (N_3814,N_685,N_74);
and U3815 (N_3815,N_1432,N_362);
nand U3816 (N_3816,N_1769,N_1820);
xnor U3817 (N_3817,N_1476,N_1195);
nand U3818 (N_3818,N_664,N_1762);
xnor U3819 (N_3819,N_1127,N_776);
or U3820 (N_3820,N_746,N_1179);
nor U3821 (N_3821,N_1331,N_1493);
and U3822 (N_3822,N_1677,N_1367);
or U3823 (N_3823,N_797,N_303);
nand U3824 (N_3824,N_1922,N_1501);
xnor U3825 (N_3825,N_1573,N_191);
and U3826 (N_3826,N_1665,N_1483);
nand U3827 (N_3827,N_964,N_1522);
or U3828 (N_3828,N_1370,N_1575);
and U3829 (N_3829,N_391,N_1889);
nand U3830 (N_3830,N_853,N_1875);
or U3831 (N_3831,N_1973,N_1029);
or U3832 (N_3832,N_89,N_65);
or U3833 (N_3833,N_548,N_145);
and U3834 (N_3834,N_460,N_1306);
nand U3835 (N_3835,N_283,N_920);
nor U3836 (N_3836,N_5,N_965);
nand U3837 (N_3837,N_1876,N_281);
nand U3838 (N_3838,N_1372,N_112);
nor U3839 (N_3839,N_1540,N_290);
xnor U3840 (N_3840,N_1691,N_1584);
or U3841 (N_3841,N_1203,N_1434);
nor U3842 (N_3842,N_394,N_1884);
and U3843 (N_3843,N_1028,N_721);
and U3844 (N_3844,N_192,N_194);
nand U3845 (N_3845,N_561,N_1253);
nand U3846 (N_3846,N_285,N_301);
nor U3847 (N_3847,N_1071,N_1514);
and U3848 (N_3848,N_970,N_178);
nor U3849 (N_3849,N_437,N_1521);
or U3850 (N_3850,N_370,N_372);
nand U3851 (N_3851,N_328,N_1762);
nor U3852 (N_3852,N_877,N_1113);
and U3853 (N_3853,N_1054,N_1523);
nand U3854 (N_3854,N_21,N_613);
xnor U3855 (N_3855,N_933,N_1203);
or U3856 (N_3856,N_1861,N_306);
and U3857 (N_3857,N_306,N_851);
nand U3858 (N_3858,N_1728,N_1568);
or U3859 (N_3859,N_1554,N_1510);
and U3860 (N_3860,N_1370,N_1398);
and U3861 (N_3861,N_14,N_980);
nand U3862 (N_3862,N_640,N_1689);
and U3863 (N_3863,N_1061,N_61);
and U3864 (N_3864,N_207,N_614);
nand U3865 (N_3865,N_1292,N_864);
nand U3866 (N_3866,N_356,N_240);
or U3867 (N_3867,N_1973,N_1425);
and U3868 (N_3868,N_623,N_1873);
xnor U3869 (N_3869,N_1835,N_860);
or U3870 (N_3870,N_1203,N_897);
nand U3871 (N_3871,N_1896,N_637);
nand U3872 (N_3872,N_1433,N_1222);
xnor U3873 (N_3873,N_630,N_1332);
nand U3874 (N_3874,N_537,N_793);
nand U3875 (N_3875,N_1988,N_874);
and U3876 (N_3876,N_1472,N_181);
and U3877 (N_3877,N_453,N_182);
and U3878 (N_3878,N_271,N_1486);
nor U3879 (N_3879,N_1304,N_1299);
nand U3880 (N_3880,N_13,N_801);
and U3881 (N_3881,N_307,N_771);
nand U3882 (N_3882,N_566,N_573);
nand U3883 (N_3883,N_776,N_1475);
xnor U3884 (N_3884,N_999,N_1070);
or U3885 (N_3885,N_299,N_887);
and U3886 (N_3886,N_769,N_533);
xor U3887 (N_3887,N_0,N_560);
nor U3888 (N_3888,N_213,N_979);
nand U3889 (N_3889,N_1440,N_418);
or U3890 (N_3890,N_716,N_820);
and U3891 (N_3891,N_941,N_929);
xor U3892 (N_3892,N_751,N_1185);
and U3893 (N_3893,N_82,N_715);
xor U3894 (N_3894,N_681,N_1691);
and U3895 (N_3895,N_216,N_294);
nand U3896 (N_3896,N_281,N_952);
and U3897 (N_3897,N_1714,N_792);
nor U3898 (N_3898,N_1644,N_1653);
nand U3899 (N_3899,N_687,N_513);
and U3900 (N_3900,N_1427,N_1094);
xor U3901 (N_3901,N_1174,N_3);
nand U3902 (N_3902,N_1680,N_1668);
xnor U3903 (N_3903,N_1024,N_936);
nand U3904 (N_3904,N_86,N_288);
nand U3905 (N_3905,N_266,N_17);
or U3906 (N_3906,N_1025,N_724);
xor U3907 (N_3907,N_1055,N_1400);
xnor U3908 (N_3908,N_46,N_1968);
nor U3909 (N_3909,N_1327,N_1047);
or U3910 (N_3910,N_1686,N_219);
nor U3911 (N_3911,N_1109,N_1641);
and U3912 (N_3912,N_90,N_5);
nand U3913 (N_3913,N_33,N_1783);
or U3914 (N_3914,N_1151,N_244);
and U3915 (N_3915,N_1948,N_609);
and U3916 (N_3916,N_398,N_297);
or U3917 (N_3917,N_1708,N_1876);
nor U3918 (N_3918,N_746,N_708);
nand U3919 (N_3919,N_606,N_1646);
and U3920 (N_3920,N_1237,N_841);
and U3921 (N_3921,N_840,N_1028);
nand U3922 (N_3922,N_1213,N_784);
nor U3923 (N_3923,N_1371,N_1225);
nand U3924 (N_3924,N_518,N_1971);
nor U3925 (N_3925,N_936,N_1429);
nor U3926 (N_3926,N_128,N_1779);
and U3927 (N_3927,N_1344,N_27);
nand U3928 (N_3928,N_287,N_1164);
xor U3929 (N_3929,N_575,N_310);
nor U3930 (N_3930,N_1135,N_169);
or U3931 (N_3931,N_1959,N_370);
or U3932 (N_3932,N_981,N_1717);
nor U3933 (N_3933,N_1223,N_1480);
nor U3934 (N_3934,N_1998,N_1250);
and U3935 (N_3935,N_1967,N_1865);
xor U3936 (N_3936,N_64,N_1875);
nand U3937 (N_3937,N_1509,N_1213);
or U3938 (N_3938,N_1751,N_93);
and U3939 (N_3939,N_1099,N_1765);
and U3940 (N_3940,N_40,N_784);
xnor U3941 (N_3941,N_981,N_1990);
and U3942 (N_3942,N_529,N_1766);
and U3943 (N_3943,N_1493,N_308);
xor U3944 (N_3944,N_211,N_1393);
or U3945 (N_3945,N_1341,N_1458);
nor U3946 (N_3946,N_1935,N_1181);
or U3947 (N_3947,N_1787,N_416);
and U3948 (N_3948,N_1108,N_1849);
nand U3949 (N_3949,N_1729,N_786);
xor U3950 (N_3950,N_335,N_11);
nor U3951 (N_3951,N_23,N_1899);
or U3952 (N_3952,N_1968,N_212);
nor U3953 (N_3953,N_1677,N_219);
or U3954 (N_3954,N_414,N_266);
xnor U3955 (N_3955,N_1789,N_336);
nor U3956 (N_3956,N_1112,N_1902);
or U3957 (N_3957,N_40,N_1486);
nor U3958 (N_3958,N_1691,N_1384);
or U3959 (N_3959,N_701,N_834);
xnor U3960 (N_3960,N_876,N_667);
nand U3961 (N_3961,N_51,N_1102);
nand U3962 (N_3962,N_1162,N_417);
or U3963 (N_3963,N_835,N_1837);
or U3964 (N_3964,N_1956,N_1214);
nand U3965 (N_3965,N_1573,N_703);
and U3966 (N_3966,N_704,N_801);
xor U3967 (N_3967,N_367,N_1314);
and U3968 (N_3968,N_1801,N_67);
and U3969 (N_3969,N_1948,N_1515);
nor U3970 (N_3970,N_1243,N_1070);
nor U3971 (N_3971,N_398,N_507);
nor U3972 (N_3972,N_934,N_148);
nor U3973 (N_3973,N_517,N_1395);
xor U3974 (N_3974,N_820,N_70);
nor U3975 (N_3975,N_604,N_1324);
xnor U3976 (N_3976,N_57,N_1377);
xnor U3977 (N_3977,N_23,N_226);
nand U3978 (N_3978,N_1289,N_435);
and U3979 (N_3979,N_123,N_1091);
nand U3980 (N_3980,N_1113,N_1539);
nor U3981 (N_3981,N_778,N_1560);
nand U3982 (N_3982,N_932,N_1348);
nor U3983 (N_3983,N_1287,N_1246);
nor U3984 (N_3984,N_1029,N_808);
nor U3985 (N_3985,N_460,N_1074);
and U3986 (N_3986,N_975,N_1715);
nor U3987 (N_3987,N_1004,N_1327);
and U3988 (N_3988,N_416,N_5);
nand U3989 (N_3989,N_1542,N_772);
nand U3990 (N_3990,N_1740,N_139);
nand U3991 (N_3991,N_1614,N_1172);
xnor U3992 (N_3992,N_861,N_1369);
nor U3993 (N_3993,N_711,N_767);
and U3994 (N_3994,N_1719,N_1983);
nor U3995 (N_3995,N_269,N_1158);
nor U3996 (N_3996,N_1782,N_1126);
and U3997 (N_3997,N_1444,N_1152);
or U3998 (N_3998,N_1229,N_960);
xor U3999 (N_3999,N_474,N_114);
nand U4000 (N_4000,N_2085,N_2857);
and U4001 (N_4001,N_3479,N_2025);
nor U4002 (N_4002,N_2839,N_3532);
nor U4003 (N_4003,N_2616,N_3014);
nor U4004 (N_4004,N_2416,N_2331);
and U4005 (N_4005,N_3525,N_2846);
nand U4006 (N_4006,N_3789,N_2958);
xnor U4007 (N_4007,N_3164,N_3410);
nor U4008 (N_4008,N_2192,N_3631);
and U4009 (N_4009,N_2594,N_3622);
nand U4010 (N_4010,N_3683,N_2008);
nand U4011 (N_4011,N_3881,N_3327);
xor U4012 (N_4012,N_3895,N_3701);
and U4013 (N_4013,N_2021,N_2893);
and U4014 (N_4014,N_2010,N_3562);
and U4015 (N_4015,N_3641,N_3768);
nor U4016 (N_4016,N_3632,N_3766);
nor U4017 (N_4017,N_2520,N_2411);
or U4018 (N_4018,N_2737,N_2926);
nor U4019 (N_4019,N_2135,N_3630);
nor U4020 (N_4020,N_3772,N_2913);
and U4021 (N_4021,N_3500,N_3537);
xor U4022 (N_4022,N_2239,N_2662);
xnor U4023 (N_4023,N_2299,N_3494);
or U4024 (N_4024,N_2775,N_3023);
nor U4025 (N_4025,N_2124,N_3288);
xnor U4026 (N_4026,N_3798,N_2671);
and U4027 (N_4027,N_2885,N_2983);
xor U4028 (N_4028,N_3841,N_3316);
and U4029 (N_4029,N_3152,N_2452);
or U4030 (N_4030,N_3922,N_3696);
nand U4031 (N_4031,N_3436,N_3963);
nand U4032 (N_4032,N_2250,N_3313);
nand U4033 (N_4033,N_2198,N_3070);
and U4034 (N_4034,N_3542,N_3967);
and U4035 (N_4035,N_3473,N_3471);
nand U4036 (N_4036,N_3433,N_3034);
nand U4037 (N_4037,N_3909,N_3364);
nor U4038 (N_4038,N_2854,N_3733);
and U4039 (N_4039,N_3634,N_3707);
and U4040 (N_4040,N_2747,N_2631);
xor U4041 (N_4041,N_3894,N_2611);
nor U4042 (N_4042,N_3348,N_3383);
nand U4043 (N_4043,N_3217,N_2308);
or U4044 (N_4044,N_3041,N_2829);
or U4045 (N_4045,N_3935,N_3816);
or U4046 (N_4046,N_2472,N_2095);
and U4047 (N_4047,N_2546,N_3178);
nand U4048 (N_4048,N_2886,N_2773);
nor U4049 (N_4049,N_2238,N_2887);
or U4050 (N_4050,N_3345,N_3510);
and U4051 (N_4051,N_3251,N_2723);
and U4052 (N_4052,N_2027,N_3516);
or U4053 (N_4053,N_3786,N_2966);
nand U4054 (N_4054,N_3310,N_3292);
or U4055 (N_4055,N_2278,N_2272);
and U4056 (N_4056,N_3547,N_2447);
and U4057 (N_4057,N_3531,N_2175);
xnor U4058 (N_4058,N_3420,N_2940);
nand U4059 (N_4059,N_3678,N_2078);
nand U4060 (N_4060,N_3872,N_2721);
or U4061 (N_4061,N_2043,N_2634);
or U4062 (N_4062,N_2202,N_3003);
or U4063 (N_4063,N_3725,N_3434);
and U4064 (N_4064,N_2882,N_2565);
nor U4065 (N_4065,N_2446,N_3151);
nand U4066 (N_4066,N_3888,N_3892);
and U4067 (N_4067,N_2637,N_3513);
xor U4068 (N_4068,N_2228,N_3394);
and U4069 (N_4069,N_2639,N_3214);
xor U4070 (N_4070,N_2449,N_2177);
nand U4071 (N_4071,N_3194,N_3447);
xor U4072 (N_4072,N_2034,N_3493);
or U4073 (N_4073,N_2211,N_2091);
or U4074 (N_4074,N_2516,N_2458);
or U4075 (N_4075,N_2699,N_2950);
and U4076 (N_4076,N_3134,N_2848);
or U4077 (N_4077,N_3769,N_3889);
and U4078 (N_4078,N_2148,N_2407);
nor U4079 (N_4079,N_3849,N_2361);
and U4080 (N_4080,N_3395,N_3893);
nor U4081 (N_4081,N_2477,N_2026);
and U4082 (N_4082,N_3486,N_2076);
or U4083 (N_4083,N_3613,N_2698);
nor U4084 (N_4084,N_3688,N_3737);
nor U4085 (N_4085,N_2469,N_2310);
nor U4086 (N_4086,N_2823,N_2767);
or U4087 (N_4087,N_3740,N_2618);
nand U4088 (N_4088,N_3643,N_3011);
and U4089 (N_4089,N_3407,N_3539);
nand U4090 (N_4090,N_3418,N_3142);
nor U4091 (N_4091,N_2867,N_3747);
nor U4092 (N_4092,N_2147,N_3211);
or U4093 (N_4093,N_3923,N_2741);
xnor U4094 (N_4094,N_2997,N_2930);
and U4095 (N_4095,N_3955,N_2931);
or U4096 (N_4096,N_3681,N_3807);
xor U4097 (N_4097,N_3148,N_3946);
nand U4098 (N_4098,N_3633,N_3903);
or U4099 (N_4099,N_2744,N_2579);
nand U4100 (N_4100,N_2113,N_2871);
xor U4101 (N_4101,N_3442,N_3022);
nand U4102 (N_4102,N_2053,N_2646);
nor U4103 (N_4103,N_2970,N_2204);
and U4104 (N_4104,N_3331,N_2367);
nor U4105 (N_4105,N_2837,N_2203);
xor U4106 (N_4106,N_3521,N_2644);
nand U4107 (N_4107,N_3049,N_3422);
and U4108 (N_4108,N_2223,N_3392);
nor U4109 (N_4109,N_2521,N_2011);
and U4110 (N_4110,N_3225,N_2197);
nor U4111 (N_4111,N_3728,N_3149);
nor U4112 (N_4112,N_3722,N_3646);
and U4113 (N_4113,N_3100,N_3937);
and U4114 (N_4114,N_2511,N_3750);
nand U4115 (N_4115,N_3748,N_2921);
nand U4116 (N_4116,N_3126,N_2051);
or U4117 (N_4117,N_2056,N_3204);
or U4118 (N_4118,N_2217,N_2083);
and U4119 (N_4119,N_2934,N_3044);
and U4120 (N_4120,N_3844,N_2112);
nor U4121 (N_4121,N_3649,N_2852);
nor U4122 (N_4122,N_3372,N_3778);
nor U4123 (N_4123,N_2720,N_3639);
or U4124 (N_4124,N_2064,N_3465);
and U4125 (N_4125,N_2879,N_2222);
nand U4126 (N_4126,N_3572,N_3197);
nand U4127 (N_4127,N_2005,N_2125);
nand U4128 (N_4128,N_3341,N_3709);
and U4129 (N_4129,N_2451,N_3424);
and U4130 (N_4130,N_3001,N_2082);
or U4131 (N_4131,N_3168,N_2249);
or U4132 (N_4132,N_3081,N_2794);
nand U4133 (N_4133,N_2398,N_2586);
or U4134 (N_4134,N_2130,N_3818);
and U4135 (N_4135,N_3915,N_2880);
nor U4136 (N_4136,N_3676,N_2589);
xnor U4137 (N_4137,N_2828,N_3721);
or U4138 (N_4138,N_3259,N_3045);
nor U4139 (N_4139,N_3851,N_3403);
xor U4140 (N_4140,N_2141,N_3947);
or U4141 (N_4141,N_3796,N_3535);
and U4142 (N_4142,N_2830,N_2975);
nor U4143 (N_4143,N_3651,N_2677);
nand U4144 (N_4144,N_2633,N_2179);
and U4145 (N_4145,N_2137,N_2971);
and U4146 (N_4146,N_3610,N_2094);
nand U4147 (N_4147,N_3891,N_2595);
nor U4148 (N_4148,N_3864,N_2136);
nor U4149 (N_4149,N_2587,N_2015);
or U4150 (N_4150,N_2001,N_2706);
xor U4151 (N_4151,N_3875,N_3674);
nor U4152 (N_4152,N_3705,N_2189);
nor U4153 (N_4153,N_2526,N_2678);
nand U4154 (N_4154,N_2332,N_3456);
and U4155 (N_4155,N_2414,N_3354);
and U4156 (N_4156,N_3555,N_3693);
nor U4157 (N_4157,N_3462,N_3557);
nor U4158 (N_4158,N_3093,N_2592);
nand U4159 (N_4159,N_3520,N_3921);
xor U4160 (N_4160,N_2075,N_3538);
and U4161 (N_4161,N_3443,N_2949);
nand U4162 (N_4162,N_3687,N_3227);
nor U4163 (N_4163,N_2626,N_2455);
and U4164 (N_4164,N_2036,N_2193);
or U4165 (N_4165,N_3363,N_2230);
nor U4166 (N_4166,N_3604,N_3644);
and U4167 (N_4167,N_3573,N_2500);
and U4168 (N_4168,N_3220,N_2717);
and U4169 (N_4169,N_2327,N_2924);
nand U4170 (N_4170,N_2743,N_3770);
nor U4171 (N_4171,N_2868,N_2870);
and U4172 (N_4172,N_3333,N_2606);
and U4173 (N_4173,N_2653,N_3458);
nand U4174 (N_4174,N_3871,N_2201);
xnor U4175 (N_4175,N_3758,N_3744);
nand U4176 (N_4176,N_3794,N_3177);
and U4177 (N_4177,N_3916,N_2935);
nor U4178 (N_4178,N_3673,N_2672);
or U4179 (N_4179,N_2263,N_3258);
nor U4180 (N_4180,N_2004,N_3317);
and U4181 (N_4181,N_3241,N_3717);
nand U4182 (N_4182,N_2369,N_3672);
nand U4183 (N_4183,N_3312,N_2922);
nor U4184 (N_4184,N_3118,N_2173);
nand U4185 (N_4185,N_2408,N_2553);
or U4186 (N_4186,N_3508,N_3847);
or U4187 (N_4187,N_2814,N_3415);
and U4188 (N_4188,N_2547,N_2302);
xor U4189 (N_4189,N_3273,N_2980);
xor U4190 (N_4190,N_3083,N_3039);
nand U4191 (N_4191,N_3397,N_2030);
or U4192 (N_4192,N_3960,N_2844);
xor U4193 (N_4193,N_2326,N_2029);
nand U4194 (N_4194,N_2480,N_2467);
nor U4195 (N_4195,N_3054,N_2896);
nor U4196 (N_4196,N_2304,N_3232);
nor U4197 (N_4197,N_2178,N_2279);
or U4198 (N_4198,N_2110,N_2253);
nor U4199 (N_4199,N_2804,N_2023);
xor U4200 (N_4200,N_2766,N_3788);
nand U4201 (N_4201,N_2769,N_3669);
and U4202 (N_4202,N_3136,N_3976);
and U4203 (N_4203,N_3635,N_3699);
and U4204 (N_4204,N_2007,N_3096);
and U4205 (N_4205,N_3529,N_2607);
nand U4206 (N_4206,N_2803,N_2615);
or U4207 (N_4207,N_3838,N_3533);
nand U4208 (N_4208,N_3412,N_2321);
and U4209 (N_4209,N_3575,N_2542);
nor U4210 (N_4210,N_3624,N_2325);
or U4211 (N_4211,N_2726,N_2000);
xnor U4212 (N_4212,N_3013,N_3839);
or U4213 (N_4213,N_2227,N_2624);
xnor U4214 (N_4214,N_3745,N_2679);
nand U4215 (N_4215,N_3086,N_2889);
nand U4216 (N_4216,N_3120,N_2777);
nand U4217 (N_4217,N_3801,N_2087);
nor U4218 (N_4218,N_3441,N_2774);
nand U4219 (N_4219,N_2295,N_3207);
nand U4220 (N_4220,N_2406,N_3250);
nor U4221 (N_4221,N_2572,N_2009);
and U4222 (N_4222,N_3075,N_3898);
nor U4223 (N_4223,N_3464,N_3668);
nand U4224 (N_4224,N_2256,N_2344);
and U4225 (N_4225,N_2658,N_2478);
nand U4226 (N_4226,N_2713,N_2667);
and U4227 (N_4227,N_3882,N_2054);
nand U4228 (N_4228,N_3591,N_3495);
xor U4229 (N_4229,N_3934,N_2465);
nand U4230 (N_4230,N_2240,N_2412);
nand U4231 (N_4231,N_2730,N_3703);
and U4232 (N_4232,N_3565,N_3492);
nor U4233 (N_4233,N_2722,N_3113);
nor U4234 (N_4234,N_2537,N_3405);
or U4235 (N_4235,N_3425,N_2641);
nor U4236 (N_4236,N_3303,N_3342);
nand U4237 (N_4237,N_3078,N_3989);
xnor U4238 (N_4238,N_3162,N_3160);
nor U4239 (N_4239,N_2786,N_2247);
nand U4240 (N_4240,N_3094,N_2994);
and U4241 (N_4241,N_3743,N_2444);
nor U4242 (N_4242,N_3460,N_2381);
or U4243 (N_4243,N_2375,N_3861);
or U4244 (N_4244,N_3427,N_2681);
nor U4245 (N_4245,N_2675,N_3732);
nor U4246 (N_4246,N_2328,N_3980);
or U4247 (N_4247,N_3180,N_2510);
or U4248 (N_4248,N_2285,N_3706);
and U4249 (N_4249,N_2895,N_3536);
nor U4250 (N_4250,N_3886,N_2476);
and U4251 (N_4251,N_2901,N_3284);
nand U4252 (N_4252,N_2066,N_3051);
nand U4253 (N_4253,N_3846,N_2735);
nand U4254 (N_4254,N_2776,N_2609);
and U4255 (N_4255,N_3131,N_3577);
nor U4256 (N_4256,N_3862,N_2359);
or U4257 (N_4257,N_3883,N_3187);
xor U4258 (N_4258,N_2787,N_2200);
and U4259 (N_4259,N_2785,N_2498);
and U4260 (N_4260,N_2961,N_2187);
and U4261 (N_4261,N_3483,N_2807);
xnor U4262 (N_4262,N_3374,N_3269);
and U4263 (N_4263,N_3652,N_2697);
and U4264 (N_4264,N_3293,N_2355);
and U4265 (N_4265,N_3519,N_3783);
xor U4266 (N_4266,N_2373,N_2676);
nor U4267 (N_4267,N_3261,N_3497);
and U4268 (N_4268,N_2170,N_2119);
nor U4269 (N_4269,N_3665,N_3514);
and U4270 (N_4270,N_2753,N_2588);
and U4271 (N_4271,N_2962,N_2733);
or U4272 (N_4272,N_2682,N_3320);
nor U4273 (N_4273,N_2567,N_2284);
nand U4274 (N_4274,N_2960,N_2540);
nand U4275 (N_4275,N_2436,N_3973);
nor U4276 (N_4276,N_3518,N_3189);
and U4277 (N_4277,N_3431,N_2802);
and U4278 (N_4278,N_2861,N_2864);
or U4279 (N_4279,N_2252,N_2625);
xnor U4280 (N_4280,N_3402,N_2292);
nand U4281 (N_4281,N_3926,N_3628);
or U4282 (N_4282,N_3522,N_2845);
xor U4283 (N_4283,N_2362,N_3977);
or U4284 (N_4284,N_2319,N_3426);
xnor U4285 (N_4285,N_3025,N_2907);
and U4286 (N_4286,N_3228,N_2352);
nand U4287 (N_4287,N_2558,N_3069);
xor U4288 (N_4288,N_3870,N_2286);
and U4289 (N_4289,N_3326,N_2665);
and U4290 (N_4290,N_3611,N_3029);
nand U4291 (N_4291,N_2499,N_3523);
and U4292 (N_4292,N_3438,N_2127);
nor U4293 (N_4293,N_2234,N_2978);
or U4294 (N_4294,N_2434,N_3863);
or U4295 (N_4295,N_2273,N_2557);
nor U4296 (N_4296,N_2300,N_2364);
xnor U4297 (N_4297,N_3620,N_2505);
and U4298 (N_4298,N_2219,N_3974);
nand U4299 (N_4299,N_3291,N_3716);
and U4300 (N_4300,N_2290,N_3362);
or U4301 (N_4301,N_3124,N_2578);
xor U4302 (N_4302,N_2397,N_2427);
or U4303 (N_4303,N_3908,N_3267);
nand U4304 (N_4304,N_3097,N_3968);
and U4305 (N_4305,N_3995,N_3820);
or U4306 (N_4306,N_3321,N_2827);
or U4307 (N_4307,N_3380,N_2789);
nor U4308 (N_4308,N_2237,N_2013);
nor U4309 (N_4309,N_2832,N_3171);
and U4310 (N_4310,N_2841,N_2663);
and U4311 (N_4311,N_2117,N_3309);
nor U4312 (N_4312,N_3393,N_3965);
nand U4313 (N_4313,N_3662,N_2162);
xor U4314 (N_4314,N_3256,N_3002);
xor U4315 (N_4315,N_3262,N_2349);
and U4316 (N_4316,N_3515,N_2335);
xor U4317 (N_4317,N_2859,N_2651);
or U4318 (N_4318,N_2372,N_2798);
and U4319 (N_4319,N_2850,N_2357);
or U4320 (N_4320,N_2655,N_2903);
nor U4321 (N_4321,N_2242,N_3808);
nor U4322 (N_4322,N_2898,N_3276);
nor U4323 (N_4323,N_3167,N_3243);
nor U4324 (N_4324,N_2339,N_3810);
and U4325 (N_4325,N_3388,N_2643);
and U4326 (N_4326,N_2153,N_3328);
or U4327 (N_4327,N_2928,N_2166);
and U4328 (N_4328,N_2261,N_3856);
nand U4329 (N_4329,N_3756,N_2002);
or U4330 (N_4330,N_3449,N_2915);
nand U4331 (N_4331,N_3245,N_2276);
and U4332 (N_4332,N_2194,N_2515);
nor U4333 (N_4333,N_3476,N_3661);
or U4334 (N_4334,N_2550,N_3586);
or U4335 (N_4335,N_2287,N_3603);
or U4336 (N_4336,N_3854,N_2825);
nor U4337 (N_4337,N_2317,N_2426);
nor U4338 (N_4338,N_3229,N_2093);
and U4339 (N_4339,N_3571,N_2418);
xnor U4340 (N_4340,N_2693,N_3887);
or U4341 (N_4341,N_3192,N_2561);
and U4342 (N_4342,N_3911,N_3108);
and U4343 (N_4343,N_3901,N_3480);
and U4344 (N_4344,N_2519,N_2851);
nor U4345 (N_4345,N_2938,N_2289);
nand U4346 (N_4346,N_3299,N_2884);
and U4347 (N_4347,N_3264,N_2435);
nor U4348 (N_4348,N_2044,N_3574);
nor U4349 (N_4349,N_2232,N_3560);
or U4350 (N_4350,N_3512,N_3485);
or U4351 (N_4351,N_3501,N_2378);
nand U4352 (N_4352,N_3457,N_2751);
or U4353 (N_4353,N_3036,N_2925);
nor U4354 (N_4354,N_2121,N_3695);
nand U4355 (N_4355,N_3691,N_3275);
or U4356 (N_4356,N_2099,N_2215);
nand U4357 (N_4357,N_2755,N_2268);
nor U4358 (N_4358,N_2405,N_3689);
nand U4359 (N_4359,N_2964,N_3742);
and U4360 (N_4360,N_3065,N_3606);
nor U4361 (N_4361,N_3082,N_2953);
nor U4362 (N_4362,N_2739,N_2486);
nor U4363 (N_4363,N_3723,N_3885);
or U4364 (N_4364,N_2251,N_3499);
and U4365 (N_4365,N_2035,N_3304);
nor U4366 (N_4366,N_2393,N_2196);
nor U4367 (N_4367,N_3027,N_2562);
and U4368 (N_4368,N_2535,N_3324);
nor U4369 (N_4369,N_3475,N_2674);
nor U4370 (N_4370,N_3592,N_3621);
nand U4371 (N_4371,N_2821,N_3637);
xor U4372 (N_4372,N_2525,N_2243);
nor U4373 (N_4373,N_3182,N_2900);
or U4374 (N_4374,N_3190,N_3230);
or U4375 (N_4375,N_2552,N_2582);
or U4376 (N_4376,N_2338,N_2188);
nand U4377 (N_4377,N_2782,N_2536);
nand U4378 (N_4378,N_2564,N_2226);
or U4379 (N_4379,N_2866,N_3379);
nand U4380 (N_4380,N_2593,N_2792);
nand U4381 (N_4381,N_3663,N_2151);
and U4382 (N_4382,N_2059,N_2298);
or U4383 (N_4383,N_3453,N_3616);
and U4384 (N_4384,N_2060,N_2784);
nand U4385 (N_4385,N_2533,N_3945);
nor U4386 (N_4386,N_3690,N_3848);
nor U4387 (N_4387,N_2098,N_3799);
nand U4388 (N_4388,N_2652,N_2779);
nor U4389 (N_4389,N_2229,N_2071);
or U4390 (N_4390,N_2993,N_3163);
or U4391 (N_4391,N_3068,N_3385);
or U4392 (N_4392,N_3066,N_3463);
nor U4393 (N_4393,N_2529,N_3140);
nand U4394 (N_4394,N_2047,N_3482);
nand U4395 (N_4395,N_3734,N_2115);
nor U4396 (N_4396,N_2718,N_2429);
or U4397 (N_4397,N_2145,N_3554);
xnor U4398 (N_4398,N_3822,N_3819);
and U4399 (N_4399,N_2580,N_2470);
or U4400 (N_4400,N_2086,N_2705);
nand U4401 (N_4401,N_3503,N_2936);
or U4402 (N_4402,N_3195,N_3138);
nand U4403 (N_4403,N_3997,N_2092);
nand U4404 (N_4404,N_3026,N_3337);
nor U4405 (N_4405,N_2968,N_3481);
nor U4406 (N_4406,N_2957,N_2635);
nand U4407 (N_4407,N_3880,N_3215);
nand U4408 (N_4408,N_3059,N_3817);
xor U4409 (N_4409,N_2568,N_2556);
nor U4410 (N_4410,N_3553,N_3580);
or U4411 (N_4411,N_3308,N_3145);
nand U4412 (N_4412,N_2692,N_3784);
nor U4413 (N_4413,N_3738,N_3409);
xnor U4414 (N_4414,N_2548,N_2384);
or U4415 (N_4415,N_2069,N_2877);
nor U4416 (N_4416,N_2809,N_2432);
nand U4417 (N_4417,N_2899,N_2576);
nand U4418 (N_4418,N_3057,N_3859);
nor U4419 (N_4419,N_2719,N_2523);
xnor U4420 (N_4420,N_3398,N_2105);
or U4421 (N_4421,N_2143,N_3594);
and U4422 (N_4422,N_2748,N_2669);
or U4423 (N_4423,N_3358,N_3660);
nor U4424 (N_4424,N_3110,N_3852);
and U4425 (N_4425,N_2758,N_2129);
and U4426 (N_4426,N_3608,N_3240);
and U4427 (N_4427,N_2150,N_2853);
nand U4428 (N_4428,N_2218,N_3546);
nand U4429 (N_4429,N_3248,N_2314);
and U4430 (N_4430,N_2538,N_2033);
and U4431 (N_4431,N_2504,N_3753);
nand U4432 (N_4432,N_2387,N_3352);
and U4433 (N_4433,N_2554,N_2383);
or U4434 (N_4434,N_2214,N_3170);
or U4435 (N_4435,N_2833,N_2664);
and U4436 (N_4436,N_3504,N_2138);
xor U4437 (N_4437,N_3985,N_2131);
nand U4438 (N_4438,N_2453,N_2297);
nand U4439 (N_4439,N_2046,N_3718);
xnor U4440 (N_4440,N_2645,N_3623);
and U4441 (N_4441,N_3414,N_3684);
and U4442 (N_4442,N_2163,N_2972);
or U4443 (N_4443,N_2947,N_3033);
nor U4444 (N_4444,N_3939,N_2600);
or U4445 (N_4445,N_2065,N_3517);
nand U4446 (N_4446,N_3824,N_2873);
or U4447 (N_4447,N_3360,N_3647);
nand U4448 (N_4448,N_3127,N_3252);
or U4449 (N_4449,N_2602,N_2495);
or U4450 (N_4450,N_2541,N_2490);
nand U4451 (N_4451,N_2591,N_2728);
xnor U4452 (N_4452,N_3419,N_2683);
or U4453 (N_4453,N_2061,N_3467);
nand U4454 (N_4454,N_3199,N_3528);
nor U4455 (N_4455,N_3158,N_2350);
nand U4456 (N_4456,N_2259,N_3930);
nand U4457 (N_4457,N_3255,N_3452);
nor U4458 (N_4458,N_2897,N_2103);
or U4459 (N_4459,N_3279,N_3836);
nand U4460 (N_4460,N_2459,N_3104);
and U4461 (N_4461,N_2530,N_3384);
nor U4462 (N_4462,N_2003,N_3376);
xor U4463 (N_4463,N_3907,N_2158);
xnor U4464 (N_4464,N_2213,N_3697);
xor U4465 (N_4465,N_3927,N_2817);
or U4466 (N_4466,N_2731,N_3077);
or U4467 (N_4467,N_2482,N_2999);
or U4468 (N_4468,N_2742,N_2759);
or U4469 (N_4469,N_2581,N_2911);
or U4470 (N_4470,N_2275,N_2241);
and U4471 (N_4471,N_2171,N_3012);
nand U4472 (N_4472,N_3835,N_2654);
or U4473 (N_4473,N_2207,N_3994);
or U4474 (N_4474,N_3566,N_3265);
or U4475 (N_4475,N_2020,N_2614);
and U4476 (N_4476,N_3727,N_3615);
and U4477 (N_4477,N_3975,N_2441);
or U4478 (N_4478,N_2695,N_2079);
or U4479 (N_4479,N_3128,N_2976);
nor U4480 (N_4480,N_2948,N_3224);
nor U4481 (N_4481,N_2878,N_2260);
nor U4482 (N_4482,N_3593,N_3246);
or U4483 (N_4483,N_3130,N_3339);
nand U4484 (N_4484,N_2544,N_2401);
or U4485 (N_4485,N_2039,N_3598);
nand U4486 (N_4486,N_3914,N_3563);
nor U4487 (N_4487,N_2167,N_3048);
nor U4488 (N_4488,N_2269,N_2800);
nor U4489 (N_4489,N_3540,N_3589);
or U4490 (N_4490,N_3842,N_2266);
nand U4491 (N_4491,N_2650,N_3857);
and U4492 (N_4492,N_3141,N_2660);
xor U4493 (N_4493,N_3607,N_3369);
and U4494 (N_4494,N_3655,N_2905);
nor U4495 (N_4495,N_2729,N_2570);
and U4496 (N_4496,N_2597,N_3448);
and U4497 (N_4497,N_3774,N_2246);
nor U4498 (N_4498,N_2771,N_2647);
nand U4499 (N_4499,N_2073,N_3496);
nand U4500 (N_4500,N_3399,N_3338);
nor U4501 (N_4501,N_3359,N_2483);
and U4502 (N_4502,N_3806,N_3585);
nor U4503 (N_4503,N_3760,N_3648);
or U4504 (N_4504,N_3349,N_3987);
and U4505 (N_4505,N_2311,N_3053);
and U4506 (N_4506,N_2710,N_2502);
nand U4507 (N_4507,N_2370,N_2734);
xnor U4508 (N_4508,N_2712,N_3103);
nor U4509 (N_4509,N_2892,N_3006);
or U4510 (N_4510,N_2123,N_3268);
nor U4511 (N_4511,N_3751,N_3387);
or U4512 (N_4512,N_2531,N_2209);
nand U4513 (N_4513,N_3642,N_2343);
and U4514 (N_4514,N_2340,N_2224);
or U4515 (N_4515,N_3306,N_2738);
nor U4516 (N_4516,N_2394,N_2090);
and U4517 (N_4517,N_2438,N_2831);
and U4518 (N_4518,N_2323,N_2174);
or U4519 (N_4519,N_2190,N_2575);
nor U4520 (N_4520,N_2354,N_2783);
nand U4521 (N_4521,N_2388,N_3368);
or U4522 (N_4522,N_2400,N_2463);
and U4523 (N_4523,N_2118,N_3855);
nand U4524 (N_4524,N_3708,N_2518);
nand U4525 (N_4525,N_3185,N_3490);
nand U4526 (N_4526,N_3831,N_2468);
nand U4527 (N_4527,N_3046,N_2428);
nor U4528 (N_4528,N_3825,N_2629);
and U4529 (N_4529,N_3294,N_2989);
nor U4530 (N_4530,N_3802,N_2684);
nor U4531 (N_4531,N_3666,N_3236);
or U4532 (N_4532,N_2439,N_3084);
nor U4533 (N_4533,N_2347,N_2670);
and U4534 (N_4534,N_3713,N_2649);
and U4535 (N_4535,N_2450,N_3114);
nand U4536 (N_4536,N_3361,N_3231);
or U4537 (N_4537,N_2780,N_3526);
nand U4538 (N_4538,N_3505,N_3670);
nor U4539 (N_4539,N_3302,N_3671);
nor U4540 (N_4540,N_2840,N_3052);
nand U4541 (N_4541,N_2371,N_2274);
nor U4542 (N_4542,N_2573,N_3263);
nor U4543 (N_4543,N_3461,N_3983);
or U4544 (N_4544,N_2822,N_2571);
nand U4545 (N_4545,N_2563,N_3730);
nor U4546 (N_4546,N_3209,N_3527);
or U4547 (N_4547,N_3430,N_3400);
and U4548 (N_4548,N_2640,N_3334);
or U4549 (N_4549,N_2981,N_2485);
nand U4550 (N_4550,N_3800,N_3986);
nand U4551 (N_4551,N_3137,N_2012);
or U4552 (N_4552,N_3809,N_2488);
xor U4553 (N_4553,N_2356,N_2305);
nand U4554 (N_4554,N_3552,N_3549);
nand U4555 (N_4555,N_3511,N_3198);
and U4556 (N_4556,N_3435,N_2790);
nand U4557 (N_4557,N_2648,N_3106);
or U4558 (N_4558,N_3455,N_3675);
and U4559 (N_4559,N_3305,N_3677);
nor U4560 (N_4560,N_2724,N_3280);
nand U4561 (N_4561,N_2967,N_2869);
nand U4562 (N_4562,N_2716,N_2599);
nor U4563 (N_4563,N_2560,N_3282);
nor U4564 (N_4564,N_2068,N_2206);
nand U4565 (N_4565,N_3404,N_2598);
nor U4566 (N_4566,N_3530,N_3123);
or U4567 (N_4567,N_3781,N_2431);
nand U4568 (N_4568,N_2132,N_2168);
or U4569 (N_4569,N_2493,N_2636);
or U4570 (N_4570,N_3401,N_2806);
or U4571 (N_4571,N_2584,N_2109);
or U4572 (N_4572,N_2032,N_2977);
and U4573 (N_4573,N_2070,N_2772);
and U4574 (N_4574,N_3984,N_2796);
nand U4575 (N_4575,N_3469,N_3823);
nor U4576 (N_4576,N_2395,N_2184);
xnor U4577 (N_4577,N_2097,N_2318);
nand U4578 (N_4578,N_3601,N_2152);
nand U4579 (N_4579,N_2927,N_2543);
nor U4580 (N_4580,N_3166,N_2404);
nand U4581 (N_4581,N_3645,N_2583);
xor U4582 (N_4582,N_2422,N_2084);
nor U4583 (N_4583,N_3558,N_2799);
nand U4584 (N_4584,N_3208,N_3218);
nor U4585 (N_4585,N_3323,N_3107);
nand U4586 (N_4586,N_3340,N_3964);
or U4587 (N_4587,N_3092,N_2180);
nand U4588 (N_4588,N_2191,N_2951);
and U4589 (N_4589,N_2933,N_2503);
or U4590 (N_4590,N_2081,N_3119);
and U4591 (N_4591,N_2623,N_2031);
nor U4592 (N_4592,N_3583,N_2306);
xor U4593 (N_4593,N_2834,N_2732);
and U4594 (N_4594,N_2826,N_2100);
nand U4595 (N_4595,N_2824,N_2916);
xor U4596 (N_4596,N_3257,N_3948);
nor U4597 (N_4597,N_3008,N_3249);
or U4598 (N_4598,N_2236,N_3640);
nand U4599 (N_4599,N_3590,N_2990);
and U4600 (N_4600,N_2159,N_2049);
nor U4601 (N_4601,N_3858,N_3949);
and U4602 (N_4602,N_3159,N_3890);
or U4603 (N_4603,N_3122,N_3919);
or U4604 (N_4604,N_3024,N_3237);
nor U4605 (N_4605,N_3843,N_2517);
nand U4606 (N_4606,N_2508,N_3588);
nor U4607 (N_4607,N_3135,N_2969);
or U4608 (N_4608,N_3277,N_2052);
nand U4609 (N_4609,N_3429,N_2858);
or U4610 (N_4610,N_3005,N_3833);
nand U4611 (N_4611,N_2496,N_3315);
nor U4612 (N_4612,N_2847,N_3154);
xor U4613 (N_4613,N_2042,N_2142);
or U4614 (N_4614,N_2756,N_3060);
nand U4615 (N_4615,N_2522,N_2855);
and U4616 (N_4616,N_2760,N_3351);
nor U4617 (N_4617,N_3715,N_3815);
xnor U4618 (N_4618,N_2257,N_3188);
nand U4619 (N_4619,N_3619,N_3010);
and U4620 (N_4620,N_3543,N_2937);
and U4621 (N_4621,N_2894,N_3929);
nand U4622 (N_4622,N_3978,N_2909);
nor U4623 (N_4623,N_3169,N_2106);
nor U4624 (N_4624,N_3776,N_3095);
or U4625 (N_4625,N_3803,N_2396);
or U4626 (N_4626,N_2425,N_3596);
nand U4627 (N_4627,N_3183,N_2420);
and U4628 (N_4628,N_3775,N_2096);
nor U4629 (N_4629,N_2018,N_3905);
and U4630 (N_4630,N_3089,N_2415);
and U4631 (N_4631,N_2291,N_2104);
nor U4632 (N_4632,N_3900,N_3150);
nor U4633 (N_4633,N_2932,N_2182);
xor U4634 (N_4634,N_3344,N_2342);
and U4635 (N_4635,N_2169,N_3869);
nand U4636 (N_4636,N_2919,N_2902);
and U4637 (N_4637,N_3981,N_3439);
nand U4638 (N_4638,N_3782,N_3396);
or U4639 (N_4639,N_3004,N_3763);
or U4640 (N_4640,N_2791,N_3191);
nor U4641 (N_4641,N_3904,N_3814);
nand U4642 (N_4642,N_3579,N_3408);
nor U4643 (N_4643,N_3686,N_3290);
nor U4644 (N_4644,N_3079,N_3437);
or U4645 (N_4645,N_2080,N_3804);
nand U4646 (N_4646,N_2638,N_3953);
and U4647 (N_4647,N_3423,N_3216);
or U4648 (N_4648,N_2939,N_2984);
or U4649 (N_4649,N_3746,N_2048);
or U4650 (N_4650,N_3381,N_3509);
nand U4651 (N_4651,N_3850,N_2315);
nand U4652 (N_4652,N_2612,N_2120);
or U4653 (N_4653,N_3332,N_2883);
nor U4654 (N_4654,N_3226,N_3478);
and U4655 (N_4655,N_3972,N_2860);
nor U4656 (N_4656,N_3726,N_3468);
nand U4657 (N_4657,N_3658,N_3285);
xor U4658 (N_4658,N_2559,N_3524);
nor U4659 (N_4659,N_2632,N_2333);
and U4660 (N_4660,N_2017,N_2494);
and U4661 (N_4661,N_3998,N_2334);
or U4662 (N_4662,N_2605,N_2891);
or U4663 (N_4663,N_3777,N_3759);
and U4664 (N_4664,N_3357,N_2233);
nand U4665 (N_4665,N_3287,N_2363);
and U4666 (N_4666,N_2849,N_2596);
nor U4667 (N_4667,N_3085,N_2808);
or U4668 (N_4668,N_3030,N_3074);
nand U4669 (N_4669,N_2154,N_3700);
or U4670 (N_4670,N_3545,N_2987);
and U4671 (N_4671,N_2836,N_2303);
or U4672 (N_4672,N_3028,N_3762);
nand U4673 (N_4673,N_3667,N_3205);
and U4674 (N_4674,N_2264,N_3550);
or U4675 (N_4675,N_3416,N_2248);
xnor U4676 (N_4676,N_2991,N_3731);
or U4677 (N_4677,N_2906,N_3470);
nor U4678 (N_4678,N_2380,N_3346);
or U4679 (N_4679,N_2077,N_2267);
nand U4680 (N_4680,N_2656,N_2793);
or U4681 (N_4681,N_2212,N_2763);
nand U4682 (N_4682,N_2377,N_3032);
or U4683 (N_4683,N_2195,N_3272);
nand U4684 (N_4684,N_3950,N_3371);
nor U4685 (N_4685,N_2382,N_3378);
and U4686 (N_4686,N_3656,N_2181);
nand U4687 (N_4687,N_3203,N_2114);
nand U4688 (N_4688,N_2471,N_3413);
nor U4689 (N_4689,N_3386,N_2986);
and U4690 (N_4690,N_2353,N_3924);
nor U4691 (N_4691,N_3971,N_3506);
and U4692 (N_4692,N_2551,N_2421);
nand U4693 (N_4693,N_3477,N_2781);
and U4694 (N_4694,N_2890,N_3682);
nand U4695 (N_4695,N_2668,N_3181);
nand U4696 (N_4696,N_3741,N_3795);
or U4697 (N_4697,N_2245,N_3319);
or U4698 (N_4698,N_2399,N_2795);
nor U4699 (N_4699,N_2040,N_2943);
nor U4700 (N_4700,N_3391,N_2464);
or U4701 (N_4701,N_3736,N_3000);
and U4702 (N_4702,N_3234,N_2622);
nand U4703 (N_4703,N_3832,N_3031);
or U4704 (N_4704,N_2574,N_3813);
and U4705 (N_4705,N_3347,N_3390);
nand U4706 (N_4706,N_2944,N_3355);
nand U4707 (N_4707,N_2700,N_3805);
and U4708 (N_4708,N_3988,N_2545);
and U4709 (N_4709,N_2424,N_2128);
and U4710 (N_4710,N_3221,N_3936);
and U4711 (N_4711,N_2041,N_2341);
nor U4712 (N_4712,N_2348,N_3176);
and U4713 (N_4713,N_2680,N_3724);
nor U4714 (N_4714,N_2155,N_3233);
nand U4715 (N_4715,N_2386,N_3445);
or U4716 (N_4716,N_3626,N_2920);
nand U4717 (N_4717,N_2133,N_3576);
and U4718 (N_4718,N_3109,N_3902);
nor U4719 (N_4719,N_3367,N_2992);
nand U4720 (N_4720,N_2417,N_2448);
or U4721 (N_4721,N_3714,N_2309);
nand U4722 (N_4722,N_3920,N_2762);
or U4723 (N_4723,N_2254,N_2176);
or U4724 (N_4724,N_2186,N_3450);
or U4725 (N_4725,N_3791,N_3692);
nand U4726 (N_4726,N_3129,N_2265);
nand U4727 (N_4727,N_3330,N_2365);
and U4728 (N_4728,N_3072,N_2351);
or U4729 (N_4729,N_2988,N_2050);
and U4730 (N_4730,N_2484,N_2569);
nor U4731 (N_4731,N_3765,N_3897);
or U4732 (N_4732,N_2628,N_3278);
and U4733 (N_4733,N_2816,N_2524);
or U4734 (N_4734,N_2281,N_3544);
nand U4735 (N_4735,N_3019,N_2457);
nand U4736 (N_4736,N_3578,N_2801);
nor U4737 (N_4737,N_3311,N_3541);
or U4738 (N_4738,N_3091,N_3432);
xnor U4739 (N_4739,N_3406,N_3389);
nand U4740 (N_4740,N_2862,N_2296);
nor U4741 (N_4741,N_3040,N_2161);
and U4742 (N_4742,N_2956,N_3173);
xor U4743 (N_4743,N_3206,N_3314);
or U4744 (N_4744,N_2045,N_2126);
or U4745 (N_4745,N_2908,N_3146);
or U4746 (N_4746,N_2872,N_3685);
nand U4747 (N_4747,N_2820,N_2262);
xnor U4748 (N_4748,N_2946,N_2630);
or U4749 (N_4749,N_2402,N_2996);
and U4750 (N_4750,N_3063,N_3764);
and U4751 (N_4751,N_2687,N_3121);
nand U4752 (N_4752,N_2604,N_2235);
or U4753 (N_4753,N_2283,N_3749);
nand U4754 (N_4754,N_3062,N_2479);
nand U4755 (N_4755,N_3155,N_2696);
xor U4756 (N_4756,N_2982,N_3719);
or U4757 (N_4757,N_2324,N_3595);
and U4758 (N_4758,N_3102,N_3382);
and U4759 (N_4759,N_2812,N_2750);
nand U4760 (N_4760,N_2838,N_3373);
nand U4761 (N_4761,N_2965,N_3829);
nor U4762 (N_4762,N_3925,N_3235);
and U4763 (N_4763,N_2691,N_3826);
nor U4764 (N_4764,N_2038,N_2139);
or U4765 (N_4765,N_3710,N_2757);
nor U4766 (N_4766,N_2199,N_3440);
and U4767 (N_4767,N_2116,N_3271);
nand U4768 (N_4768,N_2918,N_3087);
nand U4769 (N_4769,N_3153,N_2293);
nor U4770 (N_4770,N_3487,N_2815);
nor U4771 (N_4771,N_2910,N_3587);
nand U4772 (N_4772,N_3365,N_3999);
and U4773 (N_4773,N_2089,N_3990);
and U4774 (N_4774,N_2102,N_3343);
or U4775 (N_4775,N_2764,N_2481);
xnor U4776 (N_4776,N_3175,N_2244);
xnor U4777 (N_4777,N_2288,N_2221);
nor U4778 (N_4778,N_2316,N_3111);
or U4779 (N_4779,N_2385,N_3569);
nor U4780 (N_4780,N_3301,N_2403);
nand U4781 (N_4781,N_2715,N_2973);
or U4782 (N_4782,N_3720,N_2617);
and U4783 (N_4783,N_3793,N_3016);
nand U4784 (N_4784,N_3274,N_2307);
and U4785 (N_4785,N_2514,N_3172);
or U4786 (N_4786,N_2666,N_2620);
nand U4787 (N_4787,N_3067,N_3184);
and U4788 (N_4788,N_2320,N_3884);
nor U4789 (N_4789,N_2959,N_2413);
xor U4790 (N_4790,N_2754,N_3755);
xor U4791 (N_4791,N_2067,N_3098);
nand U4792 (N_4792,N_3201,N_2282);
or U4793 (N_4793,N_2346,N_3581);
nand U4794 (N_4794,N_3446,N_2497);
or U4795 (N_4795,N_3548,N_3567);
nor U4796 (N_4796,N_2874,N_2208);
nor U4797 (N_4797,N_2430,N_3599);
and U4798 (N_4798,N_2072,N_3147);
and U4799 (N_4799,N_2941,N_2513);
and U4800 (N_4800,N_2345,N_2998);
or U4801 (N_4801,N_3568,N_3296);
nor U4802 (N_4802,N_3353,N_2442);
or U4803 (N_4803,N_3350,N_2057);
nand U4804 (N_4804,N_2337,N_2006);
xor U4805 (N_4805,N_3116,N_2440);
or U4806 (N_4806,N_3238,N_2461);
nand U4807 (N_4807,N_3993,N_3298);
xor U4808 (N_4808,N_2590,N_2702);
nand U4809 (N_4809,N_3281,N_3115);
nor U4810 (N_4810,N_3502,N_2788);
nand U4811 (N_4811,N_2410,N_3223);
xor U4812 (N_4812,N_2509,N_2491);
nand U4813 (N_4813,N_3876,N_3664);
nor U4814 (N_4814,N_3827,N_3712);
and U4815 (N_4815,N_3694,N_2492);
xor U4816 (N_4816,N_3366,N_3042);
or U4817 (N_4817,N_2942,N_3679);
and U4818 (N_4818,N_3018,N_3752);
nor U4819 (N_4819,N_3488,N_3991);
xnor U4820 (N_4820,N_3099,N_2974);
and U4821 (N_4821,N_3638,N_3657);
xnor U4822 (N_4822,N_2856,N_3650);
nand U4823 (N_4823,N_2443,N_2613);
or U4824 (N_4824,N_3754,N_2376);
nor U4825 (N_4825,N_3797,N_3792);
nor U4826 (N_4826,N_3020,N_3411);
nand U4827 (N_4827,N_3729,N_2313);
nor U4828 (N_4828,N_3038,N_3867);
nand U4829 (N_4829,N_3080,N_3931);
and U4830 (N_4830,N_3954,N_2714);
nand U4831 (N_4831,N_3466,N_3056);
nand U4832 (N_4832,N_3564,N_2539);
or U4833 (N_4833,N_2528,N_2270);
or U4834 (N_4834,N_3200,N_2835);
nand U4835 (N_4835,N_2740,N_3009);
or U4836 (N_4836,N_2390,N_3771);
nand U4837 (N_4837,N_3966,N_2456);
or U4838 (N_4838,N_2619,N_2507);
and U4839 (N_4839,N_3253,N_2433);
or U4840 (N_4840,N_2144,N_2474);
or U4841 (N_4841,N_2923,N_2220);
nand U4842 (N_4842,N_3472,N_3659);
xor U4843 (N_4843,N_2423,N_3933);
and U4844 (N_4844,N_2185,N_3951);
and U4845 (N_4845,N_3117,N_2368);
nand U4846 (N_4846,N_2608,N_2985);
nand U4847 (N_4847,N_2475,N_2445);
nand U4848 (N_4848,N_2419,N_2963);
and U4849 (N_4849,N_3007,N_3112);
nor U4850 (N_4850,N_2258,N_3551);
or U4851 (N_4851,N_2694,N_2707);
nand U4852 (N_4852,N_3133,N_3830);
nand U4853 (N_4853,N_3161,N_3037);
nand U4854 (N_4854,N_3156,N_3064);
xor U4855 (N_4855,N_3017,N_2437);
xnor U4856 (N_4856,N_2865,N_3417);
and U4857 (N_4857,N_3625,N_3702);
and U4858 (N_4858,N_3356,N_3377);
or U4859 (N_4859,N_3979,N_3969);
nor U4860 (N_4860,N_2037,N_3144);
or U4861 (N_4861,N_2172,N_3101);
nand U4862 (N_4862,N_3559,N_3992);
nand U4863 (N_4863,N_3050,N_2301);
xor U4864 (N_4864,N_2810,N_2745);
and U4865 (N_4865,N_3970,N_2122);
nor U4866 (N_4866,N_3597,N_2360);
and U4867 (N_4867,N_2392,N_3561);
nand U4868 (N_4868,N_3491,N_2703);
nand U4869 (N_4869,N_2749,N_3944);
and U4870 (N_4870,N_3605,N_2255);
nor U4871 (N_4871,N_2058,N_2074);
nand U4872 (N_4872,N_3943,N_2107);
or U4873 (N_4873,N_3105,N_3600);
nor U4874 (N_4874,N_3617,N_2888);
and U4875 (N_4875,N_3773,N_3958);
nor U4876 (N_4876,N_3329,N_2690);
or U4877 (N_4877,N_3165,N_3627);
and U4878 (N_4878,N_3058,N_3035);
xor U4879 (N_4879,N_3270,N_3300);
xnor U4880 (N_4880,N_3877,N_2101);
nand U4881 (N_4881,N_3917,N_3254);
and U4882 (N_4882,N_2819,N_3193);
or U4883 (N_4883,N_3489,N_2134);
or U4884 (N_4884,N_2688,N_3484);
nor U4885 (N_4885,N_2601,N_3061);
nor U4886 (N_4886,N_3629,N_3266);
and U4887 (N_4887,N_3219,N_2642);
nor U4888 (N_4888,N_2805,N_2140);
or U4889 (N_4889,N_2391,N_2466);
xor U4890 (N_4890,N_3873,N_2627);
or U4891 (N_4891,N_2062,N_3899);
nand U4892 (N_4892,N_3015,N_2088);
nand U4893 (N_4893,N_2205,N_3244);
nand U4894 (N_4894,N_3454,N_3283);
and U4895 (N_4895,N_2954,N_3704);
xnor U4896 (N_4896,N_2875,N_2366);
and U4897 (N_4897,N_3853,N_3940);
nand U4898 (N_4898,N_3962,N_2863);
and U4899 (N_4899,N_2225,N_2330);
xor U4900 (N_4900,N_2709,N_2374);
nor U4901 (N_4901,N_3996,N_3370);
nand U4902 (N_4902,N_2160,N_2566);
or U4903 (N_4903,N_2904,N_3896);
and U4904 (N_4904,N_2462,N_3612);
or U4905 (N_4905,N_2487,N_3213);
xnor U4906 (N_4906,N_2512,N_3982);
and U4907 (N_4907,N_2165,N_3636);
or U4908 (N_4908,N_2881,N_3942);
nor U4909 (N_4909,N_2876,N_2811);
and U4910 (N_4910,N_2294,N_3459);
or U4911 (N_4911,N_3957,N_2577);
xnor U4912 (N_4912,N_2329,N_3618);
nand U4913 (N_4913,N_2657,N_3174);
nor U4914 (N_4914,N_3956,N_2473);
nor U4915 (N_4915,N_2843,N_2022);
nand U4916 (N_4916,N_2183,N_3821);
and U4917 (N_4917,N_2164,N_2725);
or U4918 (N_4918,N_3186,N_3834);
or U4919 (N_4919,N_3680,N_2686);
xor U4920 (N_4920,N_2917,N_3874);
and U4921 (N_4921,N_2979,N_2995);
or U4922 (N_4922,N_3840,N_2379);
nor U4923 (N_4923,N_2752,N_2761);
and U4924 (N_4924,N_3375,N_2016);
or U4925 (N_4925,N_3047,N_3812);
nand U4926 (N_4926,N_2146,N_3811);
and U4927 (N_4927,N_3698,N_3222);
nand U4928 (N_4928,N_3247,N_2501);
or U4929 (N_4929,N_2778,N_2312);
nand U4930 (N_4930,N_2673,N_2506);
or U4931 (N_4931,N_3556,N_3584);
or U4932 (N_4932,N_2689,N_2621);
or U4933 (N_4933,N_3910,N_2914);
or U4934 (N_4934,N_3196,N_2711);
and U4935 (N_4935,N_3602,N_2765);
and U4936 (N_4936,N_3043,N_2955);
and U4937 (N_4937,N_3322,N_3582);
nand U4938 (N_4938,N_3761,N_3073);
nor U4939 (N_4939,N_2534,N_3828);
nor U4940 (N_4940,N_3286,N_3767);
and U4941 (N_4941,N_3959,N_3421);
or U4942 (N_4942,N_2063,N_3787);
nand U4943 (N_4943,N_3428,N_2527);
or U4944 (N_4944,N_3780,N_3779);
or U4945 (N_4945,N_2019,N_3071);
xnor U4946 (N_4946,N_3336,N_2055);
nand U4947 (N_4947,N_2028,N_3918);
nor U4948 (N_4948,N_2842,N_3845);
or U4949 (N_4949,N_3866,N_2661);
nand U4950 (N_4950,N_2727,N_3132);
nor U4951 (N_4951,N_3451,N_2111);
and U4952 (N_4952,N_2231,N_3711);
or U4953 (N_4953,N_2532,N_3295);
or U4954 (N_4954,N_3952,N_3912);
nand U4955 (N_4955,N_2610,N_2685);
or U4956 (N_4956,N_2024,N_2797);
nor U4957 (N_4957,N_2277,N_3125);
nor U4958 (N_4958,N_3202,N_3297);
and U4959 (N_4959,N_2409,N_3614);
nand U4960 (N_4960,N_2912,N_2454);
nor U4961 (N_4961,N_3868,N_2358);
nor U4962 (N_4962,N_2216,N_2701);
nor U4963 (N_4963,N_3906,N_2157);
xor U4964 (N_4964,N_3837,N_2108);
or U4965 (N_4965,N_3785,N_2280);
xnor U4966 (N_4966,N_2945,N_2768);
nand U4967 (N_4967,N_2271,N_2708);
or U4968 (N_4968,N_3179,N_2585);
or U4969 (N_4969,N_3076,N_2549);
or U4970 (N_4970,N_3790,N_3318);
and U4971 (N_4971,N_3534,N_2389);
nand U4972 (N_4972,N_3474,N_2555);
nand U4973 (N_4973,N_3932,N_3444);
nor U4974 (N_4974,N_3860,N_2746);
nand U4975 (N_4975,N_3654,N_3242);
and U4976 (N_4976,N_3307,N_2489);
xnor U4977 (N_4977,N_2336,N_3735);
xor U4978 (N_4978,N_2736,N_2659);
and U4979 (N_4979,N_3913,N_2603);
nor U4980 (N_4980,N_3088,N_2210);
or U4981 (N_4981,N_2929,N_3498);
or U4982 (N_4982,N_3239,N_3143);
and U4983 (N_4983,N_2460,N_3021);
xor U4984 (N_4984,N_3210,N_3879);
and U4985 (N_4985,N_3757,N_3961);
nand U4986 (N_4986,N_3653,N_2818);
or U4987 (N_4987,N_2014,N_3335);
nor U4988 (N_4988,N_3090,N_3157);
nand U4989 (N_4989,N_3941,N_3212);
or U4990 (N_4990,N_3507,N_2149);
or U4991 (N_4991,N_2813,N_3260);
nor U4992 (N_4992,N_3865,N_3739);
nor U4993 (N_4993,N_3289,N_3938);
nand U4994 (N_4994,N_2156,N_2770);
nor U4995 (N_4995,N_2704,N_3609);
and U4996 (N_4996,N_3928,N_3139);
nor U4997 (N_4997,N_3570,N_3878);
or U4998 (N_4998,N_3055,N_2322);
nor U4999 (N_4999,N_2952,N_3325);
and U5000 (N_5000,N_2652,N_3412);
xnor U5001 (N_5001,N_3992,N_2956);
nand U5002 (N_5002,N_3598,N_2872);
and U5003 (N_5003,N_3776,N_3997);
or U5004 (N_5004,N_2053,N_3134);
nand U5005 (N_5005,N_2332,N_3466);
nor U5006 (N_5006,N_3143,N_2143);
nand U5007 (N_5007,N_2602,N_3064);
or U5008 (N_5008,N_3772,N_3728);
nor U5009 (N_5009,N_2001,N_3698);
or U5010 (N_5010,N_2203,N_2477);
nor U5011 (N_5011,N_3530,N_2898);
nand U5012 (N_5012,N_2750,N_2879);
or U5013 (N_5013,N_3528,N_3696);
or U5014 (N_5014,N_3691,N_3619);
nor U5015 (N_5015,N_2383,N_3179);
and U5016 (N_5016,N_2132,N_3348);
nand U5017 (N_5017,N_3417,N_2586);
nand U5018 (N_5018,N_3481,N_3873);
xor U5019 (N_5019,N_2761,N_2601);
nor U5020 (N_5020,N_3559,N_3176);
and U5021 (N_5021,N_3775,N_3888);
nor U5022 (N_5022,N_2407,N_2793);
xnor U5023 (N_5023,N_2167,N_3389);
and U5024 (N_5024,N_3415,N_3893);
xor U5025 (N_5025,N_3019,N_2828);
nand U5026 (N_5026,N_2777,N_3610);
and U5027 (N_5027,N_3454,N_2768);
xor U5028 (N_5028,N_3939,N_2251);
nor U5029 (N_5029,N_2496,N_2730);
or U5030 (N_5030,N_3783,N_2620);
nor U5031 (N_5031,N_2863,N_3741);
nand U5032 (N_5032,N_3285,N_2581);
nand U5033 (N_5033,N_2993,N_2986);
or U5034 (N_5034,N_3695,N_2161);
nand U5035 (N_5035,N_3997,N_3221);
or U5036 (N_5036,N_2154,N_2171);
nand U5037 (N_5037,N_3425,N_2219);
nor U5038 (N_5038,N_2179,N_2224);
and U5039 (N_5039,N_2555,N_3351);
xnor U5040 (N_5040,N_2998,N_2477);
or U5041 (N_5041,N_3485,N_2116);
nand U5042 (N_5042,N_2157,N_2958);
and U5043 (N_5043,N_2997,N_3230);
and U5044 (N_5044,N_3058,N_2346);
nand U5045 (N_5045,N_3671,N_3407);
or U5046 (N_5046,N_3905,N_2833);
nor U5047 (N_5047,N_3365,N_2848);
nor U5048 (N_5048,N_3749,N_2867);
nor U5049 (N_5049,N_2211,N_3775);
nand U5050 (N_5050,N_3979,N_3468);
and U5051 (N_5051,N_3127,N_3095);
nor U5052 (N_5052,N_2208,N_3792);
or U5053 (N_5053,N_2895,N_3810);
nand U5054 (N_5054,N_3598,N_2153);
or U5055 (N_5055,N_2049,N_2860);
nor U5056 (N_5056,N_3049,N_2418);
nand U5057 (N_5057,N_3529,N_3726);
or U5058 (N_5058,N_2005,N_3760);
nor U5059 (N_5059,N_2964,N_3948);
nor U5060 (N_5060,N_3018,N_3899);
nor U5061 (N_5061,N_2449,N_3551);
or U5062 (N_5062,N_3830,N_3402);
nand U5063 (N_5063,N_2711,N_2437);
nor U5064 (N_5064,N_2931,N_2571);
or U5065 (N_5065,N_2626,N_2321);
nand U5066 (N_5066,N_3264,N_3311);
or U5067 (N_5067,N_2315,N_2531);
nor U5068 (N_5068,N_3839,N_2626);
and U5069 (N_5069,N_3610,N_3352);
or U5070 (N_5070,N_3199,N_2799);
nor U5071 (N_5071,N_3812,N_3973);
or U5072 (N_5072,N_3949,N_3511);
or U5073 (N_5073,N_3510,N_2011);
nand U5074 (N_5074,N_2241,N_2258);
and U5075 (N_5075,N_2700,N_2159);
and U5076 (N_5076,N_2291,N_2250);
and U5077 (N_5077,N_3213,N_2591);
and U5078 (N_5078,N_2271,N_3303);
xor U5079 (N_5079,N_2004,N_2744);
nand U5080 (N_5080,N_3822,N_3309);
or U5081 (N_5081,N_2236,N_3442);
or U5082 (N_5082,N_2687,N_2635);
and U5083 (N_5083,N_3709,N_2422);
nand U5084 (N_5084,N_2473,N_2777);
or U5085 (N_5085,N_2611,N_3230);
and U5086 (N_5086,N_3609,N_3788);
nor U5087 (N_5087,N_3984,N_2358);
nand U5088 (N_5088,N_2586,N_2826);
and U5089 (N_5089,N_3297,N_3365);
and U5090 (N_5090,N_3328,N_2030);
or U5091 (N_5091,N_3796,N_2637);
nor U5092 (N_5092,N_3631,N_2286);
and U5093 (N_5093,N_2364,N_2722);
and U5094 (N_5094,N_2219,N_3018);
xor U5095 (N_5095,N_2391,N_3796);
nor U5096 (N_5096,N_2442,N_2119);
and U5097 (N_5097,N_2293,N_2062);
nor U5098 (N_5098,N_2617,N_3705);
xor U5099 (N_5099,N_3757,N_2386);
xor U5100 (N_5100,N_2272,N_2478);
nand U5101 (N_5101,N_3589,N_2888);
nor U5102 (N_5102,N_3592,N_3107);
or U5103 (N_5103,N_3125,N_2532);
nor U5104 (N_5104,N_3082,N_2310);
or U5105 (N_5105,N_3668,N_2509);
and U5106 (N_5106,N_3947,N_3446);
or U5107 (N_5107,N_3665,N_3843);
or U5108 (N_5108,N_3136,N_3112);
xnor U5109 (N_5109,N_2032,N_2742);
or U5110 (N_5110,N_2473,N_2249);
or U5111 (N_5111,N_3089,N_3184);
xnor U5112 (N_5112,N_3365,N_3926);
or U5113 (N_5113,N_2147,N_2634);
nand U5114 (N_5114,N_2419,N_2074);
nor U5115 (N_5115,N_2884,N_2885);
nand U5116 (N_5116,N_2095,N_2384);
nand U5117 (N_5117,N_2566,N_3857);
or U5118 (N_5118,N_2669,N_3558);
nor U5119 (N_5119,N_2037,N_3133);
nor U5120 (N_5120,N_2447,N_2251);
and U5121 (N_5121,N_2689,N_2669);
or U5122 (N_5122,N_2144,N_2399);
nor U5123 (N_5123,N_2134,N_3605);
nand U5124 (N_5124,N_3097,N_2501);
and U5125 (N_5125,N_2177,N_2624);
nand U5126 (N_5126,N_3939,N_2458);
nor U5127 (N_5127,N_3272,N_3035);
nor U5128 (N_5128,N_2029,N_3126);
nor U5129 (N_5129,N_2261,N_2770);
or U5130 (N_5130,N_2808,N_2405);
xor U5131 (N_5131,N_2977,N_2632);
nand U5132 (N_5132,N_3454,N_3779);
and U5133 (N_5133,N_2469,N_2621);
and U5134 (N_5134,N_2034,N_2118);
nor U5135 (N_5135,N_3527,N_2873);
xnor U5136 (N_5136,N_2410,N_2245);
or U5137 (N_5137,N_2969,N_3343);
or U5138 (N_5138,N_2406,N_2851);
and U5139 (N_5139,N_2054,N_2754);
nor U5140 (N_5140,N_3736,N_2007);
nor U5141 (N_5141,N_3487,N_2414);
or U5142 (N_5142,N_3402,N_2829);
nand U5143 (N_5143,N_2284,N_2815);
nand U5144 (N_5144,N_3331,N_3658);
or U5145 (N_5145,N_3945,N_3829);
nor U5146 (N_5146,N_3752,N_3266);
and U5147 (N_5147,N_2462,N_2602);
nand U5148 (N_5148,N_3054,N_2489);
and U5149 (N_5149,N_2606,N_3897);
nand U5150 (N_5150,N_3616,N_3142);
and U5151 (N_5151,N_3000,N_2171);
xor U5152 (N_5152,N_3505,N_2002);
nand U5153 (N_5153,N_2506,N_3900);
or U5154 (N_5154,N_2486,N_2345);
nand U5155 (N_5155,N_2996,N_2083);
nor U5156 (N_5156,N_3197,N_2218);
or U5157 (N_5157,N_3506,N_3074);
nand U5158 (N_5158,N_3794,N_3594);
nand U5159 (N_5159,N_3375,N_3853);
nand U5160 (N_5160,N_2716,N_3888);
nand U5161 (N_5161,N_3680,N_3639);
and U5162 (N_5162,N_2199,N_3056);
xor U5163 (N_5163,N_2432,N_2706);
or U5164 (N_5164,N_2645,N_2567);
or U5165 (N_5165,N_2917,N_3862);
and U5166 (N_5166,N_2055,N_3935);
xnor U5167 (N_5167,N_3051,N_3953);
nand U5168 (N_5168,N_3987,N_2232);
nand U5169 (N_5169,N_3067,N_3751);
nor U5170 (N_5170,N_3388,N_2454);
and U5171 (N_5171,N_3189,N_3366);
nor U5172 (N_5172,N_2014,N_2879);
and U5173 (N_5173,N_2942,N_3075);
nor U5174 (N_5174,N_3998,N_2734);
and U5175 (N_5175,N_3476,N_2044);
and U5176 (N_5176,N_3711,N_3015);
or U5177 (N_5177,N_2650,N_2169);
and U5178 (N_5178,N_3731,N_2555);
nand U5179 (N_5179,N_2705,N_2579);
and U5180 (N_5180,N_2620,N_3514);
xnor U5181 (N_5181,N_2435,N_2353);
nand U5182 (N_5182,N_3457,N_3099);
xor U5183 (N_5183,N_2828,N_3062);
nand U5184 (N_5184,N_2331,N_2435);
or U5185 (N_5185,N_2246,N_2034);
or U5186 (N_5186,N_3379,N_3544);
nand U5187 (N_5187,N_3161,N_2291);
or U5188 (N_5188,N_2891,N_3845);
nand U5189 (N_5189,N_2061,N_2457);
nor U5190 (N_5190,N_3617,N_3611);
and U5191 (N_5191,N_2040,N_2065);
or U5192 (N_5192,N_3693,N_2594);
and U5193 (N_5193,N_2587,N_2309);
or U5194 (N_5194,N_3849,N_2395);
xor U5195 (N_5195,N_2113,N_2338);
nor U5196 (N_5196,N_2126,N_3569);
or U5197 (N_5197,N_2284,N_3165);
nand U5198 (N_5198,N_2812,N_3055);
nor U5199 (N_5199,N_2812,N_3227);
xnor U5200 (N_5200,N_3715,N_2179);
nor U5201 (N_5201,N_2519,N_2890);
nand U5202 (N_5202,N_2626,N_2699);
or U5203 (N_5203,N_3168,N_2574);
nand U5204 (N_5204,N_3734,N_3511);
and U5205 (N_5205,N_3671,N_3767);
and U5206 (N_5206,N_2924,N_3550);
and U5207 (N_5207,N_2788,N_3271);
nand U5208 (N_5208,N_2169,N_3817);
and U5209 (N_5209,N_2941,N_2307);
or U5210 (N_5210,N_2670,N_3596);
nor U5211 (N_5211,N_3328,N_2290);
and U5212 (N_5212,N_3281,N_3514);
nand U5213 (N_5213,N_2108,N_2624);
and U5214 (N_5214,N_3416,N_3290);
or U5215 (N_5215,N_3955,N_2170);
or U5216 (N_5216,N_2679,N_2488);
or U5217 (N_5217,N_3679,N_3431);
nand U5218 (N_5218,N_2723,N_3564);
and U5219 (N_5219,N_3904,N_2220);
and U5220 (N_5220,N_2350,N_2183);
or U5221 (N_5221,N_3889,N_2648);
and U5222 (N_5222,N_2692,N_3162);
xor U5223 (N_5223,N_3441,N_3643);
nand U5224 (N_5224,N_2384,N_2683);
and U5225 (N_5225,N_2718,N_3297);
nor U5226 (N_5226,N_3748,N_2470);
nand U5227 (N_5227,N_2580,N_2781);
and U5228 (N_5228,N_3205,N_2991);
and U5229 (N_5229,N_2366,N_3045);
nand U5230 (N_5230,N_2701,N_3351);
or U5231 (N_5231,N_3202,N_3548);
nand U5232 (N_5232,N_2558,N_3278);
or U5233 (N_5233,N_3008,N_2506);
nand U5234 (N_5234,N_3162,N_2409);
and U5235 (N_5235,N_2469,N_3961);
and U5236 (N_5236,N_2450,N_2658);
nand U5237 (N_5237,N_3006,N_2073);
xnor U5238 (N_5238,N_2748,N_3895);
nor U5239 (N_5239,N_2772,N_3599);
nand U5240 (N_5240,N_3189,N_2236);
nor U5241 (N_5241,N_3040,N_2794);
nor U5242 (N_5242,N_3444,N_3165);
or U5243 (N_5243,N_2914,N_3768);
nand U5244 (N_5244,N_3861,N_3084);
nand U5245 (N_5245,N_3633,N_2979);
or U5246 (N_5246,N_2262,N_2982);
xnor U5247 (N_5247,N_3834,N_3940);
nand U5248 (N_5248,N_2671,N_3614);
and U5249 (N_5249,N_3046,N_3918);
or U5250 (N_5250,N_2871,N_3249);
or U5251 (N_5251,N_2354,N_2915);
and U5252 (N_5252,N_2053,N_3983);
nand U5253 (N_5253,N_3230,N_3104);
nor U5254 (N_5254,N_3229,N_3174);
nor U5255 (N_5255,N_3068,N_2463);
nor U5256 (N_5256,N_2315,N_2283);
nand U5257 (N_5257,N_3810,N_3212);
xnor U5258 (N_5258,N_2746,N_3333);
or U5259 (N_5259,N_3538,N_2466);
and U5260 (N_5260,N_3676,N_2411);
nand U5261 (N_5261,N_2692,N_2518);
xor U5262 (N_5262,N_3222,N_3797);
nand U5263 (N_5263,N_2292,N_3429);
nor U5264 (N_5264,N_3305,N_3795);
or U5265 (N_5265,N_3923,N_3698);
and U5266 (N_5266,N_3510,N_2079);
nor U5267 (N_5267,N_2534,N_3859);
nand U5268 (N_5268,N_2086,N_3584);
or U5269 (N_5269,N_2692,N_2032);
nand U5270 (N_5270,N_2400,N_3144);
and U5271 (N_5271,N_2733,N_3617);
nand U5272 (N_5272,N_2203,N_2570);
nand U5273 (N_5273,N_2856,N_2419);
nand U5274 (N_5274,N_2793,N_3979);
or U5275 (N_5275,N_2082,N_2784);
or U5276 (N_5276,N_2585,N_2311);
nor U5277 (N_5277,N_2945,N_3680);
xnor U5278 (N_5278,N_3725,N_2828);
nor U5279 (N_5279,N_3009,N_2478);
nand U5280 (N_5280,N_2782,N_3583);
and U5281 (N_5281,N_3032,N_3320);
nand U5282 (N_5282,N_3150,N_3330);
nand U5283 (N_5283,N_3962,N_2767);
and U5284 (N_5284,N_2212,N_2640);
nand U5285 (N_5285,N_2871,N_3382);
or U5286 (N_5286,N_2869,N_3802);
and U5287 (N_5287,N_3407,N_3762);
xnor U5288 (N_5288,N_3981,N_2072);
and U5289 (N_5289,N_2938,N_2192);
or U5290 (N_5290,N_3282,N_3843);
nor U5291 (N_5291,N_2720,N_3084);
and U5292 (N_5292,N_3213,N_2295);
and U5293 (N_5293,N_3079,N_2343);
xor U5294 (N_5294,N_2047,N_2242);
and U5295 (N_5295,N_2009,N_3851);
and U5296 (N_5296,N_3566,N_2895);
or U5297 (N_5297,N_2558,N_3509);
and U5298 (N_5298,N_2568,N_3355);
or U5299 (N_5299,N_2929,N_3369);
xor U5300 (N_5300,N_2063,N_2571);
xor U5301 (N_5301,N_2127,N_2558);
xor U5302 (N_5302,N_2011,N_3728);
or U5303 (N_5303,N_3352,N_2263);
xor U5304 (N_5304,N_3255,N_2702);
or U5305 (N_5305,N_2854,N_2005);
nand U5306 (N_5306,N_2552,N_3887);
xor U5307 (N_5307,N_3854,N_2558);
or U5308 (N_5308,N_2657,N_2547);
nor U5309 (N_5309,N_3582,N_3268);
nand U5310 (N_5310,N_3377,N_2334);
nand U5311 (N_5311,N_2589,N_2337);
or U5312 (N_5312,N_3575,N_3625);
nor U5313 (N_5313,N_3376,N_2794);
nand U5314 (N_5314,N_3759,N_2987);
and U5315 (N_5315,N_2538,N_2397);
nand U5316 (N_5316,N_3624,N_3523);
and U5317 (N_5317,N_2340,N_2538);
or U5318 (N_5318,N_2282,N_3387);
or U5319 (N_5319,N_3291,N_2238);
nand U5320 (N_5320,N_2705,N_3886);
xnor U5321 (N_5321,N_3825,N_2787);
and U5322 (N_5322,N_2765,N_3316);
or U5323 (N_5323,N_2304,N_2518);
nor U5324 (N_5324,N_2513,N_3126);
and U5325 (N_5325,N_2118,N_3874);
nor U5326 (N_5326,N_2155,N_2494);
nand U5327 (N_5327,N_3991,N_3438);
nor U5328 (N_5328,N_2185,N_2920);
xnor U5329 (N_5329,N_3743,N_2547);
nand U5330 (N_5330,N_3077,N_2091);
nand U5331 (N_5331,N_3783,N_2658);
and U5332 (N_5332,N_2125,N_2595);
or U5333 (N_5333,N_3266,N_2860);
or U5334 (N_5334,N_2329,N_2628);
nor U5335 (N_5335,N_3067,N_3504);
nand U5336 (N_5336,N_2879,N_2381);
nand U5337 (N_5337,N_2566,N_2222);
or U5338 (N_5338,N_2934,N_3283);
or U5339 (N_5339,N_3457,N_3790);
and U5340 (N_5340,N_3637,N_3171);
nor U5341 (N_5341,N_3495,N_3349);
nand U5342 (N_5342,N_2867,N_2511);
nor U5343 (N_5343,N_2875,N_3898);
nand U5344 (N_5344,N_2541,N_2352);
nand U5345 (N_5345,N_3943,N_3959);
or U5346 (N_5346,N_3535,N_3570);
nand U5347 (N_5347,N_3636,N_3151);
nand U5348 (N_5348,N_3309,N_3421);
nand U5349 (N_5349,N_3425,N_2974);
nand U5350 (N_5350,N_2453,N_3244);
nand U5351 (N_5351,N_3275,N_3766);
and U5352 (N_5352,N_2707,N_2405);
or U5353 (N_5353,N_3793,N_2647);
or U5354 (N_5354,N_2413,N_2053);
xnor U5355 (N_5355,N_2422,N_2176);
or U5356 (N_5356,N_3146,N_3678);
nor U5357 (N_5357,N_2730,N_3885);
and U5358 (N_5358,N_3194,N_2979);
nand U5359 (N_5359,N_2681,N_3800);
nor U5360 (N_5360,N_2492,N_2940);
nor U5361 (N_5361,N_3118,N_2472);
or U5362 (N_5362,N_2433,N_3611);
or U5363 (N_5363,N_2781,N_3192);
nor U5364 (N_5364,N_3768,N_3066);
and U5365 (N_5365,N_2915,N_2861);
xor U5366 (N_5366,N_3634,N_2643);
or U5367 (N_5367,N_2436,N_2128);
nand U5368 (N_5368,N_2774,N_3106);
and U5369 (N_5369,N_2665,N_2050);
or U5370 (N_5370,N_2113,N_2757);
and U5371 (N_5371,N_3155,N_3919);
and U5372 (N_5372,N_2941,N_2763);
or U5373 (N_5373,N_2055,N_2422);
and U5374 (N_5374,N_2237,N_3112);
or U5375 (N_5375,N_2277,N_3158);
nand U5376 (N_5376,N_3497,N_2123);
nand U5377 (N_5377,N_3410,N_3026);
xnor U5378 (N_5378,N_3316,N_2384);
nor U5379 (N_5379,N_3656,N_2934);
nor U5380 (N_5380,N_3502,N_3845);
and U5381 (N_5381,N_3007,N_2584);
or U5382 (N_5382,N_2285,N_3041);
and U5383 (N_5383,N_2624,N_3177);
nor U5384 (N_5384,N_2518,N_2354);
nand U5385 (N_5385,N_2688,N_2398);
or U5386 (N_5386,N_2768,N_2192);
or U5387 (N_5387,N_2494,N_3103);
xor U5388 (N_5388,N_2102,N_3945);
nand U5389 (N_5389,N_2405,N_2161);
nor U5390 (N_5390,N_2439,N_2427);
and U5391 (N_5391,N_2110,N_2902);
nand U5392 (N_5392,N_2046,N_2077);
or U5393 (N_5393,N_2687,N_2869);
and U5394 (N_5394,N_3624,N_2629);
or U5395 (N_5395,N_3306,N_2263);
and U5396 (N_5396,N_2368,N_2315);
nand U5397 (N_5397,N_2076,N_3300);
xor U5398 (N_5398,N_3540,N_3853);
xnor U5399 (N_5399,N_2046,N_2132);
or U5400 (N_5400,N_2841,N_3009);
and U5401 (N_5401,N_2501,N_3227);
nand U5402 (N_5402,N_3809,N_3770);
nor U5403 (N_5403,N_2002,N_3846);
nor U5404 (N_5404,N_2692,N_2341);
or U5405 (N_5405,N_2384,N_2860);
nand U5406 (N_5406,N_2209,N_2146);
and U5407 (N_5407,N_3220,N_3168);
nand U5408 (N_5408,N_2352,N_2166);
and U5409 (N_5409,N_2030,N_3546);
and U5410 (N_5410,N_2806,N_3645);
and U5411 (N_5411,N_2077,N_3937);
xnor U5412 (N_5412,N_2872,N_2122);
or U5413 (N_5413,N_3026,N_3615);
and U5414 (N_5414,N_3204,N_2523);
xnor U5415 (N_5415,N_3673,N_3445);
or U5416 (N_5416,N_2628,N_3558);
or U5417 (N_5417,N_2587,N_2079);
and U5418 (N_5418,N_3670,N_3860);
nor U5419 (N_5419,N_2458,N_2029);
or U5420 (N_5420,N_3819,N_2333);
or U5421 (N_5421,N_3630,N_2424);
and U5422 (N_5422,N_3289,N_3828);
or U5423 (N_5423,N_2877,N_3739);
or U5424 (N_5424,N_2992,N_3964);
nand U5425 (N_5425,N_2365,N_3851);
or U5426 (N_5426,N_3611,N_3494);
nand U5427 (N_5427,N_2041,N_2953);
nand U5428 (N_5428,N_3988,N_2671);
or U5429 (N_5429,N_3290,N_3114);
and U5430 (N_5430,N_3203,N_2799);
nand U5431 (N_5431,N_3658,N_3147);
and U5432 (N_5432,N_3903,N_3473);
or U5433 (N_5433,N_2869,N_3813);
and U5434 (N_5434,N_2203,N_2161);
nor U5435 (N_5435,N_3169,N_3810);
nor U5436 (N_5436,N_2963,N_3627);
or U5437 (N_5437,N_2969,N_3965);
nor U5438 (N_5438,N_3526,N_3662);
nand U5439 (N_5439,N_2238,N_2487);
nor U5440 (N_5440,N_2947,N_2044);
nand U5441 (N_5441,N_2360,N_2542);
or U5442 (N_5442,N_2038,N_2033);
or U5443 (N_5443,N_3808,N_2071);
and U5444 (N_5444,N_3258,N_3118);
and U5445 (N_5445,N_2819,N_3114);
xor U5446 (N_5446,N_2712,N_3483);
nor U5447 (N_5447,N_3635,N_2404);
and U5448 (N_5448,N_3750,N_3835);
nor U5449 (N_5449,N_2955,N_2641);
nand U5450 (N_5450,N_3960,N_2452);
nor U5451 (N_5451,N_3809,N_3896);
or U5452 (N_5452,N_2544,N_3864);
nor U5453 (N_5453,N_2839,N_2066);
and U5454 (N_5454,N_2214,N_3646);
and U5455 (N_5455,N_3035,N_2289);
or U5456 (N_5456,N_2775,N_2516);
nand U5457 (N_5457,N_2985,N_3183);
nand U5458 (N_5458,N_3070,N_2185);
nor U5459 (N_5459,N_2005,N_3666);
nor U5460 (N_5460,N_3359,N_3199);
and U5461 (N_5461,N_3434,N_2142);
and U5462 (N_5462,N_3801,N_3364);
and U5463 (N_5463,N_3789,N_2064);
and U5464 (N_5464,N_3425,N_2440);
or U5465 (N_5465,N_2978,N_3276);
nor U5466 (N_5466,N_3919,N_2874);
and U5467 (N_5467,N_2784,N_2243);
nor U5468 (N_5468,N_2488,N_2949);
and U5469 (N_5469,N_2336,N_3344);
nand U5470 (N_5470,N_2597,N_3026);
nor U5471 (N_5471,N_3350,N_3667);
and U5472 (N_5472,N_2211,N_2294);
xnor U5473 (N_5473,N_2199,N_2560);
nor U5474 (N_5474,N_3883,N_2704);
nor U5475 (N_5475,N_3909,N_2712);
and U5476 (N_5476,N_2745,N_3129);
nand U5477 (N_5477,N_3365,N_3874);
nand U5478 (N_5478,N_3660,N_3480);
nand U5479 (N_5479,N_2432,N_2567);
nor U5480 (N_5480,N_2999,N_3682);
and U5481 (N_5481,N_2994,N_2267);
nor U5482 (N_5482,N_3474,N_2531);
xor U5483 (N_5483,N_3614,N_2133);
nand U5484 (N_5484,N_2875,N_2299);
or U5485 (N_5485,N_2239,N_3490);
nor U5486 (N_5486,N_2991,N_3427);
nor U5487 (N_5487,N_3147,N_2600);
or U5488 (N_5488,N_2045,N_2572);
and U5489 (N_5489,N_3635,N_2001);
nor U5490 (N_5490,N_2896,N_3809);
nor U5491 (N_5491,N_2574,N_3030);
and U5492 (N_5492,N_3646,N_3464);
and U5493 (N_5493,N_2416,N_3520);
nand U5494 (N_5494,N_3480,N_3318);
nand U5495 (N_5495,N_3588,N_3749);
and U5496 (N_5496,N_3038,N_3068);
nand U5497 (N_5497,N_3035,N_3729);
xor U5498 (N_5498,N_2012,N_3864);
and U5499 (N_5499,N_3293,N_3124);
nor U5500 (N_5500,N_2349,N_2020);
xnor U5501 (N_5501,N_2802,N_2428);
and U5502 (N_5502,N_3790,N_3611);
nor U5503 (N_5503,N_3329,N_3466);
or U5504 (N_5504,N_3715,N_3280);
and U5505 (N_5505,N_2603,N_3701);
or U5506 (N_5506,N_2257,N_3327);
nand U5507 (N_5507,N_3582,N_2053);
or U5508 (N_5508,N_2795,N_3017);
nand U5509 (N_5509,N_3675,N_2757);
nand U5510 (N_5510,N_3214,N_3241);
nor U5511 (N_5511,N_2328,N_2650);
nand U5512 (N_5512,N_2915,N_3984);
and U5513 (N_5513,N_3300,N_2014);
xnor U5514 (N_5514,N_3135,N_2481);
or U5515 (N_5515,N_2181,N_3178);
nand U5516 (N_5516,N_3605,N_2222);
or U5517 (N_5517,N_3567,N_3511);
or U5518 (N_5518,N_2488,N_2135);
nand U5519 (N_5519,N_3929,N_2068);
nor U5520 (N_5520,N_2051,N_3653);
nand U5521 (N_5521,N_3807,N_3092);
nand U5522 (N_5522,N_3578,N_2201);
or U5523 (N_5523,N_2106,N_3147);
nor U5524 (N_5524,N_2533,N_3168);
and U5525 (N_5525,N_3318,N_3432);
and U5526 (N_5526,N_3850,N_3018);
nand U5527 (N_5527,N_2759,N_3803);
nand U5528 (N_5528,N_2637,N_2311);
xnor U5529 (N_5529,N_3964,N_3412);
and U5530 (N_5530,N_3607,N_3024);
nand U5531 (N_5531,N_3407,N_2292);
or U5532 (N_5532,N_2757,N_3089);
xor U5533 (N_5533,N_2127,N_3989);
nand U5534 (N_5534,N_3193,N_2578);
and U5535 (N_5535,N_3770,N_3760);
or U5536 (N_5536,N_3009,N_2606);
xor U5537 (N_5537,N_3295,N_3685);
nand U5538 (N_5538,N_2185,N_2681);
nand U5539 (N_5539,N_3149,N_2240);
nor U5540 (N_5540,N_2544,N_3689);
or U5541 (N_5541,N_3621,N_2573);
xor U5542 (N_5542,N_2778,N_3913);
nor U5543 (N_5543,N_3666,N_2762);
nand U5544 (N_5544,N_3546,N_2062);
xor U5545 (N_5545,N_3230,N_3617);
nor U5546 (N_5546,N_3043,N_3857);
or U5547 (N_5547,N_2707,N_2469);
or U5548 (N_5548,N_2828,N_3042);
and U5549 (N_5549,N_3841,N_3062);
or U5550 (N_5550,N_2007,N_2066);
nand U5551 (N_5551,N_3353,N_3492);
nand U5552 (N_5552,N_2348,N_2706);
nor U5553 (N_5553,N_3729,N_2484);
nand U5554 (N_5554,N_3639,N_3755);
or U5555 (N_5555,N_3715,N_3205);
or U5556 (N_5556,N_2875,N_2098);
xor U5557 (N_5557,N_2747,N_3749);
and U5558 (N_5558,N_2158,N_3191);
nor U5559 (N_5559,N_3096,N_3453);
or U5560 (N_5560,N_2846,N_2298);
and U5561 (N_5561,N_3330,N_2922);
or U5562 (N_5562,N_3811,N_2709);
and U5563 (N_5563,N_3347,N_2315);
nand U5564 (N_5564,N_3524,N_3168);
xnor U5565 (N_5565,N_2650,N_3083);
or U5566 (N_5566,N_2235,N_2638);
nand U5567 (N_5567,N_2470,N_2925);
or U5568 (N_5568,N_2295,N_2651);
xor U5569 (N_5569,N_2988,N_3089);
and U5570 (N_5570,N_2433,N_3823);
and U5571 (N_5571,N_2589,N_3547);
or U5572 (N_5572,N_3927,N_2562);
nor U5573 (N_5573,N_3051,N_2732);
nor U5574 (N_5574,N_3557,N_2147);
or U5575 (N_5575,N_3941,N_2084);
and U5576 (N_5576,N_3624,N_3575);
nand U5577 (N_5577,N_3387,N_2240);
or U5578 (N_5578,N_3953,N_2904);
or U5579 (N_5579,N_2278,N_3064);
nand U5580 (N_5580,N_2232,N_3918);
xor U5581 (N_5581,N_3866,N_3588);
and U5582 (N_5582,N_2388,N_2107);
and U5583 (N_5583,N_3472,N_3848);
nor U5584 (N_5584,N_3734,N_3165);
nand U5585 (N_5585,N_3194,N_3567);
and U5586 (N_5586,N_3791,N_2689);
nor U5587 (N_5587,N_3268,N_3407);
nor U5588 (N_5588,N_3512,N_2633);
and U5589 (N_5589,N_3994,N_2759);
nor U5590 (N_5590,N_2921,N_3151);
and U5591 (N_5591,N_2171,N_2327);
nand U5592 (N_5592,N_3229,N_3695);
and U5593 (N_5593,N_3392,N_2559);
and U5594 (N_5594,N_2384,N_2864);
nor U5595 (N_5595,N_2904,N_2574);
or U5596 (N_5596,N_2281,N_2463);
nor U5597 (N_5597,N_2772,N_3062);
nand U5598 (N_5598,N_3203,N_3292);
nand U5599 (N_5599,N_3968,N_2434);
nor U5600 (N_5600,N_3298,N_3623);
xor U5601 (N_5601,N_3344,N_2390);
nor U5602 (N_5602,N_2715,N_2512);
nor U5603 (N_5603,N_3741,N_3558);
nor U5604 (N_5604,N_3671,N_3691);
or U5605 (N_5605,N_2414,N_2765);
nor U5606 (N_5606,N_2754,N_3524);
and U5607 (N_5607,N_2291,N_2593);
and U5608 (N_5608,N_2562,N_3606);
nor U5609 (N_5609,N_3976,N_2581);
xor U5610 (N_5610,N_3907,N_3769);
nor U5611 (N_5611,N_2843,N_3006);
nand U5612 (N_5612,N_3263,N_3000);
nor U5613 (N_5613,N_2292,N_2522);
or U5614 (N_5614,N_3676,N_3463);
or U5615 (N_5615,N_3705,N_2634);
nor U5616 (N_5616,N_2563,N_3846);
or U5617 (N_5617,N_3707,N_3435);
xnor U5618 (N_5618,N_2256,N_3992);
or U5619 (N_5619,N_3965,N_3398);
nand U5620 (N_5620,N_3864,N_3214);
or U5621 (N_5621,N_2672,N_3815);
xor U5622 (N_5622,N_2658,N_2352);
nor U5623 (N_5623,N_3855,N_2749);
nor U5624 (N_5624,N_3384,N_3951);
nor U5625 (N_5625,N_2810,N_3582);
nand U5626 (N_5626,N_2613,N_2998);
nor U5627 (N_5627,N_2348,N_3393);
or U5628 (N_5628,N_3459,N_3488);
and U5629 (N_5629,N_3908,N_3224);
nand U5630 (N_5630,N_3231,N_3007);
nand U5631 (N_5631,N_3388,N_3099);
nand U5632 (N_5632,N_2603,N_2595);
or U5633 (N_5633,N_3812,N_3865);
xnor U5634 (N_5634,N_3793,N_3917);
and U5635 (N_5635,N_2961,N_2874);
or U5636 (N_5636,N_3650,N_2181);
nand U5637 (N_5637,N_2534,N_2878);
xnor U5638 (N_5638,N_2002,N_2169);
nor U5639 (N_5639,N_2122,N_2358);
or U5640 (N_5640,N_2554,N_3651);
and U5641 (N_5641,N_3491,N_2684);
nor U5642 (N_5642,N_2824,N_2666);
or U5643 (N_5643,N_3969,N_3677);
nor U5644 (N_5644,N_2428,N_3323);
nand U5645 (N_5645,N_3674,N_2025);
nor U5646 (N_5646,N_2104,N_2583);
xor U5647 (N_5647,N_2789,N_2555);
nand U5648 (N_5648,N_2980,N_3975);
and U5649 (N_5649,N_3405,N_2245);
xor U5650 (N_5650,N_3067,N_2793);
nand U5651 (N_5651,N_3520,N_3592);
and U5652 (N_5652,N_3554,N_2169);
and U5653 (N_5653,N_3032,N_2589);
or U5654 (N_5654,N_2067,N_3283);
xor U5655 (N_5655,N_2010,N_3197);
or U5656 (N_5656,N_3251,N_2419);
nand U5657 (N_5657,N_3817,N_3055);
nand U5658 (N_5658,N_2986,N_3661);
nand U5659 (N_5659,N_3365,N_3371);
nor U5660 (N_5660,N_2470,N_2215);
xor U5661 (N_5661,N_3827,N_3916);
nand U5662 (N_5662,N_3303,N_2321);
xor U5663 (N_5663,N_3982,N_3563);
or U5664 (N_5664,N_2628,N_3883);
and U5665 (N_5665,N_2418,N_3890);
and U5666 (N_5666,N_3131,N_2205);
and U5667 (N_5667,N_3571,N_3900);
or U5668 (N_5668,N_2085,N_2474);
or U5669 (N_5669,N_2311,N_3513);
xor U5670 (N_5670,N_2078,N_3052);
and U5671 (N_5671,N_2012,N_2410);
xor U5672 (N_5672,N_3093,N_3527);
or U5673 (N_5673,N_3010,N_2175);
nor U5674 (N_5674,N_3447,N_3378);
and U5675 (N_5675,N_2938,N_3981);
and U5676 (N_5676,N_3890,N_2837);
and U5677 (N_5677,N_3724,N_2770);
xor U5678 (N_5678,N_2814,N_3225);
nand U5679 (N_5679,N_2409,N_3818);
or U5680 (N_5680,N_2809,N_2494);
or U5681 (N_5681,N_3566,N_2818);
xor U5682 (N_5682,N_2444,N_2173);
and U5683 (N_5683,N_3405,N_2136);
or U5684 (N_5684,N_3151,N_3344);
and U5685 (N_5685,N_3605,N_2838);
and U5686 (N_5686,N_2935,N_2697);
nand U5687 (N_5687,N_2578,N_3258);
and U5688 (N_5688,N_3501,N_2005);
or U5689 (N_5689,N_3583,N_3698);
nor U5690 (N_5690,N_3752,N_3430);
or U5691 (N_5691,N_2552,N_2076);
nand U5692 (N_5692,N_3229,N_3984);
nand U5693 (N_5693,N_2530,N_3845);
xnor U5694 (N_5694,N_2272,N_2896);
nor U5695 (N_5695,N_2526,N_3082);
and U5696 (N_5696,N_2625,N_2766);
nor U5697 (N_5697,N_3215,N_2693);
nor U5698 (N_5698,N_3534,N_3890);
and U5699 (N_5699,N_3734,N_3465);
nand U5700 (N_5700,N_3614,N_2240);
and U5701 (N_5701,N_3264,N_3782);
and U5702 (N_5702,N_3143,N_2457);
nor U5703 (N_5703,N_2572,N_3628);
nand U5704 (N_5704,N_3729,N_2608);
or U5705 (N_5705,N_2443,N_3515);
nor U5706 (N_5706,N_3880,N_3652);
nand U5707 (N_5707,N_2721,N_3400);
nand U5708 (N_5708,N_2102,N_2540);
xor U5709 (N_5709,N_3290,N_2021);
and U5710 (N_5710,N_2801,N_2819);
nand U5711 (N_5711,N_2637,N_2008);
nand U5712 (N_5712,N_2226,N_3054);
nor U5713 (N_5713,N_2483,N_3479);
or U5714 (N_5714,N_3845,N_2232);
and U5715 (N_5715,N_2484,N_2368);
or U5716 (N_5716,N_3173,N_2889);
or U5717 (N_5717,N_3302,N_3598);
xnor U5718 (N_5718,N_3141,N_3341);
or U5719 (N_5719,N_3437,N_2419);
nand U5720 (N_5720,N_3898,N_3909);
and U5721 (N_5721,N_3504,N_2193);
nor U5722 (N_5722,N_2033,N_2412);
nand U5723 (N_5723,N_3784,N_3942);
or U5724 (N_5724,N_2294,N_2302);
nor U5725 (N_5725,N_2798,N_3450);
and U5726 (N_5726,N_3228,N_2491);
and U5727 (N_5727,N_3261,N_2732);
or U5728 (N_5728,N_3533,N_2845);
nand U5729 (N_5729,N_3367,N_2531);
nor U5730 (N_5730,N_3131,N_2162);
nand U5731 (N_5731,N_2106,N_3429);
nor U5732 (N_5732,N_2352,N_2409);
xnor U5733 (N_5733,N_2241,N_2572);
or U5734 (N_5734,N_3165,N_3423);
nand U5735 (N_5735,N_2088,N_3010);
and U5736 (N_5736,N_2845,N_2780);
nor U5737 (N_5737,N_3915,N_3081);
xor U5738 (N_5738,N_3369,N_2698);
xnor U5739 (N_5739,N_2883,N_2334);
nor U5740 (N_5740,N_3748,N_2784);
and U5741 (N_5741,N_3474,N_2329);
or U5742 (N_5742,N_2483,N_2503);
nand U5743 (N_5743,N_3214,N_2558);
xor U5744 (N_5744,N_2213,N_3880);
nand U5745 (N_5745,N_2058,N_3056);
or U5746 (N_5746,N_3311,N_3119);
and U5747 (N_5747,N_2793,N_3082);
xor U5748 (N_5748,N_3972,N_2805);
xor U5749 (N_5749,N_2152,N_3637);
nor U5750 (N_5750,N_3948,N_2080);
and U5751 (N_5751,N_3774,N_3249);
nor U5752 (N_5752,N_2375,N_2452);
and U5753 (N_5753,N_2247,N_2105);
nor U5754 (N_5754,N_2483,N_2545);
and U5755 (N_5755,N_2291,N_2258);
nor U5756 (N_5756,N_3485,N_3075);
and U5757 (N_5757,N_2079,N_2624);
and U5758 (N_5758,N_3619,N_3242);
nand U5759 (N_5759,N_3500,N_2117);
and U5760 (N_5760,N_2629,N_3154);
and U5761 (N_5761,N_2726,N_3772);
or U5762 (N_5762,N_2486,N_2675);
or U5763 (N_5763,N_2351,N_2429);
or U5764 (N_5764,N_2765,N_2142);
and U5765 (N_5765,N_2218,N_2821);
nor U5766 (N_5766,N_3330,N_2037);
and U5767 (N_5767,N_3852,N_3430);
nand U5768 (N_5768,N_3671,N_2094);
nor U5769 (N_5769,N_2810,N_3747);
nand U5770 (N_5770,N_2666,N_3190);
nor U5771 (N_5771,N_2261,N_2247);
or U5772 (N_5772,N_3037,N_2949);
and U5773 (N_5773,N_3715,N_3984);
nor U5774 (N_5774,N_2327,N_3042);
nor U5775 (N_5775,N_3527,N_2149);
nand U5776 (N_5776,N_3344,N_2156);
nor U5777 (N_5777,N_3512,N_3657);
nor U5778 (N_5778,N_3923,N_3663);
or U5779 (N_5779,N_2700,N_3651);
xor U5780 (N_5780,N_2577,N_3257);
and U5781 (N_5781,N_3301,N_3059);
nand U5782 (N_5782,N_2826,N_2892);
xnor U5783 (N_5783,N_3129,N_2361);
and U5784 (N_5784,N_3767,N_2205);
nor U5785 (N_5785,N_3834,N_3163);
nand U5786 (N_5786,N_3111,N_3910);
nand U5787 (N_5787,N_3418,N_2638);
or U5788 (N_5788,N_2739,N_3964);
nor U5789 (N_5789,N_2715,N_3076);
nor U5790 (N_5790,N_2959,N_3517);
and U5791 (N_5791,N_2148,N_3098);
and U5792 (N_5792,N_2715,N_3858);
nor U5793 (N_5793,N_3125,N_3297);
and U5794 (N_5794,N_2401,N_2506);
or U5795 (N_5795,N_2937,N_3961);
or U5796 (N_5796,N_2876,N_3340);
and U5797 (N_5797,N_3227,N_2714);
and U5798 (N_5798,N_2843,N_3546);
xnor U5799 (N_5799,N_3975,N_2013);
nor U5800 (N_5800,N_2188,N_2177);
nor U5801 (N_5801,N_2144,N_3450);
nor U5802 (N_5802,N_2515,N_3835);
and U5803 (N_5803,N_2979,N_2635);
and U5804 (N_5804,N_3383,N_3834);
xnor U5805 (N_5805,N_2001,N_2650);
nand U5806 (N_5806,N_2008,N_2759);
nor U5807 (N_5807,N_2019,N_3126);
and U5808 (N_5808,N_3904,N_2225);
and U5809 (N_5809,N_2789,N_2733);
nand U5810 (N_5810,N_2453,N_3068);
nand U5811 (N_5811,N_3305,N_3445);
nand U5812 (N_5812,N_3847,N_3827);
xor U5813 (N_5813,N_2326,N_3244);
nor U5814 (N_5814,N_2198,N_2452);
nor U5815 (N_5815,N_2423,N_2241);
or U5816 (N_5816,N_2815,N_3951);
or U5817 (N_5817,N_2944,N_3449);
or U5818 (N_5818,N_3223,N_3385);
xor U5819 (N_5819,N_2359,N_2903);
and U5820 (N_5820,N_2834,N_2962);
xor U5821 (N_5821,N_2609,N_2586);
nand U5822 (N_5822,N_2013,N_3895);
nand U5823 (N_5823,N_3277,N_3086);
or U5824 (N_5824,N_3519,N_3498);
nor U5825 (N_5825,N_3450,N_2804);
or U5826 (N_5826,N_2240,N_2133);
nand U5827 (N_5827,N_2949,N_2280);
and U5828 (N_5828,N_3099,N_2608);
and U5829 (N_5829,N_3020,N_2975);
nand U5830 (N_5830,N_3683,N_3155);
nand U5831 (N_5831,N_3924,N_2403);
nand U5832 (N_5832,N_3043,N_2985);
nor U5833 (N_5833,N_3749,N_3171);
and U5834 (N_5834,N_2356,N_3253);
or U5835 (N_5835,N_2953,N_2395);
and U5836 (N_5836,N_3390,N_2565);
nand U5837 (N_5837,N_3768,N_3063);
or U5838 (N_5838,N_2767,N_2909);
xor U5839 (N_5839,N_3150,N_2975);
nand U5840 (N_5840,N_2727,N_3021);
and U5841 (N_5841,N_3785,N_3655);
or U5842 (N_5842,N_2489,N_2588);
or U5843 (N_5843,N_3906,N_2317);
nor U5844 (N_5844,N_2651,N_3680);
nand U5845 (N_5845,N_2136,N_2390);
nand U5846 (N_5846,N_3785,N_2949);
or U5847 (N_5847,N_2548,N_2777);
nand U5848 (N_5848,N_2379,N_3639);
or U5849 (N_5849,N_3587,N_3603);
and U5850 (N_5850,N_3390,N_2788);
nand U5851 (N_5851,N_2116,N_3531);
or U5852 (N_5852,N_2467,N_3312);
nand U5853 (N_5853,N_3505,N_2961);
or U5854 (N_5854,N_2755,N_3218);
or U5855 (N_5855,N_3956,N_2983);
nor U5856 (N_5856,N_2421,N_3808);
and U5857 (N_5857,N_3173,N_3824);
nor U5858 (N_5858,N_2486,N_2748);
and U5859 (N_5859,N_3723,N_2795);
nor U5860 (N_5860,N_2669,N_2443);
nand U5861 (N_5861,N_2835,N_3254);
nor U5862 (N_5862,N_2733,N_2724);
or U5863 (N_5863,N_3093,N_3540);
nand U5864 (N_5864,N_3238,N_3645);
nor U5865 (N_5865,N_3246,N_2917);
or U5866 (N_5866,N_3419,N_3233);
nor U5867 (N_5867,N_2065,N_2411);
and U5868 (N_5868,N_3706,N_3710);
nor U5869 (N_5869,N_3439,N_3627);
nor U5870 (N_5870,N_2786,N_2336);
xnor U5871 (N_5871,N_2874,N_2854);
and U5872 (N_5872,N_2609,N_3826);
or U5873 (N_5873,N_3447,N_2885);
and U5874 (N_5874,N_3904,N_2064);
nand U5875 (N_5875,N_2769,N_2847);
xnor U5876 (N_5876,N_2151,N_3198);
nand U5877 (N_5877,N_3039,N_2582);
or U5878 (N_5878,N_2946,N_2290);
and U5879 (N_5879,N_2925,N_3149);
and U5880 (N_5880,N_2028,N_2932);
nor U5881 (N_5881,N_2218,N_2516);
and U5882 (N_5882,N_2642,N_2605);
and U5883 (N_5883,N_2017,N_3848);
nor U5884 (N_5884,N_2724,N_2204);
and U5885 (N_5885,N_2572,N_3225);
nor U5886 (N_5886,N_2184,N_3717);
nor U5887 (N_5887,N_3114,N_2353);
nor U5888 (N_5888,N_2614,N_2075);
xor U5889 (N_5889,N_2583,N_2714);
nor U5890 (N_5890,N_2211,N_2662);
or U5891 (N_5891,N_3178,N_2377);
nor U5892 (N_5892,N_3709,N_3285);
nand U5893 (N_5893,N_3524,N_2672);
nor U5894 (N_5894,N_2354,N_2850);
and U5895 (N_5895,N_3217,N_2372);
nor U5896 (N_5896,N_2991,N_3204);
and U5897 (N_5897,N_3188,N_3991);
nor U5898 (N_5898,N_3209,N_2100);
and U5899 (N_5899,N_2074,N_3519);
or U5900 (N_5900,N_3885,N_2141);
or U5901 (N_5901,N_3941,N_2644);
nor U5902 (N_5902,N_2567,N_2440);
nand U5903 (N_5903,N_2472,N_2859);
nor U5904 (N_5904,N_3586,N_3962);
and U5905 (N_5905,N_3979,N_2534);
or U5906 (N_5906,N_2372,N_3912);
nand U5907 (N_5907,N_2307,N_3517);
and U5908 (N_5908,N_3288,N_3278);
and U5909 (N_5909,N_2926,N_2137);
and U5910 (N_5910,N_2702,N_2803);
nand U5911 (N_5911,N_2762,N_3732);
nor U5912 (N_5912,N_2790,N_2051);
nand U5913 (N_5913,N_2333,N_2297);
and U5914 (N_5914,N_3346,N_3044);
or U5915 (N_5915,N_2746,N_3247);
and U5916 (N_5916,N_3016,N_3798);
nor U5917 (N_5917,N_3719,N_3187);
nor U5918 (N_5918,N_2645,N_2703);
xnor U5919 (N_5919,N_3306,N_2404);
xor U5920 (N_5920,N_3756,N_2287);
and U5921 (N_5921,N_2074,N_2717);
nand U5922 (N_5922,N_3333,N_2498);
and U5923 (N_5923,N_2731,N_2837);
nand U5924 (N_5924,N_3721,N_3855);
and U5925 (N_5925,N_3880,N_3199);
xor U5926 (N_5926,N_2399,N_3287);
and U5927 (N_5927,N_2698,N_2335);
and U5928 (N_5928,N_2230,N_2585);
and U5929 (N_5929,N_3106,N_3956);
nand U5930 (N_5930,N_2202,N_2427);
nor U5931 (N_5931,N_2563,N_3424);
nor U5932 (N_5932,N_3961,N_2864);
xor U5933 (N_5933,N_2163,N_2097);
xor U5934 (N_5934,N_2787,N_2920);
or U5935 (N_5935,N_3702,N_3139);
nor U5936 (N_5936,N_3648,N_3288);
and U5937 (N_5937,N_2517,N_2117);
and U5938 (N_5938,N_2538,N_2370);
nor U5939 (N_5939,N_2159,N_3795);
or U5940 (N_5940,N_2260,N_3595);
and U5941 (N_5941,N_3145,N_2990);
and U5942 (N_5942,N_2958,N_3631);
nand U5943 (N_5943,N_3751,N_3750);
or U5944 (N_5944,N_3927,N_2592);
nand U5945 (N_5945,N_2060,N_3079);
nor U5946 (N_5946,N_2045,N_3177);
and U5947 (N_5947,N_2532,N_3571);
and U5948 (N_5948,N_3386,N_2315);
nor U5949 (N_5949,N_2099,N_2649);
xnor U5950 (N_5950,N_3843,N_3025);
nand U5951 (N_5951,N_2643,N_3852);
or U5952 (N_5952,N_3321,N_3435);
and U5953 (N_5953,N_2663,N_2327);
xnor U5954 (N_5954,N_2250,N_2622);
nand U5955 (N_5955,N_2312,N_3449);
or U5956 (N_5956,N_2225,N_2713);
or U5957 (N_5957,N_2119,N_2748);
or U5958 (N_5958,N_2546,N_2944);
xnor U5959 (N_5959,N_2295,N_3991);
nor U5960 (N_5960,N_3563,N_3150);
or U5961 (N_5961,N_3859,N_3932);
or U5962 (N_5962,N_2914,N_3755);
nand U5963 (N_5963,N_2114,N_3081);
nor U5964 (N_5964,N_3914,N_3410);
nor U5965 (N_5965,N_2757,N_2187);
and U5966 (N_5966,N_3509,N_2744);
xor U5967 (N_5967,N_2128,N_2944);
nand U5968 (N_5968,N_3174,N_3916);
nor U5969 (N_5969,N_2682,N_3704);
nand U5970 (N_5970,N_3513,N_3371);
nor U5971 (N_5971,N_3194,N_3458);
xor U5972 (N_5972,N_2770,N_3037);
or U5973 (N_5973,N_3878,N_3234);
or U5974 (N_5974,N_2627,N_3842);
nor U5975 (N_5975,N_3234,N_2975);
xnor U5976 (N_5976,N_3286,N_3871);
nor U5977 (N_5977,N_3295,N_3345);
or U5978 (N_5978,N_2646,N_2354);
xor U5979 (N_5979,N_3250,N_3821);
and U5980 (N_5980,N_3251,N_3367);
and U5981 (N_5981,N_3701,N_3273);
or U5982 (N_5982,N_2715,N_3318);
nor U5983 (N_5983,N_3194,N_3233);
nand U5984 (N_5984,N_2878,N_3458);
nor U5985 (N_5985,N_2752,N_2635);
nor U5986 (N_5986,N_3036,N_3191);
and U5987 (N_5987,N_2393,N_3765);
and U5988 (N_5988,N_2442,N_3931);
or U5989 (N_5989,N_2274,N_2672);
nor U5990 (N_5990,N_3357,N_2385);
and U5991 (N_5991,N_3146,N_3855);
or U5992 (N_5992,N_3783,N_2215);
nand U5993 (N_5993,N_2626,N_3807);
and U5994 (N_5994,N_3044,N_2887);
nor U5995 (N_5995,N_3157,N_3649);
nand U5996 (N_5996,N_2850,N_2417);
nand U5997 (N_5997,N_2106,N_3048);
nor U5998 (N_5998,N_2737,N_2262);
nor U5999 (N_5999,N_2206,N_3594);
nand U6000 (N_6000,N_4218,N_4819);
or U6001 (N_6001,N_5555,N_5256);
nor U6002 (N_6002,N_5912,N_5350);
or U6003 (N_6003,N_5637,N_5651);
nor U6004 (N_6004,N_4581,N_5914);
nand U6005 (N_6005,N_5519,N_5053);
or U6006 (N_6006,N_5971,N_4281);
nand U6007 (N_6007,N_4249,N_5757);
xor U6008 (N_6008,N_4738,N_4724);
nor U6009 (N_6009,N_4144,N_4455);
xor U6010 (N_6010,N_5351,N_5685);
and U6011 (N_6011,N_5112,N_5015);
and U6012 (N_6012,N_5566,N_5771);
or U6013 (N_6013,N_5357,N_4019);
or U6014 (N_6014,N_5355,N_5412);
nand U6015 (N_6015,N_5106,N_5723);
and U6016 (N_6016,N_4418,N_4338);
nor U6017 (N_6017,N_5012,N_4464);
or U6018 (N_6018,N_5604,N_5968);
nor U6019 (N_6019,N_5255,N_4306);
nand U6020 (N_6020,N_5955,N_4305);
and U6021 (N_6021,N_4726,N_5481);
and U6022 (N_6022,N_5088,N_5742);
and U6023 (N_6023,N_4869,N_4862);
or U6024 (N_6024,N_4835,N_5185);
nand U6025 (N_6025,N_4322,N_4734);
nand U6026 (N_6026,N_5333,N_5583);
and U6027 (N_6027,N_4318,N_5608);
nor U6028 (N_6028,N_4477,N_4803);
or U6029 (N_6029,N_5774,N_5573);
nor U6030 (N_6030,N_5426,N_5375);
or U6031 (N_6031,N_5473,N_5267);
nor U6032 (N_6032,N_5219,N_5799);
nor U6033 (N_6033,N_5030,N_5992);
nand U6034 (N_6034,N_5850,N_5806);
nand U6035 (N_6035,N_4568,N_4556);
or U6036 (N_6036,N_4756,N_5014);
or U6037 (N_6037,N_5669,N_4754);
nor U6038 (N_6038,N_5849,N_4466);
and U6039 (N_6039,N_4026,N_4594);
nor U6040 (N_6040,N_4485,N_4409);
or U6041 (N_6041,N_5474,N_5092);
xnor U6042 (N_6042,N_5928,N_4105);
nor U6043 (N_6043,N_5520,N_5593);
nor U6044 (N_6044,N_4206,N_5384);
and U6045 (N_6045,N_5760,N_5073);
nor U6046 (N_6046,N_5802,N_4658);
and U6047 (N_6047,N_4312,N_5915);
or U6048 (N_6048,N_5117,N_4382);
nor U6049 (N_6049,N_5296,N_5538);
xnor U6050 (N_6050,N_5080,N_4775);
or U6051 (N_6051,N_5043,N_4171);
and U6052 (N_6052,N_5830,N_4336);
nand U6053 (N_6053,N_4173,N_4453);
nor U6054 (N_6054,N_5891,N_5901);
nor U6055 (N_6055,N_5998,N_4787);
xor U6056 (N_6056,N_5005,N_5602);
and U6057 (N_6057,N_5057,N_5562);
nor U6058 (N_6058,N_5242,N_4797);
or U6059 (N_6059,N_4555,N_4157);
nand U6060 (N_6060,N_4227,N_4744);
or U6061 (N_6061,N_4253,N_5087);
or U6062 (N_6062,N_4450,N_4930);
nor U6063 (N_6063,N_5281,N_4970);
nand U6064 (N_6064,N_5692,N_5571);
or U6065 (N_6065,N_4631,N_5151);
and U6066 (N_6066,N_5495,N_5488);
xnor U6067 (N_6067,N_4765,N_5009);
nand U6068 (N_6068,N_5887,N_5311);
or U6069 (N_6069,N_5740,N_4582);
or U6070 (N_6070,N_5622,N_5435);
nand U6071 (N_6071,N_4056,N_4152);
or U6072 (N_6072,N_4544,N_5297);
or U6073 (N_6073,N_5113,N_4510);
or U6074 (N_6074,N_4984,N_4686);
and U6075 (N_6075,N_5845,N_5455);
xnor U6076 (N_6076,N_5055,N_5721);
xnor U6077 (N_6077,N_4948,N_4628);
xnor U6078 (N_6078,N_4617,N_5741);
nor U6079 (N_6079,N_5963,N_5539);
or U6080 (N_6080,N_5874,N_4087);
xor U6081 (N_6081,N_5463,N_4843);
xnor U6082 (N_6082,N_5479,N_4012);
or U6083 (N_6083,N_5486,N_4528);
nand U6084 (N_6084,N_5527,N_4511);
xnor U6085 (N_6085,N_4127,N_5552);
nor U6086 (N_6086,N_4037,N_5205);
and U6087 (N_6087,N_4618,N_5789);
and U6088 (N_6088,N_5605,N_5938);
nor U6089 (N_6089,N_5660,N_4335);
or U6090 (N_6090,N_5973,N_4074);
nor U6091 (N_6091,N_4300,N_5490);
or U6092 (N_6092,N_5694,N_4462);
xnor U6093 (N_6093,N_4183,N_4569);
or U6094 (N_6094,N_4197,N_4494);
nor U6095 (N_6095,N_4636,N_5609);
and U6096 (N_6096,N_4264,N_5630);
nand U6097 (N_6097,N_4600,N_4616);
or U6098 (N_6098,N_5268,N_5688);
or U6099 (N_6099,N_4633,N_5542);
and U6100 (N_6100,N_5616,N_5260);
and U6101 (N_6101,N_4151,N_4910);
nor U6102 (N_6102,N_5549,N_5356);
nand U6103 (N_6103,N_5336,N_4236);
nor U6104 (N_6104,N_5244,N_5835);
and U6105 (N_6105,N_5632,N_4595);
or U6106 (N_6106,N_5946,N_5999);
and U6107 (N_6107,N_5429,N_4499);
and U6108 (N_6108,N_4325,N_4110);
or U6109 (N_6109,N_4311,N_4963);
or U6110 (N_6110,N_5229,N_5339);
or U6111 (N_6111,N_4131,N_5863);
nor U6112 (N_6112,N_5374,N_5886);
nor U6113 (N_6113,N_4760,N_5409);
nor U6114 (N_6114,N_4246,N_5642);
nor U6115 (N_6115,N_5082,N_5725);
or U6116 (N_6116,N_4924,N_5842);
xor U6117 (N_6117,N_5328,N_5294);
nand U6118 (N_6118,N_5361,N_4373);
nor U6119 (N_6119,N_5257,N_5035);
nand U6120 (N_6120,N_4199,N_5407);
nand U6121 (N_6121,N_4656,N_4178);
and U6122 (N_6122,N_5241,N_5147);
xor U6123 (N_6123,N_4530,N_5708);
and U6124 (N_6124,N_4132,N_5607);
nand U6125 (N_6125,N_5900,N_4799);
and U6126 (N_6126,N_4333,N_4412);
and U6127 (N_6127,N_5024,N_5044);
nand U6128 (N_6128,N_5293,N_4971);
xor U6129 (N_6129,N_5115,N_4863);
nor U6130 (N_6130,N_4372,N_5195);
nor U6131 (N_6131,N_5049,N_4168);
and U6132 (N_6132,N_5084,N_5516);
xnor U6133 (N_6133,N_5916,N_4039);
nor U6134 (N_6134,N_4065,N_4330);
nor U6135 (N_6135,N_4606,N_5906);
or U6136 (N_6136,N_4292,N_4534);
or U6137 (N_6137,N_4115,N_4164);
nand U6138 (N_6138,N_5981,N_5977);
nand U6139 (N_6139,N_5272,N_5840);
or U6140 (N_6140,N_5144,N_5397);
nand U6141 (N_6141,N_5653,N_5395);
or U6142 (N_6142,N_5211,N_5947);
and U6143 (N_6143,N_5780,N_4564);
or U6144 (N_6144,N_4147,N_4163);
nand U6145 (N_6145,N_4807,N_4001);
and U6146 (N_6146,N_4945,N_4410);
nor U6147 (N_6147,N_5162,N_4229);
and U6148 (N_6148,N_4624,N_4154);
nand U6149 (N_6149,N_4532,N_5331);
nor U6150 (N_6150,N_4800,N_5228);
or U6151 (N_6151,N_5169,N_4603);
or U6152 (N_6152,N_4469,N_5402);
nor U6153 (N_6153,N_4999,N_4733);
or U6154 (N_6154,N_4706,N_4166);
or U6155 (N_6155,N_5501,N_4943);
or U6156 (N_6156,N_5114,N_5003);
nand U6157 (N_6157,N_4665,N_4195);
nand U6158 (N_6158,N_5668,N_5783);
and U6159 (N_6159,N_5867,N_5366);
nor U6160 (N_6160,N_5323,N_4059);
and U6161 (N_6161,N_4830,N_5526);
and U6162 (N_6162,N_4088,N_5160);
nand U6163 (N_6163,N_4707,N_5852);
xnor U6164 (N_6164,N_5844,N_5235);
or U6165 (N_6165,N_4442,N_5624);
or U6166 (N_6166,N_4732,N_5360);
nor U6167 (N_6167,N_5793,N_4189);
nand U6168 (N_6168,N_4050,N_5039);
or U6169 (N_6169,N_4172,N_5620);
nand U6170 (N_6170,N_5826,N_5428);
nor U6171 (N_6171,N_5365,N_4885);
nand U6172 (N_6172,N_4884,N_4793);
and U6173 (N_6173,N_4233,N_4076);
nand U6174 (N_6174,N_4630,N_4145);
and U6175 (N_6175,N_5489,N_4317);
nor U6176 (N_6176,N_5439,N_5823);
nor U6177 (N_6177,N_4136,N_5274);
nand U6178 (N_6178,N_5535,N_5512);
nor U6179 (N_6179,N_4085,N_4035);
nand U6180 (N_6180,N_4276,N_4896);
nor U6181 (N_6181,N_5319,N_4991);
or U6182 (N_6182,N_4813,N_4004);
xnor U6183 (N_6183,N_5730,N_5070);
nor U6184 (N_6184,N_5478,N_4685);
nand U6185 (N_6185,N_4763,N_4722);
and U6186 (N_6186,N_4492,N_4096);
nor U6187 (N_6187,N_5989,N_5313);
xnor U6188 (N_6188,N_5058,N_5908);
nand U6189 (N_6189,N_4708,N_4586);
nand U6190 (N_6190,N_4768,N_4047);
nand U6191 (N_6191,N_4956,N_5001);
and U6192 (N_6192,N_4380,N_5770);
or U6193 (N_6193,N_4626,N_5717);
or U6194 (N_6194,N_5217,N_4950);
or U6195 (N_6195,N_5433,N_5584);
xor U6196 (N_6196,N_4424,N_5484);
or U6197 (N_6197,N_4516,N_5076);
xor U6198 (N_6198,N_5990,N_4878);
and U6199 (N_6199,N_5939,N_4831);
nand U6200 (N_6200,N_4736,N_5290);
nor U6201 (N_6201,N_5864,N_5346);
and U6202 (N_6202,N_5687,N_5019);
and U6203 (N_6203,N_4832,N_5879);
nor U6204 (N_6204,N_4653,N_5899);
xor U6205 (N_6205,N_5400,N_5672);
or U6206 (N_6206,N_4891,N_4470);
and U6207 (N_6207,N_5748,N_5872);
nor U6208 (N_6208,N_5881,N_4904);
xnor U6209 (N_6209,N_4903,N_5533);
and U6210 (N_6210,N_5031,N_5013);
nor U6211 (N_6211,N_5069,N_4279);
or U6212 (N_6212,N_4068,N_4961);
nand U6213 (N_6213,N_4941,N_4286);
nor U6214 (N_6214,N_5321,N_4451);
nand U6215 (N_6215,N_4170,N_5779);
nor U6216 (N_6216,N_4659,N_5595);
nor U6217 (N_6217,N_5784,N_5119);
nor U6218 (N_6218,N_5391,N_5421);
or U6219 (N_6219,N_4978,N_4947);
and U6220 (N_6220,N_4024,N_5875);
nor U6221 (N_6221,N_5979,N_4073);
or U6222 (N_6222,N_5695,N_5851);
nand U6223 (N_6223,N_5367,N_4875);
and U6224 (N_6224,N_5349,N_5659);
nand U6225 (N_6225,N_4901,N_4911);
nor U6226 (N_6226,N_4417,N_4124);
xor U6227 (N_6227,N_5173,N_5052);
or U6228 (N_6228,N_4866,N_5016);
nand U6229 (N_6229,N_4025,N_5657);
or U6230 (N_6230,N_4975,N_4497);
xor U6231 (N_6231,N_5270,N_4584);
and U6232 (N_6232,N_4027,N_4880);
nand U6233 (N_6233,N_5825,N_5812);
nor U6234 (N_6234,N_4690,N_4482);
or U6235 (N_6235,N_4161,N_5101);
and U6236 (N_6236,N_5329,N_5600);
nand U6237 (N_6237,N_5379,N_4585);
xor U6238 (N_6238,N_5658,N_5691);
nand U6239 (N_6239,N_4622,N_4245);
nand U6240 (N_6240,N_5085,N_4811);
nand U6241 (N_6241,N_5183,N_4357);
and U6242 (N_6242,N_5929,N_5314);
nand U6243 (N_6243,N_5332,N_5021);
and U6244 (N_6244,N_4796,N_4664);
nor U6245 (N_6245,N_4777,N_4887);
nor U6246 (N_6246,N_4208,N_5591);
nor U6247 (N_6247,N_4541,N_4965);
nand U6248 (N_6248,N_4040,N_5671);
nor U6249 (N_6249,N_5677,N_4542);
xor U6250 (N_6250,N_5203,N_5061);
and U6251 (N_6251,N_5615,N_4888);
or U6252 (N_6252,N_4996,N_4704);
nor U6253 (N_6253,N_5027,N_5824);
xor U6254 (N_6254,N_5673,N_4188);
and U6255 (N_6255,N_5233,N_5704);
and U6256 (N_6256,N_5415,N_4160);
xor U6257 (N_6257,N_5416,N_4070);
xnor U6258 (N_6258,N_5179,N_5662);
nor U6259 (N_6259,N_5305,N_4363);
nand U6260 (N_6260,N_5556,N_4551);
nand U6261 (N_6261,N_5862,N_5860);
nor U6262 (N_6262,N_4923,N_4433);
nor U6263 (N_6263,N_5337,N_5884);
and U6264 (N_6264,N_5143,N_4049);
or U6265 (N_6265,N_4812,N_4919);
xnor U6266 (N_6266,N_4436,N_4241);
nand U6267 (N_6267,N_4192,N_4444);
nor U6268 (N_6268,N_5258,N_4898);
and U6269 (N_6269,N_5347,N_5372);
xnor U6270 (N_6270,N_4590,N_4044);
and U6271 (N_6271,N_4849,N_4925);
and U6272 (N_6272,N_5964,N_4751);
and U6273 (N_6273,N_5420,N_5953);
nand U6274 (N_6274,N_5735,N_4748);
and U6275 (N_6275,N_4645,N_5759);
or U6276 (N_6276,N_5105,N_4545);
nor U6277 (N_6277,N_5686,N_4657);
nor U6278 (N_6278,N_4861,N_4016);
or U6279 (N_6279,N_4119,N_4678);
nor U6280 (N_6280,N_5978,N_5067);
nand U6281 (N_6281,N_5038,N_4562);
and U6282 (N_6282,N_4329,N_4725);
nor U6283 (N_6283,N_4829,N_5706);
nor U6284 (N_6284,N_5696,N_5292);
nor U6285 (N_6285,N_5100,N_5291);
nand U6286 (N_6286,N_4599,N_4271);
nand U6287 (N_6287,N_5588,N_4272);
and U6288 (N_6288,N_5453,N_4354);
nor U6289 (N_6289,N_4092,N_5763);
nand U6290 (N_6290,N_4993,N_5965);
nor U6291 (N_6291,N_5514,N_5800);
nand U6292 (N_6292,N_5109,N_5952);
and U6293 (N_6293,N_5747,N_4546);
or U6294 (N_6294,N_4502,N_5454);
nand U6295 (N_6295,N_4205,N_5619);
and U6296 (N_6296,N_4447,N_4902);
or U6297 (N_6297,N_5865,N_4150);
and U6298 (N_6298,N_4495,N_5425);
nor U6299 (N_6299,N_4334,N_5623);
nand U6300 (N_6300,N_4739,N_4285);
nor U6301 (N_6301,N_4086,N_5437);
nor U6302 (N_6302,N_5186,N_5189);
nand U6303 (N_6303,N_4968,N_5079);
or U6304 (N_6304,N_4596,N_4129);
or U6305 (N_6305,N_5873,N_5482);
or U6306 (N_6306,N_4366,N_5383);
nor U6307 (N_6307,N_5491,N_5712);
and U6308 (N_6308,N_4839,N_5164);
or U6309 (N_6309,N_5475,N_4431);
and U6310 (N_6310,N_5951,N_4295);
nand U6311 (N_6311,N_4121,N_5251);
nor U6312 (N_6312,N_4815,N_5132);
or U6313 (N_6313,N_5497,N_4034);
and U6314 (N_6314,N_5613,N_5983);
nor U6315 (N_6315,N_4006,N_5170);
and U6316 (N_6316,N_4109,N_4106);
or U6317 (N_6317,N_4231,N_4742);
nand U6318 (N_6318,N_4240,N_5452);
or U6319 (N_6319,N_4429,N_5046);
nor U6320 (N_6320,N_4204,N_5450);
nand U6321 (N_6321,N_5149,N_4773);
nand U6322 (N_6322,N_4142,N_4571);
nor U6323 (N_6323,N_5911,N_5335);
nor U6324 (N_6324,N_5025,N_4604);
and U6325 (N_6325,N_5166,N_5004);
xor U6326 (N_6326,N_5617,N_5643);
nand U6327 (N_6327,N_5640,N_5805);
xor U6328 (N_6328,N_4400,N_4989);
nor U6329 (N_6329,N_5062,N_5821);
or U6330 (N_6330,N_5580,N_4488);
nand U6331 (N_6331,N_5568,N_4349);
and U6332 (N_6332,N_4848,N_5744);
nor U6333 (N_6333,N_5102,N_5933);
and U6334 (N_6334,N_4360,N_5287);
or U6335 (N_6335,N_4407,N_5903);
or U6336 (N_6336,N_4883,N_4897);
nand U6337 (N_6337,N_5168,N_5813);
and U6338 (N_6338,N_4368,N_4927);
nand U6339 (N_6339,N_4261,N_5697);
or U6340 (N_6340,N_5729,N_5773);
or U6341 (N_6341,N_4364,N_5667);
or U6342 (N_6342,N_4038,N_5511);
nor U6343 (N_6343,N_5045,N_5832);
and U6344 (N_6344,N_5022,N_4610);
or U6345 (N_6345,N_4028,N_4505);
or U6346 (N_6346,N_5065,N_5072);
nor U6347 (N_6347,N_4699,N_5104);
nor U6348 (N_6348,N_5414,N_4853);
nor U6349 (N_6349,N_4340,N_5111);
and U6350 (N_6350,N_4476,N_5829);
nor U6351 (N_6351,N_5836,N_4962);
and U6352 (N_6352,N_4094,N_5140);
and U6353 (N_6353,N_4913,N_5764);
nand U6354 (N_6354,N_4438,N_5177);
nand U6355 (N_6355,N_4457,N_4611);
or U6356 (N_6356,N_5116,N_5279);
and U6357 (N_6357,N_5618,N_5344);
nand U6358 (N_6358,N_5467,N_5389);
or U6359 (N_6359,N_5107,N_5230);
nand U6360 (N_6360,N_4655,N_5804);
and U6361 (N_6361,N_4053,N_4882);
and U6362 (N_6362,N_4967,N_5392);
and U6363 (N_6363,N_4522,N_4821);
and U6364 (N_6364,N_4045,N_4274);
nand U6365 (N_6365,N_4277,N_4194);
and U6366 (N_6366,N_4779,N_5206);
or U6367 (N_6367,N_4375,N_4117);
and U6368 (N_6368,N_4212,N_5093);
xnor U6369 (N_6369,N_4940,N_5182);
nand U6370 (N_6370,N_5252,N_5212);
nand U6371 (N_6371,N_5330,N_5582);
nand U6372 (N_6372,N_5610,N_5341);
nand U6373 (N_6373,N_5577,N_4269);
nor U6374 (N_6374,N_5496,N_5834);
nor U6375 (N_6375,N_5674,N_5408);
or U6376 (N_6376,N_4077,N_5724);
nand U6377 (N_6377,N_5843,N_4123);
nor U6378 (N_6378,N_5720,N_5818);
or U6379 (N_6379,N_4203,N_4536);
nor U6380 (N_6380,N_5769,N_4439);
nor U6381 (N_6381,N_4935,N_5504);
or U6382 (N_6382,N_5307,N_5814);
and U6383 (N_6383,N_4533,N_5447);
or U6384 (N_6384,N_4638,N_5858);
xor U6385 (N_6385,N_4523,N_4851);
xor U6386 (N_6386,N_4579,N_4367);
nor U6387 (N_6387,N_5997,N_5422);
and U6388 (N_6388,N_4679,N_4767);
or U6389 (N_6389,N_4647,N_4721);
nand U6390 (N_6390,N_5299,N_4557);
nand U6391 (N_6391,N_5472,N_4817);
xnor U6392 (N_6392,N_5442,N_4654);
nor U6393 (N_6393,N_4716,N_5026);
nor U6394 (N_6394,N_5056,N_4416);
nand U6395 (N_6395,N_5959,N_5534);
nand U6396 (N_6396,N_4827,N_5011);
or U6397 (N_6397,N_4232,N_5934);
or U6398 (N_6398,N_4358,N_4507);
nor U6399 (N_6399,N_5853,N_4578);
or U6400 (N_6400,N_5731,N_5098);
and U6401 (N_6401,N_4761,N_4820);
nor U6402 (N_6402,N_4979,N_5083);
nand U6403 (N_6403,N_5153,N_4634);
or U6404 (N_6404,N_4213,N_4396);
or U6405 (N_6405,N_4251,N_4191);
xnor U6406 (N_6406,N_4886,N_5423);
xor U6407 (N_6407,N_4508,N_4003);
and U6408 (N_6408,N_4823,N_4615);
nor U6409 (N_6409,N_4671,N_5920);
and U6410 (N_6410,N_4757,N_5469);
nand U6411 (N_6411,N_4196,N_4461);
or U6412 (N_6412,N_5459,N_5171);
nand U6413 (N_6413,N_4637,N_4452);
and U6414 (N_6414,N_4465,N_5418);
nand U6415 (N_6415,N_5123,N_5572);
xor U6416 (N_6416,N_5820,N_4662);
xnor U6417 (N_6417,N_5828,N_4425);
nor U6418 (N_6418,N_4632,N_5234);
or U6419 (N_6419,N_5761,N_4969);
xor U6420 (N_6420,N_5263,N_4042);
xnor U6421 (N_6421,N_4063,N_5524);
or U6422 (N_6422,N_4928,N_4228);
nand U6423 (N_6423,N_5071,N_4609);
and U6424 (N_6424,N_5611,N_4552);
and U6425 (N_6425,N_4937,N_4022);
or U6426 (N_6426,N_4252,N_5585);
or U6427 (N_6427,N_5917,N_4352);
and U6428 (N_6428,N_4877,N_4745);
nor U6429 (N_6429,N_5334,N_4083);
or U6430 (N_6430,N_4759,N_4694);
nand U6431 (N_6431,N_4283,N_4029);
nor U6432 (N_6432,N_5184,N_4730);
and U6433 (N_6433,N_5807,N_4876);
or U6434 (N_6434,N_5340,N_5406);
nand U6435 (N_6435,N_5885,N_5448);
nand U6436 (N_6436,N_5798,N_4268);
xnor U6437 (N_6437,N_5047,N_4934);
or U6438 (N_6438,N_5654,N_5621);
nand U6439 (N_6439,N_4486,N_5443);
and U6440 (N_6440,N_4974,N_5734);
nand U6441 (N_6441,N_4390,N_4114);
nand U6442 (N_6442,N_4275,N_4512);
and U6443 (N_6443,N_5969,N_5722);
nor U6444 (N_6444,N_4247,N_4135);
xor U6445 (N_6445,N_4198,N_4009);
and U6446 (N_6446,N_5126,N_4258);
or U6447 (N_6447,N_5924,N_4791);
nor U6448 (N_6448,N_5827,N_4054);
xnor U6449 (N_6449,N_5745,N_5318);
nand U6450 (N_6450,N_5477,N_4222);
nor U6451 (N_6451,N_4855,N_5795);
nand U6452 (N_6452,N_4293,N_5096);
or U6453 (N_6453,N_5181,N_4479);
nand U6454 (N_6454,N_4155,N_5141);
nor U6455 (N_6455,N_4846,N_5427);
xnor U6456 (N_6456,N_5300,N_5778);
and U6457 (N_6457,N_4200,N_5682);
nor U6458 (N_6458,N_5493,N_4408);
or U6459 (N_6459,N_5231,N_4981);
or U6460 (N_6460,N_5750,N_5954);
and U6461 (N_6461,N_4697,N_4201);
nor U6462 (N_6462,N_4126,N_4314);
nor U6463 (N_6463,N_5711,N_4262);
and U6464 (N_6464,N_5000,N_4066);
or U6465 (N_6465,N_5308,N_5546);
and U6466 (N_6466,N_5639,N_4872);
and U6467 (N_6467,N_4792,N_4860);
nand U6468 (N_6468,N_4392,N_4795);
nand U6469 (N_6469,N_5284,N_5188);
nor U6470 (N_6470,N_5918,N_4576);
nand U6471 (N_6471,N_4822,N_5574);
nand U6472 (N_6472,N_5364,N_4879);
or U6473 (N_6473,N_5156,N_5944);
and U6474 (N_6474,N_4990,N_4642);
nor U6475 (N_6475,N_5919,N_5628);
xor U6476 (N_6476,N_5398,N_5558);
nand U6477 (N_6477,N_5180,N_4503);
nand U6478 (N_6478,N_5500,N_4426);
nor U6479 (N_6479,N_5097,N_5666);
nor U6480 (N_6480,N_5878,N_4498);
nand U6481 (N_6481,N_4321,N_4376);
nor U6482 (N_6482,N_4560,N_5578);
or U6483 (N_6483,N_5883,N_4868);
nor U6484 (N_6484,N_5316,N_5378);
or U6485 (N_6485,N_4929,N_4052);
nor U6486 (N_6486,N_5950,N_5529);
nor U6487 (N_6487,N_5129,N_4319);
nor U6488 (N_6488,N_4701,N_4675);
and U6489 (N_6489,N_5381,N_5462);
or U6490 (N_6490,N_4220,N_4509);
nand U6491 (N_6491,N_4235,N_4058);
nor U6492 (N_6492,N_5271,N_5018);
or U6493 (N_6493,N_4017,N_5131);
nor U6494 (N_6494,N_5209,N_4668);
nor U6495 (N_6495,N_4415,N_5676);
nand U6496 (N_6496,N_4982,N_5831);
nor U6497 (N_6497,N_4303,N_5785);
xnor U6498 (N_6498,N_5214,N_4339);
nand U6499 (N_6499,N_4130,N_4386);
nor U6500 (N_6500,N_5103,N_5956);
or U6501 (N_6501,N_5975,N_4575);
nand U6502 (N_6502,N_5709,N_5841);
and U6503 (N_6503,N_5994,N_4113);
nand U6504 (N_6504,N_4384,N_5320);
or U6505 (N_6505,N_5120,N_4398);
or U6506 (N_6506,N_5210,N_5394);
nand U6507 (N_6507,N_5536,N_5559);
nor U6508 (N_6508,N_5194,N_4353);
or U6509 (N_6509,N_5197,N_4825);
xor U6510 (N_6510,N_5522,N_5303);
or U6511 (N_6511,N_4755,N_4640);
and U6512 (N_6512,N_4692,N_5089);
and U6513 (N_6513,N_4750,N_5603);
or U6514 (N_6514,N_5165,N_5515);
or U6515 (N_6515,N_5438,N_5819);
nand U6516 (N_6516,N_5966,N_4071);
or U6517 (N_6517,N_4798,N_5295);
and U6518 (N_6518,N_5354,N_4445);
xnor U6519 (N_6519,N_4490,N_5767);
and U6520 (N_6520,N_5358,N_4837);
or U6521 (N_6521,N_4120,N_4583);
and U6522 (N_6522,N_5159,N_5553);
or U6523 (N_6523,N_4080,N_4938);
and U6524 (N_6524,N_5138,N_4881);
or U6525 (N_6525,N_4824,N_4521);
or U6526 (N_6526,N_5848,N_5641);
xnor U6527 (N_6527,N_5684,N_5738);
and U6528 (N_6528,N_4097,N_4500);
and U6529 (N_6529,N_5680,N_4143);
nor U6530 (N_6530,N_5543,N_5464);
nand U6531 (N_6531,N_5846,N_5974);
and U6532 (N_6532,N_4953,N_5362);
nand U6533 (N_6533,N_5207,N_4854);
or U6534 (N_6534,N_4260,N_5099);
nor U6535 (N_6535,N_5077,N_4774);
xnor U6536 (N_6536,N_4471,N_4031);
nand U6537 (N_6537,N_4958,N_5560);
nor U6538 (N_6538,N_4737,N_4781);
nand U6539 (N_6539,N_5237,N_5589);
xnor U6540 (N_6540,N_4687,N_4986);
nor U6541 (N_6541,N_5431,N_5645);
or U6542 (N_6542,N_4243,N_5910);
or U6543 (N_6543,N_4816,N_4709);
nand U6544 (N_6544,N_5074,N_5273);
or U6545 (N_6545,N_5110,N_5838);
and U6546 (N_6546,N_4298,N_4018);
nor U6547 (N_6547,N_5794,N_4081);
nor U6548 (N_6548,N_5732,N_4696);
or U6549 (N_6549,N_4346,N_4587);
xor U6550 (N_6550,N_5561,N_4972);
nor U6551 (N_6551,N_5401,N_5809);
or U6552 (N_6552,N_4501,N_5776);
nand U6553 (N_6553,N_5193,N_5090);
or U6554 (N_6554,N_4591,N_5943);
and U6555 (N_6555,N_4980,N_4146);
nor U6556 (N_6556,N_4179,N_5661);
nor U6557 (N_6557,N_4137,N_5503);
and U6558 (N_6558,N_4176,N_5957);
or U6559 (N_6559,N_4356,N_5388);
xor U6560 (N_6560,N_4931,N_5980);
or U6561 (N_6561,N_4741,N_5487);
and U6562 (N_6562,N_5282,N_4676);
nand U6563 (N_6563,N_4535,N_4496);
or U6564 (N_6564,N_5949,N_4674);
or U6565 (N_6565,N_4381,N_5936);
nor U6566 (N_6566,N_4814,N_5440);
or U6567 (N_6567,N_4964,N_4614);
or U6568 (N_6568,N_5746,N_5494);
nor U6569 (N_6569,N_5815,N_4254);
nand U6570 (N_6570,N_4859,N_5801);
nand U6571 (N_6571,N_5386,N_5118);
and U6572 (N_6572,N_4187,N_4858);
nor U6573 (N_6573,N_5064,N_4936);
and U6574 (N_6574,N_5139,N_4175);
or U6575 (N_6575,N_5163,N_4794);
or U6576 (N_6576,N_5923,N_5877);
and U6577 (N_6577,N_5648,N_5289);
or U6578 (N_6578,N_5579,N_5020);
nand U6579 (N_6579,N_4307,N_4030);
xor U6580 (N_6580,N_5663,N_4051);
xnor U6581 (N_6581,N_4723,N_5703);
or U6582 (N_6582,N_5644,N_5839);
and U6583 (N_6583,N_4939,N_4342);
and U6584 (N_6584,N_4156,N_4580);
nand U6585 (N_6585,N_4519,N_4513);
nor U6586 (N_6586,N_4036,N_5714);
and U6587 (N_6587,N_4650,N_4348);
xnor U6588 (N_6588,N_4102,N_4652);
nand U6589 (N_6589,N_4209,N_4784);
and U6590 (N_6590,N_5960,N_5649);
and U6591 (N_6591,N_5010,N_4248);
nor U6592 (N_6592,N_4284,N_4731);
and U6593 (N_6593,N_5612,N_5446);
nor U6594 (N_6594,N_4921,N_4917);
and U6595 (N_6595,N_5710,N_4627);
xnor U6596 (N_6596,N_5317,N_5218);
and U6597 (N_6597,N_4278,N_4864);
and U6598 (N_6598,N_4103,N_4377);
nor U6599 (N_6599,N_5227,N_5417);
or U6600 (N_6600,N_4565,N_4180);
xnor U6601 (N_6601,N_5240,N_4612);
and U6602 (N_6602,N_5178,N_5597);
and U6603 (N_6603,N_4639,N_4504);
nor U6604 (N_6604,N_5890,N_5816);
xnor U6605 (N_6605,N_4681,N_5909);
or U6606 (N_6606,N_5545,N_5636);
nand U6607 (N_6607,N_4244,N_4790);
and U6608 (N_6608,N_5266,N_4095);
or U6609 (N_6609,N_4711,N_4782);
or U6610 (N_6610,N_5380,N_4484);
nand U6611 (N_6611,N_4159,N_4316);
xor U6612 (N_6612,N_4857,N_4842);
or U6613 (N_6613,N_5893,N_4553);
nand U6614 (N_6614,N_5768,N_4926);
or U6615 (N_6615,N_5991,N_4021);
nor U6616 (N_6616,N_5278,N_5513);
and U6617 (N_6617,N_5895,N_5312);
xnor U6618 (N_6618,N_4440,N_5586);
nor U6619 (N_6619,N_5137,N_4976);
nand U6620 (N_6620,N_4411,N_4946);
and U6621 (N_6621,N_5876,N_5557);
or U6622 (N_6622,N_4700,N_5564);
nor U6623 (N_6623,N_5518,N_4125);
or U6624 (N_6624,N_4850,N_5525);
and U6625 (N_6625,N_5569,N_4242);
nand U6626 (N_6626,N_5817,N_5541);
xor U6627 (N_6627,N_4539,N_4537);
or U6628 (N_6628,N_5135,N_4889);
nor U6629 (N_6629,N_4383,N_4326);
and U6630 (N_6630,N_5124,N_4032);
nor U6631 (N_6631,N_5037,N_5264);
or U6632 (N_6632,N_5679,N_5249);
xor U6633 (N_6633,N_4257,N_4020);
nor U6634 (N_6634,N_5198,N_4057);
xor U6635 (N_6635,N_5376,N_5614);
or U6636 (N_6636,N_5466,N_5592);
nand U6637 (N_6637,N_4549,N_5302);
nor U6638 (N_6638,N_4301,N_5833);
nor U6639 (N_6639,N_4810,N_4660);
or U6640 (N_6640,N_5837,N_4670);
or U6641 (N_6641,N_4302,N_4370);
nor U6642 (N_6642,N_4720,N_5122);
nor U6643 (N_6643,N_4015,N_5250);
nand U6644 (N_6644,N_4573,N_4219);
or U6645 (N_6645,N_5655,N_4448);
and U6646 (N_6646,N_5032,N_4933);
nand U6647 (N_6647,N_4954,N_5468);
and U6648 (N_6648,N_5634,N_5434);
nor U6649 (N_6649,N_4635,N_5880);
and U6650 (N_6650,N_4932,N_4237);
or U6651 (N_6651,N_5325,N_5382);
nand U6652 (N_6652,N_5507,N_4294);
nor U6653 (N_6653,N_5460,N_5857);
or U6654 (N_6654,N_5436,N_4892);
nand U6655 (N_6655,N_4428,N_4153);
or U6656 (N_6656,N_5576,N_5701);
nor U6657 (N_6657,N_4836,N_4210);
nand U6658 (N_6658,N_5259,N_4548);
nand U6659 (N_6659,N_4193,N_4140);
nand U6660 (N_6660,N_5245,N_4804);
nand U6661 (N_6661,N_4432,N_5413);
or U6662 (N_6662,N_4838,N_4493);
or U6663 (N_6663,N_4141,N_4460);
and U6664 (N_6664,N_5599,N_4259);
nor U6665 (N_6665,N_5702,N_5373);
nor U6666 (N_6666,N_5733,N_5958);
and U6667 (N_6667,N_4369,N_4104);
and U6668 (N_6668,N_5199,N_5174);
nand U6669 (N_6669,N_4420,N_4414);
or U6670 (N_6670,N_5889,N_4753);
or U6671 (N_6671,N_4740,N_4374);
nor U6672 (N_6672,N_5810,N_4997);
or U6673 (N_6673,N_4365,N_5937);
nand U6674 (N_6674,N_5322,N_4952);
and U6675 (N_6675,N_4331,N_5967);
and U6676 (N_6676,N_5700,N_4515);
and U6677 (N_6677,N_4069,N_5050);
or U6678 (N_6678,N_4256,N_4265);
and U6679 (N_6679,N_4162,N_5306);
nor U6680 (N_6680,N_4865,N_4296);
or U6681 (N_6681,N_4422,N_4703);
nand U6682 (N_6682,N_4483,N_5095);
and U6683 (N_6683,N_4013,N_4920);
nor U6684 (N_6684,N_5996,N_4806);
or U6685 (N_6685,N_4717,N_4404);
nand U6686 (N_6686,N_5276,N_5066);
nand U6687 (N_6687,N_5758,N_4727);
nand U6688 (N_6688,N_5718,N_5797);
or U6689 (N_6689,N_5363,N_5130);
nand U6690 (N_6690,N_4873,N_5261);
nand U6691 (N_6691,N_4828,N_4643);
nand U6692 (N_6692,N_4060,N_4899);
nor U6693 (N_6693,N_4906,N_4572);
and U6694 (N_6694,N_5277,N_4593);
nor U6695 (N_6695,N_5715,N_5638);
or U6696 (N_6696,N_4299,N_5342);
nor U6697 (N_6697,N_4467,N_4834);
nor U6698 (N_6698,N_5796,N_5191);
nand U6699 (N_6699,N_5483,N_4138);
nor U6700 (N_6700,N_5108,N_4328);
or U6701 (N_6701,N_4267,N_5451);
nor U6702 (N_6702,N_4691,N_4567);
nor U6703 (N_6703,N_5369,N_5033);
nor U6704 (N_6704,N_5942,N_5353);
nand U6705 (N_6705,N_4315,N_5387);
or U6706 (N_6706,N_4649,N_4992);
nor U6707 (N_6707,N_5926,N_5693);
and U6708 (N_6708,N_5791,N_4847);
or U6709 (N_6709,N_4764,N_4770);
or U6710 (N_6710,N_4769,N_4239);
nand U6711 (N_6711,N_5136,N_5689);
nand U6712 (N_6712,N_4789,N_4238);
xor U6713 (N_6713,N_4000,N_4430);
nand U6714 (N_6714,N_4625,N_5775);
and U6715 (N_6715,N_5309,N_4689);
nor U6716 (N_6716,N_4561,N_4014);
nand U6717 (N_6717,N_5970,N_4900);
and U6718 (N_6718,N_5008,N_4332);
nor U6719 (N_6719,N_4402,N_4128);
nand U6720 (N_6720,N_4190,N_4666);
or U6721 (N_6721,N_4139,N_4752);
nor U6722 (N_6722,N_5925,N_4487);
or U6723 (N_6723,N_5006,N_4385);
xor U6724 (N_6724,N_5932,N_4100);
or U6725 (N_6725,N_4468,N_4091);
and U6726 (N_6726,N_5506,N_5385);
and U6727 (N_6727,N_5681,N_5498);
nor U6728 (N_6728,N_5976,N_4684);
and U6729 (N_6729,N_5158,N_4698);
xor U6730 (N_6730,N_4801,N_5216);
xnor U6731 (N_6731,N_4075,N_5458);
nor U6732 (N_6732,N_5196,N_5075);
and U6733 (N_6733,N_4995,N_5532);
and U6734 (N_6734,N_4148,N_4435);
and U6735 (N_6735,N_5059,N_4273);
or U6736 (N_6736,N_5086,N_5756);
nand U6737 (N_6737,N_4401,N_4082);
nor U6738 (N_6738,N_5719,N_5285);
xnor U6739 (N_6739,N_5224,N_4064);
xor U6740 (N_6740,N_4746,N_4350);
or U6741 (N_6741,N_5962,N_5898);
nor U6742 (N_6742,N_5461,N_4225);
or U6743 (N_6743,N_4320,N_5146);
nor U6744 (N_6744,N_5904,N_4646);
nor U6745 (N_6745,N_4270,N_5594);
or U6746 (N_6746,N_4362,N_4914);
or U6747 (N_6747,N_4559,N_4474);
or U6748 (N_6748,N_4602,N_4538);
or U6749 (N_6749,N_4688,N_5567);
nor U6750 (N_6750,N_5871,N_5528);
nor U6751 (N_6751,N_5028,N_4169);
and U6752 (N_6752,N_4207,N_4758);
nand U6753 (N_6753,N_5502,N_5961);
nand U6754 (N_6754,N_5239,N_5243);
nor U6755 (N_6755,N_4728,N_5590);
nor U6756 (N_6756,N_5781,N_4944);
or U6757 (N_6757,N_4282,N_4621);
nor U6758 (N_6758,N_5007,N_4061);
and U6759 (N_6759,N_4090,N_5921);
nand U6760 (N_6760,N_4062,N_4718);
and U6761 (N_6761,N_5656,N_4558);
or U6762 (N_6762,N_4215,N_4525);
nand U6763 (N_6763,N_5040,N_5727);
or U6764 (N_6764,N_5405,N_5897);
xor U6765 (N_6765,N_4574,N_5121);
and U6766 (N_6766,N_4518,N_5626);
nand U6767 (N_6767,N_4695,N_4735);
or U6768 (N_6768,N_5537,N_4527);
xnor U6769 (N_6769,N_5262,N_5213);
nor U6770 (N_6770,N_4918,N_4667);
nand U6771 (N_6771,N_5029,N_4184);
and U6772 (N_6772,N_4808,N_4520);
or U6773 (N_6773,N_5042,N_5902);
or U6774 (N_6774,N_4098,N_4977);
or U6775 (N_6775,N_5253,N_4449);
nand U6776 (N_6776,N_4234,N_4434);
nor U6777 (N_6777,N_4563,N_5023);
and U6778 (N_6778,N_5888,N_5172);
xor U6779 (N_6779,N_5324,N_4957);
xnor U6780 (N_6780,N_4165,N_5635);
or U6781 (N_6781,N_4719,N_4715);
nand U6782 (N_6782,N_4185,N_5587);
and U6783 (N_6783,N_4280,N_5393);
and U6784 (N_6784,N_4682,N_5948);
nand U6785 (N_6785,N_4107,N_5699);
nor U6786 (N_6786,N_4766,N_4473);
and U6787 (N_6787,N_5508,N_5664);
and U6788 (N_6788,N_4743,N_4480);
xnor U6789 (N_6789,N_4785,N_5187);
nor U6790 (N_6790,N_5531,N_4772);
and U6791 (N_6791,N_5247,N_4359);
xor U6792 (N_6792,N_5204,N_4112);
nor U6793 (N_6793,N_5254,N_4475);
xor U6794 (N_6794,N_5786,N_4592);
nor U6795 (N_6795,N_5492,N_4393);
nor U6796 (N_6796,N_5225,N_4915);
nor U6797 (N_6797,N_4405,N_5737);
or U6798 (N_6798,N_5869,N_4629);
nand U6799 (N_6799,N_4529,N_4211);
nand U6800 (N_6800,N_4472,N_4780);
and U6801 (N_6801,N_5432,N_5232);
or U6802 (N_6802,N_5128,N_5868);
nand U6803 (N_6803,N_5200,N_4693);
and U6804 (N_6804,N_4297,N_4010);
and U6805 (N_6805,N_4343,N_5505);
or U6806 (N_6806,N_4871,N_4226);
and U6807 (N_6807,N_4007,N_5551);
nand U6808 (N_6808,N_5201,N_4202);
nand U6809 (N_6809,N_4084,N_4323);
or U6810 (N_6810,N_5157,N_4710);
and U6811 (N_6811,N_4055,N_4394);
and U6812 (N_6812,N_4845,N_5326);
nor U6813 (N_6813,N_4998,N_5882);
or U6814 (N_6814,N_4341,N_5145);
nor U6815 (N_6815,N_4288,N_4454);
nand U6816 (N_6816,N_4598,N_5133);
nor U6817 (N_6817,N_4778,N_4481);
nand U6818 (N_6818,N_4387,N_4111);
nor U6819 (N_6819,N_5051,N_4223);
nor U6820 (N_6820,N_5517,N_5570);
and U6821 (N_6821,N_4023,N_4118);
nor U6822 (N_6822,N_4397,N_5288);
or U6823 (N_6823,N_4550,N_5930);
nand U6824 (N_6824,N_4702,N_4287);
xor U6825 (N_6825,N_5352,N_4217);
nor U6826 (N_6826,N_5368,N_4988);
nand U6827 (N_6827,N_4841,N_4661);
and U6828 (N_6828,N_4852,N_4391);
or U6829 (N_6829,N_4133,N_4840);
nor U6830 (N_6830,N_5220,N_4108);
or U6831 (N_6831,N_5371,N_5192);
xor U6832 (N_6832,N_4441,N_5726);
and U6833 (N_6833,N_5304,N_4762);
xnor U6834 (N_6834,N_5419,N_5444);
or U6835 (N_6835,N_5034,N_5246);
and U6836 (N_6836,N_5753,N_4826);
or U6837 (N_6837,N_4818,N_4255);
nor U6838 (N_6838,N_4949,N_4973);
nor U6839 (N_6839,N_4406,N_4399);
nor U6840 (N_6840,N_5499,N_5861);
nor U6841 (N_6841,N_5298,N_5154);
nor U6842 (N_6842,N_5931,N_4167);
nand U6843 (N_6843,N_5927,N_4916);
and U6844 (N_6844,N_5856,N_4531);
nand U6845 (N_6845,N_5142,N_5698);
xnor U6846 (N_6846,N_5208,N_4747);
nor U6847 (N_6847,N_4347,N_4543);
and U6848 (N_6848,N_5404,N_5345);
and U6849 (N_6849,N_4908,N_5202);
or U6850 (N_6850,N_5041,N_4856);
nand U6851 (N_6851,N_5441,N_5683);
nand U6852 (N_6852,N_4308,N_4570);
and U6853 (N_6853,N_5790,N_4177);
xor U6854 (N_6854,N_4079,N_5670);
or U6855 (N_6855,N_4089,N_5665);
and U6856 (N_6856,N_4266,N_5190);
or U6857 (N_6857,N_5223,N_4844);
or U6858 (N_6858,N_4008,N_5575);
nand U6859 (N_6859,N_5226,N_4786);
or U6860 (N_6860,N_4419,N_5301);
nor U6861 (N_6861,N_4771,N_5907);
nor U6862 (N_6862,N_5650,N_4378);
nor U6863 (N_6863,N_5091,N_5987);
nor U6864 (N_6864,N_4423,N_4389);
nor U6865 (N_6865,N_5854,N_5530);
xnor U6866 (N_6866,N_5913,N_4601);
or U6867 (N_6867,N_4421,N_4517);
nor U6868 (N_6868,N_5941,N_4577);
or U6869 (N_6869,N_5743,N_4588);
xor U6870 (N_6870,N_5002,N_5782);
and U6871 (N_6871,N_4478,N_5995);
nand U6872 (N_6872,N_5984,N_5762);
or U6873 (N_6873,N_5485,N_5646);
and U6874 (N_6874,N_5465,N_5036);
nor U6875 (N_6875,N_4337,N_4749);
nand U6876 (N_6876,N_4673,N_4955);
and U6877 (N_6877,N_4942,N_5480);
and U6878 (N_6878,N_5248,N_4905);
or U6879 (N_6879,N_5993,N_5054);
or U6880 (N_6880,N_5370,N_4783);
nand U6881 (N_6881,N_5134,N_5222);
and U6882 (N_6882,N_5315,N_5777);
and U6883 (N_6883,N_5176,N_5581);
or U6884 (N_6884,N_4985,N_5283);
nand U6885 (N_6885,N_5280,N_4344);
nand U6886 (N_6886,N_5627,N_4597);
nand U6887 (N_6887,N_4158,N_4078);
nand U6888 (N_6888,N_4983,N_4443);
xnor U6889 (N_6889,N_5269,N_5736);
or U6890 (N_6890,N_4712,N_5060);
nor U6891 (N_6891,N_5470,N_4867);
and U6892 (N_6892,N_5017,N_4181);
nand U6893 (N_6893,N_5081,N_4589);
xnor U6894 (N_6894,N_5598,N_5870);
nor U6895 (N_6895,N_5411,N_5221);
or U6896 (N_6896,N_4805,N_4648);
xor U6897 (N_6897,N_5792,N_4043);
nand U6898 (N_6898,N_4909,N_5238);
xor U6899 (N_6899,N_4894,N_5456);
nand U6900 (N_6900,N_5430,N_5547);
xor U6901 (N_6901,N_5631,N_5094);
xnor U6902 (N_6902,N_5523,N_5399);
or U6903 (N_6903,N_5705,N_5540);
nor U6904 (N_6904,N_4033,N_4101);
nor U6905 (N_6905,N_4987,N_4951);
nor U6906 (N_6906,N_5982,N_5625);
or U6907 (N_6907,N_5728,N_4641);
nand U6908 (N_6908,N_5521,N_4677);
xor U6909 (N_6909,N_5449,N_5338);
nor U6910 (N_6910,N_4230,N_4890);
nand U6911 (N_6911,N_5894,N_4067);
nor U6912 (N_6912,N_5675,N_4705);
or U6913 (N_6913,N_4403,N_4221);
nand U6914 (N_6914,N_4446,N_4994);
xnor U6915 (N_6915,N_4506,N_5945);
nand U6916 (N_6916,N_4619,N_5811);
xor U6917 (N_6917,N_4895,N_5565);
xor U6918 (N_6918,N_4776,N_4289);
or U6919 (N_6919,N_4002,N_4379);
xor U6920 (N_6920,N_4613,N_4250);
nand U6921 (N_6921,N_4514,N_5078);
and U6922 (N_6922,N_5127,N_5808);
nor U6923 (N_6923,N_4669,N_5476);
xnor U6924 (N_6924,N_5678,N_5690);
nand U6925 (N_6925,N_4680,N_4714);
and U6926 (N_6926,N_5390,N_5068);
and U6927 (N_6927,N_4149,N_5175);
nand U6928 (N_6928,N_4134,N_5554);
nand U6929 (N_6929,N_5548,N_4122);
nor U6930 (N_6930,N_4011,N_5847);
and U6931 (N_6931,N_4833,N_4870);
nor U6932 (N_6932,N_5988,N_5935);
nand U6933 (N_6933,N_5713,N_5788);
and U6934 (N_6934,N_4459,N_4309);
and U6935 (N_6935,N_4005,N_5410);
xor U6936 (N_6936,N_5310,N_4802);
and U6937 (N_6937,N_4186,N_4413);
xor U6938 (N_6938,N_5986,N_5985);
or U6939 (N_6939,N_5510,N_5343);
xor U6940 (N_6940,N_4361,N_4623);
nand U6941 (N_6941,N_4489,N_4620);
xor U6942 (N_6942,N_4355,N_5150);
and U6943 (N_6943,N_5167,N_5859);
nand U6944 (N_6944,N_5155,N_4809);
nand U6945 (N_6945,N_5972,N_5606);
or U6946 (N_6946,N_4313,N_5215);
and U6947 (N_6947,N_5922,N_4345);
and U6948 (N_6948,N_5772,N_4458);
or U6949 (N_6949,N_4788,N_4174);
and U6950 (N_6950,N_4291,N_4048);
nor U6951 (N_6951,N_4524,N_4310);
xor U6952 (N_6952,N_5629,N_5754);
nor U6953 (N_6953,N_4729,N_4093);
nor U6954 (N_6954,N_5327,N_4540);
nor U6955 (N_6955,N_5063,N_5866);
xor U6956 (N_6956,N_5563,N_4072);
or U6957 (N_6957,N_4099,N_4388);
or U6958 (N_6958,N_4663,N_5749);
nand U6959 (N_6959,N_5905,N_5424);
nor U6960 (N_6960,N_4547,N_5377);
or U6961 (N_6961,N_4041,N_4263);
xnor U6962 (N_6962,N_5751,N_4874);
nor U6963 (N_6963,N_4327,N_5509);
or U6964 (N_6964,N_4960,N_4437);
nor U6965 (N_6965,N_5471,N_5125);
nor U6966 (N_6966,N_5348,N_5048);
nand U6967 (N_6967,N_4922,N_4216);
or U6968 (N_6968,N_5403,N_5148);
and U6969 (N_6969,N_4427,N_5265);
nand U6970 (N_6970,N_4907,N_4395);
nor U6971 (N_6971,N_4351,N_5359);
or U6972 (N_6972,N_4893,N_5445);
nor U6973 (N_6973,N_5787,N_4182);
and U6974 (N_6974,N_4644,N_4290);
nor U6975 (N_6975,N_5544,N_4116);
nand U6976 (N_6976,N_5633,N_5892);
and U6977 (N_6977,N_4966,N_4214);
and U6978 (N_6978,N_5550,N_4566);
and U6979 (N_6979,N_4713,N_4046);
nor U6980 (N_6980,N_5940,N_5855);
nand U6981 (N_6981,N_4526,N_4463);
nand U6982 (N_6982,N_4605,N_5152);
nand U6983 (N_6983,N_5716,N_5161);
nand U6984 (N_6984,N_4324,N_4371);
and U6985 (N_6985,N_5236,N_5896);
and U6986 (N_6986,N_4456,N_4651);
nand U6987 (N_6987,N_5755,N_4683);
or U6988 (N_6988,N_5707,N_5652);
and U6989 (N_6989,N_5739,N_5822);
nor U6990 (N_6990,N_5275,N_4672);
and U6991 (N_6991,N_5766,N_5803);
or U6992 (N_6992,N_5752,N_5396);
nor U6993 (N_6993,N_4608,N_5457);
and U6994 (N_6994,N_4912,N_4554);
or U6995 (N_6995,N_5765,N_4491);
or U6996 (N_6996,N_4224,N_5286);
nor U6997 (N_6997,N_4959,N_4304);
nand U6998 (N_6998,N_4607,N_5647);
and U6999 (N_6999,N_5601,N_5596);
and U7000 (N_7000,N_5033,N_4880);
nand U7001 (N_7001,N_5572,N_5566);
nor U7002 (N_7002,N_5686,N_4637);
nand U7003 (N_7003,N_4445,N_4429);
nor U7004 (N_7004,N_4182,N_4606);
nor U7005 (N_7005,N_5870,N_4340);
nor U7006 (N_7006,N_5373,N_4769);
or U7007 (N_7007,N_4762,N_4536);
nand U7008 (N_7008,N_5793,N_5351);
nor U7009 (N_7009,N_5721,N_5002);
and U7010 (N_7010,N_4541,N_5992);
nor U7011 (N_7011,N_5177,N_4680);
xor U7012 (N_7012,N_5507,N_5381);
nand U7013 (N_7013,N_4751,N_4802);
xnor U7014 (N_7014,N_4301,N_4742);
and U7015 (N_7015,N_4914,N_5579);
and U7016 (N_7016,N_5286,N_5729);
nor U7017 (N_7017,N_5729,N_5927);
or U7018 (N_7018,N_5529,N_5757);
xor U7019 (N_7019,N_4477,N_5788);
or U7020 (N_7020,N_5069,N_4136);
and U7021 (N_7021,N_5273,N_4549);
nand U7022 (N_7022,N_5917,N_5074);
nor U7023 (N_7023,N_4811,N_5167);
xnor U7024 (N_7024,N_4193,N_5327);
nand U7025 (N_7025,N_5714,N_4863);
nand U7026 (N_7026,N_5181,N_5924);
and U7027 (N_7027,N_5884,N_4428);
nor U7028 (N_7028,N_5773,N_4063);
and U7029 (N_7029,N_5939,N_4362);
nor U7030 (N_7030,N_5714,N_4605);
or U7031 (N_7031,N_4138,N_4182);
or U7032 (N_7032,N_5426,N_5228);
nor U7033 (N_7033,N_4077,N_5589);
nor U7034 (N_7034,N_5110,N_5696);
and U7035 (N_7035,N_5944,N_4294);
nand U7036 (N_7036,N_5608,N_4014);
and U7037 (N_7037,N_4659,N_4430);
or U7038 (N_7038,N_5380,N_4621);
nand U7039 (N_7039,N_5707,N_5546);
nand U7040 (N_7040,N_4224,N_4859);
and U7041 (N_7041,N_4206,N_4632);
and U7042 (N_7042,N_5316,N_5096);
and U7043 (N_7043,N_5772,N_5388);
nor U7044 (N_7044,N_5466,N_4830);
xor U7045 (N_7045,N_4099,N_5879);
or U7046 (N_7046,N_5533,N_4473);
or U7047 (N_7047,N_5332,N_4480);
or U7048 (N_7048,N_5266,N_5329);
or U7049 (N_7049,N_4165,N_4849);
nor U7050 (N_7050,N_5529,N_4277);
or U7051 (N_7051,N_5522,N_5753);
nor U7052 (N_7052,N_5031,N_5284);
and U7053 (N_7053,N_5064,N_5865);
or U7054 (N_7054,N_4656,N_4475);
nand U7055 (N_7055,N_4251,N_4435);
nand U7056 (N_7056,N_4235,N_5969);
or U7057 (N_7057,N_4593,N_5410);
or U7058 (N_7058,N_5866,N_4361);
nand U7059 (N_7059,N_4812,N_4864);
or U7060 (N_7060,N_4554,N_4743);
xnor U7061 (N_7061,N_4002,N_4514);
nor U7062 (N_7062,N_5761,N_4323);
nor U7063 (N_7063,N_5755,N_4061);
nand U7064 (N_7064,N_4118,N_4430);
nor U7065 (N_7065,N_4018,N_4664);
nor U7066 (N_7066,N_4652,N_4294);
and U7067 (N_7067,N_4341,N_4413);
or U7068 (N_7068,N_4972,N_5779);
nor U7069 (N_7069,N_4640,N_4686);
nand U7070 (N_7070,N_4181,N_5810);
or U7071 (N_7071,N_5108,N_5677);
nand U7072 (N_7072,N_5091,N_5322);
nand U7073 (N_7073,N_5091,N_4610);
or U7074 (N_7074,N_4446,N_4584);
xnor U7075 (N_7075,N_4764,N_5185);
nor U7076 (N_7076,N_4381,N_5816);
nand U7077 (N_7077,N_5556,N_4357);
or U7078 (N_7078,N_5130,N_4549);
nor U7079 (N_7079,N_5595,N_5124);
nor U7080 (N_7080,N_4104,N_4589);
nor U7081 (N_7081,N_5275,N_5315);
or U7082 (N_7082,N_4356,N_5182);
xnor U7083 (N_7083,N_4451,N_5126);
nor U7084 (N_7084,N_4238,N_4222);
nor U7085 (N_7085,N_5515,N_4098);
nor U7086 (N_7086,N_4741,N_5222);
nand U7087 (N_7087,N_4532,N_4154);
and U7088 (N_7088,N_5235,N_4313);
nor U7089 (N_7089,N_4439,N_4432);
or U7090 (N_7090,N_4147,N_5868);
and U7091 (N_7091,N_5080,N_5473);
nand U7092 (N_7092,N_4009,N_4069);
nand U7093 (N_7093,N_4691,N_5878);
xnor U7094 (N_7094,N_5370,N_5513);
and U7095 (N_7095,N_4145,N_5923);
nand U7096 (N_7096,N_5355,N_4646);
and U7097 (N_7097,N_5341,N_5281);
xnor U7098 (N_7098,N_4487,N_5804);
or U7099 (N_7099,N_5274,N_5003);
and U7100 (N_7100,N_5397,N_4148);
nor U7101 (N_7101,N_5930,N_5524);
and U7102 (N_7102,N_4380,N_4130);
xor U7103 (N_7103,N_4859,N_4556);
nand U7104 (N_7104,N_4322,N_5384);
nor U7105 (N_7105,N_4646,N_5223);
nand U7106 (N_7106,N_4435,N_5440);
and U7107 (N_7107,N_4999,N_5795);
or U7108 (N_7108,N_4722,N_5523);
xnor U7109 (N_7109,N_5301,N_5452);
xnor U7110 (N_7110,N_4319,N_5557);
nand U7111 (N_7111,N_5064,N_4651);
nor U7112 (N_7112,N_5739,N_5126);
or U7113 (N_7113,N_5160,N_5769);
nor U7114 (N_7114,N_5524,N_4951);
nand U7115 (N_7115,N_5960,N_4828);
or U7116 (N_7116,N_4341,N_4180);
nand U7117 (N_7117,N_5326,N_4774);
nor U7118 (N_7118,N_4515,N_5379);
nor U7119 (N_7119,N_4535,N_4102);
and U7120 (N_7120,N_4794,N_4739);
nor U7121 (N_7121,N_5258,N_5213);
or U7122 (N_7122,N_5934,N_5360);
nand U7123 (N_7123,N_4997,N_5193);
and U7124 (N_7124,N_5062,N_4251);
nor U7125 (N_7125,N_4489,N_5549);
nor U7126 (N_7126,N_5092,N_5097);
nor U7127 (N_7127,N_4920,N_5807);
and U7128 (N_7128,N_5708,N_5934);
xnor U7129 (N_7129,N_4131,N_5264);
or U7130 (N_7130,N_5785,N_5157);
or U7131 (N_7131,N_5092,N_5029);
and U7132 (N_7132,N_4946,N_4663);
and U7133 (N_7133,N_4438,N_4611);
or U7134 (N_7134,N_4614,N_5347);
or U7135 (N_7135,N_5357,N_5070);
nor U7136 (N_7136,N_5943,N_4994);
and U7137 (N_7137,N_4732,N_5164);
nand U7138 (N_7138,N_5856,N_5906);
or U7139 (N_7139,N_5289,N_5724);
nor U7140 (N_7140,N_5540,N_5106);
nand U7141 (N_7141,N_4119,N_5386);
xor U7142 (N_7142,N_5352,N_5215);
and U7143 (N_7143,N_5748,N_4610);
and U7144 (N_7144,N_4919,N_4425);
and U7145 (N_7145,N_5785,N_5166);
nor U7146 (N_7146,N_5640,N_4836);
xor U7147 (N_7147,N_5821,N_4249);
or U7148 (N_7148,N_5190,N_5159);
xor U7149 (N_7149,N_4699,N_4717);
nand U7150 (N_7150,N_4957,N_5565);
and U7151 (N_7151,N_4852,N_5048);
and U7152 (N_7152,N_5022,N_4043);
xnor U7153 (N_7153,N_4710,N_5156);
nor U7154 (N_7154,N_5106,N_5096);
and U7155 (N_7155,N_4464,N_5173);
and U7156 (N_7156,N_5782,N_4042);
nand U7157 (N_7157,N_4271,N_5650);
or U7158 (N_7158,N_4455,N_4995);
or U7159 (N_7159,N_4189,N_5591);
nor U7160 (N_7160,N_4484,N_4136);
and U7161 (N_7161,N_5821,N_4981);
and U7162 (N_7162,N_4432,N_5110);
and U7163 (N_7163,N_5039,N_5574);
nand U7164 (N_7164,N_4462,N_4090);
and U7165 (N_7165,N_5471,N_4051);
nor U7166 (N_7166,N_4406,N_4470);
nand U7167 (N_7167,N_5718,N_5561);
nor U7168 (N_7168,N_4170,N_4261);
and U7169 (N_7169,N_4743,N_5069);
and U7170 (N_7170,N_5619,N_4048);
and U7171 (N_7171,N_5684,N_4796);
and U7172 (N_7172,N_5481,N_4292);
and U7173 (N_7173,N_4040,N_5712);
nor U7174 (N_7174,N_4066,N_4367);
nand U7175 (N_7175,N_5049,N_5345);
or U7176 (N_7176,N_4534,N_4435);
nand U7177 (N_7177,N_4549,N_5301);
or U7178 (N_7178,N_5387,N_4170);
or U7179 (N_7179,N_5182,N_5478);
or U7180 (N_7180,N_4836,N_4751);
or U7181 (N_7181,N_5002,N_4633);
and U7182 (N_7182,N_5642,N_4028);
or U7183 (N_7183,N_5386,N_4283);
nand U7184 (N_7184,N_4603,N_4357);
nand U7185 (N_7185,N_5061,N_5177);
or U7186 (N_7186,N_4141,N_5334);
xnor U7187 (N_7187,N_4868,N_5610);
and U7188 (N_7188,N_4223,N_4853);
and U7189 (N_7189,N_4286,N_5482);
nor U7190 (N_7190,N_5420,N_4374);
and U7191 (N_7191,N_4964,N_4908);
nand U7192 (N_7192,N_4441,N_4874);
and U7193 (N_7193,N_5547,N_4671);
nand U7194 (N_7194,N_4190,N_4162);
nand U7195 (N_7195,N_5062,N_5000);
nor U7196 (N_7196,N_4074,N_5967);
nand U7197 (N_7197,N_5765,N_4019);
nor U7198 (N_7198,N_5590,N_4328);
or U7199 (N_7199,N_5556,N_5676);
or U7200 (N_7200,N_4461,N_4888);
xor U7201 (N_7201,N_4209,N_4056);
or U7202 (N_7202,N_5529,N_4216);
nand U7203 (N_7203,N_5111,N_4316);
nor U7204 (N_7204,N_4178,N_4639);
and U7205 (N_7205,N_5059,N_5263);
nor U7206 (N_7206,N_4102,N_5657);
or U7207 (N_7207,N_4571,N_5906);
and U7208 (N_7208,N_5027,N_5813);
nor U7209 (N_7209,N_5449,N_4387);
nor U7210 (N_7210,N_5700,N_4925);
nand U7211 (N_7211,N_5930,N_4568);
or U7212 (N_7212,N_4011,N_4281);
or U7213 (N_7213,N_4279,N_5099);
xnor U7214 (N_7214,N_4178,N_5866);
and U7215 (N_7215,N_5034,N_4068);
and U7216 (N_7216,N_5145,N_4656);
and U7217 (N_7217,N_4132,N_5899);
nor U7218 (N_7218,N_4791,N_4876);
and U7219 (N_7219,N_4094,N_4040);
nand U7220 (N_7220,N_5841,N_4521);
nand U7221 (N_7221,N_4778,N_4316);
nor U7222 (N_7222,N_4464,N_5063);
or U7223 (N_7223,N_5075,N_4203);
or U7224 (N_7224,N_4176,N_4805);
or U7225 (N_7225,N_4512,N_5507);
nor U7226 (N_7226,N_4195,N_5148);
nor U7227 (N_7227,N_5485,N_4660);
nor U7228 (N_7228,N_5945,N_4979);
or U7229 (N_7229,N_4796,N_4216);
or U7230 (N_7230,N_5972,N_5588);
xnor U7231 (N_7231,N_4738,N_5926);
nor U7232 (N_7232,N_5206,N_5798);
xor U7233 (N_7233,N_4899,N_5703);
and U7234 (N_7234,N_4726,N_4164);
and U7235 (N_7235,N_5081,N_4007);
nand U7236 (N_7236,N_5404,N_5981);
and U7237 (N_7237,N_4630,N_4863);
or U7238 (N_7238,N_5317,N_5827);
or U7239 (N_7239,N_5845,N_5400);
and U7240 (N_7240,N_4333,N_4306);
and U7241 (N_7241,N_4710,N_4036);
nor U7242 (N_7242,N_4248,N_5107);
nand U7243 (N_7243,N_4091,N_4918);
or U7244 (N_7244,N_4364,N_5133);
and U7245 (N_7245,N_4896,N_5222);
and U7246 (N_7246,N_4649,N_4579);
and U7247 (N_7247,N_5027,N_5259);
and U7248 (N_7248,N_4335,N_5328);
or U7249 (N_7249,N_5856,N_4480);
nand U7250 (N_7250,N_4265,N_4104);
and U7251 (N_7251,N_5815,N_4097);
and U7252 (N_7252,N_4933,N_5566);
xor U7253 (N_7253,N_5022,N_5502);
and U7254 (N_7254,N_4382,N_5691);
or U7255 (N_7255,N_4805,N_4404);
nor U7256 (N_7256,N_4704,N_5613);
nor U7257 (N_7257,N_4266,N_5737);
and U7258 (N_7258,N_4823,N_4561);
and U7259 (N_7259,N_4528,N_4450);
and U7260 (N_7260,N_5620,N_5534);
or U7261 (N_7261,N_5880,N_4448);
nand U7262 (N_7262,N_5444,N_4354);
and U7263 (N_7263,N_4910,N_5638);
and U7264 (N_7264,N_5842,N_5090);
or U7265 (N_7265,N_5168,N_5740);
and U7266 (N_7266,N_4365,N_4018);
and U7267 (N_7267,N_4133,N_5759);
and U7268 (N_7268,N_5202,N_5493);
and U7269 (N_7269,N_5938,N_4164);
and U7270 (N_7270,N_5583,N_4836);
or U7271 (N_7271,N_5601,N_5812);
nor U7272 (N_7272,N_5930,N_4736);
and U7273 (N_7273,N_4095,N_4869);
nand U7274 (N_7274,N_5272,N_4607);
and U7275 (N_7275,N_5150,N_4696);
nor U7276 (N_7276,N_4762,N_4235);
or U7277 (N_7277,N_4410,N_5346);
and U7278 (N_7278,N_4989,N_4865);
or U7279 (N_7279,N_5713,N_4559);
and U7280 (N_7280,N_5296,N_5958);
or U7281 (N_7281,N_4085,N_5128);
or U7282 (N_7282,N_4660,N_5952);
and U7283 (N_7283,N_5152,N_4572);
nand U7284 (N_7284,N_5409,N_4532);
nor U7285 (N_7285,N_5063,N_5745);
or U7286 (N_7286,N_5548,N_5635);
nor U7287 (N_7287,N_5766,N_4050);
nor U7288 (N_7288,N_5486,N_4128);
nor U7289 (N_7289,N_5801,N_4587);
and U7290 (N_7290,N_4172,N_5614);
xnor U7291 (N_7291,N_5384,N_5580);
nand U7292 (N_7292,N_5811,N_4870);
nor U7293 (N_7293,N_5116,N_5412);
xor U7294 (N_7294,N_4046,N_4026);
and U7295 (N_7295,N_5796,N_5609);
nand U7296 (N_7296,N_4767,N_4812);
nor U7297 (N_7297,N_4531,N_5322);
nand U7298 (N_7298,N_4304,N_4966);
and U7299 (N_7299,N_4401,N_5339);
nand U7300 (N_7300,N_4787,N_4361);
or U7301 (N_7301,N_4306,N_4716);
and U7302 (N_7302,N_4602,N_5404);
or U7303 (N_7303,N_5690,N_5738);
nor U7304 (N_7304,N_4678,N_4760);
nand U7305 (N_7305,N_5987,N_5866);
or U7306 (N_7306,N_5670,N_4238);
or U7307 (N_7307,N_4700,N_4489);
nor U7308 (N_7308,N_4930,N_5684);
or U7309 (N_7309,N_4189,N_4130);
nand U7310 (N_7310,N_5135,N_4079);
nand U7311 (N_7311,N_5214,N_5907);
and U7312 (N_7312,N_5490,N_5175);
nand U7313 (N_7313,N_5419,N_4170);
nor U7314 (N_7314,N_4994,N_5114);
nor U7315 (N_7315,N_5920,N_4763);
and U7316 (N_7316,N_5879,N_5972);
or U7317 (N_7317,N_5384,N_5080);
nor U7318 (N_7318,N_5285,N_4049);
nor U7319 (N_7319,N_5529,N_5984);
nand U7320 (N_7320,N_5883,N_5230);
xor U7321 (N_7321,N_5840,N_5432);
or U7322 (N_7322,N_4613,N_5504);
xnor U7323 (N_7323,N_5264,N_5814);
and U7324 (N_7324,N_5937,N_4302);
and U7325 (N_7325,N_5983,N_5504);
nand U7326 (N_7326,N_4131,N_5395);
nor U7327 (N_7327,N_5986,N_5619);
nor U7328 (N_7328,N_5481,N_5158);
and U7329 (N_7329,N_5102,N_5422);
or U7330 (N_7330,N_5522,N_5490);
or U7331 (N_7331,N_4878,N_5880);
nand U7332 (N_7332,N_5414,N_4758);
and U7333 (N_7333,N_4990,N_5723);
and U7334 (N_7334,N_4384,N_4521);
nor U7335 (N_7335,N_4065,N_5064);
nor U7336 (N_7336,N_5391,N_5187);
or U7337 (N_7337,N_4774,N_5552);
nor U7338 (N_7338,N_4163,N_5387);
or U7339 (N_7339,N_5618,N_4855);
and U7340 (N_7340,N_4307,N_4423);
nor U7341 (N_7341,N_4611,N_5952);
and U7342 (N_7342,N_5728,N_4471);
nand U7343 (N_7343,N_5898,N_4369);
nor U7344 (N_7344,N_4272,N_5633);
and U7345 (N_7345,N_4295,N_5224);
and U7346 (N_7346,N_4015,N_4929);
or U7347 (N_7347,N_4064,N_5234);
or U7348 (N_7348,N_4760,N_5292);
or U7349 (N_7349,N_4557,N_4530);
nor U7350 (N_7350,N_5614,N_5057);
nor U7351 (N_7351,N_5499,N_4038);
nand U7352 (N_7352,N_4137,N_5087);
or U7353 (N_7353,N_5414,N_5000);
nor U7354 (N_7354,N_5322,N_5765);
and U7355 (N_7355,N_4992,N_4153);
nand U7356 (N_7356,N_5128,N_5964);
or U7357 (N_7357,N_4011,N_5094);
nand U7358 (N_7358,N_5176,N_4461);
xnor U7359 (N_7359,N_5544,N_5667);
and U7360 (N_7360,N_5719,N_4908);
nand U7361 (N_7361,N_4843,N_5983);
nor U7362 (N_7362,N_4864,N_4699);
nor U7363 (N_7363,N_5230,N_4661);
or U7364 (N_7364,N_4217,N_4351);
nor U7365 (N_7365,N_4180,N_4277);
or U7366 (N_7366,N_5071,N_5923);
nand U7367 (N_7367,N_4808,N_5196);
and U7368 (N_7368,N_5559,N_4996);
and U7369 (N_7369,N_4911,N_5110);
nor U7370 (N_7370,N_5720,N_5288);
nor U7371 (N_7371,N_4400,N_4340);
or U7372 (N_7372,N_4020,N_4614);
and U7373 (N_7373,N_5819,N_4583);
and U7374 (N_7374,N_5825,N_5916);
nor U7375 (N_7375,N_4631,N_4352);
and U7376 (N_7376,N_5487,N_5904);
nor U7377 (N_7377,N_5968,N_5834);
or U7378 (N_7378,N_4127,N_4964);
nor U7379 (N_7379,N_5121,N_5462);
nand U7380 (N_7380,N_5790,N_5559);
xnor U7381 (N_7381,N_4630,N_4008);
or U7382 (N_7382,N_4597,N_4371);
nor U7383 (N_7383,N_5590,N_5048);
and U7384 (N_7384,N_5158,N_5792);
nor U7385 (N_7385,N_5937,N_4641);
xnor U7386 (N_7386,N_5583,N_4521);
nor U7387 (N_7387,N_5088,N_5978);
nor U7388 (N_7388,N_5583,N_5965);
nor U7389 (N_7389,N_4372,N_4357);
and U7390 (N_7390,N_4036,N_5308);
nor U7391 (N_7391,N_5733,N_4805);
nand U7392 (N_7392,N_4176,N_5810);
or U7393 (N_7393,N_5812,N_4198);
nor U7394 (N_7394,N_4280,N_5961);
nand U7395 (N_7395,N_4798,N_4205);
nor U7396 (N_7396,N_4879,N_5719);
or U7397 (N_7397,N_4574,N_4187);
or U7398 (N_7398,N_4245,N_5616);
or U7399 (N_7399,N_5539,N_5202);
xor U7400 (N_7400,N_5205,N_4111);
xnor U7401 (N_7401,N_4184,N_4577);
and U7402 (N_7402,N_4054,N_5961);
and U7403 (N_7403,N_5886,N_4546);
or U7404 (N_7404,N_5642,N_5369);
nor U7405 (N_7405,N_5737,N_5330);
nand U7406 (N_7406,N_5341,N_4120);
nor U7407 (N_7407,N_4683,N_4062);
nand U7408 (N_7408,N_5053,N_5693);
nor U7409 (N_7409,N_5755,N_4777);
nor U7410 (N_7410,N_4208,N_4311);
nand U7411 (N_7411,N_5740,N_4158);
nor U7412 (N_7412,N_4988,N_4820);
nand U7413 (N_7413,N_4726,N_5532);
or U7414 (N_7414,N_5514,N_5416);
and U7415 (N_7415,N_4848,N_5590);
nor U7416 (N_7416,N_4415,N_5800);
nand U7417 (N_7417,N_4002,N_4533);
nand U7418 (N_7418,N_4802,N_4487);
and U7419 (N_7419,N_5001,N_5844);
xor U7420 (N_7420,N_4427,N_5317);
nand U7421 (N_7421,N_5796,N_4291);
nor U7422 (N_7422,N_4001,N_5318);
and U7423 (N_7423,N_5014,N_5476);
and U7424 (N_7424,N_5547,N_4832);
nor U7425 (N_7425,N_5864,N_4130);
xnor U7426 (N_7426,N_5843,N_4170);
nor U7427 (N_7427,N_4049,N_4836);
and U7428 (N_7428,N_4919,N_4746);
xnor U7429 (N_7429,N_4394,N_4843);
nand U7430 (N_7430,N_5131,N_4614);
xor U7431 (N_7431,N_5225,N_4627);
and U7432 (N_7432,N_5793,N_5943);
nand U7433 (N_7433,N_4170,N_4440);
or U7434 (N_7434,N_4681,N_4180);
or U7435 (N_7435,N_4331,N_4466);
nor U7436 (N_7436,N_5702,N_4147);
xnor U7437 (N_7437,N_4464,N_5077);
and U7438 (N_7438,N_4852,N_5004);
or U7439 (N_7439,N_5497,N_4601);
and U7440 (N_7440,N_5537,N_5281);
nor U7441 (N_7441,N_5506,N_5509);
nand U7442 (N_7442,N_4447,N_5741);
xnor U7443 (N_7443,N_4257,N_4506);
nand U7444 (N_7444,N_5518,N_4662);
and U7445 (N_7445,N_5983,N_5075);
nand U7446 (N_7446,N_5423,N_5819);
nand U7447 (N_7447,N_4606,N_4207);
or U7448 (N_7448,N_4908,N_5852);
nand U7449 (N_7449,N_5731,N_5946);
and U7450 (N_7450,N_4280,N_4625);
xnor U7451 (N_7451,N_5097,N_5371);
nor U7452 (N_7452,N_5746,N_5405);
nand U7453 (N_7453,N_4728,N_4771);
nand U7454 (N_7454,N_5079,N_5990);
and U7455 (N_7455,N_5976,N_5591);
xnor U7456 (N_7456,N_5557,N_4882);
or U7457 (N_7457,N_5921,N_4349);
and U7458 (N_7458,N_5181,N_4207);
and U7459 (N_7459,N_4044,N_4086);
or U7460 (N_7460,N_5178,N_4283);
and U7461 (N_7461,N_4741,N_4215);
or U7462 (N_7462,N_5599,N_4277);
nor U7463 (N_7463,N_5766,N_5630);
and U7464 (N_7464,N_5752,N_4431);
nand U7465 (N_7465,N_5732,N_5788);
nand U7466 (N_7466,N_5446,N_4375);
nand U7467 (N_7467,N_5136,N_4633);
and U7468 (N_7468,N_5434,N_4994);
nand U7469 (N_7469,N_5212,N_5620);
nor U7470 (N_7470,N_5817,N_5021);
nand U7471 (N_7471,N_4501,N_4589);
nand U7472 (N_7472,N_5379,N_4959);
nand U7473 (N_7473,N_4167,N_5473);
nand U7474 (N_7474,N_4203,N_4044);
nor U7475 (N_7475,N_5696,N_4227);
and U7476 (N_7476,N_5664,N_4185);
or U7477 (N_7477,N_4411,N_5319);
or U7478 (N_7478,N_4566,N_4371);
xor U7479 (N_7479,N_4060,N_5313);
nand U7480 (N_7480,N_5358,N_4484);
and U7481 (N_7481,N_5905,N_5918);
nor U7482 (N_7482,N_5894,N_5396);
and U7483 (N_7483,N_5864,N_4432);
or U7484 (N_7484,N_4892,N_4064);
or U7485 (N_7485,N_4299,N_4288);
xor U7486 (N_7486,N_4162,N_5968);
or U7487 (N_7487,N_5854,N_5688);
xnor U7488 (N_7488,N_5585,N_4137);
nor U7489 (N_7489,N_4432,N_5222);
or U7490 (N_7490,N_5668,N_4004);
nand U7491 (N_7491,N_5650,N_4031);
nand U7492 (N_7492,N_4882,N_4920);
nand U7493 (N_7493,N_4060,N_5876);
nand U7494 (N_7494,N_4885,N_5971);
nor U7495 (N_7495,N_4773,N_4272);
and U7496 (N_7496,N_4656,N_4097);
or U7497 (N_7497,N_4205,N_5009);
xnor U7498 (N_7498,N_4981,N_4506);
nand U7499 (N_7499,N_5386,N_4295);
or U7500 (N_7500,N_4835,N_4753);
nand U7501 (N_7501,N_4073,N_5097);
nand U7502 (N_7502,N_5773,N_5420);
and U7503 (N_7503,N_4008,N_5952);
nor U7504 (N_7504,N_5593,N_5131);
or U7505 (N_7505,N_5849,N_5094);
and U7506 (N_7506,N_4592,N_4587);
nand U7507 (N_7507,N_5472,N_5497);
nand U7508 (N_7508,N_4551,N_5571);
nor U7509 (N_7509,N_5408,N_5018);
and U7510 (N_7510,N_5443,N_5006);
xnor U7511 (N_7511,N_4264,N_5129);
xnor U7512 (N_7512,N_5727,N_4345);
and U7513 (N_7513,N_5893,N_4562);
or U7514 (N_7514,N_5356,N_5520);
nor U7515 (N_7515,N_4363,N_4051);
and U7516 (N_7516,N_5079,N_4360);
or U7517 (N_7517,N_5357,N_5052);
xor U7518 (N_7518,N_5604,N_5994);
xor U7519 (N_7519,N_5963,N_4980);
nand U7520 (N_7520,N_4079,N_5624);
xor U7521 (N_7521,N_5807,N_5857);
nand U7522 (N_7522,N_5404,N_5547);
and U7523 (N_7523,N_4471,N_5275);
nand U7524 (N_7524,N_4681,N_4550);
nand U7525 (N_7525,N_4606,N_5942);
nand U7526 (N_7526,N_5447,N_5046);
nor U7527 (N_7527,N_4358,N_4723);
or U7528 (N_7528,N_4340,N_5841);
nor U7529 (N_7529,N_5047,N_4275);
and U7530 (N_7530,N_4075,N_4032);
nand U7531 (N_7531,N_5634,N_5946);
nand U7532 (N_7532,N_4943,N_5950);
nor U7533 (N_7533,N_4845,N_4890);
or U7534 (N_7534,N_4125,N_4409);
xnor U7535 (N_7535,N_5759,N_4337);
nand U7536 (N_7536,N_4630,N_4258);
nor U7537 (N_7537,N_4635,N_4208);
nor U7538 (N_7538,N_4435,N_5255);
nand U7539 (N_7539,N_5709,N_4642);
xor U7540 (N_7540,N_4351,N_5587);
nand U7541 (N_7541,N_5017,N_4311);
nand U7542 (N_7542,N_4773,N_5596);
nand U7543 (N_7543,N_4613,N_4791);
nor U7544 (N_7544,N_4878,N_4381);
and U7545 (N_7545,N_4262,N_5776);
nor U7546 (N_7546,N_5927,N_5394);
nor U7547 (N_7547,N_4445,N_4579);
or U7548 (N_7548,N_4325,N_4131);
nand U7549 (N_7549,N_4148,N_5321);
nand U7550 (N_7550,N_4785,N_5061);
nor U7551 (N_7551,N_5199,N_5793);
nor U7552 (N_7552,N_5254,N_5210);
and U7553 (N_7553,N_5289,N_4990);
or U7554 (N_7554,N_4390,N_5878);
nand U7555 (N_7555,N_5800,N_4853);
and U7556 (N_7556,N_4063,N_5445);
and U7557 (N_7557,N_4984,N_4007);
nand U7558 (N_7558,N_4463,N_4450);
nor U7559 (N_7559,N_5906,N_4719);
and U7560 (N_7560,N_4596,N_5214);
xor U7561 (N_7561,N_4902,N_5719);
and U7562 (N_7562,N_4025,N_4336);
or U7563 (N_7563,N_5639,N_5129);
nand U7564 (N_7564,N_5182,N_4875);
nor U7565 (N_7565,N_4031,N_4130);
and U7566 (N_7566,N_5503,N_5192);
nand U7567 (N_7567,N_4695,N_4176);
nand U7568 (N_7568,N_5666,N_5777);
nor U7569 (N_7569,N_5996,N_4454);
nand U7570 (N_7570,N_4594,N_5412);
and U7571 (N_7571,N_4554,N_5135);
xor U7572 (N_7572,N_5282,N_4873);
or U7573 (N_7573,N_4556,N_4786);
or U7574 (N_7574,N_4942,N_5891);
nor U7575 (N_7575,N_4513,N_5438);
or U7576 (N_7576,N_5247,N_4293);
or U7577 (N_7577,N_5646,N_4785);
nand U7578 (N_7578,N_4366,N_5372);
nor U7579 (N_7579,N_5089,N_4364);
nor U7580 (N_7580,N_5632,N_5097);
nand U7581 (N_7581,N_5805,N_5978);
xnor U7582 (N_7582,N_5723,N_5194);
nand U7583 (N_7583,N_4380,N_5421);
or U7584 (N_7584,N_5114,N_4242);
or U7585 (N_7585,N_4436,N_5946);
and U7586 (N_7586,N_5636,N_4710);
nor U7587 (N_7587,N_4849,N_5538);
nor U7588 (N_7588,N_5342,N_5107);
nand U7589 (N_7589,N_4048,N_5192);
or U7590 (N_7590,N_4692,N_4177);
nor U7591 (N_7591,N_4615,N_5984);
or U7592 (N_7592,N_5925,N_5254);
or U7593 (N_7593,N_5037,N_4134);
nor U7594 (N_7594,N_4116,N_5749);
or U7595 (N_7595,N_5914,N_5741);
nand U7596 (N_7596,N_4503,N_5697);
and U7597 (N_7597,N_5789,N_4434);
nor U7598 (N_7598,N_5854,N_5396);
or U7599 (N_7599,N_5760,N_4200);
and U7600 (N_7600,N_5750,N_4282);
or U7601 (N_7601,N_5419,N_4877);
nand U7602 (N_7602,N_5552,N_4743);
nand U7603 (N_7603,N_4997,N_4725);
nand U7604 (N_7604,N_4242,N_5571);
or U7605 (N_7605,N_4093,N_4112);
or U7606 (N_7606,N_4880,N_5745);
nor U7607 (N_7607,N_4535,N_4910);
or U7608 (N_7608,N_4382,N_5236);
nor U7609 (N_7609,N_4718,N_4085);
and U7610 (N_7610,N_5603,N_4713);
xor U7611 (N_7611,N_5620,N_4900);
or U7612 (N_7612,N_5455,N_4703);
nor U7613 (N_7613,N_4124,N_4739);
and U7614 (N_7614,N_5391,N_4535);
xor U7615 (N_7615,N_4730,N_4052);
or U7616 (N_7616,N_4534,N_5998);
and U7617 (N_7617,N_5587,N_4735);
and U7618 (N_7618,N_5886,N_5562);
nand U7619 (N_7619,N_4680,N_4963);
nor U7620 (N_7620,N_5483,N_5851);
or U7621 (N_7621,N_4399,N_4766);
or U7622 (N_7622,N_5625,N_5107);
nand U7623 (N_7623,N_4015,N_5241);
nor U7624 (N_7624,N_4445,N_5781);
or U7625 (N_7625,N_4572,N_4131);
nor U7626 (N_7626,N_4339,N_4188);
xor U7627 (N_7627,N_4508,N_5330);
nor U7628 (N_7628,N_5501,N_4596);
or U7629 (N_7629,N_4078,N_4578);
xnor U7630 (N_7630,N_4095,N_5412);
nand U7631 (N_7631,N_5057,N_5435);
and U7632 (N_7632,N_5926,N_4037);
nor U7633 (N_7633,N_4436,N_4752);
nor U7634 (N_7634,N_4466,N_5864);
and U7635 (N_7635,N_4892,N_4542);
or U7636 (N_7636,N_5703,N_5401);
nor U7637 (N_7637,N_5567,N_5899);
and U7638 (N_7638,N_5063,N_5771);
or U7639 (N_7639,N_4921,N_5806);
or U7640 (N_7640,N_4082,N_5502);
and U7641 (N_7641,N_4288,N_5227);
and U7642 (N_7642,N_4355,N_5906);
nor U7643 (N_7643,N_4131,N_5591);
nand U7644 (N_7644,N_4555,N_4797);
nor U7645 (N_7645,N_5493,N_4967);
nor U7646 (N_7646,N_5895,N_5204);
and U7647 (N_7647,N_5694,N_5043);
nand U7648 (N_7648,N_5608,N_4732);
nand U7649 (N_7649,N_4859,N_5046);
and U7650 (N_7650,N_5028,N_5801);
nand U7651 (N_7651,N_5449,N_4592);
nand U7652 (N_7652,N_5873,N_4383);
and U7653 (N_7653,N_5247,N_5039);
nor U7654 (N_7654,N_5301,N_4770);
nand U7655 (N_7655,N_5301,N_4061);
and U7656 (N_7656,N_5235,N_4181);
and U7657 (N_7657,N_5920,N_4815);
and U7658 (N_7658,N_4114,N_5232);
nor U7659 (N_7659,N_5549,N_4681);
nor U7660 (N_7660,N_4493,N_4050);
and U7661 (N_7661,N_5664,N_5419);
xor U7662 (N_7662,N_5777,N_4727);
nand U7663 (N_7663,N_5278,N_4049);
and U7664 (N_7664,N_4979,N_4271);
and U7665 (N_7665,N_5202,N_4287);
or U7666 (N_7666,N_5771,N_5769);
and U7667 (N_7667,N_5480,N_5428);
nand U7668 (N_7668,N_4063,N_5142);
nor U7669 (N_7669,N_4421,N_5896);
or U7670 (N_7670,N_5073,N_5487);
nor U7671 (N_7671,N_4164,N_5264);
nor U7672 (N_7672,N_4772,N_4827);
xnor U7673 (N_7673,N_5474,N_5137);
nand U7674 (N_7674,N_5169,N_5140);
or U7675 (N_7675,N_4726,N_4946);
nor U7676 (N_7676,N_5622,N_4649);
nand U7677 (N_7677,N_4659,N_4695);
or U7678 (N_7678,N_5346,N_4751);
or U7679 (N_7679,N_5937,N_5645);
and U7680 (N_7680,N_5767,N_4168);
nor U7681 (N_7681,N_4342,N_5717);
or U7682 (N_7682,N_5297,N_4187);
or U7683 (N_7683,N_5953,N_4540);
nor U7684 (N_7684,N_4458,N_5292);
nand U7685 (N_7685,N_5603,N_4491);
or U7686 (N_7686,N_5088,N_5611);
nand U7687 (N_7687,N_4401,N_4519);
nand U7688 (N_7688,N_4462,N_5612);
nor U7689 (N_7689,N_5432,N_5230);
nor U7690 (N_7690,N_4014,N_5429);
nand U7691 (N_7691,N_4918,N_4457);
nor U7692 (N_7692,N_5956,N_4392);
or U7693 (N_7693,N_4192,N_5881);
or U7694 (N_7694,N_4652,N_4741);
nand U7695 (N_7695,N_4096,N_5201);
and U7696 (N_7696,N_5648,N_5977);
nand U7697 (N_7697,N_4980,N_5193);
and U7698 (N_7698,N_5182,N_4567);
or U7699 (N_7699,N_4084,N_4759);
nand U7700 (N_7700,N_5564,N_4383);
and U7701 (N_7701,N_5952,N_5987);
and U7702 (N_7702,N_4311,N_4561);
nand U7703 (N_7703,N_4149,N_4671);
nand U7704 (N_7704,N_4271,N_5405);
or U7705 (N_7705,N_4711,N_4357);
and U7706 (N_7706,N_5497,N_5255);
nor U7707 (N_7707,N_4564,N_4653);
nand U7708 (N_7708,N_5464,N_5108);
nor U7709 (N_7709,N_4478,N_4274);
xor U7710 (N_7710,N_4624,N_4776);
nor U7711 (N_7711,N_5819,N_4810);
nand U7712 (N_7712,N_5054,N_5818);
nor U7713 (N_7713,N_4506,N_5259);
nand U7714 (N_7714,N_5801,N_5323);
or U7715 (N_7715,N_5780,N_5428);
or U7716 (N_7716,N_4176,N_4321);
nand U7717 (N_7717,N_4442,N_5863);
xnor U7718 (N_7718,N_5013,N_4603);
nand U7719 (N_7719,N_5582,N_4257);
nor U7720 (N_7720,N_5194,N_5594);
nor U7721 (N_7721,N_5381,N_4587);
nor U7722 (N_7722,N_5720,N_4079);
nor U7723 (N_7723,N_4556,N_4114);
nand U7724 (N_7724,N_5128,N_5321);
nor U7725 (N_7725,N_4955,N_5130);
nor U7726 (N_7726,N_5852,N_5766);
xor U7727 (N_7727,N_4341,N_4651);
nand U7728 (N_7728,N_4629,N_4637);
nand U7729 (N_7729,N_4226,N_5256);
or U7730 (N_7730,N_4210,N_4688);
or U7731 (N_7731,N_4414,N_5656);
xor U7732 (N_7732,N_5320,N_5353);
and U7733 (N_7733,N_4410,N_4917);
and U7734 (N_7734,N_4430,N_5865);
nand U7735 (N_7735,N_4965,N_4710);
or U7736 (N_7736,N_5986,N_4990);
and U7737 (N_7737,N_4907,N_5875);
nor U7738 (N_7738,N_4132,N_5652);
nor U7739 (N_7739,N_4029,N_4303);
nor U7740 (N_7740,N_4292,N_5758);
or U7741 (N_7741,N_5738,N_5178);
nand U7742 (N_7742,N_5089,N_4372);
and U7743 (N_7743,N_4207,N_5135);
nor U7744 (N_7744,N_5735,N_5066);
nand U7745 (N_7745,N_4600,N_5812);
and U7746 (N_7746,N_4489,N_4976);
or U7747 (N_7747,N_4645,N_5610);
nor U7748 (N_7748,N_4289,N_4368);
nor U7749 (N_7749,N_5528,N_4033);
nand U7750 (N_7750,N_5828,N_5227);
nor U7751 (N_7751,N_5834,N_4789);
and U7752 (N_7752,N_5975,N_5008);
and U7753 (N_7753,N_4533,N_4986);
and U7754 (N_7754,N_5302,N_4227);
or U7755 (N_7755,N_5307,N_5284);
nand U7756 (N_7756,N_5028,N_4270);
or U7757 (N_7757,N_4949,N_4534);
nand U7758 (N_7758,N_5133,N_4895);
nand U7759 (N_7759,N_5624,N_4921);
nor U7760 (N_7760,N_5170,N_4625);
or U7761 (N_7761,N_4605,N_4894);
or U7762 (N_7762,N_4592,N_5006);
and U7763 (N_7763,N_5606,N_4663);
nor U7764 (N_7764,N_5686,N_4992);
nand U7765 (N_7765,N_4534,N_4699);
or U7766 (N_7766,N_4769,N_5729);
or U7767 (N_7767,N_5343,N_5983);
and U7768 (N_7768,N_5525,N_4979);
nor U7769 (N_7769,N_4650,N_5456);
nand U7770 (N_7770,N_4629,N_4702);
nor U7771 (N_7771,N_4162,N_5953);
and U7772 (N_7772,N_4787,N_5508);
or U7773 (N_7773,N_4948,N_5159);
xor U7774 (N_7774,N_5945,N_5297);
nor U7775 (N_7775,N_5912,N_4346);
nor U7776 (N_7776,N_4995,N_4537);
nand U7777 (N_7777,N_4726,N_4111);
nor U7778 (N_7778,N_4695,N_5691);
and U7779 (N_7779,N_5867,N_4840);
nor U7780 (N_7780,N_5982,N_5917);
nor U7781 (N_7781,N_4006,N_5334);
nand U7782 (N_7782,N_4973,N_5150);
nand U7783 (N_7783,N_4996,N_4398);
or U7784 (N_7784,N_5372,N_4186);
nor U7785 (N_7785,N_5663,N_4751);
nor U7786 (N_7786,N_5240,N_5568);
and U7787 (N_7787,N_4081,N_5865);
nand U7788 (N_7788,N_4546,N_5237);
nor U7789 (N_7789,N_5971,N_5767);
or U7790 (N_7790,N_4202,N_5992);
nand U7791 (N_7791,N_5968,N_5017);
or U7792 (N_7792,N_4636,N_4718);
and U7793 (N_7793,N_4985,N_4219);
nand U7794 (N_7794,N_4594,N_4373);
nand U7795 (N_7795,N_5171,N_5162);
or U7796 (N_7796,N_5409,N_4421);
nand U7797 (N_7797,N_5126,N_5348);
or U7798 (N_7798,N_4345,N_5796);
nand U7799 (N_7799,N_4680,N_5786);
nor U7800 (N_7800,N_4808,N_5452);
or U7801 (N_7801,N_4109,N_5240);
or U7802 (N_7802,N_4096,N_4771);
nand U7803 (N_7803,N_4002,N_4726);
and U7804 (N_7804,N_4272,N_5637);
nand U7805 (N_7805,N_4702,N_5259);
nor U7806 (N_7806,N_4919,N_5395);
or U7807 (N_7807,N_4049,N_4893);
xor U7808 (N_7808,N_4184,N_5994);
nand U7809 (N_7809,N_5022,N_5679);
or U7810 (N_7810,N_4401,N_5029);
or U7811 (N_7811,N_5527,N_4067);
and U7812 (N_7812,N_4597,N_4738);
nor U7813 (N_7813,N_4301,N_4442);
xnor U7814 (N_7814,N_4430,N_4366);
and U7815 (N_7815,N_4290,N_5360);
or U7816 (N_7816,N_4639,N_4193);
nor U7817 (N_7817,N_5757,N_4020);
xnor U7818 (N_7818,N_4896,N_5204);
nor U7819 (N_7819,N_4881,N_4024);
or U7820 (N_7820,N_5494,N_5364);
or U7821 (N_7821,N_4021,N_4330);
and U7822 (N_7822,N_5418,N_5280);
or U7823 (N_7823,N_4238,N_4120);
or U7824 (N_7824,N_4006,N_5986);
xor U7825 (N_7825,N_4403,N_5160);
nand U7826 (N_7826,N_5919,N_5388);
xor U7827 (N_7827,N_5202,N_4640);
xor U7828 (N_7828,N_5948,N_4473);
and U7829 (N_7829,N_5033,N_4523);
or U7830 (N_7830,N_5197,N_4777);
nand U7831 (N_7831,N_5421,N_4816);
or U7832 (N_7832,N_5540,N_5126);
and U7833 (N_7833,N_5005,N_4654);
nor U7834 (N_7834,N_5215,N_4995);
or U7835 (N_7835,N_4408,N_4482);
nand U7836 (N_7836,N_5312,N_4494);
or U7837 (N_7837,N_5320,N_5139);
nor U7838 (N_7838,N_4583,N_4308);
or U7839 (N_7839,N_4042,N_5543);
or U7840 (N_7840,N_4329,N_4574);
or U7841 (N_7841,N_4765,N_5417);
or U7842 (N_7842,N_5385,N_5987);
nor U7843 (N_7843,N_5040,N_4818);
nand U7844 (N_7844,N_5915,N_5780);
or U7845 (N_7845,N_5704,N_4567);
nand U7846 (N_7846,N_4555,N_4538);
and U7847 (N_7847,N_5457,N_5783);
and U7848 (N_7848,N_5001,N_4052);
nand U7849 (N_7849,N_4418,N_4006);
and U7850 (N_7850,N_4325,N_4040);
or U7851 (N_7851,N_4301,N_4240);
nand U7852 (N_7852,N_5771,N_5872);
nand U7853 (N_7853,N_4031,N_4763);
nand U7854 (N_7854,N_4846,N_4132);
nand U7855 (N_7855,N_4840,N_4611);
and U7856 (N_7856,N_4178,N_4599);
nand U7857 (N_7857,N_4709,N_5280);
or U7858 (N_7858,N_4789,N_4846);
or U7859 (N_7859,N_4687,N_4912);
and U7860 (N_7860,N_5706,N_5019);
nor U7861 (N_7861,N_5066,N_5730);
nor U7862 (N_7862,N_4612,N_5458);
nor U7863 (N_7863,N_5297,N_5810);
and U7864 (N_7864,N_4847,N_5131);
nand U7865 (N_7865,N_5991,N_4855);
nor U7866 (N_7866,N_5777,N_4546);
nand U7867 (N_7867,N_4111,N_5007);
xor U7868 (N_7868,N_5667,N_5605);
or U7869 (N_7869,N_4723,N_4972);
and U7870 (N_7870,N_4858,N_5627);
and U7871 (N_7871,N_5350,N_5124);
nor U7872 (N_7872,N_4100,N_5513);
or U7873 (N_7873,N_5697,N_5770);
nor U7874 (N_7874,N_5380,N_5045);
nor U7875 (N_7875,N_4853,N_5942);
or U7876 (N_7876,N_4283,N_5747);
nor U7877 (N_7877,N_4923,N_4400);
and U7878 (N_7878,N_5135,N_5080);
xnor U7879 (N_7879,N_4693,N_4556);
nand U7880 (N_7880,N_5839,N_4499);
nand U7881 (N_7881,N_4571,N_4733);
nand U7882 (N_7882,N_4486,N_5230);
nor U7883 (N_7883,N_4906,N_5612);
or U7884 (N_7884,N_5291,N_5682);
and U7885 (N_7885,N_5731,N_4543);
nand U7886 (N_7886,N_4926,N_4130);
nor U7887 (N_7887,N_4822,N_4207);
nand U7888 (N_7888,N_4064,N_5845);
nor U7889 (N_7889,N_4422,N_5168);
nand U7890 (N_7890,N_4219,N_5160);
nor U7891 (N_7891,N_4259,N_5663);
xor U7892 (N_7892,N_5864,N_4737);
and U7893 (N_7893,N_4219,N_4269);
nor U7894 (N_7894,N_5737,N_5100);
nor U7895 (N_7895,N_4588,N_4190);
nor U7896 (N_7896,N_5275,N_5948);
nand U7897 (N_7897,N_5768,N_4014);
nor U7898 (N_7898,N_4634,N_4883);
and U7899 (N_7899,N_5620,N_4863);
nor U7900 (N_7900,N_4485,N_5487);
and U7901 (N_7901,N_5513,N_4976);
nor U7902 (N_7902,N_5901,N_5491);
nand U7903 (N_7903,N_4735,N_5978);
or U7904 (N_7904,N_5132,N_5629);
or U7905 (N_7905,N_5359,N_4984);
or U7906 (N_7906,N_4811,N_5576);
and U7907 (N_7907,N_4036,N_5716);
nor U7908 (N_7908,N_4826,N_4753);
nand U7909 (N_7909,N_4161,N_4321);
xor U7910 (N_7910,N_4517,N_4732);
and U7911 (N_7911,N_5155,N_4993);
or U7912 (N_7912,N_4797,N_5192);
xnor U7913 (N_7913,N_4520,N_4207);
and U7914 (N_7914,N_4347,N_5740);
and U7915 (N_7915,N_4410,N_4541);
or U7916 (N_7916,N_5218,N_4797);
xor U7917 (N_7917,N_5166,N_4344);
or U7918 (N_7918,N_4749,N_5144);
nand U7919 (N_7919,N_4480,N_4186);
and U7920 (N_7920,N_5962,N_4932);
nor U7921 (N_7921,N_5886,N_5222);
nor U7922 (N_7922,N_4749,N_4204);
xor U7923 (N_7923,N_5956,N_5815);
or U7924 (N_7924,N_4711,N_4006);
or U7925 (N_7925,N_4105,N_5120);
nand U7926 (N_7926,N_4352,N_5561);
nor U7927 (N_7927,N_4529,N_5870);
nand U7928 (N_7928,N_5327,N_4363);
or U7929 (N_7929,N_4394,N_4252);
and U7930 (N_7930,N_5005,N_5876);
and U7931 (N_7931,N_4536,N_4409);
nand U7932 (N_7932,N_5834,N_5368);
nand U7933 (N_7933,N_5690,N_5986);
nor U7934 (N_7934,N_4160,N_4132);
and U7935 (N_7935,N_4181,N_4227);
and U7936 (N_7936,N_5752,N_4573);
xor U7937 (N_7937,N_5129,N_5181);
xnor U7938 (N_7938,N_5904,N_5533);
xnor U7939 (N_7939,N_4806,N_5625);
or U7940 (N_7940,N_5268,N_4718);
nor U7941 (N_7941,N_5690,N_5083);
or U7942 (N_7942,N_4118,N_5103);
nor U7943 (N_7943,N_5757,N_4603);
or U7944 (N_7944,N_4256,N_5879);
nor U7945 (N_7945,N_5152,N_4902);
nor U7946 (N_7946,N_4436,N_4125);
nand U7947 (N_7947,N_5600,N_5915);
nand U7948 (N_7948,N_4533,N_5324);
and U7949 (N_7949,N_4933,N_5647);
nand U7950 (N_7950,N_4208,N_5947);
xor U7951 (N_7951,N_4052,N_4844);
nor U7952 (N_7952,N_4666,N_4953);
or U7953 (N_7953,N_5850,N_4212);
nor U7954 (N_7954,N_4740,N_5340);
nor U7955 (N_7955,N_4293,N_5234);
or U7956 (N_7956,N_4440,N_5229);
xor U7957 (N_7957,N_5462,N_4812);
nand U7958 (N_7958,N_4090,N_5208);
or U7959 (N_7959,N_5742,N_5042);
nor U7960 (N_7960,N_4031,N_4266);
or U7961 (N_7961,N_4668,N_4815);
nor U7962 (N_7962,N_5560,N_4746);
and U7963 (N_7963,N_5549,N_5078);
and U7964 (N_7964,N_5033,N_5223);
nor U7965 (N_7965,N_4404,N_4999);
nand U7966 (N_7966,N_5164,N_4684);
xor U7967 (N_7967,N_4743,N_4990);
and U7968 (N_7968,N_5489,N_4817);
nand U7969 (N_7969,N_4679,N_5067);
or U7970 (N_7970,N_4739,N_4177);
nor U7971 (N_7971,N_4221,N_5743);
nand U7972 (N_7972,N_5833,N_5765);
nor U7973 (N_7973,N_5400,N_4475);
nor U7974 (N_7974,N_4950,N_5322);
or U7975 (N_7975,N_5921,N_5516);
nand U7976 (N_7976,N_4427,N_4398);
nand U7977 (N_7977,N_5008,N_4248);
or U7978 (N_7978,N_5655,N_5751);
nand U7979 (N_7979,N_5221,N_5442);
nand U7980 (N_7980,N_4906,N_5089);
and U7981 (N_7981,N_4492,N_4979);
or U7982 (N_7982,N_5474,N_5682);
nand U7983 (N_7983,N_5839,N_5603);
nand U7984 (N_7984,N_4399,N_5751);
nor U7985 (N_7985,N_4074,N_4943);
nand U7986 (N_7986,N_5971,N_5993);
xnor U7987 (N_7987,N_4094,N_5278);
nor U7988 (N_7988,N_4629,N_4022);
nor U7989 (N_7989,N_4542,N_5033);
and U7990 (N_7990,N_4120,N_4184);
nor U7991 (N_7991,N_5604,N_4777);
or U7992 (N_7992,N_5678,N_5125);
nor U7993 (N_7993,N_5104,N_4737);
or U7994 (N_7994,N_4552,N_4036);
or U7995 (N_7995,N_5347,N_4475);
and U7996 (N_7996,N_4214,N_4776);
nand U7997 (N_7997,N_4049,N_5171);
nor U7998 (N_7998,N_4497,N_4066);
and U7999 (N_7999,N_5051,N_4784);
nor U8000 (N_8000,N_6392,N_6539);
nor U8001 (N_8001,N_7126,N_7944);
or U8002 (N_8002,N_7917,N_7735);
or U8003 (N_8003,N_6360,N_6968);
and U8004 (N_8004,N_6479,N_7250);
nor U8005 (N_8005,N_6111,N_6139);
nor U8006 (N_8006,N_6918,N_7394);
and U8007 (N_8007,N_6294,N_7754);
nor U8008 (N_8008,N_7681,N_6128);
and U8009 (N_8009,N_7053,N_6009);
nand U8010 (N_8010,N_7600,N_6706);
or U8011 (N_8011,N_7379,N_7176);
or U8012 (N_8012,N_7590,N_7722);
and U8013 (N_8013,N_6816,N_7210);
nand U8014 (N_8014,N_7703,N_7784);
nor U8015 (N_8015,N_7864,N_6491);
and U8016 (N_8016,N_6789,N_7622);
nor U8017 (N_8017,N_7946,N_6316);
or U8018 (N_8018,N_6750,N_6941);
or U8019 (N_8019,N_7033,N_7064);
and U8020 (N_8020,N_7093,N_6110);
and U8021 (N_8021,N_6999,N_7903);
and U8022 (N_8022,N_7090,N_6348);
or U8023 (N_8023,N_7798,N_7593);
xor U8024 (N_8024,N_6877,N_6159);
nor U8025 (N_8025,N_6279,N_7810);
xor U8026 (N_8026,N_7206,N_6793);
nor U8027 (N_8027,N_7950,N_6622);
nand U8028 (N_8028,N_7719,N_7773);
or U8029 (N_8029,N_6486,N_7478);
nor U8030 (N_8030,N_6124,N_6383);
nor U8031 (N_8031,N_6087,N_6264);
xnor U8032 (N_8032,N_7387,N_7541);
or U8033 (N_8033,N_6621,N_6880);
nand U8034 (N_8034,N_7883,N_7862);
nand U8035 (N_8035,N_7627,N_7529);
and U8036 (N_8036,N_6059,N_7100);
nand U8037 (N_8037,N_6940,N_7503);
or U8038 (N_8038,N_6105,N_6227);
xnor U8039 (N_8039,N_6770,N_6667);
and U8040 (N_8040,N_7683,N_6642);
nor U8041 (N_8041,N_6716,N_7309);
or U8042 (N_8042,N_6946,N_7231);
nand U8043 (N_8043,N_6285,N_6885);
or U8044 (N_8044,N_7433,N_7923);
nor U8045 (N_8045,N_7385,N_7113);
and U8046 (N_8046,N_7150,N_7383);
or U8047 (N_8047,N_7269,N_7599);
or U8048 (N_8048,N_6514,N_7207);
or U8049 (N_8049,N_7438,N_6334);
xnor U8050 (N_8050,N_6363,N_7553);
xor U8051 (N_8051,N_6205,N_7768);
or U8052 (N_8052,N_7425,N_7038);
or U8053 (N_8053,N_7513,N_7500);
nand U8054 (N_8054,N_6787,N_6606);
nor U8055 (N_8055,N_7248,N_6640);
or U8056 (N_8056,N_7204,N_6577);
or U8057 (N_8057,N_6496,N_7832);
nor U8058 (N_8058,N_7502,N_7157);
or U8059 (N_8059,N_6682,N_6821);
and U8060 (N_8060,N_6112,N_6434);
and U8061 (N_8061,N_7709,N_7824);
or U8062 (N_8062,N_6118,N_7302);
or U8063 (N_8063,N_7208,N_6701);
or U8064 (N_8064,N_6472,N_6088);
nand U8065 (N_8065,N_7322,N_7332);
nor U8066 (N_8066,N_7596,N_7910);
xnor U8067 (N_8067,N_6959,N_7160);
or U8068 (N_8068,N_7898,N_6417);
xor U8069 (N_8069,N_6295,N_6546);
nand U8070 (N_8070,N_6467,N_7841);
or U8071 (N_8071,N_7548,N_6030);
nor U8072 (N_8072,N_7193,N_6977);
and U8073 (N_8073,N_7264,N_6098);
nor U8074 (N_8074,N_7510,N_6278);
nand U8075 (N_8075,N_6935,N_7254);
xnor U8076 (N_8076,N_7533,N_6757);
or U8077 (N_8077,N_7785,N_7933);
and U8078 (N_8078,N_6769,N_6488);
and U8079 (N_8079,N_7908,N_7288);
and U8080 (N_8080,N_6798,N_6876);
and U8081 (N_8081,N_6765,N_7232);
nor U8082 (N_8082,N_7902,N_7829);
nor U8083 (N_8083,N_7138,N_6567);
nand U8084 (N_8084,N_7743,N_6617);
and U8085 (N_8085,N_6201,N_6568);
nand U8086 (N_8086,N_6572,N_7581);
nor U8087 (N_8087,N_7097,N_7236);
xnor U8088 (N_8088,N_7880,N_6600);
and U8089 (N_8089,N_7489,N_6355);
nand U8090 (N_8090,N_7148,N_7293);
nor U8091 (N_8091,N_7229,N_6054);
nor U8092 (N_8092,N_6969,N_6135);
or U8093 (N_8093,N_6188,N_6748);
nor U8094 (N_8094,N_6803,N_6813);
nor U8095 (N_8095,N_7962,N_7374);
nand U8096 (N_8096,N_7457,N_6317);
xnor U8097 (N_8097,N_6326,N_6053);
nand U8098 (N_8098,N_6377,N_6198);
nor U8099 (N_8099,N_6175,N_6695);
nor U8100 (N_8100,N_7051,N_7684);
and U8101 (N_8101,N_6847,N_7114);
nand U8102 (N_8102,N_6874,N_6441);
and U8103 (N_8103,N_6257,N_7826);
nor U8104 (N_8104,N_6008,N_6504);
or U8105 (N_8105,N_6978,N_6191);
nand U8106 (N_8106,N_6819,N_6527);
and U8107 (N_8107,N_7927,N_6433);
nor U8108 (N_8108,N_6767,N_7808);
nand U8109 (N_8109,N_6996,N_6010);
xor U8110 (N_8110,N_7740,N_6861);
nor U8111 (N_8111,N_7220,N_7080);
and U8112 (N_8112,N_7105,N_6826);
nand U8113 (N_8113,N_7642,N_7377);
nand U8114 (N_8114,N_6419,N_7279);
xor U8115 (N_8115,N_7274,N_6266);
and U8116 (N_8116,N_6713,N_7532);
nand U8117 (N_8117,N_7873,N_7641);
and U8118 (N_8118,N_7865,N_7825);
or U8119 (N_8119,N_6648,N_6856);
xor U8120 (N_8120,N_6933,N_6230);
nand U8121 (N_8121,N_7414,N_7716);
nand U8122 (N_8122,N_7820,N_7911);
nand U8123 (N_8123,N_7386,N_7778);
nand U8124 (N_8124,N_6313,N_7122);
or U8125 (N_8125,N_7144,N_7119);
nor U8126 (N_8126,N_7672,N_7665);
nor U8127 (N_8127,N_7084,N_6058);
or U8128 (N_8128,N_7981,N_6980);
nor U8129 (N_8129,N_7762,N_6899);
nor U8130 (N_8130,N_6492,N_7140);
nand U8131 (N_8131,N_7247,N_7977);
nor U8132 (N_8132,N_6604,N_7850);
nor U8133 (N_8133,N_7517,N_6148);
and U8134 (N_8134,N_6714,N_7339);
or U8135 (N_8135,N_7615,N_6570);
nor U8136 (N_8136,N_7101,N_7760);
and U8137 (N_8137,N_7595,N_7586);
nand U8138 (N_8138,N_6023,N_7852);
or U8139 (N_8139,N_7062,N_7580);
or U8140 (N_8140,N_7439,N_6231);
or U8141 (N_8141,N_6049,N_7547);
or U8142 (N_8142,N_7861,N_7895);
nand U8143 (N_8143,N_7368,N_6563);
nand U8144 (N_8144,N_6209,N_6315);
and U8145 (N_8145,N_6428,N_7594);
nor U8146 (N_8146,N_7494,N_7575);
nor U8147 (N_8147,N_7801,N_7071);
and U8148 (N_8148,N_7991,N_6084);
xor U8149 (N_8149,N_6134,N_6628);
nor U8150 (N_8150,N_6415,N_7397);
nor U8151 (N_8151,N_7648,N_7240);
and U8152 (N_8152,N_7365,N_6920);
nand U8153 (N_8153,N_6371,N_6222);
nand U8154 (N_8154,N_7835,N_7437);
or U8155 (N_8155,N_7116,N_7751);
nor U8156 (N_8156,N_6709,N_6693);
nand U8157 (N_8157,N_6542,N_6443);
xor U8158 (N_8158,N_7772,N_7069);
or U8159 (N_8159,N_6760,N_6669);
and U8160 (N_8160,N_7526,N_6519);
nor U8161 (N_8161,N_7999,N_7249);
nor U8162 (N_8162,N_7166,N_6208);
and U8163 (N_8163,N_7729,N_7226);
or U8164 (N_8164,N_6248,N_7068);
or U8165 (N_8165,N_6296,N_6361);
xnor U8166 (N_8166,N_6729,N_6814);
xor U8167 (N_8167,N_7261,N_6849);
and U8168 (N_8168,N_6988,N_7731);
xor U8169 (N_8169,N_7442,N_7525);
nor U8170 (N_8170,N_7583,N_6677);
nand U8171 (N_8171,N_6138,N_6862);
nor U8172 (N_8172,N_7516,N_6903);
xor U8173 (N_8173,N_7660,N_7435);
nor U8174 (N_8174,N_7662,N_7454);
nand U8175 (N_8175,N_6218,N_7271);
nor U8176 (N_8176,N_6463,N_6283);
and U8177 (N_8177,N_7564,N_6154);
nand U8178 (N_8178,N_7334,N_6223);
and U8179 (N_8179,N_6853,N_7812);
nor U8180 (N_8180,N_6307,N_7076);
or U8181 (N_8181,N_6657,N_6906);
nor U8182 (N_8182,N_6619,N_7597);
or U8183 (N_8183,N_7380,N_7953);
or U8184 (N_8184,N_6618,N_6919);
nand U8185 (N_8185,N_7949,N_6390);
nand U8186 (N_8186,N_7049,N_6025);
nor U8187 (N_8187,N_6498,N_7321);
xor U8188 (N_8188,N_7406,N_6336);
and U8189 (N_8189,N_6343,N_7155);
nor U8190 (N_8190,N_6516,N_7693);
xor U8191 (N_8191,N_7283,N_7089);
nor U8192 (N_8192,N_6964,N_6153);
or U8193 (N_8193,N_6974,N_6900);
and U8194 (N_8194,N_7921,N_7942);
or U8195 (N_8195,N_6495,N_6471);
nand U8196 (N_8196,N_7601,N_7881);
and U8197 (N_8197,N_7614,N_7424);
nor U8198 (N_8198,N_6952,N_7882);
nor U8199 (N_8199,N_7120,N_6277);
xnor U8200 (N_8200,N_6818,N_6983);
or U8201 (N_8201,N_7694,N_7359);
or U8202 (N_8202,N_6528,N_7373);
nand U8203 (N_8203,N_7189,N_6002);
and U8204 (N_8204,N_7016,N_6200);
nor U8205 (N_8205,N_7043,N_7968);
and U8206 (N_8206,N_7849,N_6794);
nor U8207 (N_8207,N_6839,N_7984);
and U8208 (N_8208,N_7461,N_6039);
and U8209 (N_8209,N_6995,N_6302);
nor U8210 (N_8210,N_6834,N_6353);
nor U8211 (N_8211,N_6487,N_6776);
nor U8212 (N_8212,N_6203,N_7054);
nand U8213 (N_8213,N_6561,N_6210);
nand U8214 (N_8214,N_6782,N_7721);
or U8215 (N_8215,N_7156,N_7019);
nand U8216 (N_8216,N_7806,N_7096);
nand U8217 (N_8217,N_7603,N_6368);
and U8218 (N_8218,N_6115,N_6873);
nor U8219 (N_8219,N_7388,N_7788);
and U8220 (N_8220,N_7670,N_7727);
nor U8221 (N_8221,N_7707,N_6425);
xor U8222 (N_8222,N_6629,N_6631);
or U8223 (N_8223,N_7434,N_7970);
xnor U8224 (N_8224,N_6590,N_6450);
and U8225 (N_8225,N_6824,N_6897);
or U8226 (N_8226,N_6038,N_7331);
or U8227 (N_8227,N_7185,N_6435);
and U8228 (N_8228,N_7109,N_7636);
or U8229 (N_8229,N_7451,N_6364);
and U8230 (N_8230,N_7795,N_6309);
or U8231 (N_8231,N_6186,N_7780);
and U8232 (N_8232,N_6375,N_6571);
xnor U8233 (N_8233,N_6679,N_6917);
nor U8234 (N_8234,N_6276,N_6505);
nand U8235 (N_8235,N_7867,N_7147);
xnor U8236 (N_8236,N_6944,N_6595);
or U8237 (N_8237,N_6830,N_7530);
xor U8238 (N_8238,N_7871,N_7598);
nor U8239 (N_8239,N_6842,N_7037);
nor U8240 (N_8240,N_7201,N_6724);
and U8241 (N_8241,N_6651,N_6122);
xor U8242 (N_8242,N_6177,N_7017);
nand U8243 (N_8243,N_7680,N_7239);
nand U8244 (N_8244,N_7630,N_6125);
and U8245 (N_8245,N_7854,N_6020);
or U8246 (N_8246,N_6668,N_6199);
nor U8247 (N_8247,N_6187,N_7106);
or U8248 (N_8248,N_7668,N_6520);
nand U8249 (N_8249,N_7194,N_7794);
nand U8250 (N_8250,N_6120,N_6290);
or U8251 (N_8251,N_7335,N_7092);
nor U8252 (N_8252,N_6905,N_7947);
or U8253 (N_8253,N_6108,N_7487);
or U8254 (N_8254,N_6181,N_6270);
or U8255 (N_8255,N_6462,N_6066);
nor U8256 (N_8256,N_6986,N_7562);
or U8257 (N_8257,N_6144,N_7198);
xor U8258 (N_8258,N_7926,N_6344);
nor U8259 (N_8259,N_6378,N_7610);
nand U8260 (N_8260,N_7847,N_6609);
nor U8261 (N_8261,N_6687,N_7472);
nor U8262 (N_8262,N_6014,N_6453);
or U8263 (N_8263,N_6737,N_7455);
nor U8264 (N_8264,N_7845,N_6725);
nor U8265 (N_8265,N_6635,N_7522);
xor U8266 (N_8266,N_7316,N_6410);
and U8267 (N_8267,N_6678,N_7759);
and U8268 (N_8268,N_7221,N_6146);
and U8269 (N_8269,N_7624,N_6989);
and U8270 (N_8270,N_7542,N_7291);
nand U8271 (N_8271,N_6070,N_7496);
nor U8272 (N_8272,N_7919,N_7811);
or U8273 (N_8273,N_7696,N_7104);
xor U8274 (N_8274,N_6586,N_7215);
nand U8275 (N_8275,N_6216,N_7689);
or U8276 (N_8276,N_6961,N_7958);
or U8277 (N_8277,N_6473,N_6838);
nand U8278 (N_8278,N_7401,N_6573);
or U8279 (N_8279,N_7131,N_7134);
or U8280 (N_8280,N_6926,N_6015);
xnor U8281 (N_8281,N_7336,N_6632);
nor U8282 (N_8282,N_6747,N_6259);
or U8283 (N_8283,N_6575,N_7987);
or U8284 (N_8284,N_7676,N_7527);
nor U8285 (N_8285,N_7251,N_7172);
or U8286 (N_8286,N_7813,N_6396);
xnor U8287 (N_8287,N_6262,N_6207);
nor U8288 (N_8288,N_7605,N_7706);
and U8289 (N_8289,N_6720,N_6869);
or U8290 (N_8290,N_7479,N_6164);
nor U8291 (N_8291,N_7165,N_6676);
nor U8292 (N_8292,N_7197,N_6300);
or U8293 (N_8293,N_7356,N_6409);
and U8294 (N_8294,N_7007,N_6686);
nor U8295 (N_8295,N_7905,N_7514);
and U8296 (N_8296,N_7063,N_7338);
nand U8297 (N_8297,N_7545,N_7179);
and U8298 (N_8298,N_6778,N_7749);
nand U8299 (N_8299,N_7326,N_6150);
nand U8300 (N_8300,N_7475,N_6273);
and U8301 (N_8301,N_7884,N_7354);
or U8302 (N_8302,N_7554,N_6101);
or U8303 (N_8303,N_7364,N_7417);
and U8304 (N_8304,N_6734,N_7819);
and U8305 (N_8305,N_7075,N_6469);
xor U8306 (N_8306,N_7470,N_6131);
nand U8307 (N_8307,N_7918,N_6820);
nor U8308 (N_8308,N_6158,N_6797);
and U8309 (N_8309,N_6314,N_6466);
nand U8310 (N_8310,N_6909,N_7427);
and U8311 (N_8311,N_6685,N_6616);
and U8312 (N_8312,N_7961,N_6046);
and U8313 (N_8313,N_6581,N_7682);
xnor U8314 (N_8314,N_6055,N_7543);
or U8315 (N_8315,N_6241,N_6972);
nor U8316 (N_8316,N_6945,N_6949);
nor U8317 (N_8317,N_7285,N_7912);
nor U8318 (N_8318,N_6553,N_6804);
nand U8319 (N_8319,N_6416,N_7718);
and U8320 (N_8320,N_6837,N_7638);
xnor U8321 (N_8321,N_7764,N_7663);
or U8322 (N_8322,N_7159,N_6551);
or U8323 (N_8323,N_6708,N_6866);
and U8324 (N_8324,N_6073,N_6096);
xor U8325 (N_8325,N_7123,N_7639);
and U8326 (N_8326,N_6051,N_7842);
nor U8327 (N_8327,N_7536,N_6966);
and U8328 (N_8328,N_6123,N_6831);
nand U8329 (N_8329,N_7004,N_7300);
xnor U8330 (N_8330,N_6224,N_7875);
nor U8331 (N_8331,N_7544,N_6939);
or U8332 (N_8332,N_6076,N_6658);
nand U8333 (N_8333,N_7431,N_6427);
xor U8334 (N_8334,N_7402,N_6413);
nor U8335 (N_8335,N_7914,N_6745);
nand U8336 (N_8336,N_7631,N_7456);
nor U8337 (N_8337,N_7700,N_7647);
and U8338 (N_8338,N_6746,N_6502);
nand U8339 (N_8339,N_7164,N_7118);
and U8340 (N_8340,N_7899,N_6061);
nor U8341 (N_8341,N_6732,N_7015);
and U8342 (N_8342,N_7182,N_6936);
nor U8343 (N_8343,N_6050,N_6764);
nor U8344 (N_8344,N_6072,N_7606);
and U8345 (N_8345,N_6160,N_6660);
or U8346 (N_8346,N_7952,N_7688);
nand U8347 (N_8347,N_6783,N_6735);
nor U8348 (N_8348,N_7750,N_6958);
xor U8349 (N_8349,N_7256,N_7972);
or U8350 (N_8350,N_6499,N_6650);
and U8351 (N_8351,N_7242,N_6956);
and U8352 (N_8352,N_6907,N_7998);
or U8353 (N_8353,N_6557,N_7143);
nor U8354 (N_8354,N_7993,N_6942);
nor U8355 (N_8355,N_6221,N_6174);
or U8356 (N_8356,N_7538,N_6000);
nor U8357 (N_8357,N_6078,N_6235);
and U8358 (N_8358,N_6372,N_6407);
nand U8359 (N_8359,N_6109,N_6625);
or U8360 (N_8360,N_6265,N_7828);
or U8361 (N_8361,N_6069,N_6319);
nor U8362 (N_8362,N_7747,N_6696);
nor U8363 (N_8363,N_7827,N_6915);
nor U8364 (N_8364,N_7938,N_7715);
and U8365 (N_8365,N_6854,N_7151);
and U8366 (N_8366,N_7860,N_6068);
nor U8367 (N_8367,N_7506,N_6119);
nor U8368 (N_8368,N_7124,N_6057);
nand U8369 (N_8369,N_7405,N_6664);
or U8370 (N_8370,N_6460,N_6261);
nand U8371 (N_8371,N_6132,N_6848);
and U8372 (N_8372,N_6156,N_6365);
nor U8373 (N_8373,N_6385,N_7956);
or U8374 (N_8374,N_7640,N_7807);
nor U8375 (N_8375,N_6711,N_6176);
nor U8376 (N_8376,N_7960,N_6075);
or U8377 (N_8377,N_6288,N_7787);
or U8378 (N_8378,N_7419,N_6850);
and U8379 (N_8379,N_7745,N_6973);
nor U8380 (N_8380,N_6100,N_6281);
or U8381 (N_8381,N_6954,N_7102);
nand U8382 (N_8382,N_6229,N_6476);
or U8383 (N_8383,N_7979,N_6256);
nand U8384 (N_8384,N_7734,N_7499);
xor U8385 (N_8385,N_6149,N_6406);
or U8386 (N_8386,N_7704,N_7202);
or U8387 (N_8387,N_6872,N_6442);
nor U8388 (N_8388,N_6569,N_7728);
nand U8389 (N_8389,N_6901,N_6099);
nor U8390 (N_8390,N_6690,N_7428);
or U8391 (N_8391,N_7973,N_6599);
and U8392 (N_8392,N_6093,N_7649);
and U8393 (N_8393,N_7268,N_6373);
nand U8394 (N_8394,N_6532,N_6217);
and U8395 (N_8395,N_6515,N_6157);
and U8396 (N_8396,N_6928,N_6330);
and U8397 (N_8397,N_6673,N_6358);
nand U8398 (N_8398,N_6772,N_6638);
nand U8399 (N_8399,N_7679,N_7465);
or U8400 (N_8400,N_6267,N_7001);
and U8401 (N_8401,N_7619,N_6432);
nand U8402 (N_8402,N_7928,N_7410);
nor U8403 (N_8403,N_7579,N_7915);
or U8404 (N_8404,N_7152,N_6970);
and U8405 (N_8405,N_6292,N_7589);
nand U8406 (N_8406,N_7626,N_6067);
or U8407 (N_8407,N_6147,N_6547);
nand U8408 (N_8408,N_6888,N_6006);
or U8409 (N_8409,N_6998,N_7730);
nor U8410 (N_8410,N_6212,N_7078);
nand U8411 (N_8411,N_7447,N_7180);
nand U8412 (N_8412,N_7550,N_6666);
and U8413 (N_8413,N_7121,N_6846);
or U8414 (N_8414,N_6401,N_6802);
or U8415 (N_8415,N_6366,N_6751);
and U8416 (N_8416,N_7369,N_6140);
or U8417 (N_8417,N_6369,N_7146);
nand U8418 (N_8418,N_7280,N_6795);
nand U8419 (N_8419,N_6624,N_6323);
xnor U8420 (N_8420,N_7505,N_6483);
and U8421 (N_8421,N_6518,N_7382);
nand U8422 (N_8422,N_6967,N_6027);
nor U8423 (N_8423,N_7711,N_6077);
or U8424 (N_8424,N_6962,N_6056);
and U8425 (N_8425,N_7058,N_6041);
nor U8426 (N_8426,N_6328,N_7045);
and U8427 (N_8427,N_6242,N_7440);
nand U8428 (N_8428,N_6680,N_6493);
nor U8429 (N_8429,N_6934,N_6446);
nand U8430 (N_8430,N_6032,N_6605);
nand U8431 (N_8431,N_7132,N_7244);
or U8432 (N_8432,N_6858,N_6731);
nand U8433 (N_8433,N_7777,N_7994);
nor U8434 (N_8434,N_7178,N_7345);
nand U8435 (N_8435,N_7192,N_7423);
nor U8436 (N_8436,N_6937,N_7030);
and U8437 (N_8437,N_6785,N_6249);
nand U8438 (N_8438,N_7072,N_6351);
nor U8439 (N_8439,N_7422,N_6700);
nand U8440 (N_8440,N_7552,N_7349);
xor U8441 (N_8441,N_6643,N_7384);
and U8442 (N_8442,N_6219,N_6255);
and U8443 (N_8443,N_7814,N_7327);
nor U8444 (N_8444,N_6214,N_7234);
nor U8445 (N_8445,N_6386,N_7341);
and U8446 (N_8446,N_6012,N_6889);
and U8447 (N_8447,N_6552,N_7558);
or U8448 (N_8448,N_7262,N_7314);
and U8449 (N_8449,N_6984,N_7129);
nor U8450 (N_8450,N_7634,N_7817);
and U8451 (N_8451,N_6404,N_7556);
nor U8452 (N_8452,N_7246,N_6397);
nand U8453 (N_8453,N_6507,N_6444);
nand U8454 (N_8454,N_7686,N_7281);
or U8455 (N_8455,N_6091,N_6882);
and U8456 (N_8456,N_6718,N_7378);
and U8457 (N_8457,N_7413,N_7361);
nand U8458 (N_8458,N_6354,N_7395);
and U8459 (N_8459,N_7398,N_6822);
nor U8460 (N_8460,N_6168,N_7848);
or U8461 (N_8461,N_7989,N_7362);
nor U8462 (N_8462,N_7443,N_6306);
nand U8463 (N_8463,N_7408,N_6766);
nor U8464 (N_8464,N_7592,N_7888);
nor U8465 (N_8465,N_6662,N_7643);
and U8466 (N_8466,N_6195,N_7325);
xnor U8467 (N_8467,N_7879,N_7504);
nand U8468 (N_8468,N_6349,N_6759);
nor U8469 (N_8469,N_7651,N_6083);
nand U8470 (N_8470,N_6545,N_6761);
xnor U8471 (N_8471,N_6297,N_6852);
nor U8472 (N_8472,N_7652,N_7486);
and U8473 (N_8473,N_6948,N_6913);
and U8474 (N_8474,N_6284,N_7843);
or U8475 (N_8475,N_6896,N_6870);
nor U8476 (N_8476,N_6584,N_7013);
and U8477 (N_8477,N_7604,N_6688);
and U8478 (N_8478,N_6788,N_7350);
nor U8479 (N_8479,N_7789,N_7393);
nor U8480 (N_8480,N_7186,N_7870);
or U8481 (N_8481,N_7255,N_7717);
nor U8482 (N_8482,N_6163,N_6689);
nor U8483 (N_8483,N_7420,N_7524);
xnor U8484 (N_8484,N_7351,N_6021);
nor U8485 (N_8485,N_6258,N_7358);
nor U8486 (N_8486,N_7492,N_7048);
and U8487 (N_8487,N_6155,N_7429);
nor U8488 (N_8488,N_7781,N_6454);
or U8489 (N_8489,N_7432,N_7468);
or U8490 (N_8490,N_6898,N_7623);
nand U8491 (N_8491,N_7082,N_6799);
nor U8492 (N_8492,N_6141,N_7797);
or U8493 (N_8493,N_6654,N_7803);
or U8494 (N_8494,N_6845,N_6352);
or U8495 (N_8495,N_7954,N_7169);
nor U8496 (N_8496,N_7416,N_6494);
nor U8497 (N_8497,N_6768,N_6840);
xor U8498 (N_8498,N_7658,N_7653);
and U8499 (N_8499,N_7230,N_7591);
or U8500 (N_8500,N_6681,N_7705);
nor U8501 (N_8501,N_7576,N_7095);
xnor U8502 (N_8502,N_6509,N_7687);
nand U8503 (N_8503,N_6884,N_6698);
nor U8504 (N_8504,N_6929,N_6742);
nand U8505 (N_8505,N_7951,N_7929);
or U8506 (N_8506,N_7907,N_6220);
nor U8507 (N_8507,N_7853,N_7024);
or U8508 (N_8508,N_7809,N_6975);
nor U8509 (N_8509,N_7574,N_6634);
or U8510 (N_8510,N_7985,N_6851);
or U8511 (N_8511,N_6080,N_6304);
or U8512 (N_8512,N_6753,N_7876);
and U8513 (N_8513,N_6185,N_7329);
and U8514 (N_8514,N_6085,N_6311);
nor U8515 (N_8515,N_7746,N_6786);
or U8516 (N_8516,N_6591,N_7243);
nor U8517 (N_8517,N_6206,N_6033);
nor U8518 (N_8518,N_6036,N_7463);
xnor U8519 (N_8519,N_7008,N_6367);
and U8520 (N_8520,N_7702,N_6921);
and U8521 (N_8521,N_6844,N_7391);
nor U8522 (N_8522,N_6335,N_6721);
and U8523 (N_8523,N_7877,N_7618);
nor U8524 (N_8524,N_7199,N_7233);
nor U8525 (N_8525,N_6356,N_7436);
nor U8526 (N_8526,N_7978,N_7153);
nand U8527 (N_8527,N_6342,N_6792);
and U8528 (N_8528,N_7802,N_6357);
nand U8529 (N_8529,N_7671,N_6774);
or U8530 (N_8530,N_7171,N_6864);
nor U8531 (N_8531,N_6574,N_7485);
xor U8532 (N_8532,N_6272,N_6282);
or U8533 (N_8533,N_7892,N_7307);
nand U8534 (N_8534,N_6011,N_7967);
nor U8535 (N_8535,N_7257,N_7367);
nand U8536 (N_8536,N_6173,N_6533);
nor U8537 (N_8537,N_6310,N_7273);
xnor U8538 (N_8538,N_6712,N_6097);
and U8539 (N_8539,N_7790,N_7983);
nor U8540 (N_8540,N_6506,N_7612);
nor U8541 (N_8541,N_6028,N_7909);
and U8542 (N_8542,N_7036,N_7141);
nand U8543 (N_8543,N_7766,N_6512);
and U8544 (N_8544,N_6347,N_7112);
xnor U8545 (N_8545,N_6184,N_6090);
and U8546 (N_8546,N_7521,N_6904);
and U8547 (N_8547,N_7557,N_6585);
or U8548 (N_8548,N_6930,N_6420);
or U8549 (N_8549,N_6082,N_7736);
nor U8550 (N_8550,N_6308,N_7018);
nand U8551 (N_8551,N_7403,N_6979);
nor U8552 (N_8552,N_7617,N_6536);
nand U8553 (N_8553,N_6727,N_6481);
and U8554 (N_8554,N_7409,N_6908);
or U8555 (N_8555,N_6893,N_6612);
nand U8556 (N_8556,N_7426,N_7218);
nor U8557 (N_8557,N_7969,N_6412);
nor U8558 (N_8558,N_7389,N_7995);
nor U8559 (N_8559,N_7237,N_6683);
or U8560 (N_8560,N_7632,N_7173);
and U8561 (N_8561,N_7177,N_7306);
and U8562 (N_8562,N_6489,N_6268);
xor U8563 (N_8563,N_6811,N_6801);
or U8564 (N_8564,N_6548,N_6398);
xnor U8565 (N_8565,N_7059,N_6391);
or U8566 (N_8566,N_7913,N_7560);
xnor U8567 (N_8567,N_7056,N_7073);
and U8568 (N_8568,N_6923,N_7799);
nor U8569 (N_8569,N_7110,N_7471);
nand U8570 (N_8570,N_7966,N_7497);
and U8571 (N_8571,N_7028,N_6950);
and U8572 (N_8572,N_7901,N_7484);
or U8573 (N_8573,N_7066,N_7039);
xor U8574 (N_8574,N_6559,N_7948);
nor U8575 (N_8575,N_6301,N_7906);
or U8576 (N_8576,N_7343,N_6841);
and U8577 (N_8577,N_6117,N_6594);
and U8578 (N_8578,N_6287,N_7539);
and U8579 (N_8579,N_6740,N_7014);
or U8580 (N_8580,N_7200,N_7650);
nor U8581 (N_8581,N_7733,N_6603);
nor U8582 (N_8582,N_6423,N_6556);
nand U8583 (N_8583,N_6228,N_7352);
xnor U8584 (N_8584,N_6843,N_6914);
xnor U8585 (N_8585,N_7613,N_6202);
and U8586 (N_8586,N_7381,N_7213);
nand U8587 (N_8587,N_6250,N_7992);
or U8588 (N_8588,N_6647,N_7286);
nor U8589 (N_8589,N_7127,N_7277);
and U8590 (N_8590,N_7887,N_6102);
xnor U8591 (N_8591,N_7145,N_6247);
nand U8592 (N_8592,N_6812,N_6508);
nor U8593 (N_8593,N_7212,N_7863);
nor U8594 (N_8594,N_7258,N_6503);
nor U8595 (N_8595,N_6943,N_6922);
nor U8596 (N_8596,N_6395,N_7304);
and U8597 (N_8597,N_6321,N_6437);
nand U8598 (N_8598,N_7372,N_6522);
or U8599 (N_8599,N_7363,N_7139);
or U8600 (N_8600,N_6796,N_6022);
nand U8601 (N_8601,N_6531,N_7289);
xor U8602 (N_8602,N_7411,N_7055);
nand U8603 (N_8603,N_7509,N_6478);
or U8604 (N_8604,N_7566,N_6318);
nor U8605 (N_8605,N_6464,N_7869);
nand U8606 (N_8606,N_6815,N_7568);
or U8607 (N_8607,N_6388,N_6810);
or U8608 (N_8608,N_6005,N_6762);
nor U8609 (N_8609,N_6382,N_7125);
and U8610 (N_8610,N_7263,N_7834);
and U8611 (N_8611,N_7572,N_6601);
nor U8612 (N_8612,N_7238,N_6016);
or U8613 (N_8613,N_7724,N_6065);
nand U8614 (N_8614,N_6114,N_7737);
and U8615 (N_8615,N_7965,N_7301);
and U8616 (N_8616,N_6251,N_7868);
and U8617 (N_8617,N_6705,N_6894);
or U8618 (N_8618,N_6863,N_7900);
xnor U8619 (N_8619,N_7752,N_7184);
nor U8620 (N_8620,N_7836,N_6475);
nand U8621 (N_8621,N_6172,N_7009);
or U8622 (N_8622,N_7458,N_6074);
nand U8623 (N_8623,N_6610,N_7673);
or U8624 (N_8624,N_6955,N_6233);
and U8625 (N_8625,N_6675,N_7886);
and U8626 (N_8626,N_6225,N_6299);
nand U8627 (N_8627,N_6338,N_6910);
nor U8628 (N_8628,N_7855,N_6932);
xor U8629 (N_8629,N_7183,N_6468);
nand U8630 (N_8630,N_7635,N_7941);
nand U8631 (N_8631,N_6773,N_7459);
nor U8632 (N_8632,N_7034,N_7551);
and U8633 (N_8633,N_7563,N_6890);
nor U8634 (N_8634,N_7011,N_7602);
nor U8635 (N_8635,N_6560,N_6452);
nand U8636 (N_8636,N_7939,N_7081);
xnor U8637 (N_8637,N_7299,N_6013);
and U8638 (N_8638,N_7245,N_7783);
or U8639 (N_8639,N_6775,N_6674);
nand U8640 (N_8640,N_7006,N_6260);
nand U8641 (N_8641,N_6239,N_7761);
xor U8642 (N_8642,N_7937,N_7555);
nor U8643 (N_8643,N_6136,N_6589);
nor U8644 (N_8644,N_6938,N_6129);
or U8645 (N_8645,N_6438,N_7655);
nor U8646 (N_8646,N_6611,N_7010);
and U8647 (N_8647,N_6672,N_6550);
nand U8648 (N_8648,N_7698,N_7837);
nand U8649 (N_8649,N_6094,N_6728);
or U8650 (N_8650,N_6510,N_7695);
and U8651 (N_8651,N_7047,N_7086);
or U8652 (N_8652,N_7523,N_6440);
nand U8653 (N_8653,N_7430,N_6370);
or U8654 (N_8654,N_7758,N_7117);
and U8655 (N_8655,N_6133,N_7934);
or U8656 (N_8656,N_7453,N_7270);
nand U8657 (N_8657,N_6555,N_6293);
nor U8658 (N_8658,N_6582,N_7091);
and U8659 (N_8659,N_7128,N_7833);
and U8660 (N_8660,N_7450,N_7357);
and U8661 (N_8661,N_7214,N_7578);
or U8662 (N_8662,N_6661,N_7346);
or U8663 (N_8663,N_7866,N_6381);
nor U8664 (N_8664,N_6517,N_6809);
or U8665 (N_8665,N_7666,N_7130);
and U8666 (N_8666,N_7742,N_6271);
and U8667 (N_8667,N_7098,N_7032);
and U8668 (N_8668,N_7046,N_7587);
or U8669 (N_8669,N_6474,N_6245);
nand U8670 (N_8670,N_7629,N_6627);
xnor U8671 (N_8671,N_7415,N_6722);
and U8672 (N_8672,N_7107,N_7646);
nand U8673 (N_8673,N_7846,N_7508);
nand U8674 (N_8674,N_7637,N_6780);
nor U8675 (N_8675,N_7481,N_7044);
nor U8676 (N_8676,N_6730,N_7816);
nand U8677 (N_8677,N_6095,N_6543);
nor U8678 (N_8678,N_6137,N_6596);
nand U8679 (N_8679,N_7347,N_6060);
nor U8680 (N_8680,N_7943,N_6092);
and U8681 (N_8681,N_7170,N_7559);
or U8682 (N_8682,N_6192,N_6566);
or U8683 (N_8683,N_7611,N_7297);
nand U8684 (N_8684,N_7412,N_6341);
or U8685 (N_8685,N_7725,N_6564);
and U8686 (N_8686,N_6380,N_7515);
nor U8687 (N_8687,N_7421,N_7317);
or U8688 (N_8688,N_7272,N_6992);
nor U8689 (N_8689,N_6048,N_6213);
or U8690 (N_8690,N_7924,N_7616);
or U8691 (N_8691,N_6916,N_6052);
and U8692 (N_8692,N_7290,N_6710);
nor U8693 (N_8693,N_7087,N_6332);
or U8694 (N_8694,N_6501,N_6652);
or U8695 (N_8695,N_7588,N_6197);
nand U8696 (N_8696,N_6480,N_6883);
nor U8697 (N_8697,N_7195,N_6524);
nand U8698 (N_8698,N_6399,N_6449);
and U8699 (N_8699,N_6145,N_7319);
xor U8700 (N_8700,N_7577,N_6405);
nor U8701 (N_8701,N_7035,N_7821);
nand U8702 (N_8702,N_7040,N_6715);
or U8703 (N_8703,N_7320,N_6171);
nand U8704 (N_8704,N_6763,N_7894);
nand U8705 (N_8705,N_6749,N_7181);
nor U8706 (N_8706,N_6004,N_6829);
nor U8707 (N_8707,N_6752,N_6549);
nor U8708 (N_8708,N_6645,N_6040);
and U8709 (N_8709,N_6670,N_6867);
or U8710 (N_8710,N_7042,N_7466);
or U8711 (N_8711,N_7266,N_6431);
and U8712 (N_8712,N_7252,N_6162);
nor U8713 (N_8713,N_7830,N_7022);
nand U8714 (N_8714,N_7392,N_6511);
nand U8715 (N_8715,N_7756,N_6726);
nand U8716 (N_8716,N_7769,N_7371);
nand U8717 (N_8717,N_7224,N_7099);
or U8718 (N_8718,N_6630,N_6738);
nand U8719 (N_8719,N_6691,N_7491);
nor U8720 (N_8720,N_6871,N_7858);
nand U8721 (N_8721,N_6895,N_6345);
xor U8722 (N_8722,N_7697,N_6779);
and U8723 (N_8723,N_6562,N_7278);
and U8724 (N_8724,N_7460,N_6723);
nor U8725 (N_8725,N_7088,N_6121);
nand U8726 (N_8726,N_7296,N_7971);
xor U8727 (N_8727,N_6653,N_6823);
nand U8728 (N_8728,N_6754,N_6183);
nand U8729 (N_8729,N_6957,N_6459);
or U8730 (N_8730,N_7691,N_7963);
nand U8731 (N_8731,N_6692,N_7065);
and U8732 (N_8732,N_7738,N_6736);
or U8733 (N_8733,N_7253,N_7805);
nand U8734 (N_8734,N_7337,N_6400);
nor U8735 (N_8735,N_7904,N_7366);
xnor U8736 (N_8736,N_6997,N_6455);
nand U8737 (N_8737,N_6523,N_7930);
nand U8738 (N_8738,N_6659,N_6246);
nand U8739 (N_8739,N_6485,N_7077);
nand U8740 (N_8740,N_6113,N_7844);
nand U8741 (N_8741,N_7360,N_6043);
or U8742 (N_8742,N_7657,N_6018);
nor U8743 (N_8743,N_7057,N_6833);
nor U8744 (N_8744,N_7669,N_7467);
and U8745 (N_8745,N_7473,N_6331);
nand U8746 (N_8746,N_6402,N_6269);
nor U8747 (N_8747,N_6513,N_6598);
or U8748 (N_8748,N_6447,N_6490);
and U8749 (N_8749,N_6580,N_6758);
or U8750 (N_8750,N_7324,N_7893);
xnor U8751 (N_8751,N_7205,N_6805);
nand U8752 (N_8752,N_7714,N_7776);
and U8753 (N_8753,N_6971,N_7241);
nand U8754 (N_8754,N_7000,N_7774);
or U8755 (N_8755,N_7191,N_6106);
and U8756 (N_8756,N_7708,N_7275);
nand U8757 (N_8757,N_7265,N_7690);
nand U8758 (N_8758,N_7284,N_7782);
nand U8759 (N_8759,N_7050,N_7501);
nor U8760 (N_8760,N_7885,N_6588);
nor U8761 (N_8761,N_7310,N_6655);
and U8762 (N_8762,N_6702,N_7292);
and U8763 (N_8763,N_6107,N_6305);
or U8764 (N_8764,N_7223,N_6180);
nand U8765 (N_8765,N_7074,N_7585);
and U8766 (N_8766,N_7493,N_7980);
or U8767 (N_8767,N_6537,N_6865);
and U8768 (N_8768,N_6963,N_7935);
nor U8769 (N_8769,N_6878,N_6196);
or U8770 (N_8770,N_6418,N_7464);
nor U8771 (N_8771,N_6836,N_6756);
nand U8772 (N_8772,N_6924,N_6887);
or U8773 (N_8773,N_6525,N_7675);
and U8774 (N_8774,N_7897,N_7094);
nor U8775 (N_8775,N_7857,N_6339);
nand U8776 (N_8776,N_7163,N_6965);
nor U8777 (N_8777,N_7154,N_7757);
nor U8778 (N_8778,N_6019,N_6237);
nor U8779 (N_8779,N_6855,N_7026);
and U8780 (N_8780,N_6079,N_7318);
nor U8781 (N_8781,N_7303,N_7162);
nand U8782 (N_8782,N_6359,N_6807);
nand U8783 (N_8783,N_7931,N_6127);
or U8784 (N_8784,N_6376,N_7644);
nand U8785 (N_8785,N_6408,N_7328);
xnor U8786 (N_8786,N_6362,N_6178);
nor U8787 (N_8787,N_6875,N_6859);
nand U8788 (N_8788,N_7070,N_7158);
xnor U8789 (N_8789,N_7982,N_6189);
or U8790 (N_8790,N_6800,N_7027);
nor U8791 (N_8791,N_7137,N_7142);
and U8792 (N_8792,N_7399,N_6521);
or U8793 (N_8793,N_7570,N_6697);
nand U8794 (N_8794,N_7535,N_6994);
and U8795 (N_8795,N_7067,N_7997);
xnor U8796 (N_8796,N_7839,N_7800);
and U8797 (N_8797,N_7444,N_6902);
or U8798 (N_8798,N_7396,N_6671);
or U8799 (N_8799,N_6291,N_6565);
and U8800 (N_8800,N_7462,N_6182);
nor U8801 (N_8801,N_7859,N_6253);
nor U8802 (N_8802,N_7582,N_6312);
or U8803 (N_8803,N_7235,N_6327);
nand U8804 (N_8804,N_6190,N_7659);
nand U8805 (N_8805,N_6458,N_6891);
and U8806 (N_8806,N_7945,N_7108);
xor U8807 (N_8807,N_6614,N_6744);
nor U8808 (N_8808,N_6116,N_7168);
nor U8809 (N_8809,N_7677,N_6379);
and U8810 (N_8810,N_6007,N_7222);
or U8811 (N_8811,N_6037,N_7052);
and U8812 (N_8812,N_6234,N_6477);
nand U8813 (N_8813,N_7512,N_7534);
and U8814 (N_8814,N_6325,N_6063);
or U8815 (N_8815,N_6424,N_7889);
xor U8816 (N_8816,N_6835,N_7041);
nand U8817 (N_8817,N_7528,N_6592);
nor U8818 (N_8818,N_7187,N_6694);
or U8819 (N_8819,N_7840,N_6167);
and U8820 (N_8820,N_6544,N_6541);
and U8821 (N_8821,N_6142,N_7217);
nand U8822 (N_8822,N_7584,N_7540);
nor U8823 (N_8823,N_7633,N_7720);
xor U8824 (N_8824,N_7115,N_7786);
nor U8825 (N_8825,N_7446,N_7511);
nor U8826 (N_8826,N_7957,N_7804);
nand U8827 (N_8827,N_7831,N_7031);
nand U8828 (N_8828,N_6001,N_6165);
or U8829 (N_8829,N_7569,N_6329);
and U8830 (N_8830,N_7767,N_6911);
nor U8831 (N_8831,N_7196,N_7313);
xor U8832 (N_8832,N_6238,N_7449);
nand U8833 (N_8833,N_7370,N_6457);
and U8834 (N_8834,N_7308,N_7685);
and U8835 (N_8835,N_7974,N_6976);
xor U8836 (N_8836,N_7259,N_6947);
nand U8837 (N_8837,N_7664,N_7418);
or U8838 (N_8838,N_7188,N_7448);
xnor U8839 (N_8839,N_7628,N_6912);
or U8840 (N_8840,N_7770,N_7175);
and U8841 (N_8841,N_6644,N_6991);
or U8842 (N_8842,N_6806,N_7996);
nor U8843 (N_8843,N_7874,N_6857);
or U8844 (N_8844,N_6286,N_6193);
nand U8845 (N_8845,N_6583,N_6497);
xor U8846 (N_8846,N_6031,N_7507);
nand U8847 (N_8847,N_7474,N_6161);
nand U8848 (N_8848,N_7282,N_6482);
nand U8849 (N_8849,N_7856,N_7376);
or U8850 (N_8850,N_7211,N_6663);
and U8851 (N_8851,N_7771,N_7174);
and U8852 (N_8852,N_6426,N_6130);
nand U8853 (N_8853,N_7891,N_7976);
nor U8854 (N_8854,N_7342,N_7167);
or U8855 (N_8855,N_7549,N_7452);
nor U8856 (N_8856,N_7476,N_7878);
xnor U8857 (N_8857,N_7753,N_7726);
or U8858 (N_8858,N_6534,N_7561);
nor U8859 (N_8859,N_6597,N_6538);
nand U8860 (N_8860,N_6704,N_6232);
xor U8861 (N_8861,N_6064,N_6771);
and U8862 (N_8862,N_7940,N_6578);
nor U8863 (N_8863,N_6554,N_7298);
and U8864 (N_8864,N_7744,N_6026);
nand U8865 (N_8865,N_7851,N_6003);
nand U8866 (N_8866,N_6047,N_7305);
nand U8867 (N_8867,N_7815,N_6790);
or U8868 (N_8868,N_6275,N_6879);
and U8869 (N_8869,N_6615,N_6024);
or U8870 (N_8870,N_7003,N_6530);
nand U8871 (N_8871,N_7741,N_6089);
nand U8872 (N_8872,N_7988,N_6169);
nand U8873 (N_8873,N_6429,N_6280);
nor U8874 (N_8874,N_7990,N_7133);
nand U8875 (N_8875,N_7227,N_6633);
nand U8876 (N_8876,N_6333,N_6170);
nor U8877 (N_8877,N_6104,N_7025);
nand U8878 (N_8878,N_6579,N_6071);
xor U8879 (N_8879,N_6393,N_7608);
nand U8880 (N_8880,N_6244,N_7823);
and U8881 (N_8881,N_6062,N_6639);
nand U8882 (N_8882,N_6029,N_6626);
nand U8883 (N_8883,N_6985,N_6387);
or U8884 (N_8884,N_7012,N_6152);
nand U8885 (N_8885,N_7520,N_6982);
or U8886 (N_8886,N_6243,N_7872);
nand U8887 (N_8887,N_6337,N_6346);
xnor U8888 (N_8888,N_6832,N_7678);
nor U8889 (N_8889,N_6430,N_7348);
nor U8890 (N_8890,N_6422,N_6274);
nand U8891 (N_8891,N_6733,N_7763);
nand U8892 (N_8892,N_7546,N_7896);
and U8893 (N_8893,N_6322,N_7482);
and U8894 (N_8894,N_6960,N_6781);
nor U8895 (N_8895,N_7083,N_7294);
nor U8896 (N_8896,N_6825,N_6987);
nand U8897 (N_8897,N_6298,N_7021);
or U8898 (N_8898,N_6791,N_6252);
and U8899 (N_8899,N_7161,N_7955);
nor U8900 (N_8900,N_7312,N_6374);
nor U8901 (N_8901,N_6817,N_6827);
nand U8902 (N_8902,N_7739,N_6394);
xnor U8903 (N_8903,N_7323,N_6535);
or U8904 (N_8904,N_7061,N_6240);
or U8905 (N_8905,N_6868,N_6526);
nand U8906 (N_8906,N_7135,N_6350);
xnor U8907 (N_8907,N_7571,N_7219);
nor U8908 (N_8908,N_6126,N_6166);
and U8909 (N_8909,N_7667,N_6411);
and U8910 (N_8910,N_6204,N_6179);
nand U8911 (N_8911,N_7531,N_6403);
nand U8912 (N_8912,N_6439,N_7060);
or U8913 (N_8913,N_6081,N_7674);
nand U8914 (N_8914,N_6044,N_7573);
nand U8915 (N_8915,N_7103,N_6414);
or U8916 (N_8916,N_6035,N_6194);
nor U8917 (N_8917,N_6953,N_6646);
and U8918 (N_8918,N_7518,N_6086);
and U8919 (N_8919,N_6990,N_7755);
nor U8920 (N_8920,N_6461,N_7537);
or U8921 (N_8921,N_6017,N_6529);
xnor U8922 (N_8922,N_6613,N_7111);
and U8923 (N_8923,N_7620,N_7964);
and U8924 (N_8924,N_6808,N_6448);
xor U8925 (N_8925,N_6637,N_6703);
xor U8926 (N_8926,N_7723,N_7002);
nand U8927 (N_8927,N_6665,N_6741);
nor U8928 (N_8928,N_6451,N_6456);
nor U8929 (N_8929,N_6263,N_7287);
and U8930 (N_8930,N_7203,N_7692);
and U8931 (N_8931,N_7477,N_7818);
or U8932 (N_8932,N_6436,N_7490);
nand U8933 (N_8933,N_7311,N_6484);
nor U8934 (N_8934,N_7645,N_7404);
and U8935 (N_8935,N_6576,N_6254);
or U8936 (N_8936,N_7661,N_6593);
or U8937 (N_8937,N_7023,N_6981);
xnor U8938 (N_8938,N_6236,N_7779);
nor U8939 (N_8939,N_7796,N_7407);
nor U8940 (N_8940,N_7488,N_6042);
xnor U8941 (N_8941,N_7498,N_7621);
or U8942 (N_8942,N_7916,N_6500);
nand U8943 (N_8943,N_6602,N_7375);
nand U8944 (N_8944,N_7959,N_6324);
and U8945 (N_8945,N_6103,N_6558);
or U8946 (N_8946,N_7344,N_6828);
nand U8947 (N_8947,N_7029,N_7654);
nand U8948 (N_8948,N_6784,N_6886);
or U8949 (N_8949,N_7400,N_6860);
xor U8950 (N_8950,N_7190,N_7567);
nand U8951 (N_8951,N_7793,N_6211);
nor U8952 (N_8952,N_6151,N_6289);
and U8953 (N_8953,N_6719,N_7609);
nand U8954 (N_8954,N_6927,N_6034);
or U8955 (N_8955,N_6320,N_6620);
nand U8956 (N_8956,N_7656,N_6445);
and U8957 (N_8957,N_6649,N_7765);
nand U8958 (N_8958,N_7791,N_6777);
nand U8959 (N_8959,N_6684,N_7625);
and U8960 (N_8960,N_6636,N_7792);
nor U8961 (N_8961,N_6143,N_7748);
and U8962 (N_8962,N_7925,N_6892);
or U8963 (N_8963,N_7565,N_7260);
or U8964 (N_8964,N_6607,N_7975);
or U8965 (N_8965,N_6540,N_7445);
nor U8966 (N_8966,N_7333,N_7469);
or U8967 (N_8967,N_7330,N_7713);
nor U8968 (N_8968,N_6925,N_6739);
and U8969 (N_8969,N_7267,N_7519);
nand U8970 (N_8970,N_7149,N_7295);
nand U8971 (N_8971,N_7920,N_7838);
or U8972 (N_8972,N_7079,N_7936);
and U8973 (N_8973,N_7495,N_6881);
nand U8974 (N_8974,N_7441,N_7986);
xor U8975 (N_8975,N_7607,N_6707);
and U8976 (N_8976,N_7216,N_6303);
nand U8977 (N_8977,N_7315,N_6226);
nor U8978 (N_8978,N_6215,N_7701);
or U8979 (N_8979,N_7922,N_7483);
xor U8980 (N_8980,N_6743,N_7136);
or U8981 (N_8981,N_6389,N_6993);
and U8982 (N_8982,N_6931,N_6951);
or U8983 (N_8983,N_7020,N_7710);
nand U8984 (N_8984,N_7005,N_7932);
nand U8985 (N_8985,N_7225,N_6699);
nor U8986 (N_8986,N_7775,N_6045);
xor U8987 (N_8987,N_6717,N_6340);
or U8988 (N_8988,N_7276,N_7480);
xnor U8989 (N_8989,N_7353,N_6608);
xor U8990 (N_8990,N_7085,N_6421);
xnor U8991 (N_8991,N_7390,N_6656);
xor U8992 (N_8992,N_7228,N_6465);
or U8993 (N_8993,N_7732,N_6587);
or U8994 (N_8994,N_7699,N_6755);
and U8995 (N_8995,N_6623,N_7890);
or U8996 (N_8996,N_7822,N_7209);
xnor U8997 (N_8997,N_7355,N_6384);
nand U8998 (N_8998,N_7340,N_6470);
or U8999 (N_8999,N_7712,N_6641);
and U9000 (N_9000,N_6447,N_7662);
nand U9001 (N_9001,N_7470,N_6566);
xor U9002 (N_9002,N_7918,N_7464);
xor U9003 (N_9003,N_6746,N_7743);
xnor U9004 (N_9004,N_7120,N_6628);
nand U9005 (N_9005,N_6924,N_7624);
or U9006 (N_9006,N_6104,N_7267);
nor U9007 (N_9007,N_7904,N_6702);
and U9008 (N_9008,N_6001,N_7746);
nand U9009 (N_9009,N_6661,N_7296);
nand U9010 (N_9010,N_6723,N_7667);
nor U9011 (N_9011,N_6869,N_7194);
nand U9012 (N_9012,N_7143,N_6764);
and U9013 (N_9013,N_6322,N_7085);
nand U9014 (N_9014,N_6406,N_6733);
nor U9015 (N_9015,N_6966,N_6705);
or U9016 (N_9016,N_7629,N_7339);
or U9017 (N_9017,N_7783,N_7343);
or U9018 (N_9018,N_6660,N_6736);
nand U9019 (N_9019,N_7868,N_6525);
or U9020 (N_9020,N_7779,N_7125);
nor U9021 (N_9021,N_6737,N_6646);
nor U9022 (N_9022,N_7388,N_6322);
or U9023 (N_9023,N_6519,N_7598);
and U9024 (N_9024,N_6749,N_6451);
or U9025 (N_9025,N_6913,N_6497);
nand U9026 (N_9026,N_7943,N_7235);
xor U9027 (N_9027,N_7794,N_7561);
nor U9028 (N_9028,N_7975,N_6512);
and U9029 (N_9029,N_6555,N_7951);
or U9030 (N_9030,N_6965,N_7982);
nand U9031 (N_9031,N_6717,N_6853);
and U9032 (N_9032,N_7441,N_6248);
or U9033 (N_9033,N_6692,N_7294);
xnor U9034 (N_9034,N_7988,N_6371);
and U9035 (N_9035,N_7706,N_6846);
nand U9036 (N_9036,N_6490,N_6165);
nor U9037 (N_9037,N_7340,N_7384);
nor U9038 (N_9038,N_6552,N_6670);
nor U9039 (N_9039,N_6709,N_7535);
nor U9040 (N_9040,N_6991,N_7340);
nor U9041 (N_9041,N_6102,N_7845);
nor U9042 (N_9042,N_6580,N_6937);
or U9043 (N_9043,N_7551,N_7437);
and U9044 (N_9044,N_7289,N_7432);
nand U9045 (N_9045,N_7970,N_6589);
or U9046 (N_9046,N_6523,N_6351);
nor U9047 (N_9047,N_6407,N_6469);
nor U9048 (N_9048,N_6320,N_7085);
nor U9049 (N_9049,N_7085,N_6229);
or U9050 (N_9050,N_7092,N_7497);
nor U9051 (N_9051,N_7306,N_6403);
nand U9052 (N_9052,N_6893,N_7661);
nor U9053 (N_9053,N_6619,N_6913);
nor U9054 (N_9054,N_6373,N_7650);
nand U9055 (N_9055,N_7851,N_6290);
and U9056 (N_9056,N_7208,N_6823);
and U9057 (N_9057,N_6597,N_6382);
nor U9058 (N_9058,N_7740,N_7049);
or U9059 (N_9059,N_6364,N_6712);
nand U9060 (N_9060,N_6084,N_7073);
nand U9061 (N_9061,N_6488,N_7648);
nand U9062 (N_9062,N_7209,N_6783);
and U9063 (N_9063,N_7548,N_7985);
nor U9064 (N_9064,N_7743,N_7118);
and U9065 (N_9065,N_7373,N_6721);
and U9066 (N_9066,N_7348,N_7086);
or U9067 (N_9067,N_6882,N_7123);
nand U9068 (N_9068,N_6821,N_6649);
nand U9069 (N_9069,N_7908,N_7847);
or U9070 (N_9070,N_7268,N_6104);
or U9071 (N_9071,N_7753,N_7474);
nor U9072 (N_9072,N_7981,N_6477);
or U9073 (N_9073,N_7546,N_6410);
or U9074 (N_9074,N_7469,N_6778);
or U9075 (N_9075,N_7077,N_7088);
and U9076 (N_9076,N_7722,N_6841);
nand U9077 (N_9077,N_6399,N_7466);
or U9078 (N_9078,N_6707,N_7331);
or U9079 (N_9079,N_7633,N_6668);
nand U9080 (N_9080,N_6785,N_7220);
or U9081 (N_9081,N_6529,N_6575);
or U9082 (N_9082,N_7058,N_7674);
and U9083 (N_9083,N_7038,N_7841);
nor U9084 (N_9084,N_7087,N_6435);
or U9085 (N_9085,N_7878,N_7967);
or U9086 (N_9086,N_6694,N_7327);
and U9087 (N_9087,N_6878,N_7126);
or U9088 (N_9088,N_7879,N_7666);
or U9089 (N_9089,N_6949,N_6666);
nor U9090 (N_9090,N_7053,N_6482);
nand U9091 (N_9091,N_6530,N_7398);
xnor U9092 (N_9092,N_7362,N_7887);
nor U9093 (N_9093,N_7624,N_7840);
nand U9094 (N_9094,N_7812,N_7609);
nor U9095 (N_9095,N_7714,N_7193);
or U9096 (N_9096,N_6032,N_7440);
nor U9097 (N_9097,N_6120,N_6260);
nor U9098 (N_9098,N_6106,N_7053);
nor U9099 (N_9099,N_7901,N_7431);
nor U9100 (N_9100,N_6919,N_7668);
or U9101 (N_9101,N_6914,N_7683);
or U9102 (N_9102,N_7202,N_7633);
and U9103 (N_9103,N_7245,N_6025);
nor U9104 (N_9104,N_6756,N_7437);
nand U9105 (N_9105,N_6007,N_7601);
or U9106 (N_9106,N_7848,N_7583);
and U9107 (N_9107,N_6625,N_7429);
or U9108 (N_9108,N_7332,N_7405);
or U9109 (N_9109,N_7649,N_7341);
and U9110 (N_9110,N_6075,N_6833);
nor U9111 (N_9111,N_6434,N_7370);
nand U9112 (N_9112,N_6584,N_6404);
and U9113 (N_9113,N_6983,N_6900);
and U9114 (N_9114,N_7870,N_7651);
nand U9115 (N_9115,N_6480,N_7298);
nand U9116 (N_9116,N_7897,N_6068);
nor U9117 (N_9117,N_6540,N_6879);
and U9118 (N_9118,N_7925,N_7614);
nand U9119 (N_9119,N_7113,N_6729);
nor U9120 (N_9120,N_6260,N_6416);
nand U9121 (N_9121,N_6314,N_6734);
xnor U9122 (N_9122,N_6813,N_7937);
or U9123 (N_9123,N_7820,N_7382);
and U9124 (N_9124,N_7460,N_6458);
and U9125 (N_9125,N_7131,N_7281);
nand U9126 (N_9126,N_6128,N_6983);
nor U9127 (N_9127,N_6850,N_6442);
and U9128 (N_9128,N_7698,N_6569);
or U9129 (N_9129,N_6093,N_7815);
nor U9130 (N_9130,N_7515,N_6841);
and U9131 (N_9131,N_7067,N_6429);
nand U9132 (N_9132,N_7240,N_6612);
and U9133 (N_9133,N_6312,N_7408);
xnor U9134 (N_9134,N_7649,N_6077);
nand U9135 (N_9135,N_6270,N_7018);
nand U9136 (N_9136,N_7445,N_7266);
xor U9137 (N_9137,N_7366,N_7121);
nand U9138 (N_9138,N_6008,N_7724);
nand U9139 (N_9139,N_7345,N_6516);
or U9140 (N_9140,N_7125,N_6670);
and U9141 (N_9141,N_6690,N_6293);
nor U9142 (N_9142,N_7787,N_6191);
xor U9143 (N_9143,N_7783,N_7138);
nand U9144 (N_9144,N_7671,N_6204);
xor U9145 (N_9145,N_7204,N_7221);
nor U9146 (N_9146,N_7963,N_6446);
and U9147 (N_9147,N_7656,N_6030);
nor U9148 (N_9148,N_7322,N_6480);
or U9149 (N_9149,N_6456,N_6280);
xnor U9150 (N_9150,N_6423,N_6589);
nor U9151 (N_9151,N_6098,N_7248);
and U9152 (N_9152,N_7858,N_7816);
nand U9153 (N_9153,N_6635,N_6997);
nand U9154 (N_9154,N_7226,N_7103);
or U9155 (N_9155,N_6735,N_6329);
nand U9156 (N_9156,N_6383,N_6505);
or U9157 (N_9157,N_6697,N_6556);
nor U9158 (N_9158,N_6443,N_7869);
or U9159 (N_9159,N_6644,N_6965);
or U9160 (N_9160,N_6108,N_6413);
xor U9161 (N_9161,N_6331,N_7828);
and U9162 (N_9162,N_7350,N_6749);
nand U9163 (N_9163,N_6448,N_7867);
nor U9164 (N_9164,N_7480,N_6038);
xor U9165 (N_9165,N_6275,N_6065);
nor U9166 (N_9166,N_6312,N_7699);
or U9167 (N_9167,N_6518,N_7354);
nor U9168 (N_9168,N_6656,N_6596);
nor U9169 (N_9169,N_7999,N_7865);
and U9170 (N_9170,N_6829,N_7897);
xnor U9171 (N_9171,N_6318,N_6961);
and U9172 (N_9172,N_6318,N_6859);
xnor U9173 (N_9173,N_6904,N_7399);
and U9174 (N_9174,N_7210,N_6187);
or U9175 (N_9175,N_6902,N_7565);
nor U9176 (N_9176,N_7979,N_7954);
nor U9177 (N_9177,N_6842,N_7924);
or U9178 (N_9178,N_6995,N_7110);
or U9179 (N_9179,N_7397,N_6156);
nor U9180 (N_9180,N_6195,N_7227);
or U9181 (N_9181,N_6757,N_7800);
or U9182 (N_9182,N_6241,N_7794);
nand U9183 (N_9183,N_6292,N_6513);
or U9184 (N_9184,N_6515,N_7889);
nor U9185 (N_9185,N_6593,N_6714);
and U9186 (N_9186,N_7723,N_7337);
nor U9187 (N_9187,N_6760,N_6419);
or U9188 (N_9188,N_7863,N_7817);
and U9189 (N_9189,N_6244,N_7804);
nand U9190 (N_9190,N_6956,N_6639);
or U9191 (N_9191,N_6895,N_6399);
or U9192 (N_9192,N_7931,N_6187);
xor U9193 (N_9193,N_6415,N_6233);
or U9194 (N_9194,N_6062,N_7066);
nor U9195 (N_9195,N_7262,N_6826);
nand U9196 (N_9196,N_7747,N_7325);
nor U9197 (N_9197,N_6726,N_6895);
nor U9198 (N_9198,N_7450,N_7614);
or U9199 (N_9199,N_7471,N_7000);
nor U9200 (N_9200,N_7236,N_7664);
or U9201 (N_9201,N_7124,N_6520);
or U9202 (N_9202,N_6816,N_7077);
nor U9203 (N_9203,N_7720,N_6424);
nand U9204 (N_9204,N_7505,N_7711);
xnor U9205 (N_9205,N_6415,N_6929);
nor U9206 (N_9206,N_6085,N_7178);
or U9207 (N_9207,N_6815,N_6917);
nor U9208 (N_9208,N_7858,N_6793);
or U9209 (N_9209,N_6091,N_7435);
and U9210 (N_9210,N_6895,N_7006);
nand U9211 (N_9211,N_6152,N_7110);
nand U9212 (N_9212,N_6296,N_7693);
nand U9213 (N_9213,N_7193,N_7363);
nand U9214 (N_9214,N_7030,N_6620);
or U9215 (N_9215,N_6296,N_7049);
or U9216 (N_9216,N_6835,N_7397);
nand U9217 (N_9217,N_6103,N_6234);
and U9218 (N_9218,N_7184,N_7511);
or U9219 (N_9219,N_6780,N_6889);
or U9220 (N_9220,N_7797,N_7520);
and U9221 (N_9221,N_6496,N_6212);
nand U9222 (N_9222,N_7354,N_7227);
nor U9223 (N_9223,N_7878,N_6258);
xnor U9224 (N_9224,N_7043,N_7576);
or U9225 (N_9225,N_7588,N_6985);
xor U9226 (N_9226,N_7635,N_7888);
xor U9227 (N_9227,N_7706,N_6095);
or U9228 (N_9228,N_7896,N_6961);
and U9229 (N_9229,N_7837,N_6031);
or U9230 (N_9230,N_7281,N_7553);
or U9231 (N_9231,N_7047,N_6422);
or U9232 (N_9232,N_7518,N_6008);
or U9233 (N_9233,N_7516,N_7260);
or U9234 (N_9234,N_6593,N_7795);
nand U9235 (N_9235,N_6371,N_6178);
nor U9236 (N_9236,N_6832,N_7984);
and U9237 (N_9237,N_6239,N_7468);
or U9238 (N_9238,N_7434,N_7862);
nor U9239 (N_9239,N_6762,N_7004);
or U9240 (N_9240,N_6610,N_6666);
nor U9241 (N_9241,N_6066,N_6510);
xor U9242 (N_9242,N_7137,N_7750);
xnor U9243 (N_9243,N_7882,N_7424);
nor U9244 (N_9244,N_7089,N_6885);
nand U9245 (N_9245,N_7638,N_7250);
nand U9246 (N_9246,N_7940,N_6515);
nor U9247 (N_9247,N_7675,N_6921);
xor U9248 (N_9248,N_7875,N_6946);
nor U9249 (N_9249,N_7369,N_7011);
and U9250 (N_9250,N_7695,N_6202);
and U9251 (N_9251,N_6474,N_7126);
or U9252 (N_9252,N_7312,N_7733);
nor U9253 (N_9253,N_6674,N_7882);
xnor U9254 (N_9254,N_6958,N_6106);
nand U9255 (N_9255,N_6987,N_6043);
xor U9256 (N_9256,N_7502,N_6089);
nand U9257 (N_9257,N_6218,N_7718);
or U9258 (N_9258,N_6114,N_7812);
or U9259 (N_9259,N_6306,N_6275);
nor U9260 (N_9260,N_7863,N_6966);
nand U9261 (N_9261,N_6310,N_7700);
and U9262 (N_9262,N_6819,N_7047);
and U9263 (N_9263,N_6610,N_7548);
nand U9264 (N_9264,N_6127,N_7815);
nand U9265 (N_9265,N_7134,N_7641);
nand U9266 (N_9266,N_6722,N_7305);
or U9267 (N_9267,N_6772,N_6552);
nand U9268 (N_9268,N_6051,N_6409);
xnor U9269 (N_9269,N_7923,N_7067);
and U9270 (N_9270,N_7643,N_7376);
and U9271 (N_9271,N_6259,N_7315);
and U9272 (N_9272,N_7768,N_6362);
nor U9273 (N_9273,N_6659,N_7844);
nand U9274 (N_9274,N_6261,N_7128);
and U9275 (N_9275,N_7246,N_6698);
nand U9276 (N_9276,N_7575,N_6639);
or U9277 (N_9277,N_6646,N_7381);
nand U9278 (N_9278,N_6688,N_7546);
nor U9279 (N_9279,N_6430,N_6582);
and U9280 (N_9280,N_7672,N_7941);
or U9281 (N_9281,N_7715,N_7892);
or U9282 (N_9282,N_7447,N_7647);
nand U9283 (N_9283,N_6686,N_7534);
nor U9284 (N_9284,N_7305,N_7172);
or U9285 (N_9285,N_7778,N_7182);
nand U9286 (N_9286,N_6166,N_6134);
nor U9287 (N_9287,N_7934,N_7089);
nor U9288 (N_9288,N_6736,N_7138);
nand U9289 (N_9289,N_6599,N_7439);
nand U9290 (N_9290,N_7688,N_6857);
nor U9291 (N_9291,N_7050,N_6249);
nor U9292 (N_9292,N_6223,N_7536);
xnor U9293 (N_9293,N_7562,N_7786);
and U9294 (N_9294,N_7081,N_6306);
nand U9295 (N_9295,N_6289,N_6548);
and U9296 (N_9296,N_6625,N_7080);
or U9297 (N_9297,N_7935,N_6279);
and U9298 (N_9298,N_6692,N_7144);
nand U9299 (N_9299,N_6983,N_6526);
nor U9300 (N_9300,N_6079,N_7850);
nand U9301 (N_9301,N_6492,N_7615);
nor U9302 (N_9302,N_6192,N_7141);
xor U9303 (N_9303,N_7255,N_7034);
or U9304 (N_9304,N_6871,N_7953);
or U9305 (N_9305,N_7549,N_7907);
and U9306 (N_9306,N_6710,N_6170);
or U9307 (N_9307,N_6523,N_7249);
xnor U9308 (N_9308,N_7308,N_6157);
nand U9309 (N_9309,N_6591,N_7368);
or U9310 (N_9310,N_7819,N_6224);
and U9311 (N_9311,N_6812,N_6086);
xor U9312 (N_9312,N_7758,N_6867);
nand U9313 (N_9313,N_7565,N_6298);
nand U9314 (N_9314,N_6085,N_6590);
and U9315 (N_9315,N_7110,N_7524);
xor U9316 (N_9316,N_6574,N_7430);
and U9317 (N_9317,N_7463,N_6920);
and U9318 (N_9318,N_6261,N_7173);
or U9319 (N_9319,N_6815,N_6089);
nand U9320 (N_9320,N_7952,N_7627);
and U9321 (N_9321,N_6602,N_7270);
and U9322 (N_9322,N_7412,N_7917);
nand U9323 (N_9323,N_6433,N_6420);
or U9324 (N_9324,N_7361,N_7430);
and U9325 (N_9325,N_6483,N_7365);
xor U9326 (N_9326,N_7220,N_7273);
nand U9327 (N_9327,N_7101,N_6407);
and U9328 (N_9328,N_7827,N_7336);
xor U9329 (N_9329,N_6207,N_6731);
nand U9330 (N_9330,N_6918,N_7010);
or U9331 (N_9331,N_6064,N_7235);
xnor U9332 (N_9332,N_6503,N_6395);
and U9333 (N_9333,N_6434,N_7898);
nor U9334 (N_9334,N_6115,N_7427);
nand U9335 (N_9335,N_6924,N_7458);
or U9336 (N_9336,N_7672,N_6566);
nand U9337 (N_9337,N_7342,N_6090);
or U9338 (N_9338,N_7943,N_7928);
nand U9339 (N_9339,N_7362,N_7757);
and U9340 (N_9340,N_6965,N_7889);
and U9341 (N_9341,N_7201,N_6241);
nor U9342 (N_9342,N_7543,N_7395);
or U9343 (N_9343,N_7876,N_7814);
nor U9344 (N_9344,N_7823,N_6978);
nor U9345 (N_9345,N_7345,N_6346);
or U9346 (N_9346,N_6805,N_7631);
and U9347 (N_9347,N_6366,N_6814);
nor U9348 (N_9348,N_6353,N_6550);
nor U9349 (N_9349,N_7790,N_6614);
and U9350 (N_9350,N_6277,N_7461);
xnor U9351 (N_9351,N_6671,N_7429);
nand U9352 (N_9352,N_7000,N_6195);
nand U9353 (N_9353,N_6066,N_6077);
xnor U9354 (N_9354,N_7199,N_6395);
or U9355 (N_9355,N_6108,N_6170);
nand U9356 (N_9356,N_7671,N_6221);
or U9357 (N_9357,N_7737,N_7670);
xnor U9358 (N_9358,N_7654,N_6374);
xor U9359 (N_9359,N_7582,N_6327);
and U9360 (N_9360,N_7802,N_6994);
nor U9361 (N_9361,N_6922,N_6242);
or U9362 (N_9362,N_7567,N_7112);
or U9363 (N_9363,N_6889,N_7743);
nand U9364 (N_9364,N_7439,N_7576);
nor U9365 (N_9365,N_7662,N_6694);
or U9366 (N_9366,N_6646,N_7708);
and U9367 (N_9367,N_6741,N_7349);
nand U9368 (N_9368,N_7761,N_7210);
or U9369 (N_9369,N_6052,N_6705);
nor U9370 (N_9370,N_7641,N_7801);
nand U9371 (N_9371,N_7593,N_6300);
and U9372 (N_9372,N_7455,N_6801);
nand U9373 (N_9373,N_6049,N_7258);
and U9374 (N_9374,N_6344,N_7812);
nor U9375 (N_9375,N_6446,N_7007);
nand U9376 (N_9376,N_6191,N_7246);
and U9377 (N_9377,N_6050,N_7862);
xnor U9378 (N_9378,N_6242,N_7842);
or U9379 (N_9379,N_6774,N_7794);
nand U9380 (N_9380,N_6398,N_7756);
xor U9381 (N_9381,N_7029,N_7789);
or U9382 (N_9382,N_6139,N_7906);
nand U9383 (N_9383,N_7751,N_7792);
and U9384 (N_9384,N_6354,N_6712);
or U9385 (N_9385,N_7598,N_7115);
and U9386 (N_9386,N_6403,N_7123);
or U9387 (N_9387,N_6062,N_7109);
nand U9388 (N_9388,N_6722,N_7041);
nor U9389 (N_9389,N_7200,N_6415);
nor U9390 (N_9390,N_6847,N_7754);
xnor U9391 (N_9391,N_6574,N_6106);
or U9392 (N_9392,N_7794,N_7375);
and U9393 (N_9393,N_6219,N_6588);
nand U9394 (N_9394,N_7568,N_6338);
xor U9395 (N_9395,N_7866,N_6977);
or U9396 (N_9396,N_7159,N_7938);
nor U9397 (N_9397,N_6828,N_7475);
xnor U9398 (N_9398,N_6947,N_7271);
nand U9399 (N_9399,N_6495,N_6838);
and U9400 (N_9400,N_6196,N_6786);
nor U9401 (N_9401,N_7492,N_6198);
nand U9402 (N_9402,N_7636,N_6754);
nand U9403 (N_9403,N_7654,N_7847);
nand U9404 (N_9404,N_6345,N_6201);
nor U9405 (N_9405,N_6076,N_6909);
or U9406 (N_9406,N_6923,N_7717);
or U9407 (N_9407,N_7361,N_6925);
or U9408 (N_9408,N_6304,N_7700);
nand U9409 (N_9409,N_7326,N_7809);
nand U9410 (N_9410,N_6227,N_7456);
or U9411 (N_9411,N_6572,N_7671);
and U9412 (N_9412,N_6443,N_7450);
nand U9413 (N_9413,N_7268,N_7586);
nor U9414 (N_9414,N_6266,N_6003);
nor U9415 (N_9415,N_6616,N_6662);
xnor U9416 (N_9416,N_6680,N_6244);
xnor U9417 (N_9417,N_7040,N_6136);
or U9418 (N_9418,N_7627,N_6650);
or U9419 (N_9419,N_7789,N_6280);
nand U9420 (N_9420,N_7517,N_7469);
nand U9421 (N_9421,N_7659,N_7405);
and U9422 (N_9422,N_6884,N_6347);
or U9423 (N_9423,N_7378,N_6755);
nor U9424 (N_9424,N_7069,N_7634);
or U9425 (N_9425,N_6423,N_7521);
nand U9426 (N_9426,N_7887,N_6528);
nor U9427 (N_9427,N_6307,N_7788);
nor U9428 (N_9428,N_7905,N_6827);
and U9429 (N_9429,N_7763,N_7750);
nand U9430 (N_9430,N_6228,N_6374);
xor U9431 (N_9431,N_6817,N_7949);
and U9432 (N_9432,N_6430,N_7425);
nor U9433 (N_9433,N_6719,N_7524);
or U9434 (N_9434,N_6443,N_7679);
and U9435 (N_9435,N_6322,N_6091);
or U9436 (N_9436,N_6627,N_7078);
nor U9437 (N_9437,N_6869,N_6084);
and U9438 (N_9438,N_7938,N_6443);
nand U9439 (N_9439,N_7877,N_6167);
nor U9440 (N_9440,N_6837,N_7237);
nor U9441 (N_9441,N_6872,N_7798);
nor U9442 (N_9442,N_7613,N_6842);
or U9443 (N_9443,N_7921,N_6538);
nor U9444 (N_9444,N_6278,N_7822);
or U9445 (N_9445,N_7583,N_6577);
or U9446 (N_9446,N_7663,N_7109);
and U9447 (N_9447,N_7144,N_6569);
nor U9448 (N_9448,N_6292,N_6994);
nor U9449 (N_9449,N_6834,N_6078);
nand U9450 (N_9450,N_6069,N_6112);
and U9451 (N_9451,N_7847,N_7882);
or U9452 (N_9452,N_7136,N_7294);
nor U9453 (N_9453,N_7475,N_6463);
nor U9454 (N_9454,N_7253,N_6249);
nor U9455 (N_9455,N_6777,N_7424);
nand U9456 (N_9456,N_7807,N_7784);
or U9457 (N_9457,N_7333,N_7822);
nor U9458 (N_9458,N_6815,N_7720);
and U9459 (N_9459,N_6579,N_7811);
xor U9460 (N_9460,N_6008,N_7727);
and U9461 (N_9461,N_7359,N_6328);
or U9462 (N_9462,N_6671,N_6405);
or U9463 (N_9463,N_6565,N_6944);
and U9464 (N_9464,N_6884,N_7304);
nor U9465 (N_9465,N_7068,N_7493);
nand U9466 (N_9466,N_7894,N_7684);
nor U9467 (N_9467,N_7692,N_7591);
or U9468 (N_9468,N_7924,N_7957);
nor U9469 (N_9469,N_6597,N_6946);
nand U9470 (N_9470,N_7044,N_7156);
or U9471 (N_9471,N_7209,N_6114);
xnor U9472 (N_9472,N_6073,N_6149);
nand U9473 (N_9473,N_7687,N_6223);
and U9474 (N_9474,N_7650,N_7208);
nand U9475 (N_9475,N_6581,N_6477);
and U9476 (N_9476,N_6833,N_6491);
and U9477 (N_9477,N_6739,N_6611);
nor U9478 (N_9478,N_6311,N_7970);
or U9479 (N_9479,N_6817,N_6276);
nand U9480 (N_9480,N_7627,N_6091);
nor U9481 (N_9481,N_7430,N_7543);
or U9482 (N_9482,N_6016,N_6356);
xnor U9483 (N_9483,N_7485,N_6476);
or U9484 (N_9484,N_7417,N_7441);
or U9485 (N_9485,N_6673,N_6446);
or U9486 (N_9486,N_7232,N_6883);
nor U9487 (N_9487,N_6192,N_6099);
nand U9488 (N_9488,N_7163,N_7748);
nor U9489 (N_9489,N_7746,N_7327);
nor U9490 (N_9490,N_7376,N_7346);
or U9491 (N_9491,N_6435,N_7662);
and U9492 (N_9492,N_7593,N_6383);
or U9493 (N_9493,N_7422,N_6520);
or U9494 (N_9494,N_7954,N_6651);
or U9495 (N_9495,N_6462,N_6649);
nor U9496 (N_9496,N_7209,N_6767);
nand U9497 (N_9497,N_7154,N_7628);
nor U9498 (N_9498,N_6712,N_6946);
nor U9499 (N_9499,N_7084,N_7330);
or U9500 (N_9500,N_6610,N_6732);
or U9501 (N_9501,N_6403,N_6384);
nor U9502 (N_9502,N_6746,N_7547);
and U9503 (N_9503,N_6226,N_6921);
nor U9504 (N_9504,N_7019,N_7326);
nand U9505 (N_9505,N_7712,N_7749);
nand U9506 (N_9506,N_6831,N_6419);
nor U9507 (N_9507,N_6339,N_6078);
or U9508 (N_9508,N_6711,N_6865);
nor U9509 (N_9509,N_6898,N_6274);
nor U9510 (N_9510,N_7782,N_7122);
nand U9511 (N_9511,N_7551,N_7762);
nand U9512 (N_9512,N_6373,N_6201);
or U9513 (N_9513,N_7769,N_6360);
nand U9514 (N_9514,N_7570,N_6913);
and U9515 (N_9515,N_6409,N_7950);
or U9516 (N_9516,N_6056,N_6039);
or U9517 (N_9517,N_6769,N_7091);
nor U9518 (N_9518,N_7234,N_6704);
and U9519 (N_9519,N_7156,N_6327);
nor U9520 (N_9520,N_6681,N_6915);
nor U9521 (N_9521,N_7722,N_7723);
nor U9522 (N_9522,N_6999,N_7217);
and U9523 (N_9523,N_7138,N_7834);
nor U9524 (N_9524,N_7408,N_7747);
or U9525 (N_9525,N_6229,N_6509);
nand U9526 (N_9526,N_6803,N_7514);
nor U9527 (N_9527,N_7294,N_7228);
or U9528 (N_9528,N_6285,N_6356);
or U9529 (N_9529,N_7591,N_7730);
or U9530 (N_9530,N_6789,N_6892);
or U9531 (N_9531,N_6084,N_6406);
or U9532 (N_9532,N_7665,N_6018);
nor U9533 (N_9533,N_7940,N_6321);
xnor U9534 (N_9534,N_7616,N_7417);
or U9535 (N_9535,N_7500,N_7114);
and U9536 (N_9536,N_6957,N_6611);
and U9537 (N_9537,N_7238,N_7824);
nor U9538 (N_9538,N_6794,N_6218);
or U9539 (N_9539,N_7797,N_6350);
or U9540 (N_9540,N_7923,N_6114);
nor U9541 (N_9541,N_6100,N_6633);
nor U9542 (N_9542,N_7064,N_6680);
nor U9543 (N_9543,N_6305,N_7615);
or U9544 (N_9544,N_6688,N_6405);
nand U9545 (N_9545,N_6428,N_7382);
and U9546 (N_9546,N_7161,N_7585);
nor U9547 (N_9547,N_6125,N_6497);
nand U9548 (N_9548,N_7902,N_7936);
nand U9549 (N_9549,N_6645,N_7320);
or U9550 (N_9550,N_7946,N_7818);
nand U9551 (N_9551,N_7500,N_7267);
nand U9552 (N_9552,N_7430,N_6009);
nor U9553 (N_9553,N_7825,N_6145);
nor U9554 (N_9554,N_6527,N_7263);
nand U9555 (N_9555,N_7611,N_7633);
nand U9556 (N_9556,N_6840,N_6767);
nand U9557 (N_9557,N_7682,N_7279);
xnor U9558 (N_9558,N_6180,N_6984);
nor U9559 (N_9559,N_6648,N_7726);
and U9560 (N_9560,N_6462,N_7728);
xor U9561 (N_9561,N_7388,N_6946);
nor U9562 (N_9562,N_7435,N_6059);
nor U9563 (N_9563,N_7732,N_6391);
nor U9564 (N_9564,N_7494,N_6863);
nor U9565 (N_9565,N_7488,N_6667);
nand U9566 (N_9566,N_7158,N_7761);
and U9567 (N_9567,N_6809,N_6303);
or U9568 (N_9568,N_7983,N_6619);
nor U9569 (N_9569,N_7682,N_6252);
or U9570 (N_9570,N_6701,N_7888);
and U9571 (N_9571,N_7654,N_7632);
xnor U9572 (N_9572,N_7018,N_6222);
nor U9573 (N_9573,N_6680,N_7097);
or U9574 (N_9574,N_7459,N_7323);
or U9575 (N_9575,N_6169,N_6244);
nor U9576 (N_9576,N_7240,N_7311);
nand U9577 (N_9577,N_6480,N_7026);
and U9578 (N_9578,N_7777,N_6076);
or U9579 (N_9579,N_7931,N_6130);
nand U9580 (N_9580,N_7499,N_7897);
and U9581 (N_9581,N_6323,N_6917);
nor U9582 (N_9582,N_7108,N_7897);
or U9583 (N_9583,N_7188,N_7296);
xnor U9584 (N_9584,N_6610,N_7681);
and U9585 (N_9585,N_6127,N_7000);
or U9586 (N_9586,N_7156,N_7141);
nand U9587 (N_9587,N_7664,N_6711);
nor U9588 (N_9588,N_6143,N_7313);
nand U9589 (N_9589,N_6146,N_7276);
nor U9590 (N_9590,N_6998,N_7273);
nand U9591 (N_9591,N_6062,N_6371);
or U9592 (N_9592,N_6477,N_6179);
nor U9593 (N_9593,N_6291,N_6443);
nand U9594 (N_9594,N_6325,N_6575);
and U9595 (N_9595,N_6127,N_6010);
and U9596 (N_9596,N_7612,N_6825);
or U9597 (N_9597,N_6010,N_6350);
nor U9598 (N_9598,N_6387,N_7329);
nor U9599 (N_9599,N_7683,N_7650);
or U9600 (N_9600,N_6822,N_6028);
and U9601 (N_9601,N_6592,N_7582);
nor U9602 (N_9602,N_7934,N_7445);
or U9603 (N_9603,N_7945,N_7717);
xnor U9604 (N_9604,N_7965,N_7569);
nor U9605 (N_9605,N_7959,N_7441);
and U9606 (N_9606,N_6430,N_6443);
and U9607 (N_9607,N_6557,N_7216);
and U9608 (N_9608,N_7386,N_6767);
xor U9609 (N_9609,N_6571,N_6472);
xnor U9610 (N_9610,N_6232,N_7208);
or U9611 (N_9611,N_7863,N_7737);
nor U9612 (N_9612,N_7137,N_6040);
nand U9613 (N_9613,N_7864,N_6058);
and U9614 (N_9614,N_6953,N_6051);
and U9615 (N_9615,N_7505,N_7322);
nor U9616 (N_9616,N_7886,N_6465);
and U9617 (N_9617,N_7823,N_7865);
and U9618 (N_9618,N_7535,N_6381);
or U9619 (N_9619,N_6156,N_6895);
nor U9620 (N_9620,N_7984,N_6967);
or U9621 (N_9621,N_6450,N_7473);
xnor U9622 (N_9622,N_6178,N_7679);
nand U9623 (N_9623,N_7226,N_6449);
and U9624 (N_9624,N_6902,N_6778);
or U9625 (N_9625,N_6779,N_7916);
nand U9626 (N_9626,N_6793,N_6902);
nand U9627 (N_9627,N_7783,N_6268);
nor U9628 (N_9628,N_6288,N_6597);
nor U9629 (N_9629,N_7838,N_6348);
nor U9630 (N_9630,N_6479,N_6161);
and U9631 (N_9631,N_7928,N_6106);
and U9632 (N_9632,N_7934,N_6658);
or U9633 (N_9633,N_6525,N_6660);
or U9634 (N_9634,N_7525,N_7067);
or U9635 (N_9635,N_6499,N_6021);
nand U9636 (N_9636,N_6986,N_6109);
nor U9637 (N_9637,N_6967,N_6135);
or U9638 (N_9638,N_6511,N_6376);
nand U9639 (N_9639,N_6043,N_7497);
or U9640 (N_9640,N_6305,N_7737);
nor U9641 (N_9641,N_6048,N_6730);
xor U9642 (N_9642,N_6771,N_7006);
and U9643 (N_9643,N_6983,N_7966);
nor U9644 (N_9644,N_6361,N_7692);
and U9645 (N_9645,N_6772,N_6591);
or U9646 (N_9646,N_7182,N_6200);
nor U9647 (N_9647,N_6337,N_6682);
and U9648 (N_9648,N_7083,N_7033);
nand U9649 (N_9649,N_7525,N_6377);
and U9650 (N_9650,N_6118,N_6877);
xnor U9651 (N_9651,N_6448,N_6079);
nand U9652 (N_9652,N_7323,N_6864);
nand U9653 (N_9653,N_7858,N_6240);
nor U9654 (N_9654,N_7663,N_6677);
nor U9655 (N_9655,N_7033,N_7688);
nand U9656 (N_9656,N_6149,N_7158);
and U9657 (N_9657,N_7217,N_7129);
and U9658 (N_9658,N_6536,N_7511);
xnor U9659 (N_9659,N_6228,N_6032);
xnor U9660 (N_9660,N_6791,N_6972);
or U9661 (N_9661,N_6081,N_6719);
or U9662 (N_9662,N_7133,N_7144);
or U9663 (N_9663,N_7635,N_7055);
xnor U9664 (N_9664,N_6825,N_7551);
nor U9665 (N_9665,N_6183,N_6361);
xor U9666 (N_9666,N_6437,N_7476);
and U9667 (N_9667,N_6197,N_6793);
nand U9668 (N_9668,N_6683,N_7935);
nor U9669 (N_9669,N_7657,N_6738);
or U9670 (N_9670,N_6194,N_7303);
nor U9671 (N_9671,N_7713,N_7235);
or U9672 (N_9672,N_7047,N_6798);
nand U9673 (N_9673,N_7743,N_6825);
nor U9674 (N_9674,N_7397,N_6910);
or U9675 (N_9675,N_6526,N_6648);
nor U9676 (N_9676,N_7292,N_7274);
nor U9677 (N_9677,N_7634,N_6528);
nor U9678 (N_9678,N_7964,N_6836);
nand U9679 (N_9679,N_6445,N_7225);
or U9680 (N_9680,N_6954,N_6228);
or U9681 (N_9681,N_6159,N_6322);
nand U9682 (N_9682,N_7445,N_6788);
nand U9683 (N_9683,N_6838,N_6733);
nand U9684 (N_9684,N_7503,N_7142);
nor U9685 (N_9685,N_7155,N_7776);
and U9686 (N_9686,N_7220,N_7225);
nand U9687 (N_9687,N_7976,N_6621);
nor U9688 (N_9688,N_6521,N_6992);
nor U9689 (N_9689,N_6010,N_6699);
nor U9690 (N_9690,N_6523,N_6468);
nand U9691 (N_9691,N_7149,N_6590);
or U9692 (N_9692,N_7113,N_7419);
and U9693 (N_9693,N_6446,N_7596);
nor U9694 (N_9694,N_7804,N_7115);
nand U9695 (N_9695,N_7371,N_7184);
nand U9696 (N_9696,N_7043,N_7798);
and U9697 (N_9697,N_6058,N_7125);
nor U9698 (N_9698,N_6651,N_7854);
xor U9699 (N_9699,N_7935,N_6915);
or U9700 (N_9700,N_6649,N_6780);
or U9701 (N_9701,N_7123,N_6581);
nor U9702 (N_9702,N_6107,N_7556);
or U9703 (N_9703,N_7049,N_6826);
nand U9704 (N_9704,N_7812,N_6047);
nor U9705 (N_9705,N_6622,N_7321);
and U9706 (N_9706,N_7804,N_6798);
nand U9707 (N_9707,N_6547,N_6309);
nand U9708 (N_9708,N_6144,N_6346);
or U9709 (N_9709,N_6684,N_7204);
nand U9710 (N_9710,N_7230,N_7682);
and U9711 (N_9711,N_6197,N_6918);
nor U9712 (N_9712,N_7127,N_6328);
and U9713 (N_9713,N_7690,N_6414);
or U9714 (N_9714,N_7606,N_6604);
nand U9715 (N_9715,N_6423,N_6841);
xor U9716 (N_9716,N_7693,N_7200);
nand U9717 (N_9717,N_6266,N_6662);
xor U9718 (N_9718,N_7952,N_6577);
or U9719 (N_9719,N_6349,N_6316);
nand U9720 (N_9720,N_7200,N_6091);
and U9721 (N_9721,N_7289,N_6691);
and U9722 (N_9722,N_6698,N_7262);
nor U9723 (N_9723,N_6649,N_7212);
and U9724 (N_9724,N_7224,N_7164);
nor U9725 (N_9725,N_6477,N_7462);
and U9726 (N_9726,N_6171,N_7006);
nor U9727 (N_9727,N_6563,N_7903);
and U9728 (N_9728,N_7134,N_6371);
or U9729 (N_9729,N_6387,N_6432);
or U9730 (N_9730,N_7874,N_7571);
nand U9731 (N_9731,N_7364,N_6321);
xnor U9732 (N_9732,N_6182,N_6204);
and U9733 (N_9733,N_7784,N_6427);
nand U9734 (N_9734,N_7261,N_6149);
and U9735 (N_9735,N_6885,N_6365);
nand U9736 (N_9736,N_6849,N_6166);
xor U9737 (N_9737,N_7702,N_7992);
nand U9738 (N_9738,N_7020,N_7756);
nor U9739 (N_9739,N_7030,N_6246);
nand U9740 (N_9740,N_7756,N_7464);
nor U9741 (N_9741,N_7003,N_7526);
and U9742 (N_9742,N_6441,N_6855);
nor U9743 (N_9743,N_7132,N_7566);
and U9744 (N_9744,N_6091,N_7984);
nor U9745 (N_9745,N_7777,N_6918);
nand U9746 (N_9746,N_7140,N_6627);
and U9747 (N_9747,N_7524,N_7767);
nand U9748 (N_9748,N_7994,N_6468);
and U9749 (N_9749,N_6553,N_6079);
nor U9750 (N_9750,N_6489,N_6526);
nor U9751 (N_9751,N_7709,N_6623);
or U9752 (N_9752,N_7425,N_7744);
nor U9753 (N_9753,N_7308,N_6736);
xnor U9754 (N_9754,N_7612,N_6136);
and U9755 (N_9755,N_7667,N_6306);
or U9756 (N_9756,N_7785,N_6486);
nand U9757 (N_9757,N_7755,N_6279);
and U9758 (N_9758,N_7524,N_6484);
nand U9759 (N_9759,N_7469,N_7547);
nor U9760 (N_9760,N_6121,N_6266);
and U9761 (N_9761,N_7898,N_7189);
and U9762 (N_9762,N_6893,N_6824);
or U9763 (N_9763,N_6857,N_6173);
and U9764 (N_9764,N_7701,N_7853);
nor U9765 (N_9765,N_7512,N_6298);
or U9766 (N_9766,N_6988,N_7483);
and U9767 (N_9767,N_7887,N_7048);
and U9768 (N_9768,N_6362,N_6215);
or U9769 (N_9769,N_7312,N_7310);
nor U9770 (N_9770,N_6997,N_6038);
nor U9771 (N_9771,N_6998,N_7199);
nand U9772 (N_9772,N_6762,N_7916);
nor U9773 (N_9773,N_7472,N_6676);
nand U9774 (N_9774,N_7973,N_6747);
nand U9775 (N_9775,N_6227,N_7433);
and U9776 (N_9776,N_6664,N_7409);
nand U9777 (N_9777,N_7130,N_6892);
nor U9778 (N_9778,N_6541,N_7895);
nor U9779 (N_9779,N_6544,N_7928);
nand U9780 (N_9780,N_7305,N_6799);
and U9781 (N_9781,N_6781,N_7206);
and U9782 (N_9782,N_6910,N_7788);
nor U9783 (N_9783,N_6126,N_6983);
nand U9784 (N_9784,N_6987,N_7797);
xnor U9785 (N_9785,N_6692,N_6007);
and U9786 (N_9786,N_6692,N_6339);
xnor U9787 (N_9787,N_6631,N_7287);
nor U9788 (N_9788,N_7488,N_7732);
and U9789 (N_9789,N_7763,N_7846);
nand U9790 (N_9790,N_7457,N_6144);
and U9791 (N_9791,N_6147,N_7250);
or U9792 (N_9792,N_7142,N_7338);
and U9793 (N_9793,N_6676,N_6548);
xor U9794 (N_9794,N_6722,N_6381);
nor U9795 (N_9795,N_7846,N_6637);
xor U9796 (N_9796,N_6560,N_7655);
and U9797 (N_9797,N_7266,N_6733);
nor U9798 (N_9798,N_6303,N_6567);
nor U9799 (N_9799,N_7029,N_6816);
xnor U9800 (N_9800,N_7003,N_6304);
xor U9801 (N_9801,N_6192,N_6646);
and U9802 (N_9802,N_6851,N_6722);
xor U9803 (N_9803,N_7537,N_7481);
and U9804 (N_9804,N_7219,N_7562);
and U9805 (N_9805,N_6644,N_6327);
or U9806 (N_9806,N_6679,N_6356);
nand U9807 (N_9807,N_6649,N_6783);
and U9808 (N_9808,N_6390,N_6447);
and U9809 (N_9809,N_6906,N_7327);
nor U9810 (N_9810,N_6480,N_7074);
or U9811 (N_9811,N_7736,N_6033);
nand U9812 (N_9812,N_7604,N_7346);
xor U9813 (N_9813,N_6351,N_7658);
or U9814 (N_9814,N_7318,N_7600);
or U9815 (N_9815,N_6599,N_6775);
nor U9816 (N_9816,N_7271,N_6882);
or U9817 (N_9817,N_6781,N_7344);
xnor U9818 (N_9818,N_6260,N_7757);
nor U9819 (N_9819,N_7193,N_7020);
or U9820 (N_9820,N_7460,N_6598);
nand U9821 (N_9821,N_7820,N_6764);
or U9822 (N_9822,N_6541,N_7694);
or U9823 (N_9823,N_6868,N_6644);
and U9824 (N_9824,N_6399,N_7290);
nor U9825 (N_9825,N_7369,N_6389);
nor U9826 (N_9826,N_6957,N_6880);
or U9827 (N_9827,N_6701,N_7268);
and U9828 (N_9828,N_6475,N_6178);
nand U9829 (N_9829,N_7246,N_7489);
and U9830 (N_9830,N_6190,N_6399);
xnor U9831 (N_9831,N_6449,N_7257);
or U9832 (N_9832,N_6419,N_7717);
nand U9833 (N_9833,N_7880,N_7803);
xnor U9834 (N_9834,N_6426,N_6679);
or U9835 (N_9835,N_6404,N_7101);
nand U9836 (N_9836,N_7049,N_6711);
nand U9837 (N_9837,N_7720,N_7983);
nor U9838 (N_9838,N_6947,N_7517);
and U9839 (N_9839,N_6580,N_7907);
nor U9840 (N_9840,N_6476,N_7259);
or U9841 (N_9841,N_6284,N_7399);
or U9842 (N_9842,N_6907,N_7820);
or U9843 (N_9843,N_6196,N_6776);
nand U9844 (N_9844,N_7416,N_6242);
nand U9845 (N_9845,N_6877,N_7111);
or U9846 (N_9846,N_6932,N_7782);
nor U9847 (N_9847,N_7133,N_6470);
nand U9848 (N_9848,N_7186,N_6178);
xor U9849 (N_9849,N_7799,N_7686);
nor U9850 (N_9850,N_7036,N_6892);
or U9851 (N_9851,N_6442,N_7820);
and U9852 (N_9852,N_7216,N_7214);
or U9853 (N_9853,N_7824,N_6486);
nor U9854 (N_9854,N_6578,N_7822);
nand U9855 (N_9855,N_7424,N_7018);
nand U9856 (N_9856,N_7839,N_6700);
nand U9857 (N_9857,N_6577,N_7290);
and U9858 (N_9858,N_6261,N_7000);
nor U9859 (N_9859,N_6175,N_7908);
or U9860 (N_9860,N_7600,N_7311);
nor U9861 (N_9861,N_6043,N_7836);
nor U9862 (N_9862,N_6857,N_7366);
nor U9863 (N_9863,N_7183,N_6244);
nor U9864 (N_9864,N_7689,N_7494);
xnor U9865 (N_9865,N_6284,N_6586);
and U9866 (N_9866,N_6562,N_7399);
nor U9867 (N_9867,N_7014,N_6834);
or U9868 (N_9868,N_7007,N_7686);
nand U9869 (N_9869,N_7256,N_6152);
nor U9870 (N_9870,N_7017,N_7623);
nor U9871 (N_9871,N_7248,N_7310);
and U9872 (N_9872,N_6253,N_6074);
or U9873 (N_9873,N_6025,N_6101);
xnor U9874 (N_9874,N_7932,N_7845);
xnor U9875 (N_9875,N_6939,N_6533);
nand U9876 (N_9876,N_7466,N_7177);
and U9877 (N_9877,N_6071,N_7393);
nor U9878 (N_9878,N_7332,N_7251);
or U9879 (N_9879,N_7535,N_6633);
nand U9880 (N_9880,N_7283,N_7710);
and U9881 (N_9881,N_6715,N_7283);
or U9882 (N_9882,N_6241,N_6790);
or U9883 (N_9883,N_6395,N_6273);
nor U9884 (N_9884,N_7201,N_7162);
or U9885 (N_9885,N_7042,N_7950);
nor U9886 (N_9886,N_6223,N_6184);
and U9887 (N_9887,N_6790,N_7683);
and U9888 (N_9888,N_6609,N_7751);
nand U9889 (N_9889,N_7279,N_7500);
and U9890 (N_9890,N_7550,N_7489);
and U9891 (N_9891,N_7574,N_6918);
nand U9892 (N_9892,N_6793,N_6648);
nand U9893 (N_9893,N_6300,N_7175);
nor U9894 (N_9894,N_7846,N_6337);
or U9895 (N_9895,N_6315,N_6647);
and U9896 (N_9896,N_7519,N_7374);
nand U9897 (N_9897,N_6569,N_6870);
xor U9898 (N_9898,N_7781,N_6064);
or U9899 (N_9899,N_7226,N_6853);
nand U9900 (N_9900,N_6899,N_6655);
nand U9901 (N_9901,N_6303,N_7342);
and U9902 (N_9902,N_6687,N_7558);
xnor U9903 (N_9903,N_7112,N_6929);
nand U9904 (N_9904,N_6405,N_7147);
or U9905 (N_9905,N_6396,N_7822);
nand U9906 (N_9906,N_6063,N_7823);
and U9907 (N_9907,N_6107,N_6053);
or U9908 (N_9908,N_7873,N_6794);
or U9909 (N_9909,N_7027,N_6210);
and U9910 (N_9910,N_6060,N_7345);
and U9911 (N_9911,N_7855,N_6427);
nand U9912 (N_9912,N_6064,N_7667);
nor U9913 (N_9913,N_7481,N_6950);
and U9914 (N_9914,N_7544,N_7660);
nor U9915 (N_9915,N_6095,N_7827);
or U9916 (N_9916,N_7130,N_7954);
and U9917 (N_9917,N_6157,N_6951);
nor U9918 (N_9918,N_7516,N_7958);
nor U9919 (N_9919,N_6753,N_6381);
nor U9920 (N_9920,N_6359,N_7147);
and U9921 (N_9921,N_6625,N_7873);
nor U9922 (N_9922,N_6580,N_7758);
nand U9923 (N_9923,N_7004,N_6846);
nand U9924 (N_9924,N_6590,N_6683);
nand U9925 (N_9925,N_6230,N_6813);
or U9926 (N_9926,N_7553,N_7581);
nor U9927 (N_9927,N_7553,N_6481);
nor U9928 (N_9928,N_6051,N_7317);
nand U9929 (N_9929,N_7269,N_6245);
or U9930 (N_9930,N_7655,N_6594);
xnor U9931 (N_9931,N_7236,N_6429);
nor U9932 (N_9932,N_7483,N_7165);
nand U9933 (N_9933,N_7077,N_6094);
or U9934 (N_9934,N_6984,N_7844);
nand U9935 (N_9935,N_6727,N_7276);
or U9936 (N_9936,N_7814,N_6937);
nand U9937 (N_9937,N_6712,N_6499);
or U9938 (N_9938,N_6662,N_6315);
or U9939 (N_9939,N_6377,N_6554);
or U9940 (N_9940,N_7784,N_6208);
and U9941 (N_9941,N_6217,N_7925);
nor U9942 (N_9942,N_7851,N_7925);
xnor U9943 (N_9943,N_7191,N_6246);
or U9944 (N_9944,N_6223,N_7809);
or U9945 (N_9945,N_6582,N_7492);
and U9946 (N_9946,N_6165,N_6460);
or U9947 (N_9947,N_6271,N_6329);
or U9948 (N_9948,N_7990,N_7012);
and U9949 (N_9949,N_7768,N_6198);
nor U9950 (N_9950,N_7851,N_6741);
and U9951 (N_9951,N_6460,N_7187);
and U9952 (N_9952,N_7692,N_7961);
nand U9953 (N_9953,N_6798,N_7330);
nor U9954 (N_9954,N_6845,N_6699);
nor U9955 (N_9955,N_7289,N_7142);
nand U9956 (N_9956,N_7934,N_6046);
nand U9957 (N_9957,N_6191,N_6702);
xnor U9958 (N_9958,N_6421,N_7672);
and U9959 (N_9959,N_7297,N_6554);
or U9960 (N_9960,N_6155,N_7477);
or U9961 (N_9961,N_7542,N_6892);
xor U9962 (N_9962,N_7038,N_6763);
and U9963 (N_9963,N_7329,N_7809);
and U9964 (N_9964,N_6316,N_7147);
nor U9965 (N_9965,N_6638,N_7814);
or U9966 (N_9966,N_7947,N_7686);
or U9967 (N_9967,N_7553,N_6923);
or U9968 (N_9968,N_7021,N_7378);
nand U9969 (N_9969,N_6548,N_7265);
xnor U9970 (N_9970,N_7056,N_7448);
or U9971 (N_9971,N_7927,N_6187);
nand U9972 (N_9972,N_6808,N_7572);
nor U9973 (N_9973,N_7743,N_7598);
xnor U9974 (N_9974,N_7361,N_7574);
nand U9975 (N_9975,N_6131,N_6383);
nand U9976 (N_9976,N_7452,N_6020);
or U9977 (N_9977,N_6780,N_7782);
or U9978 (N_9978,N_6576,N_7003);
or U9979 (N_9979,N_7292,N_7121);
nor U9980 (N_9980,N_6014,N_6256);
xor U9981 (N_9981,N_6389,N_7937);
nor U9982 (N_9982,N_6941,N_7807);
and U9983 (N_9983,N_7681,N_6597);
and U9984 (N_9984,N_6859,N_6754);
nor U9985 (N_9985,N_7170,N_7767);
and U9986 (N_9986,N_6507,N_7244);
and U9987 (N_9987,N_7071,N_6126);
nor U9988 (N_9988,N_7804,N_6934);
or U9989 (N_9989,N_6583,N_6580);
and U9990 (N_9990,N_7495,N_6890);
or U9991 (N_9991,N_6407,N_7878);
nor U9992 (N_9992,N_7497,N_7179);
or U9993 (N_9993,N_7657,N_7543);
and U9994 (N_9994,N_7163,N_6763);
nand U9995 (N_9995,N_6575,N_6142);
nand U9996 (N_9996,N_6215,N_7430);
or U9997 (N_9997,N_6240,N_7921);
nand U9998 (N_9998,N_6450,N_6853);
or U9999 (N_9999,N_6113,N_7330);
nor U10000 (N_10000,N_8517,N_9977);
nand U10001 (N_10001,N_9883,N_8055);
or U10002 (N_10002,N_9012,N_8939);
nor U10003 (N_10003,N_9241,N_8071);
and U10004 (N_10004,N_8361,N_9824);
nand U10005 (N_10005,N_8786,N_9268);
and U10006 (N_10006,N_8058,N_8293);
nor U10007 (N_10007,N_9590,N_9013);
nand U10008 (N_10008,N_9661,N_8697);
or U10009 (N_10009,N_8513,N_8835);
and U10010 (N_10010,N_8890,N_9705);
nand U10011 (N_10011,N_9058,N_9935);
nor U10012 (N_10012,N_9919,N_9166);
or U10013 (N_10013,N_8986,N_8043);
and U10014 (N_10014,N_8026,N_9965);
xnor U10015 (N_10015,N_8805,N_9487);
and U10016 (N_10016,N_8905,N_8593);
and U10017 (N_10017,N_8191,N_8996);
nor U10018 (N_10018,N_8719,N_8211);
and U10019 (N_10019,N_8139,N_9257);
nor U10020 (N_10020,N_9776,N_8725);
nor U10021 (N_10021,N_8377,N_8126);
nand U10022 (N_10022,N_8568,N_8016);
and U10023 (N_10023,N_9056,N_8448);
nor U10024 (N_10024,N_8999,N_8707);
or U10025 (N_10025,N_9360,N_8751);
and U10026 (N_10026,N_9679,N_9745);
nand U10027 (N_10027,N_8898,N_9107);
nand U10028 (N_10028,N_8021,N_8532);
nand U10029 (N_10029,N_9535,N_8418);
nor U10030 (N_10030,N_8265,N_8533);
nor U10031 (N_10031,N_9081,N_9893);
nor U10032 (N_10032,N_8475,N_9850);
or U10033 (N_10033,N_8772,N_8696);
nand U10034 (N_10034,N_9711,N_8792);
and U10035 (N_10035,N_8557,N_8888);
xnor U10036 (N_10036,N_9440,N_9310);
nor U10037 (N_10037,N_9186,N_8777);
or U10038 (N_10038,N_8953,N_8443);
nand U10039 (N_10039,N_8669,N_9640);
nor U10040 (N_10040,N_8711,N_9109);
nand U10041 (N_10041,N_8171,N_8665);
or U10042 (N_10042,N_9915,N_9903);
nand U10043 (N_10043,N_9164,N_8210);
or U10044 (N_10044,N_8076,N_8865);
nor U10045 (N_10045,N_8342,N_8882);
nand U10046 (N_10046,N_9236,N_9541);
nor U10047 (N_10047,N_9272,N_8470);
nor U10048 (N_10048,N_9414,N_8226);
nor U10049 (N_10049,N_9890,N_9742);
nand U10050 (N_10050,N_9486,N_8212);
nand U10051 (N_10051,N_8339,N_9635);
nand U10052 (N_10052,N_9714,N_8881);
xnor U10053 (N_10053,N_8009,N_8545);
nand U10054 (N_10054,N_8283,N_8761);
xnor U10055 (N_10055,N_9558,N_9083);
nand U10056 (N_10056,N_9826,N_9697);
or U10057 (N_10057,N_8052,N_8927);
nor U10058 (N_10058,N_9684,N_9871);
and U10059 (N_10059,N_9933,N_8901);
nand U10060 (N_10060,N_9877,N_9709);
or U10061 (N_10061,N_9490,N_9795);
nor U10062 (N_10062,N_9142,N_8404);
nand U10063 (N_10063,N_8810,N_8619);
or U10064 (N_10064,N_9418,N_8208);
or U10065 (N_10065,N_9671,N_9458);
nand U10066 (N_10066,N_8731,N_8934);
nand U10067 (N_10067,N_9219,N_8913);
and U10068 (N_10068,N_9253,N_9327);
and U10069 (N_10069,N_8841,N_8040);
and U10070 (N_10070,N_9544,N_8940);
or U10071 (N_10071,N_9296,N_9834);
or U10072 (N_10072,N_9454,N_9402);
nand U10073 (N_10073,N_8842,N_9996);
nand U10074 (N_10074,N_8263,N_9080);
xnor U10075 (N_10075,N_8623,N_8867);
or U10076 (N_10076,N_8600,N_8575);
and U10077 (N_10077,N_9303,N_8896);
and U10078 (N_10078,N_9318,N_9617);
nor U10079 (N_10079,N_8745,N_8015);
or U10080 (N_10080,N_9921,N_9605);
or U10081 (N_10081,N_9132,N_8409);
or U10082 (N_10082,N_8196,N_9752);
or U10083 (N_10083,N_8231,N_8322);
nor U10084 (N_10084,N_9026,N_8968);
and U10085 (N_10085,N_9780,N_9434);
xnor U10086 (N_10086,N_9961,N_8233);
nand U10087 (N_10087,N_8437,N_9678);
nand U10088 (N_10088,N_8203,N_8702);
or U10089 (N_10089,N_9329,N_9404);
or U10090 (N_10090,N_8776,N_8417);
or U10091 (N_10091,N_9810,N_8426);
nor U10092 (N_10092,N_9205,N_8118);
or U10093 (N_10093,N_8518,N_8672);
nor U10094 (N_10094,N_9455,N_9920);
nand U10095 (N_10095,N_8523,N_8874);
nor U10096 (N_10096,N_9460,N_9981);
xnor U10097 (N_10097,N_9265,N_9672);
nor U10098 (N_10098,N_9974,N_9527);
nor U10099 (N_10099,N_9021,N_9027);
or U10100 (N_10100,N_9014,N_8784);
or U10101 (N_10101,N_8060,N_8949);
nand U10102 (N_10102,N_8027,N_9529);
xor U10103 (N_10103,N_9726,N_9936);
nor U10104 (N_10104,N_9702,N_9170);
or U10105 (N_10105,N_8394,N_9207);
or U10106 (N_10106,N_8232,N_8067);
nor U10107 (N_10107,N_9075,N_9592);
and U10108 (N_10108,N_8657,N_8400);
or U10109 (N_10109,N_8936,N_9522);
or U10110 (N_10110,N_8507,N_8257);
and U10111 (N_10111,N_8825,N_9868);
or U10112 (N_10112,N_9339,N_9864);
nand U10113 (N_10113,N_8062,N_9577);
nor U10114 (N_10114,N_9422,N_8157);
or U10115 (N_10115,N_9478,N_9618);
or U10116 (N_10116,N_9949,N_9894);
and U10117 (N_10117,N_9502,N_9523);
and U10118 (N_10118,N_9498,N_9719);
nor U10119 (N_10119,N_9284,N_8013);
xor U10120 (N_10120,N_9182,N_9861);
nor U10121 (N_10121,N_9149,N_8973);
nor U10122 (N_10122,N_9252,N_9950);
and U10123 (N_10123,N_9772,N_8469);
or U10124 (N_10124,N_8651,N_8753);
xor U10125 (N_10125,N_8634,N_8240);
and U10126 (N_10126,N_8308,N_8893);
and U10127 (N_10127,N_8653,N_8102);
nand U10128 (N_10128,N_8829,N_9443);
and U10129 (N_10129,N_8563,N_8401);
nand U10130 (N_10130,N_9054,N_8597);
or U10131 (N_10131,N_8030,N_9090);
or U10132 (N_10132,N_8536,N_9195);
or U10133 (N_10133,N_8285,N_9395);
nor U10134 (N_10134,N_8559,N_8538);
nand U10135 (N_10135,N_9214,N_9016);
xnor U10136 (N_10136,N_8641,N_9762);
or U10137 (N_10137,N_8444,N_9585);
and U10138 (N_10138,N_8331,N_8904);
and U10139 (N_10139,N_9568,N_8595);
or U10140 (N_10140,N_9774,N_9153);
and U10141 (N_10141,N_8886,N_8353);
or U10142 (N_10142,N_8255,N_8323);
and U10143 (N_10143,N_8442,N_9168);
or U10144 (N_10144,N_9701,N_8587);
nor U10145 (N_10145,N_8204,N_9955);
nand U10146 (N_10146,N_8245,N_8480);
or U10147 (N_10147,N_8650,N_8247);
or U10148 (N_10148,N_9198,N_8175);
xor U10149 (N_10149,N_8094,N_8637);
nand U10150 (N_10150,N_8487,N_8386);
nor U10151 (N_10151,N_8039,N_9513);
or U10152 (N_10152,N_8664,N_8078);
nand U10153 (N_10153,N_8717,N_8716);
or U10154 (N_10154,N_9368,N_8797);
and U10155 (N_10155,N_8820,N_9097);
nand U10156 (N_10156,N_8856,N_8161);
nor U10157 (N_10157,N_9687,N_9552);
and U10158 (N_10158,N_9157,N_9971);
and U10159 (N_10159,N_8111,N_9900);
or U10160 (N_10160,N_8685,N_9707);
nand U10161 (N_10161,N_9408,N_9323);
or U10162 (N_10162,N_9743,N_9658);
and U10163 (N_10163,N_8980,N_9730);
or U10164 (N_10164,N_8579,N_9231);
and U10165 (N_10165,N_8847,N_8871);
nand U10166 (N_10166,N_8954,N_9613);
xnor U10167 (N_10167,N_9620,N_8352);
nand U10168 (N_10168,N_9147,N_9542);
or U10169 (N_10169,N_9956,N_8433);
and U10170 (N_10170,N_9922,N_8580);
nand U10171 (N_10171,N_9556,N_8767);
nand U10172 (N_10172,N_8370,N_9423);
or U10173 (N_10173,N_8628,N_8214);
nand U10174 (N_10174,N_9447,N_8195);
nor U10175 (N_10175,N_8237,N_9904);
nor U10176 (N_10176,N_8423,N_8970);
or U10177 (N_10177,N_8610,N_8284);
nand U10178 (N_10178,N_9654,N_8706);
nand U10179 (N_10179,N_8670,N_8676);
nor U10180 (N_10180,N_9003,N_9212);
nor U10181 (N_10181,N_9341,N_9326);
and U10182 (N_10182,N_8429,N_8193);
or U10183 (N_10183,N_8292,N_8351);
nand U10184 (N_10184,N_8704,N_9985);
nand U10185 (N_10185,N_9593,N_8506);
nand U10186 (N_10186,N_9173,N_9695);
nand U10187 (N_10187,N_9238,N_8962);
or U10188 (N_10188,N_8833,N_8128);
nor U10189 (N_10189,N_8186,N_8425);
xnor U10190 (N_10190,N_9316,N_9029);
nand U10191 (N_10191,N_8919,N_8019);
nand U10192 (N_10192,N_9619,N_9978);
xor U10193 (N_10193,N_8367,N_9350);
nand U10194 (N_10194,N_9136,N_8083);
nand U10195 (N_10195,N_9713,N_9138);
xnor U10196 (N_10196,N_9218,N_8066);
and U10197 (N_10197,N_8383,N_8051);
and U10198 (N_10198,N_9706,N_9918);
xnor U10199 (N_10199,N_8869,N_8050);
nor U10200 (N_10200,N_9943,N_8047);
nor U10201 (N_10201,N_9397,N_8491);
nand U10202 (N_10202,N_9839,N_8560);
or U10203 (N_10203,N_9913,N_9651);
or U10204 (N_10204,N_8243,N_8655);
or U10205 (N_10205,N_9939,N_9446);
nor U10206 (N_10206,N_9616,N_9492);
or U10207 (N_10207,N_8765,N_8345);
xor U10208 (N_10208,N_9419,N_9531);
and U10209 (N_10209,N_8248,N_8177);
and U10210 (N_10210,N_8605,N_9823);
or U10211 (N_10211,N_9636,N_9482);
nor U10212 (N_10212,N_9938,N_9103);
nand U10213 (N_10213,N_9597,N_9630);
nor U10214 (N_10214,N_8509,N_9425);
and U10215 (N_10215,N_9537,N_9859);
or U10216 (N_10216,N_8638,N_9982);
nand U10217 (N_10217,N_8234,N_9840);
and U10218 (N_10218,N_9767,N_8863);
and U10219 (N_10219,N_9735,N_8092);
or U10220 (N_10220,N_8618,N_9332);
or U10221 (N_10221,N_8160,N_9139);
or U10222 (N_10222,N_9548,N_8225);
or U10223 (N_10223,N_8581,N_8416);
or U10224 (N_10224,N_9245,N_8872);
xnor U10225 (N_10225,N_8159,N_8238);
nand U10226 (N_10226,N_8611,N_8471);
nand U10227 (N_10227,N_9660,N_9234);
or U10228 (N_10228,N_8291,N_9357);
nand U10229 (N_10229,N_8504,N_8853);
xor U10230 (N_10230,N_9145,N_8920);
and U10231 (N_10231,N_9728,N_8304);
and U10232 (N_10232,N_8564,N_8633);
and U10233 (N_10233,N_9633,N_9768);
or U10234 (N_10234,N_9427,N_9604);
nand U10235 (N_10235,N_8995,N_9647);
and U10236 (N_10236,N_9753,N_9033);
or U10237 (N_10237,N_9415,N_9587);
and U10238 (N_10238,N_8671,N_8677);
and U10239 (N_10239,N_8174,N_9063);
or U10240 (N_10240,N_8566,N_9184);
nand U10241 (N_10241,N_8516,N_9483);
or U10242 (N_10242,N_9034,N_8802);
or U10243 (N_10243,N_9472,N_9453);
nor U10244 (N_10244,N_8738,N_8493);
or U10245 (N_10245,N_9748,N_8885);
and U10246 (N_10246,N_9030,N_9691);
xnor U10247 (N_10247,N_8054,N_8101);
nand U10248 (N_10248,N_8862,N_8024);
and U10249 (N_10249,N_8911,N_9865);
nor U10250 (N_10250,N_9796,N_9409);
and U10251 (N_10251,N_8222,N_8866);
or U10252 (N_10252,N_8722,N_8957);
nor U10253 (N_10253,N_9641,N_8680);
nor U10254 (N_10254,N_8360,N_9369);
nor U10255 (N_10255,N_8945,N_8737);
and U10256 (N_10256,N_9320,N_9151);
nand U10257 (N_10257,N_8870,N_9039);
nor U10258 (N_10258,N_9375,N_9724);
nand U10259 (N_10259,N_9932,N_8125);
nor U10260 (N_10260,N_9174,N_8556);
nor U10261 (N_10261,N_9424,N_8314);
or U10262 (N_10262,N_8044,N_9226);
and U10263 (N_10263,N_9525,N_8355);
nand U10264 (N_10264,N_9200,N_8381);
nand U10265 (N_10265,N_9511,N_9037);
xnor U10266 (N_10266,N_8780,N_8084);
nor U10267 (N_10267,N_9740,N_8700);
or U10268 (N_10268,N_8264,N_9099);
or U10269 (N_10269,N_8917,N_8915);
and U10270 (N_10270,N_8456,N_8428);
or U10271 (N_10271,N_9833,N_9975);
nor U10272 (N_10272,N_8310,N_8730);
nor U10273 (N_10273,N_9420,N_8288);
or U10274 (N_10274,N_8733,N_8976);
or U10275 (N_10275,N_8964,N_8972);
or U10276 (N_10276,N_9479,N_9550);
and U10277 (N_10277,N_9031,N_8815);
nand U10278 (N_10278,N_9841,N_8816);
and U10279 (N_10279,N_8809,N_8807);
and U10280 (N_10280,N_8567,N_8951);
and U10281 (N_10281,N_9615,N_8769);
and U10282 (N_10282,N_9637,N_8586);
nor U10283 (N_10283,N_9264,N_8817);
nor U10284 (N_10284,N_9074,N_9297);
nor U10285 (N_10285,N_8096,N_9644);
or U10286 (N_10286,N_9575,N_9643);
and U10287 (N_10287,N_9129,N_8287);
nor U10288 (N_10288,N_9788,N_8689);
nand U10289 (N_10289,N_9266,N_8390);
or U10290 (N_10290,N_9197,N_8526);
xnor U10291 (N_10291,N_9787,N_9158);
nor U10292 (N_10292,N_9650,N_8585);
nand U10293 (N_10293,N_9820,N_8132);
nor U10294 (N_10294,N_8889,N_9244);
or U10295 (N_10295,N_8299,N_9314);
and U10296 (N_10296,N_8260,N_9869);
xnor U10297 (N_10297,N_8325,N_9295);
nor U10298 (N_10298,N_8346,N_8192);
or U10299 (N_10299,N_8230,N_9354);
nor U10300 (N_10300,N_9779,N_8252);
and U10301 (N_10301,N_8691,N_8740);
xor U10302 (N_10302,N_9716,N_9829);
or U10303 (N_10303,N_9927,N_8749);
or U10304 (N_10304,N_9143,N_9925);
nand U10305 (N_10305,N_9049,N_9271);
nand U10306 (N_10306,N_8682,N_8553);
xnor U10307 (N_10307,N_9838,N_8821);
nand U10308 (N_10308,N_9516,N_8005);
nand U10309 (N_10309,N_9905,N_9737);
and U10310 (N_10310,N_8178,N_8693);
and U10311 (N_10311,N_9010,N_8922);
and U10312 (N_10312,N_8363,N_9946);
and U10313 (N_10313,N_8460,N_9328);
and U10314 (N_10314,N_8166,N_8768);
nand U10315 (N_10315,N_8272,N_8205);
nor U10316 (N_10316,N_8492,N_9365);
or U10317 (N_10317,N_8850,N_8793);
or U10318 (N_10318,N_8681,N_8510);
and U10319 (N_10319,N_9335,N_8495);
and U10320 (N_10320,N_9642,N_9356);
or U10321 (N_10321,N_9791,N_9766);
nor U10322 (N_10322,N_9972,N_9689);
nand U10323 (N_10323,N_8975,N_9108);
and U10324 (N_10324,N_9330,N_8511);
nor U10325 (N_10325,N_9607,N_9007);
or U10326 (N_10326,N_8754,N_8661);
or U10327 (N_10327,N_8946,N_9225);
nand U10328 (N_10328,N_9761,N_9601);
and U10329 (N_10329,N_8406,N_8474);
nand U10330 (N_10330,N_9065,N_9183);
nand U10331 (N_10331,N_8534,N_8734);
xor U10332 (N_10332,N_9622,N_9112);
or U10333 (N_10333,N_8337,N_9872);
nor U10334 (N_10334,N_8858,N_9733);
nand U10335 (N_10335,N_8399,N_8061);
and U10336 (N_10336,N_8723,N_9847);
nand U10337 (N_10337,N_8008,N_9576);
xor U10338 (N_10338,N_9237,N_8228);
xor U10339 (N_10339,N_8430,N_8588);
or U10340 (N_10340,N_8183,N_9690);
or U10341 (N_10341,N_9555,N_9130);
nor U10342 (N_10342,N_8535,N_9283);
or U10343 (N_10343,N_9390,N_8714);
or U10344 (N_10344,N_8663,N_8328);
nor U10345 (N_10345,N_8584,N_9385);
or U10346 (N_10346,N_9072,N_8989);
xnor U10347 (N_10347,N_8830,N_9276);
xor U10348 (N_10348,N_9274,N_8421);
nor U10349 (N_10349,N_8712,N_8477);
nand U10350 (N_10350,N_9148,N_9624);
nand U10351 (N_10351,N_8781,N_9493);
and U10352 (N_10352,N_9193,N_9746);
or U10353 (N_10353,N_8883,N_9463);
or U10354 (N_10354,N_9710,N_9573);
nor U10355 (N_10355,N_9775,N_9570);
xor U10356 (N_10356,N_8846,N_9583);
nand U10357 (N_10357,N_9300,N_9888);
nor U10358 (N_10358,N_8840,N_9902);
xor U10359 (N_10359,N_8209,N_9722);
and U10360 (N_10360,N_8652,N_9125);
xor U10361 (N_10361,N_8223,N_8916);
xor U10362 (N_10362,N_9852,N_9095);
nand U10363 (N_10363,N_9403,N_8539);
and U10364 (N_10364,N_9958,N_8899);
nor U10365 (N_10365,N_9608,N_8379);
and U10366 (N_10366,N_8318,N_8281);
nor U10367 (N_10367,N_9988,N_9844);
xor U10368 (N_10368,N_9387,N_8290);
or U10369 (N_10369,N_8582,N_8461);
and U10370 (N_10370,N_9969,N_9798);
and U10371 (N_10371,N_9700,N_9569);
nor U10372 (N_10372,N_8640,N_9298);
nand U10373 (N_10373,N_8145,N_9180);
nand U10374 (N_10374,N_8392,N_9386);
and U10375 (N_10375,N_8709,N_9634);
nand U10376 (N_10376,N_8845,N_8113);
nand U10377 (N_10377,N_9771,N_9606);
nand U10378 (N_10378,N_9289,N_9751);
and U10379 (N_10379,N_8750,N_9800);
nand U10380 (N_10380,N_9190,N_9367);
or U10381 (N_10381,N_8366,N_8520);
nand U10382 (N_10382,N_8977,N_9038);
or U10383 (N_10383,N_8427,N_8718);
and U10384 (N_10384,N_8608,N_8958);
nor U10385 (N_10385,N_8020,N_9028);
nand U10386 (N_10386,N_8173,N_9040);
nand U10387 (N_10387,N_8530,N_9596);
nand U10388 (N_10388,N_8525,N_9464);
and U10389 (N_10389,N_8278,N_8077);
nor U10390 (N_10390,N_9579,N_9741);
nand U10391 (N_10391,N_9876,N_9382);
or U10392 (N_10392,N_8578,N_8490);
nor U10393 (N_10393,N_8082,N_8453);
or U10394 (N_10394,N_8546,N_9293);
nand U10395 (N_10395,N_9947,N_8446);
nand U10396 (N_10396,N_8544,N_8993);
or U10397 (N_10397,N_9122,N_9078);
nor U10398 (N_10398,N_8667,N_8298);
or U10399 (N_10399,N_9046,N_9662);
and U10400 (N_10400,N_8569,N_9322);
or U10401 (N_10401,N_8868,N_8974);
nor U10402 (N_10402,N_9822,N_8624);
or U10403 (N_10403,N_8818,N_9441);
and U10404 (N_10404,N_8771,N_8674);
nor U10405 (N_10405,N_9280,N_8197);
nand U10406 (N_10406,N_8375,N_8476);
nor U10407 (N_10407,N_8744,N_8554);
nor U10408 (N_10408,N_8317,N_9094);
xnor U10409 (N_10409,N_9782,N_8464);
nor U10410 (N_10410,N_9899,N_8952);
or U10411 (N_10411,N_9694,N_9067);
nor U10412 (N_10412,N_8478,N_9851);
nor U10413 (N_10413,N_8282,N_8056);
nand U10414 (N_10414,N_9827,N_8130);
or U10415 (N_10415,N_8775,N_9413);
or U10416 (N_10416,N_8053,N_9417);
and U10417 (N_10417,N_9685,N_8727);
nand U10418 (N_10418,N_8256,N_8496);
and U10419 (N_10419,N_9892,N_8267);
or U10420 (N_10420,N_8156,N_9290);
and U10421 (N_10421,N_9832,N_9020);
xnor U10422 (N_10422,N_9683,N_8741);
or U10423 (N_10423,N_8782,N_9421);
nand U10424 (N_10424,N_8926,N_8420);
or U10425 (N_10425,N_8755,N_9345);
nand U10426 (N_10426,N_8108,N_9885);
nor U10427 (N_10427,N_9581,N_8105);
and U10428 (N_10428,N_8275,N_9308);
or U10429 (N_10429,N_9944,N_8449);
and U10430 (N_10430,N_9632,N_9344);
or U10431 (N_10431,N_8826,N_9061);
and U10432 (N_10432,N_9187,N_8978);
nand U10433 (N_10433,N_8022,N_8087);
nand U10434 (N_10434,N_8774,N_9018);
nor U10435 (N_10435,N_8176,N_8621);
and U10436 (N_10436,N_9305,N_8218);
and U10437 (N_10437,N_8348,N_8612);
nor U10438 (N_10438,N_8499,N_8153);
and U10439 (N_10439,N_9064,N_9873);
or U10440 (N_10440,N_8937,N_8435);
and U10441 (N_10441,N_9519,N_9278);
nor U10442 (N_10442,N_9096,N_8302);
nor U10443 (N_10443,N_8457,N_8785);
nor U10444 (N_10444,N_8141,N_8316);
or U10445 (N_10445,N_8614,N_9396);
and U10446 (N_10446,N_8037,N_8341);
xor U10447 (N_10447,N_8286,N_8935);
or U10448 (N_10448,N_9708,N_9987);
nand U10449 (N_10449,N_9496,N_9477);
or U10450 (N_10450,N_9334,N_9625);
or U10451 (N_10451,N_9858,N_9549);
or U10452 (N_10452,N_8971,N_9261);
xor U10453 (N_10453,N_8903,N_8154);
nor U10454 (N_10454,N_8541,N_9884);
nand U10455 (N_10455,N_8531,N_9783);
or U10456 (N_10456,N_8242,N_9860);
or U10457 (N_10457,N_9998,N_8017);
and U10458 (N_10458,N_8187,N_9085);
nand U10459 (N_10459,N_8548,N_8127);
xnor U10460 (N_10460,N_8837,N_8168);
and U10461 (N_10461,N_8873,N_8405);
and U10462 (N_10462,N_9870,N_8790);
or U10463 (N_10463,N_8594,N_8198);
or U10464 (N_10464,N_9718,N_8274);
and U10465 (N_10465,N_9562,N_9591);
or U10466 (N_10466,N_8483,N_8362);
nor U10467 (N_10467,N_9343,N_8190);
or U10468 (N_10468,N_8194,N_8894);
xor U10469 (N_10469,N_9437,N_8961);
or U10470 (N_10470,N_8982,N_9828);
xnor U10471 (N_10471,N_9319,N_9243);
nand U10472 (N_10472,N_8148,N_9135);
xnor U10473 (N_10473,N_8129,N_9259);
nand U10474 (N_10474,N_8142,N_9698);
nor U10475 (N_10475,N_8167,N_9373);
nor U10476 (N_10476,N_8800,N_9349);
nand U10477 (N_10477,N_8227,N_9115);
nor U10478 (N_10478,N_9355,N_9156);
nor U10479 (N_10479,N_8431,N_9940);
or U10480 (N_10480,N_9843,N_9286);
and U10481 (N_10481,N_8956,N_9948);
and U10482 (N_10482,N_9821,N_8606);
nor U10483 (N_10483,N_8561,N_8715);
and U10484 (N_10484,N_9429,N_8997);
xor U10485 (N_10485,N_9517,N_8859);
xnor U10486 (N_10486,N_8002,N_9154);
and U10487 (N_10487,N_8938,N_8397);
or U10488 (N_10488,N_9267,N_9250);
nand U10489 (N_10489,N_9655,N_9663);
and U10490 (N_10490,N_9279,N_8415);
nor U10491 (N_10491,N_9564,N_9845);
nor U10492 (N_10492,N_9008,N_8296);
nor U10493 (N_10493,N_9169,N_9676);
and U10494 (N_10494,N_9491,N_8412);
nor U10495 (N_10495,N_9374,N_8468);
nand U10496 (N_10496,N_9227,N_9677);
or U10497 (N_10497,N_9079,N_9659);
and U10498 (N_10498,N_8152,N_9804);
nor U10499 (N_10499,N_8642,N_9442);
xor U10500 (N_10500,N_9321,N_8251);
nor U10501 (N_10501,N_8843,N_8309);
or U10502 (N_10502,N_9430,N_9242);
nand U10503 (N_10503,N_8799,N_8666);
and U10504 (N_10504,N_8162,N_9240);
and U10505 (N_10505,N_9388,N_8906);
nor U10506 (N_10506,N_8109,N_8179);
nand U10507 (N_10507,N_8673,N_9407);
nand U10508 (N_10508,N_9209,N_8929);
and U10509 (N_10509,N_8006,N_9399);
nor U10510 (N_10510,N_8678,N_9215);
and U10511 (N_10511,N_8004,N_9609);
and U10512 (N_10512,N_9196,N_8447);
xor U10513 (N_10513,N_9560,N_8046);
nand U10514 (N_10514,N_9715,N_9797);
nor U10515 (N_10515,N_9664,N_9773);
nor U10516 (N_10516,N_9105,N_9536);
nand U10517 (N_10517,N_9471,N_8590);
or U10518 (N_10518,N_8647,N_9732);
nor U10519 (N_10519,N_9962,N_8220);
nor U10520 (N_10520,N_9572,N_9331);
and U10521 (N_10521,N_9333,N_8065);
nor U10522 (N_10522,N_8407,N_8912);
nand U10523 (N_10523,N_9754,N_9674);
or U10524 (N_10524,N_8644,N_8699);
nor U10525 (N_10525,N_9567,N_8963);
and U10526 (N_10526,N_8164,N_9594);
nor U10527 (N_10527,N_9191,N_8180);
and U10528 (N_10528,N_9378,N_9966);
nand U10529 (N_10529,N_9785,N_9384);
or U10530 (N_10530,N_9725,N_8434);
nand U10531 (N_10531,N_8710,N_8967);
and U10532 (N_10532,N_8549,N_8547);
nor U10533 (N_10533,N_8097,N_8705);
xor U10534 (N_10534,N_8034,N_9436);
or U10535 (N_10535,N_9468,N_9201);
xnor U10536 (N_10536,N_9992,N_8909);
or U10537 (N_10537,N_9866,N_8479);
nand U10538 (N_10538,N_9381,N_9721);
or U10539 (N_10539,N_8950,N_9489);
or U10540 (N_10540,N_9221,N_9457);
nor U10541 (N_10541,N_8551,N_9461);
xnor U10542 (N_10542,N_9340,N_9534);
and U10543 (N_10543,N_9431,N_9035);
nand U10544 (N_10544,N_8687,N_9629);
or U10545 (N_10545,N_9760,N_9547);
nand U10546 (N_10546,N_8648,N_8093);
or U10547 (N_10547,N_9526,N_8855);
nand U10548 (N_10548,N_8459,N_9287);
and U10549 (N_10549,N_9015,N_9818);
xor U10550 (N_10550,N_9769,N_8861);
nor U10551 (N_10551,N_8779,N_9133);
nand U10552 (N_10552,N_9790,N_9167);
nor U10553 (N_10553,N_9807,N_8441);
nand U10554 (N_10554,N_8679,N_9043);
nor U10555 (N_10555,N_8630,N_9055);
or U10556 (N_10556,N_9059,N_8574);
nor U10557 (N_10557,N_9400,N_9232);
xnor U10558 (N_10558,N_9627,N_9485);
or U10559 (N_10559,N_8452,N_8112);
nor U10560 (N_10560,N_9645,N_8099);
or U10561 (N_10561,N_8261,N_8729);
or U10562 (N_10562,N_9530,N_9612);
nand U10563 (N_10563,N_9066,N_8839);
and U10564 (N_10564,N_8045,N_9370);
nand U10565 (N_10565,N_9863,N_8542);
or U10566 (N_10566,N_8031,N_9896);
xor U10567 (N_10567,N_9120,N_9667);
and U10568 (N_10568,N_8570,N_8803);
or U10569 (N_10569,N_8736,N_9551);
xor U10570 (N_10570,N_9755,N_9756);
or U10571 (N_10571,N_9784,N_9467);
nor U10572 (N_10572,N_8813,N_9739);
or U10573 (N_10573,N_9192,N_9506);
and U10574 (N_10574,N_8735,N_8489);
nand U10575 (N_10575,N_8258,N_8879);
nand U10576 (N_10576,N_8081,N_8558);
nand U10577 (N_10577,N_9595,N_9539);
or U10578 (N_10578,N_9346,N_8103);
nor U10579 (N_10579,N_9494,N_8757);
nor U10580 (N_10580,N_9957,N_8907);
nand U10581 (N_10581,N_8528,N_8266);
and U10582 (N_10582,N_8206,N_9631);
and U10583 (N_10583,N_9600,N_9171);
xnor U10584 (N_10584,N_9857,N_8713);
and U10585 (N_10585,N_8981,N_9127);
xnor U10586 (N_10586,N_9348,N_9747);
or U10587 (N_10587,N_8395,N_9749);
and U10588 (N_10588,N_8854,N_8603);
nand U10589 (N_10589,N_8373,N_9614);
or U10590 (N_10590,N_8408,N_8812);
nand U10591 (N_10591,N_8508,N_8543);
nand U10592 (N_10592,N_9628,N_8380);
and U10593 (N_10593,N_8943,N_9311);
nor U10594 (N_10594,N_8616,N_8617);
nand U10595 (N_10595,N_8988,N_8656);
xor U10596 (N_10596,N_9854,N_8235);
nor U10597 (N_10597,N_8313,N_8063);
and U10598 (N_10598,N_8484,N_8042);
and U10599 (N_10599,N_9248,N_8908);
nand U10600 (N_10600,N_9366,N_8100);
nor U10601 (N_10601,N_8814,N_9830);
xnor U10602 (N_10602,N_9022,N_9497);
nand U10603 (N_10603,N_9288,N_8121);
xnor U10604 (N_10604,N_9717,N_8684);
and U10605 (N_10605,N_8064,N_8106);
nand U10606 (N_10606,N_8798,N_9586);
or U10607 (N_10607,N_9566,N_8746);
nor U10608 (N_10608,N_8521,N_9433);
or U10609 (N_10609,N_8000,N_8758);
and U10610 (N_10610,N_8789,N_9161);
and U10611 (N_10611,N_9315,N_9842);
or U10612 (N_10612,N_8703,N_8033);
nor U10613 (N_10613,N_9410,N_9216);
nand U10614 (N_10614,N_9805,N_8041);
or U10615 (N_10615,N_9809,N_9990);
nand U10616 (N_10616,N_9993,N_9131);
or U10617 (N_10617,N_8321,N_8389);
nor U10618 (N_10618,N_8763,N_9563);
xnor U10619 (N_10619,N_9603,N_9389);
and U10620 (N_10620,N_8221,N_9505);
and U10621 (N_10621,N_8933,N_8627);
nor U10622 (N_10622,N_9089,N_9210);
nand U10623 (N_10623,N_9546,N_9808);
nor U10624 (N_10624,N_8876,N_9929);
and U10625 (N_10625,N_8372,N_8199);
and U10626 (N_10626,N_8413,N_8070);
or U10627 (N_10627,N_8445,N_9571);
or U10628 (N_10628,N_9082,N_8335);
and U10629 (N_10629,N_8849,N_8398);
or U10630 (N_10630,N_9438,N_9140);
nor U10631 (N_10631,N_9336,N_8766);
nand U10632 (N_10632,N_9011,N_9474);
nor U10633 (N_10633,N_9848,N_8864);
or U10634 (N_10634,N_9897,N_9391);
nor U10635 (N_10635,N_8836,N_9393);
nor U10636 (N_10636,N_8463,N_8764);
nand U10637 (N_10637,N_9032,N_8683);
and U10638 (N_10638,N_8808,N_9891);
nor U10639 (N_10639,N_9967,N_8932);
or U10640 (N_10640,N_9758,N_8599);
or U10641 (N_10641,N_8748,N_8350);
and U10642 (N_10642,N_8137,N_9325);
and U10643 (N_10643,N_9995,N_8249);
xnor U10644 (N_10644,N_8515,N_9093);
and U10645 (N_10645,N_8979,N_9246);
nand U10646 (N_10646,N_8440,N_9657);
nor U10647 (N_10647,N_9211,N_8762);
or U10648 (N_10648,N_8991,N_9528);
xnor U10649 (N_10649,N_9765,N_9282);
or U10650 (N_10650,N_9233,N_9352);
nor U10651 (N_10651,N_8690,N_8188);
and U10652 (N_10652,N_9545,N_9509);
or U10653 (N_10653,N_8374,N_9009);
xnor U10654 (N_10654,N_8011,N_8791);
and U10655 (N_10655,N_8271,N_9285);
nand U10656 (N_10656,N_8900,N_9324);
and U10657 (N_10657,N_8823,N_8028);
or U10658 (N_10658,N_9770,N_8743);
and U10659 (N_10659,N_9481,N_9465);
or U10660 (N_10660,N_8057,N_8018);
nor U10661 (N_10661,N_8001,N_8941);
nand U10662 (N_10662,N_8320,N_8104);
nand U10663 (N_10663,N_8439,N_8794);
xnor U10664 (N_10664,N_8875,N_8801);
nor U10665 (N_10665,N_9439,N_9229);
nand U10666 (N_10666,N_9249,N_9337);
xnor U10667 (N_10667,N_8364,N_8577);
nand U10668 (N_10668,N_9459,N_8387);
or U10669 (N_10669,N_9185,N_9052);
or U10670 (N_10670,N_9559,N_9275);
and U10671 (N_10671,N_8473,N_8136);
or U10672 (N_10672,N_8306,N_8928);
nor U10673 (N_10673,N_9580,N_8910);
or U10674 (N_10674,N_9895,N_9942);
or U10675 (N_10675,N_9937,N_8326);
nor U10676 (N_10676,N_8451,N_9781);
or U10677 (N_10677,N_8819,N_8804);
nand U10678 (N_10678,N_8959,N_9867);
nand U10679 (N_10679,N_8146,N_8403);
nor U10680 (N_10680,N_8692,N_8143);
nand U10681 (N_10681,N_9362,N_9825);
and U10682 (N_10682,N_9648,N_9693);
xnor U10683 (N_10683,N_9299,N_8371);
nor U10684 (N_10684,N_9223,N_9875);
and U10685 (N_10685,N_9042,N_9908);
nand U10686 (N_10686,N_8135,N_8356);
and U10687 (N_10687,N_9006,N_9235);
and U10688 (N_10688,N_9543,N_8150);
nor U10689 (N_10689,N_8385,N_8123);
nand U10690 (N_10690,N_8778,N_8254);
nand U10691 (N_10691,N_8878,N_8280);
and U10692 (N_10692,N_9239,N_8344);
or U10693 (N_10693,N_9179,N_8122);
xor U10694 (N_10694,N_8120,N_9923);
nor U10695 (N_10695,N_8931,N_9306);
nor U10696 (N_10696,N_9053,N_9102);
xor U10697 (N_10697,N_8003,N_9561);
nor U10698 (N_10698,N_8036,N_8458);
nor U10699 (N_10699,N_8217,N_9736);
nor U10700 (N_10700,N_9675,N_9159);
and U10701 (N_10701,N_8133,N_8088);
nor U10702 (N_10702,N_9704,N_8486);
xnor U10703 (N_10703,N_8068,N_8124);
nand U10704 (N_10704,N_8987,N_9964);
and U10705 (N_10705,N_9342,N_8465);
nand U10706 (N_10706,N_8450,N_8289);
nor U10707 (N_10707,N_8357,N_8788);
nand U10708 (N_10708,N_8811,N_9598);
nor U10709 (N_10709,N_9313,N_8960);
nand U10710 (N_10710,N_9816,N_8992);
nand U10711 (N_10711,N_9889,N_9213);
nand U10712 (N_10712,N_8163,N_9669);
xnor U10713 (N_10713,N_8796,N_8241);
nor U10714 (N_10714,N_8701,N_9377);
nand U10715 (N_10715,N_9220,N_8783);
nor U10716 (N_10716,N_9398,N_9110);
nand U10717 (N_10717,N_9426,N_8887);
and U10718 (N_10718,N_9217,N_8852);
or U10719 (N_10719,N_8660,N_8613);
nor U10720 (N_10720,N_8172,N_9456);
nor U10721 (N_10721,N_9405,N_9199);
and U10722 (N_10722,N_9435,N_9815);
or U10723 (N_10723,N_9727,N_9025);
nand U10724 (N_10724,N_9160,N_8330);
xnor U10725 (N_10725,N_9358,N_8273);
and U10726 (N_10726,N_9673,N_9849);
or U10727 (N_10727,N_8075,N_8537);
nand U10728 (N_10728,N_9361,N_9394);
and U10729 (N_10729,N_8114,N_9880);
nand U10730 (N_10730,N_9688,N_9277);
nor U10731 (N_10731,N_9682,N_8411);
nor U10732 (N_10732,N_9041,N_9307);
and U10733 (N_10733,N_8918,N_9553);
or U10734 (N_10734,N_9928,N_9448);
or U10735 (N_10735,N_9638,N_8724);
and U10736 (N_10736,N_8069,N_9247);
or U10737 (N_10737,N_9162,N_8555);
xor U10738 (N_10738,N_8921,N_9137);
and U10739 (N_10739,N_8596,N_8646);
xnor U10740 (N_10740,N_9514,N_9444);
nor U10741 (N_10741,N_8454,N_9817);
and U10742 (N_10742,N_8857,N_9901);
or U10743 (N_10743,N_9835,N_8059);
nand U10744 (N_10744,N_9255,N_8119);
xnor U10745 (N_10745,N_8369,N_8576);
or U10746 (N_10746,N_8359,N_8032);
xnor U10747 (N_10747,N_8500,N_9565);
or U10748 (N_10748,N_8522,N_9005);
and U10749 (N_10749,N_8010,N_9475);
xnor U10750 (N_10750,N_9941,N_8402);
nor U10751 (N_10751,N_9230,N_8571);
nor U10752 (N_10752,N_9144,N_9836);
nor U10753 (N_10753,N_8215,N_8990);
nor U10754 (N_10754,N_9916,N_8494);
nor U10755 (N_10755,N_9379,N_8502);
nor U10756 (N_10756,N_9371,N_9799);
xor U10757 (N_10757,N_9504,N_9124);
nor U10758 (N_10758,N_9353,N_8467);
and U10759 (N_10759,N_8756,N_8828);
nand U10760 (N_10760,N_8365,N_8512);
xnor U10761 (N_10761,N_8726,N_8169);
nor U10762 (N_10762,N_8770,N_8998);
and U10763 (N_10763,N_9621,N_9924);
and U10764 (N_10764,N_8181,N_8216);
xnor U10765 (N_10765,N_9317,N_9048);
nor U10766 (N_10766,N_8472,N_9134);
nand U10767 (N_10767,N_9451,N_8115);
and U10768 (N_10768,N_8117,N_9512);
nand U10769 (N_10769,N_9188,N_9914);
or U10770 (N_10770,N_8604,N_9508);
or U10771 (N_10771,N_9855,N_9114);
nand U10772 (N_10772,N_9480,N_8025);
xnor U10773 (N_10773,N_8319,N_9101);
and U10774 (N_10774,N_8224,N_8822);
or U10775 (N_10775,N_9984,N_9602);
nor U10776 (N_10776,N_9500,N_9945);
xor U10777 (N_10777,N_9222,N_8147);
nor U10778 (N_10778,N_9254,N_9194);
nand U10779 (N_10779,N_8229,N_8388);
nand U10780 (N_10780,N_9626,N_9738);
or U10781 (N_10781,N_8649,N_9047);
nand U10782 (N_10782,N_9503,N_8824);
and U10783 (N_10783,N_9953,N_9510);
nor U10784 (N_10784,N_9045,N_8368);
nor U10785 (N_10785,N_9077,N_9068);
xnor U10786 (N_10786,N_8107,N_8012);
or U10787 (N_10787,N_9128,N_8635);
nor U10788 (N_10788,N_9126,N_8376);
or U10789 (N_10789,N_9930,N_9476);
nor U10790 (N_10790,N_9412,N_9668);
or U10791 (N_10791,N_8098,N_9520);
and U10792 (N_10792,N_9989,N_8396);
nor U10793 (N_10793,N_8688,N_8270);
and U10794 (N_10794,N_9862,N_8728);
and U10795 (N_10795,N_8422,N_9428);
nor U10796 (N_10796,N_9338,N_8481);
nor U10797 (N_10797,N_8085,N_8035);
xor U10798 (N_10798,N_8391,N_8501);
and U10799 (N_10799,N_8091,N_9177);
nor U10800 (N_10800,N_9699,N_8269);
nor U10801 (N_10801,N_9696,N_9057);
or U10802 (N_10802,N_9680,N_8253);
xor U10803 (N_10803,N_8834,N_9518);
nand U10804 (N_10804,N_9649,N_8301);
xor U10805 (N_10805,N_8089,N_9406);
and U10806 (N_10806,N_9764,N_9098);
and U10807 (N_10807,N_8694,N_9584);
or U10808 (N_10808,N_9874,N_9470);
nand U10809 (N_10809,N_9960,N_9814);
nand U10810 (N_10810,N_9639,N_8333);
nor U10811 (N_10811,N_8327,N_9819);
xor U10812 (N_10812,N_8307,N_9116);
and U10813 (N_10813,N_8332,N_8497);
or U10814 (N_10814,N_8378,N_8110);
or U10815 (N_10815,N_8438,N_8969);
nand U10816 (N_10816,N_9466,N_9588);
nor U10817 (N_10817,N_9578,N_9952);
and U10818 (N_10818,N_8349,N_8708);
and U10819 (N_10819,N_9670,N_9792);
or U10820 (N_10820,N_8029,N_9411);
and U10821 (N_10821,N_8607,N_8902);
xor U10822 (N_10822,N_9837,N_9111);
or U10823 (N_10823,N_9703,N_8895);
nor U10824 (N_10824,N_8524,N_9521);
nand U10825 (N_10825,N_9846,N_8626);
and U10826 (N_10826,N_8880,N_9106);
nand U10827 (N_10827,N_9050,N_8488);
nand U10828 (N_10828,N_8080,N_8598);
nand U10829 (N_10829,N_8806,N_9019);
and U10830 (N_10830,N_9228,N_8334);
nand U10831 (N_10831,N_9973,N_8134);
or U10832 (N_10832,N_8795,N_9881);
or U10833 (N_10833,N_9793,N_8303);
and U10834 (N_10834,N_8625,N_8049);
nand U10835 (N_10835,N_9121,N_8482);
nand U10836 (N_10836,N_8436,N_9582);
nand U10837 (N_10837,N_9269,N_8297);
or U10838 (N_10838,N_8393,N_8514);
nand U10839 (N_10839,N_9452,N_8838);
or U10840 (N_10840,N_9806,N_8170);
or U10841 (N_10841,N_9887,N_9251);
or U10842 (N_10842,N_8207,N_9113);
and U10843 (N_10843,N_9533,N_8384);
xor U10844 (N_10844,N_9886,N_9801);
and U10845 (N_10845,N_9256,N_8295);
xor U10846 (N_10846,N_9856,N_9744);
nand U10847 (N_10847,N_9104,N_9898);
or U10848 (N_10848,N_9540,N_8620);
xnor U10849 (N_10849,N_8925,N_9911);
nand U10850 (N_10850,N_9073,N_8038);
nand U10851 (N_10851,N_9507,N_9813);
or U10852 (N_10852,N_8983,N_9917);
and U10853 (N_10853,N_9646,N_9997);
and U10854 (N_10854,N_8466,N_9983);
and U10855 (N_10855,N_8300,N_9968);
and U10856 (N_10856,N_9359,N_8851);
xnor U10857 (N_10857,N_9364,N_8742);
or U10858 (N_10858,N_8831,N_9091);
or U10859 (N_10859,N_9023,N_8552);
and U10860 (N_10860,N_9260,N_8675);
xnor U10861 (N_10861,N_8219,N_8358);
or U10862 (N_10862,N_9789,N_8695);
or U10863 (N_10863,N_8632,N_8591);
and U10864 (N_10864,N_9051,N_8631);
and U10865 (N_10865,N_8144,N_9146);
and U10866 (N_10866,N_8573,N_9831);
nand U10867 (N_10867,N_9802,N_9004);
and U10868 (N_10868,N_9681,N_8095);
or U10869 (N_10869,N_9291,N_9878);
nor U10870 (N_10870,N_8592,N_9720);
nand U10871 (N_10871,N_8014,N_8503);
nand U10872 (N_10872,N_9610,N_9176);
and U10873 (N_10873,N_8155,N_8965);
and U10874 (N_10874,N_9557,N_8074);
nand U10875 (N_10875,N_9906,N_8165);
and U10876 (N_10876,N_8589,N_8897);
nand U10877 (N_10877,N_8948,N_8622);
nand U10878 (N_10878,N_9309,N_8250);
and U10879 (N_10879,N_9909,N_9163);
and U10880 (N_10880,N_9882,N_9757);
or U10881 (N_10881,N_8140,N_9189);
nor U10882 (N_10882,N_8354,N_8966);
nor U10883 (N_10883,N_9666,N_8944);
or U10884 (N_10884,N_9538,N_8659);
or U10885 (N_10885,N_8182,N_9652);
and U10886 (N_10886,N_9000,N_8924);
xor U10887 (N_10887,N_8583,N_8072);
and U10888 (N_10888,N_9723,N_9524);
and U10889 (N_10889,N_8201,N_9963);
and U10890 (N_10890,N_9495,N_9907);
nor U10891 (N_10891,N_8572,N_8860);
or U10892 (N_10892,N_8336,N_9777);
xnor U10893 (N_10893,N_9178,N_9071);
nand U10894 (N_10894,N_9999,N_8086);
nor U10895 (N_10895,N_8550,N_9304);
and U10896 (N_10896,N_8244,N_9376);
nand U10897 (N_10897,N_8151,N_9383);
or U10898 (N_10898,N_8185,N_8236);
and U10899 (N_10899,N_8827,N_9087);
nor U10900 (N_10900,N_9152,N_9270);
and U10901 (N_10901,N_9951,N_8424);
or U10902 (N_10902,N_8315,N_8615);
or U10903 (N_10903,N_8277,N_9979);
nand U10904 (N_10904,N_9202,N_8629);
or U10905 (N_10905,N_8200,N_9118);
xor U10906 (N_10906,N_9181,N_9976);
and U10907 (N_10907,N_8760,N_8294);
and U10908 (N_10908,N_8184,N_8276);
nand U10909 (N_10909,N_9811,N_8884);
nand U10910 (N_10910,N_8455,N_8787);
nand U10911 (N_10911,N_9469,N_8329);
nand U10912 (N_10912,N_9273,N_9449);
nor U10913 (N_10913,N_8562,N_9292);
nand U10914 (N_10914,N_8662,N_9653);
and U10915 (N_10915,N_9347,N_8947);
or U10916 (N_10916,N_8485,N_8686);
and U10917 (N_10917,N_9069,N_9363);
xnor U10918 (N_10918,N_9803,N_8892);
or U10919 (N_10919,N_8382,N_9954);
nor U10920 (N_10920,N_8721,N_8832);
and U10921 (N_10921,N_9623,N_9959);
or U10922 (N_10922,N_8565,N_9912);
nor U10923 (N_10923,N_8202,N_9060);
and U10924 (N_10924,N_9088,N_8007);
or U10925 (N_10925,N_9076,N_9084);
xor U10926 (N_10926,N_9501,N_8347);
nor U10927 (N_10927,N_9759,N_8877);
nor U10928 (N_10928,N_8759,N_8268);
or U10929 (N_10929,N_8149,N_9778);
nor U10930 (N_10930,N_9731,N_8994);
nand U10931 (N_10931,N_9853,N_8498);
and U10932 (N_10932,N_9910,N_9970);
and U10933 (N_10933,N_8419,N_8698);
or U10934 (N_10934,N_9001,N_9175);
or U10935 (N_10935,N_8312,N_9351);
xnor U10936 (N_10936,N_8338,N_8138);
and U10937 (N_10937,N_9763,N_9123);
and U10938 (N_10938,N_8985,N_9119);
and U10939 (N_10939,N_8752,N_9258);
xor U10940 (N_10940,N_8668,N_9665);
nand U10941 (N_10941,N_9445,N_9786);
nor U10942 (N_10942,N_8279,N_9002);
nor U10943 (N_10943,N_8246,N_9294);
and U10944 (N_10944,N_9372,N_9416);
nor U10945 (N_10945,N_9036,N_9204);
or U10946 (N_10946,N_8410,N_9656);
and U10947 (N_10947,N_8609,N_8311);
nor U10948 (N_10948,N_8519,N_9206);
nor U10949 (N_10949,N_8213,N_9599);
nand U10950 (N_10950,N_9980,N_9499);
xnor U10951 (N_10951,N_8942,N_9532);
nand U10952 (N_10952,N_8601,N_9712);
xnor U10953 (N_10953,N_8732,N_9484);
nor U10954 (N_10954,N_8343,N_9141);
and U10955 (N_10955,N_8079,N_9165);
nor U10956 (N_10956,N_9574,N_8747);
and U10957 (N_10957,N_9312,N_8462);
or U10958 (N_10958,N_8116,N_9172);
or U10959 (N_10959,N_9024,N_8654);
xor U10960 (N_10960,N_8848,N_8636);
or U10961 (N_10961,N_9062,N_9044);
nor U10962 (N_10962,N_8414,N_8259);
and U10963 (N_10963,N_8073,N_8602);
nand U10964 (N_10964,N_9750,N_8984);
nor U10965 (N_10965,N_9070,N_9208);
xor U10966 (N_10966,N_9554,N_9401);
or U10967 (N_10967,N_9462,N_9262);
nand U10968 (N_10968,N_9611,N_8158);
and U10969 (N_10969,N_9432,N_8645);
nand U10970 (N_10970,N_8189,N_8529);
or U10971 (N_10971,N_8658,N_8324);
and U10972 (N_10972,N_9931,N_8090);
and U10973 (N_10973,N_8844,N_8923);
and U10974 (N_10974,N_8891,N_9794);
nor U10975 (N_10975,N_9392,N_8305);
nor U10976 (N_10976,N_9281,N_8527);
nand U10977 (N_10977,N_9488,N_8505);
nand U10978 (N_10978,N_8639,N_9473);
nor U10979 (N_10979,N_8540,N_9729);
nor U10980 (N_10980,N_9203,N_9879);
and U10981 (N_10981,N_9926,N_9302);
nor U10982 (N_10982,N_9155,N_9986);
nor U10983 (N_10983,N_9017,N_8930);
nand U10984 (N_10984,N_9100,N_9812);
nand U10985 (N_10985,N_8048,N_9994);
and U10986 (N_10986,N_8023,N_9515);
nand U10987 (N_10987,N_9589,N_9117);
or U10988 (N_10988,N_9450,N_8914);
and U10989 (N_10989,N_9150,N_9991);
and U10990 (N_10990,N_8643,N_8955);
or U10991 (N_10991,N_8131,N_9301);
or U10992 (N_10992,N_9086,N_9934);
nand U10993 (N_10993,N_9686,N_8432);
and U10994 (N_10994,N_9692,N_8773);
nand U10995 (N_10995,N_9263,N_8720);
nand U10996 (N_10996,N_8239,N_9734);
nand U10997 (N_10997,N_8739,N_9224);
or U10998 (N_10998,N_9380,N_9092);
or U10999 (N_10999,N_8262,N_8340);
or U11000 (N_11000,N_8957,N_9102);
and U11001 (N_11001,N_9232,N_9695);
nor U11002 (N_11002,N_8513,N_9588);
nor U11003 (N_11003,N_8998,N_8229);
or U11004 (N_11004,N_8765,N_9475);
nand U11005 (N_11005,N_8594,N_8087);
and U11006 (N_11006,N_8680,N_9432);
xnor U11007 (N_11007,N_8738,N_8999);
nor U11008 (N_11008,N_8135,N_9218);
nand U11009 (N_11009,N_9773,N_8152);
and U11010 (N_11010,N_9815,N_9280);
or U11011 (N_11011,N_9370,N_9722);
and U11012 (N_11012,N_9401,N_8543);
or U11013 (N_11013,N_9667,N_9004);
or U11014 (N_11014,N_9654,N_8177);
and U11015 (N_11015,N_9571,N_8012);
and U11016 (N_11016,N_8674,N_8128);
xor U11017 (N_11017,N_9338,N_8925);
xnor U11018 (N_11018,N_9934,N_8567);
nand U11019 (N_11019,N_8160,N_8031);
xor U11020 (N_11020,N_9088,N_8091);
or U11021 (N_11021,N_9553,N_8531);
nor U11022 (N_11022,N_9115,N_8885);
nor U11023 (N_11023,N_9852,N_8691);
nand U11024 (N_11024,N_9652,N_9011);
or U11025 (N_11025,N_9395,N_9750);
nand U11026 (N_11026,N_8953,N_9815);
xnor U11027 (N_11027,N_8070,N_9574);
and U11028 (N_11028,N_9529,N_8139);
nor U11029 (N_11029,N_8217,N_9489);
nand U11030 (N_11030,N_8324,N_9889);
or U11031 (N_11031,N_9216,N_9339);
nand U11032 (N_11032,N_8277,N_9814);
nand U11033 (N_11033,N_8622,N_8338);
or U11034 (N_11034,N_9267,N_9140);
nand U11035 (N_11035,N_9891,N_8892);
xnor U11036 (N_11036,N_8174,N_9177);
and U11037 (N_11037,N_8436,N_9072);
nand U11038 (N_11038,N_9517,N_9272);
or U11039 (N_11039,N_9290,N_8051);
and U11040 (N_11040,N_8124,N_9197);
or U11041 (N_11041,N_9498,N_8403);
and U11042 (N_11042,N_9678,N_9496);
xnor U11043 (N_11043,N_8827,N_8127);
nand U11044 (N_11044,N_8968,N_8393);
nand U11045 (N_11045,N_8231,N_8949);
and U11046 (N_11046,N_8608,N_8171);
or U11047 (N_11047,N_9044,N_9316);
nor U11048 (N_11048,N_9720,N_8252);
nor U11049 (N_11049,N_8666,N_9471);
nand U11050 (N_11050,N_8413,N_8150);
and U11051 (N_11051,N_9765,N_9014);
or U11052 (N_11052,N_9396,N_8584);
xor U11053 (N_11053,N_8562,N_9455);
nor U11054 (N_11054,N_8331,N_8308);
nand U11055 (N_11055,N_8229,N_9752);
and U11056 (N_11056,N_8925,N_9123);
nor U11057 (N_11057,N_9093,N_8186);
nor U11058 (N_11058,N_8054,N_8946);
nand U11059 (N_11059,N_8499,N_8729);
nor U11060 (N_11060,N_8936,N_9146);
or U11061 (N_11061,N_8957,N_9740);
nor U11062 (N_11062,N_8139,N_9285);
xor U11063 (N_11063,N_8065,N_9300);
or U11064 (N_11064,N_8773,N_9826);
nor U11065 (N_11065,N_9997,N_9118);
or U11066 (N_11066,N_9702,N_8582);
nand U11067 (N_11067,N_9414,N_9218);
and U11068 (N_11068,N_8773,N_8324);
xnor U11069 (N_11069,N_9073,N_8603);
nor U11070 (N_11070,N_8113,N_8886);
nor U11071 (N_11071,N_9178,N_8363);
nor U11072 (N_11072,N_9576,N_9665);
nor U11073 (N_11073,N_8439,N_9995);
nor U11074 (N_11074,N_8090,N_9485);
or U11075 (N_11075,N_8690,N_8544);
xnor U11076 (N_11076,N_9378,N_8587);
nand U11077 (N_11077,N_8393,N_8462);
nor U11078 (N_11078,N_9097,N_9113);
or U11079 (N_11079,N_8981,N_8287);
or U11080 (N_11080,N_9864,N_9451);
nor U11081 (N_11081,N_9845,N_8200);
and U11082 (N_11082,N_8411,N_9884);
xnor U11083 (N_11083,N_8327,N_8876);
nand U11084 (N_11084,N_8183,N_9260);
or U11085 (N_11085,N_9995,N_9502);
nand U11086 (N_11086,N_8779,N_8228);
nor U11087 (N_11087,N_8004,N_8063);
xor U11088 (N_11088,N_9284,N_8184);
nor U11089 (N_11089,N_8906,N_9206);
nor U11090 (N_11090,N_9131,N_9941);
nor U11091 (N_11091,N_9610,N_9600);
nor U11092 (N_11092,N_9220,N_8166);
nor U11093 (N_11093,N_8173,N_9565);
xor U11094 (N_11094,N_9238,N_8232);
nor U11095 (N_11095,N_9208,N_9600);
nor U11096 (N_11096,N_9052,N_8710);
or U11097 (N_11097,N_8980,N_9584);
xor U11098 (N_11098,N_8988,N_8511);
xor U11099 (N_11099,N_9207,N_8628);
and U11100 (N_11100,N_9034,N_9024);
or U11101 (N_11101,N_8418,N_9094);
and U11102 (N_11102,N_8809,N_8778);
or U11103 (N_11103,N_9618,N_9951);
nor U11104 (N_11104,N_9804,N_8768);
nor U11105 (N_11105,N_8199,N_9549);
or U11106 (N_11106,N_8132,N_8491);
nor U11107 (N_11107,N_9483,N_9211);
and U11108 (N_11108,N_8091,N_9724);
nand U11109 (N_11109,N_8204,N_9596);
nand U11110 (N_11110,N_9143,N_8308);
xnor U11111 (N_11111,N_8406,N_9739);
xnor U11112 (N_11112,N_9431,N_8971);
nor U11113 (N_11113,N_8168,N_8413);
or U11114 (N_11114,N_9798,N_8116);
or U11115 (N_11115,N_9294,N_9812);
nor U11116 (N_11116,N_9424,N_9740);
or U11117 (N_11117,N_8653,N_9580);
nand U11118 (N_11118,N_9622,N_9364);
and U11119 (N_11119,N_9854,N_8821);
and U11120 (N_11120,N_8853,N_9624);
nand U11121 (N_11121,N_9751,N_9305);
xnor U11122 (N_11122,N_9001,N_9212);
or U11123 (N_11123,N_9438,N_8083);
nand U11124 (N_11124,N_9913,N_8882);
nor U11125 (N_11125,N_8630,N_8648);
or U11126 (N_11126,N_9758,N_9613);
or U11127 (N_11127,N_8953,N_9414);
nand U11128 (N_11128,N_9890,N_8739);
nand U11129 (N_11129,N_8717,N_9863);
or U11130 (N_11130,N_8545,N_8556);
nand U11131 (N_11131,N_8207,N_8016);
or U11132 (N_11132,N_9395,N_8727);
or U11133 (N_11133,N_8648,N_9667);
and U11134 (N_11134,N_9228,N_9126);
nand U11135 (N_11135,N_9357,N_9377);
nand U11136 (N_11136,N_9124,N_9060);
or U11137 (N_11137,N_9099,N_9581);
nor U11138 (N_11138,N_8371,N_8143);
nand U11139 (N_11139,N_9981,N_9876);
or U11140 (N_11140,N_8050,N_9256);
nand U11141 (N_11141,N_9511,N_8200);
and U11142 (N_11142,N_9522,N_8415);
or U11143 (N_11143,N_8155,N_9332);
nor U11144 (N_11144,N_9588,N_8836);
or U11145 (N_11145,N_9010,N_8479);
nor U11146 (N_11146,N_9468,N_9868);
nor U11147 (N_11147,N_9588,N_9438);
or U11148 (N_11148,N_8517,N_8166);
or U11149 (N_11149,N_9092,N_8482);
or U11150 (N_11150,N_8105,N_8647);
nor U11151 (N_11151,N_9699,N_9210);
nand U11152 (N_11152,N_8385,N_9401);
nor U11153 (N_11153,N_9699,N_8322);
or U11154 (N_11154,N_8833,N_8031);
nor U11155 (N_11155,N_9455,N_9436);
or U11156 (N_11156,N_8834,N_9413);
and U11157 (N_11157,N_8022,N_8004);
nand U11158 (N_11158,N_8147,N_8046);
or U11159 (N_11159,N_8950,N_9781);
nor U11160 (N_11160,N_9875,N_8814);
nor U11161 (N_11161,N_8079,N_8988);
nand U11162 (N_11162,N_8961,N_9651);
nor U11163 (N_11163,N_9193,N_8208);
and U11164 (N_11164,N_8225,N_9707);
xnor U11165 (N_11165,N_9617,N_8458);
xnor U11166 (N_11166,N_9715,N_9463);
or U11167 (N_11167,N_8157,N_8652);
and U11168 (N_11168,N_8753,N_8328);
or U11169 (N_11169,N_9471,N_9130);
and U11170 (N_11170,N_8411,N_9753);
and U11171 (N_11171,N_9672,N_8992);
nand U11172 (N_11172,N_8518,N_9402);
nor U11173 (N_11173,N_9043,N_8593);
nor U11174 (N_11174,N_9778,N_8645);
or U11175 (N_11175,N_9749,N_9006);
nand U11176 (N_11176,N_8935,N_9371);
xnor U11177 (N_11177,N_8300,N_8424);
and U11178 (N_11178,N_9459,N_8497);
nor U11179 (N_11179,N_9331,N_9327);
nand U11180 (N_11180,N_8354,N_9514);
nand U11181 (N_11181,N_9073,N_9285);
and U11182 (N_11182,N_9862,N_8641);
or U11183 (N_11183,N_9745,N_8384);
nor U11184 (N_11184,N_9680,N_9108);
nand U11185 (N_11185,N_9229,N_8743);
xnor U11186 (N_11186,N_8170,N_8908);
nor U11187 (N_11187,N_8456,N_9567);
or U11188 (N_11188,N_9790,N_9132);
and U11189 (N_11189,N_9802,N_9923);
nor U11190 (N_11190,N_9836,N_8148);
nor U11191 (N_11191,N_8196,N_9486);
and U11192 (N_11192,N_9827,N_9177);
or U11193 (N_11193,N_9736,N_8907);
and U11194 (N_11194,N_8782,N_9128);
or U11195 (N_11195,N_9904,N_8174);
xnor U11196 (N_11196,N_9019,N_9199);
nand U11197 (N_11197,N_9048,N_8602);
xor U11198 (N_11198,N_8955,N_8481);
or U11199 (N_11199,N_8952,N_8743);
xnor U11200 (N_11200,N_8527,N_8555);
nand U11201 (N_11201,N_8308,N_8225);
xor U11202 (N_11202,N_8272,N_9801);
nor U11203 (N_11203,N_8600,N_8954);
or U11204 (N_11204,N_8619,N_8117);
or U11205 (N_11205,N_9909,N_9921);
and U11206 (N_11206,N_9271,N_9288);
and U11207 (N_11207,N_8013,N_9739);
nand U11208 (N_11208,N_9288,N_9708);
nor U11209 (N_11209,N_8985,N_8925);
or U11210 (N_11210,N_8679,N_8614);
xnor U11211 (N_11211,N_8453,N_8152);
or U11212 (N_11212,N_8516,N_9868);
nand U11213 (N_11213,N_9683,N_8875);
nor U11214 (N_11214,N_9150,N_8272);
nand U11215 (N_11215,N_9035,N_9882);
nand U11216 (N_11216,N_9185,N_8213);
nand U11217 (N_11217,N_9687,N_8417);
nor U11218 (N_11218,N_8853,N_8959);
nor U11219 (N_11219,N_8913,N_9459);
and U11220 (N_11220,N_9205,N_9143);
and U11221 (N_11221,N_9321,N_9998);
and U11222 (N_11222,N_8870,N_8223);
or U11223 (N_11223,N_9052,N_9012);
nand U11224 (N_11224,N_9896,N_9588);
or U11225 (N_11225,N_9511,N_9080);
nand U11226 (N_11226,N_8929,N_9229);
nor U11227 (N_11227,N_8628,N_8271);
or U11228 (N_11228,N_9393,N_8084);
nor U11229 (N_11229,N_9324,N_8400);
or U11230 (N_11230,N_8958,N_9249);
and U11231 (N_11231,N_8763,N_9295);
xnor U11232 (N_11232,N_8289,N_8119);
and U11233 (N_11233,N_9520,N_8893);
or U11234 (N_11234,N_8280,N_8858);
or U11235 (N_11235,N_8179,N_9338);
xor U11236 (N_11236,N_9088,N_9252);
nor U11237 (N_11237,N_8790,N_8544);
nand U11238 (N_11238,N_8875,N_8596);
nand U11239 (N_11239,N_8883,N_8562);
and U11240 (N_11240,N_8241,N_9859);
nand U11241 (N_11241,N_8461,N_8646);
and U11242 (N_11242,N_8213,N_9130);
and U11243 (N_11243,N_9307,N_9905);
nand U11244 (N_11244,N_8520,N_9788);
and U11245 (N_11245,N_9845,N_9061);
or U11246 (N_11246,N_9211,N_8826);
nand U11247 (N_11247,N_8892,N_8095);
nand U11248 (N_11248,N_8391,N_9777);
nand U11249 (N_11249,N_8924,N_8491);
and U11250 (N_11250,N_8387,N_8533);
nor U11251 (N_11251,N_8323,N_9379);
nand U11252 (N_11252,N_8635,N_9036);
nand U11253 (N_11253,N_8455,N_8927);
or U11254 (N_11254,N_8825,N_9691);
nand U11255 (N_11255,N_8186,N_8809);
and U11256 (N_11256,N_9819,N_8250);
or U11257 (N_11257,N_8648,N_9089);
and U11258 (N_11258,N_9444,N_8806);
and U11259 (N_11259,N_9900,N_8322);
xor U11260 (N_11260,N_8723,N_9495);
nor U11261 (N_11261,N_8543,N_8787);
nand U11262 (N_11262,N_9805,N_9991);
nor U11263 (N_11263,N_8475,N_9688);
nand U11264 (N_11264,N_8129,N_9680);
nand U11265 (N_11265,N_9651,N_9381);
and U11266 (N_11266,N_8384,N_8265);
nand U11267 (N_11267,N_9756,N_9311);
xor U11268 (N_11268,N_8531,N_9847);
nand U11269 (N_11269,N_9971,N_8568);
nor U11270 (N_11270,N_9159,N_8988);
and U11271 (N_11271,N_9179,N_9953);
and U11272 (N_11272,N_8568,N_9039);
and U11273 (N_11273,N_8495,N_9282);
nor U11274 (N_11274,N_9977,N_8793);
and U11275 (N_11275,N_9740,N_9084);
nand U11276 (N_11276,N_8994,N_8991);
nand U11277 (N_11277,N_9301,N_9182);
and U11278 (N_11278,N_9542,N_8894);
and U11279 (N_11279,N_8984,N_9941);
nand U11280 (N_11280,N_9794,N_9787);
nand U11281 (N_11281,N_8798,N_9132);
nand U11282 (N_11282,N_9901,N_9852);
or U11283 (N_11283,N_8654,N_8265);
or U11284 (N_11284,N_9711,N_9279);
nand U11285 (N_11285,N_8955,N_8075);
xnor U11286 (N_11286,N_8410,N_9181);
or U11287 (N_11287,N_9925,N_8877);
nand U11288 (N_11288,N_8176,N_9993);
xor U11289 (N_11289,N_8557,N_8332);
nand U11290 (N_11290,N_8193,N_9596);
nand U11291 (N_11291,N_9142,N_9877);
nand U11292 (N_11292,N_9994,N_9889);
nor U11293 (N_11293,N_9374,N_9903);
nand U11294 (N_11294,N_8082,N_8011);
nor U11295 (N_11295,N_9234,N_9985);
nand U11296 (N_11296,N_9317,N_8033);
nor U11297 (N_11297,N_8233,N_9860);
and U11298 (N_11298,N_8194,N_8218);
nor U11299 (N_11299,N_9467,N_8463);
nand U11300 (N_11300,N_8574,N_8610);
and U11301 (N_11301,N_8405,N_8830);
or U11302 (N_11302,N_8170,N_9088);
nand U11303 (N_11303,N_8137,N_8291);
and U11304 (N_11304,N_8780,N_8598);
and U11305 (N_11305,N_9882,N_8338);
nor U11306 (N_11306,N_9342,N_8109);
nand U11307 (N_11307,N_8320,N_9575);
nand U11308 (N_11308,N_8445,N_8928);
nand U11309 (N_11309,N_9678,N_8484);
or U11310 (N_11310,N_9104,N_8719);
nand U11311 (N_11311,N_8696,N_8849);
nand U11312 (N_11312,N_9568,N_8464);
xor U11313 (N_11313,N_8207,N_9135);
xnor U11314 (N_11314,N_9629,N_9736);
and U11315 (N_11315,N_8951,N_9696);
nand U11316 (N_11316,N_8744,N_8533);
and U11317 (N_11317,N_9269,N_8788);
nand U11318 (N_11318,N_8812,N_9755);
nor U11319 (N_11319,N_9350,N_8791);
nand U11320 (N_11320,N_8171,N_8702);
xor U11321 (N_11321,N_8470,N_8906);
or U11322 (N_11322,N_9601,N_9983);
xor U11323 (N_11323,N_9883,N_9148);
and U11324 (N_11324,N_9826,N_8649);
or U11325 (N_11325,N_8907,N_9811);
or U11326 (N_11326,N_9134,N_9750);
nor U11327 (N_11327,N_9926,N_9592);
xnor U11328 (N_11328,N_9048,N_8314);
nor U11329 (N_11329,N_9834,N_8847);
nand U11330 (N_11330,N_8585,N_9697);
nor U11331 (N_11331,N_8401,N_9604);
nand U11332 (N_11332,N_8444,N_8304);
xor U11333 (N_11333,N_8537,N_8565);
nand U11334 (N_11334,N_8639,N_8112);
nor U11335 (N_11335,N_9690,N_8633);
or U11336 (N_11336,N_9755,N_8495);
nor U11337 (N_11337,N_9562,N_8078);
nor U11338 (N_11338,N_8545,N_9387);
and U11339 (N_11339,N_9982,N_8152);
nor U11340 (N_11340,N_9416,N_9561);
and U11341 (N_11341,N_8132,N_8732);
and U11342 (N_11342,N_9905,N_9723);
nand U11343 (N_11343,N_8072,N_9804);
and U11344 (N_11344,N_9426,N_9139);
nor U11345 (N_11345,N_9586,N_8276);
nor U11346 (N_11346,N_8180,N_9325);
or U11347 (N_11347,N_8534,N_8678);
xor U11348 (N_11348,N_9765,N_9373);
or U11349 (N_11349,N_9340,N_9350);
and U11350 (N_11350,N_9187,N_8860);
nor U11351 (N_11351,N_9879,N_8693);
xor U11352 (N_11352,N_8308,N_8659);
or U11353 (N_11353,N_8079,N_8407);
or U11354 (N_11354,N_8901,N_8372);
and U11355 (N_11355,N_8019,N_9856);
nand U11356 (N_11356,N_9990,N_9377);
and U11357 (N_11357,N_8608,N_8840);
xor U11358 (N_11358,N_9958,N_9631);
nand U11359 (N_11359,N_8775,N_8706);
xnor U11360 (N_11360,N_9509,N_9951);
nor U11361 (N_11361,N_9884,N_9924);
or U11362 (N_11362,N_8722,N_9540);
nand U11363 (N_11363,N_8127,N_8070);
nor U11364 (N_11364,N_8165,N_8390);
and U11365 (N_11365,N_9359,N_8512);
nand U11366 (N_11366,N_8536,N_8625);
nand U11367 (N_11367,N_8440,N_9553);
nor U11368 (N_11368,N_8381,N_8228);
or U11369 (N_11369,N_9057,N_8843);
nand U11370 (N_11370,N_9690,N_9255);
nand U11371 (N_11371,N_8919,N_9412);
nand U11372 (N_11372,N_9245,N_9887);
xor U11373 (N_11373,N_9281,N_9890);
or U11374 (N_11374,N_8897,N_8508);
xor U11375 (N_11375,N_8476,N_8101);
and U11376 (N_11376,N_9514,N_8543);
nand U11377 (N_11377,N_9869,N_9512);
and U11378 (N_11378,N_9688,N_9072);
or U11379 (N_11379,N_8983,N_8029);
nor U11380 (N_11380,N_9531,N_8303);
or U11381 (N_11381,N_8473,N_8684);
or U11382 (N_11382,N_9758,N_8170);
and U11383 (N_11383,N_8402,N_8799);
nor U11384 (N_11384,N_8318,N_8663);
nand U11385 (N_11385,N_8251,N_8436);
or U11386 (N_11386,N_8045,N_8214);
or U11387 (N_11387,N_8691,N_8917);
xor U11388 (N_11388,N_9839,N_9631);
and U11389 (N_11389,N_8068,N_9989);
xor U11390 (N_11390,N_8605,N_8750);
and U11391 (N_11391,N_9473,N_9060);
and U11392 (N_11392,N_8444,N_9339);
nand U11393 (N_11393,N_8378,N_8197);
nand U11394 (N_11394,N_9714,N_9282);
or U11395 (N_11395,N_9528,N_9633);
and U11396 (N_11396,N_9320,N_8997);
nor U11397 (N_11397,N_8827,N_9164);
nor U11398 (N_11398,N_9926,N_8648);
and U11399 (N_11399,N_8676,N_9774);
and U11400 (N_11400,N_9438,N_8502);
nand U11401 (N_11401,N_8766,N_8824);
xnor U11402 (N_11402,N_9825,N_9833);
nor U11403 (N_11403,N_9408,N_9583);
nor U11404 (N_11404,N_8051,N_8828);
and U11405 (N_11405,N_9141,N_9017);
xnor U11406 (N_11406,N_8882,N_9339);
nand U11407 (N_11407,N_9389,N_9240);
nand U11408 (N_11408,N_8867,N_9028);
xor U11409 (N_11409,N_8131,N_8468);
nand U11410 (N_11410,N_8382,N_8218);
or U11411 (N_11411,N_9438,N_8385);
xor U11412 (N_11412,N_8672,N_8571);
and U11413 (N_11413,N_9047,N_9410);
xor U11414 (N_11414,N_8632,N_8742);
and U11415 (N_11415,N_8972,N_9823);
nor U11416 (N_11416,N_9311,N_8351);
nor U11417 (N_11417,N_8226,N_9639);
or U11418 (N_11418,N_8464,N_9353);
or U11419 (N_11419,N_9895,N_8263);
or U11420 (N_11420,N_8158,N_9819);
nand U11421 (N_11421,N_8284,N_8013);
and U11422 (N_11422,N_9955,N_9024);
or U11423 (N_11423,N_9753,N_8621);
nor U11424 (N_11424,N_8023,N_9933);
and U11425 (N_11425,N_8560,N_8014);
nand U11426 (N_11426,N_8283,N_8210);
nor U11427 (N_11427,N_8014,N_8258);
xnor U11428 (N_11428,N_8699,N_9113);
nor U11429 (N_11429,N_8382,N_9446);
nor U11430 (N_11430,N_8818,N_9784);
xor U11431 (N_11431,N_9606,N_9208);
xor U11432 (N_11432,N_8771,N_9448);
nand U11433 (N_11433,N_9824,N_9784);
and U11434 (N_11434,N_9170,N_9731);
and U11435 (N_11435,N_9863,N_9130);
nor U11436 (N_11436,N_8412,N_9091);
nor U11437 (N_11437,N_8122,N_9104);
xor U11438 (N_11438,N_8629,N_8358);
nor U11439 (N_11439,N_8061,N_9324);
and U11440 (N_11440,N_8074,N_9130);
xnor U11441 (N_11441,N_9540,N_9226);
xnor U11442 (N_11442,N_9923,N_8077);
or U11443 (N_11443,N_9807,N_8576);
nand U11444 (N_11444,N_9473,N_9375);
and U11445 (N_11445,N_9271,N_8414);
nor U11446 (N_11446,N_9829,N_9487);
nor U11447 (N_11447,N_8664,N_8016);
xnor U11448 (N_11448,N_8321,N_9964);
or U11449 (N_11449,N_9383,N_8775);
nand U11450 (N_11450,N_8123,N_9971);
nand U11451 (N_11451,N_8488,N_9092);
nand U11452 (N_11452,N_8929,N_9529);
or U11453 (N_11453,N_8797,N_8472);
or U11454 (N_11454,N_9286,N_9003);
or U11455 (N_11455,N_8402,N_8156);
nor U11456 (N_11456,N_8009,N_9836);
nor U11457 (N_11457,N_9928,N_8333);
nor U11458 (N_11458,N_8309,N_9977);
nand U11459 (N_11459,N_9911,N_9015);
or U11460 (N_11460,N_9833,N_9146);
or U11461 (N_11461,N_8152,N_8508);
xnor U11462 (N_11462,N_9222,N_8315);
nor U11463 (N_11463,N_9257,N_8017);
nor U11464 (N_11464,N_8264,N_8267);
or U11465 (N_11465,N_9146,N_9390);
nor U11466 (N_11466,N_8312,N_9771);
or U11467 (N_11467,N_8430,N_9223);
or U11468 (N_11468,N_8548,N_9804);
and U11469 (N_11469,N_8721,N_9447);
or U11470 (N_11470,N_9258,N_8550);
and U11471 (N_11471,N_9010,N_9965);
and U11472 (N_11472,N_8584,N_8324);
nor U11473 (N_11473,N_8177,N_9120);
or U11474 (N_11474,N_9845,N_8483);
nor U11475 (N_11475,N_8015,N_8564);
nand U11476 (N_11476,N_8898,N_9379);
and U11477 (N_11477,N_9501,N_9786);
or U11478 (N_11478,N_9567,N_8421);
and U11479 (N_11479,N_9875,N_8485);
and U11480 (N_11480,N_9076,N_9356);
and U11481 (N_11481,N_9663,N_8300);
nand U11482 (N_11482,N_9942,N_9285);
nor U11483 (N_11483,N_9424,N_9027);
nor U11484 (N_11484,N_8630,N_9599);
nand U11485 (N_11485,N_9284,N_9477);
or U11486 (N_11486,N_8165,N_9756);
xnor U11487 (N_11487,N_9824,N_9103);
nand U11488 (N_11488,N_9284,N_9272);
nand U11489 (N_11489,N_9813,N_9827);
xnor U11490 (N_11490,N_9243,N_9299);
or U11491 (N_11491,N_9765,N_9109);
and U11492 (N_11492,N_9920,N_9188);
or U11493 (N_11493,N_8740,N_9636);
nand U11494 (N_11494,N_8243,N_9838);
and U11495 (N_11495,N_9059,N_9175);
xnor U11496 (N_11496,N_9985,N_9945);
and U11497 (N_11497,N_9808,N_8219);
or U11498 (N_11498,N_9125,N_9334);
xor U11499 (N_11499,N_9810,N_8031);
or U11500 (N_11500,N_9699,N_8248);
nor U11501 (N_11501,N_8504,N_9615);
nand U11502 (N_11502,N_9916,N_8437);
nand U11503 (N_11503,N_9311,N_8049);
or U11504 (N_11504,N_8213,N_8951);
and U11505 (N_11505,N_9505,N_8663);
nand U11506 (N_11506,N_9468,N_9606);
nor U11507 (N_11507,N_8087,N_8207);
nor U11508 (N_11508,N_9687,N_8973);
and U11509 (N_11509,N_8599,N_8303);
or U11510 (N_11510,N_9556,N_9767);
and U11511 (N_11511,N_8724,N_8467);
nand U11512 (N_11512,N_8258,N_8301);
nor U11513 (N_11513,N_8232,N_8222);
xor U11514 (N_11514,N_8085,N_8878);
and U11515 (N_11515,N_8785,N_9178);
nor U11516 (N_11516,N_9841,N_8960);
nand U11517 (N_11517,N_9193,N_8270);
nor U11518 (N_11518,N_9251,N_9553);
and U11519 (N_11519,N_9704,N_8803);
nor U11520 (N_11520,N_8303,N_9868);
nor U11521 (N_11521,N_9982,N_9828);
nor U11522 (N_11522,N_9672,N_9283);
nor U11523 (N_11523,N_8360,N_8034);
and U11524 (N_11524,N_8227,N_8698);
nand U11525 (N_11525,N_8424,N_8552);
nand U11526 (N_11526,N_9680,N_8225);
or U11527 (N_11527,N_8095,N_8789);
or U11528 (N_11528,N_9959,N_9376);
or U11529 (N_11529,N_8860,N_9042);
nand U11530 (N_11530,N_9003,N_8560);
or U11531 (N_11531,N_8687,N_8543);
or U11532 (N_11532,N_8187,N_8593);
xnor U11533 (N_11533,N_9984,N_9237);
nor U11534 (N_11534,N_9185,N_9201);
and U11535 (N_11535,N_8060,N_8502);
and U11536 (N_11536,N_9881,N_9480);
nor U11537 (N_11537,N_8269,N_9039);
nand U11538 (N_11538,N_9221,N_8073);
and U11539 (N_11539,N_9708,N_9629);
or U11540 (N_11540,N_9628,N_8114);
nor U11541 (N_11541,N_8413,N_8637);
nand U11542 (N_11542,N_9868,N_8363);
or U11543 (N_11543,N_8935,N_9791);
nor U11544 (N_11544,N_9149,N_8935);
nand U11545 (N_11545,N_8372,N_8441);
xnor U11546 (N_11546,N_8579,N_8968);
nor U11547 (N_11547,N_8954,N_9751);
and U11548 (N_11548,N_8465,N_8895);
or U11549 (N_11549,N_8264,N_9832);
nand U11550 (N_11550,N_9413,N_9446);
and U11551 (N_11551,N_8892,N_8355);
and U11552 (N_11552,N_9806,N_9274);
nor U11553 (N_11553,N_8682,N_9547);
or U11554 (N_11554,N_8355,N_8931);
nand U11555 (N_11555,N_9006,N_8923);
and U11556 (N_11556,N_8059,N_8184);
or U11557 (N_11557,N_8182,N_9952);
xor U11558 (N_11558,N_9334,N_9957);
or U11559 (N_11559,N_8295,N_9551);
or U11560 (N_11560,N_8815,N_8854);
and U11561 (N_11561,N_9738,N_8024);
nor U11562 (N_11562,N_8650,N_9145);
or U11563 (N_11563,N_9240,N_8226);
or U11564 (N_11564,N_8333,N_8796);
or U11565 (N_11565,N_8347,N_8616);
nor U11566 (N_11566,N_8476,N_8326);
xnor U11567 (N_11567,N_8532,N_8181);
and U11568 (N_11568,N_8479,N_9161);
or U11569 (N_11569,N_9460,N_9708);
nor U11570 (N_11570,N_8988,N_9232);
nor U11571 (N_11571,N_8703,N_9036);
nand U11572 (N_11572,N_8908,N_9483);
and U11573 (N_11573,N_8149,N_9643);
nand U11574 (N_11574,N_9967,N_9588);
nand U11575 (N_11575,N_8953,N_8227);
xnor U11576 (N_11576,N_9517,N_9096);
or U11577 (N_11577,N_8061,N_8953);
nor U11578 (N_11578,N_9934,N_8726);
and U11579 (N_11579,N_9103,N_9899);
nor U11580 (N_11580,N_9166,N_8414);
and U11581 (N_11581,N_8768,N_8460);
or U11582 (N_11582,N_8573,N_9996);
and U11583 (N_11583,N_9717,N_9193);
nor U11584 (N_11584,N_8383,N_8801);
or U11585 (N_11585,N_8342,N_9140);
and U11586 (N_11586,N_9978,N_8014);
nor U11587 (N_11587,N_8784,N_9873);
nand U11588 (N_11588,N_9935,N_8798);
and U11589 (N_11589,N_8029,N_8879);
nor U11590 (N_11590,N_8914,N_9681);
or U11591 (N_11591,N_9995,N_8541);
or U11592 (N_11592,N_9195,N_9161);
and U11593 (N_11593,N_8000,N_9779);
nand U11594 (N_11594,N_8415,N_8487);
nand U11595 (N_11595,N_9690,N_9821);
xor U11596 (N_11596,N_8630,N_8018);
nor U11597 (N_11597,N_8550,N_9070);
nand U11598 (N_11598,N_9572,N_9583);
or U11599 (N_11599,N_8620,N_8362);
or U11600 (N_11600,N_8800,N_8937);
nand U11601 (N_11601,N_8479,N_8834);
nand U11602 (N_11602,N_8678,N_9777);
or U11603 (N_11603,N_9341,N_8550);
or U11604 (N_11604,N_9632,N_8864);
and U11605 (N_11605,N_9768,N_9643);
nor U11606 (N_11606,N_9998,N_8085);
and U11607 (N_11607,N_8771,N_9107);
nand U11608 (N_11608,N_9176,N_9209);
nand U11609 (N_11609,N_8690,N_8306);
and U11610 (N_11610,N_8467,N_8757);
or U11611 (N_11611,N_9632,N_9392);
nand U11612 (N_11612,N_8025,N_8503);
nand U11613 (N_11613,N_8463,N_8565);
nor U11614 (N_11614,N_9620,N_8325);
nor U11615 (N_11615,N_9676,N_9764);
or U11616 (N_11616,N_9083,N_8145);
nor U11617 (N_11617,N_9274,N_8183);
and U11618 (N_11618,N_8693,N_8562);
xor U11619 (N_11619,N_9874,N_9283);
or U11620 (N_11620,N_8229,N_8913);
nand U11621 (N_11621,N_8880,N_9557);
or U11622 (N_11622,N_8072,N_8578);
nand U11623 (N_11623,N_9743,N_8872);
and U11624 (N_11624,N_8589,N_9218);
or U11625 (N_11625,N_9322,N_9406);
nand U11626 (N_11626,N_8679,N_8156);
nor U11627 (N_11627,N_9027,N_8982);
nor U11628 (N_11628,N_9539,N_9572);
and U11629 (N_11629,N_9859,N_9061);
or U11630 (N_11630,N_8702,N_9862);
and U11631 (N_11631,N_8021,N_8664);
nand U11632 (N_11632,N_9257,N_9915);
and U11633 (N_11633,N_9848,N_9082);
nand U11634 (N_11634,N_9869,N_8202);
nand U11635 (N_11635,N_8571,N_8689);
or U11636 (N_11636,N_8288,N_8790);
xnor U11637 (N_11637,N_9169,N_9801);
or U11638 (N_11638,N_8118,N_9881);
or U11639 (N_11639,N_9163,N_8639);
or U11640 (N_11640,N_9540,N_9213);
and U11641 (N_11641,N_8176,N_9391);
nand U11642 (N_11642,N_8234,N_9300);
or U11643 (N_11643,N_9386,N_9609);
and U11644 (N_11644,N_9267,N_8690);
nand U11645 (N_11645,N_9760,N_9606);
nand U11646 (N_11646,N_8907,N_9731);
nor U11647 (N_11647,N_8837,N_8169);
xnor U11648 (N_11648,N_8159,N_8527);
xnor U11649 (N_11649,N_9061,N_8248);
or U11650 (N_11650,N_8154,N_8192);
nor U11651 (N_11651,N_8034,N_9459);
nand U11652 (N_11652,N_8326,N_9310);
nor U11653 (N_11653,N_8523,N_9576);
and U11654 (N_11654,N_9656,N_8164);
nor U11655 (N_11655,N_9133,N_8682);
nand U11656 (N_11656,N_8384,N_9290);
nand U11657 (N_11657,N_9988,N_8749);
xor U11658 (N_11658,N_8841,N_9572);
and U11659 (N_11659,N_8554,N_9734);
or U11660 (N_11660,N_9916,N_9694);
nand U11661 (N_11661,N_9543,N_8670);
and U11662 (N_11662,N_8929,N_8610);
or U11663 (N_11663,N_8772,N_8135);
xor U11664 (N_11664,N_8396,N_9238);
and U11665 (N_11665,N_8120,N_9213);
and U11666 (N_11666,N_9550,N_9188);
nor U11667 (N_11667,N_8021,N_8406);
xnor U11668 (N_11668,N_8200,N_9333);
or U11669 (N_11669,N_8912,N_9037);
and U11670 (N_11670,N_8865,N_9739);
nand U11671 (N_11671,N_8641,N_8658);
xnor U11672 (N_11672,N_8056,N_9973);
and U11673 (N_11673,N_9444,N_8981);
xnor U11674 (N_11674,N_9390,N_9958);
nor U11675 (N_11675,N_8855,N_9205);
or U11676 (N_11676,N_9125,N_9076);
nor U11677 (N_11677,N_9733,N_8014);
nand U11678 (N_11678,N_8415,N_8190);
or U11679 (N_11679,N_9914,N_9241);
nor U11680 (N_11680,N_9534,N_9511);
nand U11681 (N_11681,N_8549,N_9515);
nand U11682 (N_11682,N_9740,N_8095);
nor U11683 (N_11683,N_8353,N_8199);
or U11684 (N_11684,N_9440,N_8946);
or U11685 (N_11685,N_8832,N_9515);
and U11686 (N_11686,N_9382,N_9812);
nor U11687 (N_11687,N_8003,N_9029);
or U11688 (N_11688,N_9909,N_9618);
and U11689 (N_11689,N_9683,N_8946);
and U11690 (N_11690,N_8677,N_9327);
nor U11691 (N_11691,N_9294,N_8147);
and U11692 (N_11692,N_8905,N_9688);
or U11693 (N_11693,N_8593,N_9256);
nand U11694 (N_11694,N_9584,N_9393);
and U11695 (N_11695,N_9676,N_8875);
nor U11696 (N_11696,N_8575,N_8481);
or U11697 (N_11697,N_8918,N_9589);
nand U11698 (N_11698,N_8241,N_8958);
nand U11699 (N_11699,N_9407,N_8089);
and U11700 (N_11700,N_8425,N_9822);
or U11701 (N_11701,N_9636,N_8866);
nor U11702 (N_11702,N_8778,N_8718);
or U11703 (N_11703,N_9074,N_9558);
nand U11704 (N_11704,N_8887,N_9983);
nor U11705 (N_11705,N_8839,N_8051);
nor U11706 (N_11706,N_9231,N_8887);
nand U11707 (N_11707,N_9213,N_8217);
nor U11708 (N_11708,N_8320,N_8262);
nand U11709 (N_11709,N_8817,N_8070);
nor U11710 (N_11710,N_8949,N_9695);
nor U11711 (N_11711,N_9785,N_8821);
nor U11712 (N_11712,N_9568,N_9310);
xor U11713 (N_11713,N_8665,N_8629);
nand U11714 (N_11714,N_9150,N_8867);
and U11715 (N_11715,N_8694,N_9731);
nand U11716 (N_11716,N_9769,N_9476);
nor U11717 (N_11717,N_8041,N_9415);
nor U11718 (N_11718,N_8479,N_9796);
nand U11719 (N_11719,N_9207,N_8967);
and U11720 (N_11720,N_8249,N_8089);
and U11721 (N_11721,N_8475,N_9129);
or U11722 (N_11722,N_9862,N_8009);
and U11723 (N_11723,N_9782,N_8790);
nor U11724 (N_11724,N_8421,N_9625);
and U11725 (N_11725,N_9502,N_9500);
nand U11726 (N_11726,N_8742,N_8520);
xor U11727 (N_11727,N_9828,N_9291);
nand U11728 (N_11728,N_9725,N_8781);
nand U11729 (N_11729,N_9591,N_8408);
xnor U11730 (N_11730,N_9214,N_9351);
xnor U11731 (N_11731,N_8926,N_9350);
or U11732 (N_11732,N_8984,N_8903);
or U11733 (N_11733,N_8518,N_8509);
xor U11734 (N_11734,N_8896,N_8226);
and U11735 (N_11735,N_9949,N_8169);
and U11736 (N_11736,N_9084,N_8297);
nand U11737 (N_11737,N_8199,N_8882);
or U11738 (N_11738,N_9806,N_8724);
nand U11739 (N_11739,N_9921,N_9655);
nor U11740 (N_11740,N_8087,N_8564);
and U11741 (N_11741,N_9485,N_8467);
and U11742 (N_11742,N_9878,N_9202);
nor U11743 (N_11743,N_9867,N_8775);
nor U11744 (N_11744,N_8809,N_8481);
or U11745 (N_11745,N_9467,N_8809);
nand U11746 (N_11746,N_8154,N_9243);
nand U11747 (N_11747,N_8810,N_9085);
and U11748 (N_11748,N_9494,N_8200);
or U11749 (N_11749,N_8496,N_8786);
or U11750 (N_11750,N_9296,N_9136);
xnor U11751 (N_11751,N_9002,N_8568);
and U11752 (N_11752,N_9694,N_9030);
or U11753 (N_11753,N_8649,N_8579);
nand U11754 (N_11754,N_8687,N_8452);
nor U11755 (N_11755,N_8294,N_9577);
nor U11756 (N_11756,N_9991,N_9308);
nand U11757 (N_11757,N_8409,N_8792);
or U11758 (N_11758,N_9161,N_9932);
nand U11759 (N_11759,N_8802,N_8236);
and U11760 (N_11760,N_8167,N_9210);
nor U11761 (N_11761,N_8676,N_8915);
nand U11762 (N_11762,N_8936,N_8854);
nand U11763 (N_11763,N_9845,N_9252);
nand U11764 (N_11764,N_8155,N_9766);
xnor U11765 (N_11765,N_9306,N_9590);
nand U11766 (N_11766,N_9147,N_9676);
nand U11767 (N_11767,N_8832,N_8148);
nor U11768 (N_11768,N_9445,N_9887);
nand U11769 (N_11769,N_8736,N_8561);
nand U11770 (N_11770,N_9579,N_9232);
nor U11771 (N_11771,N_8815,N_8270);
or U11772 (N_11772,N_9406,N_9293);
nand U11773 (N_11773,N_8086,N_8315);
or U11774 (N_11774,N_8050,N_8641);
xor U11775 (N_11775,N_9466,N_9282);
or U11776 (N_11776,N_9816,N_9721);
nand U11777 (N_11777,N_9570,N_8388);
and U11778 (N_11778,N_8528,N_8402);
and U11779 (N_11779,N_9348,N_8224);
or U11780 (N_11780,N_9120,N_9344);
and U11781 (N_11781,N_8191,N_8168);
nor U11782 (N_11782,N_8868,N_8720);
xor U11783 (N_11783,N_9958,N_8808);
nor U11784 (N_11784,N_8337,N_9203);
or U11785 (N_11785,N_8162,N_8057);
xor U11786 (N_11786,N_9077,N_8870);
nand U11787 (N_11787,N_8633,N_8142);
nor U11788 (N_11788,N_9145,N_9937);
xnor U11789 (N_11789,N_9776,N_8256);
and U11790 (N_11790,N_9571,N_9193);
nand U11791 (N_11791,N_8802,N_8642);
nor U11792 (N_11792,N_8808,N_8591);
or U11793 (N_11793,N_8245,N_9151);
or U11794 (N_11794,N_8994,N_9707);
nand U11795 (N_11795,N_8572,N_8008);
or U11796 (N_11796,N_8456,N_9787);
nand U11797 (N_11797,N_9398,N_9700);
nand U11798 (N_11798,N_9211,N_8935);
xnor U11799 (N_11799,N_9688,N_8015);
and U11800 (N_11800,N_8376,N_8855);
and U11801 (N_11801,N_8715,N_9230);
and U11802 (N_11802,N_8338,N_8031);
and U11803 (N_11803,N_8008,N_8273);
and U11804 (N_11804,N_8713,N_8021);
or U11805 (N_11805,N_8238,N_8588);
nand U11806 (N_11806,N_8805,N_8564);
or U11807 (N_11807,N_8076,N_9824);
nand U11808 (N_11808,N_8919,N_8179);
nand U11809 (N_11809,N_8185,N_9611);
and U11810 (N_11810,N_8226,N_8773);
nor U11811 (N_11811,N_9284,N_8789);
nor U11812 (N_11812,N_9607,N_9456);
nand U11813 (N_11813,N_9084,N_8463);
and U11814 (N_11814,N_8685,N_8480);
and U11815 (N_11815,N_8846,N_8731);
xnor U11816 (N_11816,N_8282,N_9086);
and U11817 (N_11817,N_9476,N_8086);
nor U11818 (N_11818,N_8746,N_8265);
or U11819 (N_11819,N_9006,N_9205);
or U11820 (N_11820,N_8179,N_8467);
nand U11821 (N_11821,N_8056,N_8865);
or U11822 (N_11822,N_8359,N_9130);
or U11823 (N_11823,N_9669,N_8640);
or U11824 (N_11824,N_9883,N_8800);
and U11825 (N_11825,N_9441,N_9750);
or U11826 (N_11826,N_8900,N_9208);
nor U11827 (N_11827,N_8301,N_9264);
or U11828 (N_11828,N_9414,N_9189);
xor U11829 (N_11829,N_9933,N_9379);
nand U11830 (N_11830,N_8137,N_8404);
nand U11831 (N_11831,N_8755,N_8371);
and U11832 (N_11832,N_9779,N_9776);
nand U11833 (N_11833,N_8309,N_9536);
nor U11834 (N_11834,N_9118,N_9469);
nor U11835 (N_11835,N_8957,N_8890);
or U11836 (N_11836,N_9619,N_8752);
nand U11837 (N_11837,N_9240,N_9557);
nand U11838 (N_11838,N_8017,N_8400);
nor U11839 (N_11839,N_8972,N_8199);
or U11840 (N_11840,N_8096,N_9467);
nor U11841 (N_11841,N_9426,N_8764);
and U11842 (N_11842,N_9963,N_8314);
or U11843 (N_11843,N_8462,N_9022);
and U11844 (N_11844,N_9331,N_8515);
and U11845 (N_11845,N_8542,N_9512);
xnor U11846 (N_11846,N_9805,N_8139);
or U11847 (N_11847,N_9608,N_8731);
and U11848 (N_11848,N_9319,N_8358);
xnor U11849 (N_11849,N_8139,N_9499);
and U11850 (N_11850,N_9613,N_9721);
xor U11851 (N_11851,N_8663,N_9611);
or U11852 (N_11852,N_9685,N_9414);
nand U11853 (N_11853,N_9236,N_8807);
and U11854 (N_11854,N_8624,N_8718);
nor U11855 (N_11855,N_8681,N_8508);
nor U11856 (N_11856,N_9255,N_8574);
and U11857 (N_11857,N_8818,N_8440);
nor U11858 (N_11858,N_9119,N_9096);
and U11859 (N_11859,N_9549,N_8147);
xnor U11860 (N_11860,N_8928,N_9213);
and U11861 (N_11861,N_9445,N_9973);
nor U11862 (N_11862,N_9317,N_9261);
or U11863 (N_11863,N_9629,N_9038);
nand U11864 (N_11864,N_9785,N_9862);
and U11865 (N_11865,N_8750,N_9718);
nor U11866 (N_11866,N_8845,N_9159);
nand U11867 (N_11867,N_8367,N_9740);
nor U11868 (N_11868,N_9081,N_9214);
or U11869 (N_11869,N_9871,N_8263);
and U11870 (N_11870,N_8160,N_8960);
and U11871 (N_11871,N_8113,N_9031);
nor U11872 (N_11872,N_9569,N_9748);
xnor U11873 (N_11873,N_8929,N_9770);
nand U11874 (N_11874,N_9539,N_9883);
and U11875 (N_11875,N_8243,N_9121);
or U11876 (N_11876,N_8737,N_9819);
and U11877 (N_11877,N_8385,N_8408);
nand U11878 (N_11878,N_9873,N_8600);
and U11879 (N_11879,N_9295,N_8573);
or U11880 (N_11880,N_8141,N_9414);
and U11881 (N_11881,N_9775,N_9184);
xor U11882 (N_11882,N_9392,N_9333);
and U11883 (N_11883,N_8836,N_9313);
and U11884 (N_11884,N_9733,N_9374);
or U11885 (N_11885,N_8327,N_9051);
or U11886 (N_11886,N_8119,N_8124);
xor U11887 (N_11887,N_8666,N_8341);
nand U11888 (N_11888,N_8096,N_8496);
nor U11889 (N_11889,N_8764,N_8329);
nor U11890 (N_11890,N_9214,N_8937);
or U11891 (N_11891,N_8087,N_9607);
nor U11892 (N_11892,N_9694,N_9003);
and U11893 (N_11893,N_8458,N_9744);
nand U11894 (N_11894,N_8402,N_8898);
nand U11895 (N_11895,N_9304,N_9725);
nand U11896 (N_11896,N_8393,N_9450);
or U11897 (N_11897,N_9361,N_9259);
and U11898 (N_11898,N_9397,N_9593);
or U11899 (N_11899,N_8956,N_8785);
xnor U11900 (N_11900,N_9545,N_8223);
and U11901 (N_11901,N_8487,N_8958);
and U11902 (N_11902,N_8347,N_9672);
xnor U11903 (N_11903,N_9123,N_9489);
or U11904 (N_11904,N_9448,N_9476);
nand U11905 (N_11905,N_9425,N_8733);
nor U11906 (N_11906,N_8036,N_8810);
nand U11907 (N_11907,N_8584,N_8685);
xor U11908 (N_11908,N_9317,N_8338);
nor U11909 (N_11909,N_9693,N_9027);
or U11910 (N_11910,N_9358,N_9536);
and U11911 (N_11911,N_9298,N_8754);
or U11912 (N_11912,N_9574,N_8517);
nor U11913 (N_11913,N_9151,N_9960);
nor U11914 (N_11914,N_9141,N_8510);
nand U11915 (N_11915,N_8304,N_8880);
nand U11916 (N_11916,N_9151,N_9002);
or U11917 (N_11917,N_8444,N_9769);
and U11918 (N_11918,N_9659,N_9056);
nand U11919 (N_11919,N_9947,N_8654);
and U11920 (N_11920,N_9759,N_8342);
nand U11921 (N_11921,N_9935,N_9354);
or U11922 (N_11922,N_8696,N_8822);
or U11923 (N_11923,N_9069,N_9648);
nor U11924 (N_11924,N_8401,N_8237);
nand U11925 (N_11925,N_9955,N_9609);
or U11926 (N_11926,N_8014,N_9562);
and U11927 (N_11927,N_9834,N_9146);
or U11928 (N_11928,N_8853,N_8688);
nor U11929 (N_11929,N_8657,N_9524);
and U11930 (N_11930,N_9460,N_9868);
nand U11931 (N_11931,N_9718,N_8648);
or U11932 (N_11932,N_8518,N_9477);
or U11933 (N_11933,N_8370,N_8939);
and U11934 (N_11934,N_9627,N_8920);
nand U11935 (N_11935,N_8896,N_8209);
or U11936 (N_11936,N_9650,N_9934);
and U11937 (N_11937,N_8848,N_8608);
nand U11938 (N_11938,N_8587,N_9952);
and U11939 (N_11939,N_9093,N_9760);
and U11940 (N_11940,N_9083,N_8040);
and U11941 (N_11941,N_8988,N_8052);
nand U11942 (N_11942,N_8120,N_9007);
nor U11943 (N_11943,N_9778,N_8709);
and U11944 (N_11944,N_8246,N_8567);
or U11945 (N_11945,N_8526,N_9631);
or U11946 (N_11946,N_8344,N_8096);
nor U11947 (N_11947,N_8962,N_8960);
nor U11948 (N_11948,N_8712,N_8888);
and U11949 (N_11949,N_9907,N_9523);
xor U11950 (N_11950,N_8428,N_8652);
or U11951 (N_11951,N_9744,N_8494);
nor U11952 (N_11952,N_8826,N_9849);
nand U11953 (N_11953,N_8364,N_8430);
nor U11954 (N_11954,N_8990,N_8119);
and U11955 (N_11955,N_8076,N_8693);
nor U11956 (N_11956,N_8841,N_9480);
xor U11957 (N_11957,N_8886,N_9644);
nand U11958 (N_11958,N_8916,N_9039);
nand U11959 (N_11959,N_8686,N_9561);
and U11960 (N_11960,N_9682,N_9855);
nor U11961 (N_11961,N_9092,N_8609);
or U11962 (N_11962,N_9169,N_9790);
and U11963 (N_11963,N_8923,N_8557);
xor U11964 (N_11964,N_9207,N_8349);
nand U11965 (N_11965,N_9520,N_9395);
and U11966 (N_11966,N_9037,N_8769);
nand U11967 (N_11967,N_8053,N_9063);
and U11968 (N_11968,N_8324,N_9959);
nand U11969 (N_11969,N_9174,N_9675);
or U11970 (N_11970,N_8092,N_8718);
nor U11971 (N_11971,N_8901,N_8505);
xor U11972 (N_11972,N_8664,N_9818);
xnor U11973 (N_11973,N_8552,N_9058);
and U11974 (N_11974,N_9492,N_8210);
nor U11975 (N_11975,N_8213,N_9965);
nor U11976 (N_11976,N_9076,N_9622);
or U11977 (N_11977,N_9010,N_9387);
and U11978 (N_11978,N_9245,N_8083);
and U11979 (N_11979,N_8961,N_9204);
or U11980 (N_11980,N_8746,N_8687);
or U11981 (N_11981,N_8027,N_8613);
nor U11982 (N_11982,N_8380,N_9953);
or U11983 (N_11983,N_8625,N_8840);
and U11984 (N_11984,N_9540,N_8977);
nand U11985 (N_11985,N_9517,N_8150);
nor U11986 (N_11986,N_8510,N_8237);
xnor U11987 (N_11987,N_9786,N_8080);
xor U11988 (N_11988,N_8315,N_8702);
and U11989 (N_11989,N_9787,N_9428);
xor U11990 (N_11990,N_9236,N_9063);
and U11991 (N_11991,N_8923,N_8949);
nand U11992 (N_11992,N_8503,N_9799);
nor U11993 (N_11993,N_8507,N_9846);
and U11994 (N_11994,N_9228,N_8904);
nor U11995 (N_11995,N_9012,N_8850);
nor U11996 (N_11996,N_9676,N_9718);
and U11997 (N_11997,N_9222,N_8678);
and U11998 (N_11998,N_8179,N_9358);
nor U11999 (N_11999,N_8977,N_8688);
or U12000 (N_12000,N_11057,N_10307);
and U12001 (N_12001,N_10198,N_11977);
or U12002 (N_12002,N_10124,N_10757);
or U12003 (N_12003,N_10143,N_11855);
xnor U12004 (N_12004,N_10554,N_11759);
and U12005 (N_12005,N_11271,N_10519);
or U12006 (N_12006,N_10684,N_10718);
or U12007 (N_12007,N_11648,N_10789);
and U12008 (N_12008,N_11177,N_10831);
nor U12009 (N_12009,N_11085,N_10913);
or U12010 (N_12010,N_10362,N_11055);
or U12011 (N_12011,N_10155,N_10353);
or U12012 (N_12012,N_10580,N_10659);
nor U12013 (N_12013,N_11416,N_10807);
or U12014 (N_12014,N_11273,N_10295);
and U12015 (N_12015,N_10989,N_11432);
and U12016 (N_12016,N_11487,N_10020);
or U12017 (N_12017,N_11638,N_10907);
xor U12018 (N_12018,N_10582,N_11375);
or U12019 (N_12019,N_10071,N_11576);
xor U12020 (N_12020,N_10107,N_11369);
nand U12021 (N_12021,N_11431,N_11357);
nand U12022 (N_12022,N_10940,N_11260);
xnor U12023 (N_12023,N_11790,N_10568);
and U12024 (N_12024,N_11578,N_10541);
or U12025 (N_12025,N_10750,N_11249);
or U12026 (N_12026,N_10524,N_10841);
nor U12027 (N_12027,N_11595,N_10533);
and U12028 (N_12028,N_10591,N_11963);
nand U12029 (N_12029,N_11799,N_10236);
or U12030 (N_12030,N_11291,N_11450);
xor U12031 (N_12031,N_10438,N_11142);
or U12032 (N_12032,N_10678,N_11969);
or U12033 (N_12033,N_10603,N_11635);
or U12034 (N_12034,N_11179,N_11437);
or U12035 (N_12035,N_10391,N_10703);
nor U12036 (N_12036,N_10178,N_11840);
nor U12037 (N_12037,N_10129,N_10402);
or U12038 (N_12038,N_11694,N_11022);
and U12039 (N_12039,N_10886,N_10139);
nor U12040 (N_12040,N_10982,N_10947);
and U12041 (N_12041,N_10288,N_10112);
or U12042 (N_12042,N_10342,N_10070);
and U12043 (N_12043,N_10826,N_10447);
nor U12044 (N_12044,N_11723,N_10200);
or U12045 (N_12045,N_11901,N_11821);
nand U12046 (N_12046,N_10276,N_11607);
nand U12047 (N_12047,N_11151,N_10688);
nor U12048 (N_12048,N_10279,N_10556);
xnor U12049 (N_12049,N_10477,N_11929);
nand U12050 (N_12050,N_11567,N_11039);
xor U12051 (N_12051,N_11299,N_11615);
or U12052 (N_12052,N_11767,N_11154);
nor U12053 (N_12053,N_10961,N_11235);
and U12054 (N_12054,N_11938,N_10332);
and U12055 (N_12055,N_11110,N_11372);
or U12056 (N_12056,N_10535,N_10371);
xor U12057 (N_12057,N_11051,N_10460);
nand U12058 (N_12058,N_11321,N_10270);
or U12059 (N_12059,N_11424,N_11362);
nand U12060 (N_12060,N_11891,N_10555);
or U12061 (N_12061,N_11931,N_10510);
nand U12062 (N_12062,N_11572,N_11330);
and U12063 (N_12063,N_11477,N_11614);
nor U12064 (N_12064,N_11666,N_10457);
or U12065 (N_12065,N_10628,N_11124);
or U12066 (N_12066,N_11965,N_11016);
nor U12067 (N_12067,N_10927,N_10946);
or U12068 (N_12068,N_11031,N_10220);
nor U12069 (N_12069,N_11811,N_11053);
and U12070 (N_12070,N_11815,N_11158);
and U12071 (N_12071,N_10280,N_11854);
nand U12072 (N_12072,N_10880,N_11003);
nor U12073 (N_12073,N_10035,N_11128);
or U12074 (N_12074,N_11405,N_10861);
xor U12075 (N_12075,N_11558,N_11297);
and U12076 (N_12076,N_10045,N_11820);
nor U12077 (N_12077,N_11400,N_10671);
xor U12078 (N_12078,N_10316,N_11033);
or U12079 (N_12079,N_10238,N_11340);
nand U12080 (N_12080,N_11955,N_10047);
xor U12081 (N_12081,N_11217,N_11908);
xor U12082 (N_12082,N_11333,N_11398);
nor U12083 (N_12083,N_11867,N_10144);
or U12084 (N_12084,N_10804,N_11494);
and U12085 (N_12085,N_10121,N_11749);
nor U12086 (N_12086,N_11066,N_11134);
nor U12087 (N_12087,N_11845,N_10657);
and U12088 (N_12088,N_10627,N_11644);
and U12089 (N_12089,N_11014,N_11436);
xor U12090 (N_12090,N_11247,N_11900);
or U12091 (N_12091,N_11018,N_11417);
or U12092 (N_12092,N_11985,N_11643);
or U12093 (N_12093,N_10529,N_10237);
and U12094 (N_12094,N_10226,N_10690);
nand U12095 (N_12095,N_11780,N_10348);
nor U12096 (N_12096,N_10889,N_11443);
or U12097 (N_12097,N_11859,N_10354);
or U12098 (N_12098,N_11990,N_10409);
nand U12099 (N_12099,N_10747,N_11132);
or U12100 (N_12100,N_10836,N_11603);
or U12101 (N_12101,N_11569,N_10984);
and U12102 (N_12102,N_11947,N_11617);
nand U12103 (N_12103,N_10383,N_10944);
and U12104 (N_12104,N_10033,N_10255);
xor U12105 (N_12105,N_10487,N_11981);
nand U12106 (N_12106,N_10746,N_10285);
nor U12107 (N_12107,N_11175,N_11233);
nand U12108 (N_12108,N_11789,N_11478);
or U12109 (N_12109,N_10859,N_10735);
nand U12110 (N_12110,N_10164,N_10515);
nor U12111 (N_12111,N_11147,N_11756);
nor U12112 (N_12112,N_10513,N_10117);
nor U12113 (N_12113,N_11211,N_11757);
or U12114 (N_12114,N_11536,N_10796);
nor U12115 (N_12115,N_10897,N_11633);
nor U12116 (N_12116,N_11078,N_10719);
xnor U12117 (N_12117,N_11314,N_11256);
and U12118 (N_12118,N_10809,N_10570);
nor U12119 (N_12119,N_11565,N_11678);
or U12120 (N_12120,N_10565,N_10429);
nand U12121 (N_12121,N_10712,N_11852);
and U12122 (N_12122,N_10720,N_11866);
nor U12123 (N_12123,N_11887,N_10916);
or U12124 (N_12124,N_10123,N_11924);
nor U12125 (N_12125,N_10620,N_10197);
and U12126 (N_12126,N_11302,N_10617);
nor U12127 (N_12127,N_11323,N_11542);
nand U12128 (N_12128,N_10733,N_10079);
and U12129 (N_12129,N_11038,N_11117);
and U12130 (N_12130,N_10730,N_10267);
or U12131 (N_12131,N_11379,N_10227);
nor U12132 (N_12132,N_10928,N_11155);
and U12133 (N_12133,N_10782,N_11104);
and U12134 (N_12134,N_10325,N_11539);
nand U12135 (N_12135,N_10970,N_10393);
and U12136 (N_12136,N_11704,N_10985);
xnor U12137 (N_12137,N_10696,N_11360);
and U12138 (N_12138,N_10711,N_10856);
nand U12139 (N_12139,N_10969,N_11428);
or U12140 (N_12140,N_10797,N_11515);
nor U12141 (N_12141,N_10708,N_11706);
or U12142 (N_12142,N_10072,N_10781);
nand U12143 (N_12143,N_11619,N_11599);
or U12144 (N_12144,N_11708,N_11500);
or U12145 (N_12145,N_11185,N_11309);
or U12146 (N_12146,N_10081,N_10243);
or U12147 (N_12147,N_10208,N_11327);
and U12148 (N_12148,N_10206,N_11623);
xnor U12149 (N_12149,N_11504,N_10752);
nor U12150 (N_12150,N_11153,N_10006);
or U12151 (N_12151,N_11592,N_10874);
nand U12152 (N_12152,N_11994,N_11277);
xor U12153 (N_12153,N_11168,N_10026);
nor U12154 (N_12154,N_10211,N_11076);
or U12155 (N_12155,N_11115,N_11471);
nand U12156 (N_12156,N_10249,N_11371);
and U12157 (N_12157,N_10359,N_10472);
nand U12158 (N_12158,N_11349,N_11946);
nor U12159 (N_12159,N_10415,N_11892);
and U12160 (N_12160,N_10250,N_11807);
or U12161 (N_12161,N_10904,N_10667);
nand U12162 (N_12162,N_11752,N_11758);
nand U12163 (N_12163,N_11498,N_10394);
or U12164 (N_12164,N_10286,N_10225);
and U12165 (N_12165,N_11998,N_10839);
nand U12166 (N_12166,N_10537,N_11012);
nand U12167 (N_12167,N_11102,N_10287);
and U12168 (N_12168,N_11517,N_10099);
nand U12169 (N_12169,N_11293,N_10215);
nand U12170 (N_12170,N_11275,N_11835);
nand U12171 (N_12171,N_11329,N_11916);
nand U12172 (N_12172,N_10210,N_11594);
nor U12173 (N_12173,N_10526,N_11518);
nor U12174 (N_12174,N_11566,N_11419);
nor U12175 (N_12175,N_11103,N_11898);
and U12176 (N_12176,N_10068,N_11992);
xor U12177 (N_12177,N_11818,N_11943);
xnor U12178 (N_12178,N_10523,N_11606);
nor U12179 (N_12179,N_11143,N_11034);
and U12180 (N_12180,N_10942,N_11501);
nand U12181 (N_12181,N_10340,N_11087);
nand U12182 (N_12182,N_10194,N_11182);
and U12183 (N_12183,N_11831,N_10245);
nor U12184 (N_12184,N_10407,N_10512);
and U12185 (N_12185,N_11773,N_10320);
and U12186 (N_12186,N_10461,N_11686);
nor U12187 (N_12187,N_11020,N_11363);
nand U12188 (N_12188,N_10374,N_10064);
and U12189 (N_12189,N_11396,N_11320);
nor U12190 (N_12190,N_10190,N_11681);
xor U12191 (N_12191,N_10221,N_10543);
nor U12192 (N_12192,N_10837,N_11839);
and U12193 (N_12193,N_10080,N_10097);
xnor U12194 (N_12194,N_10191,N_11613);
nand U12195 (N_12195,N_11195,N_11094);
or U12196 (N_12196,N_10488,N_10468);
xor U12197 (N_12197,N_10793,N_10399);
nor U12198 (N_12198,N_10873,N_11380);
nand U12199 (N_12199,N_10875,N_11364);
nand U12200 (N_12200,N_11684,N_10008);
or U12201 (N_12201,N_11524,N_11526);
nand U12202 (N_12202,N_10025,N_11863);
and U12203 (N_12203,N_11670,N_11682);
nor U12204 (N_12204,N_11171,N_11007);
or U12205 (N_12205,N_11342,N_11761);
nor U12206 (N_12206,N_11928,N_11527);
nor U12207 (N_12207,N_11118,N_10644);
nor U12208 (N_12208,N_10971,N_10308);
nand U12209 (N_12209,N_11590,N_10061);
xor U12210 (N_12210,N_11438,N_10923);
nor U12211 (N_12211,N_11145,N_11921);
or U12212 (N_12212,N_11164,N_10378);
nor U12213 (N_12213,N_10972,N_11934);
xnor U12214 (N_12214,N_11434,N_11668);
and U12215 (N_12215,N_10974,N_10222);
nand U12216 (N_12216,N_10436,N_11841);
nor U12217 (N_12217,N_11230,N_11970);
and U12218 (N_12218,N_11389,N_11152);
or U12219 (N_12219,N_11165,N_10463);
xnor U12220 (N_12220,N_10478,N_10729);
nor U12221 (N_12221,N_10404,N_11049);
or U12222 (N_12222,N_10410,N_11625);
and U12223 (N_12223,N_11750,N_11167);
and U12224 (N_12224,N_10187,N_10023);
nand U12225 (N_12225,N_11475,N_11785);
and U12226 (N_12226,N_11736,N_10709);
nor U12227 (N_12227,N_11203,N_11865);
and U12228 (N_12228,N_10586,N_11192);
or U12229 (N_12229,N_10778,N_10952);
nor U12230 (N_12230,N_11199,N_10284);
and U12231 (N_12231,N_11589,N_10103);
nor U12232 (N_12232,N_11043,N_10790);
or U12233 (N_12233,N_11975,N_10057);
xor U12234 (N_12234,N_10858,N_10772);
nor U12235 (N_12235,N_11739,N_10737);
and U12236 (N_12236,N_10828,N_10558);
nand U12237 (N_12237,N_10611,N_10085);
and U12238 (N_12238,N_11229,N_10993);
nand U12239 (N_12239,N_11538,N_11131);
and U12240 (N_12240,N_10815,N_11429);
and U12241 (N_12241,N_11506,N_10188);
or U12242 (N_12242,N_11270,N_11516);
nor U12243 (N_12243,N_10502,N_10641);
and U12244 (N_12244,N_11657,N_11244);
and U12245 (N_12245,N_11243,N_10967);
and U12246 (N_12246,N_11189,N_11317);
nand U12247 (N_12247,N_10717,N_11976);
or U12248 (N_12248,N_10264,N_10494);
nor U12249 (N_12249,N_10614,N_10384);
or U12250 (N_12250,N_10697,N_10365);
nand U12251 (N_12251,N_10744,N_11056);
nor U12252 (N_12252,N_10847,N_11246);
nor U12253 (N_12253,N_10299,N_11927);
nor U12254 (N_12254,N_10029,N_10086);
nand U12255 (N_12255,N_11359,N_11482);
and U12256 (N_12256,N_10272,N_11126);
or U12257 (N_12257,N_10496,N_10321);
nand U12258 (N_12258,N_10664,N_10028);
and U12259 (N_12259,N_11505,N_10643);
or U12260 (N_12260,N_10727,N_11522);
nand U12261 (N_12261,N_10052,N_10491);
and U12262 (N_12262,N_11925,N_10323);
nand U12263 (N_12263,N_11186,N_11048);
xor U12264 (N_12264,N_11441,N_10981);
nand U12265 (N_12265,N_10375,N_10260);
nor U12266 (N_12266,N_11746,N_11663);
or U12267 (N_12267,N_11823,N_11298);
and U12268 (N_12268,N_11307,N_10649);
nor U12269 (N_12269,N_10917,N_10334);
xnor U12270 (N_12270,N_10991,N_11322);
xnor U12271 (N_12271,N_10469,N_10030);
or U12272 (N_12272,N_11774,N_10193);
nand U12273 (N_12273,N_11356,N_10497);
and U12274 (N_12274,N_11305,N_10443);
nand U12275 (N_12275,N_11107,N_11991);
nor U12276 (N_12276,N_10360,N_10180);
nand U12277 (N_12277,N_11226,N_11959);
or U12278 (N_12278,N_10403,N_10130);
or U12279 (N_12279,N_11543,N_11046);
nand U12280 (N_12280,N_11636,N_10352);
nand U12281 (N_12281,N_10256,N_10743);
or U12282 (N_12282,N_11768,N_11824);
or U12283 (N_12283,N_11352,N_10585);
xor U12284 (N_12284,N_11618,N_11529);
and U12285 (N_12285,N_11328,N_10559);
or U12286 (N_12286,N_11219,N_10564);
xnor U12287 (N_12287,N_10723,N_11265);
nor U12288 (N_12288,N_11637,N_10486);
nor U12289 (N_12289,N_10275,N_11989);
and U12290 (N_12290,N_10763,N_10003);
nand U12291 (N_12291,N_10682,N_11878);
nand U12292 (N_12292,N_11097,N_11499);
or U12293 (N_12293,N_11125,N_11546);
xor U12294 (N_12294,N_10373,N_10036);
nor U12295 (N_12295,N_10490,N_10557);
nor U12296 (N_12296,N_11802,N_11972);
and U12297 (N_12297,N_11162,N_11907);
and U12298 (N_12298,N_10808,N_10259);
nand U12299 (N_12299,N_10231,N_11098);
nor U12300 (N_12300,N_11747,N_10715);
xnor U12301 (N_12301,N_11528,N_10336);
and U12302 (N_12302,N_10271,N_11806);
nor U12303 (N_12303,N_10201,N_11090);
nor U12304 (N_12304,N_10514,N_10310);
nand U12305 (N_12305,N_10141,N_11464);
and U12306 (N_12306,N_11880,N_11764);
or U12307 (N_12307,N_11511,N_10364);
xor U12308 (N_12308,N_10329,N_11279);
nor U12309 (N_12309,N_10566,N_10522);
or U12310 (N_12310,N_11734,N_10309);
or U12311 (N_12311,N_11609,N_11770);
and U12312 (N_12312,N_10199,N_11897);
xnor U12313 (N_12313,N_11601,N_11571);
and U12314 (N_12314,N_10157,N_11540);
nor U12315 (N_12315,N_11718,N_11267);
or U12316 (N_12316,N_11480,N_11714);
or U12317 (N_12317,N_10076,N_11936);
and U12318 (N_12318,N_11187,N_11732);
nand U12319 (N_12319,N_11894,N_11748);
xnor U12320 (N_12320,N_11913,N_10986);
or U12321 (N_12321,N_11476,N_11549);
or U12322 (N_12322,N_11062,N_11705);
or U12323 (N_12323,N_10749,N_11367);
nand U12324 (N_12324,N_10593,N_10319);
nor U12325 (N_12325,N_10925,N_11075);
and U12326 (N_12326,N_10297,N_11047);
or U12327 (N_12327,N_11719,N_10060);
or U12328 (N_12328,N_10527,N_11435);
nor U12329 (N_12329,N_10294,N_11834);
or U12330 (N_12330,N_10000,N_11312);
and U12331 (N_12331,N_10435,N_11030);
nand U12332 (N_12332,N_11479,N_11709);
xnor U12333 (N_12333,N_10093,N_11069);
or U12334 (N_12334,N_11001,N_11035);
and U12335 (N_12335,N_10918,N_10694);
or U12336 (N_12336,N_10864,N_10638);
and U12337 (N_12337,N_10784,N_11639);
nand U12338 (N_12338,N_10854,N_11338);
or U12339 (N_12339,N_10058,N_10964);
xnor U12340 (N_12340,N_10170,N_10168);
and U12341 (N_12341,N_11337,N_10055);
and U12342 (N_12342,N_11582,N_10147);
nand U12343 (N_12343,N_10296,N_11227);
nor U12344 (N_12344,N_10174,N_10933);
and U12345 (N_12345,N_11491,N_10489);
and U12346 (N_12346,N_11979,N_10136);
nor U12347 (N_12347,N_11869,N_10233);
or U12348 (N_12348,N_11456,N_10428);
or U12349 (N_12349,N_11454,N_10900);
or U12350 (N_12350,N_10987,N_10002);
or U12351 (N_12351,N_10774,N_11997);
xor U12352 (N_12352,N_11070,N_11870);
xor U12353 (N_12353,N_11776,N_10849);
and U12354 (N_12354,N_10962,N_10109);
or U12355 (N_12355,N_11826,N_11882);
nor U12356 (N_12356,N_11503,N_11741);
nand U12357 (N_12357,N_10909,N_11857);
nor U12358 (N_12358,N_10137,N_11906);
xnor U12359 (N_12359,N_11775,N_10695);
or U12360 (N_12360,N_10331,N_10062);
and U12361 (N_12361,N_10702,N_11508);
and U12362 (N_12362,N_11858,N_10801);
or U12363 (N_12363,N_10912,N_11514);
and U12364 (N_12364,N_10876,N_10825);
nand U12365 (N_12365,N_11054,N_11795);
nand U12366 (N_12366,N_11677,N_11485);
nand U12367 (N_12367,N_11353,N_10739);
nand U12368 (N_12368,N_10902,N_10544);
nand U12369 (N_12369,N_11206,N_10413);
nor U12370 (N_12370,N_10791,N_11220);
nor U12371 (N_12371,N_10540,N_10118);
nand U12372 (N_12372,N_11377,N_11548);
or U12373 (N_12373,N_10092,N_10878);
nand U12374 (N_12374,N_11971,N_11570);
or U12375 (N_12375,N_11272,N_11889);
nand U12376 (N_12376,N_10401,N_11250);
and U12377 (N_12377,N_11771,N_10203);
nor U12378 (N_12378,N_10012,N_11819);
and U12379 (N_12379,N_10370,N_11817);
and U12380 (N_12380,N_10376,N_10710);
and U12381 (N_12381,N_11133,N_10648);
nand U12382 (N_12382,N_10820,N_10105);
nor U12383 (N_12383,N_11285,N_10532);
nor U12384 (N_12384,N_11319,N_10623);
or U12385 (N_12385,N_11803,N_10386);
and U12386 (N_12386,N_11844,N_10098);
or U12387 (N_12387,N_10330,N_11378);
nand U12388 (N_12388,N_10425,N_10247);
or U12389 (N_12389,N_11295,N_11287);
xnor U12390 (N_12390,N_10716,N_10888);
nand U12391 (N_12391,N_10069,N_11149);
or U12392 (N_12392,N_10372,N_10606);
nor U12393 (N_12393,N_11278,N_11974);
and U12394 (N_12394,N_11507,N_11550);
or U12395 (N_12395,N_10634,N_10637);
nor U12396 (N_12396,N_10639,N_11448);
or U12397 (N_12397,N_10578,N_11061);
or U12398 (N_12398,N_11881,N_11647);
or U12399 (N_12399,N_11575,N_10630);
nor U12400 (N_12400,N_10414,N_11407);
nor U12401 (N_12401,N_11116,N_10479);
nand U12402 (N_12402,N_11208,N_10396);
nor U12403 (N_12403,N_11745,N_11995);
nand U12404 (N_12404,N_11011,N_11276);
or U12405 (N_12405,N_10453,N_11861);
xnor U12406 (N_12406,N_11720,N_11665);
nand U12407 (N_12407,N_11552,N_10369);
and U12408 (N_12408,N_10788,N_11269);
and U12409 (N_12409,N_10350,N_11346);
xor U12410 (N_12410,N_10291,N_11721);
nand U12411 (N_12411,N_11829,N_11324);
nor U12412 (N_12412,N_10417,N_10613);
nor U12413 (N_12413,N_10202,N_11577);
xor U12414 (N_12414,N_11004,N_11904);
or U12415 (N_12415,N_11395,N_10484);
nand U12416 (N_12416,N_10094,N_10914);
xnor U12417 (N_12417,N_10293,N_10663);
or U12418 (N_12418,N_11525,N_11628);
nor U12419 (N_12419,N_11213,N_11713);
nand U12420 (N_12420,N_10921,N_10465);
nand U12421 (N_12421,N_11541,N_11651);
nor U12422 (N_12422,N_10516,N_10773);
nand U12423 (N_12423,N_11455,N_11702);
and U12424 (N_12424,N_11690,N_11447);
nor U12425 (N_12425,N_11559,N_11163);
or U12426 (N_12426,N_11486,N_11851);
nor U12427 (N_12427,N_10640,N_11544);
nor U12428 (N_12428,N_10241,N_10167);
nor U12429 (N_12429,N_10761,N_10067);
or U12430 (N_12430,N_11365,N_11232);
and U12431 (N_12431,N_11326,N_10446);
nor U12432 (N_12432,N_10195,N_11311);
or U12433 (N_12433,N_10612,N_10499);
or U12434 (N_12434,N_11588,N_10467);
nand U12435 (N_12435,N_10799,N_11173);
nand U12436 (N_12436,N_10173,N_11221);
nor U12437 (N_12437,N_11041,N_11060);
nand U12438 (N_12438,N_11804,N_10834);
nand U12439 (N_12439,N_11810,N_11427);
nand U12440 (N_12440,N_10994,N_10218);
and U12441 (N_12441,N_10186,N_10009);
nor U12442 (N_12442,N_10166,N_10550);
and U12443 (N_12443,N_10592,N_11814);
nand U12444 (N_12444,N_10452,N_11953);
xnor U12445 (N_12445,N_10862,N_11877);
xor U12446 (N_12446,N_10416,N_11875);
or U12447 (N_12447,N_10951,N_10322);
or U12448 (N_12448,N_10653,N_11769);
or U12449 (N_12449,N_11473,N_10937);
and U12450 (N_12450,N_10823,N_11343);
nor U12451 (N_12451,N_11692,N_10869);
and U12452 (N_12452,N_10768,N_10775);
or U12453 (N_12453,N_11373,N_11100);
nor U12454 (N_12454,N_10482,N_11415);
and U12455 (N_12455,N_10906,N_10996);
and U12456 (N_12456,N_11032,N_10800);
and U12457 (N_12457,N_11067,N_10691);
nand U12458 (N_12458,N_10077,N_11698);
or U12459 (N_12459,N_10442,N_11290);
xnor U12460 (N_12460,N_10692,N_11876);
nor U12461 (N_12461,N_10242,N_11899);
nor U12462 (N_12462,N_11336,N_10901);
and U12463 (N_12463,N_11172,N_11557);
nor U12464 (N_12464,N_10968,N_11451);
nor U12465 (N_12465,N_10531,N_11101);
and U12466 (N_12466,N_11537,N_10935);
and U12467 (N_12467,N_10485,N_11414);
or U12468 (N_12468,N_10473,N_10736);
nand U12469 (N_12469,N_10992,N_11667);
nor U12470 (N_12470,N_11728,N_11930);
nand U12471 (N_12471,N_10213,N_11376);
and U12472 (N_12472,N_10863,N_11996);
or U12473 (N_12473,N_10207,N_11735);
nand U12474 (N_12474,N_11216,N_11509);
or U12475 (N_12475,N_10043,N_11040);
nor U12476 (N_12476,N_10915,N_10183);
or U12477 (N_12477,N_11816,N_10728);
nand U12478 (N_12478,N_10162,N_11801);
or U12479 (N_12479,N_11564,N_10795);
and U12480 (N_12480,N_11452,N_11942);
xnor U12481 (N_12481,N_10406,N_10604);
nor U12482 (N_12482,N_10848,N_11385);
or U12483 (N_12483,N_11846,N_11691);
or U12484 (N_12484,N_10884,N_10495);
nor U12485 (N_12485,N_10806,N_10941);
or U12486 (N_12486,N_10100,N_11753);
and U12487 (N_12487,N_10125,N_10274);
and U12488 (N_12488,N_10766,N_10963);
nor U12489 (N_12489,N_10379,N_10304);
and U12490 (N_12490,N_11140,N_10525);
nand U12491 (N_12491,N_10185,N_11641);
or U12492 (N_12492,N_11973,N_10281);
nand U12493 (N_12493,N_11849,N_10078);
xor U12494 (N_12494,N_11843,N_10493);
nand U12495 (N_12495,N_11630,N_11240);
or U12496 (N_12496,N_10998,N_10846);
nor U12497 (N_12497,N_11197,N_10480);
or U12498 (N_12498,N_10412,N_10054);
and U12499 (N_12499,N_10128,N_11923);
nor U12500 (N_12500,N_11632,N_11331);
xor U12501 (N_12501,N_10158,N_10905);
nand U12502 (N_12502,N_10451,N_10919);
nor U12503 (N_12503,N_11093,N_10574);
or U12504 (N_12504,N_10932,N_11042);
nand U12505 (N_12505,N_11183,N_10335);
xor U12506 (N_12506,N_11510,N_10148);
and U12507 (N_12507,N_10966,N_10344);
xor U12508 (N_12508,N_11119,N_10680);
nand U12509 (N_12509,N_11574,N_10605);
and U12510 (N_12510,N_11445,N_11710);
and U12511 (N_12511,N_11568,N_11262);
nor U12512 (N_12512,N_10707,N_11905);
xnor U12513 (N_12513,N_10654,N_11223);
or U12514 (N_12514,N_10253,N_11640);
xnor U12515 (N_12515,N_10769,N_10004);
or U12516 (N_12516,N_10855,N_11088);
or U12517 (N_12517,N_10608,N_11777);
and U12518 (N_12518,N_10224,N_10594);
xor U12519 (N_12519,N_10156,N_11987);
nand U12520 (N_12520,N_11584,N_10440);
or U12521 (N_12521,N_11896,N_10958);
or U12522 (N_12522,N_10758,N_10095);
nor U12523 (N_12523,N_11255,N_11945);
or U12524 (N_12524,N_11793,N_10871);
nand U12525 (N_12525,N_10898,N_10449);
or U12526 (N_12526,N_10381,N_11045);
xor U12527 (N_12527,N_11430,N_11341);
and U12528 (N_12528,N_10145,N_11520);
nand U12529 (N_12529,N_11727,N_10075);
nand U12530 (N_12530,N_11178,N_11248);
and U12531 (N_12531,N_11058,N_10176);
nand U12532 (N_12532,N_10034,N_11910);
nand U12533 (N_12533,N_10432,N_10018);
nand U12534 (N_12534,N_11984,N_11354);
or U12535 (N_12535,N_10508,N_11533);
nor U12536 (N_12536,N_10065,N_11962);
and U12537 (N_12537,N_11535,N_10239);
nor U12538 (N_12538,N_10324,N_10553);
nand U12539 (N_12539,N_11523,N_10596);
or U12540 (N_12540,N_11624,N_11696);
nor U12541 (N_12541,N_10929,N_11409);
nand U12542 (N_12542,N_11391,N_11086);
and U12543 (N_12543,N_11121,N_10019);
nor U12544 (N_12544,N_11237,N_11404);
or U12545 (N_12545,N_10212,N_10753);
or U12546 (N_12546,N_10363,N_11351);
or U12547 (N_12547,N_11470,N_11231);
nor U12548 (N_12548,N_10073,N_11202);
and U12549 (N_12549,N_10832,N_10411);
or U12550 (N_12550,N_11805,N_11726);
xor U12551 (N_12551,N_10785,N_11788);
or U12552 (N_12552,N_11318,N_10219);
and U12553 (N_12553,N_11457,N_11521);
nand U12554 (N_12554,N_11951,N_10651);
and U12555 (N_12555,N_10563,N_11616);
and U12556 (N_12556,N_10658,N_11680);
or U12557 (N_12557,N_10868,N_10930);
xnor U12558 (N_12558,N_11392,N_10041);
or U12559 (N_12559,N_10283,N_10705);
nor U12560 (N_12560,N_11738,N_10813);
nand U12561 (N_12561,N_11370,N_11791);
nand U12562 (N_12562,N_11646,N_10437);
nor U12563 (N_12563,N_11725,N_11700);
xnor U12564 (N_12564,N_11259,N_10341);
and U12565 (N_12565,N_10822,N_10356);
xor U12566 (N_12566,N_11872,N_10039);
and U12567 (N_12567,N_10521,N_10424);
and U12568 (N_12568,N_11920,N_10471);
or U12569 (N_12569,N_10819,N_10240);
or U12570 (N_12570,N_11822,N_10161);
and U12571 (N_12571,N_10104,N_11403);
and U12572 (N_12572,N_11672,N_10895);
nand U12573 (N_12573,N_11794,N_11109);
nor U12574 (N_12574,N_11597,N_11864);
nand U12575 (N_12575,N_11025,N_10357);
nor U12576 (N_12576,N_10439,N_11420);
or U12577 (N_12577,N_11200,N_10216);
or U12578 (N_12578,N_11028,N_10779);
nor U12579 (N_12579,N_10821,N_11687);
nand U12580 (N_12580,N_11583,N_10087);
nor U12581 (N_12581,N_11383,N_11918);
and U12582 (N_12582,N_11715,N_10385);
xor U12583 (N_12583,N_11077,N_10575);
nand U12584 (N_12584,N_10534,N_11095);
nor U12585 (N_12585,N_11661,N_10014);
nand U12586 (N_12586,N_11883,N_10151);
nor U12587 (N_12587,N_10528,N_10954);
xor U12588 (N_12588,N_10960,N_10783);
and U12589 (N_12589,N_10587,N_10433);
and U12590 (N_12590,N_11402,N_11082);
or U12591 (N_12591,N_10581,N_10679);
nor U12592 (N_12592,N_10126,N_11111);
and U12593 (N_12593,N_11873,N_10714);
nand U12594 (N_12594,N_10111,N_10405);
nand U12595 (N_12595,N_11239,N_10891);
or U12596 (N_12596,N_11621,N_11079);
nor U12597 (N_12597,N_11315,N_11381);
nand U12598 (N_12598,N_11316,N_10887);
nor U12599 (N_12599,N_10666,N_10506);
or U12600 (N_12600,N_11024,N_10475);
xor U12601 (N_12601,N_10306,N_11339);
nor U12602 (N_12602,N_10049,N_11978);
nor U12603 (N_12603,N_10500,N_11982);
nor U12604 (N_12604,N_11688,N_10108);
nor U12605 (N_12605,N_10978,N_10762);
or U12606 (N_12606,N_10976,N_11610);
nor U12607 (N_12607,N_10660,N_10462);
and U12608 (N_12608,N_10090,N_11966);
nor U12609 (N_12609,N_11941,N_10607);
or U12610 (N_12610,N_10676,N_10590);
and U12611 (N_12611,N_11611,N_10262);
and U12612 (N_12612,N_10001,N_11113);
nand U12613 (N_12613,N_10616,N_11497);
or U12614 (N_12614,N_10358,N_11159);
or U12615 (N_12615,N_10458,N_11712);
xor U12616 (N_12616,N_10091,N_11950);
nor U12617 (N_12617,N_10042,N_11605);
nand U12618 (N_12618,N_11631,N_11675);
nand U12619 (N_12619,N_11484,N_10474);
nor U12620 (N_12620,N_11210,N_11754);
nand U12621 (N_12621,N_10328,N_11252);
nand U12622 (N_12622,N_10419,N_11289);
nor U12623 (N_12623,N_11600,N_11488);
nor U12624 (N_12624,N_10498,N_10551);
or U12625 (N_12625,N_11722,N_10177);
or U12626 (N_12626,N_10507,N_10292);
nand U12627 (N_12627,N_10257,N_11903);
or U12628 (N_12628,N_11468,N_10013);
nor U12629 (N_12629,N_10102,N_10650);
xor U12630 (N_12630,N_10483,N_11926);
nand U12631 (N_12631,N_11948,N_11059);
nand U12632 (N_12632,N_11481,N_11587);
and U12633 (N_12633,N_10872,N_11361);
nand U12634 (N_12634,N_11334,N_10420);
and U12635 (N_12635,N_10421,N_11911);
nand U12636 (N_12636,N_11531,N_11645);
nor U12637 (N_12637,N_11483,N_10509);
and U12638 (N_12638,N_10084,N_11879);
nor U12639 (N_12639,N_11313,N_11837);
nor U12640 (N_12640,N_11074,N_11052);
and U12641 (N_12641,N_11813,N_10742);
nand U12642 (N_12642,N_10853,N_11655);
or U12643 (N_12643,N_10367,N_10503);
nor U12644 (N_12644,N_11689,N_11620);
nand U12645 (N_12645,N_10547,N_11830);
xnor U12646 (N_12646,N_11214,N_10444);
nor U12647 (N_12647,N_10924,N_10975);
nand U12648 (N_12648,N_10957,N_10150);
nor U12649 (N_12649,N_10973,N_10722);
and U12650 (N_12650,N_11283,N_10160);
nor U12651 (N_12651,N_11136,N_10017);
or U12652 (N_12652,N_11740,N_10127);
nand U12653 (N_12653,N_11717,N_10389);
nand U12654 (N_12654,N_11224,N_11547);
and U12655 (N_12655,N_11207,N_11669);
or U12656 (N_12656,N_10624,N_11919);
or U12657 (N_12657,N_10246,N_10244);
nor U12658 (N_12658,N_10721,N_11258);
and U12659 (N_12659,N_10894,N_11626);
and U12660 (N_12660,N_10738,N_11253);
nand U12661 (N_12661,N_10021,N_10476);
nor U12662 (N_12662,N_10686,N_11401);
nand U12663 (N_12663,N_10189,N_10179);
and U12664 (N_12664,N_10235,N_11591);
nor U12665 (N_12665,N_11236,N_10539);
and U12666 (N_12666,N_11174,N_10838);
xnor U12667 (N_12667,N_11146,N_11245);
xor U12668 (N_12668,N_11848,N_10561);
and U12669 (N_12669,N_10448,N_10995);
or U12670 (N_12670,N_10422,N_10977);
and U12671 (N_12671,N_11792,N_10120);
nand U12672 (N_12672,N_11703,N_11685);
nand U12673 (N_12673,N_10229,N_10622);
and U12674 (N_12674,N_10980,N_11444);
nand U12675 (N_12675,N_10022,N_11490);
or U12676 (N_12676,N_10171,N_10466);
nor U12677 (N_12677,N_11358,N_10318);
or U12678 (N_12678,N_10536,N_11440);
and U12679 (N_12679,N_10866,N_11386);
nor U12680 (N_12680,N_10852,N_10734);
and U12681 (N_12681,N_11397,N_10032);
or U12682 (N_12682,N_11130,N_11286);
and U12683 (N_12683,N_10520,N_10910);
nor U12684 (N_12684,N_10044,N_10192);
xnor U12685 (N_12685,N_11037,N_10726);
or U12686 (N_12686,N_11737,N_11027);
xnor U12687 (N_12687,N_11446,N_10642);
nor U12688 (N_12688,N_10530,N_11530);
or U12689 (N_12689,N_10698,N_10015);
xor U12690 (N_12690,N_11008,N_10056);
xor U12691 (N_12691,N_11015,N_10059);
nor U12692 (N_12692,N_11348,N_10811);
xnor U12693 (N_12693,N_10390,N_11274);
nand U12694 (N_12694,N_11029,N_11671);
nor U12695 (N_12695,N_11180,N_10546);
xnor U12696 (N_12696,N_10011,N_10088);
xnor U12697 (N_12697,N_10890,N_10765);
or U12698 (N_12698,N_10903,N_11763);
or U12699 (N_12699,N_11238,N_10205);
nand U12700 (N_12700,N_11091,N_11893);
or U12701 (N_12701,N_11472,N_10083);
nor U12702 (N_12702,N_10802,N_10159);
or U12703 (N_12703,N_10999,N_10922);
or U12704 (N_12704,N_11280,N_11284);
nand U12705 (N_12705,N_11886,N_10251);
nor U12706 (N_12706,N_10595,N_11006);
nor U12707 (N_12707,N_10089,N_11786);
or U12708 (N_12708,N_10610,N_10504);
xnor U12709 (N_12709,N_10833,N_11949);
or U12710 (N_12710,N_10817,N_11744);
nand U12711 (N_12711,N_11388,N_10669);
and U12712 (N_12712,N_10248,N_10602);
or U12713 (N_12713,N_10234,N_11828);
and U12714 (N_12714,N_10670,N_11308);
or U12715 (N_12715,N_10464,N_11937);
nor U12716 (N_12716,N_10050,N_10110);
nor U12717 (N_12717,N_10803,N_11551);
xor U12718 (N_12718,N_10615,N_11917);
nor U12719 (N_12719,N_10261,N_10699);
nand U12720 (N_12720,N_10798,N_10263);
nand U12721 (N_12721,N_11783,N_11598);
nor U12722 (N_12722,N_11099,N_10805);
or U12723 (N_12723,N_11652,N_10829);
and U12724 (N_12724,N_10636,N_10646);
xor U12725 (N_12725,N_11144,N_10625);
xor U12726 (N_12726,N_11241,N_11784);
nor U12727 (N_12727,N_11731,N_10885);
xnor U12728 (N_12728,N_11787,N_10492);
nand U12729 (N_12729,N_10031,N_10845);
and U12730 (N_12730,N_10600,N_11303);
and U12731 (N_12731,N_11261,N_10988);
or U12732 (N_12732,N_11555,N_11083);
nor U12733 (N_12733,N_10426,N_10584);
or U12734 (N_12734,N_10598,N_10579);
nor U12735 (N_12735,N_11755,N_11063);
or U12736 (N_12736,N_11332,N_10647);
nand U12737 (N_12737,N_11743,N_10926);
nand U12738 (N_12738,N_11585,N_11967);
nand U12739 (N_12739,N_10577,N_10301);
nor U12740 (N_12740,N_10005,N_11120);
and U12741 (N_12741,N_11563,N_10840);
or U12742 (N_12742,N_11832,N_11196);
or U12743 (N_12743,N_11825,N_11335);
or U12744 (N_12744,N_10777,N_11960);
or U12745 (N_12745,N_11656,N_11148);
or U12746 (N_12746,N_11184,N_11384);
nand U12747 (N_12747,N_11466,N_10138);
and U12748 (N_12748,N_10223,N_11304);
nor U12749 (N_12749,N_10326,N_11781);
nor U12750 (N_12750,N_10934,N_10007);
nor U12751 (N_12751,N_11129,N_11234);
and U12752 (N_12752,N_10163,N_11853);
or U12753 (N_12753,N_10258,N_10142);
or U12754 (N_12754,N_10454,N_11502);
and U12755 (N_12755,N_10754,N_10645);
nor U12756 (N_12756,N_11474,N_10333);
nor U12757 (N_12757,N_11194,N_11215);
nand U12758 (N_12758,N_10351,N_10983);
xnor U12759 (N_12759,N_11693,N_11999);
nor U12760 (N_12760,N_10787,N_10303);
or U12761 (N_12761,N_11081,N_10430);
nand U12762 (N_12762,N_11493,N_11306);
nor U12763 (N_12763,N_11105,N_11766);
and U12764 (N_12764,N_10074,N_10366);
and U12765 (N_12765,N_11833,N_10956);
and U12766 (N_12766,N_10184,N_10867);
or U12767 (N_12767,N_10441,N_10377);
or U12768 (N_12768,N_10327,N_11084);
and U12769 (N_12769,N_11127,N_11257);
nand U12770 (N_12770,N_11036,N_10794);
and U12771 (N_12771,N_11453,N_10282);
xor U12772 (N_12772,N_11426,N_11762);
and U12773 (N_12773,N_10132,N_10700);
or U12774 (N_12774,N_10689,N_10626);
and U12775 (N_12775,N_10631,N_11701);
or U12776 (N_12776,N_11495,N_10152);
and U12777 (N_12777,N_11301,N_10380);
or U12778 (N_12778,N_10016,N_11808);
xor U12779 (N_12779,N_11895,N_11458);
nor U12780 (N_12780,N_11205,N_11902);
nand U12781 (N_12781,N_11711,N_10548);
and U12782 (N_12782,N_11394,N_10748);
and U12783 (N_12783,N_11952,N_11292);
xor U12784 (N_12784,N_10214,N_11141);
nor U12785 (N_12785,N_10955,N_10741);
or U12786 (N_12786,N_10149,N_10896);
and U12787 (N_12787,N_10302,N_10300);
and U12788 (N_12788,N_10368,N_10830);
xnor U12789 (N_12789,N_10562,N_11198);
and U12790 (N_12790,N_11489,N_11137);
xor U12791 (N_12791,N_10949,N_11980);
and U12792 (N_12792,N_10153,N_10567);
xnor U12793 (N_12793,N_11596,N_11765);
nand U12794 (N_12794,N_10569,N_10814);
and U12795 (N_12795,N_10315,N_11653);
and U12796 (N_12796,N_11812,N_10134);
xnor U12797 (N_12797,N_10382,N_11838);
or U12798 (N_12798,N_11418,N_11909);
nand U12799 (N_12799,N_10674,N_10810);
nor U12800 (N_12800,N_11800,N_10675);
or U12801 (N_12801,N_10776,N_11288);
nand U12802 (N_12802,N_11190,N_11674);
nand U12803 (N_12803,N_10911,N_11425);
or U12804 (N_12804,N_11366,N_10066);
nor U12805 (N_12805,N_11602,N_11422);
and U12806 (N_12806,N_11922,N_11161);
nand U12807 (N_12807,N_10339,N_11940);
nor U12808 (N_12808,N_10842,N_10693);
and U12809 (N_12809,N_10759,N_10673);
nand U12810 (N_12810,N_10398,N_10771);
and U12811 (N_12811,N_10456,N_11554);
or U12812 (N_12812,N_10681,N_11374);
nor U12813 (N_12813,N_10943,N_11225);
nor U12814 (N_12814,N_11827,N_10632);
and U12815 (N_12815,N_10835,N_11915);
or U12816 (N_12816,N_10312,N_11492);
xnor U12817 (N_12817,N_10755,N_10953);
nor U12818 (N_12818,N_10572,N_11251);
or U12819 (N_12819,N_10950,N_11871);
nor U12820 (N_12820,N_10427,N_11850);
and U12821 (N_12821,N_11914,N_11122);
and U12822 (N_12822,N_10655,N_10082);
or U12823 (N_12823,N_10337,N_10395);
nor U12824 (N_12824,N_10844,N_11622);
and U12825 (N_12825,N_10298,N_10948);
nor U12826 (N_12826,N_11242,N_10583);
xor U12827 (N_12827,N_10588,N_10621);
or U12828 (N_12828,N_11080,N_11017);
nor U12829 (N_12829,N_10290,N_10209);
or U12830 (N_12830,N_10635,N_10146);
and U12831 (N_12831,N_11874,N_10860);
nand U12832 (N_12832,N_11193,N_10511);
or U12833 (N_12833,N_10619,N_10169);
nor U12834 (N_12834,N_11013,N_11019);
nor U12835 (N_12835,N_11108,N_10338);
nand U12836 (N_12836,N_10459,N_10347);
and U12837 (N_12837,N_10538,N_10175);
xnor U12838 (N_12838,N_11779,N_11683);
nand U12839 (N_12839,N_11460,N_11176);
xnor U12840 (N_12840,N_11772,N_11912);
nor U12841 (N_12841,N_11005,N_10571);
and U12842 (N_12842,N_10254,N_11390);
or U12843 (N_12843,N_11073,N_11222);
and U12844 (N_12844,N_10048,N_11659);
and U12845 (N_12845,N_11534,N_11662);
nor U12846 (N_12846,N_11513,N_10305);
nor U12847 (N_12847,N_11123,N_11044);
nor U12848 (N_12848,N_11170,N_11642);
and U12849 (N_12849,N_10273,N_10920);
nor U12850 (N_12850,N_11156,N_11310);
and U12851 (N_12851,N_11209,N_10549);
nand U12852 (N_12852,N_11393,N_10269);
or U12853 (N_12853,N_11885,N_10278);
nor U12854 (N_12854,N_10217,N_11344);
and U12855 (N_12855,N_11660,N_10629);
nand U12856 (N_12856,N_10053,N_11296);
or U12857 (N_12857,N_11957,N_11796);
or U12858 (N_12858,N_10725,N_10314);
xnor U12859 (N_12859,N_10724,N_10770);
nor U12860 (N_12860,N_10313,N_10731);
nor U12861 (N_12861,N_11560,N_10114);
nor U12862 (N_12862,N_11581,N_11954);
or U12863 (N_12863,N_10656,N_11462);
nand U12864 (N_12864,N_10633,N_10455);
and U12865 (N_12865,N_10140,N_11201);
nand U12866 (N_12866,N_10361,N_10470);
or U12867 (N_12867,N_11798,N_11050);
nand U12868 (N_12868,N_11697,N_10010);
nor U12869 (N_12869,N_10542,N_10388);
xnor U12870 (N_12870,N_11465,N_11573);
nor U12871 (N_12871,N_11650,N_11847);
nor U12872 (N_12872,N_11993,N_11664);
and U12873 (N_12873,N_10589,N_11135);
nand U12874 (N_12874,N_10713,N_10518);
nor U12875 (N_12875,N_11612,N_10652);
and U12876 (N_12876,N_10096,N_10687);
and U12877 (N_12877,N_11408,N_11266);
or U12878 (N_12878,N_10343,N_10576);
nor U12879 (N_12879,N_10268,N_10883);
xnor U12880 (N_12880,N_11188,N_10618);
nor U12881 (N_12881,N_10135,N_10165);
nand U12882 (N_12882,N_11092,N_10037);
xnor U12883 (N_12883,N_11707,N_10965);
nor U12884 (N_12884,N_10824,N_11423);
and U12885 (N_12885,N_11065,N_10704);
nor U12886 (N_12886,N_11695,N_10865);
nor U12887 (N_12887,N_10387,N_10818);
nor U12888 (N_12888,N_10609,N_11888);
nor U12889 (N_12889,N_10505,N_10182);
nor U12890 (N_12890,N_10545,N_10552);
or U12891 (N_12891,N_10122,N_11138);
and U12892 (N_12892,N_11459,N_10266);
or U12893 (N_12893,N_10751,N_11724);
and U12894 (N_12894,N_10277,N_10881);
nand U12895 (N_12895,N_11212,N_11649);
nor U12896 (N_12896,N_11964,N_11281);
or U12897 (N_12897,N_11986,N_10038);
or U12898 (N_12898,N_10252,N_10938);
nand U12899 (N_12899,N_11411,N_11264);
nand U12900 (N_12900,N_10997,N_11449);
nand U12901 (N_12901,N_11421,N_10434);
nand U12902 (N_12902,N_10106,N_10877);
or U12903 (N_12903,N_10851,N_11932);
nor U12904 (N_12904,N_10792,N_11935);
nor U12905 (N_12905,N_10311,N_11961);
and U12906 (N_12906,N_11561,N_10101);
nand U12907 (N_12907,N_10024,N_11345);
and U12908 (N_12908,N_11532,N_10939);
xnor U12909 (N_12909,N_10232,N_11382);
nand U12910 (N_12910,N_10706,N_11412);
and U12911 (N_12911,N_10843,N_10204);
nor U12912 (N_12912,N_11760,N_10265);
or U12913 (N_12913,N_11933,N_10780);
nor U12914 (N_12914,N_10423,N_11009);
nor U12915 (N_12915,N_10990,N_11218);
nor U12916 (N_12916,N_10113,N_10119);
and U12917 (N_12917,N_11939,N_10857);
nor U12918 (N_12918,N_11347,N_10893);
nand U12919 (N_12919,N_11469,N_11463);
nor U12920 (N_12920,N_11676,N_11579);
or U12921 (N_12921,N_10230,N_11884);
nand U12922 (N_12922,N_10397,N_11439);
nand U12923 (N_12923,N_10701,N_10740);
and U12924 (N_12924,N_10560,N_11228);
nor U12925 (N_12925,N_10400,N_11658);
xor U12926 (N_12926,N_11782,N_10959);
nand U12927 (N_12927,N_10812,N_11856);
nand U12928 (N_12928,N_11114,N_11944);
nor U12929 (N_12929,N_11467,N_11586);
nor U12930 (N_12930,N_11071,N_10850);
and U12931 (N_12931,N_11368,N_11679);
and U12932 (N_12932,N_10392,N_11556);
and U12933 (N_12933,N_11461,N_11699);
or U12934 (N_12934,N_10431,N_10672);
nor U12935 (N_12935,N_10870,N_11809);
nor U12936 (N_12936,N_10196,N_11968);
nor U12937 (N_12937,N_11629,N_11157);
and U12938 (N_12938,N_10181,N_11406);
nor U12939 (N_12939,N_10228,N_10517);
and U12940 (N_12940,N_11751,N_10289);
and U12941 (N_12941,N_11890,N_11868);
nor U12942 (N_12942,N_11191,N_11580);
nand U12943 (N_12943,N_11553,N_10349);
nand U12944 (N_12944,N_11797,N_11399);
nor U12945 (N_12945,N_10481,N_10879);
and U12946 (N_12946,N_11350,N_11410);
or U12947 (N_12947,N_10685,N_10355);
nor U12948 (N_12948,N_11654,N_11150);
nor U12949 (N_12949,N_11282,N_11355);
or U12950 (N_12950,N_11496,N_10501);
nor U12951 (N_12951,N_11010,N_10317);
xor U12952 (N_12952,N_11742,N_11593);
nor U12953 (N_12953,N_11604,N_11139);
nor U12954 (N_12954,N_10683,N_11300);
nand U12955 (N_12955,N_11112,N_10597);
or U12956 (N_12956,N_11294,N_10131);
or U12957 (N_12957,N_10931,N_11181);
nand U12958 (N_12958,N_10668,N_11545);
nor U12959 (N_12959,N_11730,N_11072);
nand U12960 (N_12960,N_11519,N_10945);
nand U12961 (N_12961,N_11325,N_10408);
nor U12962 (N_12962,N_11860,N_10450);
nand U12963 (N_12963,N_11387,N_10767);
xor U12964 (N_12964,N_10662,N_10133);
nor U12965 (N_12965,N_11021,N_11413);
xor U12966 (N_12966,N_10908,N_11002);
xnor U12967 (N_12967,N_11608,N_11160);
or U12968 (N_12968,N_10677,N_10601);
xor U12969 (N_12969,N_10445,N_10786);
nor U12970 (N_12970,N_11106,N_11263);
nand U12971 (N_12971,N_10573,N_11627);
nand U12972 (N_12972,N_10154,N_10051);
nor U12973 (N_12973,N_11958,N_11778);
and U12974 (N_12974,N_11512,N_11729);
and U12975 (N_12975,N_11716,N_11836);
nor U12976 (N_12976,N_11000,N_11254);
or U12977 (N_12977,N_10764,N_11068);
or U12978 (N_12978,N_10979,N_10756);
nor U12979 (N_12979,N_11733,N_11442);
and U12980 (N_12980,N_11634,N_11064);
and U12981 (N_12981,N_11673,N_10816);
and U12982 (N_12982,N_10745,N_10116);
nor U12983 (N_12983,N_11169,N_10760);
nand U12984 (N_12984,N_11268,N_11842);
and U12985 (N_12985,N_11988,N_11956);
and U12986 (N_12986,N_10936,N_11096);
or U12987 (N_12987,N_11089,N_10732);
or U12988 (N_12988,N_10665,N_11026);
and U12989 (N_12989,N_10040,N_10882);
xnor U12990 (N_12990,N_10661,N_11433);
nand U12991 (N_12991,N_10063,N_10599);
xor U12992 (N_12992,N_11862,N_10827);
or U12993 (N_12993,N_10346,N_10892);
and U12994 (N_12994,N_10899,N_10418);
nand U12995 (N_12995,N_10046,N_10345);
and U12996 (N_12996,N_11023,N_10172);
and U12997 (N_12997,N_11204,N_10115);
and U12998 (N_12998,N_10027,N_11983);
nor U12999 (N_12999,N_11562,N_11166);
and U13000 (N_13000,N_11907,N_10645);
nor U13001 (N_13001,N_10752,N_11925);
nor U13002 (N_13002,N_11539,N_10784);
nand U13003 (N_13003,N_11451,N_10108);
and U13004 (N_13004,N_10764,N_11653);
nor U13005 (N_13005,N_10721,N_10952);
nand U13006 (N_13006,N_10294,N_11851);
nand U13007 (N_13007,N_10924,N_10876);
nand U13008 (N_13008,N_11861,N_10805);
nor U13009 (N_13009,N_11959,N_10029);
or U13010 (N_13010,N_10346,N_11854);
nand U13011 (N_13011,N_11623,N_11740);
xor U13012 (N_13012,N_11765,N_10471);
or U13013 (N_13013,N_11667,N_10058);
xnor U13014 (N_13014,N_11614,N_11296);
nor U13015 (N_13015,N_10895,N_11829);
nor U13016 (N_13016,N_10935,N_11717);
and U13017 (N_13017,N_11578,N_11208);
or U13018 (N_13018,N_10422,N_11105);
nand U13019 (N_13019,N_10097,N_10902);
nor U13020 (N_13020,N_10669,N_11392);
and U13021 (N_13021,N_10416,N_10196);
and U13022 (N_13022,N_11981,N_10713);
and U13023 (N_13023,N_10543,N_11310);
nand U13024 (N_13024,N_11767,N_10967);
xor U13025 (N_13025,N_11053,N_10527);
nor U13026 (N_13026,N_10409,N_11225);
nand U13027 (N_13027,N_11201,N_10884);
nand U13028 (N_13028,N_11449,N_10457);
xnor U13029 (N_13029,N_10168,N_11788);
nor U13030 (N_13030,N_11888,N_11812);
xnor U13031 (N_13031,N_11111,N_10384);
nor U13032 (N_13032,N_10302,N_11572);
and U13033 (N_13033,N_11418,N_10818);
nor U13034 (N_13034,N_11961,N_10045);
nor U13035 (N_13035,N_10152,N_10662);
nor U13036 (N_13036,N_10934,N_10843);
nand U13037 (N_13037,N_11900,N_11352);
nand U13038 (N_13038,N_10067,N_10391);
nand U13039 (N_13039,N_11306,N_11323);
and U13040 (N_13040,N_11044,N_11968);
and U13041 (N_13041,N_10248,N_11280);
xor U13042 (N_13042,N_10902,N_10958);
xnor U13043 (N_13043,N_11909,N_11031);
nand U13044 (N_13044,N_11988,N_11889);
or U13045 (N_13045,N_11477,N_11206);
nand U13046 (N_13046,N_10181,N_11670);
and U13047 (N_13047,N_11713,N_11052);
or U13048 (N_13048,N_11976,N_11686);
or U13049 (N_13049,N_10718,N_10290);
nand U13050 (N_13050,N_10138,N_10554);
nand U13051 (N_13051,N_11018,N_11917);
and U13052 (N_13052,N_11651,N_11659);
nor U13053 (N_13053,N_10345,N_10929);
nor U13054 (N_13054,N_11154,N_11046);
and U13055 (N_13055,N_11366,N_10171);
or U13056 (N_13056,N_11113,N_11737);
nand U13057 (N_13057,N_11340,N_10627);
nor U13058 (N_13058,N_10204,N_10087);
nor U13059 (N_13059,N_11831,N_11452);
nor U13060 (N_13060,N_10018,N_10784);
xor U13061 (N_13061,N_11213,N_10973);
and U13062 (N_13062,N_11220,N_10966);
and U13063 (N_13063,N_11393,N_11089);
nor U13064 (N_13064,N_10529,N_10555);
and U13065 (N_13065,N_11671,N_10842);
nor U13066 (N_13066,N_10345,N_10700);
nor U13067 (N_13067,N_10105,N_10137);
nand U13068 (N_13068,N_10532,N_11306);
and U13069 (N_13069,N_11209,N_10468);
and U13070 (N_13070,N_11952,N_11902);
xor U13071 (N_13071,N_10730,N_10280);
nand U13072 (N_13072,N_11687,N_11332);
and U13073 (N_13073,N_10972,N_11756);
or U13074 (N_13074,N_10462,N_10716);
nor U13075 (N_13075,N_10319,N_11614);
nand U13076 (N_13076,N_10931,N_10723);
nor U13077 (N_13077,N_11461,N_10403);
and U13078 (N_13078,N_11152,N_11853);
or U13079 (N_13079,N_11981,N_11591);
nor U13080 (N_13080,N_11679,N_11414);
xnor U13081 (N_13081,N_10183,N_11707);
nand U13082 (N_13082,N_10786,N_11657);
nor U13083 (N_13083,N_10626,N_11705);
or U13084 (N_13084,N_10956,N_10718);
nor U13085 (N_13085,N_10620,N_10991);
xor U13086 (N_13086,N_10061,N_10831);
or U13087 (N_13087,N_11620,N_10007);
and U13088 (N_13088,N_11215,N_10679);
and U13089 (N_13089,N_11408,N_10778);
xor U13090 (N_13090,N_11231,N_11045);
or U13091 (N_13091,N_11741,N_11259);
nand U13092 (N_13092,N_11550,N_11702);
nor U13093 (N_13093,N_11654,N_11014);
nor U13094 (N_13094,N_10956,N_10073);
xor U13095 (N_13095,N_10863,N_11620);
or U13096 (N_13096,N_11899,N_10001);
xnor U13097 (N_13097,N_11197,N_10519);
nand U13098 (N_13098,N_10584,N_10759);
nor U13099 (N_13099,N_10868,N_11888);
xnor U13100 (N_13100,N_11153,N_10152);
nand U13101 (N_13101,N_10083,N_11842);
or U13102 (N_13102,N_11479,N_10269);
and U13103 (N_13103,N_11004,N_10295);
nand U13104 (N_13104,N_10416,N_11496);
nor U13105 (N_13105,N_10229,N_11066);
or U13106 (N_13106,N_11930,N_10148);
or U13107 (N_13107,N_10755,N_10186);
xor U13108 (N_13108,N_11658,N_11198);
xnor U13109 (N_13109,N_10110,N_10017);
and U13110 (N_13110,N_10406,N_11114);
and U13111 (N_13111,N_11470,N_10017);
or U13112 (N_13112,N_11161,N_11913);
or U13113 (N_13113,N_11012,N_11402);
nand U13114 (N_13114,N_11876,N_11604);
nand U13115 (N_13115,N_10366,N_10060);
and U13116 (N_13116,N_11268,N_11088);
and U13117 (N_13117,N_11919,N_10963);
xnor U13118 (N_13118,N_11552,N_10192);
or U13119 (N_13119,N_10743,N_10649);
nor U13120 (N_13120,N_11424,N_10475);
and U13121 (N_13121,N_10558,N_11980);
or U13122 (N_13122,N_11828,N_11307);
xnor U13123 (N_13123,N_10029,N_11167);
nand U13124 (N_13124,N_11900,N_11190);
and U13125 (N_13125,N_10527,N_11974);
and U13126 (N_13126,N_10941,N_10093);
or U13127 (N_13127,N_11129,N_10196);
xor U13128 (N_13128,N_10760,N_11622);
nor U13129 (N_13129,N_10410,N_10990);
and U13130 (N_13130,N_11760,N_10019);
or U13131 (N_13131,N_10657,N_10496);
or U13132 (N_13132,N_10755,N_11127);
and U13133 (N_13133,N_11520,N_11363);
or U13134 (N_13134,N_10656,N_11981);
nand U13135 (N_13135,N_11441,N_10912);
and U13136 (N_13136,N_10329,N_11952);
and U13137 (N_13137,N_10328,N_11476);
and U13138 (N_13138,N_10665,N_11574);
nand U13139 (N_13139,N_11679,N_10435);
and U13140 (N_13140,N_11571,N_10073);
nand U13141 (N_13141,N_10939,N_11344);
xnor U13142 (N_13142,N_10066,N_10079);
nand U13143 (N_13143,N_10985,N_11455);
or U13144 (N_13144,N_10058,N_11340);
xor U13145 (N_13145,N_10592,N_10070);
and U13146 (N_13146,N_11216,N_10293);
nand U13147 (N_13147,N_11329,N_10427);
or U13148 (N_13148,N_10391,N_10338);
nor U13149 (N_13149,N_10447,N_10144);
nor U13150 (N_13150,N_10326,N_11929);
and U13151 (N_13151,N_10355,N_11554);
xor U13152 (N_13152,N_10598,N_11894);
nand U13153 (N_13153,N_10567,N_10634);
xnor U13154 (N_13154,N_10553,N_10945);
nand U13155 (N_13155,N_11690,N_11674);
and U13156 (N_13156,N_11016,N_11210);
or U13157 (N_13157,N_10968,N_11793);
or U13158 (N_13158,N_11145,N_10121);
nand U13159 (N_13159,N_10662,N_11894);
nor U13160 (N_13160,N_11353,N_11484);
or U13161 (N_13161,N_10855,N_11927);
nor U13162 (N_13162,N_11221,N_11584);
or U13163 (N_13163,N_10237,N_11094);
or U13164 (N_13164,N_10078,N_10983);
and U13165 (N_13165,N_11484,N_10606);
xor U13166 (N_13166,N_10079,N_10368);
nor U13167 (N_13167,N_10822,N_10373);
nand U13168 (N_13168,N_10751,N_10590);
or U13169 (N_13169,N_11672,N_10612);
and U13170 (N_13170,N_11091,N_11073);
or U13171 (N_13171,N_10385,N_10536);
and U13172 (N_13172,N_10876,N_11578);
nor U13173 (N_13173,N_10617,N_11003);
nand U13174 (N_13174,N_10982,N_10334);
or U13175 (N_13175,N_11206,N_11664);
or U13176 (N_13176,N_10071,N_10103);
nor U13177 (N_13177,N_11654,N_10370);
or U13178 (N_13178,N_10027,N_11922);
nor U13179 (N_13179,N_10806,N_10226);
or U13180 (N_13180,N_11435,N_11754);
or U13181 (N_13181,N_10999,N_11901);
or U13182 (N_13182,N_11578,N_11543);
xor U13183 (N_13183,N_10531,N_11207);
nor U13184 (N_13184,N_10448,N_11686);
xor U13185 (N_13185,N_10534,N_10045);
or U13186 (N_13186,N_10505,N_11658);
xnor U13187 (N_13187,N_11651,N_10622);
nor U13188 (N_13188,N_11548,N_10943);
nor U13189 (N_13189,N_11687,N_11775);
nand U13190 (N_13190,N_10530,N_11595);
nand U13191 (N_13191,N_11010,N_11464);
xnor U13192 (N_13192,N_11451,N_10022);
and U13193 (N_13193,N_10295,N_11720);
nand U13194 (N_13194,N_11922,N_11442);
nor U13195 (N_13195,N_10315,N_10518);
nand U13196 (N_13196,N_11475,N_10500);
or U13197 (N_13197,N_10324,N_10980);
xor U13198 (N_13198,N_11339,N_10033);
and U13199 (N_13199,N_10726,N_10208);
and U13200 (N_13200,N_11467,N_10485);
or U13201 (N_13201,N_11017,N_11623);
nand U13202 (N_13202,N_10613,N_10133);
or U13203 (N_13203,N_11017,N_10373);
or U13204 (N_13204,N_11068,N_11713);
or U13205 (N_13205,N_11752,N_11835);
or U13206 (N_13206,N_10896,N_11129);
and U13207 (N_13207,N_11261,N_11441);
and U13208 (N_13208,N_11098,N_11395);
nand U13209 (N_13209,N_11589,N_10535);
or U13210 (N_13210,N_10684,N_11288);
xnor U13211 (N_13211,N_11016,N_11936);
nor U13212 (N_13212,N_10800,N_10531);
nor U13213 (N_13213,N_11341,N_11545);
or U13214 (N_13214,N_11741,N_10897);
xor U13215 (N_13215,N_10844,N_11954);
nor U13216 (N_13216,N_10795,N_10223);
nor U13217 (N_13217,N_10279,N_10791);
or U13218 (N_13218,N_11760,N_10995);
xor U13219 (N_13219,N_10043,N_10880);
nand U13220 (N_13220,N_10911,N_10040);
nor U13221 (N_13221,N_11152,N_11872);
nand U13222 (N_13222,N_10100,N_11884);
and U13223 (N_13223,N_10239,N_10761);
nor U13224 (N_13224,N_10091,N_10468);
or U13225 (N_13225,N_11003,N_11991);
and U13226 (N_13226,N_10599,N_10879);
nor U13227 (N_13227,N_11046,N_11890);
nor U13228 (N_13228,N_11327,N_11712);
nand U13229 (N_13229,N_11150,N_10868);
nand U13230 (N_13230,N_11436,N_10911);
nor U13231 (N_13231,N_11808,N_10680);
nand U13232 (N_13232,N_10161,N_10134);
or U13233 (N_13233,N_11639,N_11742);
nor U13234 (N_13234,N_11675,N_10572);
xnor U13235 (N_13235,N_11150,N_10920);
nand U13236 (N_13236,N_10566,N_11096);
and U13237 (N_13237,N_10529,N_11788);
and U13238 (N_13238,N_10186,N_11634);
nand U13239 (N_13239,N_11156,N_10003);
nor U13240 (N_13240,N_11392,N_11482);
or U13241 (N_13241,N_10922,N_11352);
or U13242 (N_13242,N_10505,N_11943);
nand U13243 (N_13243,N_10088,N_11774);
or U13244 (N_13244,N_10575,N_10433);
xnor U13245 (N_13245,N_10772,N_11121);
nand U13246 (N_13246,N_11928,N_10140);
xor U13247 (N_13247,N_10090,N_10066);
nor U13248 (N_13248,N_10779,N_10458);
nor U13249 (N_13249,N_10299,N_10383);
nand U13250 (N_13250,N_11464,N_11297);
nor U13251 (N_13251,N_10795,N_11412);
nand U13252 (N_13252,N_11305,N_10302);
nor U13253 (N_13253,N_11138,N_10916);
nand U13254 (N_13254,N_11122,N_11678);
or U13255 (N_13255,N_11971,N_11108);
or U13256 (N_13256,N_10698,N_11660);
or U13257 (N_13257,N_10043,N_11808);
nor U13258 (N_13258,N_10926,N_10171);
nor U13259 (N_13259,N_11842,N_11029);
and U13260 (N_13260,N_10636,N_11940);
and U13261 (N_13261,N_11696,N_10541);
and U13262 (N_13262,N_11235,N_11269);
xor U13263 (N_13263,N_11767,N_11107);
or U13264 (N_13264,N_10792,N_10751);
nor U13265 (N_13265,N_10355,N_11045);
nor U13266 (N_13266,N_11745,N_11680);
and U13267 (N_13267,N_10502,N_10979);
and U13268 (N_13268,N_11522,N_10200);
and U13269 (N_13269,N_10322,N_10800);
nor U13270 (N_13270,N_10958,N_11583);
or U13271 (N_13271,N_11317,N_11149);
xor U13272 (N_13272,N_11672,N_10616);
nand U13273 (N_13273,N_11337,N_10766);
nand U13274 (N_13274,N_10662,N_10869);
and U13275 (N_13275,N_10625,N_11607);
or U13276 (N_13276,N_11092,N_10190);
nor U13277 (N_13277,N_10364,N_10227);
nand U13278 (N_13278,N_10662,N_10437);
nand U13279 (N_13279,N_11190,N_11693);
nand U13280 (N_13280,N_10281,N_11927);
or U13281 (N_13281,N_11980,N_10871);
nor U13282 (N_13282,N_11076,N_11533);
nand U13283 (N_13283,N_11591,N_11834);
nand U13284 (N_13284,N_11480,N_11034);
and U13285 (N_13285,N_10694,N_11941);
and U13286 (N_13286,N_10882,N_10867);
nor U13287 (N_13287,N_10224,N_10421);
nand U13288 (N_13288,N_11561,N_10253);
or U13289 (N_13289,N_11924,N_11060);
nand U13290 (N_13290,N_11408,N_10006);
nor U13291 (N_13291,N_10627,N_10108);
xor U13292 (N_13292,N_11135,N_11449);
nand U13293 (N_13293,N_11974,N_11898);
nor U13294 (N_13294,N_10636,N_10274);
nor U13295 (N_13295,N_11527,N_10328);
or U13296 (N_13296,N_10646,N_10599);
or U13297 (N_13297,N_10124,N_10729);
nand U13298 (N_13298,N_11075,N_11416);
nor U13299 (N_13299,N_10459,N_11479);
nand U13300 (N_13300,N_11202,N_11873);
and U13301 (N_13301,N_10701,N_10341);
and U13302 (N_13302,N_11313,N_10013);
or U13303 (N_13303,N_11176,N_10744);
nor U13304 (N_13304,N_11734,N_10560);
and U13305 (N_13305,N_10855,N_10470);
nand U13306 (N_13306,N_10321,N_10912);
or U13307 (N_13307,N_11535,N_10300);
or U13308 (N_13308,N_10423,N_11583);
nor U13309 (N_13309,N_10045,N_11113);
nand U13310 (N_13310,N_11925,N_11768);
or U13311 (N_13311,N_11062,N_10441);
and U13312 (N_13312,N_10471,N_11926);
xnor U13313 (N_13313,N_11842,N_11545);
or U13314 (N_13314,N_11636,N_10403);
nor U13315 (N_13315,N_11708,N_11215);
or U13316 (N_13316,N_10774,N_10134);
nand U13317 (N_13317,N_10099,N_11990);
and U13318 (N_13318,N_11650,N_10613);
or U13319 (N_13319,N_11652,N_11700);
and U13320 (N_13320,N_10113,N_11148);
nor U13321 (N_13321,N_11512,N_11728);
xor U13322 (N_13322,N_11891,N_10006);
or U13323 (N_13323,N_10778,N_11562);
nand U13324 (N_13324,N_10377,N_11018);
or U13325 (N_13325,N_11948,N_11242);
nand U13326 (N_13326,N_11131,N_10119);
xor U13327 (N_13327,N_11498,N_11305);
and U13328 (N_13328,N_10180,N_10681);
xnor U13329 (N_13329,N_11247,N_11626);
nand U13330 (N_13330,N_11050,N_10130);
and U13331 (N_13331,N_10265,N_10998);
xor U13332 (N_13332,N_10639,N_10082);
xor U13333 (N_13333,N_10666,N_11383);
nor U13334 (N_13334,N_10639,N_10253);
or U13335 (N_13335,N_10972,N_10308);
or U13336 (N_13336,N_10955,N_10714);
and U13337 (N_13337,N_10828,N_11578);
nor U13338 (N_13338,N_11132,N_11419);
and U13339 (N_13339,N_11554,N_11542);
and U13340 (N_13340,N_11887,N_10703);
nand U13341 (N_13341,N_10769,N_10199);
nor U13342 (N_13342,N_11234,N_10030);
nand U13343 (N_13343,N_10395,N_11483);
nand U13344 (N_13344,N_11295,N_11891);
nor U13345 (N_13345,N_11463,N_11640);
xnor U13346 (N_13346,N_10760,N_10186);
nand U13347 (N_13347,N_11753,N_11016);
and U13348 (N_13348,N_11165,N_11428);
nand U13349 (N_13349,N_11400,N_11485);
xor U13350 (N_13350,N_10123,N_11859);
and U13351 (N_13351,N_10373,N_10251);
nand U13352 (N_13352,N_10912,N_11295);
or U13353 (N_13353,N_10005,N_11047);
or U13354 (N_13354,N_10078,N_11105);
nand U13355 (N_13355,N_10997,N_10616);
or U13356 (N_13356,N_11245,N_11879);
nor U13357 (N_13357,N_10587,N_10960);
and U13358 (N_13358,N_11417,N_10552);
or U13359 (N_13359,N_11878,N_10602);
and U13360 (N_13360,N_10117,N_11113);
nor U13361 (N_13361,N_11201,N_11551);
nor U13362 (N_13362,N_11644,N_10793);
or U13363 (N_13363,N_10899,N_11038);
nand U13364 (N_13364,N_10421,N_11655);
nand U13365 (N_13365,N_11794,N_10749);
nor U13366 (N_13366,N_10963,N_10685);
and U13367 (N_13367,N_10119,N_10111);
and U13368 (N_13368,N_10727,N_11222);
nor U13369 (N_13369,N_11476,N_10626);
nand U13370 (N_13370,N_11966,N_11589);
or U13371 (N_13371,N_10648,N_10972);
nand U13372 (N_13372,N_11241,N_11044);
or U13373 (N_13373,N_11758,N_10441);
xnor U13374 (N_13374,N_11368,N_10957);
nand U13375 (N_13375,N_11647,N_10923);
or U13376 (N_13376,N_11624,N_11490);
nor U13377 (N_13377,N_11136,N_11217);
xor U13378 (N_13378,N_10064,N_11109);
nor U13379 (N_13379,N_10747,N_10033);
or U13380 (N_13380,N_10521,N_11428);
nand U13381 (N_13381,N_10335,N_10808);
xnor U13382 (N_13382,N_10962,N_11233);
nor U13383 (N_13383,N_10491,N_11979);
or U13384 (N_13384,N_10217,N_11732);
and U13385 (N_13385,N_11746,N_11692);
or U13386 (N_13386,N_11871,N_10402);
or U13387 (N_13387,N_11344,N_11999);
nor U13388 (N_13388,N_11320,N_10270);
nor U13389 (N_13389,N_11506,N_10433);
nand U13390 (N_13390,N_11082,N_11940);
nand U13391 (N_13391,N_11362,N_11194);
nor U13392 (N_13392,N_10435,N_10111);
nand U13393 (N_13393,N_11770,N_10201);
or U13394 (N_13394,N_10714,N_11373);
and U13395 (N_13395,N_10319,N_10099);
nand U13396 (N_13396,N_11515,N_11837);
nand U13397 (N_13397,N_10943,N_11204);
or U13398 (N_13398,N_11358,N_11522);
xor U13399 (N_13399,N_10395,N_10358);
xor U13400 (N_13400,N_11988,N_10885);
and U13401 (N_13401,N_10657,N_10464);
or U13402 (N_13402,N_11119,N_10295);
xor U13403 (N_13403,N_10695,N_10501);
nand U13404 (N_13404,N_10159,N_10897);
nand U13405 (N_13405,N_10061,N_10529);
and U13406 (N_13406,N_10808,N_10591);
nand U13407 (N_13407,N_10874,N_10158);
xnor U13408 (N_13408,N_11602,N_10122);
nand U13409 (N_13409,N_10807,N_10174);
nand U13410 (N_13410,N_11958,N_10008);
nand U13411 (N_13411,N_11009,N_11047);
nand U13412 (N_13412,N_10874,N_10244);
and U13413 (N_13413,N_10807,N_10100);
or U13414 (N_13414,N_10156,N_11992);
and U13415 (N_13415,N_10427,N_10463);
nor U13416 (N_13416,N_10516,N_10857);
nand U13417 (N_13417,N_10992,N_11962);
nor U13418 (N_13418,N_10621,N_11374);
xnor U13419 (N_13419,N_11494,N_11501);
nor U13420 (N_13420,N_10816,N_11058);
or U13421 (N_13421,N_10094,N_10921);
or U13422 (N_13422,N_10750,N_10781);
xnor U13423 (N_13423,N_11745,N_11417);
nand U13424 (N_13424,N_10340,N_10431);
xnor U13425 (N_13425,N_10347,N_10351);
or U13426 (N_13426,N_10894,N_10560);
or U13427 (N_13427,N_11577,N_11119);
nand U13428 (N_13428,N_11303,N_10349);
or U13429 (N_13429,N_10048,N_10980);
or U13430 (N_13430,N_10475,N_10880);
nor U13431 (N_13431,N_11164,N_11934);
or U13432 (N_13432,N_11948,N_10749);
nor U13433 (N_13433,N_10990,N_10929);
nor U13434 (N_13434,N_10252,N_10567);
nor U13435 (N_13435,N_11741,N_10251);
or U13436 (N_13436,N_10850,N_11686);
nor U13437 (N_13437,N_10102,N_10555);
and U13438 (N_13438,N_11343,N_10336);
nor U13439 (N_13439,N_11241,N_11681);
xor U13440 (N_13440,N_10655,N_10336);
and U13441 (N_13441,N_10667,N_11933);
or U13442 (N_13442,N_11315,N_11675);
nor U13443 (N_13443,N_11504,N_11956);
nand U13444 (N_13444,N_10720,N_10079);
nand U13445 (N_13445,N_10272,N_11978);
or U13446 (N_13446,N_11785,N_10959);
nor U13447 (N_13447,N_11677,N_10721);
or U13448 (N_13448,N_10598,N_11395);
and U13449 (N_13449,N_11090,N_10876);
or U13450 (N_13450,N_11554,N_10829);
or U13451 (N_13451,N_11104,N_10978);
nor U13452 (N_13452,N_10749,N_10169);
and U13453 (N_13453,N_10007,N_11905);
nor U13454 (N_13454,N_11850,N_11499);
nand U13455 (N_13455,N_11697,N_11107);
or U13456 (N_13456,N_11805,N_10026);
and U13457 (N_13457,N_11828,N_11757);
xor U13458 (N_13458,N_11386,N_10614);
nand U13459 (N_13459,N_10971,N_10881);
nor U13460 (N_13460,N_10521,N_11414);
nor U13461 (N_13461,N_10196,N_10898);
nor U13462 (N_13462,N_10728,N_11416);
nor U13463 (N_13463,N_10781,N_11701);
nand U13464 (N_13464,N_11605,N_11895);
xor U13465 (N_13465,N_11116,N_10240);
nor U13466 (N_13466,N_11639,N_10074);
and U13467 (N_13467,N_10450,N_10576);
and U13468 (N_13468,N_11346,N_11621);
nor U13469 (N_13469,N_10546,N_11661);
or U13470 (N_13470,N_11618,N_10765);
nor U13471 (N_13471,N_11201,N_10350);
nand U13472 (N_13472,N_11864,N_11605);
or U13473 (N_13473,N_11062,N_11750);
nand U13474 (N_13474,N_11836,N_10240);
and U13475 (N_13475,N_10929,N_10420);
xnor U13476 (N_13476,N_11022,N_10758);
or U13477 (N_13477,N_11116,N_10357);
nor U13478 (N_13478,N_10117,N_11235);
or U13479 (N_13479,N_11939,N_11083);
xor U13480 (N_13480,N_11043,N_11408);
nor U13481 (N_13481,N_11739,N_10028);
nand U13482 (N_13482,N_10520,N_10084);
and U13483 (N_13483,N_11196,N_10747);
or U13484 (N_13484,N_11741,N_11575);
or U13485 (N_13485,N_10876,N_10827);
nor U13486 (N_13486,N_11786,N_10824);
or U13487 (N_13487,N_11210,N_11201);
xor U13488 (N_13488,N_10841,N_10063);
nor U13489 (N_13489,N_11962,N_11581);
nand U13490 (N_13490,N_11667,N_10283);
nor U13491 (N_13491,N_11185,N_11892);
or U13492 (N_13492,N_11322,N_11159);
or U13493 (N_13493,N_11080,N_11157);
and U13494 (N_13494,N_11077,N_10879);
nand U13495 (N_13495,N_11088,N_11766);
xor U13496 (N_13496,N_11140,N_10767);
nor U13497 (N_13497,N_11041,N_10392);
or U13498 (N_13498,N_10607,N_11046);
nand U13499 (N_13499,N_10000,N_11855);
nand U13500 (N_13500,N_11098,N_10581);
or U13501 (N_13501,N_11631,N_10799);
and U13502 (N_13502,N_11881,N_11237);
and U13503 (N_13503,N_11925,N_10395);
and U13504 (N_13504,N_10485,N_10590);
or U13505 (N_13505,N_10172,N_10159);
or U13506 (N_13506,N_11091,N_11718);
or U13507 (N_13507,N_10965,N_11488);
nor U13508 (N_13508,N_10458,N_11442);
xnor U13509 (N_13509,N_10180,N_10400);
xnor U13510 (N_13510,N_11331,N_10605);
xnor U13511 (N_13511,N_11553,N_10436);
nand U13512 (N_13512,N_10180,N_10155);
or U13513 (N_13513,N_10380,N_11451);
and U13514 (N_13514,N_10567,N_10408);
and U13515 (N_13515,N_10212,N_11924);
and U13516 (N_13516,N_10037,N_11385);
or U13517 (N_13517,N_10948,N_11209);
nand U13518 (N_13518,N_11159,N_11774);
or U13519 (N_13519,N_10716,N_11269);
nor U13520 (N_13520,N_11813,N_11189);
nor U13521 (N_13521,N_11708,N_11762);
nand U13522 (N_13522,N_11715,N_10599);
or U13523 (N_13523,N_11626,N_11227);
nor U13524 (N_13524,N_10773,N_11478);
and U13525 (N_13525,N_10919,N_11394);
xnor U13526 (N_13526,N_11312,N_10728);
xnor U13527 (N_13527,N_11830,N_11392);
nand U13528 (N_13528,N_10082,N_10006);
nand U13529 (N_13529,N_10837,N_10860);
and U13530 (N_13530,N_11972,N_10865);
nand U13531 (N_13531,N_10729,N_10056);
nor U13532 (N_13532,N_11179,N_10640);
nand U13533 (N_13533,N_11006,N_11407);
or U13534 (N_13534,N_10441,N_10224);
nand U13535 (N_13535,N_11409,N_11813);
nand U13536 (N_13536,N_11122,N_10420);
nor U13537 (N_13537,N_11515,N_11531);
and U13538 (N_13538,N_11824,N_10550);
or U13539 (N_13539,N_10208,N_11773);
or U13540 (N_13540,N_10405,N_11435);
or U13541 (N_13541,N_10009,N_10256);
and U13542 (N_13542,N_11452,N_10063);
nand U13543 (N_13543,N_11398,N_11570);
nand U13544 (N_13544,N_11658,N_11089);
or U13545 (N_13545,N_11800,N_10164);
nand U13546 (N_13546,N_10276,N_10479);
xor U13547 (N_13547,N_10998,N_10194);
nor U13548 (N_13548,N_10233,N_10900);
and U13549 (N_13549,N_11347,N_10720);
nand U13550 (N_13550,N_11807,N_11531);
nor U13551 (N_13551,N_10599,N_10243);
nor U13552 (N_13552,N_11051,N_10037);
nand U13553 (N_13553,N_10235,N_11177);
xor U13554 (N_13554,N_10625,N_10894);
or U13555 (N_13555,N_11445,N_10343);
nor U13556 (N_13556,N_10463,N_11525);
and U13557 (N_13557,N_10370,N_10931);
xor U13558 (N_13558,N_11647,N_10926);
nor U13559 (N_13559,N_11396,N_10401);
nand U13560 (N_13560,N_11116,N_11051);
nand U13561 (N_13561,N_10474,N_10143);
and U13562 (N_13562,N_10743,N_11648);
xor U13563 (N_13563,N_10714,N_11746);
nand U13564 (N_13564,N_10767,N_10318);
or U13565 (N_13565,N_10047,N_10555);
nand U13566 (N_13566,N_10702,N_11643);
and U13567 (N_13567,N_11685,N_11700);
xnor U13568 (N_13568,N_10009,N_10784);
nand U13569 (N_13569,N_11336,N_11135);
nor U13570 (N_13570,N_10352,N_10268);
or U13571 (N_13571,N_10678,N_11264);
nand U13572 (N_13572,N_10396,N_10041);
nor U13573 (N_13573,N_11357,N_10993);
or U13574 (N_13574,N_11493,N_11667);
nand U13575 (N_13575,N_10573,N_11983);
or U13576 (N_13576,N_10347,N_10068);
nor U13577 (N_13577,N_10233,N_11355);
and U13578 (N_13578,N_10073,N_11876);
nand U13579 (N_13579,N_11947,N_11997);
nor U13580 (N_13580,N_11865,N_10173);
xnor U13581 (N_13581,N_11144,N_11409);
nor U13582 (N_13582,N_10416,N_10793);
xor U13583 (N_13583,N_10428,N_10662);
xor U13584 (N_13584,N_10958,N_10916);
nand U13585 (N_13585,N_10853,N_11405);
or U13586 (N_13586,N_10258,N_11524);
and U13587 (N_13587,N_10740,N_11865);
xnor U13588 (N_13588,N_11974,N_11953);
nor U13589 (N_13589,N_11349,N_11129);
nand U13590 (N_13590,N_10900,N_10817);
nor U13591 (N_13591,N_11699,N_11619);
nand U13592 (N_13592,N_10422,N_11556);
and U13593 (N_13593,N_10512,N_10550);
nor U13594 (N_13594,N_10215,N_11905);
or U13595 (N_13595,N_11216,N_10054);
nor U13596 (N_13596,N_10307,N_11327);
nor U13597 (N_13597,N_11487,N_10277);
or U13598 (N_13598,N_11010,N_11360);
and U13599 (N_13599,N_10364,N_11187);
or U13600 (N_13600,N_11456,N_10370);
or U13601 (N_13601,N_11106,N_11737);
nand U13602 (N_13602,N_10537,N_11180);
or U13603 (N_13603,N_11103,N_10515);
xor U13604 (N_13604,N_11735,N_11026);
xnor U13605 (N_13605,N_10762,N_11575);
nand U13606 (N_13606,N_10827,N_10013);
nor U13607 (N_13607,N_10062,N_11987);
and U13608 (N_13608,N_10369,N_11838);
or U13609 (N_13609,N_10276,N_10100);
or U13610 (N_13610,N_10381,N_11912);
and U13611 (N_13611,N_11693,N_11057);
xor U13612 (N_13612,N_11968,N_10495);
nand U13613 (N_13613,N_11285,N_10158);
nand U13614 (N_13614,N_10708,N_11571);
or U13615 (N_13615,N_11312,N_10231);
nand U13616 (N_13616,N_11823,N_10197);
and U13617 (N_13617,N_10306,N_11878);
nor U13618 (N_13618,N_10557,N_11968);
or U13619 (N_13619,N_10705,N_10044);
xnor U13620 (N_13620,N_11180,N_10610);
and U13621 (N_13621,N_10477,N_10379);
and U13622 (N_13622,N_10373,N_10241);
or U13623 (N_13623,N_11131,N_10309);
and U13624 (N_13624,N_11245,N_11582);
nor U13625 (N_13625,N_11083,N_11977);
and U13626 (N_13626,N_11633,N_10277);
or U13627 (N_13627,N_11446,N_11271);
or U13628 (N_13628,N_10790,N_11070);
and U13629 (N_13629,N_11181,N_10105);
nand U13630 (N_13630,N_11195,N_10076);
or U13631 (N_13631,N_11609,N_11678);
xor U13632 (N_13632,N_10225,N_11517);
and U13633 (N_13633,N_10744,N_11211);
and U13634 (N_13634,N_11198,N_10664);
and U13635 (N_13635,N_11964,N_11081);
nand U13636 (N_13636,N_10598,N_10148);
and U13637 (N_13637,N_10529,N_11799);
nand U13638 (N_13638,N_10411,N_10012);
nor U13639 (N_13639,N_11710,N_10543);
nand U13640 (N_13640,N_10636,N_10115);
nand U13641 (N_13641,N_10919,N_10165);
xor U13642 (N_13642,N_10562,N_11327);
xnor U13643 (N_13643,N_11713,N_10082);
nand U13644 (N_13644,N_10261,N_11504);
or U13645 (N_13645,N_10415,N_11603);
xnor U13646 (N_13646,N_11929,N_10397);
and U13647 (N_13647,N_10420,N_10358);
xor U13648 (N_13648,N_11189,N_10028);
or U13649 (N_13649,N_10500,N_11398);
nand U13650 (N_13650,N_10442,N_10664);
nand U13651 (N_13651,N_11114,N_11111);
and U13652 (N_13652,N_11811,N_11336);
and U13653 (N_13653,N_11094,N_11766);
and U13654 (N_13654,N_10841,N_11062);
nor U13655 (N_13655,N_10832,N_11748);
nand U13656 (N_13656,N_10860,N_10478);
or U13657 (N_13657,N_11053,N_11821);
nor U13658 (N_13658,N_11273,N_10594);
and U13659 (N_13659,N_11218,N_11924);
nor U13660 (N_13660,N_10643,N_10658);
and U13661 (N_13661,N_10337,N_10477);
nor U13662 (N_13662,N_11786,N_11662);
nand U13663 (N_13663,N_11803,N_11736);
and U13664 (N_13664,N_10282,N_10129);
xor U13665 (N_13665,N_10879,N_11240);
nand U13666 (N_13666,N_10177,N_10580);
or U13667 (N_13667,N_10590,N_11571);
nand U13668 (N_13668,N_10212,N_10465);
or U13669 (N_13669,N_10394,N_11700);
and U13670 (N_13670,N_10801,N_11994);
xor U13671 (N_13671,N_10341,N_10982);
nor U13672 (N_13672,N_10635,N_10005);
nand U13673 (N_13673,N_10873,N_11627);
xor U13674 (N_13674,N_10452,N_10164);
and U13675 (N_13675,N_10110,N_11744);
nor U13676 (N_13676,N_10621,N_10458);
or U13677 (N_13677,N_11757,N_11873);
nand U13678 (N_13678,N_10132,N_11819);
nand U13679 (N_13679,N_10677,N_11084);
nand U13680 (N_13680,N_10009,N_10907);
nor U13681 (N_13681,N_11859,N_11168);
nor U13682 (N_13682,N_11651,N_10647);
nor U13683 (N_13683,N_11922,N_11379);
or U13684 (N_13684,N_10847,N_11444);
or U13685 (N_13685,N_11836,N_10824);
or U13686 (N_13686,N_11406,N_11311);
nand U13687 (N_13687,N_11239,N_11225);
nor U13688 (N_13688,N_11688,N_11262);
or U13689 (N_13689,N_11954,N_10155);
and U13690 (N_13690,N_11500,N_11156);
or U13691 (N_13691,N_10427,N_10303);
nand U13692 (N_13692,N_11140,N_10959);
or U13693 (N_13693,N_11398,N_10282);
and U13694 (N_13694,N_11157,N_10456);
xnor U13695 (N_13695,N_10508,N_10130);
and U13696 (N_13696,N_11883,N_10630);
nand U13697 (N_13697,N_10357,N_11333);
nor U13698 (N_13698,N_11742,N_10125);
or U13699 (N_13699,N_10973,N_10584);
or U13700 (N_13700,N_11008,N_10229);
or U13701 (N_13701,N_10272,N_10233);
nand U13702 (N_13702,N_11575,N_11259);
nor U13703 (N_13703,N_10944,N_11661);
nor U13704 (N_13704,N_10924,N_11491);
and U13705 (N_13705,N_10565,N_10078);
and U13706 (N_13706,N_11069,N_10817);
xor U13707 (N_13707,N_10730,N_11569);
nor U13708 (N_13708,N_10662,N_10414);
and U13709 (N_13709,N_10332,N_11396);
nor U13710 (N_13710,N_10483,N_10427);
nor U13711 (N_13711,N_10369,N_11958);
nand U13712 (N_13712,N_11913,N_11827);
xnor U13713 (N_13713,N_11414,N_11276);
and U13714 (N_13714,N_10804,N_11261);
xnor U13715 (N_13715,N_10421,N_10973);
nand U13716 (N_13716,N_10963,N_10217);
or U13717 (N_13717,N_10233,N_11081);
nor U13718 (N_13718,N_10965,N_10681);
or U13719 (N_13719,N_11785,N_10619);
nor U13720 (N_13720,N_10061,N_11543);
nand U13721 (N_13721,N_11587,N_10111);
and U13722 (N_13722,N_11589,N_11344);
and U13723 (N_13723,N_10590,N_11260);
or U13724 (N_13724,N_11164,N_11258);
nand U13725 (N_13725,N_10638,N_10011);
nor U13726 (N_13726,N_11439,N_10221);
xor U13727 (N_13727,N_10669,N_10515);
nor U13728 (N_13728,N_11282,N_10472);
nand U13729 (N_13729,N_11703,N_10875);
nor U13730 (N_13730,N_11217,N_11829);
xnor U13731 (N_13731,N_10805,N_10103);
and U13732 (N_13732,N_10417,N_10534);
and U13733 (N_13733,N_11755,N_11545);
nand U13734 (N_13734,N_10337,N_11565);
xor U13735 (N_13735,N_10788,N_10655);
xor U13736 (N_13736,N_10514,N_11560);
or U13737 (N_13737,N_10792,N_11998);
nand U13738 (N_13738,N_10235,N_10464);
and U13739 (N_13739,N_11857,N_10660);
nand U13740 (N_13740,N_11509,N_11649);
or U13741 (N_13741,N_10653,N_11263);
xor U13742 (N_13742,N_11032,N_10038);
and U13743 (N_13743,N_11429,N_10014);
and U13744 (N_13744,N_10486,N_10049);
or U13745 (N_13745,N_10384,N_10377);
nor U13746 (N_13746,N_10901,N_10502);
and U13747 (N_13747,N_11764,N_11651);
nand U13748 (N_13748,N_10193,N_11884);
and U13749 (N_13749,N_11357,N_11619);
and U13750 (N_13750,N_10089,N_10460);
or U13751 (N_13751,N_10951,N_10118);
nand U13752 (N_13752,N_11063,N_11497);
or U13753 (N_13753,N_11986,N_10714);
nor U13754 (N_13754,N_11610,N_11944);
or U13755 (N_13755,N_10530,N_10899);
nor U13756 (N_13756,N_11381,N_11954);
or U13757 (N_13757,N_11827,N_10317);
nor U13758 (N_13758,N_10786,N_10051);
or U13759 (N_13759,N_11440,N_10751);
or U13760 (N_13760,N_10069,N_10666);
nand U13761 (N_13761,N_10629,N_10577);
and U13762 (N_13762,N_10135,N_10868);
nor U13763 (N_13763,N_10250,N_10410);
nor U13764 (N_13764,N_10718,N_11245);
nand U13765 (N_13765,N_11410,N_10251);
and U13766 (N_13766,N_11523,N_11980);
and U13767 (N_13767,N_10046,N_11823);
nand U13768 (N_13768,N_10696,N_11344);
xor U13769 (N_13769,N_10347,N_10222);
nand U13770 (N_13770,N_11239,N_11240);
and U13771 (N_13771,N_10170,N_11396);
or U13772 (N_13772,N_11020,N_10232);
nand U13773 (N_13773,N_10328,N_11473);
or U13774 (N_13774,N_10835,N_10343);
nand U13775 (N_13775,N_10036,N_10775);
and U13776 (N_13776,N_11162,N_11056);
xor U13777 (N_13777,N_10166,N_10489);
nor U13778 (N_13778,N_10690,N_11154);
nand U13779 (N_13779,N_11410,N_11927);
nand U13780 (N_13780,N_10449,N_11143);
or U13781 (N_13781,N_11696,N_10090);
nor U13782 (N_13782,N_11311,N_11889);
and U13783 (N_13783,N_11039,N_10470);
or U13784 (N_13784,N_11324,N_10692);
and U13785 (N_13785,N_10179,N_10385);
or U13786 (N_13786,N_10031,N_11106);
nand U13787 (N_13787,N_10707,N_10763);
and U13788 (N_13788,N_11225,N_10889);
nand U13789 (N_13789,N_10973,N_10238);
and U13790 (N_13790,N_10598,N_11423);
or U13791 (N_13791,N_11296,N_10196);
nand U13792 (N_13792,N_10091,N_10907);
or U13793 (N_13793,N_11623,N_11884);
and U13794 (N_13794,N_11672,N_10742);
xnor U13795 (N_13795,N_10025,N_11443);
nand U13796 (N_13796,N_11850,N_10244);
and U13797 (N_13797,N_11958,N_10632);
nor U13798 (N_13798,N_10101,N_11730);
nand U13799 (N_13799,N_11711,N_11007);
and U13800 (N_13800,N_10114,N_11741);
and U13801 (N_13801,N_10316,N_10452);
and U13802 (N_13802,N_10289,N_10141);
nor U13803 (N_13803,N_10939,N_11882);
and U13804 (N_13804,N_10588,N_10691);
nand U13805 (N_13805,N_11386,N_11854);
and U13806 (N_13806,N_11694,N_11916);
nor U13807 (N_13807,N_10432,N_11501);
or U13808 (N_13808,N_10298,N_11064);
nand U13809 (N_13809,N_11540,N_11245);
nand U13810 (N_13810,N_11581,N_11907);
and U13811 (N_13811,N_11083,N_10201);
and U13812 (N_13812,N_10873,N_10190);
or U13813 (N_13813,N_10656,N_10983);
and U13814 (N_13814,N_10842,N_11037);
or U13815 (N_13815,N_11279,N_10034);
nand U13816 (N_13816,N_10929,N_11512);
or U13817 (N_13817,N_10688,N_11880);
or U13818 (N_13818,N_11112,N_11772);
nor U13819 (N_13819,N_11374,N_11555);
nor U13820 (N_13820,N_11600,N_11562);
or U13821 (N_13821,N_11356,N_11088);
or U13822 (N_13822,N_10523,N_11868);
or U13823 (N_13823,N_11324,N_11115);
nor U13824 (N_13824,N_11056,N_11917);
or U13825 (N_13825,N_11731,N_10187);
nor U13826 (N_13826,N_11367,N_10607);
and U13827 (N_13827,N_10218,N_11542);
nor U13828 (N_13828,N_11671,N_10399);
nand U13829 (N_13829,N_11902,N_11822);
or U13830 (N_13830,N_10132,N_11428);
and U13831 (N_13831,N_10347,N_10283);
nand U13832 (N_13832,N_11920,N_10838);
nand U13833 (N_13833,N_10749,N_10653);
nand U13834 (N_13834,N_10379,N_10197);
and U13835 (N_13835,N_10577,N_10364);
or U13836 (N_13836,N_11345,N_11398);
nor U13837 (N_13837,N_10920,N_10847);
xor U13838 (N_13838,N_11767,N_10759);
nand U13839 (N_13839,N_11819,N_10619);
xor U13840 (N_13840,N_10164,N_11358);
nor U13841 (N_13841,N_10976,N_11697);
and U13842 (N_13842,N_10024,N_10935);
nor U13843 (N_13843,N_11727,N_10387);
nor U13844 (N_13844,N_10174,N_11488);
or U13845 (N_13845,N_10335,N_11260);
nand U13846 (N_13846,N_11300,N_11870);
xor U13847 (N_13847,N_11461,N_10864);
xnor U13848 (N_13848,N_10361,N_11189);
nand U13849 (N_13849,N_10000,N_10394);
nand U13850 (N_13850,N_11710,N_11008);
or U13851 (N_13851,N_11317,N_11185);
xnor U13852 (N_13852,N_10757,N_10730);
nor U13853 (N_13853,N_11204,N_10324);
nor U13854 (N_13854,N_11035,N_11467);
or U13855 (N_13855,N_11074,N_11768);
and U13856 (N_13856,N_11321,N_10361);
and U13857 (N_13857,N_11123,N_10256);
nand U13858 (N_13858,N_11751,N_11705);
nand U13859 (N_13859,N_10686,N_10164);
or U13860 (N_13860,N_10465,N_11562);
or U13861 (N_13861,N_10521,N_11023);
nor U13862 (N_13862,N_11364,N_10985);
and U13863 (N_13863,N_11182,N_10956);
nand U13864 (N_13864,N_10033,N_10830);
xnor U13865 (N_13865,N_11122,N_11080);
nand U13866 (N_13866,N_11726,N_10197);
nor U13867 (N_13867,N_10345,N_11083);
nand U13868 (N_13868,N_11496,N_11324);
nand U13869 (N_13869,N_10002,N_11909);
nor U13870 (N_13870,N_11169,N_10405);
nor U13871 (N_13871,N_11649,N_11101);
nand U13872 (N_13872,N_10724,N_10457);
nand U13873 (N_13873,N_10487,N_10340);
nand U13874 (N_13874,N_11579,N_10091);
or U13875 (N_13875,N_11615,N_11409);
nand U13876 (N_13876,N_10634,N_10787);
nand U13877 (N_13877,N_10160,N_11293);
or U13878 (N_13878,N_11821,N_11891);
or U13879 (N_13879,N_10663,N_11398);
and U13880 (N_13880,N_10850,N_10837);
and U13881 (N_13881,N_10057,N_11232);
or U13882 (N_13882,N_10291,N_11287);
nor U13883 (N_13883,N_10949,N_11284);
nand U13884 (N_13884,N_10157,N_10812);
nand U13885 (N_13885,N_10644,N_10796);
or U13886 (N_13886,N_11315,N_11735);
or U13887 (N_13887,N_11473,N_11608);
and U13888 (N_13888,N_10583,N_10664);
and U13889 (N_13889,N_10156,N_11661);
or U13890 (N_13890,N_10115,N_11816);
nor U13891 (N_13891,N_10948,N_10174);
nand U13892 (N_13892,N_11378,N_10958);
nor U13893 (N_13893,N_10374,N_10190);
and U13894 (N_13894,N_10368,N_11330);
and U13895 (N_13895,N_11031,N_11366);
nor U13896 (N_13896,N_10929,N_11980);
or U13897 (N_13897,N_10441,N_10112);
nor U13898 (N_13898,N_11867,N_11112);
nand U13899 (N_13899,N_11190,N_11723);
nor U13900 (N_13900,N_10745,N_11932);
and U13901 (N_13901,N_11660,N_10038);
or U13902 (N_13902,N_10549,N_10461);
or U13903 (N_13903,N_10573,N_11345);
nor U13904 (N_13904,N_10758,N_11269);
or U13905 (N_13905,N_11680,N_10022);
nand U13906 (N_13906,N_11840,N_10865);
nor U13907 (N_13907,N_11584,N_11224);
and U13908 (N_13908,N_11949,N_10891);
nand U13909 (N_13909,N_10362,N_10814);
and U13910 (N_13910,N_11162,N_10571);
or U13911 (N_13911,N_10384,N_11851);
or U13912 (N_13912,N_11524,N_10709);
or U13913 (N_13913,N_11687,N_11077);
xnor U13914 (N_13914,N_11201,N_11082);
xor U13915 (N_13915,N_10163,N_10541);
and U13916 (N_13916,N_11879,N_11036);
or U13917 (N_13917,N_10413,N_11198);
nor U13918 (N_13918,N_10274,N_10884);
nand U13919 (N_13919,N_10176,N_11818);
and U13920 (N_13920,N_11849,N_10099);
xnor U13921 (N_13921,N_11694,N_11075);
or U13922 (N_13922,N_10257,N_11512);
nor U13923 (N_13923,N_10782,N_10611);
or U13924 (N_13924,N_11330,N_10052);
and U13925 (N_13925,N_11933,N_10584);
and U13926 (N_13926,N_10082,N_10979);
nand U13927 (N_13927,N_11174,N_11813);
or U13928 (N_13928,N_10342,N_11894);
nand U13929 (N_13929,N_11688,N_10416);
or U13930 (N_13930,N_10809,N_11069);
or U13931 (N_13931,N_10551,N_11059);
nor U13932 (N_13932,N_10148,N_10828);
xnor U13933 (N_13933,N_10364,N_11232);
or U13934 (N_13934,N_11753,N_11172);
nand U13935 (N_13935,N_11678,N_10036);
or U13936 (N_13936,N_10467,N_11211);
and U13937 (N_13937,N_11150,N_10533);
nand U13938 (N_13938,N_11533,N_10453);
nor U13939 (N_13939,N_10769,N_10817);
or U13940 (N_13940,N_10327,N_11946);
xnor U13941 (N_13941,N_10493,N_11984);
or U13942 (N_13942,N_11072,N_10822);
and U13943 (N_13943,N_10218,N_10111);
xnor U13944 (N_13944,N_10318,N_10203);
nor U13945 (N_13945,N_11918,N_10086);
or U13946 (N_13946,N_11156,N_10450);
or U13947 (N_13947,N_11773,N_11284);
or U13948 (N_13948,N_10450,N_10712);
or U13949 (N_13949,N_11979,N_11793);
nor U13950 (N_13950,N_10905,N_10565);
or U13951 (N_13951,N_11145,N_11013);
nand U13952 (N_13952,N_10076,N_10513);
or U13953 (N_13953,N_11167,N_10297);
and U13954 (N_13954,N_11810,N_11198);
or U13955 (N_13955,N_10966,N_11781);
nor U13956 (N_13956,N_10975,N_10237);
nand U13957 (N_13957,N_11391,N_10111);
nand U13958 (N_13958,N_11030,N_10438);
or U13959 (N_13959,N_10881,N_11571);
xnor U13960 (N_13960,N_10157,N_11922);
nand U13961 (N_13961,N_11795,N_10034);
nand U13962 (N_13962,N_11609,N_11790);
nor U13963 (N_13963,N_10689,N_10195);
or U13964 (N_13964,N_10464,N_11493);
xnor U13965 (N_13965,N_11763,N_11463);
xnor U13966 (N_13966,N_10458,N_11686);
or U13967 (N_13967,N_11867,N_11900);
nand U13968 (N_13968,N_10349,N_10267);
or U13969 (N_13969,N_10970,N_11131);
or U13970 (N_13970,N_11302,N_10491);
xor U13971 (N_13971,N_11109,N_11726);
or U13972 (N_13972,N_10997,N_11229);
nand U13973 (N_13973,N_11006,N_11023);
or U13974 (N_13974,N_11084,N_10586);
and U13975 (N_13975,N_11782,N_11437);
nand U13976 (N_13976,N_10817,N_10288);
and U13977 (N_13977,N_10968,N_11958);
and U13978 (N_13978,N_11153,N_10402);
or U13979 (N_13979,N_10224,N_10907);
nand U13980 (N_13980,N_11815,N_10934);
or U13981 (N_13981,N_11903,N_11072);
and U13982 (N_13982,N_10446,N_10624);
or U13983 (N_13983,N_11650,N_11730);
nand U13984 (N_13984,N_11923,N_11842);
xor U13985 (N_13985,N_10752,N_10064);
nor U13986 (N_13986,N_11809,N_11756);
nand U13987 (N_13987,N_10869,N_10909);
nand U13988 (N_13988,N_11131,N_11004);
and U13989 (N_13989,N_11489,N_11195);
xor U13990 (N_13990,N_10092,N_11063);
and U13991 (N_13991,N_11949,N_10878);
nand U13992 (N_13992,N_11109,N_11705);
xnor U13993 (N_13993,N_11180,N_11096);
nand U13994 (N_13994,N_11453,N_11333);
nand U13995 (N_13995,N_10282,N_11711);
nand U13996 (N_13996,N_11910,N_10098);
nand U13997 (N_13997,N_11406,N_11801);
nor U13998 (N_13998,N_10413,N_10666);
nand U13999 (N_13999,N_11606,N_11948);
nor U14000 (N_14000,N_13997,N_12060);
nor U14001 (N_14001,N_12618,N_12321);
or U14002 (N_14002,N_12304,N_12868);
nand U14003 (N_14003,N_13383,N_13066);
xor U14004 (N_14004,N_13526,N_12359);
or U14005 (N_14005,N_12463,N_13046);
and U14006 (N_14006,N_12262,N_13270);
nor U14007 (N_14007,N_13223,N_12890);
nor U14008 (N_14008,N_12358,N_13670);
nand U14009 (N_14009,N_13589,N_13178);
nand U14010 (N_14010,N_12700,N_13217);
nor U14011 (N_14011,N_12987,N_13604);
nor U14012 (N_14012,N_13434,N_12922);
or U14013 (N_14013,N_13780,N_12442);
and U14014 (N_14014,N_12169,N_12722);
nand U14015 (N_14015,N_13613,N_12324);
nor U14016 (N_14016,N_12962,N_13527);
nand U14017 (N_14017,N_13645,N_13213);
nand U14018 (N_14018,N_12325,N_12125);
nor U14019 (N_14019,N_12078,N_12456);
nand U14020 (N_14020,N_13982,N_12228);
or U14021 (N_14021,N_13584,N_13159);
nand U14022 (N_14022,N_13449,N_13784);
or U14023 (N_14023,N_13720,N_13336);
xor U14024 (N_14024,N_13629,N_12626);
xor U14025 (N_14025,N_12160,N_12167);
nand U14026 (N_14026,N_13539,N_12527);
and U14027 (N_14027,N_13960,N_13889);
nand U14028 (N_14028,N_12027,N_12586);
nor U14029 (N_14029,N_12427,N_13090);
or U14030 (N_14030,N_12180,N_12815);
and U14031 (N_14031,N_12773,N_13109);
nand U14032 (N_14032,N_12067,N_12541);
nand U14033 (N_14033,N_12149,N_12222);
nor U14034 (N_14034,N_13632,N_12485);
or U14035 (N_14035,N_13360,N_12431);
xor U14036 (N_14036,N_13320,N_13023);
and U14037 (N_14037,N_12253,N_13516);
or U14038 (N_14038,N_12942,N_13609);
nand U14039 (N_14039,N_13452,N_13549);
and U14040 (N_14040,N_13536,N_13212);
nand U14041 (N_14041,N_12164,N_12166);
or U14042 (N_14042,N_12202,N_13104);
or U14043 (N_14043,N_12246,N_13768);
and U14044 (N_14044,N_13278,N_13196);
nor U14045 (N_14045,N_13339,N_12749);
nor U14046 (N_14046,N_13332,N_13728);
nand U14047 (N_14047,N_13802,N_13369);
nand U14048 (N_14048,N_13255,N_12483);
nand U14049 (N_14049,N_12363,N_13510);
and U14050 (N_14050,N_13073,N_13863);
or U14051 (N_14051,N_12353,N_12683);
nand U14052 (N_14052,N_13558,N_13416);
xor U14053 (N_14053,N_13330,N_13357);
nand U14054 (N_14054,N_13136,N_12490);
nor U14055 (N_14055,N_13776,N_13207);
or U14056 (N_14056,N_13253,N_13752);
nand U14057 (N_14057,N_13583,N_12197);
nor U14058 (N_14058,N_12913,N_12053);
or U14059 (N_14059,N_13145,N_12404);
nand U14060 (N_14060,N_13729,N_13884);
nor U14061 (N_14061,N_13831,N_12981);
or U14062 (N_14062,N_13491,N_12388);
nor U14063 (N_14063,N_12860,N_12723);
nor U14064 (N_14064,N_13610,N_12178);
or U14065 (N_14065,N_13210,N_13545);
nand U14066 (N_14066,N_13343,N_12608);
xnor U14067 (N_14067,N_12699,N_13512);
nand U14068 (N_14068,N_13035,N_13625);
and U14069 (N_14069,N_12235,N_12903);
nand U14070 (N_14070,N_13075,N_13064);
or U14071 (N_14071,N_12924,N_12093);
or U14072 (N_14072,N_12745,N_12521);
nor U14073 (N_14073,N_13256,N_12017);
or U14074 (N_14074,N_13461,N_12571);
or U14075 (N_14075,N_12667,N_13774);
xnor U14076 (N_14076,N_13592,N_13521);
and U14077 (N_14077,N_13514,N_13171);
or U14078 (N_14078,N_12374,N_12911);
nor U14079 (N_14079,N_13546,N_13590);
nand U14080 (N_14080,N_13254,N_13303);
and U14081 (N_14081,N_13968,N_12738);
nor U14082 (N_14082,N_13081,N_13766);
nor U14083 (N_14083,N_13115,N_13707);
xor U14084 (N_14084,N_13097,N_13523);
nand U14085 (N_14085,N_12835,N_12020);
nand U14086 (N_14086,N_12518,N_12289);
or U14087 (N_14087,N_12494,N_12439);
nand U14088 (N_14088,N_13458,N_12665);
or U14089 (N_14089,N_13231,N_13849);
xor U14090 (N_14090,N_12988,N_13628);
nor U14091 (N_14091,N_12677,N_13445);
or U14092 (N_14092,N_13305,N_12550);
or U14093 (N_14093,N_12947,N_13271);
xor U14094 (N_14094,N_13448,N_12487);
nand U14095 (N_14095,N_13442,N_13074);
xor U14096 (N_14096,N_13465,N_12024);
xor U14097 (N_14097,N_13300,N_12796);
or U14098 (N_14098,N_13718,N_13499);
nand U14099 (N_14099,N_12548,N_12781);
nand U14100 (N_14100,N_13635,N_12225);
nand U14101 (N_14101,N_13500,N_13857);
and U14102 (N_14102,N_12239,N_13466);
or U14103 (N_14103,N_13597,N_13358);
nor U14104 (N_14104,N_12785,N_12214);
and U14105 (N_14105,N_13006,N_12696);
and U14106 (N_14106,N_13160,N_12399);
xor U14107 (N_14107,N_12118,N_12416);
nand U14108 (N_14108,N_12464,N_13709);
and U14109 (N_14109,N_12445,N_12173);
and U14110 (N_14110,N_13966,N_12659);
or U14111 (N_14111,N_12660,N_13887);
nor U14112 (N_14112,N_13148,N_13352);
xor U14113 (N_14113,N_13385,N_13748);
and U14114 (N_14114,N_13289,N_12418);
nand U14115 (N_14115,N_13881,N_12087);
and U14116 (N_14116,N_13276,N_12816);
nand U14117 (N_14117,N_12718,N_12443);
or U14118 (N_14118,N_12254,N_12621);
nor U14119 (N_14119,N_13475,N_12342);
or U14120 (N_14120,N_13192,N_12278);
or U14121 (N_14121,N_13436,N_12480);
or U14122 (N_14122,N_12457,N_13002);
nand U14123 (N_14123,N_13916,N_12244);
or U14124 (N_14124,N_13167,N_13076);
nand U14125 (N_14125,N_12129,N_13891);
and U14126 (N_14126,N_12127,N_12858);
nand U14127 (N_14127,N_13013,N_12838);
nand U14128 (N_14128,N_13743,N_13586);
and U14129 (N_14129,N_12831,N_12113);
nor U14130 (N_14130,N_12505,N_12146);
nor U14131 (N_14131,N_12959,N_13649);
and U14132 (N_14132,N_12467,N_12850);
xor U14133 (N_14133,N_12578,N_13415);
nor U14134 (N_14134,N_12181,N_13946);
or U14135 (N_14135,N_13754,N_13783);
or U14136 (N_14136,N_13308,N_12729);
nand U14137 (N_14137,N_12137,N_12623);
or U14138 (N_14138,N_12797,N_13390);
nor U14139 (N_14139,N_12640,N_12206);
nand U14140 (N_14140,N_12165,N_13479);
xnor U14141 (N_14141,N_13667,N_13556);
xnor U14142 (N_14142,N_12685,N_13280);
or U14143 (N_14143,N_12389,N_13812);
nor U14144 (N_14144,N_12309,N_13184);
nor U14145 (N_14145,N_12647,N_12896);
nand U14146 (N_14146,N_13298,N_12375);
or U14147 (N_14147,N_12603,N_12284);
nand U14148 (N_14148,N_12587,N_13681);
and U14149 (N_14149,N_12780,N_12282);
or U14150 (N_14150,N_13806,N_12543);
or U14151 (N_14151,N_13439,N_12465);
or U14152 (N_14152,N_12939,N_12308);
or U14153 (N_14153,N_12934,N_12866);
nand U14154 (N_14154,N_13935,N_13165);
nor U14155 (N_14155,N_13483,N_12819);
xnor U14156 (N_14156,N_12522,N_12614);
or U14157 (N_14157,N_13422,N_12386);
or U14158 (N_14158,N_12861,N_13932);
nand U14159 (N_14159,N_13325,N_13842);
and U14160 (N_14160,N_13333,N_12403);
and U14161 (N_14161,N_13984,N_13582);
nor U14162 (N_14162,N_12136,N_13092);
nand U14163 (N_14163,N_13905,N_12168);
or U14164 (N_14164,N_13426,N_12714);
nor U14165 (N_14165,N_13273,N_13474);
and U14166 (N_14166,N_12724,N_13713);
and U14167 (N_14167,N_13125,N_12744);
nand U14168 (N_14168,N_13789,N_12739);
nor U14169 (N_14169,N_13039,N_13811);
xor U14170 (N_14170,N_12596,N_12678);
or U14171 (N_14171,N_13187,N_13961);
or U14172 (N_14172,N_12430,N_13740);
or U14173 (N_14173,N_12134,N_12589);
or U14174 (N_14174,N_12591,N_13703);
nor U14175 (N_14175,N_13004,N_13532);
nor U14176 (N_14176,N_12184,N_13793);
or U14177 (N_14177,N_12385,N_12459);
and U14178 (N_14178,N_12792,N_13381);
nor U14179 (N_14179,N_12128,N_13569);
or U14180 (N_14180,N_13940,N_12142);
nor U14181 (N_14181,N_12346,N_12516);
or U14182 (N_14182,N_12095,N_12994);
or U14183 (N_14183,N_12126,N_12069);
and U14184 (N_14184,N_13991,N_13007);
and U14185 (N_14185,N_12728,N_13790);
and U14186 (N_14186,N_12867,N_13561);
or U14187 (N_14187,N_13575,N_12848);
nor U14188 (N_14188,N_12863,N_13648);
or U14189 (N_14189,N_13430,N_13211);
nor U14190 (N_14190,N_12271,N_12657);
nand U14191 (N_14191,N_12419,N_13673);
xnor U14192 (N_14192,N_13193,N_12658);
or U14193 (N_14193,N_13131,N_13833);
or U14194 (N_14194,N_12561,N_13796);
and U14195 (N_14195,N_12098,N_12566);
or U14196 (N_14196,N_13655,N_12688);
and U14197 (N_14197,N_13151,N_12472);
or U14198 (N_14198,N_12157,N_12115);
nor U14199 (N_14199,N_12805,N_13501);
xnor U14200 (N_14200,N_13118,N_12650);
or U14201 (N_14201,N_13447,N_13099);
or U14202 (N_14202,N_12758,N_13631);
xor U14203 (N_14203,N_12452,N_13990);
or U14204 (N_14204,N_12510,N_13137);
nand U14205 (N_14205,N_12140,N_13800);
nand U14206 (N_14206,N_12670,N_12899);
or U14207 (N_14207,N_12424,N_13978);
nand U14208 (N_14208,N_12662,N_13065);
nand U14209 (N_14209,N_12508,N_12967);
nor U14210 (N_14210,N_12634,N_12288);
xor U14211 (N_14211,N_13386,N_13607);
or U14212 (N_14212,N_13233,N_13660);
nand U14213 (N_14213,N_13056,N_12035);
nand U14214 (N_14214,N_13816,N_13245);
nand U14215 (N_14215,N_12022,N_12782);
and U14216 (N_14216,N_12366,N_13127);
nand U14217 (N_14217,N_12597,N_13251);
or U14218 (N_14218,N_13885,N_13967);
nor U14219 (N_14219,N_13094,N_13019);
xor U14220 (N_14220,N_12349,N_12551);
nand U14221 (N_14221,N_13457,N_12364);
nand U14222 (N_14222,N_13563,N_12393);
xnor U14223 (N_14223,N_13577,N_12847);
nand U14224 (N_14224,N_12595,N_13146);
or U14225 (N_14225,N_12094,N_13996);
and U14226 (N_14226,N_13739,N_12025);
nand U14227 (N_14227,N_12513,N_12730);
or U14228 (N_14228,N_13764,N_12074);
and U14229 (N_14229,N_12630,N_13408);
nand U14230 (N_14230,N_13181,N_13185);
or U14231 (N_14231,N_13221,N_13808);
and U14232 (N_14232,N_13825,N_13375);
or U14233 (N_14233,N_13587,N_13998);
and U14234 (N_14234,N_13071,N_13105);
nand U14235 (N_14235,N_13494,N_12061);
nor U14236 (N_14236,N_12317,N_13531);
nor U14237 (N_14237,N_13696,N_12041);
and U14238 (N_14238,N_12036,N_13888);
nand U14239 (N_14239,N_12466,N_13334);
nand U14240 (N_14240,N_13096,N_13814);
or U14241 (N_14241,N_12663,N_13611);
nand U14242 (N_14242,N_12577,N_12295);
and U14243 (N_14243,N_13620,N_13044);
or U14244 (N_14244,N_12592,N_13116);
or U14245 (N_14245,N_13172,N_12536);
and U14246 (N_14246,N_13072,N_13453);
nand U14247 (N_14247,N_13481,N_13335);
nand U14248 (N_14248,N_12798,N_13355);
and U14249 (N_14249,N_12016,N_12365);
nor U14250 (N_14250,N_12776,N_13043);
and U14251 (N_14251,N_12382,N_13508);
and U14252 (N_14252,N_13683,N_13286);
nand U14253 (N_14253,N_12904,N_13674);
and U14254 (N_14254,N_12175,N_13837);
nor U14255 (N_14255,N_12671,N_13139);
and U14256 (N_14256,N_13511,N_13183);
nor U14257 (N_14257,N_13818,N_12477);
nor U14258 (N_14258,N_13003,N_12644);
and U14259 (N_14259,N_12669,N_13147);
and U14260 (N_14260,N_13287,N_12379);
and U14261 (N_14261,N_12664,N_12279);
nor U14262 (N_14262,N_13867,N_13626);
or U14263 (N_14263,N_12322,N_13656);
or U14264 (N_14264,N_12361,N_12726);
nand U14265 (N_14265,N_13898,N_13711);
or U14266 (N_14266,N_12555,N_13755);
nand U14267 (N_14267,N_12461,N_13069);
xnor U14268 (N_14268,N_12841,N_13896);
or U14269 (N_14269,N_12769,N_13292);
or U14270 (N_14270,N_13679,N_12190);
and U14271 (N_14271,N_13809,N_12559);
nand U14272 (N_14272,N_13522,N_13637);
or U14273 (N_14273,N_12676,N_13269);
or U14274 (N_14274,N_12232,N_12408);
nand U14275 (N_14275,N_13395,N_13082);
and U14276 (N_14276,N_12192,N_12145);
and U14277 (N_14277,N_12938,N_13616);
and U14278 (N_14278,N_12417,N_12252);
nor U14279 (N_14279,N_12802,N_13150);
nand U14280 (N_14280,N_12207,N_13744);
or U14281 (N_14281,N_12048,N_12553);
nor U14282 (N_14282,N_12707,N_12743);
and U14283 (N_14283,N_13588,N_12809);
xor U14284 (N_14284,N_13591,N_12854);
nand U14285 (N_14285,N_13686,N_13624);
nor U14286 (N_14286,N_12096,N_12444);
nand U14287 (N_14287,N_12919,N_13701);
nand U14288 (N_14288,N_12901,N_13432);
nand U14289 (N_14289,N_13959,N_12152);
or U14290 (N_14290,N_13574,N_12538);
and U14291 (N_14291,N_12898,N_13142);
nand U14292 (N_14292,N_12932,N_13573);
or U14293 (N_14293,N_13214,N_12983);
and U14294 (N_14294,N_12557,N_12562);
nor U14295 (N_14295,N_13020,N_13845);
and U14296 (N_14296,N_12090,N_12935);
or U14297 (N_14297,N_12189,N_12693);
and U14298 (N_14298,N_12766,N_12478);
nor U14299 (N_14299,N_12493,N_13643);
nor U14300 (N_14300,N_13197,N_12238);
nor U14301 (N_14301,N_13612,N_13232);
nand U14302 (N_14302,N_12303,N_12423);
nor U14303 (N_14303,N_13454,N_12121);
nand U14304 (N_14304,N_13994,N_13409);
and U14305 (N_14305,N_12196,N_12545);
nor U14306 (N_14306,N_12381,N_13509);
nand U14307 (N_14307,N_12679,N_13909);
nand U14308 (N_14308,N_12920,N_13528);
nand U14309 (N_14309,N_13282,N_13429);
nor U14310 (N_14310,N_12992,N_12208);
and U14311 (N_14311,N_12892,N_13040);
nand U14312 (N_14312,N_13451,N_12409);
nand U14313 (N_14313,N_12791,N_13566);
nand U14314 (N_14314,N_12611,N_12187);
and U14315 (N_14315,N_12514,N_13858);
nor U14316 (N_14316,N_12641,N_13440);
nor U14317 (N_14317,N_12736,N_12391);
nor U14318 (N_14318,N_13893,N_12043);
and U14319 (N_14319,N_12627,N_13042);
or U14320 (N_14320,N_12383,N_13987);
nor U14321 (N_14321,N_12199,N_12229);
and U14322 (N_14322,N_13782,N_12139);
and U14323 (N_14323,N_12205,N_13850);
xnor U14324 (N_14324,N_13053,N_13706);
and U14325 (N_14325,N_13306,N_13410);
and U14326 (N_14326,N_12446,N_12582);
or U14327 (N_14327,N_12112,N_13560);
nor U14328 (N_14328,N_13659,N_12908);
nor U14329 (N_14329,N_13011,N_12120);
nor U14330 (N_14330,N_13699,N_13562);
nand U14331 (N_14331,N_13767,N_13769);
or U14332 (N_14332,N_12742,N_13249);
nand U14333 (N_14333,N_12400,N_12661);
or U14334 (N_14334,N_13952,N_12666);
nor U14335 (N_14335,N_13162,N_12059);
and U14336 (N_14336,N_13277,N_12500);
or U14337 (N_14337,N_12130,N_13698);
and U14338 (N_14338,N_13661,N_13133);
nor U14339 (N_14339,N_12148,N_13702);
or U14340 (N_14340,N_13433,N_13021);
nand U14341 (N_14341,N_12684,N_13851);
xnor U14342 (N_14342,N_13377,N_13051);
nor U14343 (N_14343,N_12865,N_12633);
and U14344 (N_14344,N_12945,N_13741);
nand U14345 (N_14345,N_13403,N_13024);
nor U14346 (N_14346,N_12930,N_12948);
or U14347 (N_14347,N_12198,N_13423);
xor U14348 (N_14348,N_13775,N_13398);
xnor U14349 (N_14349,N_13394,N_12620);
and U14350 (N_14350,N_13484,N_12006);
nor U14351 (N_14351,N_13174,N_13224);
xnor U14352 (N_14352,N_13977,N_13126);
and U14353 (N_14353,N_13937,N_12989);
nand U14354 (N_14354,N_12927,N_13406);
or U14355 (N_14355,N_12843,N_12572);
and U14356 (N_14356,N_13954,N_12014);
or U14357 (N_14357,N_13387,N_13870);
nor U14358 (N_14358,N_13919,N_12818);
or U14359 (N_14359,N_12610,N_13762);
or U14360 (N_14360,N_12925,N_12268);
xor U14361 (N_14361,N_12846,N_12646);
or U14362 (N_14362,N_12021,N_13459);
nor U14363 (N_14363,N_12715,N_12387);
nor U14364 (N_14364,N_12682,N_12328);
and U14365 (N_14365,N_13163,N_13319);
or U14366 (N_14366,N_13008,N_13951);
and U14367 (N_14367,N_13314,N_13313);
or U14368 (N_14368,N_13302,N_13949);
nand U14369 (N_14369,N_13926,N_12171);
and U14370 (N_14370,N_13520,N_13640);
and U14371 (N_14371,N_13446,N_12732);
or U14372 (N_14372,N_13176,N_13288);
nor U14373 (N_14373,N_13882,N_12885);
nand U14374 (N_14374,N_13291,N_12836);
nor U14375 (N_14375,N_12470,N_13747);
nand U14376 (N_14376,N_13931,N_12471);
or U14377 (N_14377,N_13839,N_13719);
or U14378 (N_14378,N_13450,N_12263);
nand U14379 (N_14379,N_12294,N_12921);
nand U14380 (N_14380,N_12585,N_12906);
and U14381 (N_14381,N_12499,N_13751);
or U14382 (N_14382,N_13363,N_12751);
xor U14383 (N_14383,N_12344,N_12762);
or U14384 (N_14384,N_13853,N_12694);
nor U14385 (N_14385,N_12757,N_12928);
nand U14386 (N_14386,N_12425,N_12250);
and U14387 (N_14387,N_12691,N_13027);
and U14388 (N_14388,N_12712,N_13441);
nand U14389 (N_14389,N_12631,N_12489);
nand U14390 (N_14390,N_12045,N_13274);
or U14391 (N_14391,N_12497,N_12576);
or U14392 (N_14392,N_13324,N_13792);
nor U14393 (N_14393,N_12568,N_13567);
xor U14394 (N_14394,N_13157,N_13402);
or U14395 (N_14395,N_12291,N_12170);
or U14396 (N_14396,N_12909,N_12259);
nand U14397 (N_14397,N_13515,N_12186);
nand U14398 (N_14398,N_13258,N_12554);
or U14399 (N_14399,N_12434,N_13061);
and U14400 (N_14400,N_12918,N_12428);
xor U14401 (N_14401,N_13689,N_12486);
or U14402 (N_14402,N_12750,N_12255);
xnor U14403 (N_14403,N_13555,N_13206);
and U14404 (N_14404,N_13399,N_12237);
nand U14405 (N_14405,N_12032,N_13602);
or U14406 (N_14406,N_12042,N_13285);
and U14407 (N_14407,N_13149,N_13397);
or U14408 (N_14408,N_13414,N_13503);
and U14409 (N_14409,N_13999,N_13144);
nor U14410 (N_14410,N_13830,N_12954);
and U14411 (N_14411,N_12355,N_13936);
nand U14412 (N_14412,N_12803,N_12265);
nor U14413 (N_14413,N_13140,N_13529);
or U14414 (N_14414,N_12855,N_12135);
or U14415 (N_14415,N_13283,N_13693);
or U14416 (N_14416,N_13930,N_12639);
or U14417 (N_14417,N_12143,N_12037);
and U14418 (N_14418,N_13067,N_13943);
nor U14419 (N_14419,N_13322,N_12377);
nor U14420 (N_14420,N_12302,N_12062);
or U14421 (N_14421,N_13017,N_13524);
nand U14422 (N_14422,N_13950,N_12804);
nor U14423 (N_14423,N_13664,N_12329);
or U14424 (N_14424,N_12929,N_12055);
xnor U14425 (N_14425,N_13407,N_12507);
and U14426 (N_14426,N_13871,N_12097);
and U14427 (N_14427,N_13756,N_12300);
nand U14428 (N_14428,N_12869,N_13370);
or U14429 (N_14429,N_13770,N_12356);
nor U14430 (N_14430,N_13252,N_12001);
nand U14431 (N_14431,N_12673,N_13261);
nor U14432 (N_14432,N_12706,N_12454);
nor U14433 (N_14433,N_12231,N_13022);
nand U14434 (N_14434,N_13041,N_12220);
and U14435 (N_14435,N_13878,N_12549);
or U14436 (N_14436,N_12213,N_13921);
or U14437 (N_14437,N_13963,N_13141);
and U14438 (N_14438,N_13903,N_12542);
nor U14439 (N_14439,N_13034,N_12458);
or U14440 (N_14440,N_13102,N_13129);
nand U14441 (N_14441,N_12319,N_13724);
nand U14442 (N_14442,N_13691,N_13259);
and U14443 (N_14443,N_13257,N_12982);
and U14444 (N_14444,N_12331,N_12984);
or U14445 (N_14445,N_12569,N_12811);
and U14446 (N_14446,N_13715,N_12241);
or U14447 (N_14447,N_12871,N_13376);
nor U14448 (N_14448,N_12827,N_12267);
or U14449 (N_14449,N_12488,N_12974);
nand U14450 (N_14450,N_12635,N_12720);
and U14451 (N_14451,N_12313,N_12537);
nand U14452 (N_14452,N_13411,N_13089);
nand U14453 (N_14453,N_12484,N_13988);
nor U14454 (N_14454,N_12789,N_13964);
nand U14455 (N_14455,N_12420,N_13110);
and U14456 (N_14456,N_13480,N_12065);
nand U14457 (N_14457,N_12971,N_13123);
nor U14458 (N_14458,N_12011,N_13828);
xor U14459 (N_14459,N_13914,N_13838);
nor U14460 (N_14460,N_13606,N_13507);
xor U14461 (N_14461,N_13883,N_12943);
nand U14462 (N_14462,N_13578,N_12102);
and U14463 (N_14463,N_13331,N_13902);
nand U14464 (N_14464,N_13361,N_12645);
nand U14465 (N_14465,N_13682,N_13009);
or U14466 (N_14466,N_12216,N_13247);
nor U14467 (N_14467,N_13974,N_13899);
nand U14468 (N_14468,N_13485,N_12575);
nand U14469 (N_14469,N_12524,N_13840);
nor U14470 (N_14470,N_13704,N_13490);
and U14471 (N_14471,N_12234,N_12002);
or U14472 (N_14472,N_13543,N_12138);
xnor U14473 (N_14473,N_12031,N_12539);
nand U14474 (N_14474,N_12799,N_12900);
and U14475 (N_14475,N_13367,N_12713);
or U14476 (N_14476,N_12248,N_12005);
nor U14477 (N_14477,N_12710,N_13976);
nor U14478 (N_14478,N_13362,N_12509);
xnor U14479 (N_14479,N_13267,N_12793);
nor U14480 (N_14480,N_12975,N_13164);
and U14481 (N_14481,N_12453,N_13345);
and U14482 (N_14482,N_13564,N_12607);
nand U14483 (N_14483,N_12450,N_13834);
nand U14484 (N_14484,N_13264,N_13855);
and U14485 (N_14485,N_12777,N_13248);
nor U14486 (N_14486,N_13551,N_13552);
nand U14487 (N_14487,N_12986,N_12089);
and U14488 (N_14488,N_12612,N_12695);
xnor U14489 (N_14489,N_12958,N_12339);
nor U14490 (N_14490,N_13347,N_12264);
nor U14491 (N_14491,N_12680,N_12912);
or U14492 (N_14492,N_12656,N_13981);
nand U14493 (N_14493,N_13969,N_13063);
or U14494 (N_14494,N_12277,N_13675);
nand U14495 (N_14495,N_13242,N_13737);
nor U14496 (N_14496,N_13486,N_13424);
and U14497 (N_14497,N_13904,N_12637);
xnor U14498 (N_14498,N_12163,N_13716);
xor U14499 (N_14499,N_12226,N_13677);
nor U14500 (N_14500,N_13841,N_12523);
and U14501 (N_14501,N_12598,N_13900);
xor U14502 (N_14502,N_12162,N_12099);
nand U14503 (N_14503,N_12654,N_13986);
nor U14504 (N_14504,N_13239,N_12413);
and U14505 (N_14505,N_13498,N_13568);
and U14506 (N_14506,N_13128,N_12159);
nand U14507 (N_14507,N_12049,N_12506);
nor U14508 (N_14508,N_13908,N_13487);
xor U14509 (N_14509,N_12917,N_12100);
and U14510 (N_14510,N_13638,N_13070);
or U14511 (N_14511,N_13615,N_13879);
and U14512 (N_14512,N_13340,N_13079);
and U14513 (N_14513,N_13712,N_12979);
nand U14514 (N_14514,N_12312,N_12448);
and U14515 (N_14515,N_12643,N_12340);
xor U14516 (N_14516,N_13208,N_12996);
xnor U14517 (N_14517,N_13685,N_12083);
and U14518 (N_14518,N_12606,N_13797);
nand U14519 (N_14519,N_13835,N_12533);
or U14520 (N_14520,N_13112,N_12937);
nor U14521 (N_14521,N_13294,N_12108);
xnor U14522 (N_14522,N_13570,N_12840);
nor U14523 (N_14523,N_13262,N_12886);
nor U14524 (N_14524,N_13642,N_12857);
and U14525 (N_14525,N_13846,N_12622);
nor U14526 (N_14526,N_12481,N_13464);
nand U14527 (N_14527,N_12086,N_13894);
or U14528 (N_14528,N_13103,N_12786);
nor U14529 (N_14529,N_12370,N_13323);
or U14530 (N_14530,N_12822,N_13438);
nand U14531 (N_14531,N_13238,N_13230);
nor U14532 (N_14532,N_12352,N_12028);
or U14533 (N_14533,N_12956,N_13418);
and U14534 (N_14534,N_13753,N_12151);
nand U14535 (N_14535,N_13874,N_12335);
nor U14536 (N_14536,N_13634,N_13062);
nor U14537 (N_14537,N_13920,N_13463);
nand U14538 (N_14538,N_13692,N_13098);
nor U14539 (N_14539,N_12296,N_13572);
nor U14540 (N_14540,N_12556,N_12649);
or U14541 (N_14541,N_13156,N_13618);
nand U14542 (N_14542,N_12949,N_12012);
nand U14543 (N_14543,N_13651,N_12795);
or U14544 (N_14544,N_12891,N_12498);
nand U14545 (N_14545,N_13456,N_13001);
nor U14546 (N_14546,N_13665,N_12546);
nand U14547 (N_14547,N_12106,N_12251);
nand U14548 (N_14548,N_12188,N_12000);
or U14549 (N_14549,N_12740,N_13392);
nor U14550 (N_14550,N_13372,N_13316);
or U14551 (N_14551,N_12046,N_12004);
nand U14552 (N_14552,N_12201,N_13823);
nor U14553 (N_14553,N_13813,N_12287);
nand U14554 (N_14554,N_13731,N_13557);
and U14555 (N_14555,N_12877,N_13668);
and U14556 (N_14556,N_12878,N_13650);
or U14557 (N_14557,N_13865,N_12570);
nand U14558 (N_14558,N_12357,N_12301);
or U14559 (N_14559,N_12950,N_13281);
nand U14560 (N_14560,N_13947,N_13925);
or U14561 (N_14561,N_12915,N_13084);
or U14562 (N_14562,N_13836,N_12601);
and U14563 (N_14563,N_12088,N_13945);
and U14564 (N_14564,N_12642,N_12310);
xor U14565 (N_14565,N_12870,N_13721);
xor U14566 (N_14566,N_13311,N_13733);
or U14567 (N_14567,N_12619,N_13540);
or U14568 (N_14568,N_13215,N_12479);
or U14569 (N_14569,N_12422,N_13518);
or U14570 (N_14570,N_12995,N_13906);
nand U14571 (N_14571,N_12574,N_13653);
and U14572 (N_14572,N_12648,N_13191);
nor U14573 (N_14573,N_13437,N_12475);
xnor U14574 (N_14574,N_13965,N_13505);
nor U14575 (N_14575,N_13944,N_12674);
nand U14576 (N_14576,N_12985,N_12764);
and U14577 (N_14577,N_12668,N_12193);
nand U14578 (N_14578,N_12672,N_12072);
or U14579 (N_14579,N_13493,N_12155);
nand U14580 (N_14580,N_12305,N_12734);
and U14581 (N_14581,N_13389,N_12839);
nor U14582 (N_14582,N_13260,N_13732);
and U14583 (N_14583,N_12275,N_13860);
or U14584 (N_14584,N_12775,N_13055);
nor U14585 (N_14585,N_12211,N_13293);
and U14586 (N_14586,N_13772,N_13033);
or U14587 (N_14587,N_13177,N_13473);
and U14588 (N_14588,N_13832,N_13471);
and U14589 (N_14589,N_12412,N_12690);
or U14590 (N_14590,N_12039,N_13843);
xnor U14591 (N_14591,N_12013,N_13296);
nand U14592 (N_14592,N_12874,N_13472);
nand U14593 (N_14593,N_12194,N_12082);
nand U14594 (N_14594,N_13227,N_13749);
and U14595 (N_14595,N_12580,N_12689);
and U14596 (N_14596,N_13344,N_12584);
or U14597 (N_14597,N_12204,N_13220);
or U14598 (N_14598,N_13085,N_13596);
nor U14599 (N_14599,N_12274,N_12092);
nand U14600 (N_14600,N_13873,N_13576);
nor U14601 (N_14601,N_13087,N_13057);
or U14602 (N_14602,N_12019,N_12426);
or U14603 (N_14603,N_12276,N_12038);
nor U14604 (N_14604,N_12999,N_12054);
and U14605 (N_14605,N_13821,N_12285);
or U14606 (N_14606,N_13297,N_12156);
xnor U14607 (N_14607,N_13382,N_13530);
and U14608 (N_14608,N_12859,N_13186);
nand U14609 (N_14609,N_13600,N_13400);
and U14610 (N_14610,N_12968,N_12600);
nand U14611 (N_14611,N_12185,N_13517);
xnor U14612 (N_14612,N_12754,N_13844);
or U14613 (N_14613,N_13117,N_12405);
and U14614 (N_14614,N_12070,N_13378);
and U14615 (N_14615,N_12398,N_13219);
or U14616 (N_14616,N_13026,N_12842);
nand U14617 (N_14617,N_12107,N_13083);
nor U14618 (N_14618,N_12105,N_12825);
and U14619 (N_14619,N_13785,N_13497);
and U14620 (N_14620,N_13955,N_12273);
nand U14621 (N_14621,N_13496,N_12883);
and U14622 (N_14622,N_12298,N_13787);
and U14623 (N_14623,N_12636,N_12091);
nor U14624 (N_14624,N_13666,N_13166);
nor U14625 (N_14625,N_12583,N_12535);
nand U14626 (N_14626,N_13179,N_13658);
nand U14627 (N_14627,N_12830,N_13153);
xor U14628 (N_14628,N_12941,N_12821);
and U14629 (N_14629,N_13550,N_12887);
nor U14630 (N_14630,N_12755,N_13773);
and U14631 (N_14631,N_12397,N_12501);
and U14632 (N_14632,N_12200,N_12057);
nand U14633 (N_14633,N_13143,N_13348);
nor U14634 (N_14634,N_13236,N_13805);
and U14635 (N_14635,N_13121,N_12299);
and U14636 (N_14636,N_13310,N_13985);
nand U14637 (N_14637,N_13605,N_13771);
nor U14638 (N_14638,N_13815,N_12526);
xor U14639 (N_14639,N_12852,N_12703);
nand U14640 (N_14640,N_12052,N_13337);
and U14641 (N_14641,N_13924,N_13091);
or U14642 (N_14642,N_13939,N_12931);
nor U14643 (N_14643,N_13199,N_13354);
and U14644 (N_14644,N_12727,N_12392);
or U14645 (N_14645,N_13875,N_12747);
or U14646 (N_14646,N_12801,N_12015);
nor U14647 (N_14647,N_12632,N_13868);
xnor U14648 (N_14648,N_12495,N_13373);
and U14649 (N_14649,N_12761,N_12980);
nand U14650 (N_14650,N_13723,N_13404);
nand U14651 (N_14651,N_13763,N_13190);
nor U14652 (N_14652,N_13353,N_13405);
nor U14653 (N_14653,N_12469,N_12236);
nand U14654 (N_14654,N_12297,N_12212);
nand U14655 (N_14655,N_12474,N_13396);
nor U14656 (N_14656,N_12023,N_13717);
or U14657 (N_14657,N_12316,N_12429);
nor U14658 (N_14658,N_13130,N_12829);
or U14659 (N_14659,N_12407,N_13015);
and U14660 (N_14660,N_12249,N_12368);
nand U14661 (N_14661,N_13469,N_12652);
nor U14662 (N_14662,N_12628,N_12354);
and U14663 (N_14663,N_13781,N_13478);
and U14664 (N_14664,N_12336,N_13803);
nand U14665 (N_14665,N_13745,N_13016);
nand U14666 (N_14666,N_13047,N_12117);
nand U14667 (N_14667,N_13533,N_13864);
or U14668 (N_14668,N_12376,N_13080);
or U14669 (N_14669,N_13972,N_12079);
or U14670 (N_14670,N_13700,N_12064);
or U14671 (N_14671,N_12864,N_12122);
nor U14672 (N_14672,N_13161,N_12348);
xnor U14673 (N_14673,N_13106,N_12116);
and U14674 (N_14674,N_12326,N_12176);
or U14675 (N_14675,N_13266,N_13758);
or U14676 (N_14676,N_13927,N_13122);
xor U14677 (N_14677,N_12944,N_13519);
or U14678 (N_14678,N_12373,N_13170);
nand U14679 (N_14679,N_13036,N_12884);
nor U14680 (N_14680,N_12759,N_12063);
or U14681 (N_14681,N_12991,N_12602);
or U14682 (N_14682,N_13048,N_13488);
and U14683 (N_14683,N_12615,N_13537);
nor U14684 (N_14684,N_12077,N_12763);
and U14685 (N_14685,N_13694,N_13856);
or U14686 (N_14686,N_13958,N_13054);
or U14687 (N_14687,N_12905,N_12965);
nor U14688 (N_14688,N_13427,N_12579);
and U14689 (N_14689,N_12050,N_12334);
xor U14690 (N_14690,N_12504,N_12402);
or U14691 (N_14691,N_13180,N_12182);
nand U14692 (N_14692,N_12940,N_12191);
and U14693 (N_14693,N_13359,N_13200);
or U14694 (N_14694,N_12812,N_13327);
and U14695 (N_14695,N_12735,N_13710);
and U14696 (N_14696,N_13736,N_12851);
xor U14697 (N_14697,N_12698,N_13134);
and U14698 (N_14698,N_13598,N_13804);
and U14699 (N_14699,N_12411,N_13971);
xor U14700 (N_14700,N_13617,N_12433);
nand U14701 (N_14701,N_12496,N_13005);
xor U14702 (N_14702,N_13506,N_12040);
nor U14703 (N_14703,N_13750,N_12401);
nand U14704 (N_14704,N_12068,N_12880);
nor U14705 (N_14705,N_13045,N_13746);
and U14706 (N_14706,N_13435,N_12209);
xnor U14707 (N_14707,N_13364,N_13077);
xnor U14708 (N_14708,N_12460,N_13279);
and U14709 (N_14709,N_13272,N_12227);
nand U14710 (N_14710,N_12765,N_13910);
nor U14711 (N_14711,N_12692,N_12315);
nor U14712 (N_14712,N_13237,N_12964);
or U14713 (N_14713,N_13209,N_12770);
or U14714 (N_14714,N_12823,N_12369);
and U14715 (N_14715,N_13579,N_12283);
nor U14716 (N_14716,N_13687,N_12963);
nor U14717 (N_14717,N_13801,N_12378);
or U14718 (N_14718,N_12593,N_13847);
or U14719 (N_14719,N_13688,N_13321);
or U14720 (N_14720,N_13204,N_13038);
or U14721 (N_14721,N_13012,N_13205);
nor U14722 (N_14722,N_13371,N_13680);
nand U14723 (N_14723,N_12826,N_12779);
or U14724 (N_14724,N_13032,N_13890);
nand U14725 (N_14725,N_12952,N_13810);
nor U14726 (N_14726,N_13243,N_13482);
nor U14727 (N_14727,N_13135,N_12716);
or U14728 (N_14728,N_13349,N_12421);
xor U14729 (N_14729,N_12756,N_13827);
nand U14730 (N_14730,N_13970,N_12174);
or U14731 (N_14731,N_12144,N_13817);
and U14732 (N_14732,N_13795,N_12882);
nor U14733 (N_14733,N_12010,N_12243);
and U14734 (N_14734,N_13695,N_13595);
nand U14735 (N_14735,N_12990,N_12753);
and U14736 (N_14736,N_12110,N_13368);
nand U14737 (N_14737,N_12629,N_12210);
or U14738 (N_14738,N_12560,N_12888);
or U14739 (N_14739,N_13554,N_12977);
and U14740 (N_14740,N_12733,N_12910);
and U14741 (N_14741,N_12123,N_13462);
xor U14742 (N_14742,N_12834,N_13938);
and U14743 (N_14743,N_12007,N_13738);
and U14744 (N_14744,N_12085,N_13068);
nand U14745 (N_14745,N_12103,N_12923);
nand U14746 (N_14746,N_13307,N_12158);
nand U14747 (N_14747,N_13284,N_13662);
nand U14748 (N_14748,N_12462,N_12717);
and U14749 (N_14749,N_12697,N_12306);
and U14750 (N_14750,N_13862,N_13492);
nor U14751 (N_14751,N_13608,N_13263);
or U14752 (N_14752,N_13443,N_12993);
xor U14753 (N_14753,N_12338,N_13684);
nor U14754 (N_14754,N_13541,N_12814);
nor U14755 (N_14755,N_13107,N_12147);
nand U14756 (N_14756,N_13168,N_12828);
nor U14757 (N_14757,N_12257,N_13412);
or U14758 (N_14758,N_12837,N_13824);
or U14759 (N_14759,N_13861,N_13194);
or U14760 (N_14760,N_12768,N_13124);
nand U14761 (N_14761,N_13268,N_13657);
nor U14762 (N_14762,N_13934,N_12111);
nor U14763 (N_14763,N_12217,N_12953);
nand U14764 (N_14764,N_13078,N_13593);
nor U14765 (N_14765,N_12879,N_13705);
and U14766 (N_14766,N_12741,N_13941);
nand U14767 (N_14767,N_12788,N_12150);
xnor U14768 (N_14768,N_13759,N_13413);
nor U14769 (N_14769,N_13095,N_13299);
and U14770 (N_14770,N_13502,N_12807);
or U14771 (N_14771,N_13929,N_13989);
nand U14772 (N_14772,N_13467,N_13535);
and U14773 (N_14773,N_12708,N_13100);
nor U14774 (N_14774,N_12058,N_12330);
nand U14775 (N_14775,N_12337,N_13633);
xnor U14776 (N_14776,N_13290,N_13820);
nand U14777 (N_14777,N_13779,N_13309);
or U14778 (N_14778,N_13169,N_13419);
nor U14779 (N_14779,N_12760,N_12311);
nor U14780 (N_14780,N_12653,N_12902);
nand U14781 (N_14781,N_13571,N_12820);
nand U14782 (N_14782,N_13052,N_13742);
and U14783 (N_14783,N_12705,N_12183);
and U14784 (N_14784,N_12347,N_12512);
nor U14785 (N_14785,N_13644,N_12655);
or U14786 (N_14786,N_13678,N_12519);
nand U14787 (N_14787,N_12709,N_12415);
and U14788 (N_14788,N_13697,N_12436);
nor U14789 (N_14789,N_12447,N_13059);
nor U14790 (N_14790,N_12810,N_13859);
or U14791 (N_14791,N_13948,N_12172);
xor U14792 (N_14792,N_13646,N_12746);
xor U14793 (N_14793,N_13581,N_13630);
and U14794 (N_14794,N_12529,N_12783);
and U14795 (N_14795,N_12233,N_12350);
or U14796 (N_14796,N_13246,N_12307);
nand U14797 (N_14797,N_12540,N_13778);
nor U14798 (N_14798,N_12245,N_12737);
or U14799 (N_14799,N_12367,N_12056);
or U14800 (N_14800,N_12018,N_12266);
nor U14801 (N_14801,N_12161,N_12808);
nor U14802 (N_14802,N_12875,N_13922);
nand U14803 (N_14803,N_13599,N_12895);
nand U14804 (N_14804,N_13559,N_12362);
xor U14805 (N_14805,N_13086,N_12437);
nor U14806 (N_14806,N_13477,N_13565);
nor U14807 (N_14807,N_13235,N_13585);
nand U14808 (N_14808,N_13425,N_12075);
nor U14809 (N_14809,N_13388,N_13158);
and U14810 (N_14810,N_12711,N_13119);
and U14811 (N_14811,N_13799,N_13663);
nor U14812 (N_14812,N_12515,N_12482);
nor U14813 (N_14813,N_13962,N_13923);
or U14814 (N_14814,N_13953,N_12558);
or U14815 (N_14815,N_13201,N_13928);
xor U14816 (N_14816,N_12520,N_12517);
or U14817 (N_14817,N_13101,N_12893);
and U14818 (N_14818,N_13636,N_13050);
nand U14819 (N_14819,N_13421,N_12414);
nor U14820 (N_14820,N_12573,N_12616);
and U14821 (N_14821,N_13726,N_12372);
nor U14822 (N_14822,N_13647,N_13730);
nand U14823 (N_14823,N_12449,N_12380);
xor U14824 (N_14824,N_12876,N_12153);
or U14825 (N_14825,N_12790,N_12476);
and U14826 (N_14826,N_13794,N_13229);
nand U14827 (N_14827,N_12907,N_13428);
or U14828 (N_14828,N_13341,N_13895);
or U14829 (N_14829,N_12511,N_12124);
nand U14830 (N_14830,N_13619,N_13892);
and U14831 (N_14831,N_12532,N_13058);
and U14832 (N_14832,N_13195,N_12787);
or U14833 (N_14833,N_13791,N_13877);
nand U14834 (N_14834,N_12223,N_12686);
nand U14835 (N_14835,N_13049,N_13203);
nor U14836 (N_14836,N_12528,N_13000);
nor U14837 (N_14837,N_12258,N_12563);
nand U14838 (N_14838,N_13228,N_13725);
or U14839 (N_14839,N_13444,N_12609);
xnor U14840 (N_14840,N_13544,N_13460);
or U14841 (N_14841,N_12395,N_12332);
xor U14842 (N_14842,N_13244,N_12976);
xor U14843 (N_14843,N_12084,N_12473);
nand U14844 (N_14844,N_13060,N_13886);
nor U14845 (N_14845,N_13315,N_12926);
xnor U14846 (N_14846,N_13391,N_12752);
xnor U14847 (N_14847,N_13876,N_12581);
nand U14848 (N_14848,N_12438,N_12856);
or U14849 (N_14849,N_12534,N_12406);
or U14850 (N_14850,N_12552,N_13132);
nor U14851 (N_14851,N_12873,N_13234);
nand U14852 (N_14852,N_12073,N_13872);
or U14853 (N_14853,N_12955,N_13603);
nor U14854 (N_14854,N_12966,N_13975);
nor U14855 (N_14855,N_12293,N_12154);
nor U14856 (N_14856,N_13973,N_12345);
and U14857 (N_14857,N_13495,N_13351);
nor U14858 (N_14858,N_13028,N_13880);
and U14859 (N_14859,N_12051,N_13108);
nand U14860 (N_14860,N_13708,N_12468);
and U14861 (N_14861,N_13761,N_13913);
or U14862 (N_14862,N_12030,N_12599);
nand U14863 (N_14863,N_12390,N_13525);
or U14864 (N_14864,N_13317,N_12960);
xnor U14865 (N_14865,N_13942,N_12384);
and U14866 (N_14866,N_13240,N_13328);
or U14867 (N_14867,N_13983,N_13111);
and U14868 (N_14868,N_12101,N_12894);
nand U14869 (N_14869,N_12605,N_12327);
and U14870 (N_14870,N_12230,N_13379);
or U14871 (N_14871,N_13553,N_13601);
and U14872 (N_14872,N_12961,N_12224);
and U14873 (N_14873,N_12503,N_12784);
or U14874 (N_14874,N_12119,N_12195);
nor U14875 (N_14875,N_13338,N_13807);
and U14876 (N_14876,N_12933,N_13025);
nor U14877 (N_14877,N_13401,N_12725);
nor U14878 (N_14878,N_12721,N_12881);
and U14879 (N_14879,N_12071,N_12177);
and U14880 (N_14880,N_13326,N_13907);
and U14881 (N_14881,N_13622,N_13265);
xnor U14882 (N_14882,N_12131,N_13854);
and U14883 (N_14883,N_13734,N_12286);
and U14884 (N_14884,N_12104,N_12853);
and U14885 (N_14885,N_13241,N_13917);
nand U14886 (N_14886,N_12916,N_13829);
nor U14887 (N_14887,N_12281,N_13547);
nor U14888 (N_14888,N_13275,N_12033);
nor U14889 (N_14889,N_12394,N_13225);
nor U14890 (N_14890,N_12604,N_13014);
nor U14891 (N_14891,N_13614,N_12806);
nor U14892 (N_14892,N_12624,N_12441);
or U14893 (N_14893,N_12003,N_12292);
or U14894 (N_14894,N_13030,N_13714);
nor U14895 (N_14895,N_12849,N_13010);
nand U14896 (N_14896,N_13915,N_12491);
or U14897 (N_14897,N_13979,N_13852);
nor U14898 (N_14898,N_13654,N_12280);
xor U14899 (N_14899,N_12767,N_13798);
or U14900 (N_14900,N_13911,N_12371);
nand U14901 (N_14901,N_13417,N_13318);
xnor U14902 (N_14902,N_13350,N_12824);
or U14903 (N_14903,N_13152,N_12675);
nand U14904 (N_14904,N_13672,N_13202);
or U14905 (N_14905,N_13594,N_12034);
nand U14906 (N_14906,N_12080,N_12270);
nand U14907 (N_14907,N_13476,N_13765);
or U14908 (N_14908,N_13897,N_13468);
xor U14909 (N_14909,N_12972,N_12455);
or U14910 (N_14910,N_12133,N_12862);
nand U14911 (N_14911,N_12731,N_12704);
and U14912 (N_14912,N_13869,N_12590);
nand U14913 (N_14913,N_13623,N_13652);
or U14914 (N_14914,N_13018,N_12360);
nand U14915 (N_14915,N_12719,N_13580);
and U14916 (N_14916,N_12771,N_12613);
and U14917 (N_14917,N_12969,N_12008);
and U14918 (N_14918,N_12845,N_13250);
nand U14919 (N_14919,N_12817,N_13669);
nand U14920 (N_14920,N_13957,N_13114);
nor U14921 (N_14921,N_13866,N_12998);
or U14922 (N_14922,N_13393,N_13980);
nand U14923 (N_14923,N_12567,N_12221);
and U14924 (N_14924,N_12897,N_12564);
nor U14925 (N_14925,N_13786,N_13222);
or U14926 (N_14926,N_12530,N_12813);
and U14927 (N_14927,N_12625,N_13470);
or U14928 (N_14928,N_13722,N_13777);
or U14929 (N_14929,N_12951,N_13819);
and U14930 (N_14930,N_12651,N_13301);
nand U14931 (N_14931,N_13154,N_12081);
xnor U14932 (N_14932,N_12440,N_13956);
or U14933 (N_14933,N_13788,N_12044);
nor U14934 (N_14934,N_13216,N_13182);
or U14935 (N_14935,N_12970,N_12066);
nand U14936 (N_14936,N_12256,N_12778);
nand U14937 (N_14937,N_13189,N_12290);
or U14938 (N_14938,N_12702,N_13175);
xnor U14939 (N_14939,N_12774,N_13031);
nor U14940 (N_14940,N_13365,N_12109);
xnor U14941 (N_14941,N_12565,N_12318);
nand U14942 (N_14942,N_13992,N_12544);
nand U14943 (N_14943,N_13504,N_13312);
or U14944 (N_14944,N_13671,N_13639);
or U14945 (N_14945,N_12978,N_13621);
nor U14946 (N_14946,N_12973,N_13088);
nor U14947 (N_14947,N_12748,N_12396);
xnor U14948 (N_14948,N_12314,N_13384);
nand U14949 (N_14949,N_12492,N_13380);
nand U14950 (N_14950,N_13676,N_13366);
nand U14951 (N_14951,N_13155,N_12333);
and U14952 (N_14952,N_12320,N_12179);
nor U14953 (N_14953,N_13912,N_12141);
xnor U14954 (N_14954,N_12272,N_13304);
and U14955 (N_14955,N_12617,N_12215);
nand U14956 (N_14956,N_13218,N_12219);
and U14957 (N_14957,N_12681,N_12114);
and U14958 (N_14958,N_12547,N_12047);
nor U14959 (N_14959,N_12914,N_13198);
or U14960 (N_14960,N_13420,N_13548);
nand U14961 (N_14961,N_13727,N_13822);
nand U14962 (N_14962,N_13029,N_13542);
nand U14963 (N_14963,N_13431,N_12525);
xor U14964 (N_14964,N_13346,N_13489);
and U14965 (N_14965,N_12638,N_13513);
xor U14966 (N_14966,N_13993,N_13188);
nor U14967 (N_14967,N_13455,N_12029);
or U14968 (N_14968,N_13037,N_13329);
nor U14969 (N_14969,N_12832,N_12260);
and U14970 (N_14970,N_13113,N_13918);
nand U14971 (N_14971,N_12203,N_13735);
and U14972 (N_14972,N_12701,N_13295);
nand U14973 (N_14973,N_12594,N_13641);
or U14974 (N_14974,N_13093,N_12343);
and U14975 (N_14975,N_12341,N_13995);
xor U14976 (N_14976,N_12026,N_12872);
nor U14977 (N_14977,N_13757,N_12410);
or U14978 (N_14978,N_12772,N_12247);
nor U14979 (N_14979,N_13374,N_12242);
or U14980 (N_14980,N_12889,N_12687);
nand U14981 (N_14981,N_13138,N_12009);
nand U14982 (N_14982,N_12800,N_13826);
or U14983 (N_14983,N_12936,N_12240);
and U14984 (N_14984,N_13356,N_12269);
and U14985 (N_14985,N_12957,N_12351);
nand U14986 (N_14986,N_12261,N_13120);
nand U14987 (N_14987,N_13901,N_12844);
nand U14988 (N_14988,N_13627,N_13534);
nand U14989 (N_14989,N_12323,N_13226);
xor U14990 (N_14990,N_13342,N_13848);
or U14991 (N_14991,N_13538,N_12132);
nor U14992 (N_14992,N_12502,N_12218);
nor U14993 (N_14993,N_13933,N_12833);
nand U14994 (N_14994,N_12076,N_12451);
or U14995 (N_14995,N_12794,N_13760);
nor U14996 (N_14996,N_13690,N_12997);
and U14997 (N_14997,N_12432,N_12588);
and U14998 (N_14998,N_12435,N_12531);
nand U14999 (N_14999,N_12946,N_13173);
nor U15000 (N_15000,N_13972,N_13674);
nand U15001 (N_15001,N_12656,N_13727);
or U15002 (N_15002,N_12463,N_12495);
nand U15003 (N_15003,N_12047,N_12165);
nor U15004 (N_15004,N_13008,N_12115);
xnor U15005 (N_15005,N_12773,N_12741);
nor U15006 (N_15006,N_13008,N_13707);
xor U15007 (N_15007,N_12270,N_12399);
and U15008 (N_15008,N_13709,N_13392);
and U15009 (N_15009,N_13473,N_12738);
nand U15010 (N_15010,N_12905,N_12080);
or U15011 (N_15011,N_12709,N_12520);
or U15012 (N_15012,N_13704,N_12806);
nor U15013 (N_15013,N_13062,N_13834);
or U15014 (N_15014,N_13162,N_13673);
or U15015 (N_15015,N_12719,N_12103);
nand U15016 (N_15016,N_13734,N_13878);
xnor U15017 (N_15017,N_13262,N_13766);
nor U15018 (N_15018,N_12782,N_12331);
nand U15019 (N_15019,N_13392,N_13922);
or U15020 (N_15020,N_12147,N_12974);
and U15021 (N_15021,N_13344,N_12481);
xnor U15022 (N_15022,N_12790,N_13621);
nand U15023 (N_15023,N_12254,N_13810);
nand U15024 (N_15024,N_13733,N_12073);
xnor U15025 (N_15025,N_12456,N_12529);
and U15026 (N_15026,N_12499,N_12203);
or U15027 (N_15027,N_13492,N_12406);
nand U15028 (N_15028,N_13219,N_12952);
and U15029 (N_15029,N_13181,N_12295);
and U15030 (N_15030,N_13240,N_12468);
nor U15031 (N_15031,N_12548,N_13852);
nor U15032 (N_15032,N_13941,N_13449);
nor U15033 (N_15033,N_12446,N_12036);
or U15034 (N_15034,N_12105,N_13944);
or U15035 (N_15035,N_13756,N_12281);
or U15036 (N_15036,N_12651,N_13825);
and U15037 (N_15037,N_12680,N_12399);
and U15038 (N_15038,N_13319,N_12845);
nor U15039 (N_15039,N_12724,N_12069);
nand U15040 (N_15040,N_13732,N_12294);
xor U15041 (N_15041,N_12073,N_12671);
and U15042 (N_15042,N_13135,N_12706);
nand U15043 (N_15043,N_12726,N_12079);
nand U15044 (N_15044,N_12782,N_12406);
and U15045 (N_15045,N_13701,N_12231);
and U15046 (N_15046,N_12706,N_12402);
nand U15047 (N_15047,N_13228,N_12236);
and U15048 (N_15048,N_12975,N_13830);
nor U15049 (N_15049,N_13882,N_13879);
and U15050 (N_15050,N_12298,N_12311);
or U15051 (N_15051,N_13493,N_12396);
nand U15052 (N_15052,N_12892,N_13027);
and U15053 (N_15053,N_13945,N_12622);
or U15054 (N_15054,N_12663,N_13921);
or U15055 (N_15055,N_12605,N_12716);
nor U15056 (N_15056,N_13817,N_13666);
and U15057 (N_15057,N_13933,N_12617);
xor U15058 (N_15058,N_13473,N_12577);
xnor U15059 (N_15059,N_13405,N_12899);
nand U15060 (N_15060,N_12195,N_12042);
and U15061 (N_15061,N_13945,N_13698);
or U15062 (N_15062,N_12544,N_12730);
and U15063 (N_15063,N_12572,N_13046);
nand U15064 (N_15064,N_12486,N_13217);
nor U15065 (N_15065,N_13407,N_13615);
or U15066 (N_15066,N_13707,N_13674);
and U15067 (N_15067,N_12903,N_12113);
nor U15068 (N_15068,N_13583,N_13595);
and U15069 (N_15069,N_12916,N_13068);
and U15070 (N_15070,N_13510,N_12991);
and U15071 (N_15071,N_13291,N_12378);
nand U15072 (N_15072,N_13106,N_12235);
xor U15073 (N_15073,N_13638,N_13628);
and U15074 (N_15074,N_12986,N_13899);
nor U15075 (N_15075,N_12364,N_12316);
nor U15076 (N_15076,N_13795,N_12629);
and U15077 (N_15077,N_13329,N_13944);
or U15078 (N_15078,N_12799,N_13537);
nand U15079 (N_15079,N_13222,N_12425);
or U15080 (N_15080,N_13172,N_12713);
nor U15081 (N_15081,N_13193,N_12734);
xnor U15082 (N_15082,N_12187,N_13882);
and U15083 (N_15083,N_13322,N_12248);
and U15084 (N_15084,N_12895,N_12523);
nand U15085 (N_15085,N_12058,N_13769);
or U15086 (N_15086,N_12205,N_12394);
or U15087 (N_15087,N_13332,N_12892);
nor U15088 (N_15088,N_12553,N_12710);
and U15089 (N_15089,N_12312,N_12718);
nand U15090 (N_15090,N_13608,N_12762);
xnor U15091 (N_15091,N_13034,N_13210);
nand U15092 (N_15092,N_12021,N_12912);
or U15093 (N_15093,N_13553,N_12495);
nand U15094 (N_15094,N_12821,N_13993);
nand U15095 (N_15095,N_13065,N_13717);
nand U15096 (N_15096,N_12749,N_12471);
xnor U15097 (N_15097,N_13567,N_12024);
and U15098 (N_15098,N_13699,N_12252);
nand U15099 (N_15099,N_12541,N_13701);
and U15100 (N_15100,N_13166,N_12745);
or U15101 (N_15101,N_12699,N_13967);
nor U15102 (N_15102,N_12345,N_12179);
or U15103 (N_15103,N_12483,N_13946);
and U15104 (N_15104,N_13994,N_13299);
nand U15105 (N_15105,N_13118,N_12422);
or U15106 (N_15106,N_13049,N_12848);
nand U15107 (N_15107,N_12539,N_13171);
xor U15108 (N_15108,N_12956,N_13936);
and U15109 (N_15109,N_12098,N_13534);
nand U15110 (N_15110,N_12331,N_12029);
nand U15111 (N_15111,N_12435,N_12161);
and U15112 (N_15112,N_12400,N_13861);
or U15113 (N_15113,N_12992,N_12617);
or U15114 (N_15114,N_13999,N_12783);
nor U15115 (N_15115,N_13888,N_12225);
nor U15116 (N_15116,N_12955,N_12048);
nand U15117 (N_15117,N_13218,N_12689);
nor U15118 (N_15118,N_13282,N_12332);
and U15119 (N_15119,N_13399,N_13350);
xnor U15120 (N_15120,N_13162,N_13713);
or U15121 (N_15121,N_12030,N_13345);
xnor U15122 (N_15122,N_12459,N_12530);
nand U15123 (N_15123,N_12099,N_13715);
nand U15124 (N_15124,N_12942,N_13896);
and U15125 (N_15125,N_12574,N_12059);
or U15126 (N_15126,N_12523,N_13006);
or U15127 (N_15127,N_12578,N_13573);
nand U15128 (N_15128,N_12579,N_13834);
and U15129 (N_15129,N_12124,N_12969);
or U15130 (N_15130,N_12025,N_13084);
nand U15131 (N_15131,N_12065,N_13986);
or U15132 (N_15132,N_13696,N_13289);
or U15133 (N_15133,N_13423,N_13283);
nor U15134 (N_15134,N_13863,N_12155);
nand U15135 (N_15135,N_13366,N_12490);
nor U15136 (N_15136,N_13722,N_12820);
or U15137 (N_15137,N_13967,N_13855);
and U15138 (N_15138,N_12442,N_13436);
nor U15139 (N_15139,N_13658,N_12649);
and U15140 (N_15140,N_13288,N_12455);
nor U15141 (N_15141,N_12449,N_12024);
nand U15142 (N_15142,N_12265,N_13861);
and U15143 (N_15143,N_13565,N_13571);
and U15144 (N_15144,N_12696,N_13232);
or U15145 (N_15145,N_12563,N_12562);
or U15146 (N_15146,N_13308,N_13457);
and U15147 (N_15147,N_13048,N_13492);
nor U15148 (N_15148,N_13259,N_12431);
or U15149 (N_15149,N_12321,N_12088);
and U15150 (N_15150,N_13214,N_13533);
or U15151 (N_15151,N_12281,N_12900);
nor U15152 (N_15152,N_13324,N_12730);
or U15153 (N_15153,N_12918,N_12326);
and U15154 (N_15154,N_12306,N_13086);
nand U15155 (N_15155,N_12811,N_12211);
or U15156 (N_15156,N_12593,N_13254);
or U15157 (N_15157,N_13469,N_13231);
nand U15158 (N_15158,N_13564,N_12804);
nand U15159 (N_15159,N_13786,N_12981);
or U15160 (N_15160,N_13512,N_12835);
or U15161 (N_15161,N_12349,N_12622);
nand U15162 (N_15162,N_12629,N_13051);
nand U15163 (N_15163,N_13525,N_13813);
and U15164 (N_15164,N_13861,N_12968);
and U15165 (N_15165,N_13582,N_12788);
and U15166 (N_15166,N_13924,N_13885);
or U15167 (N_15167,N_13711,N_12896);
nand U15168 (N_15168,N_13863,N_12085);
nand U15169 (N_15169,N_12271,N_12582);
nand U15170 (N_15170,N_13668,N_13788);
and U15171 (N_15171,N_13361,N_12124);
nand U15172 (N_15172,N_12485,N_13163);
nor U15173 (N_15173,N_12296,N_13603);
or U15174 (N_15174,N_12620,N_13950);
and U15175 (N_15175,N_12488,N_12496);
xnor U15176 (N_15176,N_12219,N_12063);
and U15177 (N_15177,N_12796,N_12482);
xnor U15178 (N_15178,N_12882,N_13104);
or U15179 (N_15179,N_13761,N_13511);
nand U15180 (N_15180,N_13226,N_12341);
nand U15181 (N_15181,N_13580,N_13473);
nor U15182 (N_15182,N_13688,N_13257);
or U15183 (N_15183,N_12059,N_12877);
nand U15184 (N_15184,N_13966,N_12223);
and U15185 (N_15185,N_12472,N_13098);
and U15186 (N_15186,N_12256,N_13088);
or U15187 (N_15187,N_12590,N_12500);
nand U15188 (N_15188,N_13805,N_13846);
or U15189 (N_15189,N_13383,N_13774);
and U15190 (N_15190,N_12315,N_12316);
nor U15191 (N_15191,N_12423,N_13409);
or U15192 (N_15192,N_13588,N_13662);
nor U15193 (N_15193,N_13569,N_13765);
or U15194 (N_15194,N_13090,N_12037);
and U15195 (N_15195,N_13078,N_12447);
xnor U15196 (N_15196,N_12349,N_12281);
and U15197 (N_15197,N_13362,N_13125);
nand U15198 (N_15198,N_13311,N_12850);
nand U15199 (N_15199,N_12832,N_13861);
nand U15200 (N_15200,N_13378,N_13215);
or U15201 (N_15201,N_13103,N_12105);
nor U15202 (N_15202,N_12419,N_12111);
nand U15203 (N_15203,N_13155,N_13265);
nand U15204 (N_15204,N_12600,N_12051);
and U15205 (N_15205,N_13621,N_13734);
nand U15206 (N_15206,N_12833,N_12176);
nand U15207 (N_15207,N_13179,N_12760);
and U15208 (N_15208,N_13182,N_12448);
nor U15209 (N_15209,N_13705,N_12728);
nor U15210 (N_15210,N_12787,N_12373);
xnor U15211 (N_15211,N_12670,N_13710);
nor U15212 (N_15212,N_12711,N_12440);
nand U15213 (N_15213,N_12053,N_13429);
or U15214 (N_15214,N_13468,N_12192);
xnor U15215 (N_15215,N_13369,N_12433);
and U15216 (N_15216,N_12418,N_12575);
and U15217 (N_15217,N_12372,N_13140);
nor U15218 (N_15218,N_13896,N_12843);
or U15219 (N_15219,N_13555,N_13630);
nor U15220 (N_15220,N_13477,N_12289);
and U15221 (N_15221,N_12859,N_12235);
nor U15222 (N_15222,N_12688,N_12058);
nor U15223 (N_15223,N_13981,N_12832);
or U15224 (N_15224,N_13445,N_13709);
nor U15225 (N_15225,N_13268,N_13210);
nand U15226 (N_15226,N_12972,N_12421);
or U15227 (N_15227,N_13091,N_12106);
nor U15228 (N_15228,N_13202,N_12290);
and U15229 (N_15229,N_13682,N_12621);
and U15230 (N_15230,N_13954,N_12684);
or U15231 (N_15231,N_13463,N_12514);
nor U15232 (N_15232,N_13559,N_13343);
and U15233 (N_15233,N_13049,N_13453);
and U15234 (N_15234,N_12115,N_13771);
nand U15235 (N_15235,N_12188,N_12989);
and U15236 (N_15236,N_13013,N_13863);
or U15237 (N_15237,N_13006,N_12947);
and U15238 (N_15238,N_13325,N_13340);
nand U15239 (N_15239,N_12352,N_13051);
or U15240 (N_15240,N_12540,N_12496);
and U15241 (N_15241,N_12083,N_12064);
nand U15242 (N_15242,N_12152,N_13237);
nor U15243 (N_15243,N_13416,N_12333);
or U15244 (N_15244,N_12866,N_13097);
nand U15245 (N_15245,N_12088,N_12853);
nand U15246 (N_15246,N_13457,N_13437);
or U15247 (N_15247,N_13979,N_13607);
nor U15248 (N_15248,N_12844,N_13227);
xor U15249 (N_15249,N_12482,N_12038);
or U15250 (N_15250,N_12210,N_13550);
nand U15251 (N_15251,N_13921,N_13609);
xor U15252 (N_15252,N_12963,N_12025);
nand U15253 (N_15253,N_13091,N_13363);
nand U15254 (N_15254,N_13135,N_12822);
and U15255 (N_15255,N_12647,N_12545);
and U15256 (N_15256,N_12060,N_13058);
nor U15257 (N_15257,N_12686,N_13095);
xor U15258 (N_15258,N_13351,N_13952);
and U15259 (N_15259,N_12280,N_12800);
xor U15260 (N_15260,N_12586,N_13417);
nand U15261 (N_15261,N_13123,N_13943);
nor U15262 (N_15262,N_12441,N_13798);
or U15263 (N_15263,N_12651,N_13692);
and U15264 (N_15264,N_13575,N_13319);
and U15265 (N_15265,N_12168,N_13743);
or U15266 (N_15266,N_13022,N_13098);
nand U15267 (N_15267,N_12372,N_12971);
nand U15268 (N_15268,N_13832,N_12851);
nor U15269 (N_15269,N_13444,N_13902);
or U15270 (N_15270,N_12646,N_13231);
and U15271 (N_15271,N_12319,N_13230);
and U15272 (N_15272,N_12978,N_12070);
nor U15273 (N_15273,N_13808,N_13282);
nor U15274 (N_15274,N_13707,N_12104);
and U15275 (N_15275,N_13984,N_13349);
or U15276 (N_15276,N_12302,N_12506);
nand U15277 (N_15277,N_13214,N_12254);
nor U15278 (N_15278,N_13380,N_12915);
and U15279 (N_15279,N_12832,N_12719);
nor U15280 (N_15280,N_13025,N_12374);
xor U15281 (N_15281,N_12608,N_12302);
and U15282 (N_15282,N_12206,N_12223);
or U15283 (N_15283,N_13840,N_12622);
or U15284 (N_15284,N_13899,N_13107);
xor U15285 (N_15285,N_13231,N_12776);
nand U15286 (N_15286,N_13680,N_13689);
and U15287 (N_15287,N_13464,N_13434);
and U15288 (N_15288,N_12172,N_12060);
and U15289 (N_15289,N_12901,N_12080);
xor U15290 (N_15290,N_13912,N_13504);
or U15291 (N_15291,N_13461,N_12712);
nor U15292 (N_15292,N_13953,N_13163);
nor U15293 (N_15293,N_12955,N_13641);
xor U15294 (N_15294,N_13885,N_12046);
and U15295 (N_15295,N_13121,N_12885);
nor U15296 (N_15296,N_13340,N_13135);
nor U15297 (N_15297,N_12895,N_13893);
or U15298 (N_15298,N_13137,N_13880);
or U15299 (N_15299,N_13989,N_12572);
or U15300 (N_15300,N_13962,N_13448);
nand U15301 (N_15301,N_13482,N_13065);
and U15302 (N_15302,N_13903,N_13182);
nand U15303 (N_15303,N_12947,N_12349);
or U15304 (N_15304,N_13277,N_12901);
nor U15305 (N_15305,N_12689,N_13806);
and U15306 (N_15306,N_13898,N_12962);
nand U15307 (N_15307,N_13546,N_13003);
and U15308 (N_15308,N_12992,N_13963);
nand U15309 (N_15309,N_13127,N_12315);
nand U15310 (N_15310,N_13726,N_13768);
nor U15311 (N_15311,N_13712,N_13645);
or U15312 (N_15312,N_13516,N_12795);
nor U15313 (N_15313,N_12035,N_13185);
nand U15314 (N_15314,N_12678,N_12501);
and U15315 (N_15315,N_12238,N_13627);
xnor U15316 (N_15316,N_13186,N_12249);
or U15317 (N_15317,N_12413,N_13292);
nand U15318 (N_15318,N_12778,N_12987);
and U15319 (N_15319,N_12506,N_13629);
nand U15320 (N_15320,N_12561,N_12402);
or U15321 (N_15321,N_13842,N_13708);
nand U15322 (N_15322,N_13239,N_13907);
and U15323 (N_15323,N_12553,N_13825);
and U15324 (N_15324,N_13671,N_12601);
nand U15325 (N_15325,N_13103,N_13922);
or U15326 (N_15326,N_12718,N_13053);
nand U15327 (N_15327,N_13303,N_13762);
or U15328 (N_15328,N_13084,N_13737);
nand U15329 (N_15329,N_12169,N_12634);
nor U15330 (N_15330,N_13782,N_12095);
nand U15331 (N_15331,N_13870,N_12900);
and U15332 (N_15332,N_13190,N_13599);
nand U15333 (N_15333,N_12926,N_12522);
and U15334 (N_15334,N_12304,N_12060);
or U15335 (N_15335,N_13639,N_12113);
nor U15336 (N_15336,N_13831,N_12277);
and U15337 (N_15337,N_13325,N_12339);
nor U15338 (N_15338,N_12463,N_12607);
and U15339 (N_15339,N_13903,N_13524);
or U15340 (N_15340,N_13662,N_13181);
nand U15341 (N_15341,N_12586,N_12680);
nor U15342 (N_15342,N_12238,N_13227);
or U15343 (N_15343,N_12391,N_12033);
nor U15344 (N_15344,N_13640,N_12716);
nor U15345 (N_15345,N_13515,N_13022);
nand U15346 (N_15346,N_12794,N_12144);
nand U15347 (N_15347,N_12886,N_12276);
or U15348 (N_15348,N_13110,N_13921);
nor U15349 (N_15349,N_12729,N_13805);
nor U15350 (N_15350,N_13516,N_13202);
nor U15351 (N_15351,N_13593,N_12987);
nand U15352 (N_15352,N_13183,N_12698);
nor U15353 (N_15353,N_13681,N_12736);
nand U15354 (N_15354,N_13624,N_13261);
or U15355 (N_15355,N_13495,N_12435);
or U15356 (N_15356,N_12389,N_13197);
nor U15357 (N_15357,N_13420,N_12340);
nor U15358 (N_15358,N_12431,N_13075);
nor U15359 (N_15359,N_13524,N_13180);
or U15360 (N_15360,N_12794,N_13307);
or U15361 (N_15361,N_12395,N_12220);
and U15362 (N_15362,N_12472,N_13746);
and U15363 (N_15363,N_12934,N_13933);
or U15364 (N_15364,N_12262,N_12450);
and U15365 (N_15365,N_12701,N_13610);
nor U15366 (N_15366,N_12994,N_12718);
xor U15367 (N_15367,N_12903,N_12989);
nand U15368 (N_15368,N_13045,N_12553);
or U15369 (N_15369,N_12901,N_12071);
nor U15370 (N_15370,N_12395,N_13066);
or U15371 (N_15371,N_13006,N_13083);
nor U15372 (N_15372,N_12536,N_13543);
nor U15373 (N_15373,N_12369,N_13375);
nand U15374 (N_15374,N_13476,N_12880);
and U15375 (N_15375,N_13619,N_13884);
nand U15376 (N_15376,N_12304,N_12195);
and U15377 (N_15377,N_13610,N_12300);
nand U15378 (N_15378,N_13450,N_13176);
and U15379 (N_15379,N_13206,N_12508);
or U15380 (N_15380,N_12289,N_13305);
or U15381 (N_15381,N_13775,N_13677);
nor U15382 (N_15382,N_13167,N_12191);
xnor U15383 (N_15383,N_12064,N_12716);
and U15384 (N_15384,N_12793,N_13921);
and U15385 (N_15385,N_12567,N_13678);
and U15386 (N_15386,N_12174,N_12296);
or U15387 (N_15387,N_12219,N_13831);
and U15388 (N_15388,N_12747,N_12830);
nand U15389 (N_15389,N_13842,N_13333);
and U15390 (N_15390,N_12154,N_12140);
nand U15391 (N_15391,N_12616,N_13319);
nor U15392 (N_15392,N_13790,N_13471);
or U15393 (N_15393,N_13655,N_13644);
or U15394 (N_15394,N_12445,N_12221);
or U15395 (N_15395,N_13900,N_13048);
nor U15396 (N_15396,N_12881,N_12752);
nand U15397 (N_15397,N_12186,N_13411);
nor U15398 (N_15398,N_12807,N_13726);
nand U15399 (N_15399,N_13304,N_13628);
xor U15400 (N_15400,N_12792,N_13396);
nand U15401 (N_15401,N_12306,N_13355);
or U15402 (N_15402,N_13758,N_12276);
nand U15403 (N_15403,N_13966,N_12448);
xor U15404 (N_15404,N_13129,N_13336);
and U15405 (N_15405,N_12003,N_12653);
nor U15406 (N_15406,N_13664,N_12318);
nor U15407 (N_15407,N_13441,N_13960);
nand U15408 (N_15408,N_12599,N_12886);
and U15409 (N_15409,N_12918,N_13531);
and U15410 (N_15410,N_13908,N_13583);
nor U15411 (N_15411,N_12160,N_13926);
and U15412 (N_15412,N_12827,N_13423);
and U15413 (N_15413,N_13075,N_12652);
nor U15414 (N_15414,N_12527,N_12643);
nor U15415 (N_15415,N_13335,N_12136);
xor U15416 (N_15416,N_12039,N_12380);
and U15417 (N_15417,N_13336,N_12272);
or U15418 (N_15418,N_12822,N_12417);
nand U15419 (N_15419,N_12552,N_12753);
or U15420 (N_15420,N_12658,N_12310);
nor U15421 (N_15421,N_12009,N_13891);
nand U15422 (N_15422,N_13495,N_12907);
or U15423 (N_15423,N_13149,N_13704);
and U15424 (N_15424,N_12801,N_13339);
or U15425 (N_15425,N_12752,N_12017);
nor U15426 (N_15426,N_12876,N_13174);
nor U15427 (N_15427,N_13814,N_12041);
nor U15428 (N_15428,N_13586,N_13335);
or U15429 (N_15429,N_13410,N_13383);
or U15430 (N_15430,N_13291,N_12825);
and U15431 (N_15431,N_13616,N_13494);
xnor U15432 (N_15432,N_12008,N_12278);
and U15433 (N_15433,N_12446,N_12739);
xor U15434 (N_15434,N_13406,N_12074);
nor U15435 (N_15435,N_12646,N_13019);
nand U15436 (N_15436,N_13570,N_12074);
or U15437 (N_15437,N_13288,N_12631);
or U15438 (N_15438,N_13326,N_12232);
xor U15439 (N_15439,N_12752,N_12758);
nand U15440 (N_15440,N_12282,N_12426);
nor U15441 (N_15441,N_12794,N_13613);
nand U15442 (N_15442,N_13712,N_12918);
nor U15443 (N_15443,N_13862,N_13041);
or U15444 (N_15444,N_13330,N_12947);
and U15445 (N_15445,N_13302,N_12623);
and U15446 (N_15446,N_13733,N_13551);
nand U15447 (N_15447,N_13288,N_12898);
xnor U15448 (N_15448,N_13176,N_12262);
and U15449 (N_15449,N_13510,N_12626);
and U15450 (N_15450,N_12773,N_13743);
or U15451 (N_15451,N_12121,N_13216);
nand U15452 (N_15452,N_12092,N_13862);
xnor U15453 (N_15453,N_13803,N_12148);
or U15454 (N_15454,N_12223,N_13632);
nand U15455 (N_15455,N_12338,N_12881);
and U15456 (N_15456,N_13054,N_13804);
nand U15457 (N_15457,N_13864,N_12284);
nand U15458 (N_15458,N_13433,N_12709);
or U15459 (N_15459,N_12550,N_12099);
nand U15460 (N_15460,N_13918,N_12996);
nand U15461 (N_15461,N_13583,N_12781);
xor U15462 (N_15462,N_13928,N_12135);
or U15463 (N_15463,N_12269,N_13688);
xnor U15464 (N_15464,N_12973,N_13518);
and U15465 (N_15465,N_13348,N_13999);
or U15466 (N_15466,N_13769,N_13611);
nand U15467 (N_15467,N_12179,N_13977);
nor U15468 (N_15468,N_12116,N_13420);
nand U15469 (N_15469,N_13185,N_13104);
xor U15470 (N_15470,N_13977,N_13226);
or U15471 (N_15471,N_13736,N_12399);
or U15472 (N_15472,N_12783,N_13746);
nand U15473 (N_15473,N_13742,N_12135);
and U15474 (N_15474,N_13949,N_13304);
xnor U15475 (N_15475,N_13291,N_12089);
nand U15476 (N_15476,N_12482,N_12104);
and U15477 (N_15477,N_13710,N_13072);
and U15478 (N_15478,N_13078,N_12665);
and U15479 (N_15479,N_13708,N_13620);
xnor U15480 (N_15480,N_13418,N_13106);
nor U15481 (N_15481,N_12304,N_12344);
nor U15482 (N_15482,N_12384,N_13526);
and U15483 (N_15483,N_13730,N_12321);
or U15484 (N_15484,N_12809,N_12100);
and U15485 (N_15485,N_13201,N_12816);
or U15486 (N_15486,N_13282,N_12616);
nor U15487 (N_15487,N_13702,N_13003);
and U15488 (N_15488,N_13197,N_13542);
nand U15489 (N_15489,N_12046,N_12853);
or U15490 (N_15490,N_13283,N_13448);
and U15491 (N_15491,N_13290,N_13053);
nor U15492 (N_15492,N_12644,N_13412);
and U15493 (N_15493,N_12573,N_12862);
and U15494 (N_15494,N_12983,N_13166);
nand U15495 (N_15495,N_12002,N_12676);
nand U15496 (N_15496,N_13723,N_12059);
xnor U15497 (N_15497,N_13385,N_13823);
nor U15498 (N_15498,N_13920,N_13366);
or U15499 (N_15499,N_13260,N_12239);
or U15500 (N_15500,N_12414,N_13062);
and U15501 (N_15501,N_12131,N_13194);
and U15502 (N_15502,N_12295,N_13214);
or U15503 (N_15503,N_13374,N_12178);
and U15504 (N_15504,N_13131,N_13256);
or U15505 (N_15505,N_12952,N_12018);
nand U15506 (N_15506,N_13403,N_13057);
or U15507 (N_15507,N_13988,N_12742);
and U15508 (N_15508,N_13448,N_12549);
and U15509 (N_15509,N_12314,N_13632);
and U15510 (N_15510,N_13060,N_13884);
nand U15511 (N_15511,N_13149,N_12027);
or U15512 (N_15512,N_12280,N_13268);
xor U15513 (N_15513,N_13099,N_13112);
nand U15514 (N_15514,N_13876,N_12487);
xor U15515 (N_15515,N_13632,N_12519);
nor U15516 (N_15516,N_13741,N_13299);
or U15517 (N_15517,N_12111,N_12812);
and U15518 (N_15518,N_12469,N_13511);
and U15519 (N_15519,N_13727,N_13486);
nand U15520 (N_15520,N_12732,N_12706);
nor U15521 (N_15521,N_12266,N_13567);
nor U15522 (N_15522,N_12317,N_13684);
and U15523 (N_15523,N_13653,N_13119);
or U15524 (N_15524,N_13821,N_13848);
nor U15525 (N_15525,N_12899,N_13330);
xor U15526 (N_15526,N_13029,N_13667);
and U15527 (N_15527,N_13211,N_12688);
nor U15528 (N_15528,N_13071,N_13035);
nand U15529 (N_15529,N_12529,N_13812);
and U15530 (N_15530,N_13849,N_12797);
xor U15531 (N_15531,N_13498,N_12332);
nand U15532 (N_15532,N_12403,N_13651);
nand U15533 (N_15533,N_13695,N_13575);
nor U15534 (N_15534,N_12625,N_12455);
nand U15535 (N_15535,N_13769,N_13956);
nor U15536 (N_15536,N_13755,N_12735);
and U15537 (N_15537,N_13818,N_12816);
nor U15538 (N_15538,N_12664,N_12380);
nor U15539 (N_15539,N_12917,N_12653);
or U15540 (N_15540,N_13421,N_12961);
or U15541 (N_15541,N_12720,N_13692);
nor U15542 (N_15542,N_13058,N_12835);
or U15543 (N_15543,N_13117,N_13982);
or U15544 (N_15544,N_13004,N_12969);
and U15545 (N_15545,N_13691,N_13415);
and U15546 (N_15546,N_13855,N_12171);
or U15547 (N_15547,N_13381,N_12910);
or U15548 (N_15548,N_12596,N_12297);
or U15549 (N_15549,N_13665,N_13891);
nand U15550 (N_15550,N_13080,N_12507);
and U15551 (N_15551,N_13728,N_12504);
or U15552 (N_15552,N_12857,N_12418);
or U15553 (N_15553,N_13115,N_12102);
or U15554 (N_15554,N_12115,N_13189);
or U15555 (N_15555,N_12635,N_12281);
or U15556 (N_15556,N_13049,N_12992);
nor U15557 (N_15557,N_12197,N_13061);
nor U15558 (N_15558,N_12071,N_13866);
nor U15559 (N_15559,N_12966,N_13426);
nor U15560 (N_15560,N_13040,N_12038);
xor U15561 (N_15561,N_12754,N_13877);
nand U15562 (N_15562,N_12472,N_12381);
or U15563 (N_15563,N_12185,N_13708);
and U15564 (N_15564,N_12453,N_13448);
or U15565 (N_15565,N_12050,N_12395);
nand U15566 (N_15566,N_13093,N_12173);
and U15567 (N_15567,N_13130,N_12844);
nor U15568 (N_15568,N_13168,N_13334);
nor U15569 (N_15569,N_12076,N_12999);
nor U15570 (N_15570,N_13545,N_13387);
nand U15571 (N_15571,N_13408,N_13444);
xor U15572 (N_15572,N_13166,N_13696);
or U15573 (N_15573,N_13955,N_12733);
nor U15574 (N_15574,N_13075,N_13691);
or U15575 (N_15575,N_13569,N_13410);
nand U15576 (N_15576,N_13951,N_13016);
or U15577 (N_15577,N_13844,N_13611);
nor U15578 (N_15578,N_13505,N_13158);
or U15579 (N_15579,N_12402,N_12812);
or U15580 (N_15580,N_12337,N_12780);
or U15581 (N_15581,N_12755,N_12968);
xor U15582 (N_15582,N_13607,N_12875);
nand U15583 (N_15583,N_13092,N_12550);
xor U15584 (N_15584,N_12625,N_13149);
or U15585 (N_15585,N_13596,N_13791);
nand U15586 (N_15586,N_13507,N_12703);
nand U15587 (N_15587,N_13881,N_12634);
and U15588 (N_15588,N_13995,N_12997);
nand U15589 (N_15589,N_13383,N_13764);
and U15590 (N_15590,N_12927,N_12125);
nor U15591 (N_15591,N_13274,N_13443);
nor U15592 (N_15592,N_13301,N_13056);
and U15593 (N_15593,N_13928,N_12368);
nor U15594 (N_15594,N_13495,N_12905);
or U15595 (N_15595,N_13156,N_13561);
xnor U15596 (N_15596,N_13152,N_12930);
and U15597 (N_15597,N_12720,N_12307);
nand U15598 (N_15598,N_13191,N_13121);
nand U15599 (N_15599,N_13317,N_12099);
or U15600 (N_15600,N_13195,N_12805);
and U15601 (N_15601,N_13099,N_13468);
nor U15602 (N_15602,N_13641,N_12857);
nand U15603 (N_15603,N_13877,N_12225);
and U15604 (N_15604,N_12856,N_12827);
nor U15605 (N_15605,N_12106,N_12154);
nand U15606 (N_15606,N_13071,N_13723);
nor U15607 (N_15607,N_12738,N_12613);
nand U15608 (N_15608,N_12641,N_12596);
or U15609 (N_15609,N_12296,N_13537);
and U15610 (N_15610,N_12103,N_12336);
xnor U15611 (N_15611,N_13247,N_12236);
xnor U15612 (N_15612,N_13653,N_12150);
nor U15613 (N_15613,N_12886,N_13820);
and U15614 (N_15614,N_13985,N_13329);
nor U15615 (N_15615,N_13627,N_13490);
xor U15616 (N_15616,N_12643,N_12651);
nor U15617 (N_15617,N_13635,N_12703);
xor U15618 (N_15618,N_13022,N_13107);
nor U15619 (N_15619,N_13036,N_13130);
nand U15620 (N_15620,N_13123,N_13306);
and U15621 (N_15621,N_12010,N_12669);
or U15622 (N_15622,N_12913,N_13016);
nand U15623 (N_15623,N_13194,N_13500);
or U15624 (N_15624,N_12941,N_13467);
and U15625 (N_15625,N_12224,N_13664);
nand U15626 (N_15626,N_13295,N_12716);
nor U15627 (N_15627,N_12275,N_13423);
xnor U15628 (N_15628,N_13131,N_12830);
or U15629 (N_15629,N_13962,N_12173);
or U15630 (N_15630,N_13804,N_12065);
nor U15631 (N_15631,N_13483,N_12672);
nor U15632 (N_15632,N_12598,N_12786);
nor U15633 (N_15633,N_13825,N_13818);
nor U15634 (N_15634,N_13391,N_13551);
or U15635 (N_15635,N_13341,N_12137);
nor U15636 (N_15636,N_12386,N_13912);
nor U15637 (N_15637,N_12138,N_12750);
or U15638 (N_15638,N_13834,N_13698);
or U15639 (N_15639,N_13646,N_13551);
nor U15640 (N_15640,N_12450,N_13327);
or U15641 (N_15641,N_12318,N_12831);
nand U15642 (N_15642,N_12945,N_12954);
or U15643 (N_15643,N_13629,N_13917);
nand U15644 (N_15644,N_13282,N_13627);
or U15645 (N_15645,N_12297,N_12663);
and U15646 (N_15646,N_13565,N_13999);
nand U15647 (N_15647,N_13957,N_12314);
nand U15648 (N_15648,N_12066,N_12269);
nor U15649 (N_15649,N_12213,N_13588);
nand U15650 (N_15650,N_13600,N_12211);
or U15651 (N_15651,N_13824,N_12076);
nor U15652 (N_15652,N_12010,N_12146);
and U15653 (N_15653,N_13205,N_12016);
nor U15654 (N_15654,N_13353,N_12173);
xnor U15655 (N_15655,N_12102,N_12396);
nor U15656 (N_15656,N_12591,N_12660);
nor U15657 (N_15657,N_13471,N_12431);
or U15658 (N_15658,N_12866,N_12214);
and U15659 (N_15659,N_12439,N_13342);
nand U15660 (N_15660,N_13076,N_12532);
and U15661 (N_15661,N_13574,N_12721);
or U15662 (N_15662,N_12512,N_13261);
nor U15663 (N_15663,N_12283,N_13938);
and U15664 (N_15664,N_12769,N_13745);
and U15665 (N_15665,N_12875,N_12167);
or U15666 (N_15666,N_13443,N_13857);
nand U15667 (N_15667,N_12023,N_13766);
or U15668 (N_15668,N_12102,N_13307);
nor U15669 (N_15669,N_13774,N_12944);
nand U15670 (N_15670,N_13148,N_12404);
nand U15671 (N_15671,N_12969,N_12902);
nor U15672 (N_15672,N_12877,N_13540);
nand U15673 (N_15673,N_13645,N_13286);
nor U15674 (N_15674,N_12948,N_12899);
xnor U15675 (N_15675,N_12001,N_13962);
nand U15676 (N_15676,N_13869,N_12777);
nand U15677 (N_15677,N_12055,N_13007);
or U15678 (N_15678,N_13695,N_13667);
nand U15679 (N_15679,N_13899,N_12449);
or U15680 (N_15680,N_12793,N_12800);
nand U15681 (N_15681,N_13989,N_12287);
or U15682 (N_15682,N_12227,N_13638);
and U15683 (N_15683,N_13854,N_12270);
or U15684 (N_15684,N_12051,N_12890);
nor U15685 (N_15685,N_13119,N_13284);
xnor U15686 (N_15686,N_13138,N_12828);
nor U15687 (N_15687,N_12279,N_12707);
nand U15688 (N_15688,N_13394,N_13245);
or U15689 (N_15689,N_13850,N_13022);
nand U15690 (N_15690,N_12971,N_13208);
or U15691 (N_15691,N_12195,N_12666);
nor U15692 (N_15692,N_12761,N_12874);
and U15693 (N_15693,N_12641,N_13515);
and U15694 (N_15694,N_12414,N_13975);
and U15695 (N_15695,N_12949,N_12784);
and U15696 (N_15696,N_12673,N_13709);
nor U15697 (N_15697,N_13984,N_12204);
nor U15698 (N_15698,N_12777,N_13086);
nor U15699 (N_15699,N_12790,N_13851);
and U15700 (N_15700,N_13223,N_13806);
xnor U15701 (N_15701,N_12055,N_12676);
xor U15702 (N_15702,N_12164,N_12220);
and U15703 (N_15703,N_13766,N_12502);
and U15704 (N_15704,N_13444,N_12528);
nand U15705 (N_15705,N_12356,N_12691);
xnor U15706 (N_15706,N_12564,N_13441);
nand U15707 (N_15707,N_13413,N_12884);
xnor U15708 (N_15708,N_12545,N_12292);
nor U15709 (N_15709,N_12764,N_13425);
or U15710 (N_15710,N_12019,N_13143);
nand U15711 (N_15711,N_12386,N_13876);
or U15712 (N_15712,N_12612,N_12487);
nand U15713 (N_15713,N_13599,N_13228);
nand U15714 (N_15714,N_12868,N_13062);
or U15715 (N_15715,N_13081,N_13249);
and U15716 (N_15716,N_13415,N_13758);
nor U15717 (N_15717,N_13753,N_13835);
and U15718 (N_15718,N_12306,N_13280);
and U15719 (N_15719,N_13586,N_13552);
nand U15720 (N_15720,N_12283,N_12818);
nand U15721 (N_15721,N_13582,N_13887);
and U15722 (N_15722,N_12154,N_12935);
and U15723 (N_15723,N_13633,N_13749);
and U15724 (N_15724,N_13521,N_13318);
xnor U15725 (N_15725,N_13726,N_12503);
or U15726 (N_15726,N_13975,N_12485);
and U15727 (N_15727,N_13294,N_13099);
nor U15728 (N_15728,N_13353,N_13248);
nand U15729 (N_15729,N_12373,N_12383);
nor U15730 (N_15730,N_12009,N_12076);
nand U15731 (N_15731,N_13252,N_12098);
nand U15732 (N_15732,N_12688,N_12548);
or U15733 (N_15733,N_13137,N_12653);
xor U15734 (N_15734,N_13261,N_13342);
or U15735 (N_15735,N_12110,N_13631);
or U15736 (N_15736,N_12366,N_13470);
xnor U15737 (N_15737,N_12869,N_13445);
nand U15738 (N_15738,N_13288,N_13658);
nand U15739 (N_15739,N_13376,N_12151);
and U15740 (N_15740,N_13188,N_13945);
nand U15741 (N_15741,N_13939,N_13454);
nor U15742 (N_15742,N_13985,N_13327);
nor U15743 (N_15743,N_13760,N_13323);
and U15744 (N_15744,N_13093,N_13469);
or U15745 (N_15745,N_12887,N_12615);
xor U15746 (N_15746,N_13432,N_13509);
nand U15747 (N_15747,N_13330,N_12185);
and U15748 (N_15748,N_12778,N_13756);
and U15749 (N_15749,N_13270,N_12006);
nand U15750 (N_15750,N_13021,N_12929);
or U15751 (N_15751,N_12359,N_13877);
xor U15752 (N_15752,N_12232,N_12865);
nand U15753 (N_15753,N_12822,N_13383);
xnor U15754 (N_15754,N_13325,N_13310);
nor U15755 (N_15755,N_13519,N_13193);
or U15756 (N_15756,N_12790,N_13005);
nand U15757 (N_15757,N_13601,N_13642);
or U15758 (N_15758,N_12620,N_12611);
xnor U15759 (N_15759,N_13658,N_12439);
or U15760 (N_15760,N_12199,N_13967);
nand U15761 (N_15761,N_12076,N_13434);
nand U15762 (N_15762,N_13915,N_12290);
nand U15763 (N_15763,N_12219,N_13024);
or U15764 (N_15764,N_12227,N_13308);
nor U15765 (N_15765,N_13687,N_13269);
or U15766 (N_15766,N_12759,N_12804);
or U15767 (N_15767,N_12273,N_12377);
and U15768 (N_15768,N_12920,N_12375);
nand U15769 (N_15769,N_13869,N_13755);
and U15770 (N_15770,N_13937,N_12016);
nor U15771 (N_15771,N_13070,N_12262);
and U15772 (N_15772,N_13247,N_13141);
xor U15773 (N_15773,N_12422,N_13717);
nand U15774 (N_15774,N_12414,N_12377);
and U15775 (N_15775,N_12986,N_13588);
nand U15776 (N_15776,N_13676,N_12686);
nor U15777 (N_15777,N_12373,N_13972);
and U15778 (N_15778,N_12547,N_12293);
and U15779 (N_15779,N_13341,N_13827);
nand U15780 (N_15780,N_12606,N_12930);
nand U15781 (N_15781,N_13234,N_12860);
and U15782 (N_15782,N_13797,N_13784);
or U15783 (N_15783,N_12946,N_12300);
or U15784 (N_15784,N_13827,N_13140);
xor U15785 (N_15785,N_13443,N_13991);
nor U15786 (N_15786,N_12130,N_12860);
xnor U15787 (N_15787,N_13598,N_13703);
nand U15788 (N_15788,N_12207,N_12156);
nor U15789 (N_15789,N_12215,N_13058);
xnor U15790 (N_15790,N_13880,N_13397);
nor U15791 (N_15791,N_12425,N_13287);
nand U15792 (N_15792,N_13733,N_13222);
nand U15793 (N_15793,N_12598,N_13376);
nor U15794 (N_15794,N_13053,N_12889);
or U15795 (N_15795,N_12235,N_13914);
or U15796 (N_15796,N_13174,N_13717);
nor U15797 (N_15797,N_12222,N_13013);
and U15798 (N_15798,N_12820,N_13279);
or U15799 (N_15799,N_13392,N_13246);
nor U15800 (N_15800,N_13055,N_13111);
and U15801 (N_15801,N_12295,N_13615);
nand U15802 (N_15802,N_12071,N_13594);
or U15803 (N_15803,N_12352,N_12183);
nor U15804 (N_15804,N_13193,N_12114);
nand U15805 (N_15805,N_12739,N_12653);
and U15806 (N_15806,N_13678,N_13278);
and U15807 (N_15807,N_13164,N_12819);
nand U15808 (N_15808,N_12594,N_13084);
and U15809 (N_15809,N_13939,N_13065);
and U15810 (N_15810,N_12288,N_13215);
nand U15811 (N_15811,N_12450,N_12999);
xnor U15812 (N_15812,N_13515,N_13981);
or U15813 (N_15813,N_13104,N_13828);
nor U15814 (N_15814,N_12192,N_12438);
or U15815 (N_15815,N_12764,N_13143);
xor U15816 (N_15816,N_12983,N_12729);
nand U15817 (N_15817,N_12884,N_12549);
nor U15818 (N_15818,N_12725,N_12098);
nand U15819 (N_15819,N_13028,N_12307);
or U15820 (N_15820,N_13051,N_12228);
or U15821 (N_15821,N_12435,N_12767);
or U15822 (N_15822,N_13393,N_12944);
nand U15823 (N_15823,N_13052,N_13229);
or U15824 (N_15824,N_12546,N_13383);
nor U15825 (N_15825,N_12737,N_12705);
nand U15826 (N_15826,N_12194,N_13844);
and U15827 (N_15827,N_12380,N_12264);
nand U15828 (N_15828,N_12284,N_12185);
and U15829 (N_15829,N_12408,N_12894);
and U15830 (N_15830,N_13052,N_12189);
xor U15831 (N_15831,N_13129,N_13690);
nand U15832 (N_15832,N_12268,N_12432);
nand U15833 (N_15833,N_12270,N_13979);
nand U15834 (N_15834,N_13392,N_13374);
nand U15835 (N_15835,N_13292,N_12157);
nor U15836 (N_15836,N_12268,N_12185);
nand U15837 (N_15837,N_12188,N_12614);
nor U15838 (N_15838,N_13529,N_12562);
nand U15839 (N_15839,N_12331,N_12063);
and U15840 (N_15840,N_13539,N_13421);
or U15841 (N_15841,N_13200,N_13879);
and U15842 (N_15842,N_12740,N_13133);
or U15843 (N_15843,N_12645,N_12708);
and U15844 (N_15844,N_13604,N_12236);
nor U15845 (N_15845,N_13443,N_13678);
or U15846 (N_15846,N_13962,N_13729);
nand U15847 (N_15847,N_12916,N_12394);
nor U15848 (N_15848,N_12107,N_12870);
nor U15849 (N_15849,N_13743,N_12288);
nor U15850 (N_15850,N_12633,N_13985);
xor U15851 (N_15851,N_13236,N_12505);
nand U15852 (N_15852,N_12630,N_13327);
nor U15853 (N_15853,N_12730,N_13984);
xnor U15854 (N_15854,N_13994,N_12178);
and U15855 (N_15855,N_13415,N_12883);
nand U15856 (N_15856,N_13232,N_12379);
or U15857 (N_15857,N_13836,N_13151);
and U15858 (N_15858,N_12933,N_13650);
xor U15859 (N_15859,N_13707,N_12297);
nor U15860 (N_15860,N_12122,N_12473);
nor U15861 (N_15861,N_13482,N_13976);
and U15862 (N_15862,N_12630,N_13265);
nand U15863 (N_15863,N_13814,N_13143);
or U15864 (N_15864,N_13831,N_12896);
and U15865 (N_15865,N_13537,N_12300);
nor U15866 (N_15866,N_12354,N_12274);
nand U15867 (N_15867,N_13472,N_12414);
nand U15868 (N_15868,N_12188,N_13738);
nand U15869 (N_15869,N_12587,N_12289);
xnor U15870 (N_15870,N_12487,N_12103);
xor U15871 (N_15871,N_12570,N_13951);
nand U15872 (N_15872,N_13449,N_12711);
nor U15873 (N_15873,N_12438,N_13903);
xor U15874 (N_15874,N_12281,N_12297);
or U15875 (N_15875,N_13138,N_12248);
and U15876 (N_15876,N_12834,N_12978);
and U15877 (N_15877,N_13727,N_12405);
or U15878 (N_15878,N_12668,N_12895);
or U15879 (N_15879,N_13303,N_13923);
or U15880 (N_15880,N_12404,N_13554);
xnor U15881 (N_15881,N_12432,N_12369);
and U15882 (N_15882,N_12240,N_12910);
or U15883 (N_15883,N_13422,N_13094);
and U15884 (N_15884,N_13717,N_12356);
nand U15885 (N_15885,N_13635,N_12642);
xor U15886 (N_15886,N_13024,N_12371);
or U15887 (N_15887,N_12592,N_12953);
or U15888 (N_15888,N_13025,N_13420);
nand U15889 (N_15889,N_13381,N_13690);
nor U15890 (N_15890,N_13338,N_13689);
nand U15891 (N_15891,N_13631,N_12005);
nand U15892 (N_15892,N_13686,N_13863);
and U15893 (N_15893,N_13008,N_13791);
or U15894 (N_15894,N_13380,N_13157);
nand U15895 (N_15895,N_13057,N_12248);
xnor U15896 (N_15896,N_13326,N_12434);
and U15897 (N_15897,N_13663,N_12485);
and U15898 (N_15898,N_13471,N_13100);
nand U15899 (N_15899,N_13629,N_12689);
nor U15900 (N_15900,N_13882,N_12200);
and U15901 (N_15901,N_13959,N_13179);
nand U15902 (N_15902,N_12779,N_13788);
nand U15903 (N_15903,N_12648,N_13950);
and U15904 (N_15904,N_13114,N_13977);
nand U15905 (N_15905,N_13279,N_12178);
and U15906 (N_15906,N_13565,N_13725);
or U15907 (N_15907,N_13953,N_12665);
xnor U15908 (N_15908,N_13470,N_13028);
and U15909 (N_15909,N_12683,N_12782);
and U15910 (N_15910,N_13380,N_13384);
or U15911 (N_15911,N_12778,N_13430);
nor U15912 (N_15912,N_12022,N_13351);
or U15913 (N_15913,N_13062,N_12111);
and U15914 (N_15914,N_13837,N_12353);
or U15915 (N_15915,N_12411,N_13868);
nor U15916 (N_15916,N_12310,N_13774);
nor U15917 (N_15917,N_12043,N_12798);
nor U15918 (N_15918,N_12554,N_12730);
nor U15919 (N_15919,N_13489,N_12706);
nand U15920 (N_15920,N_13690,N_13804);
xnor U15921 (N_15921,N_13024,N_12760);
and U15922 (N_15922,N_13524,N_12402);
nand U15923 (N_15923,N_13497,N_12029);
or U15924 (N_15924,N_13331,N_13706);
nand U15925 (N_15925,N_12451,N_13878);
nor U15926 (N_15926,N_13459,N_12206);
xor U15927 (N_15927,N_12959,N_13679);
and U15928 (N_15928,N_13040,N_13530);
or U15929 (N_15929,N_13120,N_12400);
nor U15930 (N_15930,N_12578,N_13047);
nor U15931 (N_15931,N_12072,N_13635);
nor U15932 (N_15932,N_12191,N_12164);
nand U15933 (N_15933,N_12120,N_12813);
nand U15934 (N_15934,N_12345,N_13741);
or U15935 (N_15935,N_12983,N_12785);
nand U15936 (N_15936,N_12369,N_13288);
and U15937 (N_15937,N_13053,N_12273);
nor U15938 (N_15938,N_12030,N_12362);
nor U15939 (N_15939,N_12618,N_12480);
and U15940 (N_15940,N_12331,N_13095);
or U15941 (N_15941,N_12853,N_13837);
and U15942 (N_15942,N_13201,N_12739);
nor U15943 (N_15943,N_13708,N_13210);
xnor U15944 (N_15944,N_13001,N_12514);
nor U15945 (N_15945,N_12036,N_12340);
or U15946 (N_15946,N_12293,N_13889);
nand U15947 (N_15947,N_13429,N_13487);
xnor U15948 (N_15948,N_12023,N_12391);
or U15949 (N_15949,N_12224,N_13696);
or U15950 (N_15950,N_12627,N_12266);
and U15951 (N_15951,N_12922,N_12217);
nand U15952 (N_15952,N_13560,N_13831);
nor U15953 (N_15953,N_13375,N_13744);
nand U15954 (N_15954,N_12490,N_13813);
or U15955 (N_15955,N_13533,N_13390);
nor U15956 (N_15956,N_13319,N_13389);
nand U15957 (N_15957,N_12883,N_13647);
nor U15958 (N_15958,N_12114,N_13897);
or U15959 (N_15959,N_12393,N_13857);
nor U15960 (N_15960,N_13097,N_13945);
and U15961 (N_15961,N_12110,N_13480);
and U15962 (N_15962,N_12250,N_13445);
and U15963 (N_15963,N_13373,N_12456);
nand U15964 (N_15964,N_12516,N_13445);
xnor U15965 (N_15965,N_12277,N_13903);
nand U15966 (N_15966,N_13247,N_12494);
nor U15967 (N_15967,N_13720,N_12704);
nand U15968 (N_15968,N_13442,N_13740);
and U15969 (N_15969,N_12500,N_13288);
and U15970 (N_15970,N_13599,N_13528);
nand U15971 (N_15971,N_12019,N_13827);
nand U15972 (N_15972,N_13657,N_12457);
or U15973 (N_15973,N_13514,N_13130);
and U15974 (N_15974,N_12324,N_12037);
or U15975 (N_15975,N_13639,N_13273);
nor U15976 (N_15976,N_13410,N_13424);
and U15977 (N_15977,N_12180,N_13375);
nand U15978 (N_15978,N_13458,N_13085);
or U15979 (N_15979,N_12216,N_13076);
or U15980 (N_15980,N_12385,N_12919);
xnor U15981 (N_15981,N_12730,N_12903);
or U15982 (N_15982,N_12864,N_13374);
and U15983 (N_15983,N_12524,N_12052);
xor U15984 (N_15984,N_13522,N_13639);
nor U15985 (N_15985,N_13391,N_13650);
nand U15986 (N_15986,N_13160,N_13411);
nor U15987 (N_15987,N_12079,N_13488);
xnor U15988 (N_15988,N_12497,N_13260);
nand U15989 (N_15989,N_13572,N_12337);
or U15990 (N_15990,N_12540,N_13048);
nand U15991 (N_15991,N_12015,N_12402);
nor U15992 (N_15992,N_13794,N_13409);
or U15993 (N_15993,N_13169,N_13669);
and U15994 (N_15994,N_12066,N_13117);
nor U15995 (N_15995,N_13856,N_12975);
nand U15996 (N_15996,N_12131,N_13860);
nor U15997 (N_15997,N_13017,N_13114);
and U15998 (N_15998,N_13455,N_12953);
or U15999 (N_15999,N_13356,N_12281);
xnor U16000 (N_16000,N_14961,N_14756);
and U16001 (N_16001,N_15767,N_15028);
nand U16002 (N_16002,N_15919,N_14579);
and U16003 (N_16003,N_15838,N_15494);
and U16004 (N_16004,N_14947,N_15759);
and U16005 (N_16005,N_14030,N_15887);
nor U16006 (N_16006,N_15289,N_14470);
nand U16007 (N_16007,N_15492,N_15757);
nand U16008 (N_16008,N_14158,N_15634);
xor U16009 (N_16009,N_15804,N_15422);
or U16010 (N_16010,N_14498,N_15642);
nand U16011 (N_16011,N_15976,N_14363);
or U16012 (N_16012,N_15936,N_15091);
nand U16013 (N_16013,N_14207,N_14502);
nand U16014 (N_16014,N_14668,N_14051);
xnor U16015 (N_16015,N_15139,N_14737);
nor U16016 (N_16016,N_14827,N_15453);
nor U16017 (N_16017,N_15507,N_15533);
nor U16018 (N_16018,N_14707,N_14350);
xor U16019 (N_16019,N_14681,N_15032);
nor U16020 (N_16020,N_14073,N_14962);
nand U16021 (N_16021,N_14763,N_15275);
nor U16022 (N_16022,N_14764,N_15914);
and U16023 (N_16023,N_14314,N_14919);
and U16024 (N_16024,N_15077,N_15547);
or U16025 (N_16025,N_15538,N_15308);
nor U16026 (N_16026,N_14289,N_14606);
and U16027 (N_16027,N_14824,N_14679);
nor U16028 (N_16028,N_15482,N_15956);
nor U16029 (N_16029,N_14615,N_14375);
nor U16030 (N_16030,N_14297,N_15774);
and U16031 (N_16031,N_14166,N_14012);
nor U16032 (N_16032,N_15543,N_14123);
and U16033 (N_16033,N_14813,N_15444);
nor U16034 (N_16034,N_14230,N_15886);
nor U16035 (N_16035,N_15400,N_15729);
nand U16036 (N_16036,N_14234,N_14743);
nand U16037 (N_16037,N_14674,N_15655);
nand U16038 (N_16038,N_15063,N_14370);
or U16039 (N_16039,N_14432,N_14990);
and U16040 (N_16040,N_14277,N_15626);
nor U16041 (N_16041,N_14496,N_14634);
xnor U16042 (N_16042,N_15391,N_15302);
or U16043 (N_16043,N_15163,N_15814);
or U16044 (N_16044,N_14165,N_15145);
nor U16045 (N_16045,N_14531,N_14902);
and U16046 (N_16046,N_14630,N_14141);
nand U16047 (N_16047,N_14362,N_14868);
and U16048 (N_16048,N_15446,N_14759);
or U16049 (N_16049,N_14895,N_14656);
nor U16050 (N_16050,N_14617,N_15932);
and U16051 (N_16051,N_15604,N_14105);
or U16052 (N_16052,N_15281,N_15044);
and U16053 (N_16053,N_15342,N_14768);
nand U16054 (N_16054,N_14677,N_15871);
or U16055 (N_16055,N_14908,N_15349);
xor U16056 (N_16056,N_14678,N_15094);
nand U16057 (N_16057,N_15640,N_14042);
or U16058 (N_16058,N_15466,N_14089);
and U16059 (N_16059,N_14332,N_14811);
or U16060 (N_16060,N_14407,N_14875);
or U16061 (N_16061,N_15568,N_15065);
and U16062 (N_16062,N_14406,N_15361);
nand U16063 (N_16063,N_15898,N_15001);
nor U16064 (N_16064,N_15389,N_14561);
xnor U16065 (N_16065,N_15068,N_14219);
and U16066 (N_16066,N_15980,N_14456);
or U16067 (N_16067,N_15676,N_15681);
or U16068 (N_16068,N_15500,N_14146);
or U16069 (N_16069,N_14083,N_14680);
nor U16070 (N_16070,N_14322,N_14433);
nor U16071 (N_16071,N_15020,N_14003);
nand U16072 (N_16072,N_15786,N_14575);
nor U16073 (N_16073,N_14608,N_15623);
and U16074 (N_16074,N_14514,N_15504);
xor U16075 (N_16075,N_15196,N_15419);
or U16076 (N_16076,N_14556,N_14356);
or U16077 (N_16077,N_15917,N_14404);
nor U16078 (N_16078,N_15114,N_15645);
nor U16079 (N_16079,N_15227,N_15599);
and U16080 (N_16080,N_15692,N_14592);
and U16081 (N_16081,N_15570,N_15230);
nor U16082 (N_16082,N_14955,N_14929);
or U16083 (N_16083,N_14671,N_14390);
or U16084 (N_16084,N_14121,N_14884);
or U16085 (N_16085,N_15356,N_14348);
or U16086 (N_16086,N_15884,N_15141);
nor U16087 (N_16087,N_14582,N_14232);
or U16088 (N_16088,N_15684,N_14388);
nor U16089 (N_16089,N_15637,N_14347);
and U16090 (N_16090,N_15474,N_14437);
nor U16091 (N_16091,N_15173,N_15407);
and U16092 (N_16092,N_15732,N_14274);
or U16093 (N_16093,N_15841,N_15123);
or U16094 (N_16094,N_14765,N_15140);
or U16095 (N_16095,N_14292,N_14488);
or U16096 (N_16096,N_14562,N_14978);
or U16097 (N_16097,N_14966,N_14174);
and U16098 (N_16098,N_15095,N_14021);
or U16099 (N_16099,N_15338,N_15221);
nand U16100 (N_16100,N_14068,N_14914);
nor U16101 (N_16101,N_14633,N_15927);
xor U16102 (N_16102,N_15172,N_15184);
nor U16103 (N_16103,N_15495,N_14169);
and U16104 (N_16104,N_14381,N_14031);
nand U16105 (N_16105,N_14983,N_14129);
or U16106 (N_16106,N_15499,N_15788);
or U16107 (N_16107,N_15084,N_15042);
and U16108 (N_16108,N_15475,N_14980);
nor U16109 (N_16109,N_14741,N_14610);
and U16110 (N_16110,N_15742,N_14076);
and U16111 (N_16111,N_15376,N_15697);
xnor U16112 (N_16112,N_15341,N_14593);
nor U16113 (N_16113,N_14410,N_15987);
or U16114 (N_16114,N_15049,N_14518);
nand U16115 (N_16115,N_14070,N_14194);
nor U16116 (N_16116,N_15970,N_15563);
xnor U16117 (N_16117,N_15310,N_14760);
or U16118 (N_16118,N_14327,N_15487);
nand U16119 (N_16119,N_14913,N_15279);
nor U16120 (N_16120,N_14310,N_14171);
nand U16121 (N_16121,N_15022,N_15188);
nand U16122 (N_16122,N_14443,N_15229);
and U16123 (N_16123,N_15519,N_14584);
nor U16124 (N_16124,N_15392,N_15307);
nand U16125 (N_16125,N_15223,N_15778);
nor U16126 (N_16126,N_14773,N_14215);
nand U16127 (N_16127,N_14001,N_15268);
nor U16128 (N_16128,N_14689,N_15910);
nand U16129 (N_16129,N_14987,N_14863);
nor U16130 (N_16130,N_14134,N_15581);
nor U16131 (N_16131,N_14936,N_14039);
nand U16132 (N_16132,N_15794,N_14871);
or U16133 (N_16133,N_15964,N_14300);
and U16134 (N_16134,N_15561,N_14816);
nand U16135 (N_16135,N_14874,N_14452);
nand U16136 (N_16136,N_14211,N_14270);
or U16137 (N_16137,N_15263,N_14035);
nor U16138 (N_16138,N_14798,N_15282);
nor U16139 (N_16139,N_15240,N_14503);
or U16140 (N_16140,N_15710,N_15434);
nand U16141 (N_16141,N_14355,N_15408);
nor U16142 (N_16142,N_14185,N_14571);
nor U16143 (N_16143,N_14053,N_14711);
and U16144 (N_16144,N_15923,N_14702);
nand U16145 (N_16145,N_15251,N_14724);
nand U16146 (N_16146,N_15336,N_15206);
nor U16147 (N_16147,N_14264,N_14534);
or U16148 (N_16148,N_15174,N_14117);
nor U16149 (N_16149,N_15217,N_14436);
nor U16150 (N_16150,N_14500,N_14393);
xor U16151 (N_16151,N_15860,N_14049);
nand U16152 (N_16152,N_14576,N_15238);
and U16153 (N_16153,N_15702,N_14193);
or U16154 (N_16154,N_15369,N_14590);
or U16155 (N_16155,N_14081,N_15394);
nand U16156 (N_16156,N_15505,N_15802);
nand U16157 (N_16157,N_14563,N_14434);
nand U16158 (N_16158,N_15573,N_15854);
nand U16159 (N_16159,N_15317,N_14027);
and U16160 (N_16160,N_14646,N_15214);
nor U16161 (N_16161,N_15806,N_15647);
and U16162 (N_16162,N_14361,N_15678);
and U16163 (N_16163,N_15993,N_15904);
and U16164 (N_16164,N_14014,N_15508);
nor U16165 (N_16165,N_15971,N_15087);
and U16166 (N_16166,N_15824,N_14682);
and U16167 (N_16167,N_14537,N_14334);
nor U16168 (N_16168,N_15200,N_15579);
or U16169 (N_16169,N_14420,N_14530);
nand U16170 (N_16170,N_15189,N_15406);
nor U16171 (N_16171,N_14916,N_14609);
nor U16172 (N_16172,N_14542,N_15630);
and U16173 (N_16173,N_14687,N_15056);
nor U16174 (N_16174,N_14308,N_14795);
and U16175 (N_16175,N_15447,N_15479);
nor U16176 (N_16176,N_14387,N_14822);
or U16177 (N_16177,N_15975,N_14898);
nor U16178 (N_16178,N_15602,N_14323);
xor U16179 (N_16179,N_15117,N_15705);
nor U16180 (N_16180,N_15823,N_14440);
or U16181 (N_16181,N_14170,N_15297);
and U16182 (N_16182,N_14360,N_15764);
and U16183 (N_16183,N_14047,N_15986);
nand U16184 (N_16184,N_14940,N_15513);
nor U16185 (N_16185,N_15978,N_14541);
or U16186 (N_16186,N_15018,N_15339);
and U16187 (N_16187,N_14907,N_14447);
nor U16188 (N_16188,N_14048,N_15252);
and U16189 (N_16189,N_14302,N_15286);
or U16190 (N_16190,N_14621,N_15512);
nor U16191 (N_16191,N_14739,N_15261);
nand U16192 (N_16192,N_14338,N_15826);
nand U16193 (N_16193,N_14629,N_14993);
xnor U16194 (N_16194,N_15578,N_15365);
or U16195 (N_16195,N_15734,N_15291);
nor U16196 (N_16196,N_14754,N_15878);
and U16197 (N_16197,N_15869,N_15137);
nand U16198 (N_16198,N_14623,N_14945);
nand U16199 (N_16199,N_15690,N_15663);
nor U16200 (N_16200,N_15309,N_15435);
or U16201 (N_16201,N_14934,N_14192);
xor U16202 (N_16202,N_15799,N_14212);
or U16203 (N_16203,N_14142,N_14915);
nor U16204 (N_16204,N_15785,N_14830);
nor U16205 (N_16205,N_14365,N_15484);
nor U16206 (N_16206,N_15059,N_15709);
and U16207 (N_16207,N_14971,N_15190);
nand U16208 (N_16208,N_14717,N_14122);
xnor U16209 (N_16209,N_15670,N_15329);
nand U16210 (N_16210,N_14368,N_15193);
or U16211 (N_16211,N_15074,N_14278);
nor U16212 (N_16212,N_15235,N_15704);
nand U16213 (N_16213,N_15575,N_14311);
or U16214 (N_16214,N_15314,N_14226);
nor U16215 (N_16215,N_15582,N_14402);
and U16216 (N_16216,N_14451,N_15572);
or U16217 (N_16217,N_14112,N_14793);
nand U16218 (N_16218,N_14878,N_14482);
and U16219 (N_16219,N_15565,N_14660);
or U16220 (N_16220,N_14897,N_14599);
and U16221 (N_16221,N_15585,N_15038);
or U16222 (N_16222,N_14869,N_15649);
or U16223 (N_16223,N_15344,N_15070);
nand U16224 (N_16224,N_14565,N_14927);
or U16225 (N_16225,N_15384,N_15102);
and U16226 (N_16226,N_14886,N_15366);
nand U16227 (N_16227,N_14742,N_15320);
nor U16228 (N_16228,N_14719,N_15693);
nor U16229 (N_16229,N_14789,N_14011);
or U16230 (N_16230,N_15559,N_14686);
nor U16231 (N_16231,N_15187,N_15061);
nand U16232 (N_16232,N_15107,N_14981);
or U16233 (N_16233,N_14631,N_14034);
and U16234 (N_16234,N_14342,N_14135);
nor U16235 (N_16235,N_15280,N_15201);
or U16236 (N_16236,N_15592,N_15008);
nor U16237 (N_16237,N_15560,N_15237);
and U16238 (N_16238,N_15873,N_15371);
or U16239 (N_16239,N_14844,N_14823);
xor U16240 (N_16240,N_15192,N_14239);
nand U16241 (N_16241,N_15925,N_14540);
nand U16242 (N_16242,N_15766,N_14849);
xor U16243 (N_16243,N_15161,N_14516);
and U16244 (N_16244,N_15821,N_15135);
and U16245 (N_16245,N_15072,N_14168);
nand U16246 (N_16246,N_14473,N_14797);
nand U16247 (N_16247,N_15333,N_14603);
nand U16248 (N_16248,N_14800,N_14507);
nand U16249 (N_16249,N_15820,N_15829);
nor U16250 (N_16250,N_15224,N_15103);
nor U16251 (N_16251,N_15959,N_15451);
or U16252 (N_16252,N_14524,N_15058);
or U16253 (N_16253,N_15553,N_15773);
and U16254 (N_16254,N_14956,N_15834);
nor U16255 (N_16255,N_14727,N_14517);
xor U16256 (N_16256,N_14474,N_15298);
nand U16257 (N_16257,N_14029,N_14377);
nand U16258 (N_16258,N_14512,N_14358);
and U16259 (N_16259,N_15427,N_14326);
and U16260 (N_16260,N_14731,N_15374);
nand U16261 (N_16261,N_15946,N_14810);
or U16262 (N_16262,N_15675,N_15777);
and U16263 (N_16263,N_15737,N_14072);
and U16264 (N_16264,N_15536,N_15597);
nand U16265 (N_16265,N_15381,N_14832);
and U16266 (N_16266,N_14475,N_14803);
and U16267 (N_16267,N_14700,N_14380);
nand U16268 (N_16268,N_14867,N_15567);
nor U16269 (N_16269,N_14179,N_15480);
nand U16270 (N_16270,N_14228,N_14222);
or U16271 (N_16271,N_14002,N_14588);
and U16272 (N_16272,N_14062,N_14325);
nand U16273 (N_16273,N_15246,N_15701);
and U16274 (N_16274,N_14263,N_15832);
or U16275 (N_16275,N_15088,N_15177);
and U16276 (N_16276,N_14244,N_15648);
nor U16277 (N_16277,N_14779,N_14113);
nand U16278 (N_16278,N_14722,N_14735);
nand U16279 (N_16279,N_15706,N_14762);
or U16280 (N_16280,N_15111,N_15194);
nor U16281 (N_16281,N_15358,N_15875);
nand U16282 (N_16282,N_15528,N_14594);
xor U16283 (N_16283,N_14152,N_14710);
nor U16284 (N_16284,N_14831,N_15907);
and U16285 (N_16285,N_14783,N_14359);
and U16286 (N_16286,N_15283,N_14213);
and U16287 (N_16287,N_15254,N_14706);
or U16288 (N_16288,N_15347,N_14885);
or U16289 (N_16289,N_15885,N_14801);
xor U16290 (N_16290,N_14665,N_15036);
or U16291 (N_16291,N_15698,N_14748);
and U16292 (N_16292,N_15324,N_14218);
nor U16293 (N_16293,N_15541,N_15781);
nor U16294 (N_16294,N_15149,N_15746);
and U16295 (N_16295,N_14843,N_14953);
nand U16296 (N_16296,N_14412,N_14196);
or U16297 (N_16297,N_15784,N_14840);
nor U16298 (N_16298,N_15245,N_15849);
and U16299 (N_16299,N_14495,N_14111);
and U16300 (N_16300,N_14837,N_15856);
or U16301 (N_16301,N_15301,N_14604);
and U16302 (N_16302,N_15362,N_14970);
nand U16303 (N_16303,N_15656,N_15954);
or U16304 (N_16304,N_14125,N_15273);
or U16305 (N_16305,N_14544,N_15468);
and U16306 (N_16306,N_15127,N_14619);
xnor U16307 (N_16307,N_15464,N_14890);
nand U16308 (N_16308,N_14371,N_14769);
or U16309 (N_16309,N_15580,N_14454);
and U16310 (N_16310,N_15285,N_14572);
xnor U16311 (N_16311,N_14964,N_15712);
or U16312 (N_16312,N_14835,N_15981);
nand U16313 (N_16313,N_14613,N_14648);
nand U16314 (N_16314,N_14161,N_14600);
and U16315 (N_16315,N_14464,N_14386);
or U16316 (N_16316,N_15544,N_14357);
or U16317 (N_16317,N_14257,N_14643);
and U16318 (N_16318,N_14805,N_14785);
xor U16319 (N_16319,N_15164,N_14792);
and U16320 (N_16320,N_14189,N_15731);
nand U16321 (N_16321,N_14519,N_15311);
or U16322 (N_16322,N_15379,N_15303);
and U16323 (N_16323,N_14344,N_14296);
nand U16324 (N_16324,N_15319,N_15334);
nand U16325 (N_16325,N_15169,N_14016);
xor U16326 (N_16326,N_14972,N_15598);
or U16327 (N_16327,N_15352,N_15894);
xor U16328 (N_16328,N_15724,N_14336);
nor U16329 (N_16329,N_15006,N_15614);
and U16330 (N_16330,N_15234,N_14261);
nand U16331 (N_16331,N_15958,N_15934);
nand U16332 (N_16332,N_14243,N_14578);
nand U16333 (N_16333,N_14143,N_14485);
or U16334 (N_16334,N_15753,N_15048);
nor U16335 (N_16335,N_14490,N_14399);
or U16336 (N_16336,N_14108,N_14777);
and U16337 (N_16337,N_15853,N_15079);
or U16338 (N_16338,N_14538,N_15158);
or U16339 (N_16339,N_14431,N_15514);
or U16340 (N_16340,N_14557,N_14715);
nor U16341 (N_16341,N_14397,N_14683);
or U16342 (N_16342,N_14909,N_15331);
and U16343 (N_16343,N_14351,N_15714);
xor U16344 (N_16344,N_15481,N_14667);
and U16345 (N_16345,N_15857,N_15034);
nor U16346 (N_16346,N_14893,N_15168);
and U16347 (N_16347,N_15299,N_14231);
and U16348 (N_16348,N_15638,N_15616);
and U16349 (N_16349,N_15160,N_15862);
and U16350 (N_16350,N_14267,N_15920);
nor U16351 (N_16351,N_14664,N_14471);
nand U16352 (N_16352,N_14254,N_15052);
nand U16353 (N_16353,N_14761,N_14223);
xnor U16354 (N_16354,N_15636,N_14271);
nor U16355 (N_16355,N_14333,N_14088);
nand U16356 (N_16356,N_14453,N_15571);
and U16357 (N_16357,N_14820,N_15534);
xnor U16358 (N_16358,N_15325,N_15618);
nor U16359 (N_16359,N_15467,N_15968);
or U16360 (N_16360,N_15888,N_15688);
and U16361 (N_16361,N_14494,N_14533);
and U16362 (N_16362,N_14558,N_15367);
nor U16363 (N_16363,N_15625,N_15249);
nor U16364 (N_16364,N_14888,N_14589);
and U16365 (N_16365,N_15557,N_14852);
and U16366 (N_16366,N_14637,N_15780);
nand U16367 (N_16367,N_15798,N_15205);
nand U16368 (N_16368,N_15040,N_14635);
nor U16369 (N_16369,N_14501,N_15691);
nor U16370 (N_16370,N_15574,N_14476);
nand U16371 (N_16371,N_15113,N_14612);
nor U16372 (N_16372,N_15726,N_14045);
or U16373 (N_16373,N_14992,N_15902);
and U16374 (N_16374,N_14734,N_15522);
nand U16375 (N_16375,N_15353,N_15312);
and U16376 (N_16376,N_14199,N_15743);
nor U16377 (N_16377,N_14509,N_15321);
nand U16378 (N_16378,N_14391,N_15540);
nand U16379 (N_16379,N_14180,N_14726);
or U16380 (N_16380,N_14255,N_15428);
nor U16381 (N_16381,N_14305,N_15905);
and U16382 (N_16382,N_14233,N_14266);
and U16383 (N_16383,N_15085,N_15431);
or U16384 (N_16384,N_15754,N_14703);
or U16385 (N_16385,N_15098,N_14836);
and U16386 (N_16386,N_14118,N_15996);
and U16387 (N_16387,N_14596,N_15866);
and U16388 (N_16388,N_14627,N_15868);
nand U16389 (N_16389,N_15387,N_15372);
xnor U16390 (N_16390,N_15207,N_15432);
nand U16391 (N_16391,N_15835,N_14618);
or U16392 (N_16392,N_15232,N_15488);
or U16393 (N_16393,N_15222,N_14780);
and U16394 (N_16394,N_14303,N_15782);
nand U16395 (N_16395,N_14708,N_15659);
or U16396 (N_16396,N_14006,N_14282);
nand U16397 (N_16397,N_14197,N_14238);
or U16398 (N_16398,N_14786,N_15792);
nand U16399 (N_16399,N_15236,N_14175);
nand U16400 (N_16400,N_14106,N_15666);
or U16401 (N_16401,N_14137,N_14713);
nor U16402 (N_16402,N_15672,N_15765);
nor U16403 (N_16403,N_14546,N_14466);
nand U16404 (N_16404,N_15953,N_14120);
nand U16405 (N_16405,N_14896,N_15524);
nand U16406 (N_16406,N_14060,N_14932);
and U16407 (N_16407,N_15345,N_15459);
and U16408 (N_16408,N_15015,N_14550);
nand U16409 (N_16409,N_15787,N_14644);
and U16410 (N_16410,N_14144,N_15346);
nand U16411 (N_16411,N_15287,N_14017);
nand U16412 (N_16412,N_14744,N_15855);
and U16413 (N_16413,N_14632,N_15607);
nor U16414 (N_16414,N_14862,N_15092);
and U16415 (N_16415,N_14791,N_15191);
xnor U16416 (N_16416,N_15941,N_15497);
and U16417 (N_16417,N_14173,N_15219);
nor U16418 (N_16418,N_15807,N_14625);
or U16419 (N_16419,N_14221,N_15972);
and U16420 (N_16420,N_14647,N_15119);
nand U16421 (N_16421,N_15639,N_14382);
nand U16422 (N_16422,N_14845,N_14906);
nand U16423 (N_16423,N_14392,N_14236);
or U16424 (N_16424,N_15348,N_15491);
or U16425 (N_16425,N_14285,N_14973);
and U16426 (N_16426,N_15937,N_14979);
nor U16427 (N_16427,N_14809,N_15673);
nand U16428 (N_16428,N_14901,N_15775);
nand U16429 (N_16429,N_14442,N_15703);
or U16430 (N_16430,N_15892,N_15667);
nand U16431 (N_16431,N_14115,N_14057);
or U16432 (N_16432,N_15967,N_14484);
nor U16433 (N_16433,N_14652,N_15859);
and U16434 (N_16434,N_14772,N_15498);
or U16435 (N_16435,N_15116,N_15393);
and U16436 (N_16436,N_15450,N_14438);
and U16437 (N_16437,N_14952,N_15526);
xor U16438 (N_16438,N_14650,N_14986);
xnor U16439 (N_16439,N_14937,N_15099);
or U16440 (N_16440,N_15906,N_15723);
nand U16441 (N_16441,N_15741,N_15262);
xor U16442 (N_16442,N_14879,N_14425);
or U16443 (N_16443,N_14776,N_14547);
xor U16444 (N_16444,N_15537,N_15082);
nor U16445 (N_16445,N_15760,N_14128);
or U16446 (N_16446,N_15183,N_14567);
nand U16447 (N_16447,N_14782,N_14299);
nand U16448 (N_16448,N_15373,N_14833);
and U16449 (N_16449,N_14994,N_15118);
nor U16450 (N_16450,N_15550,N_14138);
or U16451 (N_16451,N_14692,N_15564);
nor U16452 (N_16452,N_15430,N_15783);
nor U16453 (N_16453,N_15109,N_14080);
or U16454 (N_16454,N_15576,N_15748);
or U16455 (N_16455,N_15083,N_14753);
and U16456 (N_16456,N_15086,N_15259);
or U16457 (N_16457,N_15555,N_15828);
nand U16458 (N_16458,N_14153,N_15961);
nor U16459 (N_16459,N_14227,N_15461);
nor U16460 (N_16460,N_15231,N_14341);
nor U16461 (N_16461,N_15415,N_14904);
and U16462 (N_16462,N_15606,N_14976);
nor U16463 (N_16463,N_15031,N_14784);
and U16464 (N_16464,N_15050,N_14020);
nor U16465 (N_16465,N_14499,N_15097);
or U16466 (N_16466,N_15962,N_15157);
nor U16467 (N_16467,N_15005,N_15628);
nand U16468 (N_16468,N_14419,N_14718);
nand U16469 (N_16469,N_14639,N_14167);
xnor U16470 (N_16470,N_14926,N_15617);
and U16471 (N_16471,N_15162,N_15277);
or U16472 (N_16472,N_15674,N_14781);
xor U16473 (N_16473,N_15002,N_15182);
or U16474 (N_16474,N_14394,N_15150);
and U16475 (N_16475,N_15605,N_14237);
or U16476 (N_16476,N_15694,N_14935);
and U16477 (N_16477,N_14384,N_15715);
and U16478 (N_16478,N_14688,N_15912);
and U16479 (N_16479,N_14939,N_15985);
or U16480 (N_16480,N_14838,N_15827);
nor U16481 (N_16481,N_15176,N_14424);
or U16482 (N_16482,N_15405,N_14676);
and U16483 (N_16483,N_15654,N_14046);
or U16484 (N_16484,N_14188,N_15944);
nand U16485 (N_16485,N_14555,N_14864);
nand U16486 (N_16486,N_14241,N_14699);
and U16487 (N_16487,N_14999,N_14367);
nor U16488 (N_16488,N_15969,N_15256);
and U16489 (N_16489,N_15877,N_14249);
nand U16490 (N_16490,N_14529,N_15896);
nor U16491 (N_16491,N_14131,N_14696);
xnor U16492 (N_16492,N_15292,N_14551);
and U16493 (N_16493,N_15115,N_14284);
xor U16494 (N_16494,N_14510,N_14250);
xnor U16495 (N_16495,N_15876,N_15752);
or U16496 (N_16496,N_14891,N_14214);
and U16497 (N_16497,N_15426,N_15745);
nand U16498 (N_16498,N_15621,N_15523);
nor U16499 (N_16499,N_14005,N_15845);
nor U16500 (N_16500,N_14008,N_14353);
or U16501 (N_16501,N_14661,N_14821);
nor U16502 (N_16502,N_14790,N_14787);
and U16503 (N_16503,N_14204,N_15390);
nand U16504 (N_16504,N_14828,N_15651);
nor U16505 (N_16505,N_15076,N_14467);
or U16506 (N_16506,N_14581,N_14252);
or U16507 (N_16507,N_15641,N_15449);
and U16508 (N_16508,N_14505,N_14082);
and U16509 (N_16509,N_14441,N_14881);
nor U16510 (N_16510,N_15913,N_14957);
xor U16511 (N_16511,N_15984,N_14497);
nor U16512 (N_16512,N_15590,N_15558);
nor U16513 (N_16513,N_14587,N_14463);
or U16514 (N_16514,N_14577,N_14877);
nor U16515 (N_16515,N_15661,N_14938);
nand U16516 (N_16516,N_15198,N_15057);
nand U16517 (N_16517,N_15288,N_15813);
xor U16518 (N_16518,N_15411,N_14092);
nor U16519 (N_16519,N_15916,N_15518);
nand U16520 (N_16520,N_15529,N_14435);
or U16521 (N_16521,N_15202,N_15239);
xnor U16522 (N_16522,N_15211,N_15593);
or U16523 (N_16523,N_15226,N_15758);
nor U16524 (N_16524,N_15151,N_15359);
nor U16525 (N_16525,N_14974,N_14922);
nor U16526 (N_16526,N_15768,N_15465);
nor U16527 (N_16527,N_15134,N_14094);
or U16528 (N_16528,N_15947,N_15772);
nor U16529 (N_16529,N_15382,N_14493);
and U16530 (N_16530,N_15600,N_14685);
xor U16531 (N_16531,N_14948,N_15552);
or U16532 (N_16532,N_14069,N_15511);
nand U16533 (N_16533,N_14693,N_15989);
nand U16534 (N_16534,N_15053,N_14190);
nor U16535 (N_16535,N_14855,N_15270);
and U16536 (N_16536,N_14260,N_14931);
xor U16537 (N_16537,N_15250,N_15532);
nor U16538 (N_16538,N_15403,N_14658);
nand U16539 (N_16539,N_14468,N_15110);
and U16540 (N_16540,N_15062,N_14149);
nor U16541 (N_16541,N_14923,N_15306);
and U16542 (N_16542,N_15165,N_14548);
nor U16543 (N_16543,N_15900,N_14208);
or U16544 (N_16544,N_14585,N_14829);
nor U16545 (N_16545,N_15588,N_14924);
or U16546 (N_16546,N_14422,N_14071);
and U16547 (N_16547,N_15619,N_15003);
nand U16548 (N_16548,N_14900,N_15462);
and U16549 (N_16549,N_15148,N_15883);
nand U16550 (N_16550,N_15895,N_14598);
or U16551 (N_16551,N_14858,N_15197);
and U16552 (N_16552,N_15433,N_15974);
and U16553 (N_16553,N_15893,N_15327);
nand U16554 (N_16554,N_14988,N_14943);
nand U16555 (N_16555,N_15485,N_14229);
nor U16556 (N_16556,N_15404,N_14489);
and U16557 (N_16557,N_14995,N_14009);
nor U16558 (N_16558,N_15368,N_15833);
nor U16559 (N_16559,N_14860,N_15370);
or U16560 (N_16560,N_14345,N_14670);
nor U16561 (N_16561,N_14705,N_15997);
and U16562 (N_16562,N_14186,N_15472);
xor U16563 (N_16563,N_14918,N_14155);
nor U16564 (N_16564,N_15490,N_14492);
nand U16565 (N_16565,N_14164,N_14091);
nand U16566 (N_16566,N_14657,N_15650);
and U16567 (N_16567,N_15520,N_14217);
and U16568 (N_16568,N_14626,N_15750);
and U16569 (N_16569,N_14815,N_14889);
or U16570 (N_16570,N_15837,N_14449);
nor U16571 (N_16571,N_15973,N_14767);
or U16572 (N_16572,N_15041,N_15736);
nor U16573 (N_16573,N_14328,N_15965);
or U16574 (N_16574,N_15903,N_15680);
nand U16575 (N_16575,N_14411,N_15313);
or U16576 (N_16576,N_14535,N_14032);
and U16577 (N_16577,N_14066,N_14522);
or U16578 (N_16578,N_15412,N_14448);
or U16579 (N_16579,N_15351,N_14873);
or U16580 (N_16580,N_14000,N_14007);
or U16581 (N_16581,N_14651,N_14101);
nor U16582 (N_16582,N_14145,N_15594);
or U16583 (N_16583,N_15000,N_15029);
nand U16584 (N_16584,N_15587,N_14569);
nand U16585 (N_16585,N_15548,N_14628);
and U16586 (N_16586,N_15846,N_14714);
nor U16587 (N_16587,N_14812,N_14084);
and U16588 (N_16588,N_14574,N_15023);
and U16589 (N_16589,N_14774,N_14601);
nand U16590 (N_16590,N_15867,N_15874);
nor U16591 (N_16591,N_14851,N_14320);
nand U16592 (N_16592,N_15897,N_14573);
nand U16593 (N_16593,N_15128,N_14818);
nor U16594 (N_16594,N_14894,N_15330);
nor U16595 (N_16595,N_15566,N_15677);
and U16596 (N_16596,N_14736,N_14364);
or U16597 (N_16597,N_15093,N_14758);
nor U16598 (N_16598,N_15635,N_15398);
nor U16599 (N_16599,N_14695,N_14251);
and U16600 (N_16600,N_14887,N_15720);
xor U16601 (N_16601,N_15943,N_14265);
nand U16602 (N_16602,N_14694,N_14025);
nor U16603 (N_16603,N_14775,N_14675);
or U16604 (N_16604,N_15771,N_15452);
nand U16605 (N_16605,N_14160,N_15125);
nand U16606 (N_16606,N_15457,N_15631);
nand U16607 (N_16607,N_14200,N_14749);
nor U16608 (N_16608,N_14064,N_15421);
nand U16609 (N_16609,N_15138,N_14010);
nor U16610 (N_16610,N_15458,N_15181);
or U16611 (N_16611,N_14872,N_14794);
and U16612 (N_16612,N_14421,N_14487);
nor U16613 (N_16613,N_14814,N_15931);
nand U16614 (N_16614,N_15646,N_14486);
or U16615 (N_16615,N_15890,N_14024);
nand U16616 (N_16616,N_15662,N_15999);
xnor U16617 (N_16617,N_15027,N_15928);
nand U16618 (N_16618,N_14480,N_14564);
nand U16619 (N_16619,N_14099,N_14645);
nand U16620 (N_16620,N_15318,N_15535);
nor U16621 (N_16621,N_14899,N_14352);
and U16622 (N_16622,N_15763,N_14324);
nand U16623 (N_16623,N_15510,N_15952);
or U16624 (N_16624,N_15940,N_14659);
xor U16625 (N_16625,N_15159,N_15143);
and U16626 (N_16626,N_14376,N_14426);
or U16627 (N_16627,N_14147,N_15721);
and U16628 (N_16628,N_15296,N_15879);
and U16629 (N_16629,N_15611,N_15033);
nor U16630 (N_16630,N_14459,N_15470);
and U16631 (N_16631,N_15696,N_15210);
xnor U16632 (N_16632,N_15901,N_14056);
xor U16633 (N_16633,N_15355,N_14156);
nor U16634 (N_16634,N_14090,N_14330);
nor U16635 (N_16635,N_15615,N_15589);
nand U16636 (N_16636,N_14245,N_14738);
nand U16637 (N_16637,N_15386,N_15443);
xnor U16638 (N_16638,N_15870,N_15248);
or U16639 (N_16639,N_14354,N_15881);
or U16640 (N_16640,N_14036,N_14469);
nor U16641 (N_16641,N_15501,N_15562);
nand U16642 (N_16642,N_14925,N_15489);
nor U16643 (N_16643,N_15257,N_14033);
and U16644 (N_16644,N_14553,N_15009);
or U16645 (N_16645,N_15284,N_15708);
nor U16646 (N_16646,N_14903,N_15013);
nor U16647 (N_16647,N_15808,N_15601);
nor U16648 (N_16648,N_14752,N_14315);
xnor U16649 (N_16649,N_14181,N_14826);
xor U16650 (N_16650,N_14413,N_15689);
nor U16651 (N_16651,N_14817,N_14378);
and U16652 (N_16652,N_15471,N_15979);
or U16653 (N_16653,N_14026,N_15749);
nand U16654 (N_16654,N_15328,N_15112);
and U16655 (N_16655,N_14847,N_14097);
or U16656 (N_16656,N_15418,N_14054);
nand U16657 (N_16657,N_14834,N_15429);
nand U16658 (N_16658,N_15586,N_15016);
and U16659 (N_16659,N_15209,N_15735);
or U16660 (N_16660,N_15025,N_15679);
and U16661 (N_16661,N_15395,N_14242);
and U16662 (N_16662,N_15454,N_15469);
nor U16663 (N_16663,N_15945,N_14162);
or U16664 (N_16664,N_14246,N_15195);
and U16665 (N_16665,N_14605,N_14527);
xor U16666 (N_16666,N_15122,N_14697);
and U16667 (N_16667,N_14018,N_14611);
nor U16668 (N_16668,N_15055,N_15990);
and U16669 (N_16669,N_14290,N_15744);
nand U16670 (N_16670,N_14636,N_15542);
or U16671 (N_16671,N_15424,N_15998);
and U16672 (N_16672,N_15067,N_14159);
nor U16673 (N_16673,N_14093,N_14415);
and U16674 (N_16674,N_14306,N_14318);
nor U16675 (N_16675,N_15266,N_14766);
or U16676 (N_16676,N_14523,N_14954);
or U16677 (N_16677,N_15258,N_14150);
xor U16678 (N_16678,N_14771,N_14220);
and U16679 (N_16679,N_14876,N_14086);
xor U16680 (N_16680,N_15699,N_15612);
and U16681 (N_16681,N_14457,N_15010);
nand U16682 (N_16682,N_14136,N_14969);
nor U16683 (N_16683,N_14124,N_14807);
and U16684 (N_16684,N_15208,N_15687);
xor U16685 (N_16685,N_14850,N_15043);
or U16686 (N_16686,N_15793,N_15899);
nand U16687 (N_16687,N_14728,N_14079);
nand U16688 (N_16688,N_14478,N_14998);
or U16689 (N_16689,N_15521,N_14865);
or U16690 (N_16690,N_14272,N_15801);
or U16691 (N_16691,N_15213,N_15241);
nand U16692 (N_16692,N_15955,N_14317);
nand U16693 (N_16693,N_15154,N_15761);
nor U16694 (N_16694,N_14712,N_15445);
and U16695 (N_16695,N_15762,N_14205);
and U16696 (N_16696,N_15531,N_14732);
nand U16697 (N_16697,N_15340,N_14154);
nand U16698 (N_16698,N_15991,N_15515);
xor U16699 (N_16699,N_15274,N_15120);
nand U16700 (N_16700,N_14526,N_15478);
and U16701 (N_16701,N_15096,N_15717);
nand U16702 (N_16702,N_14975,N_15212);
or U16703 (N_16703,N_15839,N_15819);
nor U16704 (N_16704,N_14508,N_14279);
or U16705 (N_16705,N_15622,N_15933);
nand U16706 (N_16706,N_14959,N_14933);
nor U16707 (N_16707,N_14163,N_14116);
or U16708 (N_16708,N_15218,N_14319);
or U16709 (N_16709,N_15803,N_14506);
xnor U16710 (N_16710,N_14460,N_15994);
nor U16711 (N_16711,N_14414,N_15982);
nand U16712 (N_16712,N_14946,N_14740);
or U16713 (N_16713,N_15397,N_14177);
nor U16714 (N_16714,N_14210,N_14806);
nor U16715 (N_16715,N_14624,N_14942);
or U16716 (N_16716,N_15822,N_15725);
nor U16717 (N_16717,N_15078,N_15583);
or U16718 (N_16718,N_14883,N_14515);
and U16719 (N_16719,N_15305,N_14770);
nand U16720 (N_16720,N_15409,N_15108);
or U16721 (N_16721,N_14912,N_14416);
nand U16722 (N_16722,N_14335,N_15858);
nor U16723 (N_16723,N_15942,N_14023);
and U16724 (N_16724,N_14653,N_15315);
nor U16725 (N_16725,N_15106,N_15142);
and U16726 (N_16726,N_14745,N_14930);
nor U16727 (N_16727,N_15035,N_14642);
or U16728 (N_16728,N_14235,N_15755);
nor U16729 (N_16729,N_14198,N_15121);
and U16730 (N_16730,N_15323,N_15388);
and U16731 (N_16731,N_15610,N_14096);
nand U16732 (N_16732,N_15326,N_15045);
xnor U16733 (N_16733,N_14951,N_15882);
and U16734 (N_16734,N_14055,N_15438);
nor U16735 (N_16735,N_14178,N_15620);
and U16736 (N_16736,N_14968,N_15131);
nor U16737 (N_16737,N_14640,N_14545);
nor U16738 (N_16738,N_14427,N_14050);
nor U16739 (N_16739,N_14398,N_15378);
nand U16740 (N_16740,N_15683,N_14127);
or U16741 (N_16741,N_15051,N_15530);
xnor U16742 (N_16742,N_15516,N_14077);
or U16743 (N_16743,N_14859,N_14846);
nand U16744 (N_16744,N_15260,N_15842);
nand U16745 (N_16745,N_14802,N_15880);
or U16746 (N_16746,N_15436,N_15228);
and U16747 (N_16747,N_15652,N_15643);
nand U16748 (N_16748,N_15830,N_15037);
or U16749 (N_16749,N_15950,N_15441);
nor U16750 (N_16750,N_15335,N_14110);
and U16751 (N_16751,N_15609,N_14291);
nand U16752 (N_16752,N_14157,N_14015);
and U16753 (N_16753,N_14880,N_14977);
xor U16754 (N_16754,N_14458,N_14857);
or U16755 (N_16755,N_14288,N_14552);
nand U16756 (N_16756,N_15496,N_14799);
nand U16757 (N_16757,N_15350,N_15957);
and U16758 (N_16758,N_15805,N_15756);
nor U16759 (N_16759,N_14400,N_14216);
or U16760 (N_16760,N_15242,N_15278);
nand U16761 (N_16761,N_14504,N_15167);
or U16762 (N_16762,N_15300,N_15477);
and U16763 (N_16763,N_14401,N_15591);
nor U16764 (N_16764,N_14984,N_15073);
nor U16765 (N_16765,N_15437,N_15420);
nor U16766 (N_16766,N_15152,N_15414);
nand U16767 (N_16767,N_14041,N_15080);
nor U16768 (N_16768,N_15225,N_14958);
or U16769 (N_16769,N_15847,N_15439);
and U16770 (N_16770,N_15977,N_15843);
and U16771 (N_16771,N_15243,N_14521);
nor U16772 (N_16772,N_15136,N_14481);
and U16773 (N_16773,N_14989,N_15493);
or U16774 (N_16774,N_14586,N_14132);
or U16775 (N_16775,N_14882,N_14662);
or U16776 (N_16776,N_15460,N_14087);
xor U16777 (N_16777,N_15014,N_14349);
nand U16778 (N_16778,N_14848,N_15665);
nor U16779 (N_16779,N_15722,N_15247);
nand U16780 (N_16780,N_15921,N_15809);
nor U16781 (N_16781,N_14294,N_15081);
nand U16782 (N_16782,N_15264,N_14059);
xor U16783 (N_16783,N_14037,N_14098);
nand U16784 (N_16784,N_14176,N_15713);
or U16785 (N_16785,N_14418,N_15271);
nor U16786 (N_16786,N_14408,N_14248);
nor U16787 (N_16787,N_14729,N_15199);
nor U16788 (N_16788,N_15132,N_14465);
nor U16789 (N_16789,N_15004,N_15316);
xor U16790 (N_16790,N_15354,N_14366);
and U16791 (N_16791,N_15026,N_14280);
or U16792 (N_16792,N_15337,N_14140);
nor U16793 (N_16793,N_15790,N_15019);
nor U16794 (N_16794,N_15304,N_15385);
nor U16795 (N_16795,N_15423,N_14472);
xnor U16796 (N_16796,N_14067,N_15831);
xnor U16797 (N_16797,N_14013,N_14905);
or U16798 (N_16798,N_14139,N_14372);
or U16799 (N_16799,N_15908,N_14554);
and U16800 (N_16800,N_14119,N_14841);
or U16801 (N_16801,N_14455,N_14491);
nand U16802 (N_16802,N_14395,N_14316);
nor U16803 (N_16803,N_14591,N_15682);
nor U16804 (N_16804,N_15818,N_14423);
and U16805 (N_16805,N_15030,N_15658);
nor U16806 (N_16806,N_14259,N_14172);
xor U16807 (N_16807,N_15178,N_14183);
or U16808 (N_16808,N_15624,N_14329);
nor U16809 (N_16809,N_15608,N_14304);
nor U16810 (N_16810,N_14532,N_14191);
xor U16811 (N_16811,N_15769,N_15863);
or U16812 (N_16812,N_14960,N_14701);
and U16813 (N_16813,N_15938,N_15632);
nor U16814 (N_16814,N_14690,N_15269);
nor U16815 (N_16815,N_14911,N_14374);
or U16816 (N_16816,N_15517,N_15613);
nand U16817 (N_16817,N_15546,N_14287);
nor U16818 (N_16818,N_14275,N_14133);
or U16819 (N_16819,N_15545,N_15506);
or U16820 (N_16820,N_15539,N_15046);
nand U16821 (N_16821,N_15105,N_15011);
nor U16822 (N_16822,N_14570,N_15294);
nor U16823 (N_16823,N_15090,N_14061);
or U16824 (N_16824,N_15144,N_15852);
xor U16825 (N_16825,N_14963,N_14654);
nor U16826 (N_16826,N_15779,N_14704);
and U16827 (N_16827,N_14583,N_15918);
or U16828 (N_16828,N_15629,N_14684);
nand U16829 (N_16829,N_15939,N_14539);
nand U16830 (N_16830,N_14383,N_15817);
or U16831 (N_16831,N_14461,N_14309);
and U16832 (N_16832,N_14040,N_14331);
nand U16833 (N_16833,N_15669,N_14733);
and U16834 (N_16834,N_14450,N_15848);
xnor U16835 (N_16835,N_15402,N_14669);
nand U16836 (N_16836,N_15844,N_15812);
or U16837 (N_16837,N_14663,N_15811);
nand U16838 (N_16838,N_14614,N_15153);
and U16839 (N_16839,N_14751,N_15644);
or U16840 (N_16840,N_15377,N_14543);
and U16841 (N_16841,N_14343,N_15276);
nand U16842 (N_16842,N_14038,N_14597);
nand U16843 (N_16843,N_14281,N_14276);
nor U16844 (N_16844,N_14825,N_14808);
or U16845 (N_16845,N_14483,N_14985);
nand U16846 (N_16846,N_15791,N_14253);
and U16847 (N_16847,N_15463,N_14536);
and U16848 (N_16848,N_15146,N_15664);
and U16849 (N_16849,N_14560,N_15101);
nor U16850 (N_16850,N_14107,N_14409);
nor U16851 (N_16851,N_15089,N_14301);
and U16852 (N_16852,N_14063,N_14616);
or U16853 (N_16853,N_14991,N_14870);
or U16854 (N_16854,N_15375,N_14723);
xnor U16855 (N_16855,N_15739,N_14258);
nand U16856 (N_16856,N_14725,N_15155);
and U16857 (N_16857,N_15728,N_14866);
nor U16858 (N_16858,N_15066,N_15416);
nand U16859 (N_16859,N_15865,N_15966);
nor U16860 (N_16860,N_14445,N_15718);
or U16861 (N_16861,N_15130,N_15872);
or U16862 (N_16862,N_15751,N_14602);
or U16863 (N_16863,N_14528,N_14804);
or U16864 (N_16864,N_15383,N_14209);
nor U16865 (N_16865,N_14385,N_15700);
nor U16866 (N_16866,N_15012,N_14513);
xor U16867 (N_16867,N_14607,N_14273);
nor U16868 (N_16868,N_15797,N_14861);
xnor U16869 (N_16869,N_14206,N_15983);
nand U16870 (N_16870,N_14379,N_14949);
xnor U16871 (N_16871,N_15727,N_14337);
and U16872 (N_16872,N_14085,N_15525);
and U16873 (N_16873,N_14339,N_14672);
and U16874 (N_16874,N_14187,N_14716);
and U16875 (N_16875,N_14996,N_15627);
or U16876 (N_16876,N_15686,N_14346);
or U16877 (N_16877,N_14321,N_14917);
and U16878 (N_16878,N_15596,N_14103);
and U16879 (N_16879,N_15864,N_14444);
nand U16880 (N_16880,N_15401,N_15060);
nor U16881 (N_16881,N_15740,N_15915);
nand U16882 (N_16882,N_14389,N_14201);
or U16883 (N_16883,N_15364,N_15995);
or U16884 (N_16884,N_15502,N_14058);
or U16885 (N_16885,N_14655,N_14074);
nor U16886 (N_16886,N_15911,N_15551);
and U16887 (N_16887,N_14965,N_15216);
and U16888 (N_16888,N_15473,N_15800);
nand U16889 (N_16889,N_15603,N_14709);
and U16890 (N_16890,N_15175,N_14778);
nand U16891 (N_16891,N_14620,N_14755);
nand U16892 (N_16892,N_15100,N_15795);
and U16893 (N_16893,N_15360,N_14078);
or U16894 (N_16894,N_15960,N_15413);
nand U16895 (N_16895,N_15124,N_15738);
nand U16896 (N_16896,N_14638,N_14247);
or U16897 (N_16897,N_14417,N_15255);
nor U16898 (N_16898,N_15935,N_15549);
or U16899 (N_16899,N_14910,N_15442);
or U16900 (N_16900,N_14566,N_14295);
and U16901 (N_16901,N_14446,N_15156);
nand U16902 (N_16902,N_14720,N_15440);
xnor U16903 (N_16903,N_15527,N_15069);
or U16904 (N_16904,N_14479,N_15064);
and U16905 (N_16905,N_14293,N_15695);
nor U16906 (N_16906,N_14746,N_15951);
nor U16907 (N_16907,N_14549,N_14439);
nand U16908 (N_16908,N_14307,N_14796);
and U16909 (N_16909,N_15929,N_15825);
nor U16910 (N_16910,N_14148,N_14195);
or U16911 (N_16911,N_15129,N_15399);
or U16912 (N_16912,N_14819,N_15071);
xor U16913 (N_16913,N_15024,N_14182);
nor U16914 (N_16914,N_15924,N_15179);
and U16915 (N_16915,N_15357,N_14520);
xor U16916 (N_16916,N_15380,N_14698);
and U16917 (N_16917,N_15180,N_15909);
and U16918 (N_16918,N_14429,N_14286);
or U16919 (N_16919,N_15126,N_14854);
and U16920 (N_16920,N_15410,N_15949);
nor U16921 (N_16921,N_15963,N_14405);
nand U16922 (N_16922,N_14202,N_14856);
or U16923 (N_16923,N_14920,N_14941);
and U16924 (N_16924,N_14666,N_15244);
or U16925 (N_16925,N_14595,N_15891);
nand U16926 (N_16926,N_15657,N_14559);
and U16927 (N_16927,N_15290,N_15836);
or U16928 (N_16928,N_14462,N_14065);
nor U16929 (N_16929,N_15322,N_15711);
or U16930 (N_16930,N_15253,N_15047);
nor U16931 (N_16931,N_15861,N_14396);
nor U16932 (N_16932,N_14104,N_14028);
and U16933 (N_16933,N_15417,N_15483);
nand U16934 (N_16934,N_15293,N_14525);
or U16935 (N_16935,N_15233,N_14673);
nand U16936 (N_16936,N_15265,N_15166);
xor U16937 (N_16937,N_15815,N_14019);
xnor U16938 (N_16938,N_14256,N_15685);
nand U16939 (N_16939,N_14004,N_15017);
or U16940 (N_16940,N_14477,N_15716);
nor U16941 (N_16941,N_15133,N_15204);
xor U16942 (N_16942,N_15577,N_14950);
nor U16943 (N_16943,N_14967,N_15455);
nand U16944 (N_16944,N_14839,N_15448);
xor U16945 (N_16945,N_15554,N_15816);
nor U16946 (N_16946,N_14283,N_15796);
or U16947 (N_16947,N_15789,N_15486);
xnor U16948 (N_16948,N_14842,N_14691);
nor U16949 (N_16949,N_15730,N_14369);
or U16950 (N_16950,N_14100,N_14312);
nand U16951 (N_16951,N_15747,N_14649);
nand U16952 (N_16952,N_14373,N_15203);
nand U16953 (N_16953,N_14130,N_14403);
and U16954 (N_16954,N_14109,N_14428);
nor U16955 (N_16955,N_15988,N_14095);
and U16956 (N_16956,N_15733,N_14944);
and U16957 (N_16957,N_14203,N_15668);
nor U16958 (N_16958,N_15343,N_15850);
nand U16959 (N_16959,N_15186,N_14853);
nor U16960 (N_16960,N_14184,N_14730);
nor U16961 (N_16961,N_14747,N_14043);
xor U16962 (N_16962,N_14757,N_15295);
nor U16963 (N_16963,N_14224,N_14892);
or U16964 (N_16964,N_15889,N_15456);
or U16965 (N_16965,N_14997,N_15170);
and U16966 (N_16966,N_15476,N_15556);
and U16967 (N_16967,N_15810,N_15776);
and U16968 (N_16968,N_15569,N_15503);
nand U16969 (N_16969,N_15633,N_14340);
and U16970 (N_16970,N_15584,N_14269);
and U16971 (N_16971,N_14430,N_14622);
nand U16972 (N_16972,N_14982,N_15707);
and U16973 (N_16973,N_14225,N_14928);
nand U16974 (N_16974,N_14721,N_15653);
nand U16975 (N_16975,N_14262,N_15425);
or U16976 (N_16976,N_15220,N_15948);
or U16977 (N_16977,N_15363,N_15770);
nor U16978 (N_16978,N_14022,N_15851);
xor U16979 (N_16979,N_14641,N_14921);
and U16980 (N_16980,N_15104,N_14240);
nor U16981 (N_16981,N_14268,N_15054);
and U16982 (N_16982,N_15171,N_14568);
and U16983 (N_16983,N_14511,N_14044);
and U16984 (N_16984,N_15509,N_14313);
and U16985 (N_16985,N_14750,N_15840);
nor U16986 (N_16986,N_14075,N_15185);
xor U16987 (N_16987,N_15021,N_15992);
or U16988 (N_16988,N_15215,N_15007);
and U16989 (N_16989,N_15075,N_15719);
and U16990 (N_16990,N_15930,N_15922);
and U16991 (N_16991,N_15147,N_15272);
or U16992 (N_16992,N_15671,N_15660);
or U16993 (N_16993,N_15039,N_14580);
and U16994 (N_16994,N_15595,N_14102);
nand U16995 (N_16995,N_14788,N_14151);
nor U16996 (N_16996,N_15926,N_15267);
or U16997 (N_16997,N_14052,N_14126);
or U16998 (N_16998,N_14114,N_15396);
nor U16999 (N_16999,N_14298,N_15332);
or U17000 (N_17000,N_14206,N_14662);
nor U17001 (N_17001,N_15496,N_15830);
nor U17002 (N_17002,N_15032,N_15577);
xnor U17003 (N_17003,N_14790,N_14640);
nand U17004 (N_17004,N_15128,N_14327);
nand U17005 (N_17005,N_15656,N_15067);
or U17006 (N_17006,N_14925,N_14322);
nor U17007 (N_17007,N_15757,N_15396);
or U17008 (N_17008,N_15342,N_14352);
or U17009 (N_17009,N_15066,N_15256);
and U17010 (N_17010,N_15631,N_14732);
and U17011 (N_17011,N_14400,N_15126);
and U17012 (N_17012,N_14478,N_15412);
and U17013 (N_17013,N_15631,N_15721);
nand U17014 (N_17014,N_14452,N_14691);
nand U17015 (N_17015,N_14235,N_15633);
and U17016 (N_17016,N_15605,N_15077);
nand U17017 (N_17017,N_14744,N_15604);
nor U17018 (N_17018,N_15101,N_15147);
and U17019 (N_17019,N_14482,N_14553);
and U17020 (N_17020,N_14684,N_14232);
and U17021 (N_17021,N_14046,N_15755);
nor U17022 (N_17022,N_14873,N_15596);
or U17023 (N_17023,N_15706,N_14705);
or U17024 (N_17024,N_14432,N_15005);
nor U17025 (N_17025,N_15632,N_15132);
nor U17026 (N_17026,N_14907,N_14340);
or U17027 (N_17027,N_14439,N_15886);
and U17028 (N_17028,N_14782,N_15459);
nand U17029 (N_17029,N_14419,N_15606);
nand U17030 (N_17030,N_15607,N_15289);
or U17031 (N_17031,N_14353,N_15579);
nand U17032 (N_17032,N_14078,N_15703);
and U17033 (N_17033,N_15717,N_15132);
and U17034 (N_17034,N_15824,N_15864);
nand U17035 (N_17035,N_14569,N_14963);
or U17036 (N_17036,N_15806,N_15598);
nand U17037 (N_17037,N_15086,N_15493);
or U17038 (N_17038,N_15869,N_15228);
nor U17039 (N_17039,N_15953,N_14494);
and U17040 (N_17040,N_14498,N_14176);
or U17041 (N_17041,N_15776,N_14562);
nand U17042 (N_17042,N_15561,N_15880);
or U17043 (N_17043,N_14147,N_14122);
or U17044 (N_17044,N_14955,N_15861);
nor U17045 (N_17045,N_14283,N_15281);
xnor U17046 (N_17046,N_15660,N_15341);
and U17047 (N_17047,N_14158,N_15580);
and U17048 (N_17048,N_14579,N_14456);
nand U17049 (N_17049,N_15584,N_15429);
nand U17050 (N_17050,N_14573,N_15973);
or U17051 (N_17051,N_14619,N_15246);
nor U17052 (N_17052,N_14346,N_14186);
or U17053 (N_17053,N_14023,N_14566);
and U17054 (N_17054,N_14381,N_14795);
or U17055 (N_17055,N_14760,N_15818);
and U17056 (N_17056,N_14542,N_14832);
and U17057 (N_17057,N_14907,N_15969);
and U17058 (N_17058,N_15419,N_14433);
nor U17059 (N_17059,N_14020,N_14886);
or U17060 (N_17060,N_14241,N_14763);
nor U17061 (N_17061,N_15449,N_15702);
and U17062 (N_17062,N_14296,N_15031);
or U17063 (N_17063,N_15590,N_15155);
and U17064 (N_17064,N_15102,N_15878);
and U17065 (N_17065,N_14692,N_14367);
nand U17066 (N_17066,N_15450,N_14428);
and U17067 (N_17067,N_15402,N_14877);
xnor U17068 (N_17068,N_15431,N_15303);
and U17069 (N_17069,N_14337,N_14090);
and U17070 (N_17070,N_14794,N_15533);
nor U17071 (N_17071,N_14887,N_15076);
or U17072 (N_17072,N_15505,N_15957);
and U17073 (N_17073,N_15668,N_14533);
nand U17074 (N_17074,N_14678,N_14797);
and U17075 (N_17075,N_15289,N_14021);
nand U17076 (N_17076,N_15269,N_15159);
and U17077 (N_17077,N_15973,N_14734);
and U17078 (N_17078,N_14822,N_15400);
xnor U17079 (N_17079,N_14388,N_14465);
nor U17080 (N_17080,N_15015,N_15455);
and U17081 (N_17081,N_14916,N_15636);
nand U17082 (N_17082,N_14548,N_14905);
or U17083 (N_17083,N_15223,N_15003);
nor U17084 (N_17084,N_14855,N_15386);
nand U17085 (N_17085,N_14632,N_15940);
and U17086 (N_17086,N_15982,N_14188);
or U17087 (N_17087,N_14278,N_14698);
nand U17088 (N_17088,N_15134,N_15678);
and U17089 (N_17089,N_15288,N_15583);
nand U17090 (N_17090,N_15080,N_15651);
nor U17091 (N_17091,N_15761,N_15669);
nor U17092 (N_17092,N_14852,N_14405);
or U17093 (N_17093,N_14114,N_15988);
and U17094 (N_17094,N_15888,N_15020);
nor U17095 (N_17095,N_14273,N_14173);
or U17096 (N_17096,N_15497,N_15835);
and U17097 (N_17097,N_14856,N_15815);
nand U17098 (N_17098,N_15658,N_15344);
xor U17099 (N_17099,N_15814,N_14075);
or U17100 (N_17100,N_15248,N_14651);
or U17101 (N_17101,N_15452,N_14993);
nor U17102 (N_17102,N_14857,N_15840);
nand U17103 (N_17103,N_15857,N_15570);
and U17104 (N_17104,N_14182,N_14326);
nor U17105 (N_17105,N_15548,N_15744);
nor U17106 (N_17106,N_14955,N_15151);
and U17107 (N_17107,N_15377,N_14264);
and U17108 (N_17108,N_15411,N_14844);
nand U17109 (N_17109,N_15013,N_14647);
or U17110 (N_17110,N_15956,N_14098);
or U17111 (N_17111,N_14143,N_15807);
or U17112 (N_17112,N_15863,N_14371);
nor U17113 (N_17113,N_14229,N_14829);
or U17114 (N_17114,N_15811,N_15187);
nand U17115 (N_17115,N_15918,N_14651);
nand U17116 (N_17116,N_15676,N_15095);
and U17117 (N_17117,N_15906,N_15102);
nor U17118 (N_17118,N_14811,N_15829);
xor U17119 (N_17119,N_14705,N_15376);
or U17120 (N_17120,N_15971,N_14270);
and U17121 (N_17121,N_14777,N_15663);
or U17122 (N_17122,N_14125,N_14162);
nand U17123 (N_17123,N_14657,N_15024);
or U17124 (N_17124,N_15964,N_15024);
nand U17125 (N_17125,N_14790,N_14823);
and U17126 (N_17126,N_15208,N_15374);
and U17127 (N_17127,N_15134,N_14311);
and U17128 (N_17128,N_15360,N_15382);
xnor U17129 (N_17129,N_15248,N_15031);
or U17130 (N_17130,N_14233,N_14416);
or U17131 (N_17131,N_14842,N_15739);
nand U17132 (N_17132,N_15962,N_15503);
nand U17133 (N_17133,N_15619,N_15809);
nor U17134 (N_17134,N_14614,N_15680);
nand U17135 (N_17135,N_14949,N_14134);
and U17136 (N_17136,N_14537,N_15920);
and U17137 (N_17137,N_14669,N_14469);
or U17138 (N_17138,N_14807,N_14157);
or U17139 (N_17139,N_15857,N_15804);
or U17140 (N_17140,N_15075,N_14188);
nand U17141 (N_17141,N_15078,N_15561);
nand U17142 (N_17142,N_15535,N_14262);
and U17143 (N_17143,N_15056,N_15819);
nor U17144 (N_17144,N_15001,N_15351);
nand U17145 (N_17145,N_14097,N_15905);
or U17146 (N_17146,N_15775,N_15137);
and U17147 (N_17147,N_15359,N_15702);
xor U17148 (N_17148,N_15131,N_14348);
nand U17149 (N_17149,N_15296,N_15121);
xor U17150 (N_17150,N_14559,N_14500);
nand U17151 (N_17151,N_15491,N_14075);
or U17152 (N_17152,N_15490,N_14702);
and U17153 (N_17153,N_15688,N_15792);
nand U17154 (N_17154,N_14353,N_14489);
nor U17155 (N_17155,N_15377,N_15773);
nor U17156 (N_17156,N_15363,N_15284);
or U17157 (N_17157,N_15303,N_15762);
or U17158 (N_17158,N_15135,N_14906);
or U17159 (N_17159,N_14286,N_14030);
or U17160 (N_17160,N_15301,N_15456);
and U17161 (N_17161,N_14884,N_15638);
and U17162 (N_17162,N_14517,N_14443);
nor U17163 (N_17163,N_15558,N_14531);
xnor U17164 (N_17164,N_14713,N_14551);
or U17165 (N_17165,N_14265,N_14673);
nor U17166 (N_17166,N_15689,N_14834);
nor U17167 (N_17167,N_14488,N_15173);
or U17168 (N_17168,N_15194,N_15969);
nand U17169 (N_17169,N_15134,N_14973);
xor U17170 (N_17170,N_14385,N_15093);
nor U17171 (N_17171,N_15987,N_15878);
nor U17172 (N_17172,N_14340,N_15991);
or U17173 (N_17173,N_14472,N_14054);
nor U17174 (N_17174,N_14956,N_14251);
nand U17175 (N_17175,N_14567,N_15229);
or U17176 (N_17176,N_15732,N_14946);
or U17177 (N_17177,N_14040,N_15487);
xnor U17178 (N_17178,N_15645,N_15364);
nand U17179 (N_17179,N_14291,N_14185);
nand U17180 (N_17180,N_15206,N_14632);
xnor U17181 (N_17181,N_14912,N_15487);
xor U17182 (N_17182,N_15415,N_15943);
xor U17183 (N_17183,N_15267,N_14268);
nor U17184 (N_17184,N_14594,N_14800);
or U17185 (N_17185,N_15054,N_14167);
or U17186 (N_17186,N_15787,N_14279);
and U17187 (N_17187,N_15176,N_14032);
and U17188 (N_17188,N_14083,N_14531);
or U17189 (N_17189,N_14976,N_14969);
nand U17190 (N_17190,N_14498,N_14537);
or U17191 (N_17191,N_14382,N_15992);
or U17192 (N_17192,N_14266,N_15303);
or U17193 (N_17193,N_14385,N_15470);
or U17194 (N_17194,N_15698,N_15840);
and U17195 (N_17195,N_14406,N_15031);
or U17196 (N_17196,N_14770,N_15183);
and U17197 (N_17197,N_14727,N_14997);
nand U17198 (N_17198,N_14158,N_15795);
or U17199 (N_17199,N_14817,N_14778);
nor U17200 (N_17200,N_15219,N_14521);
nand U17201 (N_17201,N_14500,N_15897);
or U17202 (N_17202,N_14343,N_14867);
nor U17203 (N_17203,N_14299,N_14563);
xnor U17204 (N_17204,N_14421,N_14370);
nor U17205 (N_17205,N_14991,N_15084);
nor U17206 (N_17206,N_14144,N_15742);
nand U17207 (N_17207,N_15049,N_14926);
nand U17208 (N_17208,N_15998,N_15848);
nor U17209 (N_17209,N_15100,N_15403);
nor U17210 (N_17210,N_14865,N_14770);
nor U17211 (N_17211,N_14287,N_14897);
xnor U17212 (N_17212,N_15655,N_14318);
nand U17213 (N_17213,N_15088,N_15854);
nand U17214 (N_17214,N_14628,N_15479);
and U17215 (N_17215,N_15067,N_15799);
nand U17216 (N_17216,N_15619,N_15232);
nor U17217 (N_17217,N_15984,N_15661);
nor U17218 (N_17218,N_15971,N_15184);
and U17219 (N_17219,N_14705,N_15024);
nor U17220 (N_17220,N_14486,N_15197);
or U17221 (N_17221,N_15096,N_14058);
nor U17222 (N_17222,N_15571,N_14077);
or U17223 (N_17223,N_15551,N_15559);
xnor U17224 (N_17224,N_14153,N_14958);
xnor U17225 (N_17225,N_14301,N_15970);
nand U17226 (N_17226,N_15240,N_14833);
xor U17227 (N_17227,N_14380,N_14744);
nor U17228 (N_17228,N_14738,N_15292);
xnor U17229 (N_17229,N_15118,N_15556);
nor U17230 (N_17230,N_15641,N_14512);
or U17231 (N_17231,N_15910,N_15122);
and U17232 (N_17232,N_14078,N_14666);
xnor U17233 (N_17233,N_14066,N_15422);
xnor U17234 (N_17234,N_15463,N_15980);
or U17235 (N_17235,N_15832,N_15917);
or U17236 (N_17236,N_14252,N_14869);
or U17237 (N_17237,N_15068,N_15039);
or U17238 (N_17238,N_15739,N_15547);
or U17239 (N_17239,N_14651,N_14671);
nor U17240 (N_17240,N_15864,N_14347);
nor U17241 (N_17241,N_14308,N_14645);
nand U17242 (N_17242,N_14567,N_15803);
or U17243 (N_17243,N_15254,N_14243);
or U17244 (N_17244,N_14801,N_14067);
nand U17245 (N_17245,N_14296,N_15975);
nor U17246 (N_17246,N_14374,N_14301);
nand U17247 (N_17247,N_14421,N_15657);
or U17248 (N_17248,N_15745,N_15247);
nor U17249 (N_17249,N_14581,N_15975);
or U17250 (N_17250,N_15226,N_15608);
xor U17251 (N_17251,N_15431,N_14004);
and U17252 (N_17252,N_15649,N_14052);
nor U17253 (N_17253,N_15534,N_15393);
nand U17254 (N_17254,N_14804,N_14378);
and U17255 (N_17255,N_14876,N_15730);
or U17256 (N_17256,N_14060,N_15403);
nor U17257 (N_17257,N_15207,N_14090);
or U17258 (N_17258,N_15233,N_15992);
or U17259 (N_17259,N_14417,N_15985);
nor U17260 (N_17260,N_15160,N_14801);
and U17261 (N_17261,N_15644,N_15371);
nand U17262 (N_17262,N_15490,N_14663);
or U17263 (N_17263,N_14342,N_14649);
and U17264 (N_17264,N_14496,N_15796);
and U17265 (N_17265,N_14384,N_15316);
xnor U17266 (N_17266,N_14937,N_14351);
and U17267 (N_17267,N_14508,N_14193);
nor U17268 (N_17268,N_15512,N_14767);
and U17269 (N_17269,N_14532,N_14750);
or U17270 (N_17270,N_14640,N_15986);
or U17271 (N_17271,N_15951,N_14817);
nor U17272 (N_17272,N_15481,N_15619);
nand U17273 (N_17273,N_14246,N_14662);
nand U17274 (N_17274,N_15190,N_14269);
nand U17275 (N_17275,N_15598,N_15764);
nor U17276 (N_17276,N_14475,N_15880);
or U17277 (N_17277,N_15418,N_14618);
nand U17278 (N_17278,N_15045,N_15398);
or U17279 (N_17279,N_14205,N_14931);
or U17280 (N_17280,N_15830,N_14089);
nor U17281 (N_17281,N_14513,N_14419);
xnor U17282 (N_17282,N_15277,N_14635);
nand U17283 (N_17283,N_15824,N_15595);
nor U17284 (N_17284,N_15087,N_15710);
nor U17285 (N_17285,N_14394,N_14277);
nand U17286 (N_17286,N_15939,N_14816);
nand U17287 (N_17287,N_15235,N_14612);
and U17288 (N_17288,N_15939,N_14362);
and U17289 (N_17289,N_15900,N_14827);
or U17290 (N_17290,N_15703,N_14237);
and U17291 (N_17291,N_14561,N_14069);
and U17292 (N_17292,N_14392,N_15484);
or U17293 (N_17293,N_15466,N_14628);
and U17294 (N_17294,N_14227,N_14119);
nor U17295 (N_17295,N_15963,N_15585);
xnor U17296 (N_17296,N_15381,N_15204);
nand U17297 (N_17297,N_15756,N_14584);
or U17298 (N_17298,N_15656,N_14334);
and U17299 (N_17299,N_15131,N_15948);
xor U17300 (N_17300,N_14053,N_14537);
or U17301 (N_17301,N_15874,N_15169);
xnor U17302 (N_17302,N_14372,N_15365);
nand U17303 (N_17303,N_14287,N_15121);
and U17304 (N_17304,N_15787,N_15349);
and U17305 (N_17305,N_15581,N_14675);
and U17306 (N_17306,N_15323,N_14404);
nor U17307 (N_17307,N_14774,N_15464);
and U17308 (N_17308,N_15383,N_14321);
xnor U17309 (N_17309,N_14391,N_15058);
and U17310 (N_17310,N_15200,N_15749);
xnor U17311 (N_17311,N_14311,N_15548);
and U17312 (N_17312,N_15087,N_15084);
nand U17313 (N_17313,N_15315,N_15376);
nand U17314 (N_17314,N_15009,N_15573);
and U17315 (N_17315,N_15407,N_14796);
or U17316 (N_17316,N_15783,N_14430);
nor U17317 (N_17317,N_14507,N_15286);
and U17318 (N_17318,N_14372,N_15680);
nor U17319 (N_17319,N_14026,N_14935);
or U17320 (N_17320,N_15815,N_15069);
nand U17321 (N_17321,N_15212,N_15673);
xor U17322 (N_17322,N_14883,N_15543);
nor U17323 (N_17323,N_15208,N_15591);
nand U17324 (N_17324,N_15833,N_15401);
or U17325 (N_17325,N_15975,N_15724);
nand U17326 (N_17326,N_15136,N_14208);
or U17327 (N_17327,N_14608,N_14741);
nor U17328 (N_17328,N_15274,N_15776);
nor U17329 (N_17329,N_14743,N_14813);
xor U17330 (N_17330,N_14483,N_15348);
and U17331 (N_17331,N_14043,N_15423);
and U17332 (N_17332,N_14538,N_15821);
and U17333 (N_17333,N_14549,N_14179);
nand U17334 (N_17334,N_14087,N_15981);
xor U17335 (N_17335,N_15020,N_14765);
nor U17336 (N_17336,N_15738,N_14687);
nand U17337 (N_17337,N_14157,N_15584);
xor U17338 (N_17338,N_15247,N_14867);
or U17339 (N_17339,N_15371,N_15333);
nor U17340 (N_17340,N_14173,N_14427);
nor U17341 (N_17341,N_15705,N_14205);
xor U17342 (N_17342,N_15629,N_15364);
and U17343 (N_17343,N_15881,N_15075);
or U17344 (N_17344,N_14237,N_14397);
or U17345 (N_17345,N_15123,N_14901);
and U17346 (N_17346,N_14615,N_15612);
and U17347 (N_17347,N_14368,N_15367);
or U17348 (N_17348,N_14330,N_14590);
nor U17349 (N_17349,N_15207,N_14093);
and U17350 (N_17350,N_14782,N_14331);
nor U17351 (N_17351,N_14443,N_15508);
and U17352 (N_17352,N_14974,N_14962);
nor U17353 (N_17353,N_15400,N_15623);
xor U17354 (N_17354,N_15407,N_15020);
nand U17355 (N_17355,N_15395,N_14650);
nand U17356 (N_17356,N_15265,N_14795);
nand U17357 (N_17357,N_14682,N_14017);
nor U17358 (N_17358,N_15563,N_15035);
xnor U17359 (N_17359,N_15129,N_15935);
nand U17360 (N_17360,N_14650,N_15265);
nor U17361 (N_17361,N_15360,N_15260);
nor U17362 (N_17362,N_14752,N_14521);
nand U17363 (N_17363,N_14106,N_15367);
nor U17364 (N_17364,N_15073,N_14308);
and U17365 (N_17365,N_14771,N_14200);
nand U17366 (N_17366,N_14769,N_15080);
or U17367 (N_17367,N_14075,N_14421);
nand U17368 (N_17368,N_15389,N_14671);
or U17369 (N_17369,N_15248,N_14342);
and U17370 (N_17370,N_14171,N_14474);
xnor U17371 (N_17371,N_14198,N_14514);
or U17372 (N_17372,N_15298,N_15955);
and U17373 (N_17373,N_14543,N_15063);
and U17374 (N_17374,N_15881,N_15271);
nor U17375 (N_17375,N_15904,N_15744);
or U17376 (N_17376,N_15621,N_15646);
and U17377 (N_17377,N_14413,N_14212);
or U17378 (N_17378,N_14977,N_14249);
and U17379 (N_17379,N_14250,N_14376);
nand U17380 (N_17380,N_15988,N_15241);
and U17381 (N_17381,N_14378,N_14459);
or U17382 (N_17382,N_14216,N_14222);
and U17383 (N_17383,N_15441,N_14629);
nand U17384 (N_17384,N_14595,N_14714);
or U17385 (N_17385,N_14602,N_15392);
nand U17386 (N_17386,N_15956,N_15990);
or U17387 (N_17387,N_14674,N_15181);
nor U17388 (N_17388,N_14257,N_14261);
xor U17389 (N_17389,N_14529,N_14791);
and U17390 (N_17390,N_15797,N_15674);
and U17391 (N_17391,N_15799,N_14767);
nor U17392 (N_17392,N_15740,N_15751);
and U17393 (N_17393,N_14213,N_15216);
or U17394 (N_17394,N_15043,N_14962);
nand U17395 (N_17395,N_14108,N_15439);
nor U17396 (N_17396,N_14645,N_15802);
nor U17397 (N_17397,N_14612,N_14169);
nor U17398 (N_17398,N_14352,N_15307);
nand U17399 (N_17399,N_14913,N_15474);
or U17400 (N_17400,N_15250,N_14323);
nor U17401 (N_17401,N_15920,N_14562);
or U17402 (N_17402,N_14498,N_15417);
nand U17403 (N_17403,N_15404,N_15761);
or U17404 (N_17404,N_14731,N_15888);
and U17405 (N_17405,N_15679,N_14389);
nor U17406 (N_17406,N_14236,N_14174);
nor U17407 (N_17407,N_14627,N_14021);
or U17408 (N_17408,N_15739,N_15897);
nand U17409 (N_17409,N_15442,N_14093);
and U17410 (N_17410,N_14143,N_15375);
and U17411 (N_17411,N_14822,N_15969);
and U17412 (N_17412,N_15343,N_14873);
xnor U17413 (N_17413,N_14294,N_14653);
or U17414 (N_17414,N_14542,N_14739);
nand U17415 (N_17415,N_15206,N_14697);
and U17416 (N_17416,N_14006,N_15422);
and U17417 (N_17417,N_14935,N_14991);
nand U17418 (N_17418,N_15510,N_14982);
or U17419 (N_17419,N_15058,N_14320);
nor U17420 (N_17420,N_14339,N_15136);
nor U17421 (N_17421,N_15751,N_15358);
xnor U17422 (N_17422,N_14084,N_14566);
or U17423 (N_17423,N_15381,N_14177);
or U17424 (N_17424,N_15359,N_15945);
nor U17425 (N_17425,N_15288,N_14321);
or U17426 (N_17426,N_15434,N_14810);
or U17427 (N_17427,N_14676,N_14301);
nand U17428 (N_17428,N_15208,N_15013);
or U17429 (N_17429,N_14956,N_14199);
xor U17430 (N_17430,N_15073,N_15883);
nor U17431 (N_17431,N_15892,N_14612);
nor U17432 (N_17432,N_14876,N_14087);
and U17433 (N_17433,N_14588,N_14680);
and U17434 (N_17434,N_14893,N_15094);
and U17435 (N_17435,N_14543,N_14221);
or U17436 (N_17436,N_14094,N_15659);
or U17437 (N_17437,N_15268,N_15831);
nand U17438 (N_17438,N_15551,N_14951);
nand U17439 (N_17439,N_14493,N_14514);
nor U17440 (N_17440,N_14009,N_14790);
nor U17441 (N_17441,N_14495,N_14585);
nor U17442 (N_17442,N_14263,N_15198);
nand U17443 (N_17443,N_15037,N_15531);
and U17444 (N_17444,N_14921,N_15075);
nor U17445 (N_17445,N_14479,N_15465);
and U17446 (N_17446,N_15302,N_15764);
xnor U17447 (N_17447,N_15542,N_14610);
nor U17448 (N_17448,N_15547,N_15603);
xnor U17449 (N_17449,N_15831,N_15978);
nor U17450 (N_17450,N_14201,N_14035);
or U17451 (N_17451,N_14168,N_14738);
nand U17452 (N_17452,N_14288,N_15863);
nor U17453 (N_17453,N_15992,N_15186);
and U17454 (N_17454,N_14704,N_15850);
nand U17455 (N_17455,N_15974,N_14723);
and U17456 (N_17456,N_14857,N_14996);
nor U17457 (N_17457,N_14516,N_15665);
nand U17458 (N_17458,N_14709,N_15388);
or U17459 (N_17459,N_14607,N_14505);
and U17460 (N_17460,N_14821,N_14925);
nor U17461 (N_17461,N_15980,N_14599);
and U17462 (N_17462,N_14977,N_14969);
nor U17463 (N_17463,N_14914,N_15716);
or U17464 (N_17464,N_14457,N_14517);
or U17465 (N_17465,N_14362,N_14819);
nand U17466 (N_17466,N_14232,N_14212);
nor U17467 (N_17467,N_14691,N_14181);
nor U17468 (N_17468,N_14319,N_15604);
and U17469 (N_17469,N_15901,N_14165);
nor U17470 (N_17470,N_15036,N_14151);
nand U17471 (N_17471,N_14481,N_15106);
and U17472 (N_17472,N_14418,N_14124);
or U17473 (N_17473,N_14688,N_15031);
xnor U17474 (N_17474,N_15841,N_14311);
and U17475 (N_17475,N_15291,N_15410);
or U17476 (N_17476,N_15926,N_14412);
and U17477 (N_17477,N_14640,N_14866);
nand U17478 (N_17478,N_14008,N_14834);
xor U17479 (N_17479,N_15516,N_15665);
or U17480 (N_17480,N_15111,N_14044);
xor U17481 (N_17481,N_14096,N_14899);
nor U17482 (N_17482,N_15962,N_15208);
and U17483 (N_17483,N_14596,N_15012);
nor U17484 (N_17484,N_15140,N_14278);
nand U17485 (N_17485,N_15786,N_15751);
xor U17486 (N_17486,N_15144,N_14389);
nand U17487 (N_17487,N_14831,N_14256);
nand U17488 (N_17488,N_14669,N_14618);
nor U17489 (N_17489,N_15281,N_14462);
nor U17490 (N_17490,N_15110,N_15436);
and U17491 (N_17491,N_14916,N_15882);
nor U17492 (N_17492,N_15689,N_14251);
or U17493 (N_17493,N_15513,N_15255);
xor U17494 (N_17494,N_15744,N_14620);
or U17495 (N_17495,N_15679,N_14253);
and U17496 (N_17496,N_15918,N_15776);
or U17497 (N_17497,N_14731,N_14750);
nand U17498 (N_17498,N_14130,N_14428);
xor U17499 (N_17499,N_14994,N_15286);
and U17500 (N_17500,N_15128,N_15856);
and U17501 (N_17501,N_15272,N_15711);
and U17502 (N_17502,N_14968,N_15685);
or U17503 (N_17503,N_14646,N_15983);
nand U17504 (N_17504,N_15527,N_14815);
and U17505 (N_17505,N_15305,N_14488);
nand U17506 (N_17506,N_14864,N_15346);
xnor U17507 (N_17507,N_15197,N_14926);
or U17508 (N_17508,N_15800,N_15357);
nand U17509 (N_17509,N_15764,N_15668);
and U17510 (N_17510,N_15650,N_15214);
nand U17511 (N_17511,N_14241,N_15795);
or U17512 (N_17512,N_14345,N_15814);
and U17513 (N_17513,N_14676,N_15349);
or U17514 (N_17514,N_14451,N_14586);
and U17515 (N_17515,N_15867,N_15651);
and U17516 (N_17516,N_15897,N_14468);
or U17517 (N_17517,N_15537,N_15996);
and U17518 (N_17518,N_15489,N_14756);
nand U17519 (N_17519,N_15751,N_14661);
or U17520 (N_17520,N_14667,N_14993);
and U17521 (N_17521,N_15715,N_15132);
or U17522 (N_17522,N_14801,N_14501);
nand U17523 (N_17523,N_14219,N_14490);
or U17524 (N_17524,N_14657,N_15472);
or U17525 (N_17525,N_15596,N_14038);
nor U17526 (N_17526,N_15202,N_15091);
and U17527 (N_17527,N_14715,N_14778);
xor U17528 (N_17528,N_14413,N_15918);
and U17529 (N_17529,N_15057,N_14496);
xor U17530 (N_17530,N_14069,N_15162);
nand U17531 (N_17531,N_14523,N_14829);
and U17532 (N_17532,N_15973,N_15959);
nand U17533 (N_17533,N_14863,N_15598);
nand U17534 (N_17534,N_15963,N_14300);
and U17535 (N_17535,N_14587,N_14056);
nand U17536 (N_17536,N_14394,N_14373);
and U17537 (N_17537,N_15780,N_14840);
and U17538 (N_17538,N_14990,N_15061);
or U17539 (N_17539,N_14307,N_15025);
or U17540 (N_17540,N_15776,N_14038);
nor U17541 (N_17541,N_15545,N_14120);
nand U17542 (N_17542,N_15824,N_15144);
and U17543 (N_17543,N_14623,N_15369);
nor U17544 (N_17544,N_14384,N_15042);
nand U17545 (N_17545,N_14190,N_15668);
or U17546 (N_17546,N_14809,N_15927);
and U17547 (N_17547,N_14318,N_14048);
or U17548 (N_17548,N_14021,N_15819);
and U17549 (N_17549,N_15917,N_14357);
nand U17550 (N_17550,N_14024,N_15082);
nor U17551 (N_17551,N_14163,N_14751);
nor U17552 (N_17552,N_15937,N_15502);
or U17553 (N_17553,N_15657,N_14207);
nand U17554 (N_17554,N_14918,N_14929);
or U17555 (N_17555,N_14472,N_15143);
nand U17556 (N_17556,N_15224,N_14640);
or U17557 (N_17557,N_14905,N_15487);
and U17558 (N_17558,N_14420,N_14570);
or U17559 (N_17559,N_15210,N_15105);
nor U17560 (N_17560,N_14658,N_14026);
nor U17561 (N_17561,N_14027,N_15684);
nor U17562 (N_17562,N_14654,N_15941);
nand U17563 (N_17563,N_14600,N_14173);
or U17564 (N_17564,N_15855,N_14654);
or U17565 (N_17565,N_15021,N_14017);
and U17566 (N_17566,N_14531,N_14021);
and U17567 (N_17567,N_15589,N_15171);
nor U17568 (N_17568,N_15116,N_15459);
and U17569 (N_17569,N_14757,N_14892);
or U17570 (N_17570,N_14221,N_14961);
and U17571 (N_17571,N_14678,N_15802);
nand U17572 (N_17572,N_14699,N_14382);
nand U17573 (N_17573,N_15908,N_14388);
or U17574 (N_17574,N_15835,N_14785);
nor U17575 (N_17575,N_14325,N_15862);
nand U17576 (N_17576,N_15413,N_15920);
nand U17577 (N_17577,N_14809,N_15354);
and U17578 (N_17578,N_14843,N_15563);
or U17579 (N_17579,N_15552,N_15036);
xnor U17580 (N_17580,N_15860,N_14044);
or U17581 (N_17581,N_14961,N_15607);
nor U17582 (N_17582,N_14640,N_14574);
and U17583 (N_17583,N_15285,N_15305);
and U17584 (N_17584,N_15732,N_15553);
nand U17585 (N_17585,N_14243,N_15774);
or U17586 (N_17586,N_14313,N_15931);
nand U17587 (N_17587,N_14010,N_14487);
xor U17588 (N_17588,N_15198,N_15729);
nor U17589 (N_17589,N_14469,N_15641);
nand U17590 (N_17590,N_14885,N_14413);
or U17591 (N_17591,N_15377,N_15689);
nor U17592 (N_17592,N_14037,N_14735);
or U17593 (N_17593,N_14803,N_15730);
nand U17594 (N_17594,N_14187,N_14490);
and U17595 (N_17595,N_15842,N_14758);
and U17596 (N_17596,N_14928,N_15552);
and U17597 (N_17597,N_15483,N_14778);
or U17598 (N_17598,N_14266,N_15833);
nor U17599 (N_17599,N_14162,N_15485);
nor U17600 (N_17600,N_15080,N_14672);
nor U17601 (N_17601,N_15513,N_14728);
or U17602 (N_17602,N_14128,N_14513);
and U17603 (N_17603,N_15232,N_15196);
xor U17604 (N_17604,N_15282,N_14819);
and U17605 (N_17605,N_14834,N_14869);
xnor U17606 (N_17606,N_15363,N_15473);
and U17607 (N_17607,N_15920,N_14333);
xnor U17608 (N_17608,N_14276,N_14397);
nand U17609 (N_17609,N_15244,N_15449);
nand U17610 (N_17610,N_14656,N_15228);
or U17611 (N_17611,N_14597,N_15449);
xor U17612 (N_17612,N_15598,N_15340);
and U17613 (N_17613,N_15521,N_14698);
and U17614 (N_17614,N_14140,N_15485);
or U17615 (N_17615,N_14959,N_15234);
xor U17616 (N_17616,N_15354,N_15281);
nor U17617 (N_17617,N_15019,N_14128);
or U17618 (N_17618,N_14554,N_14698);
nand U17619 (N_17619,N_14113,N_15662);
and U17620 (N_17620,N_15988,N_14917);
and U17621 (N_17621,N_14595,N_14887);
nor U17622 (N_17622,N_15496,N_14845);
nor U17623 (N_17623,N_15024,N_14902);
xor U17624 (N_17624,N_15315,N_14225);
nand U17625 (N_17625,N_14528,N_14489);
nor U17626 (N_17626,N_14526,N_14853);
and U17627 (N_17627,N_14059,N_14505);
nand U17628 (N_17628,N_15858,N_15792);
and U17629 (N_17629,N_14413,N_14117);
xor U17630 (N_17630,N_15357,N_14627);
xnor U17631 (N_17631,N_15870,N_14430);
nand U17632 (N_17632,N_15105,N_15774);
nor U17633 (N_17633,N_14043,N_15729);
nor U17634 (N_17634,N_15978,N_14157);
and U17635 (N_17635,N_15973,N_14642);
nand U17636 (N_17636,N_14975,N_14996);
nand U17637 (N_17637,N_14713,N_15614);
nand U17638 (N_17638,N_14789,N_15854);
or U17639 (N_17639,N_14249,N_14379);
and U17640 (N_17640,N_15173,N_15466);
nor U17641 (N_17641,N_15849,N_14980);
nand U17642 (N_17642,N_14607,N_15309);
and U17643 (N_17643,N_15682,N_15335);
or U17644 (N_17644,N_15677,N_14955);
and U17645 (N_17645,N_14864,N_14999);
and U17646 (N_17646,N_15336,N_15779);
or U17647 (N_17647,N_14070,N_14253);
or U17648 (N_17648,N_14010,N_15649);
or U17649 (N_17649,N_15310,N_14631);
nor U17650 (N_17650,N_15342,N_15663);
or U17651 (N_17651,N_15474,N_14482);
nor U17652 (N_17652,N_15922,N_15536);
or U17653 (N_17653,N_14601,N_15308);
nand U17654 (N_17654,N_14660,N_15027);
or U17655 (N_17655,N_15585,N_15652);
xor U17656 (N_17656,N_15163,N_15984);
and U17657 (N_17657,N_15824,N_14679);
nand U17658 (N_17658,N_14859,N_14185);
or U17659 (N_17659,N_15193,N_14604);
and U17660 (N_17660,N_14150,N_15657);
nand U17661 (N_17661,N_15216,N_14421);
and U17662 (N_17662,N_15184,N_15160);
nand U17663 (N_17663,N_14870,N_14645);
nand U17664 (N_17664,N_14514,N_14640);
and U17665 (N_17665,N_15559,N_15554);
nand U17666 (N_17666,N_15589,N_15064);
nor U17667 (N_17667,N_14470,N_14141);
or U17668 (N_17668,N_14065,N_15413);
nor U17669 (N_17669,N_15807,N_14789);
or U17670 (N_17670,N_14203,N_14513);
and U17671 (N_17671,N_15921,N_14525);
nand U17672 (N_17672,N_15458,N_15844);
and U17673 (N_17673,N_15929,N_15464);
or U17674 (N_17674,N_15545,N_14002);
nand U17675 (N_17675,N_14680,N_15171);
nand U17676 (N_17676,N_14904,N_14814);
nor U17677 (N_17677,N_15076,N_14872);
nand U17678 (N_17678,N_14593,N_14216);
and U17679 (N_17679,N_15730,N_15870);
and U17680 (N_17680,N_14577,N_15316);
or U17681 (N_17681,N_14092,N_14144);
nor U17682 (N_17682,N_15912,N_14302);
or U17683 (N_17683,N_14854,N_15611);
and U17684 (N_17684,N_15331,N_15090);
or U17685 (N_17685,N_15290,N_14477);
and U17686 (N_17686,N_14584,N_15415);
or U17687 (N_17687,N_14844,N_15342);
nor U17688 (N_17688,N_15379,N_15841);
nor U17689 (N_17689,N_14092,N_14213);
nor U17690 (N_17690,N_14126,N_15560);
or U17691 (N_17691,N_14982,N_14479);
nor U17692 (N_17692,N_15133,N_15023);
and U17693 (N_17693,N_14033,N_15556);
nor U17694 (N_17694,N_15394,N_15416);
nand U17695 (N_17695,N_14505,N_14523);
or U17696 (N_17696,N_14258,N_14893);
or U17697 (N_17697,N_15713,N_14428);
or U17698 (N_17698,N_15912,N_15957);
nor U17699 (N_17699,N_15928,N_14058);
xnor U17700 (N_17700,N_14886,N_14810);
nand U17701 (N_17701,N_15414,N_15517);
nand U17702 (N_17702,N_14869,N_14790);
nor U17703 (N_17703,N_15352,N_14532);
nand U17704 (N_17704,N_14237,N_14417);
nor U17705 (N_17705,N_15073,N_15550);
nand U17706 (N_17706,N_15475,N_15849);
nor U17707 (N_17707,N_15576,N_14697);
nor U17708 (N_17708,N_15064,N_14488);
or U17709 (N_17709,N_14657,N_14053);
nor U17710 (N_17710,N_15102,N_14046);
xor U17711 (N_17711,N_15318,N_14834);
nand U17712 (N_17712,N_14017,N_15434);
nand U17713 (N_17713,N_14067,N_14582);
or U17714 (N_17714,N_14888,N_14846);
or U17715 (N_17715,N_15087,N_14273);
nand U17716 (N_17716,N_15653,N_15677);
or U17717 (N_17717,N_14926,N_14887);
or U17718 (N_17718,N_14762,N_14689);
and U17719 (N_17719,N_14908,N_15671);
or U17720 (N_17720,N_14311,N_15286);
nor U17721 (N_17721,N_15022,N_14308);
or U17722 (N_17722,N_15974,N_14712);
nand U17723 (N_17723,N_14918,N_15046);
nor U17724 (N_17724,N_15746,N_14953);
or U17725 (N_17725,N_15749,N_15723);
or U17726 (N_17726,N_14015,N_15929);
and U17727 (N_17727,N_14946,N_14596);
or U17728 (N_17728,N_14660,N_14982);
nor U17729 (N_17729,N_15379,N_15659);
and U17730 (N_17730,N_15468,N_14841);
nor U17731 (N_17731,N_15358,N_14086);
and U17732 (N_17732,N_14796,N_15280);
or U17733 (N_17733,N_15670,N_14489);
or U17734 (N_17734,N_15836,N_14709);
or U17735 (N_17735,N_15337,N_14535);
or U17736 (N_17736,N_14590,N_14576);
nand U17737 (N_17737,N_14962,N_15187);
and U17738 (N_17738,N_15360,N_14326);
nand U17739 (N_17739,N_15593,N_14348);
or U17740 (N_17740,N_14308,N_14740);
or U17741 (N_17741,N_15808,N_15205);
nor U17742 (N_17742,N_15655,N_14731);
and U17743 (N_17743,N_15130,N_15449);
and U17744 (N_17744,N_14908,N_15795);
or U17745 (N_17745,N_14669,N_15566);
nor U17746 (N_17746,N_15660,N_15106);
xnor U17747 (N_17747,N_15258,N_15597);
or U17748 (N_17748,N_14449,N_14045);
nor U17749 (N_17749,N_15177,N_14228);
nor U17750 (N_17750,N_14756,N_15599);
or U17751 (N_17751,N_15977,N_15663);
nor U17752 (N_17752,N_14431,N_14077);
nand U17753 (N_17753,N_15500,N_15895);
nor U17754 (N_17754,N_15578,N_14849);
and U17755 (N_17755,N_15984,N_15394);
nor U17756 (N_17756,N_14691,N_15265);
or U17757 (N_17757,N_14563,N_14306);
nand U17758 (N_17758,N_14139,N_15678);
and U17759 (N_17759,N_15857,N_15309);
nor U17760 (N_17760,N_15372,N_14653);
and U17761 (N_17761,N_15924,N_15066);
or U17762 (N_17762,N_14445,N_15611);
or U17763 (N_17763,N_14704,N_15199);
and U17764 (N_17764,N_15723,N_14633);
and U17765 (N_17765,N_15822,N_15260);
and U17766 (N_17766,N_14456,N_14306);
or U17767 (N_17767,N_15959,N_15900);
nor U17768 (N_17768,N_15821,N_14914);
nand U17769 (N_17769,N_15344,N_15926);
nor U17770 (N_17770,N_15624,N_15006);
xnor U17771 (N_17771,N_14987,N_15623);
and U17772 (N_17772,N_15988,N_14418);
or U17773 (N_17773,N_14161,N_15869);
or U17774 (N_17774,N_14351,N_14058);
and U17775 (N_17775,N_15637,N_15776);
nor U17776 (N_17776,N_14003,N_15445);
and U17777 (N_17777,N_14454,N_14886);
nor U17778 (N_17778,N_15101,N_14367);
and U17779 (N_17779,N_14680,N_15181);
xnor U17780 (N_17780,N_15627,N_15215);
and U17781 (N_17781,N_14576,N_15965);
nand U17782 (N_17782,N_15938,N_15141);
and U17783 (N_17783,N_15210,N_15253);
or U17784 (N_17784,N_15864,N_14748);
and U17785 (N_17785,N_14326,N_14299);
xor U17786 (N_17786,N_14250,N_14303);
and U17787 (N_17787,N_14907,N_14159);
nor U17788 (N_17788,N_15990,N_15553);
nand U17789 (N_17789,N_15551,N_15436);
nor U17790 (N_17790,N_14006,N_14895);
nor U17791 (N_17791,N_15282,N_14605);
nor U17792 (N_17792,N_14458,N_14420);
nor U17793 (N_17793,N_15605,N_14773);
and U17794 (N_17794,N_14959,N_15922);
and U17795 (N_17795,N_14944,N_14114);
and U17796 (N_17796,N_14427,N_15723);
and U17797 (N_17797,N_14472,N_15872);
nor U17798 (N_17798,N_14898,N_14291);
or U17799 (N_17799,N_15189,N_15076);
nor U17800 (N_17800,N_14744,N_14402);
nor U17801 (N_17801,N_15080,N_15535);
nand U17802 (N_17802,N_15341,N_14936);
or U17803 (N_17803,N_15240,N_15320);
and U17804 (N_17804,N_15840,N_14563);
xor U17805 (N_17805,N_15695,N_15184);
and U17806 (N_17806,N_15449,N_14315);
nand U17807 (N_17807,N_15035,N_15433);
and U17808 (N_17808,N_14645,N_14742);
nor U17809 (N_17809,N_14565,N_15187);
nand U17810 (N_17810,N_15269,N_14896);
nand U17811 (N_17811,N_15157,N_15708);
nand U17812 (N_17812,N_15469,N_14010);
nand U17813 (N_17813,N_15643,N_14079);
nand U17814 (N_17814,N_15589,N_14618);
xnor U17815 (N_17815,N_15548,N_14533);
nor U17816 (N_17816,N_15017,N_14225);
or U17817 (N_17817,N_14961,N_14003);
and U17818 (N_17818,N_15218,N_14518);
or U17819 (N_17819,N_15728,N_14780);
nor U17820 (N_17820,N_14742,N_14776);
and U17821 (N_17821,N_15486,N_14924);
and U17822 (N_17822,N_15593,N_15751);
xnor U17823 (N_17823,N_15817,N_14475);
or U17824 (N_17824,N_15327,N_15746);
xnor U17825 (N_17825,N_15703,N_14788);
and U17826 (N_17826,N_15114,N_15634);
or U17827 (N_17827,N_15665,N_14151);
and U17828 (N_17828,N_15805,N_14827);
nand U17829 (N_17829,N_14497,N_14543);
nor U17830 (N_17830,N_14691,N_14151);
and U17831 (N_17831,N_14095,N_14024);
or U17832 (N_17832,N_15469,N_14524);
nor U17833 (N_17833,N_15723,N_14789);
and U17834 (N_17834,N_14685,N_15656);
nand U17835 (N_17835,N_15460,N_14897);
or U17836 (N_17836,N_15813,N_15623);
nand U17837 (N_17837,N_14016,N_15971);
or U17838 (N_17838,N_15229,N_15647);
nand U17839 (N_17839,N_14699,N_15553);
nor U17840 (N_17840,N_15323,N_15345);
xor U17841 (N_17841,N_14586,N_15612);
xnor U17842 (N_17842,N_14531,N_14098);
nor U17843 (N_17843,N_15447,N_15829);
and U17844 (N_17844,N_14574,N_15312);
nand U17845 (N_17845,N_14592,N_15486);
nand U17846 (N_17846,N_15837,N_14852);
nand U17847 (N_17847,N_15075,N_15194);
or U17848 (N_17848,N_14811,N_14940);
nand U17849 (N_17849,N_14201,N_14134);
nor U17850 (N_17850,N_14294,N_14208);
nand U17851 (N_17851,N_15260,N_15063);
and U17852 (N_17852,N_14989,N_14134);
or U17853 (N_17853,N_14193,N_14791);
and U17854 (N_17854,N_15908,N_15585);
nor U17855 (N_17855,N_15944,N_14881);
and U17856 (N_17856,N_15576,N_15886);
and U17857 (N_17857,N_14158,N_14004);
nand U17858 (N_17858,N_15863,N_15412);
or U17859 (N_17859,N_14070,N_14532);
or U17860 (N_17860,N_15282,N_15408);
or U17861 (N_17861,N_14238,N_14168);
xor U17862 (N_17862,N_14824,N_14547);
or U17863 (N_17863,N_15334,N_14921);
or U17864 (N_17864,N_14844,N_15048);
and U17865 (N_17865,N_15321,N_14012);
nand U17866 (N_17866,N_15590,N_15982);
nor U17867 (N_17867,N_15348,N_15649);
and U17868 (N_17868,N_14550,N_14091);
and U17869 (N_17869,N_14032,N_14340);
and U17870 (N_17870,N_15149,N_14291);
or U17871 (N_17871,N_14834,N_14050);
and U17872 (N_17872,N_14705,N_14415);
or U17873 (N_17873,N_15784,N_15462);
nor U17874 (N_17874,N_15103,N_15496);
nand U17875 (N_17875,N_15240,N_14877);
nand U17876 (N_17876,N_14176,N_14378);
or U17877 (N_17877,N_14064,N_14861);
nand U17878 (N_17878,N_15070,N_14129);
nor U17879 (N_17879,N_15501,N_15057);
nand U17880 (N_17880,N_14720,N_15627);
and U17881 (N_17881,N_15929,N_14522);
or U17882 (N_17882,N_14518,N_14544);
or U17883 (N_17883,N_14272,N_14313);
or U17884 (N_17884,N_14034,N_15658);
or U17885 (N_17885,N_14862,N_15824);
nor U17886 (N_17886,N_14855,N_15550);
nor U17887 (N_17887,N_14371,N_14501);
and U17888 (N_17888,N_14208,N_14073);
or U17889 (N_17889,N_14418,N_15383);
xnor U17890 (N_17890,N_14484,N_14791);
and U17891 (N_17891,N_15115,N_14795);
and U17892 (N_17892,N_14864,N_15567);
or U17893 (N_17893,N_14206,N_14223);
or U17894 (N_17894,N_15823,N_15158);
nor U17895 (N_17895,N_14436,N_14472);
or U17896 (N_17896,N_15676,N_15379);
or U17897 (N_17897,N_15360,N_14725);
nand U17898 (N_17898,N_14801,N_15456);
and U17899 (N_17899,N_15779,N_14458);
nand U17900 (N_17900,N_14863,N_15251);
or U17901 (N_17901,N_15495,N_15176);
nor U17902 (N_17902,N_14567,N_14059);
nor U17903 (N_17903,N_15183,N_15489);
xor U17904 (N_17904,N_14348,N_15098);
nor U17905 (N_17905,N_15815,N_15249);
nand U17906 (N_17906,N_15378,N_14086);
or U17907 (N_17907,N_15626,N_14267);
nor U17908 (N_17908,N_15175,N_14680);
nor U17909 (N_17909,N_14203,N_15722);
or U17910 (N_17910,N_15273,N_14009);
xnor U17911 (N_17911,N_15488,N_15571);
nand U17912 (N_17912,N_15657,N_15975);
nor U17913 (N_17913,N_15833,N_14924);
and U17914 (N_17914,N_14313,N_15493);
nand U17915 (N_17915,N_14882,N_14579);
nor U17916 (N_17916,N_14408,N_14123);
nor U17917 (N_17917,N_15332,N_15642);
nand U17918 (N_17918,N_14331,N_15252);
nor U17919 (N_17919,N_14706,N_14132);
or U17920 (N_17920,N_15586,N_14499);
or U17921 (N_17921,N_14162,N_14255);
nand U17922 (N_17922,N_14347,N_14341);
and U17923 (N_17923,N_14489,N_14837);
nor U17924 (N_17924,N_15087,N_15883);
nor U17925 (N_17925,N_15383,N_15988);
and U17926 (N_17926,N_15911,N_14405);
and U17927 (N_17927,N_14000,N_15363);
and U17928 (N_17928,N_15542,N_15867);
or U17929 (N_17929,N_15354,N_15440);
nor U17930 (N_17930,N_14973,N_15373);
xnor U17931 (N_17931,N_15397,N_14435);
xnor U17932 (N_17932,N_15302,N_15491);
nand U17933 (N_17933,N_15674,N_14198);
or U17934 (N_17934,N_15840,N_15794);
nor U17935 (N_17935,N_15386,N_15288);
xnor U17936 (N_17936,N_14556,N_15761);
nand U17937 (N_17937,N_15364,N_14470);
nor U17938 (N_17938,N_15396,N_15574);
and U17939 (N_17939,N_15472,N_15420);
or U17940 (N_17940,N_14293,N_15136);
and U17941 (N_17941,N_15809,N_15354);
or U17942 (N_17942,N_15373,N_15040);
and U17943 (N_17943,N_15927,N_14214);
or U17944 (N_17944,N_14747,N_15574);
nor U17945 (N_17945,N_15312,N_15738);
xor U17946 (N_17946,N_14710,N_14930);
nor U17947 (N_17947,N_14773,N_15726);
nor U17948 (N_17948,N_15928,N_15484);
nor U17949 (N_17949,N_15747,N_14683);
nand U17950 (N_17950,N_14680,N_14058);
and U17951 (N_17951,N_15813,N_14885);
nor U17952 (N_17952,N_15801,N_14911);
nor U17953 (N_17953,N_15311,N_15224);
nor U17954 (N_17954,N_14732,N_15248);
xor U17955 (N_17955,N_15860,N_15433);
and U17956 (N_17956,N_14065,N_15414);
and U17957 (N_17957,N_14195,N_15674);
and U17958 (N_17958,N_15707,N_14637);
or U17959 (N_17959,N_15052,N_15678);
or U17960 (N_17960,N_14352,N_14302);
and U17961 (N_17961,N_15818,N_14000);
or U17962 (N_17962,N_14112,N_15922);
nor U17963 (N_17963,N_15558,N_14679);
nor U17964 (N_17964,N_15531,N_14821);
and U17965 (N_17965,N_14947,N_15664);
and U17966 (N_17966,N_15175,N_15834);
nor U17967 (N_17967,N_14499,N_14921);
and U17968 (N_17968,N_14105,N_15170);
and U17969 (N_17969,N_14756,N_14487);
or U17970 (N_17970,N_15946,N_15047);
nor U17971 (N_17971,N_15062,N_14882);
nand U17972 (N_17972,N_14068,N_14588);
or U17973 (N_17973,N_15032,N_15443);
or U17974 (N_17974,N_15679,N_15361);
or U17975 (N_17975,N_14195,N_14521);
nor U17976 (N_17976,N_15925,N_14922);
nor U17977 (N_17977,N_14919,N_14269);
and U17978 (N_17978,N_15081,N_15975);
nor U17979 (N_17979,N_14879,N_15522);
xor U17980 (N_17980,N_15304,N_15846);
or U17981 (N_17981,N_15201,N_14180);
xor U17982 (N_17982,N_15014,N_14144);
or U17983 (N_17983,N_15779,N_15569);
xnor U17984 (N_17984,N_15081,N_14603);
or U17985 (N_17985,N_14160,N_14620);
nor U17986 (N_17986,N_15663,N_15873);
or U17987 (N_17987,N_15767,N_14272);
and U17988 (N_17988,N_15442,N_14024);
or U17989 (N_17989,N_14082,N_14575);
nor U17990 (N_17990,N_14527,N_15848);
and U17991 (N_17991,N_14459,N_15767);
and U17992 (N_17992,N_15034,N_15740);
xor U17993 (N_17993,N_14192,N_14311);
or U17994 (N_17994,N_15311,N_14082);
and U17995 (N_17995,N_15732,N_15315);
nor U17996 (N_17996,N_14944,N_14099);
xor U17997 (N_17997,N_14569,N_14362);
nor U17998 (N_17998,N_14581,N_15100);
nor U17999 (N_17999,N_15888,N_15458);
xor U18000 (N_18000,N_16004,N_17155);
nor U18001 (N_18001,N_17369,N_16276);
nor U18002 (N_18002,N_16355,N_16128);
nor U18003 (N_18003,N_16149,N_17136);
or U18004 (N_18004,N_17187,N_17833);
or U18005 (N_18005,N_17065,N_17826);
and U18006 (N_18006,N_17810,N_16471);
and U18007 (N_18007,N_17754,N_17710);
xor U18008 (N_18008,N_16227,N_17540);
or U18009 (N_18009,N_16479,N_17918);
nand U18010 (N_18010,N_17657,N_16602);
xnor U18011 (N_18011,N_16343,N_16719);
and U18012 (N_18012,N_17956,N_16409);
and U18013 (N_18013,N_17153,N_16302);
and U18014 (N_18014,N_16356,N_16671);
and U18015 (N_18015,N_17167,N_17024);
or U18016 (N_18016,N_16436,N_17890);
nor U18017 (N_18017,N_16920,N_17950);
and U18018 (N_18018,N_17711,N_17888);
nand U18019 (N_18019,N_17862,N_16491);
xor U18020 (N_18020,N_17249,N_16451);
and U18021 (N_18021,N_17329,N_17993);
nor U18022 (N_18022,N_16617,N_16572);
or U18023 (N_18023,N_17893,N_16812);
nor U18024 (N_18024,N_17855,N_17449);
and U18025 (N_18025,N_17482,N_16999);
and U18026 (N_18026,N_16929,N_17177);
nand U18027 (N_18027,N_17995,N_16291);
or U18028 (N_18028,N_17870,N_17849);
xor U18029 (N_18029,N_16477,N_16133);
nor U18030 (N_18030,N_16412,N_17234);
or U18031 (N_18031,N_16712,N_16434);
nor U18032 (N_18032,N_16124,N_16605);
nand U18033 (N_18033,N_17029,N_16126);
nand U18034 (N_18034,N_16410,N_17007);
nand U18035 (N_18035,N_16567,N_16936);
nand U18036 (N_18036,N_17878,N_16918);
nand U18037 (N_18037,N_17083,N_16281);
xnor U18038 (N_18038,N_17420,N_17931);
and U18039 (N_18039,N_16688,N_16545);
xor U18040 (N_18040,N_16352,N_16770);
or U18041 (N_18041,N_17905,N_17084);
nand U18042 (N_18042,N_17182,N_16831);
and U18043 (N_18043,N_17027,N_17533);
xnor U18044 (N_18044,N_16098,N_17543);
nand U18045 (N_18045,N_16317,N_17267);
or U18046 (N_18046,N_16954,N_17583);
nand U18047 (N_18047,N_17159,N_16984);
nor U18048 (N_18048,N_16253,N_16199);
and U18049 (N_18049,N_17464,N_17097);
nand U18050 (N_18050,N_16201,N_16060);
and U18051 (N_18051,N_16368,N_16297);
xor U18052 (N_18052,N_17410,N_16686);
nand U18053 (N_18053,N_16312,N_16123);
or U18054 (N_18054,N_16768,N_17506);
and U18055 (N_18055,N_16767,N_17842);
or U18056 (N_18056,N_17627,N_17118);
nor U18057 (N_18057,N_17185,N_16233);
nor U18058 (N_18058,N_17593,N_17953);
nor U18059 (N_18059,N_16463,N_16131);
or U18060 (N_18060,N_16484,N_16868);
nand U18061 (N_18061,N_17815,N_16928);
nand U18062 (N_18062,N_17792,N_17689);
or U18063 (N_18063,N_16525,N_17474);
nor U18064 (N_18064,N_17417,N_16906);
nand U18065 (N_18065,N_16594,N_17020);
xor U18066 (N_18066,N_17203,N_16910);
or U18067 (N_18067,N_17477,N_16092);
nor U18068 (N_18068,N_17618,N_16109);
and U18069 (N_18069,N_16922,N_16592);
nor U18070 (N_18070,N_16483,N_17515);
and U18071 (N_18071,N_16962,N_17491);
or U18072 (N_18072,N_17392,N_17762);
nor U18073 (N_18073,N_16258,N_17478);
or U18074 (N_18074,N_16859,N_16216);
nor U18075 (N_18075,N_17693,N_16304);
or U18076 (N_18076,N_17812,N_17850);
nand U18077 (N_18077,N_17753,N_17158);
or U18078 (N_18078,N_16667,N_16170);
and U18079 (N_18079,N_16673,N_16137);
nand U18080 (N_18080,N_16626,N_16951);
xor U18081 (N_18081,N_17735,N_16727);
nor U18082 (N_18082,N_16053,N_17493);
xnor U18083 (N_18083,N_16518,N_17816);
or U18084 (N_18084,N_17462,N_17713);
and U18085 (N_18085,N_16827,N_16158);
and U18086 (N_18086,N_17977,N_17082);
xor U18087 (N_18087,N_17052,N_16474);
nand U18088 (N_18088,N_16566,N_16457);
or U18089 (N_18089,N_16786,N_17384);
or U18090 (N_18090,N_16705,N_16959);
or U18091 (N_18091,N_17922,N_16584);
and U18092 (N_18092,N_16665,N_16238);
and U18093 (N_18093,N_17759,N_16653);
nor U18094 (N_18094,N_17643,N_17039);
or U18095 (N_18095,N_17312,N_17916);
nor U18096 (N_18096,N_17419,N_17990);
or U18097 (N_18097,N_16998,N_16424);
or U18098 (N_18098,N_17373,N_16174);
nand U18099 (N_18099,N_16492,N_17952);
nand U18100 (N_18100,N_17614,N_17201);
nand U18101 (N_18101,N_17205,N_17736);
or U18102 (N_18102,N_16988,N_16037);
nand U18103 (N_18103,N_17925,N_17740);
and U18104 (N_18104,N_17585,N_16386);
nor U18105 (N_18105,N_17926,N_17824);
and U18106 (N_18106,N_17920,N_17220);
and U18107 (N_18107,N_16777,N_17265);
xor U18108 (N_18108,N_17380,N_17929);
or U18109 (N_18109,N_16274,N_16269);
and U18110 (N_18110,N_16441,N_17231);
or U18111 (N_18111,N_17194,N_17649);
xnor U18112 (N_18112,N_16361,N_16250);
nand U18113 (N_18113,N_16257,N_17786);
nand U18114 (N_18114,N_16075,N_17761);
xnor U18115 (N_18115,N_16469,N_16862);
nor U18116 (N_18116,N_17733,N_17268);
and U18117 (N_18117,N_17741,N_17914);
and U18118 (N_18118,N_16817,N_17058);
nor U18119 (N_18119,N_16325,N_16314);
nand U18120 (N_18120,N_16609,N_17398);
or U18121 (N_18121,N_16919,N_17919);
nand U18122 (N_18122,N_17121,N_16108);
nor U18123 (N_18123,N_16077,N_17688);
or U18124 (N_18124,N_17257,N_17322);
or U18125 (N_18125,N_16578,N_16366);
nand U18126 (N_18126,N_17588,N_16025);
or U18127 (N_18127,N_17061,N_16947);
or U18128 (N_18128,N_17293,N_16877);
and U18129 (N_18129,N_17228,N_17610);
nand U18130 (N_18130,N_17938,N_17747);
or U18131 (N_18131,N_16086,N_16809);
nand U18132 (N_18132,N_16308,N_16007);
and U18133 (N_18133,N_16526,N_16198);
or U18134 (N_18134,N_16121,N_17756);
and U18135 (N_18135,N_16421,N_17031);
xor U18136 (N_18136,N_16327,N_16520);
nor U18137 (N_18137,N_16587,N_16563);
or U18138 (N_18138,N_17250,N_17484);
xnor U18139 (N_18139,N_16209,N_16689);
nor U18140 (N_18140,N_16618,N_17361);
or U18141 (N_18141,N_17105,N_16989);
and U18142 (N_18142,N_16094,N_17086);
xnor U18143 (N_18143,N_17366,N_16042);
and U18144 (N_18144,N_16925,N_17615);
nor U18145 (N_18145,N_17758,N_16502);
nor U18146 (N_18146,N_16582,N_16608);
nor U18147 (N_18147,N_17828,N_16071);
and U18148 (N_18148,N_17433,N_17143);
nand U18149 (N_18149,N_16405,N_16960);
nor U18150 (N_18150,N_17655,N_16437);
or U18151 (N_18151,N_16600,N_17139);
nand U18152 (N_18152,N_17067,N_17056);
nand U18153 (N_18153,N_17080,N_16443);
and U18154 (N_18154,N_16277,N_17854);
and U18155 (N_18155,N_17161,N_16548);
and U18156 (N_18156,N_16850,N_17718);
nor U18157 (N_18157,N_17880,N_17604);
and U18158 (N_18158,N_16569,N_17690);
and U18159 (N_18159,N_17912,N_16334);
and U18160 (N_18160,N_16338,N_17276);
and U18161 (N_18161,N_17004,N_17012);
or U18162 (N_18162,N_16958,N_16800);
nand U18163 (N_18163,N_17275,N_17383);
xor U18164 (N_18164,N_17064,N_16535);
or U18165 (N_18165,N_17387,N_16478);
nand U18166 (N_18166,N_16461,N_16691);
xnor U18167 (N_18167,N_17856,N_16397);
or U18168 (N_18168,N_16139,N_17566);
xor U18169 (N_18169,N_16011,N_16547);
or U18170 (N_18170,N_17882,N_17575);
and U18171 (N_18171,N_17994,N_16829);
xor U18172 (N_18172,N_16555,N_17089);
nand U18173 (N_18173,N_16177,N_16083);
and U18174 (N_18174,N_16903,N_16728);
nand U18175 (N_18175,N_17793,N_16486);
nand U18176 (N_18176,N_16481,N_16814);
and U18177 (N_18177,N_16035,N_17364);
nand U18178 (N_18178,N_16046,N_16305);
and U18179 (N_18179,N_17242,N_16666);
nand U18180 (N_18180,N_17094,N_16008);
and U18181 (N_18181,N_16684,N_17138);
nor U18182 (N_18182,N_16242,N_17126);
xor U18183 (N_18183,N_17490,N_16280);
nand U18184 (N_18184,N_17318,N_16839);
nand U18185 (N_18185,N_17670,N_17987);
nand U18186 (N_18186,N_16031,N_16351);
or U18187 (N_18187,N_17451,N_16232);
and U18188 (N_18188,N_17869,N_16400);
nor U18189 (N_18189,N_17653,N_16805);
or U18190 (N_18190,N_17054,N_16625);
and U18191 (N_18191,N_16278,N_16841);
nor U18192 (N_18192,N_17986,N_16023);
or U18193 (N_18193,N_16911,N_17306);
xnor U18194 (N_18194,N_17134,N_17283);
and U18195 (N_18195,N_16119,N_16869);
nor U18196 (N_18196,N_16726,N_16021);
or U18197 (N_18197,N_17144,N_17011);
and U18198 (N_18198,N_16235,N_16265);
and U18199 (N_18199,N_17014,N_17394);
and U18200 (N_18200,N_17487,N_17367);
nand U18201 (N_18201,N_17211,N_17715);
nor U18202 (N_18202,N_17519,N_16210);
and U18203 (N_18203,N_17598,N_16788);
nor U18204 (N_18204,N_17001,N_17036);
and U18205 (N_18205,N_17866,N_17556);
and U18206 (N_18206,N_16465,N_17620);
or U18207 (N_18207,N_16980,N_17915);
xnor U18208 (N_18208,N_16524,N_16058);
or U18209 (N_18209,N_16480,N_17692);
nand U18210 (N_18210,N_17349,N_17208);
nor U18211 (N_18211,N_17040,N_17189);
and U18212 (N_18212,N_17281,N_17179);
xnor U18213 (N_18213,N_16044,N_16082);
nand U18214 (N_18214,N_17513,N_16136);
and U18215 (N_18215,N_17418,N_17055);
or U18216 (N_18216,N_16428,N_17791);
nor U18217 (N_18217,N_16835,N_16791);
nor U18218 (N_18218,N_17965,N_16896);
nand U18219 (N_18219,N_16715,N_17483);
or U18220 (N_18220,N_17647,N_16837);
or U18221 (N_18221,N_17215,N_16380);
or U18222 (N_18222,N_17512,N_17796);
or U18223 (N_18223,N_16144,N_16818);
and U18224 (N_18224,N_16010,N_17353);
and U18225 (N_18225,N_17101,N_16738);
and U18226 (N_18226,N_17823,N_17725);
or U18227 (N_18227,N_16806,N_17835);
nand U18228 (N_18228,N_17272,N_16912);
or U18229 (N_18229,N_17169,N_16861);
and U18230 (N_18230,N_16532,N_17386);
or U18231 (N_18231,N_17579,N_16493);
and U18232 (N_18232,N_16141,N_17949);
or U18233 (N_18233,N_17877,N_16435);
nor U18234 (N_18234,N_16203,N_17181);
and U18235 (N_18235,N_16773,N_17681);
nor U18236 (N_18236,N_16760,N_17184);
and U18237 (N_18237,N_17340,N_17156);
and U18238 (N_18238,N_17180,N_16716);
nor U18239 (N_18239,N_17534,N_16544);
nand U18240 (N_18240,N_16654,N_16255);
nor U18241 (N_18241,N_17437,N_17957);
and U18242 (N_18242,N_16677,N_17291);
and U18243 (N_18243,N_17175,N_16458);
and U18244 (N_18244,N_16781,N_17428);
or U18245 (N_18245,N_16374,N_17269);
nand U18246 (N_18246,N_16268,N_16372);
nand U18247 (N_18247,N_17675,N_16658);
nand U18248 (N_18248,N_17038,N_16482);
nand U18249 (N_18249,N_16485,N_17172);
and U18250 (N_18250,N_17465,N_16442);
or U18251 (N_18251,N_16192,N_17171);
xor U18252 (N_18252,N_17974,N_16403);
and U18253 (N_18253,N_16766,N_16935);
or U18254 (N_18254,N_16634,N_16891);
nor U18255 (N_18255,N_17438,N_16117);
nand U18256 (N_18256,N_16615,N_17308);
nand U18257 (N_18257,N_16650,N_17382);
and U18258 (N_18258,N_16236,N_16224);
and U18259 (N_18259,N_17385,N_17699);
nor U18260 (N_18260,N_17109,N_17219);
nor U18261 (N_18261,N_16455,N_16759);
and U18262 (N_18262,N_17648,N_17897);
nor U18263 (N_18263,N_17261,N_17602);
nor U18264 (N_18264,N_17680,N_17818);
nand U18265 (N_18265,N_17424,N_16294);
nor U18266 (N_18266,N_17430,N_16659);
xor U18267 (N_18267,N_17650,N_17459);
nand U18268 (N_18268,N_17396,N_17537);
nand U18269 (N_18269,N_16783,N_16142);
and U18270 (N_18270,N_16106,N_16262);
nand U18271 (N_18271,N_17522,N_17445);
xor U18272 (N_18272,N_16976,N_17313);
and U18273 (N_18273,N_17875,N_17496);
or U18274 (N_18274,N_16337,N_17633);
xor U18275 (N_18275,N_16769,N_17334);
or U18276 (N_18276,N_17873,N_17881);
nand U18277 (N_18277,N_16709,N_16620);
and U18278 (N_18278,N_17190,N_17998);
and U18279 (N_18279,N_17685,N_16764);
or U18280 (N_18280,N_17391,N_16849);
xor U18281 (N_18281,N_16494,N_16881);
or U18282 (N_18282,N_16822,N_17243);
or U18283 (N_18283,N_17296,N_17018);
nor U18284 (N_18284,N_17037,N_16840);
or U18285 (N_18285,N_17421,N_16702);
nand U18286 (N_18286,N_16059,N_17750);
and U18287 (N_18287,N_16225,N_16807);
or U18288 (N_18288,N_17597,N_17573);
or U18289 (N_18289,N_17489,N_17365);
and U18290 (N_18290,N_16576,N_16798);
nor U18291 (N_18291,N_16054,N_17034);
or U18292 (N_18292,N_17235,N_17840);
xor U18293 (N_18293,N_17299,N_16176);
or U18294 (N_18294,N_16687,N_17102);
nor U18295 (N_18295,N_16105,N_17623);
nand U18296 (N_18296,N_16181,N_17698);
nand U18297 (N_18297,N_16145,N_17017);
or U18298 (N_18298,N_17775,N_16631);
nor U18299 (N_18299,N_17608,N_17645);
nor U18300 (N_18300,N_17485,N_17502);
nor U18301 (N_18301,N_17589,N_16826);
nand U18302 (N_18302,N_16241,N_16821);
nor U18303 (N_18303,N_17968,N_16874);
and U18304 (N_18304,N_16186,N_17431);
and U18305 (N_18305,N_17578,N_16857);
nand U18306 (N_18306,N_17729,N_16762);
nand U18307 (N_18307,N_16699,N_16604);
nand U18308 (N_18308,N_16401,N_16032);
nand U18309 (N_18309,N_16462,N_17586);
nor U18310 (N_18310,N_17411,N_16758);
nor U18311 (N_18311,N_17193,N_16730);
nand U18312 (N_18312,N_17284,N_16089);
or U18313 (N_18313,N_17510,N_16034);
or U18314 (N_18314,N_16636,N_17830);
or U18315 (N_18315,N_16516,N_16901);
xnor U18316 (N_18316,N_17148,N_16944);
nor U18317 (N_18317,N_16554,N_17825);
nand U18318 (N_18318,N_17572,N_16744);
and U18319 (N_18319,N_16793,N_17996);
nor U18320 (N_18320,N_17457,N_17884);
nand U18321 (N_18321,N_16398,N_16694);
and U18322 (N_18322,N_17936,N_17595);
or U18323 (N_18323,N_16995,N_17051);
and U18324 (N_18324,N_17476,N_16217);
nand U18325 (N_18325,N_16301,N_16447);
and U18326 (N_18326,N_17811,N_16022);
xnor U18327 (N_18327,N_16140,N_16848);
nor U18328 (N_18328,N_16539,N_16395);
and U18329 (N_18329,N_17731,N_16103);
xnor U18330 (N_18330,N_17722,N_17630);
or U18331 (N_18331,N_17637,N_16514);
and U18332 (N_18332,N_16155,N_17352);
and U18333 (N_18333,N_17258,N_17934);
nand U18334 (N_18334,N_16266,N_16003);
or U18335 (N_18335,N_16440,N_16858);
xor U18336 (N_18336,N_17016,N_17133);
or U18337 (N_18337,N_17617,N_16866);
nand U18338 (N_18338,N_17805,N_16949);
or U18339 (N_18339,N_17135,N_17665);
or U18340 (N_18340,N_16175,N_17605);
and U18341 (N_18341,N_16571,N_16924);
nor U18342 (N_18342,N_16369,N_16416);
and U18343 (N_18343,N_17541,N_17568);
nand U18344 (N_18344,N_16348,N_16336);
and U18345 (N_18345,N_17677,N_16711);
and U18346 (N_18346,N_17246,N_17471);
nand U18347 (N_18347,N_16680,N_16212);
nand U18348 (N_18348,N_17393,N_16052);
and U18349 (N_18349,N_16472,N_16391);
nand U18350 (N_18350,N_17708,N_17638);
and U18351 (N_18351,N_16580,N_16107);
nand U18352 (N_18352,N_17535,N_17661);
or U18353 (N_18353,N_16973,N_16639);
nor U18354 (N_18354,N_16956,N_17834);
nor U18355 (N_18355,N_16797,N_16990);
nor U18356 (N_18356,N_17239,N_16595);
and U18357 (N_18357,N_16038,N_17434);
nand U18358 (N_18358,N_16487,N_16432);
or U18359 (N_18359,N_16088,N_17204);
or U18360 (N_18360,N_16193,N_16873);
xnor U18361 (N_18361,N_16638,N_17071);
or U18362 (N_18362,N_17821,N_17100);
nand U18363 (N_18363,N_17344,N_17323);
or U18364 (N_18364,N_17277,N_16245);
nand U18365 (N_18365,N_16231,N_17043);
xor U18366 (N_18366,N_17846,N_16794);
and U18367 (N_18367,N_16847,N_16838);
or U18368 (N_18368,N_16836,N_16568);
nor U18369 (N_18369,N_17966,N_16741);
or U18370 (N_18370,N_16414,N_16606);
nor U18371 (N_18371,N_16200,N_16413);
nand U18372 (N_18372,N_16444,N_17160);
nor U18373 (N_18373,N_16473,N_17274);
nor U18374 (N_18374,N_17456,N_17137);
nand U18375 (N_18375,N_16187,N_16725);
and U18376 (N_18376,N_16254,N_16603);
xnor U18377 (N_18377,N_17152,N_17724);
xnor U18378 (N_18378,N_17302,N_16860);
and U18379 (N_18379,N_16698,N_17224);
nor U18380 (N_18380,N_16382,N_17427);
or U18381 (N_18381,N_16162,N_17678);
and U18382 (N_18382,N_16496,N_17790);
nand U18383 (N_18383,N_17889,N_16701);
nand U18384 (N_18384,N_17173,N_16195);
xor U18385 (N_18385,N_17902,N_17795);
nor U18386 (N_18386,N_17492,N_17737);
and U18387 (N_18387,N_16674,N_17165);
nor U18388 (N_18388,N_16977,N_17348);
nor U18389 (N_18389,N_16940,N_17806);
or U18390 (N_18390,N_16523,N_16081);
nor U18391 (N_18391,N_17959,N_16510);
nor U18392 (N_18392,N_16130,N_17282);
nand U18393 (N_18393,N_16994,N_17788);
nor U18394 (N_18394,N_17720,N_16460);
xnor U18395 (N_18395,N_17113,N_16331);
or U18396 (N_18396,N_17009,N_16497);
nand U18397 (N_18397,N_16830,N_17444);
xnor U18398 (N_18398,N_17975,N_17210);
nor U18399 (N_18399,N_17749,N_17030);
or U18400 (N_18400,N_16904,N_16855);
and U18401 (N_18401,N_16470,N_17813);
or U18402 (N_18402,N_16808,N_16865);
or U18403 (N_18403,N_17196,N_17524);
and U18404 (N_18404,N_16772,N_16115);
or U18405 (N_18405,N_17454,N_17801);
nand U18406 (N_18406,N_16828,N_17378);
xnor U18407 (N_18407,N_16870,N_17755);
or U18408 (N_18408,N_17532,N_17049);
and U18409 (N_18409,N_16371,N_17738);
nor U18410 (N_18410,N_16067,N_17028);
xor U18411 (N_18411,N_17178,N_16915);
or U18412 (N_18412,N_17943,N_16878);
nand U18413 (N_18413,N_16310,N_17885);
nor U18414 (N_18414,N_17229,N_17797);
or U18415 (N_18415,N_16282,N_17576);
or U18416 (N_18416,N_16965,N_16168);
nor U18417 (N_18417,N_17023,N_17695);
nor U18418 (N_18418,N_16512,N_17553);
nor U18419 (N_18419,N_16407,N_16450);
nand U18420 (N_18420,N_16047,N_16279);
nand U18421 (N_18421,N_17860,N_16341);
and U18422 (N_18422,N_17984,N_16426);
or U18423 (N_18423,N_17745,N_17551);
nor U18424 (N_18424,N_16926,N_16663);
or U18425 (N_18425,N_17145,N_16295);
nor U18426 (N_18426,N_16459,N_17317);
and U18427 (N_18427,N_16289,N_17958);
nor U18428 (N_18428,N_16953,N_17819);
or U18429 (N_18429,N_17191,N_17259);
and U18430 (N_18430,N_16261,N_16466);
nand U18431 (N_18431,N_16591,N_16880);
nor U18432 (N_18432,N_17504,N_16013);
nor U18433 (N_18433,N_17904,N_17587);
and U18434 (N_18434,N_16775,N_16795);
and U18435 (N_18435,N_17115,N_17560);
nand U18436 (N_18436,N_17442,N_17538);
or U18437 (N_18437,N_17714,N_16952);
or U18438 (N_18438,N_16737,N_16854);
nand U18439 (N_18439,N_16589,N_16160);
or U18440 (N_18440,N_16394,N_16681);
nor U18441 (N_18441,N_16153,N_16986);
and U18442 (N_18442,N_16419,N_16757);
or U18443 (N_18443,N_16693,N_17486);
or U18444 (N_18444,N_16641,N_17426);
and U18445 (N_18445,N_17423,N_16649);
nand U18446 (N_18446,N_16888,N_17542);
or U18447 (N_18447,N_16074,N_16430);
or U18448 (N_18448,N_16307,N_16601);
nand U18449 (N_18449,N_17707,N_16364);
nand U18450 (N_18450,N_16118,N_16933);
nor U18451 (N_18451,N_16070,N_16884);
nand U18452 (N_18452,N_17044,N_17748);
or U18453 (N_18453,N_17271,N_17400);
xor U18454 (N_18454,N_17784,N_16498);
or U18455 (N_18455,N_17127,N_17500);
and U18456 (N_18456,N_16101,N_17170);
or U18457 (N_18457,N_17646,N_16296);
or U18458 (N_18458,N_17961,N_17622);
and U18459 (N_18459,N_16541,N_17076);
and U18460 (N_18460,N_17319,N_17116);
and U18461 (N_18461,N_17886,N_16100);
and U18462 (N_18462,N_16495,N_17085);
xnor U18463 (N_18463,N_17660,N_16825);
nor U18464 (N_18464,N_17599,N_17436);
or U18465 (N_18465,N_17453,N_16561);
nor U18466 (N_18466,N_17081,N_17728);
or U18467 (N_18467,N_16230,N_16246);
nand U18468 (N_18468,N_16152,N_17983);
nand U18469 (N_18469,N_16420,N_17946);
or U18470 (N_18470,N_16347,N_17499);
nor U18471 (N_18471,N_16064,N_16894);
or U18472 (N_18472,N_17694,N_16506);
or U18473 (N_18473,N_16755,N_16887);
or U18474 (N_18474,N_17651,N_17358);
nand U18475 (N_18475,N_16189,N_17088);
nor U18476 (N_18476,N_16752,N_16226);
and U18477 (N_18477,N_17321,N_17221);
and U18478 (N_18478,N_16646,N_17666);
nor U18479 (N_18479,N_16528,N_16599);
nand U18480 (N_18480,N_17783,N_16562);
or U18481 (N_18481,N_17612,N_16964);
or U18482 (N_18482,N_17174,N_17331);
xor U18483 (N_18483,N_16550,N_16536);
nor U18484 (N_18484,N_16742,N_16662);
or U18485 (N_18485,N_17095,N_17377);
nor U18486 (N_18486,N_17472,N_16522);
and U18487 (N_18487,N_17429,N_17752);
nand U18488 (N_18488,N_17624,N_16527);
and U18489 (N_18489,N_16288,N_17458);
and U18490 (N_18490,N_16196,N_16629);
nand U18491 (N_18491,N_16057,N_16027);
nand U18492 (N_18492,N_16570,N_16796);
and U18493 (N_18493,N_17676,N_16283);
and U18494 (N_18494,N_16350,N_17820);
xor U18495 (N_18495,N_16000,N_17997);
nor U18496 (N_18496,N_17656,N_16670);
xnor U18497 (N_18497,N_17894,N_17923);
nand U18498 (N_18498,N_16375,N_16218);
nand U18499 (N_18499,N_17119,N_16834);
and U18500 (N_18500,N_16202,N_17481);
or U18501 (N_18501,N_16036,N_17335);
nand U18502 (N_18502,N_17917,N_16116);
and U18503 (N_18503,N_17407,N_17843);
and U18504 (N_18504,N_16389,N_17764);
or U18505 (N_18505,N_17600,N_16621);
nor U18506 (N_18506,N_17683,N_16543);
or U18507 (N_18507,N_17213,N_17360);
xor U18508 (N_18508,N_17351,N_16132);
nor U18509 (N_18509,N_16504,N_17955);
xor U18510 (N_18510,N_17941,N_16624);
nand U18511 (N_18511,N_16722,N_17552);
xor U18512 (N_18512,N_16648,N_17721);
nand U18513 (N_18513,N_17425,N_17516);
and U18514 (N_18514,N_16360,N_17763);
nand U18515 (N_18515,N_16747,N_16789);
nor U18516 (N_18516,N_17558,N_17526);
or U18517 (N_18517,N_17899,N_17839);
nor U18518 (N_18518,N_17757,N_16320);
nand U18519 (N_18519,N_16824,N_16889);
or U18520 (N_18520,N_16503,N_16204);
xor U18521 (N_18521,N_16384,N_16538);
and U18522 (N_18522,N_16078,N_17000);
and U18523 (N_18523,N_16322,N_16971);
or U18524 (N_18524,N_16438,N_17129);
or U18525 (N_18525,N_16614,N_16785);
xnor U18526 (N_18526,N_16417,N_17070);
nor U18527 (N_18527,N_16087,N_17976);
nand U18528 (N_18528,N_17562,N_17404);
nand U18529 (N_18529,N_17853,N_16549);
nor U18530 (N_18530,N_17503,N_17932);
and U18531 (N_18531,N_17960,N_17285);
xor U18532 (N_18532,N_17908,N_17536);
or U18533 (N_18533,N_16357,N_16963);
xnor U18534 (N_18534,N_16220,N_16387);
or U18535 (N_18535,N_16640,N_17671);
nand U18536 (N_18536,N_17769,N_17789);
and U18537 (N_18537,N_17460,N_16736);
or U18538 (N_18538,N_17021,N_16367);
nand U18539 (N_18539,N_17314,N_16390);
xor U18540 (N_18540,N_16345,N_17947);
or U18541 (N_18541,N_16937,N_16733);
nor U18542 (N_18542,N_17214,N_17794);
nand U18543 (N_18543,N_16819,N_16406);
and U18544 (N_18544,N_17868,N_17495);
or U18545 (N_18545,N_16340,N_17050);
nand U18546 (N_18546,N_17898,N_17123);
nand U18547 (N_18547,N_16802,N_16063);
and U18548 (N_18548,N_16173,N_16875);
nand U18549 (N_18549,N_16359,N_17609);
nor U18550 (N_18550,N_17644,N_17570);
nand U18551 (N_18551,N_16206,N_16851);
and U18552 (N_18552,N_16607,N_16264);
or U18553 (N_18553,N_17149,N_16180);
and U18554 (N_18554,N_16972,N_17117);
nor U18555 (N_18555,N_17026,N_16154);
or U18556 (N_18556,N_17232,N_16511);
nand U18557 (N_18557,N_17703,N_17217);
nor U18558 (N_18558,N_16590,N_17874);
nand U18559 (N_18559,N_16734,N_16981);
xnor U18560 (N_18560,N_17700,N_17778);
or U18561 (N_18561,N_16721,N_17980);
nor U18562 (N_18562,N_16319,N_17531);
nor U18563 (N_18563,N_16260,N_16761);
or U18564 (N_18564,N_16586,N_16392);
nand U18565 (N_18565,N_17327,N_17973);
nand U18566 (N_18566,N_16095,N_16610);
nand U18567 (N_18567,N_17225,N_16914);
nand U18568 (N_18568,N_16537,N_17892);
and U18569 (N_18569,N_16051,N_16784);
xor U18570 (N_18570,N_17337,N_17937);
nand U18571 (N_18571,N_17252,N_17350);
nor U18572 (N_18572,N_17525,N_16685);
nand U18573 (N_18573,N_16751,N_17262);
nor U18574 (N_18574,N_17667,N_16191);
or U18575 (N_18575,N_17292,N_16970);
xnor U18576 (N_18576,N_16656,N_16778);
xor U18577 (N_18577,N_17230,N_17412);
nand U18578 (N_18578,N_17046,N_16707);
and U18579 (N_18579,N_16967,N_17865);
and U18580 (N_18580,N_17470,N_17362);
nand U18581 (N_18581,N_16239,N_17363);
xor U18582 (N_18582,N_16913,N_16678);
and U18583 (N_18583,N_16879,N_17408);
and U18584 (N_18584,N_17452,N_17379);
nor U18585 (N_18585,N_16222,N_16790);
nor U18586 (N_18586,N_17832,N_17057);
and U18587 (N_18587,N_17183,N_16710);
xnor U18588 (N_18588,N_16553,N_17785);
nor U18589 (N_18589,N_16339,N_16135);
xnor U18590 (N_18590,N_16185,N_16433);
and U18591 (N_18591,N_17212,N_17910);
nor U18592 (N_18592,N_17569,N_17041);
nor U18593 (N_18593,N_17371,N_16006);
nor U18594 (N_18594,N_17305,N_17900);
nor U18595 (N_18595,N_16270,N_17090);
nand U18596 (N_18596,N_16692,N_16598);
and U18597 (N_18597,N_17945,N_16779);
nand U18598 (N_18598,N_17078,N_17963);
nor U18599 (N_18599,N_16069,N_17682);
or U18600 (N_18600,N_16745,N_16311);
and U18601 (N_18601,N_16134,N_16040);
or U18602 (N_18602,N_16138,N_16682);
and U18603 (N_18603,N_17142,N_16771);
nand U18604 (N_18604,N_16012,N_16365);
nand U18605 (N_18605,N_16765,N_17227);
nor U18606 (N_18606,N_16731,N_16184);
nand U18607 (N_18607,N_16002,N_17466);
nand U18608 (N_18608,N_17130,N_16574);
xor U18609 (N_18609,N_17896,N_17216);
and U18610 (N_18610,N_17019,N_16718);
nor U18611 (N_18611,N_17032,N_16229);
or U18612 (N_18612,N_16056,N_16985);
or U18613 (N_18613,N_16300,N_17132);
nor U18614 (N_18614,N_17341,N_17206);
or U18615 (N_18615,N_17837,N_17176);
or U18616 (N_18616,N_16756,N_17399);
xor U18617 (N_18617,N_16507,N_16157);
nor U18618 (N_18618,N_16321,N_16431);
and U18619 (N_18619,N_17072,N_16943);
and U18620 (N_18620,N_17131,N_16323);
xor U18621 (N_18621,N_17103,N_16695);
or U18622 (N_18622,N_17841,N_16743);
or U18623 (N_18623,N_16696,N_16163);
xnor U18624 (N_18624,N_16735,N_16801);
nand U18625 (N_18625,N_17592,N_17577);
or U18626 (N_18626,N_17505,N_17287);
nand U18627 (N_18627,N_17851,N_17798);
nand U18628 (N_18628,N_17767,N_17518);
nor U18629 (N_18629,N_17858,N_17290);
nand U18630 (N_18630,N_17218,N_17236);
or U18631 (N_18631,N_16146,N_16946);
or U18632 (N_18632,N_16585,N_17469);
nand U18633 (N_18633,N_17732,N_17726);
xnor U18634 (N_18634,N_16577,N_17356);
or U18635 (N_18635,N_16679,N_16517);
nand U18636 (N_18636,N_17202,N_16558);
or U18637 (N_18637,N_17260,N_17546);
nand U18638 (N_18638,N_17802,N_17091);
xnor U18639 (N_18639,N_16324,N_17629);
nor U18640 (N_18640,N_17280,N_16697);
nand U18641 (N_18641,N_16373,N_17852);
and U18642 (N_18642,N_16275,N_17188);
nand U18643 (N_18643,N_17059,N_17008);
nor U18644 (N_18644,N_17375,N_17047);
nor U18645 (N_18645,N_16418,N_16408);
nor U18646 (N_18646,N_17372,N_17942);
nand U18647 (N_18647,N_16112,N_16645);
nor U18648 (N_18648,N_16713,N_16039);
or U18649 (N_18649,N_17836,N_17370);
or U18650 (N_18650,N_16293,N_17529);
and U18651 (N_18651,N_16613,N_17374);
or U18652 (N_18652,N_16706,N_16156);
nand U18653 (N_18653,N_17247,N_16513);
or U18654 (N_18654,N_17530,N_17780);
nor U18655 (N_18655,N_17406,N_16197);
nor U18656 (N_18656,N_17359,N_16248);
nor U18657 (N_18657,N_16931,N_16363);
nor U18658 (N_18658,N_17376,N_16328);
or U18659 (N_18659,N_16628,N_17122);
nor U18660 (N_18660,N_17982,N_17035);
or U18661 (N_18661,N_16723,N_16564);
or U18662 (N_18662,N_17557,N_16968);
nor U18663 (N_18663,N_17799,N_17092);
nor U18664 (N_18664,N_16941,N_17422);
and U18665 (N_18665,N_17010,N_17971);
or U18666 (N_18666,N_17523,N_17978);
and U18667 (N_18667,N_17300,N_17539);
and U18668 (N_18668,N_16644,N_17601);
nand U18669 (N_18669,N_17672,N_17548);
and U18670 (N_18670,N_16732,N_17613);
and U18671 (N_18671,N_16273,N_16179);
or U18672 (N_18672,N_16445,N_16096);
nor U18673 (N_18673,N_16381,N_16183);
or U18674 (N_18674,N_17626,N_16353);
nand U18675 (N_18675,N_17042,N_17497);
nor U18676 (N_18676,N_17120,N_17099);
and U18677 (N_18677,N_17565,N_17207);
nand U18678 (N_18678,N_17093,N_17416);
and U18679 (N_18679,N_17111,N_16099);
nand U18680 (N_18680,N_16263,N_17867);
and U18681 (N_18681,N_17628,N_17809);
nand U18682 (N_18682,N_17684,N_16642);
or U18683 (N_18683,N_16127,N_16439);
xor U18684 (N_18684,N_16344,N_16508);
or U18685 (N_18685,N_17706,N_17075);
nor U18686 (N_18686,N_16704,N_17871);
nand U18687 (N_18687,N_17582,N_16883);
or U18688 (N_18688,N_16425,N_17940);
and U18689 (N_18689,N_17447,N_17625);
and U18690 (N_18690,N_17414,N_16676);
nor U18691 (N_18691,N_16423,N_17669);
and U18692 (N_18692,N_17347,N_17872);
nand U18693 (N_18693,N_16332,N_17108);
nor U18694 (N_18694,N_16024,N_16110);
nand U18695 (N_18695,N_16739,N_16531);
nor U18696 (N_18696,N_16637,N_17621);
or U18697 (N_18697,N_16867,N_17804);
and U18698 (N_18698,N_16475,N_16895);
nor U18699 (N_18699,N_17697,N_17087);
nor U18700 (N_18700,N_17709,N_17413);
and U18701 (N_18701,N_17068,N_17163);
nand U18702 (N_18702,N_16660,N_17632);
or U18703 (N_18703,N_17332,N_17555);
or U18704 (N_18704,N_17197,N_17594);
nor U18705 (N_18705,N_16017,N_16905);
and U18706 (N_18706,N_17686,N_16316);
nor U18707 (N_18707,N_16557,N_16893);
nor U18708 (N_18708,N_17635,N_16076);
and U18709 (N_18709,N_16820,N_16073);
nand U18710 (N_18710,N_17355,N_16534);
and U18711 (N_18711,N_16593,N_17473);
nor U18712 (N_18712,N_17079,N_17005);
and U18713 (N_18713,N_16551,N_17981);
nor U18714 (N_18714,N_17616,N_17550);
or U18715 (N_18715,N_17668,N_17066);
nand U18716 (N_18716,N_16930,N_17554);
and U18717 (N_18717,N_16393,N_16740);
and U18718 (N_18718,N_17226,N_16313);
nand U18719 (N_18719,N_17822,N_17480);
or U18720 (N_18720,N_17567,N_17125);
nor U18721 (N_18721,N_16856,N_17003);
or U18722 (N_18722,N_16996,N_17654);
nor U18723 (N_18723,N_17186,N_16376);
nand U18724 (N_18724,N_17301,N_16945);
nor U18725 (N_18725,N_17346,N_16214);
nor U18726 (N_18726,N_16252,N_17584);
nand U18727 (N_18727,N_17488,N_17859);
nor U18728 (N_18728,N_17831,N_16787);
xnor U18729 (N_18729,N_17402,N_17405);
nor U18730 (N_18730,N_17991,N_17520);
nand U18731 (N_18731,N_16188,N_16111);
xor U18732 (N_18732,N_16249,N_17664);
xnor U18733 (N_18733,N_17164,N_16041);
and U18734 (N_18734,N_17124,N_17343);
nand U18735 (N_18735,N_17766,N_16240);
nor U18736 (N_18736,N_17443,N_16652);
or U18737 (N_18737,N_16846,N_17463);
nand U18738 (N_18738,N_16983,N_16961);
nor U18739 (N_18739,N_17954,N_17288);
nor U18740 (N_18740,N_17106,N_16090);
nand U18741 (N_18741,N_17596,N_17508);
or U18742 (N_18742,N_16243,N_16890);
or U18743 (N_18743,N_17639,N_16259);
nor U18744 (N_18744,N_16190,N_16427);
nor U18745 (N_18745,N_17256,N_16616);
nand U18746 (N_18746,N_17141,N_16396);
and U18747 (N_18747,N_17527,N_16048);
or U18748 (N_18748,N_16164,N_17511);
nor U18749 (N_18749,N_17739,N_17642);
xnor U18750 (N_18750,N_16515,N_16228);
or U18751 (N_18751,N_16244,N_17307);
nor U18752 (N_18752,N_17320,N_16633);
and U18753 (N_18753,N_16647,N_17006);
or U18754 (N_18754,N_16488,N_17251);
or U18755 (N_18755,N_17827,N_16882);
and U18756 (N_18756,N_17845,N_17704);
or U18757 (N_18757,N_16690,N_16066);
and U18758 (N_18758,N_17295,N_16729);
nor U18759 (N_18759,N_17328,N_16182);
nor U18760 (N_18760,N_16596,N_16309);
nor U18761 (N_18761,N_16597,N_17776);
xnor U18762 (N_18762,N_16521,N_17450);
or U18763 (N_18763,N_17921,N_17544);
nor U18764 (N_18764,N_16724,N_16533);
or U18765 (N_18765,N_16863,N_17110);
nor U18766 (N_18766,N_16501,N_16151);
nor U18767 (N_18767,N_17401,N_16955);
and U18768 (N_18768,N_16546,N_16664);
xnor U18769 (N_18769,N_16815,N_16091);
nand U18770 (N_18770,N_16842,N_16299);
nand U18771 (N_18771,N_17388,N_17479);
and U18772 (N_18772,N_16560,N_17659);
or U18773 (N_18773,N_17330,N_16542);
or U18774 (N_18774,N_16285,N_17002);
nor U18775 (N_18775,N_17368,N_16530);
or U18776 (N_18776,N_17240,N_16476);
xor U18777 (N_18777,N_17838,N_16899);
nor U18778 (N_18778,N_17712,N_17662);
or U18779 (N_18779,N_17304,N_16030);
or U18780 (N_18780,N_17760,N_16383);
nor U18781 (N_18781,N_16832,N_17439);
nor U18782 (N_18782,N_17774,N_16982);
nor U18783 (N_18783,N_17342,N_16627);
nor U18784 (N_18784,N_17636,N_17564);
nand U18785 (N_18785,N_16330,N_17409);
xnor U18786 (N_18786,N_16385,N_16404);
or U18787 (N_18787,N_16104,N_17033);
nor U18788 (N_18788,N_16916,N_17782);
nand U18789 (N_18789,N_16306,N_16446);
or U18790 (N_18790,N_17244,N_16247);
and U18791 (N_18791,N_16573,N_16234);
or U18792 (N_18792,N_17254,N_16015);
and U18793 (N_18793,N_17951,N_17611);
nand U18794 (N_18794,N_17972,N_17333);
and U18795 (N_18795,N_17389,N_16774);
or U18796 (N_18796,N_17357,N_17603);
or U18797 (N_18797,N_16050,N_17390);
and U18798 (N_18798,N_16886,N_17864);
nand U18799 (N_18799,N_17415,N_17746);
and U18800 (N_18800,N_17857,N_16068);
xor U18801 (N_18801,N_16872,N_17705);
and U18802 (N_18802,N_17803,N_16748);
and U18803 (N_18803,N_17273,N_17967);
and U18804 (N_18804,N_17013,N_16675);
nor U18805 (N_18805,N_17509,N_17772);
and U18806 (N_18806,N_16362,N_17238);
nor U18807 (N_18807,N_17468,N_16354);
xnor U18808 (N_18808,N_16559,N_17069);
and U18809 (N_18809,N_16272,N_16211);
or U18810 (N_18810,N_17716,N_17563);
and U18811 (N_18811,N_17717,N_16552);
nand U18812 (N_18812,N_16966,N_16178);
or U18813 (N_18813,N_16456,N_17310);
nor U18814 (N_18814,N_17547,N_16172);
or U18815 (N_18815,N_17279,N_17992);
nand U18816 (N_18816,N_17829,N_16026);
or U18817 (N_18817,N_16975,N_16237);
nand U18818 (N_18818,N_16084,N_17985);
or U18819 (N_18819,N_17222,N_17549);
and U18820 (N_18820,N_16065,N_16018);
or U18821 (N_18821,N_16978,N_16746);
nand U18822 (N_18822,N_17264,N_16062);
nand U18823 (N_18823,N_16754,N_16208);
and U18824 (N_18824,N_16061,N_16448);
nand U18825 (N_18825,N_16284,N_17844);
and U18826 (N_18826,N_17198,N_16669);
or U18827 (N_18827,N_17847,N_16780);
nand U18828 (N_18828,N_16898,N_17879);
nand U18829 (N_18829,N_17652,N_16902);
nand U18830 (N_18830,N_17999,N_17861);
or U18831 (N_18831,N_16969,N_17025);
or U18832 (N_18832,N_16668,N_17195);
nor U18833 (N_18833,N_17580,N_16415);
nor U18834 (N_18834,N_17751,N_17199);
and U18835 (N_18835,N_17098,N_17640);
nor U18836 (N_18836,N_16612,N_16529);
and U18837 (N_18837,N_16776,N_16346);
and U18838 (N_18838,N_17435,N_16055);
xnor U18839 (N_18839,N_17607,N_17237);
nand U18840 (N_18840,N_17315,N_16150);
or U18841 (N_18841,N_17933,N_16939);
nand U18842 (N_18842,N_17154,N_17521);
or U18843 (N_18843,N_17631,N_16932);
nor U18844 (N_18844,N_17338,N_17663);
nor U18845 (N_18845,N_17336,N_17658);
nor U18846 (N_18846,N_17887,N_16097);
and U18847 (N_18847,N_16672,N_17316);
nand U18848 (N_18848,N_16519,N_16388);
or U18849 (N_18849,N_16588,N_17808);
and U18850 (N_18850,N_16950,N_17781);
or U18851 (N_18851,N_16500,N_16490);
nand U18852 (N_18852,N_17911,N_17517);
and U18853 (N_18853,N_16708,N_16703);
nor U18854 (N_18854,N_16120,N_16147);
or U18855 (N_18855,N_17903,N_16810);
or U18856 (N_18856,N_16657,N_17157);
nand U18857 (N_18857,N_16329,N_17255);
nor U18858 (N_18858,N_16166,N_17077);
and U18859 (N_18859,N_17048,N_16750);
and U18860 (N_18860,N_16556,N_16864);
or U18861 (N_18861,N_16792,N_17514);
nor U18862 (N_18862,N_17311,N_16079);
xor U18863 (N_18863,N_16816,N_17209);
or U18864 (N_18864,N_16974,N_17494);
xnor U18865 (N_18865,N_16993,N_16651);
and U18866 (N_18866,N_16871,N_16900);
or U18867 (N_18867,N_16683,N_17297);
or U18868 (N_18868,N_16452,N_17528);
nor U18869 (N_18869,N_16581,N_17673);
nand U18870 (N_18870,N_17817,N_17876);
or U18871 (N_18871,N_16449,N_16049);
or U18872 (N_18872,N_16028,N_16213);
or U18873 (N_18873,N_16934,N_17270);
nand U18874 (N_18874,N_16540,N_17467);
nor U18875 (N_18875,N_16635,N_16399);
nand U18876 (N_18876,N_17166,N_16303);
or U18877 (N_18877,N_17962,N_16113);
nor U18878 (N_18878,N_16072,N_17970);
nor U18879 (N_18879,N_17906,N_16923);
xor U18880 (N_18880,N_17935,N_17581);
or U18881 (N_18881,N_16169,N_16326);
nand U18882 (N_18882,N_17104,N_16619);
and U18883 (N_18883,N_17107,N_17619);
nor U18884 (N_18884,N_16043,N_17475);
and U18885 (N_18885,N_16632,N_16813);
xor U18886 (N_18886,N_17895,N_17162);
xor U18887 (N_18887,N_17719,N_17324);
nand U18888 (N_18888,N_17989,N_16803);
and U18889 (N_18889,N_17073,N_16853);
and U18890 (N_18890,N_17114,N_17432);
xnor U18891 (N_18891,N_16271,N_16763);
nand U18892 (N_18892,N_17948,N_17771);
or U18893 (N_18893,N_17223,N_16979);
and U18894 (N_18894,N_17150,N_17128);
or U18895 (N_18895,N_16378,N_16379);
nand U18896 (N_18896,N_16844,N_17606);
nand U18897 (N_18897,N_17944,N_17015);
nor U18898 (N_18898,N_17590,N_16287);
or U18899 (N_18899,N_16505,N_16655);
or U18900 (N_18900,N_16897,N_17498);
nor U18901 (N_18901,N_16009,N_17787);
nand U18902 (N_18902,N_17200,N_17779);
or U18903 (N_18903,N_16267,N_16948);
xor U18904 (N_18904,N_16333,N_16093);
nand U18905 (N_18905,N_17192,N_16167);
and U18906 (N_18906,N_17687,N_16909);
xor U18907 (N_18907,N_16714,N_17339);
nand U18908 (N_18908,N_17045,N_16927);
nand U18909 (N_18909,N_16422,N_16129);
or U18910 (N_18910,N_17696,N_17807);
nor U18911 (N_18911,N_16661,N_17325);
and U18912 (N_18912,N_16080,N_17063);
nand U18913 (N_18913,N_17863,N_17734);
nor U18914 (N_18914,N_17448,N_17294);
or U18915 (N_18915,N_17233,N_16298);
nor U18916 (N_18916,N_17765,N_16782);
nand U18917 (N_18917,N_16005,N_17245);
nand U18918 (N_18918,N_17691,N_17913);
nand U18919 (N_18919,N_16499,N_17303);
or U18920 (N_18920,N_16045,N_17743);
and U18921 (N_18921,N_17266,N_17702);
nor U18922 (N_18922,N_17927,N_17988);
and U18923 (N_18923,N_16161,N_16290);
nor U18924 (N_18924,N_16467,N_16143);
and U18925 (N_18925,N_16700,N_16720);
and U18926 (N_18926,N_16335,N_17814);
xor U18927 (N_18927,N_17507,N_16622);
nand U18928 (N_18928,N_16016,N_17440);
nor U18929 (N_18929,N_16159,N_17248);
xor U18930 (N_18930,N_17545,N_17298);
or U18931 (N_18931,N_17289,N_16623);
nand U18932 (N_18932,N_17909,N_17112);
xor U18933 (N_18933,N_17730,N_17773);
nand U18934 (N_18934,N_17770,N_16643);
or U18935 (N_18935,N_16876,N_16102);
nor U18936 (N_18936,N_17559,N_16630);
or U18937 (N_18937,N_17561,N_16221);
and U18938 (N_18938,N_16125,N_17634);
and U18939 (N_18939,N_17241,N_17446);
nor U18940 (N_18940,N_17395,N_16468);
or U18941 (N_18941,N_17964,N_17907);
xor U18942 (N_18942,N_16342,N_16992);
xnor U18943 (N_18943,N_16122,N_17096);
nor U18944 (N_18944,N_16171,N_16165);
nand U18945 (N_18945,N_17461,N_17744);
and U18946 (N_18946,N_16205,N_16251);
and U18947 (N_18947,N_17060,N_16019);
and U18948 (N_18948,N_16454,N_17674);
nand U18949 (N_18949,N_16942,N_16256);
nor U18950 (N_18950,N_17168,N_17140);
nor U18951 (N_18951,N_17151,N_17074);
or U18952 (N_18952,N_17924,N_16429);
nand U18953 (N_18953,N_16997,N_16717);
or U18954 (N_18954,N_17969,N_16014);
or U18955 (N_18955,N_16907,N_16843);
or U18956 (N_18956,N_16085,N_16223);
and U18957 (N_18957,N_16885,N_16489);
xor U18958 (N_18958,N_17727,N_17278);
xnor U18959 (N_18959,N_16453,N_16852);
nand U18960 (N_18960,N_17891,N_16349);
and U18961 (N_18961,N_17930,N_17286);
xnor U18962 (N_18962,N_17263,N_17939);
or U18963 (N_18963,N_16318,N_17381);
xor U18964 (N_18964,N_16377,N_16833);
or U18965 (N_18965,N_16509,N_17883);
nor U18966 (N_18966,N_16114,N_16286);
or U18967 (N_18967,N_17253,N_16749);
or U18968 (N_18968,N_16938,N_16811);
or U18969 (N_18969,N_16565,N_17501);
and U18970 (N_18970,N_17354,N_17928);
xnor U18971 (N_18971,N_16219,N_16029);
xnor U18972 (N_18972,N_16411,N_16402);
and U18973 (N_18973,N_17147,N_16917);
and U18974 (N_18974,N_16987,N_16033);
or U18975 (N_18975,N_16611,N_17848);
nand U18976 (N_18976,N_17146,N_17571);
nor U18977 (N_18977,N_16908,N_16957);
or U18978 (N_18978,N_16799,N_17053);
nand U18979 (N_18979,N_16148,N_16020);
nor U18980 (N_18980,N_17441,N_16892);
and U18981 (N_18981,N_16991,N_17403);
or U18982 (N_18982,N_16464,N_16845);
nor U18983 (N_18983,N_17742,N_16575);
nor U18984 (N_18984,N_17062,N_16215);
nand U18985 (N_18985,N_17679,N_16370);
nor U18986 (N_18986,N_17800,N_16823);
or U18987 (N_18987,N_17768,N_16921);
and U18988 (N_18988,N_17641,N_16804);
or U18989 (N_18989,N_17979,N_17723);
or U18990 (N_18990,N_16001,N_17901);
nor U18991 (N_18991,N_17345,N_17574);
and U18992 (N_18992,N_17022,N_17701);
and U18993 (N_18993,N_16358,N_17777);
xor U18994 (N_18994,N_16579,N_16583);
or U18995 (N_18995,N_16292,N_17397);
nor U18996 (N_18996,N_17309,N_17326);
nor U18997 (N_18997,N_16207,N_16753);
xor U18998 (N_18998,N_17455,N_17591);
nor U18999 (N_18999,N_16315,N_16194);
nor U19000 (N_19000,N_17298,N_16970);
nand U19001 (N_19001,N_16966,N_16136);
nor U19002 (N_19002,N_17184,N_16750);
nor U19003 (N_19003,N_16881,N_17491);
and U19004 (N_19004,N_16017,N_16790);
nor U19005 (N_19005,N_17244,N_17337);
or U19006 (N_19006,N_17519,N_17081);
and U19007 (N_19007,N_16536,N_17944);
xnor U19008 (N_19008,N_16109,N_17355);
and U19009 (N_19009,N_17729,N_17935);
and U19010 (N_19010,N_16841,N_17253);
nand U19011 (N_19011,N_16919,N_17543);
nor U19012 (N_19012,N_16676,N_16342);
or U19013 (N_19013,N_17029,N_17504);
nor U19014 (N_19014,N_16151,N_17709);
and U19015 (N_19015,N_17025,N_16216);
nand U19016 (N_19016,N_16374,N_17125);
and U19017 (N_19017,N_16788,N_17198);
nand U19018 (N_19018,N_17393,N_16755);
or U19019 (N_19019,N_16299,N_17013);
nor U19020 (N_19020,N_17257,N_16899);
nand U19021 (N_19021,N_17860,N_17958);
xor U19022 (N_19022,N_17254,N_17385);
or U19023 (N_19023,N_17607,N_16651);
xor U19024 (N_19024,N_16368,N_17108);
xnor U19025 (N_19025,N_17896,N_17007);
or U19026 (N_19026,N_16081,N_17546);
nor U19027 (N_19027,N_16931,N_17053);
and U19028 (N_19028,N_16083,N_17186);
and U19029 (N_19029,N_17006,N_16347);
and U19030 (N_19030,N_17864,N_17484);
or U19031 (N_19031,N_16717,N_17201);
or U19032 (N_19032,N_16202,N_17216);
and U19033 (N_19033,N_17040,N_16008);
nor U19034 (N_19034,N_17968,N_16668);
nor U19035 (N_19035,N_17598,N_17538);
or U19036 (N_19036,N_17016,N_17203);
nor U19037 (N_19037,N_17177,N_17272);
and U19038 (N_19038,N_16472,N_16454);
nand U19039 (N_19039,N_17757,N_17067);
xor U19040 (N_19040,N_17988,N_16701);
or U19041 (N_19041,N_16488,N_17052);
nand U19042 (N_19042,N_17096,N_16492);
or U19043 (N_19043,N_16278,N_16186);
xor U19044 (N_19044,N_17500,N_16075);
xor U19045 (N_19045,N_16924,N_17065);
xnor U19046 (N_19046,N_16602,N_16840);
nor U19047 (N_19047,N_16743,N_16299);
nor U19048 (N_19048,N_17762,N_17111);
nand U19049 (N_19049,N_17307,N_17689);
or U19050 (N_19050,N_16659,N_17508);
or U19051 (N_19051,N_17413,N_16723);
nand U19052 (N_19052,N_16087,N_17807);
or U19053 (N_19053,N_16171,N_17484);
and U19054 (N_19054,N_16939,N_17651);
nor U19055 (N_19055,N_17200,N_16553);
nor U19056 (N_19056,N_16903,N_16570);
nand U19057 (N_19057,N_16592,N_16933);
or U19058 (N_19058,N_16165,N_17826);
nand U19059 (N_19059,N_17355,N_16633);
or U19060 (N_19060,N_17680,N_16722);
nand U19061 (N_19061,N_16247,N_17365);
nor U19062 (N_19062,N_17893,N_16434);
and U19063 (N_19063,N_17899,N_16015);
nand U19064 (N_19064,N_17284,N_16795);
nor U19065 (N_19065,N_17278,N_16017);
xnor U19066 (N_19066,N_17094,N_17915);
xor U19067 (N_19067,N_16854,N_17589);
and U19068 (N_19068,N_17254,N_16269);
and U19069 (N_19069,N_16418,N_17748);
and U19070 (N_19070,N_16978,N_16497);
xor U19071 (N_19071,N_16646,N_16819);
nand U19072 (N_19072,N_17727,N_17298);
nand U19073 (N_19073,N_17186,N_17266);
nand U19074 (N_19074,N_16404,N_17976);
nor U19075 (N_19075,N_16992,N_16755);
and U19076 (N_19076,N_16832,N_17371);
and U19077 (N_19077,N_16004,N_17599);
nand U19078 (N_19078,N_16316,N_17512);
or U19079 (N_19079,N_16344,N_17130);
xnor U19080 (N_19080,N_16008,N_17447);
xor U19081 (N_19081,N_17054,N_17852);
nor U19082 (N_19082,N_17554,N_16286);
or U19083 (N_19083,N_16193,N_16619);
or U19084 (N_19084,N_17902,N_16504);
nor U19085 (N_19085,N_17670,N_17402);
nor U19086 (N_19086,N_16455,N_17818);
or U19087 (N_19087,N_17491,N_17082);
and U19088 (N_19088,N_17656,N_16773);
and U19089 (N_19089,N_16906,N_16142);
nor U19090 (N_19090,N_16220,N_17053);
xnor U19091 (N_19091,N_16794,N_16770);
xnor U19092 (N_19092,N_16640,N_17260);
nand U19093 (N_19093,N_16066,N_16259);
or U19094 (N_19094,N_17945,N_16612);
nor U19095 (N_19095,N_16465,N_16276);
and U19096 (N_19096,N_16542,N_16130);
nand U19097 (N_19097,N_16522,N_17952);
xnor U19098 (N_19098,N_17907,N_16010);
and U19099 (N_19099,N_17685,N_17938);
or U19100 (N_19100,N_16548,N_16550);
nand U19101 (N_19101,N_16382,N_16925);
and U19102 (N_19102,N_17969,N_16183);
nand U19103 (N_19103,N_16266,N_16567);
nand U19104 (N_19104,N_17927,N_16273);
and U19105 (N_19105,N_17674,N_17658);
nor U19106 (N_19106,N_16465,N_16547);
or U19107 (N_19107,N_17307,N_17438);
xor U19108 (N_19108,N_17676,N_16830);
and U19109 (N_19109,N_16834,N_16826);
or U19110 (N_19110,N_17241,N_16748);
nor U19111 (N_19111,N_17109,N_16159);
or U19112 (N_19112,N_16014,N_16570);
xnor U19113 (N_19113,N_17786,N_17184);
nor U19114 (N_19114,N_16562,N_17736);
or U19115 (N_19115,N_16979,N_16420);
nor U19116 (N_19116,N_16513,N_17599);
and U19117 (N_19117,N_17294,N_16699);
xnor U19118 (N_19118,N_16313,N_17049);
or U19119 (N_19119,N_17087,N_17719);
nor U19120 (N_19120,N_17946,N_16951);
and U19121 (N_19121,N_17919,N_17242);
and U19122 (N_19122,N_17383,N_16262);
or U19123 (N_19123,N_17619,N_17993);
or U19124 (N_19124,N_16251,N_16867);
nand U19125 (N_19125,N_16825,N_17514);
or U19126 (N_19126,N_16799,N_16365);
nand U19127 (N_19127,N_16383,N_17674);
or U19128 (N_19128,N_16585,N_17572);
and U19129 (N_19129,N_17353,N_17061);
or U19130 (N_19130,N_17488,N_16690);
xor U19131 (N_19131,N_16634,N_16000);
xnor U19132 (N_19132,N_16877,N_16551);
nand U19133 (N_19133,N_17346,N_17065);
or U19134 (N_19134,N_17720,N_16770);
nand U19135 (N_19135,N_16388,N_17248);
or U19136 (N_19136,N_17972,N_16942);
and U19137 (N_19137,N_17408,N_16719);
or U19138 (N_19138,N_16541,N_17983);
or U19139 (N_19139,N_17261,N_17927);
xor U19140 (N_19140,N_16633,N_16578);
or U19141 (N_19141,N_17552,N_16491);
and U19142 (N_19142,N_17738,N_17829);
nand U19143 (N_19143,N_17489,N_17864);
and U19144 (N_19144,N_17082,N_17469);
xnor U19145 (N_19145,N_16933,N_17168);
nor U19146 (N_19146,N_16049,N_16753);
nor U19147 (N_19147,N_16561,N_17006);
xor U19148 (N_19148,N_17900,N_17441);
nand U19149 (N_19149,N_16012,N_17125);
nor U19150 (N_19150,N_17240,N_16873);
nor U19151 (N_19151,N_17322,N_16000);
nor U19152 (N_19152,N_16128,N_16385);
or U19153 (N_19153,N_17739,N_16536);
or U19154 (N_19154,N_16896,N_17714);
or U19155 (N_19155,N_17813,N_16430);
nor U19156 (N_19156,N_17955,N_16521);
or U19157 (N_19157,N_17116,N_17803);
or U19158 (N_19158,N_16162,N_16450);
nand U19159 (N_19159,N_17465,N_16850);
nor U19160 (N_19160,N_16208,N_16317);
and U19161 (N_19161,N_16233,N_16299);
nand U19162 (N_19162,N_17535,N_17492);
or U19163 (N_19163,N_17925,N_16982);
xnor U19164 (N_19164,N_17437,N_16995);
and U19165 (N_19165,N_17275,N_17691);
and U19166 (N_19166,N_16943,N_17309);
or U19167 (N_19167,N_17256,N_16872);
or U19168 (N_19168,N_17984,N_16276);
nand U19169 (N_19169,N_16161,N_16074);
or U19170 (N_19170,N_16261,N_16696);
nor U19171 (N_19171,N_16462,N_17140);
nor U19172 (N_19172,N_16728,N_17197);
nor U19173 (N_19173,N_17435,N_16697);
nand U19174 (N_19174,N_17560,N_16374);
nand U19175 (N_19175,N_17581,N_16589);
and U19176 (N_19176,N_16365,N_17353);
nand U19177 (N_19177,N_16761,N_16384);
or U19178 (N_19178,N_17787,N_16700);
xor U19179 (N_19179,N_17421,N_17317);
nor U19180 (N_19180,N_17852,N_16430);
or U19181 (N_19181,N_16933,N_17119);
and U19182 (N_19182,N_16064,N_16903);
and U19183 (N_19183,N_17354,N_16357);
nor U19184 (N_19184,N_17656,N_17871);
xnor U19185 (N_19185,N_16484,N_16724);
nand U19186 (N_19186,N_17184,N_16764);
nor U19187 (N_19187,N_17931,N_16021);
or U19188 (N_19188,N_16383,N_17027);
nand U19189 (N_19189,N_17583,N_17750);
and U19190 (N_19190,N_17706,N_16645);
nor U19191 (N_19191,N_16062,N_17291);
nor U19192 (N_19192,N_17939,N_16200);
nor U19193 (N_19193,N_17223,N_16665);
or U19194 (N_19194,N_16466,N_17255);
or U19195 (N_19195,N_17337,N_17205);
or U19196 (N_19196,N_17750,N_17417);
or U19197 (N_19197,N_16944,N_16530);
and U19198 (N_19198,N_16618,N_16398);
and U19199 (N_19199,N_17190,N_17225);
nand U19200 (N_19200,N_17367,N_16200);
and U19201 (N_19201,N_16172,N_17087);
or U19202 (N_19202,N_16629,N_17586);
and U19203 (N_19203,N_16465,N_17721);
and U19204 (N_19204,N_16296,N_17441);
nand U19205 (N_19205,N_16837,N_17256);
or U19206 (N_19206,N_16419,N_16227);
and U19207 (N_19207,N_17427,N_16665);
or U19208 (N_19208,N_17364,N_16291);
nand U19209 (N_19209,N_16645,N_16299);
or U19210 (N_19210,N_16072,N_16135);
nand U19211 (N_19211,N_17791,N_17189);
and U19212 (N_19212,N_16773,N_17184);
nor U19213 (N_19213,N_17952,N_17393);
or U19214 (N_19214,N_16773,N_17694);
xor U19215 (N_19215,N_16715,N_17789);
nor U19216 (N_19216,N_16370,N_16244);
or U19217 (N_19217,N_17325,N_16979);
nor U19218 (N_19218,N_17354,N_17707);
or U19219 (N_19219,N_17943,N_17362);
and U19220 (N_19220,N_17178,N_17374);
or U19221 (N_19221,N_17818,N_17356);
or U19222 (N_19222,N_16297,N_17219);
nor U19223 (N_19223,N_17345,N_17023);
nor U19224 (N_19224,N_16221,N_17370);
and U19225 (N_19225,N_17065,N_16638);
xor U19226 (N_19226,N_17264,N_17241);
nor U19227 (N_19227,N_17288,N_16284);
xnor U19228 (N_19228,N_16156,N_17882);
or U19229 (N_19229,N_17878,N_16936);
nand U19230 (N_19230,N_17911,N_17636);
nor U19231 (N_19231,N_16787,N_17961);
and U19232 (N_19232,N_16057,N_17530);
nand U19233 (N_19233,N_16614,N_16504);
xor U19234 (N_19234,N_17678,N_16519);
or U19235 (N_19235,N_17131,N_17200);
nor U19236 (N_19236,N_17339,N_17241);
and U19237 (N_19237,N_16899,N_17416);
or U19238 (N_19238,N_17378,N_17690);
nand U19239 (N_19239,N_17274,N_17616);
nor U19240 (N_19240,N_17653,N_17844);
or U19241 (N_19241,N_17114,N_17154);
or U19242 (N_19242,N_16453,N_16407);
and U19243 (N_19243,N_16871,N_17935);
nand U19244 (N_19244,N_16899,N_16306);
nor U19245 (N_19245,N_16123,N_16885);
and U19246 (N_19246,N_17426,N_17390);
nor U19247 (N_19247,N_17428,N_17726);
and U19248 (N_19248,N_16853,N_16969);
and U19249 (N_19249,N_16533,N_16593);
and U19250 (N_19250,N_16650,N_16046);
xnor U19251 (N_19251,N_16597,N_16367);
and U19252 (N_19252,N_17710,N_17383);
nand U19253 (N_19253,N_17741,N_17522);
or U19254 (N_19254,N_16166,N_17711);
and U19255 (N_19255,N_17116,N_17235);
and U19256 (N_19256,N_16249,N_16600);
or U19257 (N_19257,N_17649,N_16130);
nand U19258 (N_19258,N_16244,N_16493);
and U19259 (N_19259,N_16895,N_17261);
or U19260 (N_19260,N_16331,N_16407);
and U19261 (N_19261,N_16323,N_17961);
or U19262 (N_19262,N_17346,N_17316);
nand U19263 (N_19263,N_16224,N_17463);
or U19264 (N_19264,N_16056,N_17873);
and U19265 (N_19265,N_16608,N_16324);
or U19266 (N_19266,N_16913,N_17934);
nand U19267 (N_19267,N_17426,N_17921);
nand U19268 (N_19268,N_17674,N_17394);
nor U19269 (N_19269,N_17147,N_16836);
nand U19270 (N_19270,N_16135,N_17290);
nand U19271 (N_19271,N_17883,N_17552);
and U19272 (N_19272,N_17363,N_16483);
and U19273 (N_19273,N_17637,N_16013);
and U19274 (N_19274,N_17587,N_16884);
and U19275 (N_19275,N_16224,N_17949);
or U19276 (N_19276,N_17268,N_17933);
nor U19277 (N_19277,N_17655,N_17524);
and U19278 (N_19278,N_17894,N_17436);
nand U19279 (N_19279,N_16776,N_16924);
nor U19280 (N_19280,N_17546,N_17787);
and U19281 (N_19281,N_16804,N_17450);
nor U19282 (N_19282,N_16178,N_17713);
and U19283 (N_19283,N_17266,N_17066);
or U19284 (N_19284,N_16883,N_17019);
nand U19285 (N_19285,N_17106,N_17769);
nor U19286 (N_19286,N_16162,N_16856);
nor U19287 (N_19287,N_17984,N_16388);
nand U19288 (N_19288,N_17066,N_17977);
or U19289 (N_19289,N_16393,N_17903);
or U19290 (N_19290,N_17922,N_17393);
or U19291 (N_19291,N_17336,N_16949);
and U19292 (N_19292,N_16386,N_17709);
and U19293 (N_19293,N_16330,N_17170);
and U19294 (N_19294,N_16720,N_17786);
nand U19295 (N_19295,N_16847,N_16383);
and U19296 (N_19296,N_16594,N_16439);
xor U19297 (N_19297,N_17042,N_16495);
or U19298 (N_19298,N_17117,N_17566);
and U19299 (N_19299,N_17706,N_17295);
and U19300 (N_19300,N_17836,N_17447);
or U19301 (N_19301,N_16188,N_16285);
and U19302 (N_19302,N_16390,N_16816);
and U19303 (N_19303,N_16834,N_16865);
or U19304 (N_19304,N_16678,N_17572);
nand U19305 (N_19305,N_16713,N_17280);
or U19306 (N_19306,N_16071,N_16332);
nor U19307 (N_19307,N_17614,N_16245);
or U19308 (N_19308,N_16046,N_16055);
nor U19309 (N_19309,N_16775,N_17091);
nor U19310 (N_19310,N_16426,N_17185);
nor U19311 (N_19311,N_16469,N_16845);
and U19312 (N_19312,N_16854,N_16581);
nor U19313 (N_19313,N_16459,N_17262);
and U19314 (N_19314,N_16143,N_17097);
xnor U19315 (N_19315,N_16253,N_16758);
and U19316 (N_19316,N_16038,N_16292);
and U19317 (N_19317,N_16728,N_16573);
nand U19318 (N_19318,N_16531,N_17515);
or U19319 (N_19319,N_17567,N_17879);
and U19320 (N_19320,N_17916,N_16221);
nand U19321 (N_19321,N_16912,N_16309);
or U19322 (N_19322,N_17251,N_17727);
nor U19323 (N_19323,N_16870,N_17426);
or U19324 (N_19324,N_17825,N_16842);
nor U19325 (N_19325,N_17590,N_17340);
nor U19326 (N_19326,N_17137,N_16365);
or U19327 (N_19327,N_16187,N_17684);
nand U19328 (N_19328,N_16007,N_16531);
and U19329 (N_19329,N_17780,N_16419);
nand U19330 (N_19330,N_16510,N_17641);
or U19331 (N_19331,N_17473,N_17713);
nand U19332 (N_19332,N_17931,N_17191);
nand U19333 (N_19333,N_17715,N_17818);
nand U19334 (N_19334,N_17230,N_17356);
or U19335 (N_19335,N_16871,N_17754);
and U19336 (N_19336,N_16789,N_16503);
nand U19337 (N_19337,N_16214,N_16423);
nand U19338 (N_19338,N_17837,N_16501);
and U19339 (N_19339,N_16550,N_17037);
nand U19340 (N_19340,N_16671,N_17304);
and U19341 (N_19341,N_17769,N_16168);
or U19342 (N_19342,N_17838,N_16459);
nand U19343 (N_19343,N_17719,N_16727);
xnor U19344 (N_19344,N_17176,N_17941);
nand U19345 (N_19345,N_17090,N_16969);
xor U19346 (N_19346,N_16363,N_17781);
nand U19347 (N_19347,N_17139,N_16094);
and U19348 (N_19348,N_16541,N_16077);
nand U19349 (N_19349,N_16313,N_16728);
nand U19350 (N_19350,N_17774,N_16178);
and U19351 (N_19351,N_16866,N_16852);
nor U19352 (N_19352,N_17245,N_17891);
or U19353 (N_19353,N_17014,N_17974);
and U19354 (N_19354,N_17637,N_17522);
and U19355 (N_19355,N_16383,N_17743);
and U19356 (N_19356,N_17773,N_17876);
nor U19357 (N_19357,N_16299,N_16807);
xor U19358 (N_19358,N_17696,N_17970);
and U19359 (N_19359,N_17474,N_17357);
and U19360 (N_19360,N_16876,N_16973);
nand U19361 (N_19361,N_17077,N_16778);
and U19362 (N_19362,N_17699,N_16589);
and U19363 (N_19363,N_16794,N_17020);
nor U19364 (N_19364,N_16511,N_17086);
nor U19365 (N_19365,N_17465,N_16487);
nand U19366 (N_19366,N_17867,N_17586);
xnor U19367 (N_19367,N_17130,N_16300);
or U19368 (N_19368,N_17909,N_16099);
and U19369 (N_19369,N_16223,N_17626);
and U19370 (N_19370,N_16235,N_17267);
or U19371 (N_19371,N_16158,N_16699);
nor U19372 (N_19372,N_16194,N_16461);
and U19373 (N_19373,N_17507,N_16624);
or U19374 (N_19374,N_16789,N_16966);
nand U19375 (N_19375,N_17412,N_16566);
nand U19376 (N_19376,N_17384,N_17714);
or U19377 (N_19377,N_17542,N_16552);
or U19378 (N_19378,N_17413,N_16887);
or U19379 (N_19379,N_17311,N_16135);
nand U19380 (N_19380,N_16662,N_16339);
or U19381 (N_19381,N_17094,N_16085);
nand U19382 (N_19382,N_16234,N_16757);
nand U19383 (N_19383,N_17230,N_16343);
and U19384 (N_19384,N_17876,N_16514);
nand U19385 (N_19385,N_17251,N_16569);
and U19386 (N_19386,N_17220,N_16565);
nor U19387 (N_19387,N_16813,N_17098);
or U19388 (N_19388,N_17426,N_16943);
nor U19389 (N_19389,N_17874,N_16400);
and U19390 (N_19390,N_16991,N_17539);
nand U19391 (N_19391,N_17547,N_16352);
xnor U19392 (N_19392,N_16450,N_17101);
nand U19393 (N_19393,N_16903,N_17348);
and U19394 (N_19394,N_16350,N_17472);
or U19395 (N_19395,N_17109,N_17851);
nor U19396 (N_19396,N_17439,N_17377);
xnor U19397 (N_19397,N_16525,N_16139);
or U19398 (N_19398,N_17893,N_16145);
nor U19399 (N_19399,N_17567,N_16014);
or U19400 (N_19400,N_16293,N_16345);
xor U19401 (N_19401,N_17408,N_17047);
nor U19402 (N_19402,N_17711,N_16463);
nor U19403 (N_19403,N_16106,N_16107);
xor U19404 (N_19404,N_17462,N_17966);
nor U19405 (N_19405,N_16071,N_17022);
xnor U19406 (N_19406,N_16858,N_16970);
xnor U19407 (N_19407,N_17726,N_17080);
or U19408 (N_19408,N_16404,N_16021);
and U19409 (N_19409,N_17629,N_16832);
xnor U19410 (N_19410,N_16733,N_16138);
nand U19411 (N_19411,N_17823,N_17329);
xor U19412 (N_19412,N_16269,N_16874);
nor U19413 (N_19413,N_16912,N_16625);
or U19414 (N_19414,N_17858,N_17766);
nor U19415 (N_19415,N_16573,N_16098);
and U19416 (N_19416,N_17997,N_16667);
and U19417 (N_19417,N_17224,N_17565);
or U19418 (N_19418,N_16889,N_17456);
nand U19419 (N_19419,N_17746,N_17718);
nor U19420 (N_19420,N_17473,N_16087);
or U19421 (N_19421,N_16745,N_17019);
xnor U19422 (N_19422,N_17976,N_16252);
xor U19423 (N_19423,N_16210,N_17597);
xnor U19424 (N_19424,N_16326,N_16404);
nor U19425 (N_19425,N_16700,N_17918);
or U19426 (N_19426,N_17897,N_17431);
nor U19427 (N_19427,N_16261,N_17157);
nand U19428 (N_19428,N_16622,N_16777);
nor U19429 (N_19429,N_16394,N_17292);
and U19430 (N_19430,N_16986,N_16801);
and U19431 (N_19431,N_17031,N_17980);
and U19432 (N_19432,N_16410,N_16926);
nand U19433 (N_19433,N_16238,N_17480);
nor U19434 (N_19434,N_16819,N_16953);
nor U19435 (N_19435,N_16556,N_16320);
nor U19436 (N_19436,N_16054,N_17885);
nand U19437 (N_19437,N_17143,N_17117);
or U19438 (N_19438,N_16517,N_16544);
or U19439 (N_19439,N_16633,N_16359);
or U19440 (N_19440,N_17886,N_16707);
and U19441 (N_19441,N_16472,N_17124);
nor U19442 (N_19442,N_17900,N_16751);
nand U19443 (N_19443,N_17852,N_16840);
xnor U19444 (N_19444,N_16593,N_16832);
nor U19445 (N_19445,N_17269,N_17005);
nor U19446 (N_19446,N_16505,N_16025);
nor U19447 (N_19447,N_16673,N_17674);
nand U19448 (N_19448,N_17659,N_16744);
and U19449 (N_19449,N_16873,N_16020);
and U19450 (N_19450,N_16538,N_17299);
nand U19451 (N_19451,N_17925,N_17329);
xor U19452 (N_19452,N_16832,N_17372);
or U19453 (N_19453,N_17623,N_16775);
or U19454 (N_19454,N_17712,N_16013);
or U19455 (N_19455,N_16446,N_16724);
or U19456 (N_19456,N_17612,N_16726);
nor U19457 (N_19457,N_16439,N_16015);
nand U19458 (N_19458,N_16948,N_16517);
nor U19459 (N_19459,N_16866,N_16268);
nor U19460 (N_19460,N_17499,N_16950);
nor U19461 (N_19461,N_17278,N_17045);
nand U19462 (N_19462,N_16374,N_16721);
and U19463 (N_19463,N_16471,N_17774);
nand U19464 (N_19464,N_17574,N_17986);
xnor U19465 (N_19465,N_17118,N_17379);
nor U19466 (N_19466,N_16392,N_16699);
or U19467 (N_19467,N_17250,N_16237);
nand U19468 (N_19468,N_17926,N_16399);
and U19469 (N_19469,N_17001,N_17654);
nand U19470 (N_19470,N_16332,N_16564);
and U19471 (N_19471,N_16931,N_17173);
and U19472 (N_19472,N_16409,N_16152);
and U19473 (N_19473,N_16266,N_16757);
nand U19474 (N_19474,N_17702,N_16333);
nor U19475 (N_19475,N_17033,N_17632);
or U19476 (N_19476,N_16045,N_17902);
nand U19477 (N_19477,N_16549,N_16006);
and U19478 (N_19478,N_16901,N_17124);
xnor U19479 (N_19479,N_16289,N_16916);
or U19480 (N_19480,N_16475,N_17794);
and U19481 (N_19481,N_17815,N_17982);
or U19482 (N_19482,N_17621,N_17328);
nor U19483 (N_19483,N_17906,N_16345);
or U19484 (N_19484,N_17684,N_17341);
or U19485 (N_19485,N_17556,N_17879);
xor U19486 (N_19486,N_16598,N_16331);
nor U19487 (N_19487,N_17358,N_16287);
or U19488 (N_19488,N_16298,N_17594);
and U19489 (N_19489,N_16953,N_17862);
or U19490 (N_19490,N_17240,N_16840);
nand U19491 (N_19491,N_17685,N_16685);
nor U19492 (N_19492,N_16909,N_16851);
nor U19493 (N_19493,N_16230,N_17801);
nand U19494 (N_19494,N_16383,N_17433);
xnor U19495 (N_19495,N_16652,N_17618);
xnor U19496 (N_19496,N_16565,N_16765);
or U19497 (N_19497,N_16775,N_16495);
nand U19498 (N_19498,N_17219,N_16643);
and U19499 (N_19499,N_16755,N_17001);
or U19500 (N_19500,N_17622,N_17819);
nand U19501 (N_19501,N_17858,N_16745);
or U19502 (N_19502,N_16239,N_16165);
or U19503 (N_19503,N_16400,N_16152);
nor U19504 (N_19504,N_16626,N_17891);
nor U19505 (N_19505,N_16135,N_17509);
nand U19506 (N_19506,N_17147,N_17407);
nand U19507 (N_19507,N_17058,N_16266);
nor U19508 (N_19508,N_17104,N_16470);
nor U19509 (N_19509,N_17183,N_17763);
or U19510 (N_19510,N_16723,N_16181);
and U19511 (N_19511,N_17027,N_17861);
nor U19512 (N_19512,N_16419,N_17347);
nor U19513 (N_19513,N_16949,N_16840);
and U19514 (N_19514,N_16376,N_17961);
or U19515 (N_19515,N_17285,N_16865);
or U19516 (N_19516,N_17895,N_16005);
nor U19517 (N_19517,N_16753,N_17554);
xor U19518 (N_19518,N_16311,N_17767);
or U19519 (N_19519,N_17210,N_16950);
nor U19520 (N_19520,N_17354,N_17483);
or U19521 (N_19521,N_16560,N_16734);
or U19522 (N_19522,N_16478,N_16054);
nor U19523 (N_19523,N_16494,N_16410);
or U19524 (N_19524,N_16598,N_17974);
xnor U19525 (N_19525,N_16151,N_17115);
and U19526 (N_19526,N_16598,N_17495);
nor U19527 (N_19527,N_17731,N_17000);
nor U19528 (N_19528,N_16241,N_16786);
xor U19529 (N_19529,N_16790,N_16118);
xnor U19530 (N_19530,N_17190,N_16625);
or U19531 (N_19531,N_17144,N_17571);
and U19532 (N_19532,N_17702,N_16329);
or U19533 (N_19533,N_17270,N_17548);
nor U19534 (N_19534,N_17275,N_17495);
and U19535 (N_19535,N_16950,N_16332);
and U19536 (N_19536,N_16248,N_16302);
or U19537 (N_19537,N_16391,N_16575);
and U19538 (N_19538,N_16967,N_16366);
nor U19539 (N_19539,N_16333,N_16339);
or U19540 (N_19540,N_17366,N_16644);
xor U19541 (N_19541,N_17487,N_17683);
or U19542 (N_19542,N_17444,N_17241);
nand U19543 (N_19543,N_17095,N_16787);
xor U19544 (N_19544,N_16421,N_17029);
nor U19545 (N_19545,N_16977,N_16369);
nand U19546 (N_19546,N_16667,N_17759);
or U19547 (N_19547,N_17604,N_17561);
or U19548 (N_19548,N_16752,N_17781);
and U19549 (N_19549,N_16948,N_16230);
and U19550 (N_19550,N_17535,N_16940);
nor U19551 (N_19551,N_17157,N_17570);
or U19552 (N_19552,N_16587,N_16633);
or U19553 (N_19553,N_16237,N_16791);
or U19554 (N_19554,N_16496,N_16627);
nor U19555 (N_19555,N_16867,N_16028);
and U19556 (N_19556,N_17792,N_16738);
nand U19557 (N_19557,N_17288,N_16928);
or U19558 (N_19558,N_17963,N_17033);
and U19559 (N_19559,N_16328,N_16231);
nor U19560 (N_19560,N_17691,N_16696);
or U19561 (N_19561,N_16259,N_17071);
nor U19562 (N_19562,N_17342,N_17954);
xnor U19563 (N_19563,N_16513,N_17404);
xor U19564 (N_19564,N_16702,N_16475);
nor U19565 (N_19565,N_16499,N_17462);
or U19566 (N_19566,N_16772,N_17801);
and U19567 (N_19567,N_17684,N_16806);
nor U19568 (N_19568,N_17311,N_16429);
and U19569 (N_19569,N_16199,N_16925);
and U19570 (N_19570,N_17061,N_16527);
nor U19571 (N_19571,N_16477,N_17905);
and U19572 (N_19572,N_16228,N_16972);
nor U19573 (N_19573,N_16884,N_16367);
nor U19574 (N_19574,N_17266,N_16776);
nand U19575 (N_19575,N_16066,N_17275);
nor U19576 (N_19576,N_17398,N_17725);
nand U19577 (N_19577,N_17535,N_17466);
nand U19578 (N_19578,N_17796,N_17836);
nand U19579 (N_19579,N_16604,N_16422);
xor U19580 (N_19580,N_17165,N_17633);
or U19581 (N_19581,N_17132,N_16476);
or U19582 (N_19582,N_16430,N_16084);
and U19583 (N_19583,N_17352,N_17451);
or U19584 (N_19584,N_17621,N_16198);
or U19585 (N_19585,N_16452,N_17730);
and U19586 (N_19586,N_16782,N_17002);
and U19587 (N_19587,N_16403,N_17402);
nor U19588 (N_19588,N_16139,N_17477);
nor U19589 (N_19589,N_17828,N_16008);
nand U19590 (N_19590,N_17760,N_16318);
and U19591 (N_19591,N_17320,N_17228);
and U19592 (N_19592,N_16386,N_17200);
nor U19593 (N_19593,N_17742,N_16149);
nand U19594 (N_19594,N_16186,N_16881);
or U19595 (N_19595,N_17839,N_17125);
and U19596 (N_19596,N_17457,N_17152);
nor U19597 (N_19597,N_17150,N_16463);
or U19598 (N_19598,N_16995,N_16124);
nor U19599 (N_19599,N_17844,N_16556);
nand U19600 (N_19600,N_16485,N_17626);
and U19601 (N_19601,N_17204,N_17036);
nand U19602 (N_19602,N_17582,N_16741);
or U19603 (N_19603,N_16475,N_16462);
nor U19604 (N_19604,N_17962,N_17253);
and U19605 (N_19605,N_16707,N_17793);
nor U19606 (N_19606,N_17832,N_16459);
and U19607 (N_19607,N_16534,N_17545);
nand U19608 (N_19608,N_17998,N_16862);
or U19609 (N_19609,N_16272,N_16347);
and U19610 (N_19610,N_17432,N_16147);
nor U19611 (N_19611,N_17407,N_17462);
nor U19612 (N_19612,N_17194,N_17255);
or U19613 (N_19613,N_17550,N_17309);
xnor U19614 (N_19614,N_16259,N_16675);
or U19615 (N_19615,N_17173,N_16234);
xnor U19616 (N_19616,N_16721,N_16438);
nand U19617 (N_19617,N_17436,N_17288);
nor U19618 (N_19618,N_17763,N_16145);
nor U19619 (N_19619,N_17200,N_16135);
or U19620 (N_19620,N_16901,N_16361);
xnor U19621 (N_19621,N_16319,N_17790);
nand U19622 (N_19622,N_17825,N_16862);
nor U19623 (N_19623,N_17886,N_17630);
or U19624 (N_19624,N_17585,N_16662);
and U19625 (N_19625,N_17621,N_17182);
nand U19626 (N_19626,N_16136,N_16857);
or U19627 (N_19627,N_16723,N_17388);
nor U19628 (N_19628,N_16694,N_17667);
or U19629 (N_19629,N_16308,N_16433);
nor U19630 (N_19630,N_17227,N_16414);
nand U19631 (N_19631,N_16988,N_17623);
nor U19632 (N_19632,N_16202,N_16938);
or U19633 (N_19633,N_16307,N_17849);
nor U19634 (N_19634,N_16386,N_17190);
and U19635 (N_19635,N_17320,N_17694);
nand U19636 (N_19636,N_16993,N_17883);
nand U19637 (N_19637,N_16341,N_17354);
nand U19638 (N_19638,N_16344,N_16440);
xor U19639 (N_19639,N_17842,N_17024);
or U19640 (N_19640,N_17637,N_16259);
or U19641 (N_19641,N_17747,N_16613);
nand U19642 (N_19642,N_16656,N_17396);
or U19643 (N_19643,N_17841,N_16411);
nor U19644 (N_19644,N_16397,N_17785);
nor U19645 (N_19645,N_17478,N_17232);
xor U19646 (N_19646,N_17760,N_16473);
nor U19647 (N_19647,N_16235,N_16187);
or U19648 (N_19648,N_16621,N_16658);
nand U19649 (N_19649,N_17295,N_16572);
and U19650 (N_19650,N_17384,N_17469);
nor U19651 (N_19651,N_16178,N_17175);
nand U19652 (N_19652,N_17798,N_16864);
xor U19653 (N_19653,N_16496,N_16037);
or U19654 (N_19654,N_16821,N_17983);
or U19655 (N_19655,N_16115,N_17771);
and U19656 (N_19656,N_16128,N_16737);
nor U19657 (N_19657,N_17224,N_17188);
xnor U19658 (N_19658,N_16235,N_16531);
nor U19659 (N_19659,N_17660,N_17943);
nor U19660 (N_19660,N_17652,N_16821);
xnor U19661 (N_19661,N_16327,N_17171);
or U19662 (N_19662,N_17688,N_16559);
or U19663 (N_19663,N_17359,N_17788);
nor U19664 (N_19664,N_16745,N_16716);
or U19665 (N_19665,N_17707,N_16362);
nand U19666 (N_19666,N_17195,N_17520);
or U19667 (N_19667,N_16840,N_16271);
or U19668 (N_19668,N_16397,N_16606);
nand U19669 (N_19669,N_17620,N_17889);
nand U19670 (N_19670,N_17616,N_17885);
or U19671 (N_19671,N_17134,N_17186);
and U19672 (N_19672,N_16770,N_16153);
nor U19673 (N_19673,N_16146,N_16274);
or U19674 (N_19674,N_16947,N_16695);
or U19675 (N_19675,N_17840,N_16845);
or U19676 (N_19676,N_16891,N_17840);
nand U19677 (N_19677,N_16290,N_16193);
nand U19678 (N_19678,N_16484,N_16011);
nor U19679 (N_19679,N_16082,N_17116);
and U19680 (N_19680,N_16192,N_17448);
nand U19681 (N_19681,N_17826,N_17261);
nand U19682 (N_19682,N_17977,N_16878);
xor U19683 (N_19683,N_17885,N_16972);
and U19684 (N_19684,N_16923,N_16108);
or U19685 (N_19685,N_16060,N_16453);
nor U19686 (N_19686,N_16221,N_17009);
or U19687 (N_19687,N_16485,N_17418);
or U19688 (N_19688,N_17939,N_16631);
or U19689 (N_19689,N_17056,N_16063);
nor U19690 (N_19690,N_16729,N_16138);
nor U19691 (N_19691,N_17980,N_16002);
and U19692 (N_19692,N_16997,N_17868);
or U19693 (N_19693,N_17509,N_17248);
or U19694 (N_19694,N_17327,N_16337);
and U19695 (N_19695,N_16278,N_16482);
or U19696 (N_19696,N_16797,N_16060);
or U19697 (N_19697,N_17249,N_17050);
and U19698 (N_19698,N_17203,N_17249);
nor U19699 (N_19699,N_16555,N_17065);
and U19700 (N_19700,N_16674,N_16447);
nand U19701 (N_19701,N_17723,N_17942);
or U19702 (N_19702,N_16910,N_17330);
and U19703 (N_19703,N_17159,N_17112);
nand U19704 (N_19704,N_17549,N_17665);
nand U19705 (N_19705,N_17172,N_17773);
nor U19706 (N_19706,N_16919,N_16454);
or U19707 (N_19707,N_17815,N_16469);
nand U19708 (N_19708,N_17586,N_17866);
nor U19709 (N_19709,N_16538,N_17576);
or U19710 (N_19710,N_17414,N_17953);
nand U19711 (N_19711,N_16794,N_16520);
xnor U19712 (N_19712,N_17168,N_16688);
or U19713 (N_19713,N_16274,N_16807);
or U19714 (N_19714,N_16169,N_16909);
xor U19715 (N_19715,N_16506,N_17355);
and U19716 (N_19716,N_16575,N_17777);
nand U19717 (N_19717,N_16221,N_16814);
nor U19718 (N_19718,N_17328,N_17390);
nand U19719 (N_19719,N_16527,N_16777);
nand U19720 (N_19720,N_16967,N_16921);
nand U19721 (N_19721,N_17526,N_17118);
nand U19722 (N_19722,N_16217,N_16371);
and U19723 (N_19723,N_16503,N_16656);
xor U19724 (N_19724,N_16616,N_16827);
nor U19725 (N_19725,N_16828,N_17680);
nor U19726 (N_19726,N_17159,N_16908);
nor U19727 (N_19727,N_17527,N_16345);
and U19728 (N_19728,N_17069,N_16297);
nand U19729 (N_19729,N_17785,N_17450);
and U19730 (N_19730,N_17781,N_16537);
nand U19731 (N_19731,N_17784,N_17480);
nor U19732 (N_19732,N_17704,N_16876);
or U19733 (N_19733,N_17071,N_17972);
nor U19734 (N_19734,N_16830,N_16451);
nor U19735 (N_19735,N_16075,N_17655);
nand U19736 (N_19736,N_17221,N_16871);
xnor U19737 (N_19737,N_17887,N_16203);
or U19738 (N_19738,N_17963,N_17495);
or U19739 (N_19739,N_16725,N_17044);
nor U19740 (N_19740,N_17472,N_17177);
nor U19741 (N_19741,N_17701,N_16353);
and U19742 (N_19742,N_17225,N_16667);
nor U19743 (N_19743,N_16801,N_17279);
or U19744 (N_19744,N_16393,N_17101);
nor U19745 (N_19745,N_17322,N_17182);
or U19746 (N_19746,N_16411,N_17059);
or U19747 (N_19747,N_17440,N_16134);
nor U19748 (N_19748,N_16689,N_17122);
and U19749 (N_19749,N_16180,N_17620);
nor U19750 (N_19750,N_16363,N_17117);
and U19751 (N_19751,N_16842,N_16110);
and U19752 (N_19752,N_16556,N_17734);
nand U19753 (N_19753,N_17222,N_16285);
nand U19754 (N_19754,N_16693,N_16571);
xnor U19755 (N_19755,N_17477,N_16003);
nor U19756 (N_19756,N_16101,N_16189);
or U19757 (N_19757,N_17088,N_17246);
and U19758 (N_19758,N_17005,N_16770);
and U19759 (N_19759,N_17074,N_16644);
and U19760 (N_19760,N_16361,N_17999);
nand U19761 (N_19761,N_16097,N_16266);
or U19762 (N_19762,N_16642,N_17914);
and U19763 (N_19763,N_16991,N_16734);
nand U19764 (N_19764,N_16558,N_16660);
nand U19765 (N_19765,N_16070,N_16487);
and U19766 (N_19766,N_17885,N_16895);
and U19767 (N_19767,N_16832,N_17183);
xnor U19768 (N_19768,N_17051,N_17247);
nand U19769 (N_19769,N_17248,N_17633);
nor U19770 (N_19770,N_16493,N_17075);
xor U19771 (N_19771,N_16031,N_16989);
nor U19772 (N_19772,N_16957,N_17730);
nor U19773 (N_19773,N_17971,N_17489);
nor U19774 (N_19774,N_16532,N_17814);
or U19775 (N_19775,N_17696,N_17931);
and U19776 (N_19776,N_16823,N_17325);
nor U19777 (N_19777,N_16265,N_16611);
and U19778 (N_19778,N_17300,N_16633);
nand U19779 (N_19779,N_17463,N_16476);
nand U19780 (N_19780,N_16359,N_17246);
or U19781 (N_19781,N_16323,N_17975);
or U19782 (N_19782,N_17473,N_16221);
nor U19783 (N_19783,N_16731,N_17927);
nor U19784 (N_19784,N_17650,N_17945);
nand U19785 (N_19785,N_17928,N_17029);
or U19786 (N_19786,N_17319,N_17529);
nor U19787 (N_19787,N_17027,N_16487);
nor U19788 (N_19788,N_16284,N_16213);
nor U19789 (N_19789,N_17600,N_17416);
nor U19790 (N_19790,N_16918,N_17939);
nor U19791 (N_19791,N_16140,N_16665);
nand U19792 (N_19792,N_17354,N_16664);
nor U19793 (N_19793,N_17957,N_16176);
and U19794 (N_19794,N_17430,N_17706);
or U19795 (N_19795,N_17530,N_17829);
nor U19796 (N_19796,N_16951,N_16804);
nor U19797 (N_19797,N_17593,N_17346);
and U19798 (N_19798,N_17959,N_16126);
or U19799 (N_19799,N_16512,N_17101);
xor U19800 (N_19800,N_16818,N_17204);
nor U19801 (N_19801,N_16029,N_16289);
and U19802 (N_19802,N_16903,N_16367);
or U19803 (N_19803,N_16106,N_17236);
xor U19804 (N_19804,N_16643,N_16078);
xor U19805 (N_19805,N_16929,N_17329);
and U19806 (N_19806,N_16027,N_17557);
xnor U19807 (N_19807,N_16183,N_16186);
or U19808 (N_19808,N_17913,N_16590);
nor U19809 (N_19809,N_17026,N_17231);
or U19810 (N_19810,N_16948,N_16726);
xor U19811 (N_19811,N_17278,N_17842);
nor U19812 (N_19812,N_16461,N_16577);
nor U19813 (N_19813,N_16964,N_16311);
nand U19814 (N_19814,N_16419,N_17084);
or U19815 (N_19815,N_17361,N_17215);
nor U19816 (N_19816,N_17433,N_16518);
or U19817 (N_19817,N_17614,N_17107);
or U19818 (N_19818,N_17519,N_16027);
xor U19819 (N_19819,N_16658,N_17051);
xor U19820 (N_19820,N_17536,N_16313);
and U19821 (N_19821,N_16874,N_17244);
and U19822 (N_19822,N_17567,N_16078);
or U19823 (N_19823,N_16472,N_17811);
and U19824 (N_19824,N_17245,N_16384);
nand U19825 (N_19825,N_17995,N_16079);
nand U19826 (N_19826,N_16899,N_16650);
nor U19827 (N_19827,N_17554,N_16598);
nor U19828 (N_19828,N_17272,N_17485);
and U19829 (N_19829,N_16457,N_16760);
nor U19830 (N_19830,N_17422,N_17850);
and U19831 (N_19831,N_16868,N_17052);
nand U19832 (N_19832,N_16717,N_17315);
nand U19833 (N_19833,N_17491,N_17328);
nand U19834 (N_19834,N_17368,N_16392);
nand U19835 (N_19835,N_17964,N_16277);
nand U19836 (N_19836,N_16359,N_16539);
and U19837 (N_19837,N_17654,N_16507);
xor U19838 (N_19838,N_16560,N_16776);
nor U19839 (N_19839,N_17034,N_17289);
or U19840 (N_19840,N_16263,N_17205);
and U19841 (N_19841,N_17960,N_17495);
xor U19842 (N_19842,N_17923,N_16565);
nor U19843 (N_19843,N_16344,N_16118);
nand U19844 (N_19844,N_16644,N_16202);
nor U19845 (N_19845,N_16089,N_17074);
nor U19846 (N_19846,N_17480,N_16856);
or U19847 (N_19847,N_17433,N_16755);
and U19848 (N_19848,N_17052,N_17718);
xor U19849 (N_19849,N_17645,N_17123);
xor U19850 (N_19850,N_17206,N_16951);
nand U19851 (N_19851,N_17597,N_16538);
nand U19852 (N_19852,N_17597,N_17171);
nand U19853 (N_19853,N_17413,N_16194);
and U19854 (N_19854,N_16840,N_17970);
nor U19855 (N_19855,N_17927,N_16477);
nor U19856 (N_19856,N_17315,N_17986);
nor U19857 (N_19857,N_17483,N_17171);
or U19858 (N_19858,N_16300,N_16101);
or U19859 (N_19859,N_17752,N_16826);
nor U19860 (N_19860,N_17405,N_16848);
and U19861 (N_19861,N_17395,N_17558);
nand U19862 (N_19862,N_16463,N_16028);
nor U19863 (N_19863,N_17360,N_17945);
nor U19864 (N_19864,N_17112,N_16394);
nor U19865 (N_19865,N_17717,N_16085);
nor U19866 (N_19866,N_16716,N_17186);
xor U19867 (N_19867,N_17814,N_17304);
nor U19868 (N_19868,N_16524,N_17863);
nor U19869 (N_19869,N_16839,N_16686);
and U19870 (N_19870,N_17422,N_16357);
or U19871 (N_19871,N_17682,N_16646);
nand U19872 (N_19872,N_17030,N_17051);
nand U19873 (N_19873,N_16994,N_17745);
nand U19874 (N_19874,N_17712,N_16903);
or U19875 (N_19875,N_17876,N_17389);
and U19876 (N_19876,N_17942,N_17479);
nand U19877 (N_19877,N_17493,N_16616);
and U19878 (N_19878,N_16601,N_16063);
nand U19879 (N_19879,N_16132,N_17069);
nand U19880 (N_19880,N_17993,N_17105);
or U19881 (N_19881,N_17105,N_16903);
or U19882 (N_19882,N_16756,N_17769);
xor U19883 (N_19883,N_17003,N_16609);
or U19884 (N_19884,N_17548,N_17914);
and U19885 (N_19885,N_17267,N_17745);
nor U19886 (N_19886,N_17131,N_16492);
nand U19887 (N_19887,N_16828,N_17962);
and U19888 (N_19888,N_17953,N_17682);
and U19889 (N_19889,N_17078,N_17606);
and U19890 (N_19890,N_17990,N_17213);
or U19891 (N_19891,N_17748,N_16350);
and U19892 (N_19892,N_16321,N_17326);
nor U19893 (N_19893,N_16784,N_16768);
or U19894 (N_19894,N_16902,N_17138);
or U19895 (N_19895,N_17158,N_16335);
or U19896 (N_19896,N_17723,N_17221);
and U19897 (N_19897,N_16357,N_17472);
nand U19898 (N_19898,N_16601,N_17479);
nand U19899 (N_19899,N_16624,N_16011);
and U19900 (N_19900,N_17662,N_17675);
nand U19901 (N_19901,N_17841,N_17129);
or U19902 (N_19902,N_17903,N_17772);
nand U19903 (N_19903,N_17484,N_16931);
and U19904 (N_19904,N_17624,N_17280);
nand U19905 (N_19905,N_17835,N_16789);
nor U19906 (N_19906,N_16323,N_16343);
nand U19907 (N_19907,N_16302,N_16361);
nor U19908 (N_19908,N_16706,N_16527);
and U19909 (N_19909,N_17754,N_16329);
or U19910 (N_19910,N_17390,N_16682);
nand U19911 (N_19911,N_17650,N_17460);
and U19912 (N_19912,N_16000,N_16608);
or U19913 (N_19913,N_17982,N_16067);
and U19914 (N_19914,N_17354,N_17015);
nor U19915 (N_19915,N_16479,N_16330);
and U19916 (N_19916,N_16847,N_17997);
and U19917 (N_19917,N_17867,N_16390);
nor U19918 (N_19918,N_16417,N_17967);
or U19919 (N_19919,N_17929,N_17464);
or U19920 (N_19920,N_17921,N_16809);
or U19921 (N_19921,N_16868,N_16783);
nand U19922 (N_19922,N_16810,N_17897);
or U19923 (N_19923,N_16451,N_17927);
or U19924 (N_19924,N_16120,N_16552);
or U19925 (N_19925,N_16736,N_16780);
xnor U19926 (N_19926,N_17042,N_17494);
nand U19927 (N_19927,N_16471,N_16287);
nor U19928 (N_19928,N_17015,N_16797);
nor U19929 (N_19929,N_16962,N_16624);
nor U19930 (N_19930,N_17699,N_17693);
nand U19931 (N_19931,N_16699,N_16517);
nor U19932 (N_19932,N_16224,N_16180);
or U19933 (N_19933,N_16810,N_16097);
or U19934 (N_19934,N_17377,N_17120);
or U19935 (N_19935,N_17470,N_17229);
or U19936 (N_19936,N_17314,N_17977);
nand U19937 (N_19937,N_16268,N_17531);
or U19938 (N_19938,N_17024,N_16858);
nand U19939 (N_19939,N_17425,N_17387);
and U19940 (N_19940,N_17593,N_17185);
and U19941 (N_19941,N_17083,N_17360);
nor U19942 (N_19942,N_17207,N_17745);
xnor U19943 (N_19943,N_16974,N_16437);
or U19944 (N_19944,N_16674,N_17280);
xnor U19945 (N_19945,N_17345,N_17167);
nand U19946 (N_19946,N_16769,N_17142);
or U19947 (N_19947,N_17890,N_17807);
nand U19948 (N_19948,N_16395,N_16145);
nor U19949 (N_19949,N_16583,N_17721);
or U19950 (N_19950,N_17910,N_17028);
nor U19951 (N_19951,N_17316,N_16112);
nand U19952 (N_19952,N_16691,N_16681);
nor U19953 (N_19953,N_17898,N_16752);
nand U19954 (N_19954,N_17189,N_16194);
nor U19955 (N_19955,N_16640,N_16921);
and U19956 (N_19956,N_17325,N_16626);
nor U19957 (N_19957,N_16299,N_17554);
nor U19958 (N_19958,N_17085,N_16890);
nor U19959 (N_19959,N_17759,N_16219);
and U19960 (N_19960,N_17216,N_17879);
and U19961 (N_19961,N_16857,N_16542);
nor U19962 (N_19962,N_17682,N_17281);
nor U19963 (N_19963,N_17506,N_16074);
or U19964 (N_19964,N_16563,N_17518);
nor U19965 (N_19965,N_16561,N_17072);
and U19966 (N_19966,N_17174,N_17007);
nor U19967 (N_19967,N_16687,N_16357);
or U19968 (N_19968,N_16363,N_17988);
xnor U19969 (N_19969,N_17441,N_16346);
and U19970 (N_19970,N_17693,N_17273);
and U19971 (N_19971,N_16835,N_17274);
or U19972 (N_19972,N_17388,N_17912);
and U19973 (N_19973,N_16224,N_16756);
nand U19974 (N_19974,N_16852,N_16182);
or U19975 (N_19975,N_16990,N_16605);
nand U19976 (N_19976,N_16598,N_16682);
nand U19977 (N_19977,N_16839,N_16496);
or U19978 (N_19978,N_16874,N_17882);
or U19979 (N_19979,N_17772,N_16402);
or U19980 (N_19980,N_16807,N_17288);
or U19981 (N_19981,N_17250,N_16466);
xor U19982 (N_19982,N_17017,N_17737);
nand U19983 (N_19983,N_17848,N_17731);
or U19984 (N_19984,N_17490,N_17523);
or U19985 (N_19985,N_16783,N_17177);
or U19986 (N_19986,N_17483,N_16199);
xor U19987 (N_19987,N_17752,N_16384);
or U19988 (N_19988,N_17416,N_16710);
and U19989 (N_19989,N_17822,N_16480);
or U19990 (N_19990,N_17626,N_17547);
and U19991 (N_19991,N_16656,N_17921);
and U19992 (N_19992,N_16544,N_17619);
and U19993 (N_19993,N_17414,N_17857);
or U19994 (N_19994,N_16169,N_17460);
nand U19995 (N_19995,N_17248,N_17620);
or U19996 (N_19996,N_16359,N_16564);
and U19997 (N_19997,N_17278,N_17900);
or U19998 (N_19998,N_17749,N_17687);
nor U19999 (N_19999,N_16480,N_16236);
nor UO_0 (O_0,N_19624,N_18267);
xnor UO_1 (O_1,N_18105,N_19644);
nor UO_2 (O_2,N_18152,N_19241);
nand UO_3 (O_3,N_18485,N_18935);
nand UO_4 (O_4,N_18753,N_18334);
nor UO_5 (O_5,N_18398,N_18986);
or UO_6 (O_6,N_18900,N_19317);
nor UO_7 (O_7,N_18418,N_19980);
and UO_8 (O_8,N_19877,N_19627);
xor UO_9 (O_9,N_19991,N_18716);
or UO_10 (O_10,N_19947,N_19708);
or UO_11 (O_11,N_18280,N_19550);
nand UO_12 (O_12,N_18841,N_18144);
and UO_13 (O_13,N_18588,N_19191);
xnor UO_14 (O_14,N_19066,N_19019);
nand UO_15 (O_15,N_19999,N_18960);
nand UO_16 (O_16,N_19207,N_18168);
nand UO_17 (O_17,N_18577,N_19400);
xor UO_18 (O_18,N_18374,N_18030);
or UO_19 (O_19,N_18563,N_18145);
and UO_20 (O_20,N_18958,N_18008);
or UO_21 (O_21,N_19145,N_18993);
nand UO_22 (O_22,N_18221,N_19985);
nor UO_23 (O_23,N_18681,N_19628);
nand UO_24 (O_24,N_18430,N_19919);
xor UO_25 (O_25,N_18165,N_19106);
xor UO_26 (O_26,N_19322,N_19717);
nor UO_27 (O_27,N_18099,N_18747);
nand UO_28 (O_28,N_19170,N_19719);
and UO_29 (O_29,N_18862,N_18797);
or UO_30 (O_30,N_18112,N_18714);
nor UO_31 (O_31,N_18414,N_19753);
nor UO_32 (O_32,N_19871,N_18306);
xor UO_33 (O_33,N_18157,N_18452);
nand UO_34 (O_34,N_18939,N_18799);
nor UO_35 (O_35,N_18938,N_19598);
nand UO_36 (O_36,N_19101,N_19950);
and UO_37 (O_37,N_19316,N_18239);
and UO_38 (O_38,N_19928,N_18863);
nand UO_39 (O_39,N_18096,N_19039);
xor UO_40 (O_40,N_19920,N_19357);
nor UO_41 (O_41,N_18216,N_18825);
nand UO_42 (O_42,N_19164,N_18219);
nor UO_43 (O_43,N_18416,N_19970);
xor UO_44 (O_44,N_19132,N_19288);
and UO_45 (O_45,N_18864,N_18609);
xor UO_46 (O_46,N_18730,N_19802);
and UO_47 (O_47,N_19757,N_18352);
nand UO_48 (O_48,N_19245,N_18164);
or UO_49 (O_49,N_18220,N_18976);
or UO_50 (O_50,N_19833,N_19477);
or UO_51 (O_51,N_19792,N_18394);
xor UO_52 (O_52,N_18372,N_18495);
nand UO_53 (O_53,N_18957,N_19325);
xnor UO_54 (O_54,N_18576,N_19058);
and UO_55 (O_55,N_18916,N_18901);
and UO_56 (O_56,N_19309,N_18843);
or UO_57 (O_57,N_18003,N_18400);
or UO_58 (O_58,N_18422,N_19760);
nand UO_59 (O_59,N_19895,N_18455);
or UO_60 (O_60,N_19275,N_18535);
xnor UO_61 (O_61,N_18579,N_18460);
or UO_62 (O_62,N_18290,N_19763);
and UO_63 (O_63,N_18572,N_19825);
or UO_64 (O_64,N_19687,N_18650);
nor UO_65 (O_65,N_18189,N_19829);
and UO_66 (O_66,N_19846,N_19018);
or UO_67 (O_67,N_19184,N_19027);
nor UO_68 (O_68,N_18929,N_19501);
or UO_69 (O_69,N_19386,N_19777);
nand UO_70 (O_70,N_19102,N_19848);
nor UO_71 (O_71,N_19755,N_19218);
nand UO_72 (O_72,N_19032,N_18540);
nor UO_73 (O_73,N_19674,N_19390);
nand UO_74 (O_74,N_19479,N_18432);
nand UO_75 (O_75,N_19087,N_19989);
xnor UO_76 (O_76,N_19748,N_19124);
xnor UO_77 (O_77,N_19197,N_18885);
nand UO_78 (O_78,N_19650,N_18312);
xnor UO_79 (O_79,N_19817,N_19455);
and UO_80 (O_80,N_18234,N_18982);
or UO_81 (O_81,N_18205,N_18971);
or UO_82 (O_82,N_18440,N_19125);
and UO_83 (O_83,N_19751,N_18243);
xor UO_84 (O_84,N_18270,N_18343);
or UO_85 (O_85,N_19156,N_19348);
and UO_86 (O_86,N_19403,N_18402);
and UO_87 (O_87,N_19744,N_18437);
or UO_88 (O_88,N_18025,N_18151);
and UO_89 (O_89,N_19352,N_19045);
or UO_90 (O_90,N_19063,N_18693);
nor UO_91 (O_91,N_19503,N_18685);
or UO_92 (O_92,N_19508,N_19269);
and UO_93 (O_93,N_19319,N_19556);
and UO_94 (O_94,N_18710,N_19810);
or UO_95 (O_95,N_19169,N_19922);
nor UO_96 (O_96,N_18072,N_19535);
nor UO_97 (O_97,N_18889,N_19399);
or UO_98 (O_98,N_18739,N_18257);
nor UO_99 (O_99,N_19016,N_19375);
or UO_100 (O_100,N_18664,N_18984);
and UO_101 (O_101,N_18170,N_19559);
or UO_102 (O_102,N_19187,N_19144);
nand UO_103 (O_103,N_19362,N_19216);
nand UO_104 (O_104,N_19704,N_19858);
or UO_105 (O_105,N_19179,N_19664);
or UO_106 (O_106,N_18926,N_19140);
nand UO_107 (O_107,N_19213,N_18904);
xnor UO_108 (O_108,N_18148,N_18052);
and UO_109 (O_109,N_19982,N_18087);
nand UO_110 (O_110,N_18210,N_18264);
nand UO_111 (O_111,N_19294,N_18631);
nand UO_112 (O_112,N_19521,N_19229);
xnor UO_113 (O_113,N_18712,N_19026);
xnor UO_114 (O_114,N_19017,N_19461);
and UO_115 (O_115,N_18829,N_19192);
and UO_116 (O_116,N_18659,N_18071);
xnor UO_117 (O_117,N_18750,N_18634);
or UO_118 (O_118,N_19404,N_18925);
and UO_119 (O_119,N_18042,N_18606);
xor UO_120 (O_120,N_18698,N_19849);
and UO_121 (O_121,N_18847,N_18447);
nand UO_122 (O_122,N_19252,N_19996);
or UO_123 (O_123,N_19548,N_18263);
nand UO_124 (O_124,N_19631,N_19803);
or UO_125 (O_125,N_19790,N_18855);
nor UO_126 (O_126,N_19021,N_19932);
xor UO_127 (O_127,N_18842,N_19212);
nor UO_128 (O_128,N_18187,N_19028);
nor UO_129 (O_129,N_18442,N_19617);
nand UO_130 (O_130,N_19366,N_18590);
nand UO_131 (O_131,N_19287,N_18200);
nor UO_132 (O_132,N_19551,N_19733);
nand UO_133 (O_133,N_19234,N_18496);
nor UO_134 (O_134,N_19669,N_19117);
and UO_135 (O_135,N_19129,N_19769);
and UO_136 (O_136,N_19020,N_19844);
nor UO_137 (O_137,N_19202,N_18601);
nand UO_138 (O_138,N_18456,N_18793);
and UO_139 (O_139,N_19707,N_18504);
nand UO_140 (O_140,N_19998,N_19268);
nand UO_141 (O_141,N_18751,N_19797);
nor UO_142 (O_142,N_19861,N_18011);
and UO_143 (O_143,N_19310,N_18537);
nand UO_144 (O_144,N_19343,N_18344);
nor UO_145 (O_145,N_19385,N_18526);
or UO_146 (O_146,N_18467,N_18019);
or UO_147 (O_147,N_18380,N_19429);
or UO_148 (O_148,N_19141,N_18918);
nor UO_149 (O_149,N_19783,N_19110);
nand UO_150 (O_150,N_19804,N_18330);
or UO_151 (O_151,N_19564,N_18992);
and UO_152 (O_152,N_18840,N_18801);
xnor UO_153 (O_153,N_18018,N_18834);
or UO_154 (O_154,N_19055,N_19199);
and UO_155 (O_155,N_19302,N_18283);
and UO_156 (O_156,N_19206,N_18922);
nor UO_157 (O_157,N_19166,N_18819);
nor UO_158 (O_158,N_19887,N_19577);
nor UO_159 (O_159,N_18788,N_19281);
and UO_160 (O_160,N_19115,N_18644);
and UO_161 (O_161,N_18106,N_19839);
xor UO_162 (O_162,N_19364,N_19636);
nor UO_163 (O_163,N_18180,N_18009);
nand UO_164 (O_164,N_19023,N_18636);
nand UO_165 (O_165,N_18082,N_18331);
and UO_166 (O_166,N_18176,N_18907);
and UO_167 (O_167,N_18779,N_19258);
nor UO_168 (O_168,N_18622,N_19370);
nor UO_169 (O_169,N_18552,N_19040);
nand UO_170 (O_170,N_18014,N_18530);
and UO_171 (O_171,N_18230,N_18359);
xnor UO_172 (O_172,N_18109,N_19750);
xor UO_173 (O_173,N_19711,N_18260);
or UO_174 (O_174,N_19138,N_18120);
xnor UO_175 (O_175,N_18208,N_18651);
nor UO_176 (O_176,N_18272,N_18034);
nand UO_177 (O_177,N_19558,N_18369);
nand UO_178 (O_178,N_19318,N_19189);
nor UO_179 (O_179,N_18684,N_19057);
nand UO_180 (O_180,N_18241,N_18502);
or UO_181 (O_181,N_19091,N_19933);
nand UO_182 (O_182,N_19464,N_19897);
nor UO_183 (O_183,N_18893,N_19475);
nand UO_184 (O_184,N_19183,N_18229);
and UO_185 (O_185,N_19542,N_19648);
or UO_186 (O_186,N_19034,N_19690);
and UO_187 (O_187,N_19038,N_19538);
or UO_188 (O_188,N_19705,N_19983);
nand UO_189 (O_189,N_19340,N_19754);
xor UO_190 (O_190,N_19271,N_18253);
nand UO_191 (O_191,N_18817,N_18131);
and UO_192 (O_192,N_19824,N_19360);
nor UO_193 (O_193,N_19620,N_18875);
and UO_194 (O_194,N_19075,N_19356);
nand UO_195 (O_195,N_19250,N_19642);
and UO_196 (O_196,N_19693,N_18118);
and UO_197 (O_197,N_19766,N_19762);
nand UO_198 (O_198,N_19159,N_18068);
or UO_199 (O_199,N_18757,N_18608);
and UO_200 (O_200,N_18408,N_19622);
or UO_201 (O_201,N_19579,N_19767);
or UO_202 (O_202,N_19863,N_18020);
nand UO_203 (O_203,N_18409,N_18128);
nand UO_204 (O_204,N_19435,N_19675);
or UO_205 (O_205,N_19379,N_18902);
xor UO_206 (O_206,N_19300,N_18655);
or UO_207 (O_207,N_19473,N_19181);
or UO_208 (O_208,N_18340,N_18026);
nor UO_209 (O_209,N_19296,N_18326);
or UO_210 (O_210,N_18878,N_18173);
and UO_211 (O_211,N_18356,N_18881);
xnor UO_212 (O_212,N_18249,N_18484);
and UO_213 (O_213,N_18110,N_19489);
and UO_214 (O_214,N_18813,N_18679);
nor UO_215 (O_215,N_19255,N_18182);
nand UO_216 (O_216,N_19806,N_18259);
nor UO_217 (O_217,N_18091,N_19314);
nand UO_218 (O_218,N_18621,N_18088);
xor UO_219 (O_219,N_18669,N_19634);
nand UO_220 (O_220,N_19328,N_18930);
nand UO_221 (O_221,N_18764,N_18532);
or UO_222 (O_222,N_19517,N_19505);
nor UO_223 (O_223,N_18490,N_19772);
xnor UO_224 (O_224,N_18574,N_19198);
nor UO_225 (O_225,N_18955,N_18748);
nand UO_226 (O_226,N_18420,N_19632);
or UO_227 (O_227,N_18245,N_18472);
nand UO_228 (O_228,N_18541,N_18001);
nand UO_229 (O_229,N_19469,N_18171);
or UO_230 (O_230,N_18016,N_18097);
nand UO_231 (O_231,N_19257,N_18774);
and UO_232 (O_232,N_18232,N_19222);
or UO_233 (O_233,N_18479,N_18617);
and UO_234 (O_234,N_18972,N_19085);
nand UO_235 (O_235,N_18752,N_18155);
nor UO_236 (O_236,N_18375,N_18589);
and UO_237 (O_237,N_19937,N_19789);
and UO_238 (O_238,N_19780,N_19731);
nor UO_239 (O_239,N_18564,N_19941);
and UO_240 (O_240,N_18293,N_19714);
nand UO_241 (O_241,N_18395,N_19527);
or UO_242 (O_242,N_18592,N_18523);
nand UO_243 (O_243,N_19478,N_19420);
nand UO_244 (O_244,N_18027,N_19363);
xor UO_245 (O_245,N_19158,N_18427);
or UO_246 (O_246,N_19977,N_18159);
nand UO_247 (O_247,N_18199,N_19807);
nor UO_248 (O_248,N_18554,N_19630);
nand UO_249 (O_249,N_18510,N_18158);
or UO_250 (O_250,N_19436,N_18836);
and UO_251 (O_251,N_19580,N_19217);
and UO_252 (O_252,N_19889,N_19280);
nor UO_253 (O_253,N_18499,N_19745);
xnor UO_254 (O_254,N_18154,N_19080);
nand UO_255 (O_255,N_18401,N_19872);
nor UO_256 (O_256,N_19532,N_19912);
xor UO_257 (O_257,N_18461,N_19666);
nand UO_258 (O_258,N_19741,N_18419);
and UO_259 (O_259,N_19326,N_18193);
nor UO_260 (O_260,N_18879,N_19694);
and UO_261 (O_261,N_18141,N_19393);
nor UO_262 (O_262,N_18130,N_18524);
nand UO_263 (O_263,N_18913,N_19232);
nor UO_264 (O_264,N_19852,N_19530);
xnor UO_265 (O_265,N_19367,N_19938);
nor UO_266 (O_266,N_19112,N_19312);
and UO_267 (O_267,N_19226,N_19729);
and UO_268 (O_268,N_19842,N_18873);
nand UO_269 (O_269,N_19256,N_19108);
nor UO_270 (O_270,N_18791,N_19832);
nor UO_271 (O_271,N_18543,N_19380);
or UO_272 (O_272,N_18464,N_18877);
or UO_273 (O_273,N_18040,N_18597);
nand UO_274 (O_274,N_18423,N_18119);
nand UO_275 (O_275,N_18772,N_18818);
and UO_276 (O_276,N_19174,N_19796);
nand UO_277 (O_277,N_19595,N_19820);
or UO_278 (O_278,N_18487,N_19692);
and UO_279 (O_279,N_19487,N_18048);
and UO_280 (O_280,N_19452,N_19361);
or UO_281 (O_281,N_19458,N_18161);
nand UO_282 (O_282,N_18188,N_19954);
nor UO_283 (O_283,N_18575,N_19917);
or UO_284 (O_284,N_18546,N_19210);
xor UO_285 (O_285,N_18251,N_19531);
and UO_286 (O_286,N_18560,N_19481);
or UO_287 (O_287,N_19981,N_19702);
nor UO_288 (O_288,N_19180,N_19637);
and UO_289 (O_289,N_18392,N_19134);
xor UO_290 (O_290,N_19022,N_18318);
or UO_291 (O_291,N_19495,N_19406);
or UO_292 (O_292,N_19685,N_19960);
xnor UO_293 (O_293,N_18620,N_19823);
nor UO_294 (O_294,N_18827,N_18246);
or UO_295 (O_295,N_19862,N_18429);
nor UO_296 (O_296,N_18682,N_18613);
or UO_297 (O_297,N_18433,N_19143);
or UO_298 (O_298,N_18782,N_18800);
xor UO_299 (O_299,N_19378,N_19907);
or UO_300 (O_300,N_18185,N_19573);
xor UO_301 (O_301,N_18022,N_19446);
nor UO_302 (O_302,N_18652,N_19486);
or UO_303 (O_303,N_18921,N_18727);
nand UO_304 (O_304,N_18327,N_18905);
xor UO_305 (O_305,N_19683,N_18874);
and UO_306 (O_306,N_18458,N_18163);
and UO_307 (O_307,N_19060,N_19740);
xor UO_308 (O_308,N_19453,N_19279);
nor UO_309 (O_309,N_18421,N_18987);
nor UO_310 (O_310,N_18985,N_19405);
and UO_311 (O_311,N_19968,N_19805);
or UO_312 (O_312,N_19868,N_18903);
nand UO_313 (O_313,N_19249,N_19522);
or UO_314 (O_314,N_19539,N_19801);
xor UO_315 (O_315,N_19493,N_19335);
nand UO_316 (O_316,N_19883,N_18697);
or UO_317 (O_317,N_19044,N_18288);
and UO_318 (O_318,N_19761,N_19261);
xor UO_319 (O_319,N_19082,N_19822);
or UO_320 (O_320,N_19944,N_18102);
xnor UO_321 (O_321,N_19866,N_19052);
nand UO_322 (O_322,N_18990,N_19195);
or UO_323 (O_323,N_18630,N_18505);
and UO_324 (O_324,N_18528,N_18517);
and UO_325 (O_325,N_18337,N_19787);
and UO_326 (O_326,N_18302,N_18122);
and UO_327 (O_327,N_18067,N_19840);
nand UO_328 (O_328,N_18107,N_18624);
or UO_329 (O_329,N_19643,N_18196);
nor UO_330 (O_330,N_18722,N_19609);
and UO_331 (O_331,N_19054,N_18483);
or UO_332 (O_332,N_19553,N_19886);
or UO_333 (O_333,N_19788,N_19209);
nand UO_334 (O_334,N_19472,N_19836);
nor UO_335 (O_335,N_19738,N_18133);
nor UO_336 (O_336,N_18850,N_18226);
and UO_337 (O_337,N_18217,N_18694);
nand UO_338 (O_338,N_18339,N_19875);
or UO_339 (O_339,N_19163,N_18053);
and UO_340 (O_340,N_18470,N_18041);
xor UO_341 (O_341,N_18095,N_19888);
and UO_342 (O_342,N_18671,N_18775);
nor UO_343 (O_343,N_18043,N_18077);
nor UO_344 (O_344,N_19572,N_19333);
nor UO_345 (O_345,N_19071,N_19396);
xor UO_346 (O_346,N_19086,N_19838);
nor UO_347 (O_347,N_19172,N_18397);
xnor UO_348 (O_348,N_19419,N_18376);
and UO_349 (O_349,N_19515,N_19597);
nand UO_350 (O_350,N_18811,N_19306);
and UO_351 (O_351,N_18810,N_19381);
nand UO_352 (O_352,N_19905,N_19953);
or UO_353 (O_353,N_18600,N_18323);
nand UO_354 (O_354,N_19149,N_19392);
or UO_355 (O_355,N_19915,N_18305);
and UO_356 (O_356,N_19560,N_19388);
and UO_357 (O_357,N_19518,N_18688);
and UO_358 (O_358,N_19646,N_19682);
and UO_359 (O_359,N_18462,N_18478);
nor UO_360 (O_360,N_19695,N_18941);
or UO_361 (O_361,N_18177,N_18521);
nand UO_362 (O_362,N_18911,N_19710);
nor UO_363 (O_363,N_19662,N_19847);
nor UO_364 (O_364,N_19677,N_19881);
or UO_365 (O_365,N_19655,N_18645);
nand UO_366 (O_366,N_18435,N_18709);
nand UO_367 (O_367,N_18227,N_19430);
and UO_368 (O_368,N_18127,N_18508);
nor UO_369 (O_369,N_19334,N_18762);
nand UO_370 (O_370,N_19010,N_19373);
or UO_371 (O_371,N_18968,N_19809);
nor UO_372 (O_372,N_19421,N_18950);
and UO_373 (O_373,N_19483,N_19774);
nand UO_374 (O_374,N_19735,N_18247);
or UO_375 (O_375,N_18823,N_19602);
nand UO_376 (O_376,N_18673,N_19074);
nor UO_377 (O_377,N_19526,N_18197);
nand UO_378 (O_378,N_19504,N_18884);
nand UO_379 (O_379,N_19752,N_19387);
or UO_380 (O_380,N_19200,N_18770);
nand UO_381 (O_381,N_19837,N_19908);
nor UO_382 (O_382,N_18755,N_18399);
nor UO_383 (O_383,N_19676,N_19921);
and UO_384 (O_384,N_18861,N_19194);
nand UO_385 (O_385,N_18733,N_19005);
nor UO_386 (O_386,N_19147,N_18568);
or UO_387 (O_387,N_19476,N_19537);
or UO_388 (O_388,N_18999,N_18277);
nor UO_389 (O_389,N_19460,N_18663);
and UO_390 (O_390,N_18013,N_19165);
and UO_391 (O_391,N_19499,N_18284);
or UO_392 (O_392,N_18776,N_18927);
nor UO_393 (O_393,N_18045,N_18648);
nor UO_394 (O_394,N_19984,N_18509);
and UO_395 (O_395,N_19377,N_19128);
nand UO_396 (O_396,N_18953,N_19700);
nor UO_397 (O_397,N_18482,N_19480);
and UO_398 (O_398,N_19465,N_18808);
and UO_399 (O_399,N_19699,N_19546);
nand UO_400 (O_400,N_19013,N_18743);
and UO_401 (O_401,N_18010,N_19555);
nor UO_402 (O_402,N_19509,N_18285);
nor UO_403 (O_403,N_19819,N_18691);
xnor UO_404 (O_404,N_19047,N_18179);
and UO_405 (O_405,N_19413,N_18868);
nand UO_406 (O_406,N_19374,N_19976);
nand UO_407 (O_407,N_18599,N_19437);
or UO_408 (O_408,N_18281,N_19732);
or UO_409 (O_409,N_18700,N_19168);
and UO_410 (O_410,N_19860,N_18769);
and UO_411 (O_411,N_18704,N_19657);
or UO_412 (O_412,N_18718,N_18357);
or UO_413 (O_413,N_18493,N_19898);
or UO_414 (O_414,N_19089,N_18591);
and UO_415 (O_415,N_18598,N_18135);
nand UO_416 (O_416,N_18821,N_18844);
nand UO_417 (O_417,N_19845,N_18974);
nand UO_418 (O_418,N_18500,N_19408);
and UO_419 (O_419,N_19350,N_18551);
nand UO_420 (O_420,N_18961,N_18956);
or UO_421 (O_421,N_19069,N_18728);
xor UO_422 (O_422,N_19812,N_18086);
nor UO_423 (O_423,N_19974,N_19625);
xor UO_424 (O_424,N_18345,N_18846);
and UO_425 (O_425,N_19791,N_19282);
and UO_426 (O_426,N_18996,N_18944);
nand UO_427 (O_427,N_18906,N_18289);
nand UO_428 (O_428,N_18428,N_18760);
or UO_429 (O_429,N_19581,N_19899);
nand UO_430 (O_430,N_19092,N_18705);
nor UO_431 (O_431,N_19177,N_19094);
or UO_432 (O_432,N_18307,N_19656);
and UO_433 (O_433,N_19447,N_18054);
or UO_434 (O_434,N_18471,N_19449);
nand UO_435 (O_435,N_18894,N_18824);
or UO_436 (O_436,N_19185,N_19545);
nor UO_437 (O_437,N_18124,N_18434);
and UO_438 (O_438,N_18798,N_19369);
nand UO_439 (O_439,N_18108,N_18237);
nor UO_440 (O_440,N_19633,N_18181);
and UO_441 (O_441,N_18963,N_19304);
or UO_442 (O_442,N_18732,N_19186);
nor UO_443 (O_443,N_18544,N_18256);
nand UO_444 (O_444,N_19412,N_19652);
nand UO_445 (O_445,N_18058,N_19994);
or UO_446 (O_446,N_18450,N_19301);
nand UO_447 (O_447,N_19104,N_18269);
nor UO_448 (O_448,N_18023,N_19415);
nor UO_449 (O_449,N_19418,N_19488);
nand UO_450 (O_450,N_18550,N_19036);
nand UO_451 (O_451,N_19389,N_19441);
or UO_452 (O_452,N_18790,N_18852);
or UO_453 (O_453,N_18366,N_19709);
or UO_454 (O_454,N_18300,N_18931);
and UO_455 (O_455,N_18585,N_19339);
or UO_456 (O_456,N_19660,N_18211);
and UO_457 (O_457,N_19720,N_19874);
nor UO_458 (O_458,N_19414,N_18514);
or UO_459 (O_459,N_19613,N_19629);
nand UO_460 (O_460,N_19703,N_18276);
nor UO_461 (O_461,N_19240,N_18379);
nand UO_462 (O_462,N_19397,N_19337);
nor UO_463 (O_463,N_18898,N_19965);
xor UO_464 (O_464,N_19457,N_19482);
nor UO_465 (O_465,N_18275,N_18194);
and UO_466 (O_466,N_18024,N_18677);
and UO_467 (O_467,N_19997,N_18153);
nand UO_468 (O_468,N_19943,N_19030);
or UO_469 (O_469,N_18268,N_19565);
nor UO_470 (O_470,N_19203,N_19891);
nor UO_471 (O_471,N_18315,N_18804);
nor UO_472 (O_472,N_19879,N_18890);
nor UO_473 (O_473,N_19076,N_18166);
or UO_474 (O_474,N_19680,N_18384);
and UO_475 (O_475,N_19583,N_18362);
nand UO_476 (O_476,N_19211,N_18977);
nor UO_477 (O_477,N_18954,N_19594);
nor UO_478 (O_478,N_18547,N_18527);
nand UO_479 (O_479,N_19315,N_19885);
nor UO_480 (O_480,N_19893,N_19127);
nor UO_481 (O_481,N_18069,N_18492);
nor UO_482 (O_482,N_18582,N_18571);
nand UO_483 (O_483,N_19113,N_18035);
nor UO_484 (O_484,N_19121,N_19549);
and UO_485 (O_485,N_18477,N_18596);
or UO_486 (O_486,N_18914,N_19067);
or UO_487 (O_487,N_19064,N_18413);
nand UO_488 (O_488,N_19365,N_18883);
or UO_489 (O_489,N_18676,N_18468);
nand UO_490 (O_490,N_18474,N_19585);
and UO_491 (O_491,N_18311,N_19940);
nand UO_492 (O_492,N_18191,N_19041);
or UO_493 (O_493,N_19118,N_19230);
and UO_494 (O_494,N_18796,N_18876);
and UO_495 (O_495,N_19284,N_18007);
or UO_496 (O_496,N_19519,N_18389);
xnor UO_497 (O_497,N_18887,N_19821);
and UO_498 (O_498,N_18126,N_19313);
and UO_499 (O_499,N_18335,N_18933);
nand UO_500 (O_500,N_18192,N_19649);
and UO_501 (O_501,N_18602,N_18132);
nand UO_502 (O_502,N_18578,N_18888);
nand UO_503 (O_503,N_18431,N_18316);
nor UO_504 (O_504,N_18417,N_18851);
and UO_505 (O_505,N_18329,N_18279);
nor UO_506 (O_506,N_18489,N_18573);
and UO_507 (O_507,N_18235,N_18962);
xnor UO_508 (O_508,N_19721,N_18129);
and UO_509 (O_509,N_18425,N_18101);
or UO_510 (O_510,N_18396,N_18480);
and UO_511 (O_511,N_19081,N_19093);
nand UO_512 (O_512,N_18081,N_18565);
or UO_513 (O_513,N_18250,N_19969);
nand UO_514 (O_514,N_19894,N_18539);
or UO_515 (O_515,N_18642,N_18794);
nand UO_516 (O_516,N_18294,N_19610);
xor UO_517 (O_517,N_18076,N_18463);
nand UO_518 (O_518,N_19835,N_18353);
nor UO_519 (O_519,N_19554,N_19114);
nand UO_520 (O_520,N_19424,N_18966);
nand UO_521 (O_521,N_18780,N_19496);
nand UO_522 (O_522,N_18032,N_18661);
and UO_523 (O_523,N_18498,N_19658);
nand UO_524 (O_524,N_18777,N_19090);
and UO_525 (O_525,N_19971,N_18328);
xor UO_526 (O_526,N_18178,N_19758);
or UO_527 (O_527,N_18839,N_18637);
and UO_528 (O_528,N_19247,N_18321);
nand UO_529 (O_529,N_18497,N_19000);
and UO_530 (O_530,N_19528,N_18789);
xnor UO_531 (O_531,N_19474,N_18857);
nand UO_532 (O_532,N_19150,N_19135);
xor UO_533 (O_533,N_18997,N_19670);
and UO_534 (O_534,N_18632,N_19914);
nand UO_535 (O_535,N_19608,N_18454);
xor UO_536 (O_536,N_19736,N_18717);
nand UO_537 (O_537,N_19043,N_18981);
and UO_538 (O_538,N_18292,N_18570);
nor UO_539 (O_539,N_18448,N_19193);
xnor UO_540 (O_540,N_19428,N_18908);
nand UO_541 (O_541,N_19471,N_18970);
or UO_542 (O_542,N_19966,N_18723);
or UO_543 (O_543,N_18856,N_18618);
nor UO_544 (O_544,N_19401,N_18869);
and UO_545 (O_545,N_18299,N_19663);
or UO_546 (O_546,N_19841,N_18657);
xor UO_547 (O_547,N_19952,N_18529);
or UO_548 (O_548,N_19228,N_19342);
and UO_549 (O_549,N_18545,N_19688);
or UO_550 (O_550,N_19239,N_18218);
or UO_551 (O_551,N_18021,N_18265);
nand UO_552 (O_552,N_18365,N_18858);
and UO_553 (O_553,N_18093,N_19065);
and UO_554 (O_554,N_19492,N_18503);
or UO_555 (O_555,N_19934,N_18703);
or UO_556 (O_556,N_18314,N_19718);
and UO_557 (O_557,N_19451,N_18767);
or UO_558 (O_558,N_19723,N_19990);
or UO_559 (O_559,N_18886,N_19095);
nand UO_560 (O_560,N_18342,N_19376);
nand UO_561 (O_561,N_19267,N_19502);
nor UO_562 (O_562,N_19524,N_18140);
and UO_563 (O_563,N_19830,N_18946);
xor UO_564 (O_564,N_19715,N_19726);
nand UO_565 (O_565,N_19238,N_19615);
nand UO_566 (O_566,N_19859,N_19619);
nand UO_567 (O_567,N_18803,N_19248);
or UO_568 (O_568,N_18763,N_18046);
xor UO_569 (O_569,N_18920,N_18382);
nor UO_570 (O_570,N_18724,N_18715);
and UO_571 (O_571,N_19568,N_19099);
nor UO_572 (O_572,N_19167,N_19563);
or UO_573 (O_573,N_18765,N_18203);
and UO_574 (O_574,N_19616,N_19870);
and UO_575 (O_575,N_18457,N_18802);
nor UO_576 (O_576,N_18333,N_18988);
nor UO_577 (O_577,N_18297,N_18786);
and UO_578 (O_578,N_19208,N_19768);
nand UO_579 (O_579,N_19259,N_19109);
xnor UO_580 (O_580,N_18809,N_18518);
or UO_581 (O_581,N_18084,N_18006);
and UO_582 (O_582,N_18731,N_19426);
xor UO_583 (O_583,N_18860,N_19993);
xor UO_584 (O_584,N_19463,N_19440);
or UO_585 (O_585,N_18261,N_18945);
xor UO_586 (O_586,N_18228,N_18542);
nor UO_587 (O_587,N_19586,N_19697);
nand UO_588 (O_588,N_19146,N_19442);
nand UO_589 (O_589,N_19773,N_18947);
xor UO_590 (O_590,N_18866,N_19407);
and UO_591 (O_591,N_19864,N_19347);
and UO_592 (O_592,N_19225,N_18360);
and UO_593 (O_593,N_19588,N_18626);
nand UO_594 (O_594,N_18057,N_19264);
nand UO_595 (O_595,N_18744,N_18346);
and UO_596 (O_596,N_19025,N_19851);
nor UO_597 (O_597,N_18737,N_19794);
nand UO_598 (O_598,N_19679,N_19651);
nand UO_599 (O_599,N_18473,N_18160);
xor UO_600 (O_600,N_18038,N_19084);
or UO_601 (O_601,N_18405,N_19285);
or UO_602 (O_602,N_19297,N_18680);
and UO_603 (O_603,N_19765,N_19684);
and UO_604 (O_604,N_18867,N_18361);
nor UO_605 (O_605,N_18494,N_19635);
nand UO_606 (O_606,N_18167,N_18262);
nand UO_607 (O_607,N_18978,N_19311);
nand UO_608 (O_608,N_19979,N_18699);
and UO_609 (O_609,N_18089,N_18002);
or UO_610 (O_610,N_18004,N_19730);
nor UO_611 (O_611,N_19265,N_19278);
nor UO_612 (O_612,N_19584,N_19223);
xnor UO_613 (O_613,N_18139,N_19798);
or UO_614 (O_614,N_18951,N_19884);
nor UO_615 (O_615,N_18363,N_19432);
and UO_616 (O_616,N_19614,N_18548);
nor UO_617 (O_617,N_18792,N_19048);
or UO_618 (O_618,N_19541,N_19438);
xor UO_619 (O_619,N_19592,N_19799);
or UO_620 (O_620,N_19959,N_19330);
xnor UO_621 (O_621,N_19698,N_19951);
xnor UO_622 (O_622,N_18146,N_19749);
or UO_623 (O_623,N_19254,N_19273);
nor UO_624 (O_624,N_19828,N_19712);
or UO_625 (O_625,N_18062,N_19681);
nor UO_626 (O_626,N_19498,N_19004);
nand UO_627 (O_627,N_19910,N_18441);
or UO_628 (O_628,N_18936,N_18520);
and UO_629 (O_629,N_18134,N_18795);
or UO_630 (O_630,N_18892,N_19778);
xor UO_631 (O_631,N_18781,N_19640);
xor UO_632 (O_632,N_18662,N_19272);
and UO_633 (O_633,N_18721,N_18686);
and UO_634 (O_634,N_18449,N_18895);
or UO_635 (O_635,N_18853,N_18967);
and UO_636 (O_636,N_19507,N_18942);
nor UO_637 (O_637,N_18561,N_19439);
nor UO_638 (O_638,N_18633,N_18627);
or UO_639 (O_639,N_18103,N_19942);
nor UO_640 (O_640,N_19024,N_19484);
and UO_641 (O_641,N_18629,N_18183);
nand UO_642 (O_642,N_18481,N_18531);
nand UO_643 (O_643,N_18117,N_18643);
nand UO_644 (O_644,N_18015,N_18604);
and UO_645 (O_645,N_18092,N_19260);
nand UO_646 (O_646,N_19151,N_19882);
or UO_647 (O_647,N_19596,N_18949);
and UO_648 (O_648,N_18121,N_19547);
nor UO_649 (O_649,N_19987,N_18443);
or UO_650 (O_650,N_18501,N_19814);
nor UO_651 (O_651,N_19611,N_18212);
or UO_652 (O_652,N_19188,N_18989);
and UO_653 (O_653,N_18784,N_18924);
nor UO_654 (O_654,N_19050,N_18534);
and UO_655 (O_655,N_18224,N_19665);
or UO_656 (O_656,N_19756,N_18031);
nand UO_657 (O_657,N_19911,N_18934);
nand UO_658 (O_658,N_19470,N_19062);
xnor UO_659 (O_659,N_19701,N_19345);
nand UO_660 (O_660,N_18538,N_18513);
or UO_661 (O_661,N_18298,N_18583);
or UO_662 (O_662,N_19601,N_18309);
nor UO_663 (O_663,N_18845,N_18386);
nor UO_664 (O_664,N_18085,N_18998);
xor UO_665 (O_665,N_18355,N_19800);
nor UO_666 (O_666,N_18675,N_18778);
or UO_667 (O_667,N_18388,N_19963);
nor UO_668 (O_668,N_19672,N_19382);
and UO_669 (O_669,N_18507,N_18274);
nor UO_670 (O_670,N_19536,N_19713);
and UO_671 (O_671,N_18735,N_19160);
nor UO_672 (O_672,N_19737,N_19119);
and UO_673 (O_673,N_19575,N_18415);
nor UO_674 (O_674,N_18184,N_18668);
and UO_675 (O_675,N_18713,N_19371);
nand UO_676 (O_676,N_18113,N_19626);
or UO_677 (O_677,N_19001,N_18766);
or UO_678 (O_678,N_18351,N_18815);
or UO_679 (O_679,N_19283,N_18201);
nor UO_680 (O_680,N_19227,N_18658);
or UO_681 (O_681,N_18749,N_19014);
or UO_682 (O_682,N_19638,N_19604);
or UO_683 (O_683,N_18348,N_19603);
nor UO_684 (O_684,N_18785,N_19880);
nand UO_685 (O_685,N_19173,N_19571);
and UO_686 (O_686,N_18653,N_18061);
nor UO_687 (O_687,N_19253,N_19321);
nor UO_688 (O_688,N_19368,N_19243);
and UO_689 (O_689,N_18116,N_18783);
or UO_690 (O_690,N_19949,N_18320);
nor UO_691 (O_691,N_19097,N_18407);
nor UO_692 (O_692,N_19834,N_18910);
and UO_693 (O_693,N_19853,N_18980);
nor UO_694 (O_694,N_19423,N_19511);
and UO_695 (O_695,N_19154,N_18258);
nand UO_696 (O_696,N_19009,N_18254);
or UO_697 (O_697,N_18142,N_18486);
and UO_698 (O_698,N_19290,N_19231);
and UO_699 (O_699,N_19896,N_19002);
nor UO_700 (O_700,N_18341,N_18896);
nand UO_701 (O_701,N_18640,N_19576);
and UO_702 (O_702,N_18665,N_18738);
or UO_703 (O_703,N_18325,N_19037);
or UO_704 (O_704,N_18138,N_18696);
and UO_705 (O_705,N_18169,N_19878);
nand UO_706 (O_706,N_18317,N_19490);
nand UO_707 (O_707,N_18952,N_19291);
and UO_708 (O_708,N_18319,N_19667);
nor UO_709 (O_709,N_19759,N_18595);
nor UO_710 (O_710,N_18940,N_18605);
or UO_711 (O_711,N_18580,N_19327);
and UO_712 (O_712,N_18937,N_18702);
or UO_713 (O_713,N_19454,N_19513);
or UO_714 (O_714,N_18029,N_18198);
nand UO_715 (O_715,N_18005,N_19402);
nand UO_716 (O_716,N_18377,N_19190);
or UO_717 (O_717,N_19305,N_19384);
nor UO_718 (O_718,N_19235,N_18973);
and UO_719 (O_719,N_19689,N_18549);
and UO_720 (O_720,N_19372,N_19122);
nand UO_721 (O_721,N_19587,N_18059);
xnor UO_722 (O_722,N_19865,N_18928);
or UO_723 (O_723,N_18516,N_19988);
nand UO_724 (O_724,N_18625,N_18060);
nor UO_725 (O_725,N_19103,N_19175);
nor UO_726 (O_726,N_18286,N_18238);
nor UO_727 (O_727,N_19612,N_19925);
nor UO_728 (O_728,N_19552,N_19236);
nand UO_729 (O_729,N_18725,N_18707);
xnor UO_730 (O_730,N_19107,N_19338);
and UO_731 (O_731,N_18787,N_18623);
and UO_732 (O_732,N_18047,N_18553);
xnor UO_733 (O_733,N_19892,N_18304);
or UO_734 (O_734,N_19332,N_18872);
and UO_735 (O_735,N_19569,N_19843);
nand UO_736 (O_736,N_19341,N_18090);
and UO_737 (O_737,N_18865,N_18063);
or UO_738 (O_738,N_19901,N_19171);
xnor UO_739 (O_739,N_18049,N_18584);
nor UO_740 (O_740,N_19425,N_19456);
nand UO_741 (O_741,N_18364,N_18255);
xor UO_742 (O_742,N_19068,N_18332);
and UO_743 (O_743,N_19678,N_18078);
nand UO_744 (O_744,N_19485,N_19246);
or UO_745 (O_745,N_18436,N_19012);
or UO_746 (O_746,N_18125,N_19274);
nand UO_747 (O_747,N_19540,N_18837);
and UO_748 (O_748,N_19747,N_18701);
and UO_749 (O_749,N_18909,N_18079);
xnor UO_750 (O_750,N_18354,N_18266);
or UO_751 (O_751,N_18943,N_19033);
or UO_752 (O_752,N_19355,N_19153);
or UO_753 (O_753,N_19929,N_18066);
nand UO_754 (O_754,N_19204,N_18206);
nand UO_755 (O_755,N_19599,N_19520);
and UO_756 (O_756,N_19398,N_19764);
and UO_757 (O_757,N_19346,N_19467);
nor UO_758 (O_758,N_18438,N_18073);
nor UO_759 (O_759,N_19641,N_18033);
xor UO_760 (O_760,N_18773,N_19395);
nor UO_761 (O_761,N_18162,N_18562);
or UO_762 (O_762,N_19590,N_19056);
nand UO_763 (O_763,N_18756,N_19042);
nor UO_764 (O_764,N_19410,N_18871);
or UO_765 (O_765,N_19046,N_18612);
nor UO_766 (O_766,N_18759,N_18740);
xor UO_767 (O_767,N_18512,N_18036);
or UO_768 (O_768,N_18816,N_18880);
or UO_769 (O_769,N_18557,N_18322);
and UO_770 (O_770,N_18519,N_18708);
nor UO_771 (O_771,N_19079,N_18581);
nand UO_772 (O_772,N_18959,N_18248);
nand UO_773 (O_773,N_18385,N_18639);
nor UO_774 (O_774,N_18439,N_18805);
nand UO_775 (O_775,N_18174,N_19299);
and UO_776 (O_776,N_18368,N_19434);
nand UO_777 (O_777,N_18424,N_18558);
xnor UO_778 (O_778,N_18635,N_18614);
or UO_779 (O_779,N_18282,N_18336);
xor UO_780 (O_780,N_19433,N_18273);
nand UO_781 (O_781,N_18736,N_19293);
or UO_782 (O_782,N_19645,N_19251);
nand UO_783 (O_783,N_19450,N_18536);
nand UO_784 (O_784,N_18807,N_19725);
or UO_785 (O_785,N_19939,N_19529);
xnor UO_786 (O_786,N_19148,N_19961);
and UO_787 (O_787,N_19059,N_18912);
xnor UO_788 (O_788,N_19739,N_19123);
or UO_789 (O_789,N_19935,N_18603);
or UO_790 (O_790,N_18806,N_18393);
nor UO_791 (O_791,N_18511,N_19722);
nor UO_792 (O_792,N_19262,N_19131);
xor UO_793 (O_793,N_19237,N_18683);
and UO_794 (O_794,N_19409,N_18371);
or UO_795 (O_795,N_18295,N_18186);
nand UO_796 (O_796,N_18969,N_18055);
and UO_797 (O_797,N_18349,N_18403);
nand UO_798 (O_798,N_18689,N_18204);
nand UO_799 (O_799,N_19978,N_19582);
or UO_800 (O_800,N_19785,N_19161);
nand UO_801 (O_801,N_19443,N_19734);
nor UO_802 (O_802,N_18000,N_18051);
nor UO_803 (O_803,N_18308,N_19775);
or UO_804 (O_804,N_19647,N_19533);
xnor UO_805 (O_805,N_19525,N_19233);
nand UO_806 (O_806,N_19973,N_19867);
nor UO_807 (O_807,N_19926,N_19006);
nand UO_808 (O_808,N_19813,N_18706);
or UO_809 (O_809,N_18695,N_18587);
nand UO_810 (O_810,N_19956,N_19011);
and UO_811 (O_811,N_19359,N_18115);
and UO_812 (O_812,N_19781,N_18338);
nand UO_813 (O_813,N_19696,N_19639);
nor UO_814 (O_814,N_18252,N_18666);
or UO_815 (O_815,N_19931,N_18692);
nor UO_816 (O_816,N_19557,N_19854);
or UO_817 (O_817,N_18826,N_18225);
or UO_818 (O_818,N_18240,N_19606);
nor UO_819 (O_819,N_18244,N_18619);
nand UO_820 (O_820,N_18991,N_19574);
or UO_821 (O_821,N_19303,N_19972);
xnor UO_822 (O_822,N_19100,N_19220);
nor UO_823 (O_823,N_19219,N_18446);
or UO_824 (O_824,N_19323,N_18100);
nor UO_825 (O_825,N_19818,N_19105);
nor UO_826 (O_826,N_19909,N_18207);
or UO_827 (O_827,N_18291,N_19605);
xnor UO_828 (O_828,N_19728,N_19902);
or UO_829 (O_829,N_19826,N_19083);
nand UO_830 (O_830,N_19008,N_18975);
or UO_831 (O_831,N_19623,N_18324);
or UO_832 (O_832,N_19459,N_19242);
or UO_833 (O_833,N_18832,N_19743);
and UO_834 (O_834,N_19876,N_19673);
and UO_835 (O_835,N_19215,N_19600);
nor UO_836 (O_836,N_19468,N_19088);
and UO_837 (O_837,N_18761,N_18383);
and UO_838 (O_838,N_19955,N_18964);
or UO_839 (O_839,N_19621,N_19566);
and UO_840 (O_840,N_18854,N_19126);
nand UO_841 (O_841,N_19292,N_19742);
xnor UO_842 (O_842,N_19986,N_18746);
nor UO_843 (O_843,N_19431,N_18995);
and UO_844 (O_844,N_19072,N_19654);
nand UO_845 (O_845,N_18726,N_18350);
nand UO_846 (O_846,N_19182,N_18410);
and UO_847 (O_847,N_19686,N_18838);
and UO_848 (O_848,N_18719,N_19077);
nor UO_849 (O_849,N_19827,N_18381);
nor UO_850 (O_850,N_19567,N_19793);
nor UO_851 (O_851,N_19706,N_19591);
xnor UO_852 (O_852,N_19771,N_18044);
and UO_853 (O_853,N_18242,N_19924);
or UO_854 (O_854,N_18236,N_19967);
nand UO_855 (O_855,N_18453,N_18660);
or UO_856 (O_856,N_19422,N_19178);
nor UO_857 (O_857,N_19831,N_18406);
nor UO_858 (O_858,N_18754,N_18915);
nor UO_859 (O_859,N_19096,N_19716);
or UO_860 (O_860,N_19927,N_18771);
and UO_861 (O_861,N_18303,N_19136);
or UO_862 (O_862,N_18149,N_18525);
and UO_863 (O_863,N_18948,N_19512);
or UO_864 (O_864,N_19266,N_18233);
and UO_865 (O_865,N_19462,N_19383);
nor UO_866 (O_866,N_19816,N_18175);
xnor UO_867 (O_867,N_19196,N_19962);
nor UO_868 (O_868,N_19276,N_18301);
and UO_869 (O_869,N_19214,N_18074);
and UO_870 (O_870,N_19349,N_19811);
and UO_871 (O_871,N_18567,N_19270);
or UO_872 (O_872,N_18555,N_18687);
or UO_873 (O_873,N_18094,N_19111);
nor UO_874 (O_874,N_18678,N_18469);
nor UO_875 (O_875,N_18039,N_19351);
nand UO_876 (O_876,N_19916,N_19975);
nor UO_877 (O_877,N_19244,N_19331);
or UO_878 (O_878,N_19691,N_19007);
nand UO_879 (O_879,N_19906,N_18411);
and UO_880 (O_880,N_18848,N_19116);
nor UO_881 (O_881,N_18147,N_19391);
nand UO_882 (O_882,N_19776,N_18213);
nand UO_883 (O_883,N_18459,N_18367);
or UO_884 (O_884,N_18711,N_19120);
nor UO_885 (O_885,N_19494,N_19945);
nor UO_886 (O_886,N_19857,N_19277);
or UO_887 (O_887,N_18313,N_19155);
nor UO_888 (O_888,N_19795,N_18412);
nand UO_889 (O_889,N_19671,N_18656);
nor UO_890 (O_890,N_19510,N_19035);
or UO_891 (O_891,N_18559,N_19903);
and UO_892 (O_892,N_18820,N_18870);
nor UO_893 (O_893,N_18390,N_19534);
or UO_894 (O_894,N_19668,N_19133);
or UO_895 (O_895,N_19263,N_18720);
or UO_896 (O_896,N_19221,N_18607);
nand UO_897 (O_897,N_18822,N_18037);
and UO_898 (O_898,N_19070,N_19593);
xnor UO_899 (O_899,N_19516,N_18064);
or UO_900 (O_900,N_18506,N_19411);
nor UO_901 (O_901,N_18647,N_19746);
xnor UO_902 (O_902,N_19500,N_19344);
nand UO_903 (O_903,N_19957,N_19354);
xor UO_904 (O_904,N_19031,N_18195);
xnor UO_905 (O_905,N_19779,N_19900);
nor UO_906 (O_906,N_18065,N_19307);
nor UO_907 (O_907,N_18891,N_19324);
and UO_908 (O_908,N_18070,N_18104);
nand UO_909 (O_909,N_19784,N_19448);
and UO_910 (O_910,N_18214,N_18616);
nor UO_911 (O_911,N_19157,N_18172);
or UO_912 (O_912,N_18859,N_18391);
nor UO_913 (O_913,N_19873,N_18586);
nor UO_914 (O_914,N_18745,N_18491);
and UO_915 (O_915,N_19358,N_19444);
or UO_916 (O_916,N_18690,N_18814);
or UO_917 (O_917,N_19051,N_19770);
and UO_918 (O_918,N_18641,N_18649);
nand UO_919 (O_919,N_19727,N_18137);
nand UO_920 (O_920,N_19286,N_19946);
or UO_921 (O_921,N_18287,N_18923);
xnor UO_922 (O_922,N_19923,N_18615);
nor UO_923 (O_923,N_19417,N_18919);
nand UO_924 (O_924,N_18370,N_19201);
or UO_925 (O_925,N_18734,N_18404);
and UO_926 (O_926,N_18310,N_19497);
and UO_927 (O_927,N_18899,N_19562);
nand UO_928 (O_928,N_18638,N_18445);
xnor UO_929 (O_929,N_18768,N_18835);
nand UO_930 (O_930,N_19514,N_18741);
xnor UO_931 (O_931,N_18674,N_19003);
or UO_932 (O_932,N_18882,N_19394);
xnor UO_933 (O_933,N_19913,N_18111);
and UO_934 (O_934,N_18667,N_19298);
nand UO_935 (O_935,N_18465,N_19176);
and UO_936 (O_936,N_18296,N_18729);
nand UO_937 (O_937,N_18028,N_18114);
nand UO_938 (O_938,N_18050,N_19815);
nor UO_939 (O_939,N_18358,N_18917);
or UO_940 (O_940,N_18515,N_19139);
nor UO_941 (O_941,N_18080,N_19607);
and UO_942 (O_942,N_18994,N_19992);
nor UO_943 (O_943,N_19289,N_19137);
and UO_944 (O_944,N_18849,N_18672);
nand UO_945 (O_945,N_19053,N_19856);
nand UO_946 (O_946,N_18812,N_19618);
nand UO_947 (O_947,N_19570,N_19098);
and UO_948 (O_948,N_18533,N_18347);
or UO_949 (O_949,N_19659,N_19336);
nand UO_950 (O_950,N_19130,N_18654);
nand UO_951 (O_951,N_19782,N_19152);
and UO_952 (O_952,N_18136,N_18566);
xnor UO_953 (O_953,N_18123,N_19427);
nand UO_954 (O_954,N_19724,N_19049);
and UO_955 (O_955,N_18083,N_18387);
and UO_956 (O_956,N_19205,N_18979);
and UO_957 (O_957,N_19589,N_18830);
nor UO_958 (O_958,N_18075,N_18444);
and UO_959 (O_959,N_19561,N_18222);
and UO_960 (O_960,N_18897,N_19061);
nor UO_961 (O_961,N_18426,N_19029);
or UO_962 (O_962,N_19918,N_18209);
nand UO_963 (O_963,N_18378,N_18831);
xor UO_964 (O_964,N_19995,N_19506);
or UO_965 (O_965,N_19958,N_18628);
nor UO_966 (O_966,N_19416,N_19295);
or UO_967 (O_967,N_18758,N_19578);
or UO_968 (O_968,N_19015,N_18223);
and UO_969 (O_969,N_18983,N_19162);
or UO_970 (O_970,N_19904,N_18278);
nand UO_971 (O_971,N_19078,N_19466);
xnor UO_972 (O_972,N_19661,N_19142);
nor UO_973 (O_973,N_19523,N_19964);
xnor UO_974 (O_974,N_18190,N_18742);
nand UO_975 (O_975,N_18610,N_19329);
nand UO_976 (O_976,N_18646,N_19445);
and UO_977 (O_977,N_18150,N_19543);
nand UO_978 (O_978,N_18828,N_19224);
or UO_979 (O_979,N_19491,N_18231);
nor UO_980 (O_980,N_18932,N_19544);
nand UO_981 (O_981,N_18215,N_18593);
and UO_982 (O_982,N_18556,N_19808);
nor UO_983 (O_983,N_18012,N_18476);
nand UO_984 (O_984,N_18670,N_18098);
nand UO_985 (O_985,N_18056,N_18569);
xor UO_986 (O_986,N_19930,N_18833);
nand UO_987 (O_987,N_19320,N_18475);
nor UO_988 (O_988,N_18271,N_19855);
nor UO_989 (O_989,N_19653,N_18156);
xnor UO_990 (O_990,N_19073,N_19308);
nand UO_991 (O_991,N_19948,N_18017);
nor UO_992 (O_992,N_19850,N_19353);
nor UO_993 (O_993,N_18594,N_18611);
nand UO_994 (O_994,N_18143,N_18202);
xnor UO_995 (O_995,N_19786,N_18965);
nand UO_996 (O_996,N_18451,N_18488);
or UO_997 (O_997,N_18373,N_18522);
nand UO_998 (O_998,N_19869,N_19890);
nand UO_999 (O_999,N_18466,N_19936);
and UO_1000 (O_1000,N_18223,N_18439);
xor UO_1001 (O_1001,N_19834,N_18012);
nor UO_1002 (O_1002,N_18742,N_18782);
or UO_1003 (O_1003,N_19821,N_18964);
xnor UO_1004 (O_1004,N_18827,N_19296);
xor UO_1005 (O_1005,N_18658,N_19012);
or UO_1006 (O_1006,N_18818,N_19221);
and UO_1007 (O_1007,N_18279,N_19646);
xor UO_1008 (O_1008,N_18866,N_18312);
and UO_1009 (O_1009,N_19419,N_18056);
or UO_1010 (O_1010,N_18054,N_18714);
nor UO_1011 (O_1011,N_19590,N_18224);
or UO_1012 (O_1012,N_18938,N_18019);
and UO_1013 (O_1013,N_19018,N_19747);
and UO_1014 (O_1014,N_18273,N_19762);
xnor UO_1015 (O_1015,N_18628,N_18637);
nor UO_1016 (O_1016,N_18566,N_19930);
nor UO_1017 (O_1017,N_18087,N_19099);
nor UO_1018 (O_1018,N_18167,N_19603);
nand UO_1019 (O_1019,N_19518,N_19490);
nand UO_1020 (O_1020,N_18403,N_19829);
and UO_1021 (O_1021,N_19731,N_18090);
nand UO_1022 (O_1022,N_19477,N_19244);
nand UO_1023 (O_1023,N_19004,N_18858);
or UO_1024 (O_1024,N_19786,N_18325);
nor UO_1025 (O_1025,N_19077,N_18451);
and UO_1026 (O_1026,N_18199,N_19155);
xor UO_1027 (O_1027,N_18539,N_18172);
nor UO_1028 (O_1028,N_19189,N_19756);
nor UO_1029 (O_1029,N_18778,N_18155);
xor UO_1030 (O_1030,N_18546,N_18320);
or UO_1031 (O_1031,N_18771,N_18401);
nand UO_1032 (O_1032,N_19567,N_18854);
and UO_1033 (O_1033,N_18481,N_19419);
xor UO_1034 (O_1034,N_18752,N_19929);
or UO_1035 (O_1035,N_18278,N_19656);
nand UO_1036 (O_1036,N_19238,N_19122);
nand UO_1037 (O_1037,N_18761,N_18987);
and UO_1038 (O_1038,N_19847,N_18687);
and UO_1039 (O_1039,N_18064,N_19846);
or UO_1040 (O_1040,N_18606,N_18219);
or UO_1041 (O_1041,N_19496,N_19674);
nand UO_1042 (O_1042,N_19400,N_18933);
nand UO_1043 (O_1043,N_18276,N_18300);
or UO_1044 (O_1044,N_19237,N_18628);
nor UO_1045 (O_1045,N_18334,N_19444);
or UO_1046 (O_1046,N_19212,N_19135);
and UO_1047 (O_1047,N_19529,N_19625);
nor UO_1048 (O_1048,N_18334,N_18941);
and UO_1049 (O_1049,N_18123,N_19818);
or UO_1050 (O_1050,N_18807,N_18089);
xnor UO_1051 (O_1051,N_18235,N_19219);
or UO_1052 (O_1052,N_18860,N_18609);
nand UO_1053 (O_1053,N_19262,N_18763);
nor UO_1054 (O_1054,N_18459,N_19109);
and UO_1055 (O_1055,N_18001,N_19301);
or UO_1056 (O_1056,N_19691,N_18162);
or UO_1057 (O_1057,N_18132,N_19757);
nand UO_1058 (O_1058,N_18864,N_18001);
and UO_1059 (O_1059,N_18013,N_19338);
or UO_1060 (O_1060,N_19002,N_19508);
or UO_1061 (O_1061,N_18712,N_19013);
nand UO_1062 (O_1062,N_18235,N_18408);
or UO_1063 (O_1063,N_18411,N_19714);
nor UO_1064 (O_1064,N_18114,N_18112);
or UO_1065 (O_1065,N_19940,N_18055);
and UO_1066 (O_1066,N_19248,N_18231);
and UO_1067 (O_1067,N_18166,N_19973);
nor UO_1068 (O_1068,N_18870,N_18930);
and UO_1069 (O_1069,N_19297,N_19960);
or UO_1070 (O_1070,N_19524,N_18818);
and UO_1071 (O_1071,N_19644,N_18297);
or UO_1072 (O_1072,N_18477,N_18626);
xnor UO_1073 (O_1073,N_19544,N_19168);
nor UO_1074 (O_1074,N_18525,N_19363);
nor UO_1075 (O_1075,N_19512,N_19391);
xor UO_1076 (O_1076,N_18232,N_18964);
or UO_1077 (O_1077,N_18242,N_18944);
or UO_1078 (O_1078,N_18858,N_19242);
or UO_1079 (O_1079,N_19496,N_19554);
nand UO_1080 (O_1080,N_18735,N_18516);
and UO_1081 (O_1081,N_18474,N_18325);
or UO_1082 (O_1082,N_19712,N_19736);
or UO_1083 (O_1083,N_18598,N_19256);
nor UO_1084 (O_1084,N_19729,N_18512);
nor UO_1085 (O_1085,N_18855,N_19170);
nand UO_1086 (O_1086,N_18847,N_18966);
or UO_1087 (O_1087,N_18438,N_19009);
or UO_1088 (O_1088,N_19360,N_18125);
and UO_1089 (O_1089,N_18457,N_19739);
nand UO_1090 (O_1090,N_18672,N_19325);
or UO_1091 (O_1091,N_18852,N_18130);
nor UO_1092 (O_1092,N_19519,N_19155);
xnor UO_1093 (O_1093,N_19574,N_18063);
nand UO_1094 (O_1094,N_19526,N_19825);
nand UO_1095 (O_1095,N_19900,N_18285);
nor UO_1096 (O_1096,N_19493,N_19560);
nand UO_1097 (O_1097,N_18307,N_19396);
nor UO_1098 (O_1098,N_18814,N_18936);
xor UO_1099 (O_1099,N_18758,N_18713);
nand UO_1100 (O_1100,N_19919,N_18156);
nor UO_1101 (O_1101,N_18065,N_18977);
nor UO_1102 (O_1102,N_18326,N_19020);
xnor UO_1103 (O_1103,N_19099,N_19282);
and UO_1104 (O_1104,N_18442,N_19730);
or UO_1105 (O_1105,N_19784,N_19444);
and UO_1106 (O_1106,N_19342,N_18578);
and UO_1107 (O_1107,N_18921,N_18003);
or UO_1108 (O_1108,N_19204,N_19757);
and UO_1109 (O_1109,N_19680,N_18587);
nor UO_1110 (O_1110,N_18467,N_18495);
nand UO_1111 (O_1111,N_19231,N_18853);
or UO_1112 (O_1112,N_19354,N_19280);
nand UO_1113 (O_1113,N_19624,N_18543);
nand UO_1114 (O_1114,N_19363,N_18314);
and UO_1115 (O_1115,N_19155,N_19467);
and UO_1116 (O_1116,N_19713,N_18509);
or UO_1117 (O_1117,N_19086,N_19958);
nand UO_1118 (O_1118,N_19536,N_18613);
nand UO_1119 (O_1119,N_18340,N_19346);
or UO_1120 (O_1120,N_19173,N_19387);
or UO_1121 (O_1121,N_18461,N_19823);
nor UO_1122 (O_1122,N_18403,N_18952);
and UO_1123 (O_1123,N_19373,N_19792);
and UO_1124 (O_1124,N_19639,N_18202);
and UO_1125 (O_1125,N_18974,N_18881);
nor UO_1126 (O_1126,N_19205,N_19245);
and UO_1127 (O_1127,N_18999,N_19066);
nand UO_1128 (O_1128,N_19760,N_18151);
nand UO_1129 (O_1129,N_18396,N_18562);
nor UO_1130 (O_1130,N_19730,N_19205);
and UO_1131 (O_1131,N_18648,N_18249);
nor UO_1132 (O_1132,N_19918,N_18717);
nor UO_1133 (O_1133,N_19593,N_19685);
and UO_1134 (O_1134,N_18069,N_18081);
nor UO_1135 (O_1135,N_19664,N_18867);
or UO_1136 (O_1136,N_18205,N_19975);
and UO_1137 (O_1137,N_19611,N_18718);
or UO_1138 (O_1138,N_18616,N_19219);
nor UO_1139 (O_1139,N_19321,N_19020);
xor UO_1140 (O_1140,N_19457,N_18485);
nand UO_1141 (O_1141,N_19784,N_19533);
and UO_1142 (O_1142,N_18813,N_19790);
and UO_1143 (O_1143,N_18976,N_18874);
and UO_1144 (O_1144,N_18819,N_18001);
and UO_1145 (O_1145,N_18514,N_19446);
nor UO_1146 (O_1146,N_18444,N_18551);
nor UO_1147 (O_1147,N_19584,N_18382);
nand UO_1148 (O_1148,N_19235,N_18432);
and UO_1149 (O_1149,N_19637,N_18161);
nand UO_1150 (O_1150,N_19889,N_19269);
nor UO_1151 (O_1151,N_18646,N_19672);
and UO_1152 (O_1152,N_19373,N_18635);
or UO_1153 (O_1153,N_18276,N_18466);
nor UO_1154 (O_1154,N_19750,N_18496);
nor UO_1155 (O_1155,N_18385,N_18161);
nand UO_1156 (O_1156,N_19582,N_18240);
and UO_1157 (O_1157,N_19226,N_18889);
nor UO_1158 (O_1158,N_18355,N_19786);
or UO_1159 (O_1159,N_18074,N_19207);
nand UO_1160 (O_1160,N_18357,N_19176);
nand UO_1161 (O_1161,N_18477,N_19227);
or UO_1162 (O_1162,N_19367,N_19686);
and UO_1163 (O_1163,N_19306,N_19799);
and UO_1164 (O_1164,N_19755,N_19238);
or UO_1165 (O_1165,N_19290,N_18744);
and UO_1166 (O_1166,N_19189,N_18014);
and UO_1167 (O_1167,N_19024,N_19705);
and UO_1168 (O_1168,N_18556,N_18569);
and UO_1169 (O_1169,N_19409,N_19571);
nand UO_1170 (O_1170,N_18266,N_19931);
or UO_1171 (O_1171,N_19296,N_18776);
or UO_1172 (O_1172,N_19859,N_19413);
and UO_1173 (O_1173,N_18509,N_19224);
nor UO_1174 (O_1174,N_19176,N_18287);
xor UO_1175 (O_1175,N_18801,N_19514);
or UO_1176 (O_1176,N_19461,N_18599);
and UO_1177 (O_1177,N_18958,N_18956);
xnor UO_1178 (O_1178,N_19168,N_19068);
nand UO_1179 (O_1179,N_19941,N_18228);
nor UO_1180 (O_1180,N_19923,N_19409);
nand UO_1181 (O_1181,N_18718,N_18679);
nand UO_1182 (O_1182,N_18538,N_18134);
nor UO_1183 (O_1183,N_18067,N_19930);
and UO_1184 (O_1184,N_19018,N_19282);
nor UO_1185 (O_1185,N_19608,N_18009);
or UO_1186 (O_1186,N_19839,N_19233);
xnor UO_1187 (O_1187,N_18325,N_18286);
and UO_1188 (O_1188,N_19329,N_19388);
nand UO_1189 (O_1189,N_19034,N_19028);
nand UO_1190 (O_1190,N_18344,N_18416);
or UO_1191 (O_1191,N_19375,N_18672);
and UO_1192 (O_1192,N_19895,N_19433);
nor UO_1193 (O_1193,N_19036,N_18111);
nand UO_1194 (O_1194,N_19932,N_19552);
nand UO_1195 (O_1195,N_18359,N_19435);
nand UO_1196 (O_1196,N_18143,N_19187);
or UO_1197 (O_1197,N_18904,N_19841);
or UO_1198 (O_1198,N_19446,N_19117);
xor UO_1199 (O_1199,N_18096,N_18749);
nand UO_1200 (O_1200,N_19470,N_18873);
and UO_1201 (O_1201,N_19798,N_19629);
or UO_1202 (O_1202,N_18468,N_18136);
nor UO_1203 (O_1203,N_19072,N_18226);
nand UO_1204 (O_1204,N_19684,N_18209);
and UO_1205 (O_1205,N_19994,N_19034);
nand UO_1206 (O_1206,N_18070,N_18866);
and UO_1207 (O_1207,N_19859,N_18565);
and UO_1208 (O_1208,N_18754,N_18766);
or UO_1209 (O_1209,N_18261,N_19021);
nor UO_1210 (O_1210,N_18745,N_19874);
xor UO_1211 (O_1211,N_18408,N_18386);
nor UO_1212 (O_1212,N_18862,N_18659);
xnor UO_1213 (O_1213,N_18706,N_18334);
xor UO_1214 (O_1214,N_19910,N_19407);
xnor UO_1215 (O_1215,N_18472,N_18803);
nor UO_1216 (O_1216,N_19480,N_18050);
or UO_1217 (O_1217,N_18268,N_19933);
nor UO_1218 (O_1218,N_19041,N_18627);
xor UO_1219 (O_1219,N_18753,N_18997);
nor UO_1220 (O_1220,N_18632,N_18363);
or UO_1221 (O_1221,N_18762,N_19416);
nor UO_1222 (O_1222,N_18585,N_18488);
nor UO_1223 (O_1223,N_18438,N_18657);
or UO_1224 (O_1224,N_18474,N_18852);
nor UO_1225 (O_1225,N_18384,N_18561);
or UO_1226 (O_1226,N_19575,N_19113);
nand UO_1227 (O_1227,N_18252,N_18040);
or UO_1228 (O_1228,N_19817,N_18920);
or UO_1229 (O_1229,N_18903,N_18152);
nand UO_1230 (O_1230,N_19565,N_19772);
and UO_1231 (O_1231,N_19438,N_19859);
or UO_1232 (O_1232,N_19114,N_19940);
and UO_1233 (O_1233,N_18134,N_18144);
xnor UO_1234 (O_1234,N_18519,N_18671);
or UO_1235 (O_1235,N_19729,N_19770);
and UO_1236 (O_1236,N_18975,N_19465);
nand UO_1237 (O_1237,N_19762,N_18432);
nand UO_1238 (O_1238,N_19283,N_18401);
and UO_1239 (O_1239,N_19176,N_19316);
and UO_1240 (O_1240,N_19715,N_19740);
nor UO_1241 (O_1241,N_19859,N_18190);
or UO_1242 (O_1242,N_19924,N_18314);
or UO_1243 (O_1243,N_18887,N_18274);
xnor UO_1244 (O_1244,N_18406,N_18838);
nor UO_1245 (O_1245,N_18658,N_18576);
nand UO_1246 (O_1246,N_18052,N_18638);
nor UO_1247 (O_1247,N_18775,N_19801);
nor UO_1248 (O_1248,N_19789,N_18408);
nand UO_1249 (O_1249,N_18936,N_19278);
nor UO_1250 (O_1250,N_18680,N_18912);
nand UO_1251 (O_1251,N_19948,N_18877);
nor UO_1252 (O_1252,N_18010,N_18495);
xor UO_1253 (O_1253,N_18923,N_19784);
nand UO_1254 (O_1254,N_19785,N_19813);
and UO_1255 (O_1255,N_19834,N_19766);
or UO_1256 (O_1256,N_18828,N_18642);
or UO_1257 (O_1257,N_19481,N_18835);
nor UO_1258 (O_1258,N_18701,N_18558);
nor UO_1259 (O_1259,N_18636,N_19552);
or UO_1260 (O_1260,N_19277,N_18551);
or UO_1261 (O_1261,N_19806,N_18260);
nor UO_1262 (O_1262,N_18015,N_19151);
and UO_1263 (O_1263,N_18646,N_18554);
nand UO_1264 (O_1264,N_19665,N_18849);
or UO_1265 (O_1265,N_19288,N_19424);
and UO_1266 (O_1266,N_19054,N_18863);
or UO_1267 (O_1267,N_18534,N_19557);
nand UO_1268 (O_1268,N_18686,N_19647);
or UO_1269 (O_1269,N_19284,N_19944);
nand UO_1270 (O_1270,N_19095,N_18181);
or UO_1271 (O_1271,N_19094,N_19485);
and UO_1272 (O_1272,N_19869,N_19221);
nand UO_1273 (O_1273,N_18027,N_18884);
and UO_1274 (O_1274,N_19224,N_19276);
nand UO_1275 (O_1275,N_18360,N_18995);
or UO_1276 (O_1276,N_18122,N_19194);
nor UO_1277 (O_1277,N_19951,N_19216);
and UO_1278 (O_1278,N_19373,N_18036);
or UO_1279 (O_1279,N_18157,N_18966);
and UO_1280 (O_1280,N_19584,N_18092);
nor UO_1281 (O_1281,N_19291,N_18362);
nor UO_1282 (O_1282,N_19448,N_19397);
and UO_1283 (O_1283,N_19373,N_18648);
nor UO_1284 (O_1284,N_19542,N_19309);
nand UO_1285 (O_1285,N_18486,N_19566);
or UO_1286 (O_1286,N_19925,N_18890);
xor UO_1287 (O_1287,N_18256,N_19924);
nor UO_1288 (O_1288,N_19804,N_18875);
nor UO_1289 (O_1289,N_19439,N_18024);
nand UO_1290 (O_1290,N_18461,N_19668);
nand UO_1291 (O_1291,N_19801,N_18488);
nand UO_1292 (O_1292,N_19002,N_18496);
or UO_1293 (O_1293,N_19694,N_18351);
or UO_1294 (O_1294,N_18458,N_18697);
xnor UO_1295 (O_1295,N_19740,N_19352);
or UO_1296 (O_1296,N_18205,N_18136);
nor UO_1297 (O_1297,N_18368,N_19958);
and UO_1298 (O_1298,N_19837,N_19865);
or UO_1299 (O_1299,N_18472,N_19830);
or UO_1300 (O_1300,N_19913,N_19459);
xor UO_1301 (O_1301,N_18154,N_18312);
and UO_1302 (O_1302,N_18841,N_18533);
and UO_1303 (O_1303,N_19123,N_19936);
or UO_1304 (O_1304,N_18861,N_19008);
nor UO_1305 (O_1305,N_19617,N_18481);
nand UO_1306 (O_1306,N_18004,N_19280);
nand UO_1307 (O_1307,N_18246,N_19833);
nand UO_1308 (O_1308,N_18951,N_18972);
or UO_1309 (O_1309,N_19569,N_18280);
or UO_1310 (O_1310,N_18593,N_19767);
xnor UO_1311 (O_1311,N_19274,N_19473);
nand UO_1312 (O_1312,N_19548,N_18515);
nor UO_1313 (O_1313,N_18137,N_19243);
and UO_1314 (O_1314,N_18964,N_19535);
and UO_1315 (O_1315,N_18704,N_18542);
xnor UO_1316 (O_1316,N_19772,N_18906);
xor UO_1317 (O_1317,N_18325,N_19356);
nand UO_1318 (O_1318,N_18882,N_19252);
and UO_1319 (O_1319,N_18050,N_18057);
nand UO_1320 (O_1320,N_18453,N_19670);
or UO_1321 (O_1321,N_18670,N_19170);
or UO_1322 (O_1322,N_19974,N_18255);
or UO_1323 (O_1323,N_18037,N_18133);
nand UO_1324 (O_1324,N_18514,N_19789);
or UO_1325 (O_1325,N_18016,N_18363);
and UO_1326 (O_1326,N_18196,N_18321);
nor UO_1327 (O_1327,N_18627,N_18074);
or UO_1328 (O_1328,N_19357,N_18505);
nand UO_1329 (O_1329,N_19538,N_18634);
or UO_1330 (O_1330,N_18416,N_19591);
and UO_1331 (O_1331,N_19815,N_19457);
and UO_1332 (O_1332,N_19814,N_19241);
xor UO_1333 (O_1333,N_19870,N_19001);
and UO_1334 (O_1334,N_18480,N_19386);
nand UO_1335 (O_1335,N_18772,N_18812);
or UO_1336 (O_1336,N_19207,N_18267);
nand UO_1337 (O_1337,N_19142,N_18507);
or UO_1338 (O_1338,N_18785,N_18999);
nor UO_1339 (O_1339,N_18479,N_19580);
xor UO_1340 (O_1340,N_19596,N_19870);
nor UO_1341 (O_1341,N_18974,N_18554);
and UO_1342 (O_1342,N_19851,N_19448);
xnor UO_1343 (O_1343,N_18636,N_18494);
xnor UO_1344 (O_1344,N_18748,N_19771);
nor UO_1345 (O_1345,N_18786,N_18261);
xor UO_1346 (O_1346,N_19949,N_18613);
nand UO_1347 (O_1347,N_19175,N_18317);
and UO_1348 (O_1348,N_18591,N_19727);
nor UO_1349 (O_1349,N_18303,N_18749);
nor UO_1350 (O_1350,N_18076,N_18489);
and UO_1351 (O_1351,N_19047,N_19139);
nor UO_1352 (O_1352,N_18982,N_19149);
nor UO_1353 (O_1353,N_18866,N_18104);
nand UO_1354 (O_1354,N_18205,N_19825);
or UO_1355 (O_1355,N_18305,N_18325);
nor UO_1356 (O_1356,N_18134,N_19781);
xnor UO_1357 (O_1357,N_19478,N_18514);
or UO_1358 (O_1358,N_19696,N_19559);
xor UO_1359 (O_1359,N_19844,N_19395);
or UO_1360 (O_1360,N_19583,N_19677);
nand UO_1361 (O_1361,N_19229,N_19195);
or UO_1362 (O_1362,N_19031,N_18863);
or UO_1363 (O_1363,N_19818,N_19729);
nand UO_1364 (O_1364,N_18668,N_18660);
nor UO_1365 (O_1365,N_19112,N_19462);
nand UO_1366 (O_1366,N_18941,N_19783);
nor UO_1367 (O_1367,N_18614,N_18997);
nor UO_1368 (O_1368,N_18650,N_19440);
or UO_1369 (O_1369,N_18839,N_19085);
xnor UO_1370 (O_1370,N_18147,N_18752);
nand UO_1371 (O_1371,N_18305,N_19211);
and UO_1372 (O_1372,N_19067,N_19376);
and UO_1373 (O_1373,N_18307,N_18679);
nor UO_1374 (O_1374,N_19326,N_19030);
or UO_1375 (O_1375,N_18879,N_19201);
and UO_1376 (O_1376,N_18549,N_19196);
or UO_1377 (O_1377,N_19747,N_18637);
nand UO_1378 (O_1378,N_19005,N_18857);
nand UO_1379 (O_1379,N_18015,N_19820);
or UO_1380 (O_1380,N_19772,N_19649);
xor UO_1381 (O_1381,N_18326,N_19810);
xnor UO_1382 (O_1382,N_18454,N_18236);
or UO_1383 (O_1383,N_19818,N_18159);
and UO_1384 (O_1384,N_19628,N_18180);
or UO_1385 (O_1385,N_18740,N_18577);
nor UO_1386 (O_1386,N_19328,N_18388);
and UO_1387 (O_1387,N_18929,N_19284);
and UO_1388 (O_1388,N_19249,N_19471);
and UO_1389 (O_1389,N_18349,N_19020);
nor UO_1390 (O_1390,N_19539,N_19659);
nand UO_1391 (O_1391,N_18496,N_18322);
and UO_1392 (O_1392,N_18822,N_19720);
nor UO_1393 (O_1393,N_18419,N_19542);
xnor UO_1394 (O_1394,N_18122,N_19196);
or UO_1395 (O_1395,N_19913,N_18761);
or UO_1396 (O_1396,N_19848,N_19806);
or UO_1397 (O_1397,N_18531,N_19907);
xor UO_1398 (O_1398,N_19765,N_18452);
nor UO_1399 (O_1399,N_18557,N_18121);
or UO_1400 (O_1400,N_18841,N_18600);
and UO_1401 (O_1401,N_18110,N_18517);
nor UO_1402 (O_1402,N_19261,N_19146);
and UO_1403 (O_1403,N_19202,N_18004);
nor UO_1404 (O_1404,N_19468,N_19234);
xor UO_1405 (O_1405,N_19372,N_19933);
nand UO_1406 (O_1406,N_19718,N_18383);
nand UO_1407 (O_1407,N_18798,N_18753);
and UO_1408 (O_1408,N_18596,N_18833);
xnor UO_1409 (O_1409,N_18995,N_18159);
or UO_1410 (O_1410,N_18993,N_19731);
nand UO_1411 (O_1411,N_18715,N_19807);
nand UO_1412 (O_1412,N_19410,N_19498);
or UO_1413 (O_1413,N_19607,N_19093);
xnor UO_1414 (O_1414,N_18659,N_18992);
and UO_1415 (O_1415,N_18284,N_18041);
and UO_1416 (O_1416,N_19513,N_18023);
and UO_1417 (O_1417,N_18772,N_19822);
nor UO_1418 (O_1418,N_19915,N_19580);
xor UO_1419 (O_1419,N_19803,N_18339);
and UO_1420 (O_1420,N_19046,N_18252);
nor UO_1421 (O_1421,N_18475,N_19793);
nand UO_1422 (O_1422,N_19903,N_19279);
or UO_1423 (O_1423,N_18307,N_18619);
and UO_1424 (O_1424,N_19583,N_19746);
and UO_1425 (O_1425,N_18978,N_19687);
and UO_1426 (O_1426,N_18970,N_18179);
or UO_1427 (O_1427,N_19019,N_19865);
nor UO_1428 (O_1428,N_19903,N_18451);
or UO_1429 (O_1429,N_18660,N_19848);
and UO_1430 (O_1430,N_19978,N_18026);
nor UO_1431 (O_1431,N_18593,N_18272);
nor UO_1432 (O_1432,N_19735,N_19461);
or UO_1433 (O_1433,N_18870,N_18931);
and UO_1434 (O_1434,N_19488,N_18527);
xor UO_1435 (O_1435,N_18258,N_18350);
or UO_1436 (O_1436,N_19145,N_18225);
or UO_1437 (O_1437,N_18315,N_18743);
nor UO_1438 (O_1438,N_18721,N_19043);
nor UO_1439 (O_1439,N_18435,N_19400);
and UO_1440 (O_1440,N_18035,N_19882);
or UO_1441 (O_1441,N_19131,N_19402);
or UO_1442 (O_1442,N_19703,N_19084);
or UO_1443 (O_1443,N_19062,N_18074);
or UO_1444 (O_1444,N_18938,N_19089);
xnor UO_1445 (O_1445,N_19560,N_19867);
xnor UO_1446 (O_1446,N_18131,N_19271);
nor UO_1447 (O_1447,N_18916,N_18206);
or UO_1448 (O_1448,N_18221,N_19008);
or UO_1449 (O_1449,N_19711,N_18686);
and UO_1450 (O_1450,N_19081,N_18841);
nor UO_1451 (O_1451,N_18175,N_18268);
nand UO_1452 (O_1452,N_19982,N_19374);
and UO_1453 (O_1453,N_18320,N_18282);
or UO_1454 (O_1454,N_18833,N_18856);
and UO_1455 (O_1455,N_19313,N_18952);
or UO_1456 (O_1456,N_19632,N_18707);
nor UO_1457 (O_1457,N_19872,N_18392);
nor UO_1458 (O_1458,N_19231,N_19789);
xnor UO_1459 (O_1459,N_18333,N_18868);
nand UO_1460 (O_1460,N_18785,N_19015);
nor UO_1461 (O_1461,N_19715,N_18715);
xor UO_1462 (O_1462,N_18076,N_18318);
nor UO_1463 (O_1463,N_19837,N_18791);
and UO_1464 (O_1464,N_18478,N_18581);
and UO_1465 (O_1465,N_18304,N_18274);
nand UO_1466 (O_1466,N_19236,N_18974);
nor UO_1467 (O_1467,N_19925,N_19857);
xnor UO_1468 (O_1468,N_18994,N_19763);
nor UO_1469 (O_1469,N_19462,N_19610);
xor UO_1470 (O_1470,N_19053,N_18696);
and UO_1471 (O_1471,N_18696,N_19820);
and UO_1472 (O_1472,N_19388,N_19806);
or UO_1473 (O_1473,N_18733,N_18548);
or UO_1474 (O_1474,N_18502,N_19981);
nor UO_1475 (O_1475,N_19925,N_19998);
or UO_1476 (O_1476,N_18232,N_19228);
or UO_1477 (O_1477,N_19297,N_19303);
and UO_1478 (O_1478,N_18654,N_19705);
and UO_1479 (O_1479,N_18410,N_19465);
or UO_1480 (O_1480,N_19114,N_19708);
and UO_1481 (O_1481,N_19334,N_18083);
nand UO_1482 (O_1482,N_18872,N_18102);
nand UO_1483 (O_1483,N_18587,N_19685);
nor UO_1484 (O_1484,N_18256,N_18800);
nor UO_1485 (O_1485,N_19605,N_19380);
and UO_1486 (O_1486,N_18979,N_18639);
and UO_1487 (O_1487,N_19478,N_19638);
and UO_1488 (O_1488,N_19116,N_18161);
and UO_1489 (O_1489,N_19753,N_18498);
and UO_1490 (O_1490,N_19985,N_19603);
or UO_1491 (O_1491,N_19448,N_19376);
or UO_1492 (O_1492,N_19995,N_19387);
or UO_1493 (O_1493,N_19774,N_19418);
or UO_1494 (O_1494,N_18223,N_18981);
and UO_1495 (O_1495,N_18410,N_19672);
or UO_1496 (O_1496,N_18922,N_19619);
and UO_1497 (O_1497,N_19089,N_19355);
and UO_1498 (O_1498,N_19319,N_19923);
nand UO_1499 (O_1499,N_19866,N_18723);
xnor UO_1500 (O_1500,N_18784,N_19440);
nor UO_1501 (O_1501,N_18157,N_19043);
or UO_1502 (O_1502,N_19210,N_19940);
or UO_1503 (O_1503,N_18642,N_19751);
or UO_1504 (O_1504,N_18524,N_19005);
nor UO_1505 (O_1505,N_19522,N_18996);
nand UO_1506 (O_1506,N_19707,N_19354);
or UO_1507 (O_1507,N_18261,N_19803);
or UO_1508 (O_1508,N_18452,N_18492);
xnor UO_1509 (O_1509,N_19967,N_19365);
nor UO_1510 (O_1510,N_19081,N_18652);
nor UO_1511 (O_1511,N_18891,N_19271);
and UO_1512 (O_1512,N_18906,N_19534);
nand UO_1513 (O_1513,N_19604,N_18593);
nor UO_1514 (O_1514,N_19112,N_18544);
xnor UO_1515 (O_1515,N_19161,N_19902);
nor UO_1516 (O_1516,N_19370,N_19935);
nand UO_1517 (O_1517,N_18326,N_19241);
and UO_1518 (O_1518,N_19769,N_19687);
nor UO_1519 (O_1519,N_18145,N_18253);
and UO_1520 (O_1520,N_19109,N_18356);
nand UO_1521 (O_1521,N_19195,N_19510);
and UO_1522 (O_1522,N_19815,N_18960);
and UO_1523 (O_1523,N_18862,N_18411);
and UO_1524 (O_1524,N_19942,N_19744);
and UO_1525 (O_1525,N_19831,N_18060);
or UO_1526 (O_1526,N_19729,N_18364);
nand UO_1527 (O_1527,N_19040,N_19971);
or UO_1528 (O_1528,N_19478,N_18610);
and UO_1529 (O_1529,N_18874,N_18919);
and UO_1530 (O_1530,N_19761,N_19440);
nor UO_1531 (O_1531,N_19652,N_19646);
or UO_1532 (O_1532,N_18027,N_18732);
and UO_1533 (O_1533,N_19084,N_18937);
nand UO_1534 (O_1534,N_19621,N_18969);
nor UO_1535 (O_1535,N_19774,N_18938);
nor UO_1536 (O_1536,N_19680,N_18222);
nand UO_1537 (O_1537,N_18826,N_19991);
nand UO_1538 (O_1538,N_18345,N_18543);
nand UO_1539 (O_1539,N_19017,N_18467);
or UO_1540 (O_1540,N_19418,N_18416);
nand UO_1541 (O_1541,N_18870,N_18315);
and UO_1542 (O_1542,N_19300,N_19153);
nand UO_1543 (O_1543,N_18595,N_18801);
nand UO_1544 (O_1544,N_18516,N_19606);
or UO_1545 (O_1545,N_19080,N_18080);
nor UO_1546 (O_1546,N_19807,N_19133);
and UO_1547 (O_1547,N_19910,N_19865);
or UO_1548 (O_1548,N_18377,N_18755);
nand UO_1549 (O_1549,N_19423,N_19252);
or UO_1550 (O_1550,N_18243,N_18875);
or UO_1551 (O_1551,N_18996,N_19215);
or UO_1552 (O_1552,N_19606,N_19023);
nand UO_1553 (O_1553,N_18067,N_18118);
nor UO_1554 (O_1554,N_18255,N_19273);
nor UO_1555 (O_1555,N_19009,N_19776);
or UO_1556 (O_1556,N_18871,N_18380);
or UO_1557 (O_1557,N_18134,N_18626);
nor UO_1558 (O_1558,N_19594,N_18680);
and UO_1559 (O_1559,N_19740,N_19402);
nand UO_1560 (O_1560,N_18808,N_19872);
nor UO_1561 (O_1561,N_19407,N_18793);
xor UO_1562 (O_1562,N_19949,N_18980);
or UO_1563 (O_1563,N_18057,N_18229);
xor UO_1564 (O_1564,N_18661,N_18829);
nand UO_1565 (O_1565,N_19084,N_19112);
nor UO_1566 (O_1566,N_18208,N_19899);
nand UO_1567 (O_1567,N_18407,N_18654);
nor UO_1568 (O_1568,N_18947,N_19401);
or UO_1569 (O_1569,N_18849,N_18208);
xor UO_1570 (O_1570,N_18822,N_19648);
and UO_1571 (O_1571,N_19942,N_19896);
or UO_1572 (O_1572,N_18266,N_18442);
nand UO_1573 (O_1573,N_19672,N_19446);
and UO_1574 (O_1574,N_18318,N_18763);
or UO_1575 (O_1575,N_18391,N_18862);
and UO_1576 (O_1576,N_19519,N_18444);
and UO_1577 (O_1577,N_19272,N_19047);
nor UO_1578 (O_1578,N_19410,N_18779);
and UO_1579 (O_1579,N_19849,N_18487);
nand UO_1580 (O_1580,N_19930,N_19622);
and UO_1581 (O_1581,N_19359,N_19206);
and UO_1582 (O_1582,N_19998,N_18697);
nor UO_1583 (O_1583,N_18152,N_19105);
and UO_1584 (O_1584,N_18396,N_19848);
or UO_1585 (O_1585,N_18360,N_19879);
xor UO_1586 (O_1586,N_19952,N_19748);
nor UO_1587 (O_1587,N_18648,N_19575);
nor UO_1588 (O_1588,N_19321,N_19519);
nor UO_1589 (O_1589,N_18143,N_19576);
or UO_1590 (O_1590,N_19431,N_19394);
or UO_1591 (O_1591,N_18524,N_18387);
or UO_1592 (O_1592,N_18727,N_18048);
and UO_1593 (O_1593,N_18953,N_18658);
and UO_1594 (O_1594,N_18350,N_19155);
or UO_1595 (O_1595,N_18027,N_19776);
or UO_1596 (O_1596,N_19862,N_18815);
nor UO_1597 (O_1597,N_19876,N_19312);
nor UO_1598 (O_1598,N_19378,N_19761);
and UO_1599 (O_1599,N_18205,N_18864);
nand UO_1600 (O_1600,N_19714,N_18704);
or UO_1601 (O_1601,N_18111,N_18850);
nor UO_1602 (O_1602,N_19348,N_19685);
and UO_1603 (O_1603,N_19052,N_18117);
xor UO_1604 (O_1604,N_18693,N_18421);
or UO_1605 (O_1605,N_18808,N_18548);
or UO_1606 (O_1606,N_18495,N_19998);
and UO_1607 (O_1607,N_18642,N_19972);
nand UO_1608 (O_1608,N_18329,N_18859);
nor UO_1609 (O_1609,N_18358,N_19284);
or UO_1610 (O_1610,N_19869,N_18637);
or UO_1611 (O_1611,N_18809,N_18657);
or UO_1612 (O_1612,N_18084,N_19879);
and UO_1613 (O_1613,N_19992,N_18126);
nand UO_1614 (O_1614,N_19982,N_19753);
and UO_1615 (O_1615,N_19322,N_18588);
or UO_1616 (O_1616,N_18935,N_18090);
xor UO_1617 (O_1617,N_18034,N_19787);
or UO_1618 (O_1618,N_18745,N_19335);
nor UO_1619 (O_1619,N_18977,N_19332);
nor UO_1620 (O_1620,N_18535,N_18185);
nand UO_1621 (O_1621,N_19204,N_18297);
or UO_1622 (O_1622,N_18224,N_18765);
or UO_1623 (O_1623,N_19028,N_19812);
nor UO_1624 (O_1624,N_18207,N_18198);
xor UO_1625 (O_1625,N_18576,N_19276);
nand UO_1626 (O_1626,N_18499,N_18285);
or UO_1627 (O_1627,N_18909,N_18948);
nor UO_1628 (O_1628,N_19952,N_19309);
nor UO_1629 (O_1629,N_18929,N_19935);
and UO_1630 (O_1630,N_19525,N_19728);
or UO_1631 (O_1631,N_19794,N_19752);
xor UO_1632 (O_1632,N_19391,N_18628);
nor UO_1633 (O_1633,N_19729,N_19263);
nor UO_1634 (O_1634,N_19826,N_19760);
nand UO_1635 (O_1635,N_19893,N_19848);
or UO_1636 (O_1636,N_19461,N_19284);
xor UO_1637 (O_1637,N_19027,N_19982);
xnor UO_1638 (O_1638,N_19380,N_18871);
nor UO_1639 (O_1639,N_18545,N_19549);
nor UO_1640 (O_1640,N_19225,N_18913);
xnor UO_1641 (O_1641,N_19014,N_18371);
or UO_1642 (O_1642,N_18316,N_18528);
or UO_1643 (O_1643,N_18471,N_19844);
or UO_1644 (O_1644,N_18547,N_19025);
or UO_1645 (O_1645,N_19470,N_19593);
or UO_1646 (O_1646,N_18332,N_18441);
and UO_1647 (O_1647,N_19092,N_19509);
or UO_1648 (O_1648,N_18034,N_19765);
nand UO_1649 (O_1649,N_18548,N_19810);
nand UO_1650 (O_1650,N_18324,N_18184);
nand UO_1651 (O_1651,N_19169,N_19971);
or UO_1652 (O_1652,N_19567,N_19533);
nand UO_1653 (O_1653,N_18279,N_18720);
or UO_1654 (O_1654,N_18720,N_18474);
nand UO_1655 (O_1655,N_19817,N_18567);
nand UO_1656 (O_1656,N_19863,N_19445);
nor UO_1657 (O_1657,N_19510,N_18513);
and UO_1658 (O_1658,N_19691,N_19682);
nand UO_1659 (O_1659,N_19213,N_18868);
or UO_1660 (O_1660,N_18660,N_19393);
and UO_1661 (O_1661,N_19106,N_19021);
or UO_1662 (O_1662,N_18977,N_19803);
and UO_1663 (O_1663,N_18419,N_19977);
or UO_1664 (O_1664,N_19620,N_19872);
nand UO_1665 (O_1665,N_19591,N_18333);
xor UO_1666 (O_1666,N_18498,N_19534);
and UO_1667 (O_1667,N_18770,N_19474);
nor UO_1668 (O_1668,N_19544,N_19810);
or UO_1669 (O_1669,N_18817,N_19328);
or UO_1670 (O_1670,N_18748,N_18413);
nand UO_1671 (O_1671,N_18905,N_18456);
and UO_1672 (O_1672,N_19665,N_19237);
nor UO_1673 (O_1673,N_19364,N_18226);
nand UO_1674 (O_1674,N_18811,N_18235);
or UO_1675 (O_1675,N_18430,N_19869);
nand UO_1676 (O_1676,N_19603,N_19610);
nor UO_1677 (O_1677,N_18195,N_19466);
and UO_1678 (O_1678,N_19350,N_19854);
nand UO_1679 (O_1679,N_19968,N_18637);
nand UO_1680 (O_1680,N_18351,N_18378);
or UO_1681 (O_1681,N_18528,N_18334);
or UO_1682 (O_1682,N_18177,N_19612);
nor UO_1683 (O_1683,N_18092,N_18578);
nor UO_1684 (O_1684,N_19068,N_18874);
and UO_1685 (O_1685,N_18188,N_18721);
or UO_1686 (O_1686,N_19835,N_18962);
or UO_1687 (O_1687,N_18584,N_19470);
nand UO_1688 (O_1688,N_18865,N_19833);
nand UO_1689 (O_1689,N_18892,N_19116);
or UO_1690 (O_1690,N_19893,N_18757);
or UO_1691 (O_1691,N_18875,N_18123);
nand UO_1692 (O_1692,N_19538,N_18490);
nand UO_1693 (O_1693,N_19841,N_19995);
nand UO_1694 (O_1694,N_18095,N_19872);
nor UO_1695 (O_1695,N_18216,N_19677);
nor UO_1696 (O_1696,N_19777,N_19119);
or UO_1697 (O_1697,N_18430,N_19301);
nand UO_1698 (O_1698,N_18798,N_19012);
xnor UO_1699 (O_1699,N_18586,N_18934);
nor UO_1700 (O_1700,N_18822,N_19153);
and UO_1701 (O_1701,N_18753,N_18326);
or UO_1702 (O_1702,N_19970,N_19753);
and UO_1703 (O_1703,N_19967,N_18415);
and UO_1704 (O_1704,N_19295,N_18313);
or UO_1705 (O_1705,N_19725,N_18013);
or UO_1706 (O_1706,N_18620,N_18704);
and UO_1707 (O_1707,N_18785,N_18392);
and UO_1708 (O_1708,N_18549,N_19556);
or UO_1709 (O_1709,N_19135,N_18412);
nand UO_1710 (O_1710,N_18773,N_18595);
or UO_1711 (O_1711,N_18596,N_18869);
and UO_1712 (O_1712,N_18518,N_19827);
nor UO_1713 (O_1713,N_19271,N_18002);
and UO_1714 (O_1714,N_19773,N_18738);
nand UO_1715 (O_1715,N_19287,N_19081);
or UO_1716 (O_1716,N_19214,N_18378);
nor UO_1717 (O_1717,N_19792,N_18884);
nand UO_1718 (O_1718,N_19622,N_19392);
xor UO_1719 (O_1719,N_18022,N_19748);
xnor UO_1720 (O_1720,N_19201,N_18247);
xor UO_1721 (O_1721,N_19892,N_18916);
or UO_1722 (O_1722,N_18938,N_19977);
and UO_1723 (O_1723,N_18726,N_19747);
nand UO_1724 (O_1724,N_18210,N_18176);
xor UO_1725 (O_1725,N_19372,N_19959);
or UO_1726 (O_1726,N_18843,N_19369);
nand UO_1727 (O_1727,N_19414,N_18354);
and UO_1728 (O_1728,N_18480,N_18655);
or UO_1729 (O_1729,N_19149,N_19933);
nand UO_1730 (O_1730,N_18016,N_18336);
and UO_1731 (O_1731,N_18438,N_19993);
and UO_1732 (O_1732,N_18576,N_18774);
nor UO_1733 (O_1733,N_19933,N_18773);
xor UO_1734 (O_1734,N_18650,N_19992);
or UO_1735 (O_1735,N_19639,N_19487);
or UO_1736 (O_1736,N_18785,N_18794);
or UO_1737 (O_1737,N_19066,N_19061);
and UO_1738 (O_1738,N_19522,N_19568);
and UO_1739 (O_1739,N_19220,N_18151);
nor UO_1740 (O_1740,N_18897,N_19845);
and UO_1741 (O_1741,N_19331,N_19692);
and UO_1742 (O_1742,N_18266,N_18226);
nor UO_1743 (O_1743,N_18979,N_19100);
xor UO_1744 (O_1744,N_18190,N_18475);
nand UO_1745 (O_1745,N_18959,N_18000);
nor UO_1746 (O_1746,N_18803,N_18390);
xnor UO_1747 (O_1747,N_18285,N_18215);
nand UO_1748 (O_1748,N_18677,N_18614);
and UO_1749 (O_1749,N_18387,N_19051);
or UO_1750 (O_1750,N_18507,N_19134);
nand UO_1751 (O_1751,N_18725,N_19216);
or UO_1752 (O_1752,N_18042,N_19994);
and UO_1753 (O_1753,N_18538,N_19284);
or UO_1754 (O_1754,N_18347,N_18953);
and UO_1755 (O_1755,N_18199,N_18259);
and UO_1756 (O_1756,N_19442,N_19057);
or UO_1757 (O_1757,N_19039,N_19310);
nand UO_1758 (O_1758,N_19390,N_18118);
nor UO_1759 (O_1759,N_19247,N_18776);
nand UO_1760 (O_1760,N_18033,N_18177);
or UO_1761 (O_1761,N_18043,N_18341);
and UO_1762 (O_1762,N_19661,N_19904);
nand UO_1763 (O_1763,N_18474,N_19380);
nand UO_1764 (O_1764,N_19199,N_18391);
xor UO_1765 (O_1765,N_19496,N_18287);
nor UO_1766 (O_1766,N_19804,N_19219);
and UO_1767 (O_1767,N_18984,N_18989);
nand UO_1768 (O_1768,N_18885,N_19209);
nor UO_1769 (O_1769,N_18456,N_19772);
nor UO_1770 (O_1770,N_19598,N_18884);
and UO_1771 (O_1771,N_18221,N_19498);
or UO_1772 (O_1772,N_19542,N_18950);
or UO_1773 (O_1773,N_19670,N_19433);
or UO_1774 (O_1774,N_19285,N_19449);
and UO_1775 (O_1775,N_18946,N_19609);
and UO_1776 (O_1776,N_18268,N_19554);
and UO_1777 (O_1777,N_19840,N_18541);
and UO_1778 (O_1778,N_18416,N_19520);
nor UO_1779 (O_1779,N_19039,N_18613);
nand UO_1780 (O_1780,N_18832,N_18902);
nand UO_1781 (O_1781,N_18927,N_19593);
nor UO_1782 (O_1782,N_18446,N_19679);
or UO_1783 (O_1783,N_18063,N_18602);
or UO_1784 (O_1784,N_18492,N_18111);
or UO_1785 (O_1785,N_19902,N_18465);
xnor UO_1786 (O_1786,N_19887,N_18802);
xnor UO_1787 (O_1787,N_18715,N_19215);
nor UO_1788 (O_1788,N_19262,N_18421);
nand UO_1789 (O_1789,N_19669,N_19968);
or UO_1790 (O_1790,N_18520,N_19415);
nor UO_1791 (O_1791,N_18573,N_18396);
or UO_1792 (O_1792,N_19587,N_19205);
nor UO_1793 (O_1793,N_18176,N_18567);
or UO_1794 (O_1794,N_18279,N_19309);
nor UO_1795 (O_1795,N_19601,N_18122);
or UO_1796 (O_1796,N_19524,N_19908);
nor UO_1797 (O_1797,N_19299,N_19991);
nand UO_1798 (O_1798,N_19972,N_18737);
nand UO_1799 (O_1799,N_19565,N_18293);
xor UO_1800 (O_1800,N_18720,N_18241);
nor UO_1801 (O_1801,N_19917,N_18495);
nor UO_1802 (O_1802,N_19240,N_18704);
and UO_1803 (O_1803,N_18636,N_18964);
nand UO_1804 (O_1804,N_19685,N_18535);
or UO_1805 (O_1805,N_19170,N_18063);
nand UO_1806 (O_1806,N_18086,N_19377);
nand UO_1807 (O_1807,N_19298,N_18282);
nand UO_1808 (O_1808,N_19560,N_18733);
and UO_1809 (O_1809,N_19041,N_19045);
and UO_1810 (O_1810,N_18988,N_19579);
nor UO_1811 (O_1811,N_18042,N_18967);
or UO_1812 (O_1812,N_18481,N_18442);
nand UO_1813 (O_1813,N_18453,N_18279);
xnor UO_1814 (O_1814,N_19323,N_19947);
or UO_1815 (O_1815,N_18709,N_18646);
or UO_1816 (O_1816,N_19866,N_19027);
nand UO_1817 (O_1817,N_19047,N_19171);
xor UO_1818 (O_1818,N_19901,N_18391);
or UO_1819 (O_1819,N_18819,N_19429);
xor UO_1820 (O_1820,N_18643,N_19901);
and UO_1821 (O_1821,N_18921,N_19072);
nand UO_1822 (O_1822,N_19716,N_18938);
nor UO_1823 (O_1823,N_18254,N_18427);
nor UO_1824 (O_1824,N_18610,N_18285);
nand UO_1825 (O_1825,N_18470,N_19842);
and UO_1826 (O_1826,N_18153,N_18251);
and UO_1827 (O_1827,N_18982,N_18782);
or UO_1828 (O_1828,N_18113,N_19582);
and UO_1829 (O_1829,N_18724,N_19373);
nand UO_1830 (O_1830,N_19757,N_19325);
and UO_1831 (O_1831,N_19314,N_19603);
nand UO_1832 (O_1832,N_18085,N_19215);
nand UO_1833 (O_1833,N_19884,N_18956);
and UO_1834 (O_1834,N_19473,N_18224);
and UO_1835 (O_1835,N_18901,N_19692);
and UO_1836 (O_1836,N_19673,N_18323);
nor UO_1837 (O_1837,N_19230,N_19735);
and UO_1838 (O_1838,N_18897,N_18896);
nand UO_1839 (O_1839,N_18478,N_18533);
xnor UO_1840 (O_1840,N_19559,N_18607);
and UO_1841 (O_1841,N_19445,N_18025);
nand UO_1842 (O_1842,N_18730,N_18468);
nor UO_1843 (O_1843,N_19512,N_19853);
and UO_1844 (O_1844,N_18663,N_18269);
xor UO_1845 (O_1845,N_19197,N_18967);
and UO_1846 (O_1846,N_18775,N_18001);
or UO_1847 (O_1847,N_19281,N_18974);
or UO_1848 (O_1848,N_18061,N_19510);
or UO_1849 (O_1849,N_19461,N_18345);
and UO_1850 (O_1850,N_18300,N_19926);
or UO_1851 (O_1851,N_18517,N_18527);
nor UO_1852 (O_1852,N_19068,N_19243);
or UO_1853 (O_1853,N_18813,N_19567);
nor UO_1854 (O_1854,N_19899,N_18296);
nor UO_1855 (O_1855,N_19469,N_19367);
and UO_1856 (O_1856,N_19351,N_18115);
or UO_1857 (O_1857,N_19794,N_18416);
and UO_1858 (O_1858,N_19296,N_18398);
and UO_1859 (O_1859,N_18604,N_18235);
or UO_1860 (O_1860,N_18721,N_18122);
nor UO_1861 (O_1861,N_19322,N_19801);
nand UO_1862 (O_1862,N_19634,N_18503);
or UO_1863 (O_1863,N_19395,N_18617);
and UO_1864 (O_1864,N_19577,N_18396);
or UO_1865 (O_1865,N_19650,N_19353);
nand UO_1866 (O_1866,N_18031,N_19494);
and UO_1867 (O_1867,N_18675,N_18138);
xor UO_1868 (O_1868,N_19001,N_19488);
nand UO_1869 (O_1869,N_19868,N_18666);
nand UO_1870 (O_1870,N_18379,N_19407);
and UO_1871 (O_1871,N_19956,N_18308);
xor UO_1872 (O_1872,N_18590,N_18921);
nor UO_1873 (O_1873,N_18544,N_19624);
or UO_1874 (O_1874,N_19850,N_19872);
nor UO_1875 (O_1875,N_18560,N_19614);
nor UO_1876 (O_1876,N_19485,N_19125);
or UO_1877 (O_1877,N_18768,N_18471);
nor UO_1878 (O_1878,N_19328,N_18810);
or UO_1879 (O_1879,N_18537,N_19833);
nand UO_1880 (O_1880,N_19372,N_18343);
or UO_1881 (O_1881,N_18427,N_18009);
or UO_1882 (O_1882,N_18147,N_18711);
or UO_1883 (O_1883,N_19882,N_19808);
nor UO_1884 (O_1884,N_19016,N_19918);
or UO_1885 (O_1885,N_19315,N_19880);
nand UO_1886 (O_1886,N_19170,N_18297);
nand UO_1887 (O_1887,N_18431,N_18662);
nor UO_1888 (O_1888,N_18818,N_18561);
or UO_1889 (O_1889,N_19770,N_18360);
nor UO_1890 (O_1890,N_19372,N_18177);
and UO_1891 (O_1891,N_19521,N_19570);
nor UO_1892 (O_1892,N_18839,N_18316);
nand UO_1893 (O_1893,N_19145,N_19141);
or UO_1894 (O_1894,N_18917,N_18480);
and UO_1895 (O_1895,N_18931,N_19724);
and UO_1896 (O_1896,N_18538,N_18505);
or UO_1897 (O_1897,N_18919,N_19789);
and UO_1898 (O_1898,N_19981,N_18127);
and UO_1899 (O_1899,N_19027,N_18419);
nor UO_1900 (O_1900,N_18446,N_18170);
nand UO_1901 (O_1901,N_19830,N_18455);
nand UO_1902 (O_1902,N_19571,N_19014);
nand UO_1903 (O_1903,N_18137,N_19065);
nand UO_1904 (O_1904,N_18005,N_19331);
nor UO_1905 (O_1905,N_18047,N_19777);
or UO_1906 (O_1906,N_18767,N_19728);
nor UO_1907 (O_1907,N_19973,N_18127);
xnor UO_1908 (O_1908,N_18976,N_19854);
nand UO_1909 (O_1909,N_18480,N_18161);
and UO_1910 (O_1910,N_19610,N_18820);
xnor UO_1911 (O_1911,N_18105,N_19832);
and UO_1912 (O_1912,N_18805,N_18848);
and UO_1913 (O_1913,N_19441,N_19564);
nand UO_1914 (O_1914,N_19308,N_19804);
nand UO_1915 (O_1915,N_19570,N_19717);
or UO_1916 (O_1916,N_19700,N_18794);
nand UO_1917 (O_1917,N_18709,N_19200);
and UO_1918 (O_1918,N_19903,N_18782);
and UO_1919 (O_1919,N_19793,N_18726);
nand UO_1920 (O_1920,N_19090,N_19593);
nor UO_1921 (O_1921,N_18448,N_18465);
or UO_1922 (O_1922,N_19203,N_18796);
nand UO_1923 (O_1923,N_18725,N_18060);
or UO_1924 (O_1924,N_18205,N_18272);
or UO_1925 (O_1925,N_18631,N_19567);
or UO_1926 (O_1926,N_19893,N_18132);
nor UO_1927 (O_1927,N_19689,N_18974);
and UO_1928 (O_1928,N_18305,N_19006);
nand UO_1929 (O_1929,N_19298,N_18168);
xnor UO_1930 (O_1930,N_19024,N_18793);
or UO_1931 (O_1931,N_19238,N_18862);
and UO_1932 (O_1932,N_18294,N_19904);
or UO_1933 (O_1933,N_18622,N_19927);
nand UO_1934 (O_1934,N_19052,N_18368);
nand UO_1935 (O_1935,N_18412,N_19647);
or UO_1936 (O_1936,N_18621,N_18917);
nand UO_1937 (O_1937,N_19528,N_19084);
nor UO_1938 (O_1938,N_18556,N_18030);
nor UO_1939 (O_1939,N_18794,N_18947);
and UO_1940 (O_1940,N_19073,N_19182);
nor UO_1941 (O_1941,N_18968,N_19813);
nand UO_1942 (O_1942,N_18163,N_19344);
nand UO_1943 (O_1943,N_19352,N_19173);
and UO_1944 (O_1944,N_19775,N_18106);
and UO_1945 (O_1945,N_19036,N_18808);
nand UO_1946 (O_1946,N_19157,N_19192);
or UO_1947 (O_1947,N_19376,N_19527);
or UO_1948 (O_1948,N_18091,N_18636);
and UO_1949 (O_1949,N_19439,N_18188);
nor UO_1950 (O_1950,N_19536,N_19775);
nand UO_1951 (O_1951,N_19045,N_19318);
xnor UO_1952 (O_1952,N_18052,N_19672);
and UO_1953 (O_1953,N_18197,N_19323);
xnor UO_1954 (O_1954,N_19559,N_18898);
xor UO_1955 (O_1955,N_19809,N_19094);
nand UO_1956 (O_1956,N_19696,N_18327);
or UO_1957 (O_1957,N_18068,N_18940);
nand UO_1958 (O_1958,N_18281,N_19379);
nor UO_1959 (O_1959,N_19405,N_19836);
nand UO_1960 (O_1960,N_18594,N_18220);
nor UO_1961 (O_1961,N_18322,N_18223);
nand UO_1962 (O_1962,N_19848,N_18946);
and UO_1963 (O_1963,N_18458,N_19609);
and UO_1964 (O_1964,N_19562,N_19125);
nor UO_1965 (O_1965,N_19636,N_18815);
and UO_1966 (O_1966,N_19839,N_18777);
and UO_1967 (O_1967,N_19556,N_18809);
nand UO_1968 (O_1968,N_19979,N_18595);
or UO_1969 (O_1969,N_18258,N_19773);
and UO_1970 (O_1970,N_18598,N_19456);
nand UO_1971 (O_1971,N_19893,N_19605);
xor UO_1972 (O_1972,N_18672,N_19087);
xor UO_1973 (O_1973,N_18045,N_19942);
xor UO_1974 (O_1974,N_18639,N_19108);
or UO_1975 (O_1975,N_19257,N_19452);
or UO_1976 (O_1976,N_19460,N_19532);
nor UO_1977 (O_1977,N_19186,N_19532);
nor UO_1978 (O_1978,N_19259,N_18074);
xnor UO_1979 (O_1979,N_19623,N_18132);
nor UO_1980 (O_1980,N_18758,N_19985);
and UO_1981 (O_1981,N_18908,N_18963);
nand UO_1982 (O_1982,N_18444,N_19497);
nor UO_1983 (O_1983,N_18979,N_19943);
nand UO_1984 (O_1984,N_18667,N_18485);
and UO_1985 (O_1985,N_19695,N_18500);
nand UO_1986 (O_1986,N_18046,N_18097);
and UO_1987 (O_1987,N_19926,N_19174);
nand UO_1988 (O_1988,N_19236,N_19307);
nor UO_1989 (O_1989,N_19101,N_18404);
nor UO_1990 (O_1990,N_18025,N_18001);
nor UO_1991 (O_1991,N_18383,N_18285);
xor UO_1992 (O_1992,N_19141,N_18763);
or UO_1993 (O_1993,N_19744,N_18656);
or UO_1994 (O_1994,N_18671,N_19770);
nand UO_1995 (O_1995,N_19648,N_18517);
xor UO_1996 (O_1996,N_18111,N_19922);
nor UO_1997 (O_1997,N_19153,N_19943);
nor UO_1998 (O_1998,N_19108,N_19043);
and UO_1999 (O_1999,N_19806,N_18310);
or UO_2000 (O_2000,N_19785,N_19990);
nand UO_2001 (O_2001,N_19275,N_19232);
and UO_2002 (O_2002,N_18648,N_19901);
or UO_2003 (O_2003,N_19541,N_19790);
nand UO_2004 (O_2004,N_19838,N_19784);
or UO_2005 (O_2005,N_18911,N_18041);
nand UO_2006 (O_2006,N_18805,N_18419);
xor UO_2007 (O_2007,N_19138,N_19337);
and UO_2008 (O_2008,N_18393,N_18336);
or UO_2009 (O_2009,N_19856,N_19880);
nor UO_2010 (O_2010,N_19412,N_18379);
or UO_2011 (O_2011,N_19079,N_19164);
xor UO_2012 (O_2012,N_18136,N_19069);
nand UO_2013 (O_2013,N_19386,N_19893);
and UO_2014 (O_2014,N_18454,N_19862);
nor UO_2015 (O_2015,N_19197,N_18260);
or UO_2016 (O_2016,N_18320,N_19788);
and UO_2017 (O_2017,N_18451,N_18818);
nor UO_2018 (O_2018,N_18351,N_18011);
and UO_2019 (O_2019,N_18453,N_18190);
nor UO_2020 (O_2020,N_19902,N_18513);
and UO_2021 (O_2021,N_19477,N_19483);
and UO_2022 (O_2022,N_18929,N_18570);
nor UO_2023 (O_2023,N_19056,N_19424);
or UO_2024 (O_2024,N_19725,N_18568);
nor UO_2025 (O_2025,N_19211,N_19117);
and UO_2026 (O_2026,N_18773,N_19725);
nand UO_2027 (O_2027,N_18719,N_18385);
nor UO_2028 (O_2028,N_18504,N_18619);
nor UO_2029 (O_2029,N_18194,N_19955);
nor UO_2030 (O_2030,N_19931,N_18902);
and UO_2031 (O_2031,N_19193,N_18966);
nand UO_2032 (O_2032,N_18584,N_19649);
and UO_2033 (O_2033,N_19874,N_18733);
xnor UO_2034 (O_2034,N_18718,N_19319);
nor UO_2035 (O_2035,N_19889,N_19027);
or UO_2036 (O_2036,N_19837,N_18136);
nor UO_2037 (O_2037,N_19830,N_18944);
nand UO_2038 (O_2038,N_18308,N_19439);
nor UO_2039 (O_2039,N_19292,N_19524);
nand UO_2040 (O_2040,N_19332,N_18502);
nand UO_2041 (O_2041,N_19137,N_19084);
nor UO_2042 (O_2042,N_18946,N_18864);
nor UO_2043 (O_2043,N_18478,N_18199);
nor UO_2044 (O_2044,N_19254,N_19388);
and UO_2045 (O_2045,N_18956,N_19430);
and UO_2046 (O_2046,N_18633,N_19653);
and UO_2047 (O_2047,N_19956,N_18979);
or UO_2048 (O_2048,N_18667,N_19189);
nand UO_2049 (O_2049,N_18220,N_19395);
xor UO_2050 (O_2050,N_19981,N_19254);
and UO_2051 (O_2051,N_18082,N_19017);
or UO_2052 (O_2052,N_19132,N_19940);
nand UO_2053 (O_2053,N_18887,N_19640);
xnor UO_2054 (O_2054,N_18909,N_19332);
nor UO_2055 (O_2055,N_18273,N_19616);
xor UO_2056 (O_2056,N_19991,N_19789);
nor UO_2057 (O_2057,N_18868,N_18247);
nand UO_2058 (O_2058,N_19737,N_18968);
xnor UO_2059 (O_2059,N_18029,N_18601);
nor UO_2060 (O_2060,N_19483,N_18182);
nor UO_2061 (O_2061,N_18016,N_18391);
nor UO_2062 (O_2062,N_19260,N_19718);
nand UO_2063 (O_2063,N_18220,N_18154);
nand UO_2064 (O_2064,N_18539,N_19020);
nor UO_2065 (O_2065,N_19531,N_19100);
or UO_2066 (O_2066,N_19677,N_19958);
nor UO_2067 (O_2067,N_19339,N_19017);
nor UO_2068 (O_2068,N_19441,N_19881);
nand UO_2069 (O_2069,N_19148,N_19312);
or UO_2070 (O_2070,N_18264,N_19261);
nand UO_2071 (O_2071,N_19275,N_18170);
nand UO_2072 (O_2072,N_18284,N_19596);
and UO_2073 (O_2073,N_19783,N_18109);
xnor UO_2074 (O_2074,N_19355,N_18419);
xor UO_2075 (O_2075,N_19727,N_18905);
nand UO_2076 (O_2076,N_18847,N_18629);
and UO_2077 (O_2077,N_18951,N_19858);
and UO_2078 (O_2078,N_18057,N_19194);
or UO_2079 (O_2079,N_19574,N_18073);
nor UO_2080 (O_2080,N_18529,N_18052);
or UO_2081 (O_2081,N_19958,N_19974);
nand UO_2082 (O_2082,N_18513,N_19924);
and UO_2083 (O_2083,N_19351,N_19622);
and UO_2084 (O_2084,N_19381,N_19363);
and UO_2085 (O_2085,N_19168,N_19427);
nor UO_2086 (O_2086,N_19916,N_18984);
xor UO_2087 (O_2087,N_18654,N_19929);
and UO_2088 (O_2088,N_18012,N_18468);
nand UO_2089 (O_2089,N_18484,N_19576);
and UO_2090 (O_2090,N_19247,N_18224);
nor UO_2091 (O_2091,N_18371,N_18775);
nor UO_2092 (O_2092,N_19314,N_19845);
or UO_2093 (O_2093,N_18938,N_19561);
or UO_2094 (O_2094,N_19404,N_18236);
or UO_2095 (O_2095,N_19792,N_18738);
and UO_2096 (O_2096,N_19344,N_19316);
nor UO_2097 (O_2097,N_19080,N_18414);
and UO_2098 (O_2098,N_18782,N_18562);
nand UO_2099 (O_2099,N_18749,N_18130);
nor UO_2100 (O_2100,N_19311,N_19842);
nand UO_2101 (O_2101,N_19061,N_19386);
and UO_2102 (O_2102,N_18373,N_19903);
or UO_2103 (O_2103,N_19389,N_18858);
nor UO_2104 (O_2104,N_18972,N_19672);
and UO_2105 (O_2105,N_19516,N_18818);
nor UO_2106 (O_2106,N_19430,N_18657);
nand UO_2107 (O_2107,N_19132,N_18101);
and UO_2108 (O_2108,N_18169,N_18656);
nor UO_2109 (O_2109,N_18995,N_19927);
or UO_2110 (O_2110,N_19240,N_18089);
or UO_2111 (O_2111,N_19078,N_19580);
or UO_2112 (O_2112,N_19820,N_19670);
or UO_2113 (O_2113,N_18210,N_18311);
nand UO_2114 (O_2114,N_18871,N_19489);
and UO_2115 (O_2115,N_18903,N_18790);
nor UO_2116 (O_2116,N_19971,N_19240);
nor UO_2117 (O_2117,N_18794,N_18561);
or UO_2118 (O_2118,N_18973,N_19955);
or UO_2119 (O_2119,N_18857,N_19404);
nor UO_2120 (O_2120,N_18612,N_18858);
nand UO_2121 (O_2121,N_18111,N_18502);
xor UO_2122 (O_2122,N_18068,N_18455);
and UO_2123 (O_2123,N_19976,N_18004);
nand UO_2124 (O_2124,N_19002,N_19182);
nor UO_2125 (O_2125,N_18179,N_19144);
nand UO_2126 (O_2126,N_19198,N_18025);
nor UO_2127 (O_2127,N_18244,N_18193);
and UO_2128 (O_2128,N_18639,N_18306);
and UO_2129 (O_2129,N_18211,N_18861);
nand UO_2130 (O_2130,N_19170,N_18879);
nor UO_2131 (O_2131,N_19424,N_18317);
xnor UO_2132 (O_2132,N_18896,N_18056);
nand UO_2133 (O_2133,N_18406,N_19810);
or UO_2134 (O_2134,N_18660,N_18754);
or UO_2135 (O_2135,N_18272,N_18628);
nor UO_2136 (O_2136,N_19997,N_18920);
nand UO_2137 (O_2137,N_19958,N_19385);
nand UO_2138 (O_2138,N_18589,N_19679);
nor UO_2139 (O_2139,N_19754,N_18543);
nand UO_2140 (O_2140,N_19539,N_19034);
nand UO_2141 (O_2141,N_19186,N_18988);
nand UO_2142 (O_2142,N_18797,N_19016);
and UO_2143 (O_2143,N_18864,N_18532);
nor UO_2144 (O_2144,N_18087,N_19097);
nand UO_2145 (O_2145,N_18931,N_18491);
nor UO_2146 (O_2146,N_18026,N_19428);
and UO_2147 (O_2147,N_19686,N_19244);
nor UO_2148 (O_2148,N_19941,N_19897);
nand UO_2149 (O_2149,N_19542,N_19949);
nor UO_2150 (O_2150,N_19761,N_18472);
nor UO_2151 (O_2151,N_19237,N_18238);
nor UO_2152 (O_2152,N_19835,N_19751);
nor UO_2153 (O_2153,N_18486,N_19012);
and UO_2154 (O_2154,N_18815,N_18282);
nor UO_2155 (O_2155,N_19330,N_18954);
or UO_2156 (O_2156,N_19544,N_19434);
and UO_2157 (O_2157,N_19964,N_19531);
or UO_2158 (O_2158,N_19935,N_19655);
nand UO_2159 (O_2159,N_19032,N_18645);
and UO_2160 (O_2160,N_19322,N_19745);
or UO_2161 (O_2161,N_18933,N_18345);
and UO_2162 (O_2162,N_19258,N_18579);
nor UO_2163 (O_2163,N_18473,N_19077);
nand UO_2164 (O_2164,N_18048,N_19032);
or UO_2165 (O_2165,N_18581,N_18188);
nand UO_2166 (O_2166,N_19062,N_19179);
and UO_2167 (O_2167,N_18279,N_19673);
or UO_2168 (O_2168,N_19539,N_19268);
and UO_2169 (O_2169,N_18413,N_19715);
or UO_2170 (O_2170,N_19456,N_19607);
or UO_2171 (O_2171,N_18449,N_19126);
nor UO_2172 (O_2172,N_19933,N_19622);
xor UO_2173 (O_2173,N_18549,N_19178);
xnor UO_2174 (O_2174,N_19990,N_18007);
nor UO_2175 (O_2175,N_18785,N_19933);
and UO_2176 (O_2176,N_18716,N_19669);
and UO_2177 (O_2177,N_18970,N_18653);
nor UO_2178 (O_2178,N_19678,N_18808);
nor UO_2179 (O_2179,N_18717,N_18640);
nor UO_2180 (O_2180,N_18515,N_18607);
xnor UO_2181 (O_2181,N_19517,N_19734);
xor UO_2182 (O_2182,N_18449,N_19361);
nor UO_2183 (O_2183,N_18857,N_19970);
nand UO_2184 (O_2184,N_18651,N_19781);
and UO_2185 (O_2185,N_18811,N_19032);
and UO_2186 (O_2186,N_19542,N_19796);
nor UO_2187 (O_2187,N_18422,N_18087);
nor UO_2188 (O_2188,N_18930,N_19091);
xor UO_2189 (O_2189,N_19371,N_18882);
xor UO_2190 (O_2190,N_18452,N_19709);
nor UO_2191 (O_2191,N_19512,N_19948);
or UO_2192 (O_2192,N_18261,N_19429);
and UO_2193 (O_2193,N_19528,N_18884);
xnor UO_2194 (O_2194,N_19435,N_18773);
and UO_2195 (O_2195,N_18389,N_18122);
or UO_2196 (O_2196,N_18004,N_19393);
or UO_2197 (O_2197,N_19749,N_18877);
xnor UO_2198 (O_2198,N_19852,N_19379);
or UO_2199 (O_2199,N_19721,N_18564);
or UO_2200 (O_2200,N_19214,N_18014);
nand UO_2201 (O_2201,N_19147,N_18588);
or UO_2202 (O_2202,N_18138,N_19022);
nand UO_2203 (O_2203,N_18032,N_18607);
or UO_2204 (O_2204,N_19362,N_18233);
and UO_2205 (O_2205,N_18571,N_18304);
nor UO_2206 (O_2206,N_18159,N_18089);
nor UO_2207 (O_2207,N_19962,N_18573);
and UO_2208 (O_2208,N_19310,N_18611);
and UO_2209 (O_2209,N_18552,N_19805);
and UO_2210 (O_2210,N_19531,N_19521);
nand UO_2211 (O_2211,N_19853,N_18885);
and UO_2212 (O_2212,N_18489,N_19630);
and UO_2213 (O_2213,N_18948,N_19610);
nand UO_2214 (O_2214,N_19927,N_19239);
nand UO_2215 (O_2215,N_18721,N_18343);
and UO_2216 (O_2216,N_18955,N_19732);
and UO_2217 (O_2217,N_19593,N_18979);
nand UO_2218 (O_2218,N_19719,N_18910);
and UO_2219 (O_2219,N_19034,N_18977);
and UO_2220 (O_2220,N_19401,N_18687);
nor UO_2221 (O_2221,N_19861,N_18398);
nand UO_2222 (O_2222,N_19067,N_19419);
and UO_2223 (O_2223,N_18107,N_19192);
xor UO_2224 (O_2224,N_19469,N_18369);
or UO_2225 (O_2225,N_18156,N_19096);
and UO_2226 (O_2226,N_19221,N_19538);
and UO_2227 (O_2227,N_19650,N_19294);
nor UO_2228 (O_2228,N_19811,N_18689);
nor UO_2229 (O_2229,N_19373,N_19953);
nor UO_2230 (O_2230,N_18045,N_18415);
nor UO_2231 (O_2231,N_19964,N_18857);
and UO_2232 (O_2232,N_19736,N_19113);
nor UO_2233 (O_2233,N_18060,N_18845);
or UO_2234 (O_2234,N_19805,N_19090);
and UO_2235 (O_2235,N_18540,N_18863);
nand UO_2236 (O_2236,N_19049,N_18852);
nor UO_2237 (O_2237,N_18580,N_19626);
nand UO_2238 (O_2238,N_18898,N_19869);
xor UO_2239 (O_2239,N_19640,N_19878);
nand UO_2240 (O_2240,N_19893,N_19299);
or UO_2241 (O_2241,N_19225,N_19477);
or UO_2242 (O_2242,N_19582,N_19888);
and UO_2243 (O_2243,N_19110,N_18091);
nor UO_2244 (O_2244,N_18385,N_18567);
xnor UO_2245 (O_2245,N_18326,N_18566);
nand UO_2246 (O_2246,N_18624,N_18789);
nor UO_2247 (O_2247,N_18321,N_18610);
or UO_2248 (O_2248,N_19781,N_19215);
nand UO_2249 (O_2249,N_19330,N_19742);
nor UO_2250 (O_2250,N_19562,N_19464);
nand UO_2251 (O_2251,N_19518,N_19714);
and UO_2252 (O_2252,N_19127,N_19548);
xnor UO_2253 (O_2253,N_19918,N_19559);
nand UO_2254 (O_2254,N_19187,N_18063);
nor UO_2255 (O_2255,N_18515,N_18854);
nor UO_2256 (O_2256,N_19789,N_19139);
or UO_2257 (O_2257,N_18853,N_18633);
and UO_2258 (O_2258,N_19082,N_18955);
nor UO_2259 (O_2259,N_18410,N_19445);
and UO_2260 (O_2260,N_18226,N_19980);
nand UO_2261 (O_2261,N_19462,N_19778);
and UO_2262 (O_2262,N_18677,N_19408);
or UO_2263 (O_2263,N_19935,N_19095);
xor UO_2264 (O_2264,N_18759,N_18015);
nor UO_2265 (O_2265,N_19283,N_18864);
and UO_2266 (O_2266,N_18876,N_18388);
or UO_2267 (O_2267,N_18976,N_19747);
or UO_2268 (O_2268,N_19952,N_18582);
nor UO_2269 (O_2269,N_19110,N_19174);
and UO_2270 (O_2270,N_18991,N_19681);
or UO_2271 (O_2271,N_19188,N_18999);
nor UO_2272 (O_2272,N_18971,N_19142);
nand UO_2273 (O_2273,N_18590,N_19446);
or UO_2274 (O_2274,N_18029,N_19165);
nand UO_2275 (O_2275,N_19160,N_18323);
or UO_2276 (O_2276,N_18788,N_19803);
nor UO_2277 (O_2277,N_19179,N_18145);
or UO_2278 (O_2278,N_18511,N_19675);
nor UO_2279 (O_2279,N_18740,N_18368);
nor UO_2280 (O_2280,N_19909,N_18427);
nor UO_2281 (O_2281,N_18899,N_18740);
nor UO_2282 (O_2282,N_18074,N_18329);
xor UO_2283 (O_2283,N_18237,N_18347);
or UO_2284 (O_2284,N_19845,N_18183);
and UO_2285 (O_2285,N_18386,N_18956);
nand UO_2286 (O_2286,N_18831,N_18076);
and UO_2287 (O_2287,N_19920,N_18184);
nand UO_2288 (O_2288,N_18907,N_18296);
or UO_2289 (O_2289,N_18467,N_18527);
nand UO_2290 (O_2290,N_19946,N_19943);
nor UO_2291 (O_2291,N_19073,N_18485);
xor UO_2292 (O_2292,N_19907,N_18444);
xnor UO_2293 (O_2293,N_19211,N_19893);
nand UO_2294 (O_2294,N_19400,N_19463);
nor UO_2295 (O_2295,N_19271,N_18058);
nand UO_2296 (O_2296,N_18341,N_19720);
and UO_2297 (O_2297,N_19724,N_19067);
and UO_2298 (O_2298,N_18798,N_19227);
or UO_2299 (O_2299,N_18052,N_19131);
nor UO_2300 (O_2300,N_19195,N_18113);
nor UO_2301 (O_2301,N_19130,N_18074);
or UO_2302 (O_2302,N_19215,N_18562);
and UO_2303 (O_2303,N_18053,N_18113);
or UO_2304 (O_2304,N_19884,N_19637);
nand UO_2305 (O_2305,N_19853,N_19814);
or UO_2306 (O_2306,N_18010,N_19851);
or UO_2307 (O_2307,N_19976,N_19452);
nor UO_2308 (O_2308,N_19713,N_19703);
nor UO_2309 (O_2309,N_19116,N_18869);
or UO_2310 (O_2310,N_19522,N_18287);
and UO_2311 (O_2311,N_18560,N_19814);
xor UO_2312 (O_2312,N_18514,N_18431);
and UO_2313 (O_2313,N_18134,N_18730);
and UO_2314 (O_2314,N_19734,N_19671);
nand UO_2315 (O_2315,N_18994,N_19775);
and UO_2316 (O_2316,N_18563,N_18768);
nor UO_2317 (O_2317,N_18480,N_19863);
or UO_2318 (O_2318,N_19400,N_18418);
nand UO_2319 (O_2319,N_19263,N_18112);
and UO_2320 (O_2320,N_18041,N_19680);
nor UO_2321 (O_2321,N_18252,N_19600);
nor UO_2322 (O_2322,N_18623,N_19830);
nor UO_2323 (O_2323,N_18083,N_19945);
and UO_2324 (O_2324,N_19032,N_19180);
and UO_2325 (O_2325,N_18803,N_19554);
nand UO_2326 (O_2326,N_18865,N_18739);
or UO_2327 (O_2327,N_18172,N_18504);
nand UO_2328 (O_2328,N_19637,N_19422);
and UO_2329 (O_2329,N_19975,N_18510);
and UO_2330 (O_2330,N_19784,N_19327);
nand UO_2331 (O_2331,N_19915,N_19690);
or UO_2332 (O_2332,N_19430,N_19922);
nand UO_2333 (O_2333,N_18765,N_18151);
nor UO_2334 (O_2334,N_18236,N_18638);
and UO_2335 (O_2335,N_19629,N_18190);
or UO_2336 (O_2336,N_18114,N_19801);
or UO_2337 (O_2337,N_18169,N_19105);
nor UO_2338 (O_2338,N_18536,N_18685);
or UO_2339 (O_2339,N_18220,N_19116);
and UO_2340 (O_2340,N_19720,N_18082);
and UO_2341 (O_2341,N_19331,N_19950);
and UO_2342 (O_2342,N_18071,N_18476);
nand UO_2343 (O_2343,N_18523,N_18437);
nand UO_2344 (O_2344,N_18236,N_19239);
nand UO_2345 (O_2345,N_19291,N_19665);
nand UO_2346 (O_2346,N_18722,N_19562);
or UO_2347 (O_2347,N_18415,N_18754);
or UO_2348 (O_2348,N_18292,N_18869);
nor UO_2349 (O_2349,N_19746,N_19100);
nor UO_2350 (O_2350,N_18309,N_18208);
nand UO_2351 (O_2351,N_19071,N_18209);
or UO_2352 (O_2352,N_18987,N_18510);
and UO_2353 (O_2353,N_19946,N_18918);
xnor UO_2354 (O_2354,N_19693,N_18309);
nor UO_2355 (O_2355,N_19972,N_18074);
nor UO_2356 (O_2356,N_19354,N_19009);
or UO_2357 (O_2357,N_18005,N_18564);
nand UO_2358 (O_2358,N_19045,N_19540);
and UO_2359 (O_2359,N_19677,N_18024);
or UO_2360 (O_2360,N_18261,N_19397);
nor UO_2361 (O_2361,N_19558,N_18707);
or UO_2362 (O_2362,N_19719,N_18528);
nor UO_2363 (O_2363,N_19345,N_19961);
nor UO_2364 (O_2364,N_19544,N_18580);
or UO_2365 (O_2365,N_18605,N_18972);
nand UO_2366 (O_2366,N_18939,N_18005);
nor UO_2367 (O_2367,N_18806,N_18495);
and UO_2368 (O_2368,N_18597,N_18263);
nor UO_2369 (O_2369,N_18167,N_18655);
xor UO_2370 (O_2370,N_19406,N_19989);
and UO_2371 (O_2371,N_18710,N_18584);
or UO_2372 (O_2372,N_19889,N_18078);
and UO_2373 (O_2373,N_18954,N_19235);
and UO_2374 (O_2374,N_18605,N_19050);
nand UO_2375 (O_2375,N_18651,N_19729);
and UO_2376 (O_2376,N_18798,N_18674);
nor UO_2377 (O_2377,N_18908,N_18017);
and UO_2378 (O_2378,N_19440,N_18804);
nand UO_2379 (O_2379,N_19592,N_19239);
or UO_2380 (O_2380,N_18723,N_19099);
nand UO_2381 (O_2381,N_19541,N_18584);
nor UO_2382 (O_2382,N_19356,N_18753);
and UO_2383 (O_2383,N_18107,N_19178);
xnor UO_2384 (O_2384,N_18897,N_19112);
and UO_2385 (O_2385,N_18003,N_18119);
xor UO_2386 (O_2386,N_18796,N_19454);
or UO_2387 (O_2387,N_19587,N_19985);
nand UO_2388 (O_2388,N_19173,N_18534);
xor UO_2389 (O_2389,N_19686,N_18864);
or UO_2390 (O_2390,N_18618,N_18818);
or UO_2391 (O_2391,N_19521,N_18695);
or UO_2392 (O_2392,N_18583,N_18038);
nor UO_2393 (O_2393,N_18948,N_18531);
nor UO_2394 (O_2394,N_19582,N_18620);
nor UO_2395 (O_2395,N_19611,N_18155);
or UO_2396 (O_2396,N_19267,N_19563);
and UO_2397 (O_2397,N_19895,N_18573);
and UO_2398 (O_2398,N_18214,N_19609);
and UO_2399 (O_2399,N_19958,N_19051);
nor UO_2400 (O_2400,N_19494,N_19898);
nand UO_2401 (O_2401,N_19758,N_19020);
and UO_2402 (O_2402,N_19248,N_19495);
and UO_2403 (O_2403,N_19178,N_19964);
nor UO_2404 (O_2404,N_18077,N_18272);
or UO_2405 (O_2405,N_18714,N_18500);
nor UO_2406 (O_2406,N_19125,N_19247);
nand UO_2407 (O_2407,N_19933,N_19595);
or UO_2408 (O_2408,N_18172,N_18036);
or UO_2409 (O_2409,N_18355,N_19382);
or UO_2410 (O_2410,N_18423,N_19718);
xor UO_2411 (O_2411,N_18906,N_19427);
and UO_2412 (O_2412,N_19810,N_18225);
and UO_2413 (O_2413,N_18539,N_19721);
or UO_2414 (O_2414,N_19482,N_18815);
nand UO_2415 (O_2415,N_19628,N_18700);
nand UO_2416 (O_2416,N_19633,N_18509);
nor UO_2417 (O_2417,N_19133,N_18165);
nor UO_2418 (O_2418,N_18038,N_18703);
nor UO_2419 (O_2419,N_19036,N_18422);
nand UO_2420 (O_2420,N_19259,N_19421);
or UO_2421 (O_2421,N_18992,N_18113);
or UO_2422 (O_2422,N_18429,N_19846);
nand UO_2423 (O_2423,N_18221,N_18368);
nor UO_2424 (O_2424,N_19342,N_19879);
nand UO_2425 (O_2425,N_19020,N_19530);
nand UO_2426 (O_2426,N_19756,N_19423);
nor UO_2427 (O_2427,N_19036,N_19105);
nand UO_2428 (O_2428,N_19448,N_18930);
or UO_2429 (O_2429,N_19331,N_19636);
xnor UO_2430 (O_2430,N_18344,N_19184);
nor UO_2431 (O_2431,N_18834,N_18988);
nor UO_2432 (O_2432,N_19347,N_18580);
xor UO_2433 (O_2433,N_18181,N_18361);
and UO_2434 (O_2434,N_19596,N_19959);
and UO_2435 (O_2435,N_19051,N_18114);
nand UO_2436 (O_2436,N_18935,N_18289);
nor UO_2437 (O_2437,N_19584,N_19860);
nor UO_2438 (O_2438,N_19534,N_19099);
nand UO_2439 (O_2439,N_19286,N_19737);
nand UO_2440 (O_2440,N_19511,N_18458);
or UO_2441 (O_2441,N_18109,N_19778);
or UO_2442 (O_2442,N_18579,N_18633);
xor UO_2443 (O_2443,N_18859,N_18875);
xor UO_2444 (O_2444,N_18203,N_18220);
or UO_2445 (O_2445,N_19765,N_18812);
nand UO_2446 (O_2446,N_19845,N_18511);
nand UO_2447 (O_2447,N_18049,N_19221);
nor UO_2448 (O_2448,N_18269,N_18270);
and UO_2449 (O_2449,N_19894,N_19549);
and UO_2450 (O_2450,N_18624,N_18168);
xor UO_2451 (O_2451,N_18966,N_19421);
nand UO_2452 (O_2452,N_18370,N_19017);
or UO_2453 (O_2453,N_19109,N_18379);
nand UO_2454 (O_2454,N_18372,N_19339);
or UO_2455 (O_2455,N_18277,N_18057);
nand UO_2456 (O_2456,N_19650,N_19038);
xor UO_2457 (O_2457,N_19476,N_19355);
and UO_2458 (O_2458,N_19725,N_18044);
or UO_2459 (O_2459,N_19096,N_18427);
nor UO_2460 (O_2460,N_19322,N_18980);
or UO_2461 (O_2461,N_19277,N_19701);
or UO_2462 (O_2462,N_18110,N_18016);
nand UO_2463 (O_2463,N_18678,N_19331);
nor UO_2464 (O_2464,N_18303,N_18861);
nor UO_2465 (O_2465,N_19717,N_18987);
nor UO_2466 (O_2466,N_19798,N_18566);
or UO_2467 (O_2467,N_19663,N_18232);
xor UO_2468 (O_2468,N_19255,N_18348);
and UO_2469 (O_2469,N_19939,N_19150);
and UO_2470 (O_2470,N_18671,N_19655);
nand UO_2471 (O_2471,N_18246,N_18442);
xor UO_2472 (O_2472,N_19330,N_19307);
nand UO_2473 (O_2473,N_18743,N_18555);
or UO_2474 (O_2474,N_18496,N_19192);
nor UO_2475 (O_2475,N_19711,N_19323);
xnor UO_2476 (O_2476,N_19541,N_19547);
nand UO_2477 (O_2477,N_18332,N_19599);
nand UO_2478 (O_2478,N_19705,N_19387);
nand UO_2479 (O_2479,N_19328,N_18935);
xnor UO_2480 (O_2480,N_18841,N_19684);
or UO_2481 (O_2481,N_18377,N_19368);
or UO_2482 (O_2482,N_18968,N_19193);
xnor UO_2483 (O_2483,N_18807,N_18637);
and UO_2484 (O_2484,N_18352,N_19604);
nand UO_2485 (O_2485,N_18143,N_18917);
nand UO_2486 (O_2486,N_18484,N_18020);
and UO_2487 (O_2487,N_19555,N_18236);
nand UO_2488 (O_2488,N_19421,N_19584);
nand UO_2489 (O_2489,N_18564,N_18116);
and UO_2490 (O_2490,N_18976,N_19538);
and UO_2491 (O_2491,N_19723,N_18112);
nor UO_2492 (O_2492,N_18521,N_19093);
xnor UO_2493 (O_2493,N_19965,N_18556);
nor UO_2494 (O_2494,N_18903,N_18845);
nor UO_2495 (O_2495,N_19185,N_19085);
nor UO_2496 (O_2496,N_19317,N_19217);
xor UO_2497 (O_2497,N_19092,N_18575);
and UO_2498 (O_2498,N_19404,N_19503);
and UO_2499 (O_2499,N_18932,N_18513);
endmodule