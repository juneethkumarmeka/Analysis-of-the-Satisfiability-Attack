module basic_750_5000_1000_10_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_620,In_399);
or U1 (N_1,In_400,In_632);
nor U2 (N_2,In_681,In_116);
or U3 (N_3,In_146,In_120);
nor U4 (N_4,In_520,In_32);
or U5 (N_5,In_584,In_442);
nor U6 (N_6,In_179,In_588);
nand U7 (N_7,In_30,In_445);
nand U8 (N_8,In_69,In_614);
or U9 (N_9,In_309,In_211);
nand U10 (N_10,In_176,In_200);
nand U11 (N_11,In_271,In_175);
or U12 (N_12,In_367,In_21);
or U13 (N_13,In_297,In_745);
nor U14 (N_14,In_368,In_523);
nand U15 (N_15,In_487,In_645);
nand U16 (N_16,In_42,In_383);
nor U17 (N_17,In_391,In_37);
nand U18 (N_18,In_464,In_561);
nand U19 (N_19,In_371,In_551);
nor U20 (N_20,In_448,In_119);
nand U21 (N_21,In_98,In_246);
nor U22 (N_22,In_337,In_601);
and U23 (N_23,In_52,In_743);
or U24 (N_24,In_629,In_259);
nand U25 (N_25,In_344,In_83);
and U26 (N_26,In_335,In_555);
nand U27 (N_27,In_392,In_115);
xnor U28 (N_28,In_612,In_708);
nand U29 (N_29,In_690,In_247);
nor U30 (N_30,In_231,In_53);
or U31 (N_31,In_587,In_536);
and U32 (N_32,In_689,In_10);
or U33 (N_33,In_703,In_502);
nand U34 (N_34,In_133,In_623);
nand U35 (N_35,In_333,In_222);
and U36 (N_36,In_132,In_78);
or U37 (N_37,In_552,In_699);
nand U38 (N_38,In_171,In_504);
or U39 (N_39,In_67,In_44);
or U40 (N_40,In_479,In_16);
nand U41 (N_41,In_204,In_616);
and U42 (N_42,In_99,In_294);
and U43 (N_43,In_62,In_596);
nand U44 (N_44,In_111,In_118);
nand U45 (N_45,In_2,In_109);
and U46 (N_46,In_291,In_156);
or U47 (N_47,In_624,In_726);
or U48 (N_48,In_0,In_286);
or U49 (N_49,In_379,In_595);
or U50 (N_50,In_355,In_700);
and U51 (N_51,In_470,In_518);
nor U52 (N_52,In_573,In_480);
nor U53 (N_53,In_427,In_729);
and U54 (N_54,In_388,In_138);
xor U55 (N_55,In_321,In_610);
nand U56 (N_56,In_134,In_112);
and U57 (N_57,In_477,In_419);
or U58 (N_58,In_190,In_542);
nand U59 (N_59,In_178,In_695);
nand U60 (N_60,In_26,In_356);
nor U61 (N_61,In_611,In_72);
nor U62 (N_62,In_251,In_346);
and U63 (N_63,In_507,In_4);
nand U64 (N_64,In_710,In_339);
nand U65 (N_65,In_205,In_409);
nand U66 (N_66,In_221,In_385);
nand U67 (N_67,In_510,In_27);
nor U68 (N_68,In_415,In_455);
nor U69 (N_69,In_151,In_663);
and U70 (N_70,In_563,In_357);
nor U71 (N_71,In_272,In_397);
and U72 (N_72,In_471,In_217);
and U73 (N_73,In_287,In_433);
nor U74 (N_74,In_631,In_13);
or U75 (N_75,In_342,In_64);
nand U76 (N_76,In_264,In_48);
and U77 (N_77,In_312,In_240);
nor U78 (N_78,In_3,In_716);
or U79 (N_79,In_589,In_336);
and U80 (N_80,In_664,In_489);
and U81 (N_81,In_239,In_674);
and U82 (N_82,In_500,In_150);
nor U83 (N_83,In_575,In_401);
or U84 (N_84,In_642,In_43);
nand U85 (N_85,In_332,In_659);
and U86 (N_86,In_672,In_11);
nand U87 (N_87,In_39,In_665);
xor U88 (N_88,In_256,In_328);
nor U89 (N_89,In_582,In_57);
nand U90 (N_90,In_84,In_526);
or U91 (N_91,In_378,In_538);
nand U92 (N_92,In_432,In_640);
nand U93 (N_93,In_124,In_651);
nand U94 (N_94,In_34,In_511);
nor U95 (N_95,In_531,In_698);
or U96 (N_96,In_412,In_714);
nand U97 (N_97,In_130,In_254);
and U98 (N_98,In_330,In_723);
and U99 (N_99,In_566,In_186);
and U100 (N_100,In_19,In_216);
and U101 (N_101,In_313,In_686);
or U102 (N_102,In_506,In_576);
and U103 (N_103,In_281,In_476);
and U104 (N_104,In_436,In_189);
nor U105 (N_105,In_474,In_530);
nor U106 (N_106,In_375,In_425);
nand U107 (N_107,In_349,In_565);
xor U108 (N_108,In_300,In_331);
nor U109 (N_109,In_418,In_381);
nor U110 (N_110,In_396,In_517);
nand U111 (N_111,In_22,In_524);
or U112 (N_112,In_707,In_647);
or U113 (N_113,In_194,In_282);
or U114 (N_114,In_258,In_157);
nand U115 (N_115,In_302,In_586);
and U116 (N_116,In_634,In_577);
and U117 (N_117,In_75,In_492);
nand U118 (N_118,In_145,In_718);
and U119 (N_119,In_261,In_311);
nand U120 (N_120,In_546,In_456);
or U121 (N_121,In_210,In_416);
and U122 (N_122,In_354,In_613);
and U123 (N_123,In_110,In_428);
nor U124 (N_124,In_318,In_508);
and U125 (N_125,In_528,In_557);
nor U126 (N_126,In_225,In_424);
nor U127 (N_127,In_56,In_715);
and U128 (N_128,In_503,In_574);
and U129 (N_129,In_376,In_618);
or U130 (N_130,In_420,In_550);
and U131 (N_131,In_564,In_267);
nand U132 (N_132,In_82,In_403);
and U133 (N_133,In_314,In_630);
and U134 (N_134,In_541,In_276);
or U135 (N_135,In_114,In_701);
or U136 (N_136,In_547,In_209);
nor U137 (N_137,In_235,In_724);
and U138 (N_138,In_369,In_705);
nand U139 (N_139,In_158,In_148);
nor U140 (N_140,In_554,In_91);
and U141 (N_141,In_320,In_633);
or U142 (N_142,In_439,In_55);
nor U143 (N_143,In_285,In_627);
nor U144 (N_144,In_741,In_603);
and U145 (N_145,In_213,In_232);
or U146 (N_146,In_41,In_636);
or U147 (N_147,In_556,In_545);
nand U148 (N_148,In_70,In_174);
and U149 (N_149,In_182,In_660);
or U150 (N_150,In_458,In_126);
nor U151 (N_151,In_599,In_341);
nand U152 (N_152,In_402,In_713);
or U153 (N_153,In_417,In_527);
and U154 (N_154,In_410,In_180);
nand U155 (N_155,In_35,In_384);
or U156 (N_156,In_277,In_571);
and U157 (N_157,In_14,In_80);
nor U158 (N_158,In_693,In_165);
or U159 (N_159,In_467,In_496);
and U160 (N_160,In_387,In_366);
and U161 (N_161,In_350,In_658);
nor U162 (N_162,In_275,In_441);
nor U163 (N_163,In_63,In_47);
or U164 (N_164,In_308,In_404);
or U165 (N_165,In_516,In_656);
nand U166 (N_166,In_65,In_137);
and U167 (N_167,In_602,In_533);
nand U168 (N_168,In_485,In_499);
or U169 (N_169,In_461,In_365);
nand U170 (N_170,In_229,In_74);
nand U171 (N_171,In_242,In_495);
nand U172 (N_172,In_394,In_347);
nor U173 (N_173,In_568,In_236);
nand U174 (N_174,In_559,In_592);
and U175 (N_175,In_682,In_649);
and U176 (N_176,In_326,In_666);
and U177 (N_177,In_208,In_426);
or U178 (N_178,In_299,In_289);
or U179 (N_179,In_744,In_278);
and U180 (N_180,In_621,In_459);
nand U181 (N_181,In_730,In_478);
or U182 (N_182,In_735,In_683);
or U183 (N_183,In_23,In_702);
and U184 (N_184,In_548,In_40);
or U185 (N_185,In_226,In_188);
and U186 (N_186,In_58,In_214);
or U187 (N_187,In_494,In_722);
nand U188 (N_188,In_532,In_155);
nand U189 (N_189,In_628,In_351);
nor U190 (N_190,In_49,In_28);
nor U191 (N_191,In_739,In_319);
and U192 (N_192,In_173,In_431);
and U193 (N_193,In_227,In_212);
and U194 (N_194,In_583,In_626);
and U195 (N_195,In_688,In_102);
nand U196 (N_196,In_484,In_562);
nand U197 (N_197,In_680,In_590);
or U198 (N_198,In_169,In_668);
nand U199 (N_199,In_315,In_373);
and U200 (N_200,In_260,In_619);
and U201 (N_201,In_594,In_296);
nor U202 (N_202,In_20,In_421);
and U203 (N_203,In_73,In_482);
nand U204 (N_204,In_199,In_706);
and U205 (N_205,In_121,In_529);
and U206 (N_206,In_444,In_125);
nand U207 (N_207,In_206,In_184);
nand U208 (N_208,In_87,In_717);
nand U209 (N_209,In_544,In_446);
and U210 (N_210,In_244,In_678);
nor U211 (N_211,In_360,In_152);
and U212 (N_212,In_304,In_234);
nand U213 (N_213,In_105,In_740);
and U214 (N_214,In_60,In_560);
nand U215 (N_215,In_273,In_488);
or U216 (N_216,In_68,In_736);
nor U217 (N_217,In_661,In_59);
and U218 (N_218,In_465,In_293);
and U219 (N_219,In_719,In_238);
nand U220 (N_220,In_593,In_66);
nor U221 (N_221,In_18,In_475);
nor U222 (N_222,In_306,In_692);
nand U223 (N_223,In_728,In_606);
nor U224 (N_224,In_737,In_650);
or U225 (N_225,In_389,In_746);
or U226 (N_226,In_472,In_501);
and U227 (N_227,In_525,In_274);
and U228 (N_228,In_691,In_248);
or U229 (N_229,In_162,In_71);
nand U230 (N_230,In_654,In_377);
and U231 (N_231,In_100,In_245);
nand U232 (N_232,In_519,In_514);
xor U233 (N_233,In_197,In_352);
or U234 (N_234,In_581,In_423);
nand U235 (N_235,In_372,In_51);
nor U236 (N_236,In_295,In_604);
nor U237 (N_237,In_440,In_644);
and U238 (N_238,In_280,In_748);
and U239 (N_239,In_522,In_405);
or U240 (N_240,In_535,In_742);
or U241 (N_241,In_580,In_453);
nor U242 (N_242,In_224,In_370);
or U243 (N_243,In_615,In_268);
and U244 (N_244,In_639,In_725);
nor U245 (N_245,In_657,In_81);
or U246 (N_246,In_608,In_288);
nand U247 (N_247,In_648,In_720);
and U248 (N_248,In_407,In_679);
and U249 (N_249,In_727,In_414);
nor U250 (N_250,In_153,In_600);
or U251 (N_251,In_325,In_24);
nor U252 (N_252,In_122,In_343);
nand U253 (N_253,In_164,In_185);
nor U254 (N_254,In_662,In_486);
nor U255 (N_255,In_358,In_90);
nand U256 (N_256,In_572,In_435);
nand U257 (N_257,In_127,In_643);
nand U258 (N_258,In_107,In_452);
or U259 (N_259,In_187,In_215);
nor U260 (N_260,In_732,In_29);
nand U261 (N_261,In_512,In_298);
nand U262 (N_262,In_135,In_443);
xor U263 (N_263,In_144,In_270);
or U264 (N_264,In_709,In_143);
or U265 (N_265,In_635,In_374);
and U266 (N_266,In_45,In_540);
nor U267 (N_267,In_36,In_46);
nand U268 (N_268,In_31,In_327);
nor U269 (N_269,In_266,In_466);
and U270 (N_270,In_323,In_322);
nand U271 (N_271,In_283,In_223);
or U272 (N_272,In_451,In_413);
nand U273 (N_273,In_95,In_93);
nor U274 (N_274,In_578,In_198);
or U275 (N_275,In_104,In_290);
nor U276 (N_276,In_734,In_422);
nor U277 (N_277,In_509,In_625);
or U278 (N_278,In_203,In_671);
nand U279 (N_279,In_361,In_33);
nor U280 (N_280,In_228,In_738);
nand U281 (N_281,In_303,In_353);
nand U282 (N_282,In_136,In_468);
nor U283 (N_283,In_598,In_348);
and U284 (N_284,In_233,In_123);
or U285 (N_285,In_25,In_670);
nor U286 (N_286,In_605,In_345);
or U287 (N_287,In_617,In_38);
nand U288 (N_288,In_324,In_310);
or U289 (N_289,In_597,In_570);
nand U290 (N_290,In_430,In_17);
or U291 (N_291,In_159,In_638);
nor U292 (N_292,In_237,In_667);
nor U293 (N_293,In_641,In_493);
nand U294 (N_294,In_301,In_129);
nand U295 (N_295,In_307,In_305);
nand U296 (N_296,In_89,In_12);
nand U297 (N_297,In_257,In_106);
nor U298 (N_298,In_97,In_147);
nor U299 (N_299,In_195,In_646);
or U300 (N_300,In_279,In_149);
or U301 (N_301,In_607,In_449);
nand U302 (N_302,In_386,In_408);
nor U303 (N_303,In_398,In_481);
nand U304 (N_304,In_50,In_543);
or U305 (N_305,In_553,In_637);
nand U306 (N_306,In_167,In_96);
nor U307 (N_307,In_491,In_177);
nor U308 (N_308,In_202,In_362);
nor U309 (N_309,In_549,In_539);
xnor U310 (N_310,In_673,In_498);
nand U311 (N_311,In_463,In_515);
nor U312 (N_312,In_250,In_61);
nand U313 (N_313,In_382,In_54);
or U314 (N_314,In_450,In_207);
or U315 (N_315,In_7,In_141);
or U316 (N_316,In_696,In_163);
nor U317 (N_317,In_329,In_569);
and U318 (N_318,In_128,In_334);
and U319 (N_319,In_558,In_168);
nor U320 (N_320,In_469,In_166);
nor U321 (N_321,In_196,In_731);
and U322 (N_322,In_139,In_269);
and U323 (N_323,In_170,In_521);
nor U324 (N_324,In_395,In_181);
nand U325 (N_325,In_76,In_359);
nor U326 (N_326,In_6,In_241);
nand U327 (N_327,In_317,In_192);
nor U328 (N_328,In_191,In_8);
nor U329 (N_329,In_117,In_460);
and U330 (N_330,In_103,In_406);
nand U331 (N_331,In_101,In_437);
or U332 (N_332,In_434,In_497);
or U333 (N_333,In_140,In_652);
and U334 (N_334,In_363,In_622);
nor U335 (N_335,In_220,In_537);
nor U336 (N_336,In_201,In_160);
nor U337 (N_337,In_711,In_534);
or U338 (N_338,In_88,In_142);
or U339 (N_339,In_108,In_697);
or U340 (N_340,In_438,In_687);
nand U341 (N_341,In_15,In_94);
nand U342 (N_342,In_249,In_77);
or U343 (N_343,In_721,In_655);
or U344 (N_344,In_364,In_712);
nor U345 (N_345,In_505,In_243);
nor U346 (N_346,In_747,In_172);
nor U347 (N_347,In_653,In_230);
or U348 (N_348,In_684,In_9);
and U349 (N_349,In_457,In_393);
and U350 (N_350,In_113,In_131);
nor U351 (N_351,In_609,In_447);
and U352 (N_352,In_579,In_677);
nand U353 (N_353,In_5,In_316);
or U354 (N_354,In_340,In_292);
nand U355 (N_355,In_462,In_429);
nand U356 (N_356,In_704,In_483);
nor U357 (N_357,In_490,In_473);
or U358 (N_358,In_86,In_685);
or U359 (N_359,In_161,In_585);
nand U360 (N_360,In_380,In_154);
and U361 (N_361,In_255,In_253);
nand U362 (N_362,In_454,In_262);
nor U363 (N_363,In_749,In_252);
or U364 (N_364,In_675,In_219);
nand U365 (N_365,In_733,In_1);
nand U366 (N_366,In_218,In_338);
and U367 (N_367,In_513,In_92);
nor U368 (N_368,In_85,In_265);
or U369 (N_369,In_694,In_390);
or U370 (N_370,In_183,In_567);
or U371 (N_371,In_79,In_591);
nand U372 (N_372,In_263,In_411);
or U373 (N_373,In_193,In_669);
or U374 (N_374,In_284,In_676);
nand U375 (N_375,In_671,In_653);
nor U376 (N_376,In_535,In_685);
nand U377 (N_377,In_172,In_729);
nor U378 (N_378,In_503,In_193);
and U379 (N_379,In_182,In_493);
or U380 (N_380,In_691,In_130);
or U381 (N_381,In_507,In_583);
nand U382 (N_382,In_151,In_56);
nor U383 (N_383,In_518,In_91);
nand U384 (N_384,In_85,In_526);
nor U385 (N_385,In_448,In_732);
nor U386 (N_386,In_738,In_400);
nor U387 (N_387,In_279,In_376);
nand U388 (N_388,In_669,In_662);
nor U389 (N_389,In_441,In_231);
nor U390 (N_390,In_450,In_560);
or U391 (N_391,In_341,In_188);
nand U392 (N_392,In_391,In_256);
or U393 (N_393,In_453,In_36);
nor U394 (N_394,In_20,In_556);
nand U395 (N_395,In_320,In_65);
nor U396 (N_396,In_631,In_269);
nand U397 (N_397,In_404,In_385);
nor U398 (N_398,In_326,In_463);
nor U399 (N_399,In_567,In_395);
or U400 (N_400,In_376,In_268);
xnor U401 (N_401,In_373,In_509);
nor U402 (N_402,In_523,In_464);
nor U403 (N_403,In_308,In_286);
or U404 (N_404,In_504,In_226);
nor U405 (N_405,In_408,In_59);
nor U406 (N_406,In_434,In_441);
xnor U407 (N_407,In_363,In_159);
nand U408 (N_408,In_15,In_160);
and U409 (N_409,In_549,In_598);
and U410 (N_410,In_127,In_505);
and U411 (N_411,In_141,In_346);
or U412 (N_412,In_739,In_232);
nor U413 (N_413,In_450,In_203);
or U414 (N_414,In_645,In_38);
and U415 (N_415,In_572,In_674);
xor U416 (N_416,In_171,In_274);
or U417 (N_417,In_681,In_401);
and U418 (N_418,In_531,In_386);
and U419 (N_419,In_255,In_500);
and U420 (N_420,In_394,In_564);
and U421 (N_421,In_404,In_118);
nor U422 (N_422,In_645,In_202);
or U423 (N_423,In_515,In_206);
or U424 (N_424,In_528,In_197);
nor U425 (N_425,In_534,In_540);
nand U426 (N_426,In_719,In_714);
and U427 (N_427,In_363,In_131);
or U428 (N_428,In_330,In_77);
and U429 (N_429,In_708,In_600);
nand U430 (N_430,In_114,In_154);
or U431 (N_431,In_280,In_715);
nor U432 (N_432,In_460,In_178);
and U433 (N_433,In_440,In_62);
nand U434 (N_434,In_166,In_229);
and U435 (N_435,In_298,In_357);
or U436 (N_436,In_102,In_74);
nor U437 (N_437,In_277,In_291);
xnor U438 (N_438,In_85,In_1);
and U439 (N_439,In_316,In_191);
or U440 (N_440,In_740,In_301);
nor U441 (N_441,In_81,In_214);
nor U442 (N_442,In_709,In_678);
nand U443 (N_443,In_399,In_648);
nor U444 (N_444,In_279,In_232);
nand U445 (N_445,In_353,In_130);
and U446 (N_446,In_30,In_102);
nand U447 (N_447,In_367,In_84);
nor U448 (N_448,In_139,In_110);
nor U449 (N_449,In_373,In_736);
xor U450 (N_450,In_718,In_309);
and U451 (N_451,In_127,In_556);
or U452 (N_452,In_144,In_535);
nor U453 (N_453,In_302,In_287);
and U454 (N_454,In_249,In_661);
nor U455 (N_455,In_529,In_431);
nor U456 (N_456,In_676,In_331);
nand U457 (N_457,In_359,In_610);
nand U458 (N_458,In_456,In_30);
xor U459 (N_459,In_207,In_543);
and U460 (N_460,In_589,In_135);
nand U461 (N_461,In_313,In_463);
or U462 (N_462,In_260,In_634);
nor U463 (N_463,In_353,In_380);
or U464 (N_464,In_139,In_128);
and U465 (N_465,In_199,In_521);
and U466 (N_466,In_732,In_345);
nor U467 (N_467,In_127,In_500);
and U468 (N_468,In_667,In_77);
or U469 (N_469,In_649,In_177);
nand U470 (N_470,In_493,In_656);
or U471 (N_471,In_107,In_346);
nand U472 (N_472,In_356,In_588);
nand U473 (N_473,In_289,In_81);
nor U474 (N_474,In_1,In_213);
and U475 (N_475,In_561,In_298);
or U476 (N_476,In_253,In_224);
or U477 (N_477,In_172,In_519);
and U478 (N_478,In_425,In_467);
nor U479 (N_479,In_118,In_123);
or U480 (N_480,In_132,In_134);
or U481 (N_481,In_265,In_214);
xor U482 (N_482,In_657,In_380);
and U483 (N_483,In_257,In_391);
and U484 (N_484,In_224,In_305);
nor U485 (N_485,In_138,In_586);
or U486 (N_486,In_303,In_31);
nand U487 (N_487,In_86,In_558);
nor U488 (N_488,In_741,In_460);
or U489 (N_489,In_55,In_289);
nand U490 (N_490,In_660,In_366);
or U491 (N_491,In_120,In_25);
and U492 (N_492,In_703,In_283);
and U493 (N_493,In_106,In_673);
or U494 (N_494,In_217,In_194);
and U495 (N_495,In_449,In_495);
nor U496 (N_496,In_466,In_25);
and U497 (N_497,In_212,In_607);
or U498 (N_498,In_481,In_8);
nor U499 (N_499,In_684,In_545);
and U500 (N_500,N_17,N_202);
nand U501 (N_501,N_372,N_322);
and U502 (N_502,N_146,N_136);
nor U503 (N_503,N_487,N_426);
nor U504 (N_504,N_294,N_227);
and U505 (N_505,N_381,N_199);
nand U506 (N_506,N_210,N_88);
nand U507 (N_507,N_339,N_392);
nand U508 (N_508,N_6,N_296);
or U509 (N_509,N_469,N_463);
nand U510 (N_510,N_348,N_117);
nand U511 (N_511,N_442,N_72);
or U512 (N_512,N_404,N_456);
nand U513 (N_513,N_179,N_100);
xnor U514 (N_514,N_47,N_375);
xnor U515 (N_515,N_422,N_63);
and U516 (N_516,N_32,N_309);
nor U517 (N_517,N_174,N_145);
nor U518 (N_518,N_219,N_259);
nor U519 (N_519,N_396,N_376);
and U520 (N_520,N_112,N_14);
and U521 (N_521,N_495,N_25);
xnor U522 (N_522,N_19,N_450);
or U523 (N_523,N_382,N_29);
nand U524 (N_524,N_153,N_474);
nand U525 (N_525,N_143,N_308);
nor U526 (N_526,N_85,N_147);
and U527 (N_527,N_111,N_81);
and U528 (N_528,N_283,N_353);
and U529 (N_529,N_346,N_340);
and U530 (N_530,N_104,N_21);
nand U531 (N_531,N_78,N_189);
or U532 (N_532,N_443,N_394);
or U533 (N_533,N_238,N_180);
and U534 (N_534,N_278,N_126);
nor U535 (N_535,N_395,N_218);
or U536 (N_536,N_53,N_192);
nand U537 (N_537,N_31,N_256);
or U538 (N_538,N_436,N_142);
or U539 (N_539,N_137,N_217);
and U540 (N_540,N_282,N_234);
nand U541 (N_541,N_452,N_9);
nand U542 (N_542,N_352,N_252);
nor U543 (N_543,N_141,N_359);
and U544 (N_544,N_447,N_203);
nand U545 (N_545,N_285,N_48);
nand U546 (N_546,N_247,N_99);
and U547 (N_547,N_35,N_267);
and U548 (N_548,N_454,N_11);
xnor U549 (N_549,N_451,N_7);
nor U550 (N_550,N_354,N_249);
and U551 (N_551,N_39,N_480);
or U552 (N_552,N_440,N_304);
nor U553 (N_553,N_57,N_50);
nor U554 (N_554,N_338,N_60);
nand U555 (N_555,N_277,N_321);
nand U556 (N_556,N_272,N_411);
and U557 (N_557,N_260,N_41);
nand U558 (N_558,N_151,N_478);
nand U559 (N_559,N_434,N_211);
nor U560 (N_560,N_163,N_423);
nor U561 (N_561,N_242,N_369);
nor U562 (N_562,N_318,N_453);
and U563 (N_563,N_313,N_264);
or U564 (N_564,N_403,N_168);
or U565 (N_565,N_162,N_20);
or U566 (N_566,N_129,N_86);
and U567 (N_567,N_213,N_248);
and U568 (N_568,N_62,N_430);
and U569 (N_569,N_470,N_262);
or U570 (N_570,N_108,N_171);
and U571 (N_571,N_459,N_297);
nor U572 (N_572,N_386,N_55);
or U573 (N_573,N_204,N_87);
nand U574 (N_574,N_188,N_43);
nor U575 (N_575,N_84,N_82);
nand U576 (N_576,N_274,N_131);
and U577 (N_577,N_127,N_388);
nand U578 (N_578,N_161,N_128);
nand U579 (N_579,N_377,N_184);
nand U580 (N_580,N_327,N_45);
nand U581 (N_581,N_428,N_245);
and U582 (N_582,N_221,N_330);
and U583 (N_583,N_114,N_150);
nor U584 (N_584,N_389,N_152);
xor U585 (N_585,N_149,N_130);
or U586 (N_586,N_1,N_26);
nand U587 (N_587,N_97,N_408);
nor U588 (N_588,N_457,N_483);
and U589 (N_589,N_125,N_374);
and U590 (N_590,N_244,N_455);
xnor U591 (N_591,N_183,N_44);
nand U592 (N_592,N_79,N_134);
nor U593 (N_593,N_276,N_431);
nand U594 (N_594,N_64,N_305);
nor U595 (N_595,N_226,N_177);
xor U596 (N_596,N_186,N_323);
nor U597 (N_597,N_89,N_121);
nor U598 (N_598,N_233,N_361);
nand U599 (N_599,N_257,N_448);
nand U600 (N_600,N_75,N_413);
xor U601 (N_601,N_397,N_194);
nand U602 (N_602,N_466,N_176);
and U603 (N_603,N_228,N_132);
nor U604 (N_604,N_206,N_419);
nand U605 (N_605,N_412,N_358);
xnor U606 (N_606,N_182,N_3);
or U607 (N_607,N_387,N_239);
and U608 (N_608,N_328,N_356);
nand U609 (N_609,N_401,N_498);
nand U610 (N_610,N_109,N_307);
and U611 (N_611,N_298,N_342);
and U612 (N_612,N_406,N_52);
or U613 (N_613,N_123,N_200);
nand U614 (N_614,N_326,N_230);
nand U615 (N_615,N_421,N_461);
nor U616 (N_616,N_98,N_236);
or U617 (N_617,N_347,N_435);
xor U618 (N_618,N_493,N_336);
or U619 (N_619,N_362,N_140);
or U620 (N_620,N_301,N_254);
and U621 (N_621,N_488,N_207);
and U622 (N_622,N_280,N_289);
and U623 (N_623,N_222,N_22);
nor U624 (N_624,N_178,N_16);
or U625 (N_625,N_420,N_159);
nor U626 (N_626,N_391,N_209);
or U627 (N_627,N_23,N_148);
nor U628 (N_628,N_497,N_485);
and U629 (N_629,N_5,N_324);
and U630 (N_630,N_165,N_351);
xor U631 (N_631,N_445,N_317);
and U632 (N_632,N_92,N_360);
nand U633 (N_633,N_311,N_292);
nand U634 (N_634,N_122,N_441);
nand U635 (N_635,N_286,N_429);
nand U636 (N_636,N_0,N_74);
xor U637 (N_637,N_172,N_258);
nor U638 (N_638,N_287,N_281);
nor U639 (N_639,N_494,N_49);
nand U640 (N_640,N_490,N_385);
nor U641 (N_641,N_458,N_61);
and U642 (N_642,N_365,N_471);
or U643 (N_643,N_415,N_270);
nor U644 (N_644,N_341,N_299);
nor U645 (N_645,N_93,N_373);
or U646 (N_646,N_95,N_366);
nor U647 (N_647,N_349,N_246);
nor U648 (N_648,N_473,N_118);
nand U649 (N_649,N_193,N_479);
nor U650 (N_650,N_157,N_329);
and U651 (N_651,N_59,N_208);
nor U652 (N_652,N_390,N_198);
nor U653 (N_653,N_486,N_417);
nor U654 (N_654,N_144,N_400);
nand U655 (N_655,N_187,N_215);
or U656 (N_656,N_379,N_170);
or U657 (N_657,N_51,N_164);
nand U658 (N_658,N_224,N_83);
nand U659 (N_659,N_36,N_139);
or U660 (N_660,N_472,N_2);
and U661 (N_661,N_433,N_476);
nand U662 (N_662,N_34,N_438);
or U663 (N_663,N_464,N_425);
and U664 (N_664,N_12,N_462);
or U665 (N_665,N_70,N_124);
nand U666 (N_666,N_195,N_10);
or U667 (N_667,N_237,N_439);
and U668 (N_668,N_467,N_316);
nand U669 (N_669,N_197,N_335);
nor U670 (N_670,N_27,N_231);
or U671 (N_671,N_266,N_71);
or U672 (N_672,N_155,N_302);
and U673 (N_673,N_491,N_409);
or U674 (N_674,N_255,N_371);
nand U675 (N_675,N_468,N_378);
and U676 (N_676,N_80,N_268);
nand U677 (N_677,N_235,N_333);
xnor U678 (N_678,N_398,N_119);
nor U679 (N_679,N_477,N_24);
nor U680 (N_680,N_28,N_69);
nor U681 (N_681,N_320,N_407);
xor U682 (N_682,N_444,N_295);
and U683 (N_683,N_229,N_68);
nand U684 (N_684,N_135,N_275);
or U685 (N_685,N_482,N_261);
nor U686 (N_686,N_38,N_363);
nor U687 (N_687,N_185,N_383);
nand U688 (N_688,N_263,N_300);
nor U689 (N_689,N_113,N_418);
nor U690 (N_690,N_288,N_279);
nor U691 (N_691,N_67,N_331);
nor U692 (N_692,N_103,N_223);
nand U693 (N_693,N_460,N_465);
or U694 (N_694,N_18,N_427);
and U695 (N_695,N_56,N_332);
or U696 (N_696,N_30,N_399);
or U697 (N_697,N_115,N_156);
nor U698 (N_698,N_107,N_66);
and U699 (N_699,N_205,N_496);
nand U700 (N_700,N_303,N_293);
or U701 (N_701,N_290,N_33);
or U702 (N_702,N_265,N_492);
and U703 (N_703,N_484,N_350);
and U704 (N_704,N_344,N_232);
nor U705 (N_705,N_173,N_76);
or U706 (N_706,N_91,N_273);
or U707 (N_707,N_158,N_481);
nor U708 (N_708,N_410,N_169);
and U709 (N_709,N_15,N_437);
or U710 (N_710,N_345,N_120);
nand U711 (N_711,N_4,N_343);
nand U712 (N_712,N_46,N_116);
nor U713 (N_713,N_106,N_319);
nand U714 (N_714,N_402,N_37);
nand U715 (N_715,N_73,N_380);
or U716 (N_716,N_40,N_414);
nor U717 (N_717,N_475,N_310);
or U718 (N_718,N_196,N_271);
or U719 (N_719,N_384,N_240);
and U720 (N_720,N_489,N_101);
and U721 (N_721,N_102,N_96);
nand U722 (N_722,N_243,N_337);
or U723 (N_723,N_191,N_212);
or U724 (N_724,N_190,N_133);
nor U725 (N_725,N_367,N_214);
nand U726 (N_726,N_253,N_94);
nand U727 (N_727,N_370,N_250);
nand U728 (N_728,N_241,N_446);
nor U729 (N_729,N_216,N_105);
or U730 (N_730,N_499,N_225);
and U731 (N_731,N_90,N_8);
or U732 (N_732,N_54,N_167);
nand U733 (N_733,N_269,N_325);
nor U734 (N_734,N_77,N_355);
and U735 (N_735,N_284,N_13);
nor U736 (N_736,N_160,N_181);
nand U737 (N_737,N_315,N_291);
nor U738 (N_738,N_312,N_201);
or U739 (N_739,N_65,N_334);
nor U740 (N_740,N_424,N_175);
or U741 (N_741,N_357,N_364);
nor U742 (N_742,N_251,N_138);
or U743 (N_743,N_416,N_166);
nor U744 (N_744,N_154,N_58);
nor U745 (N_745,N_306,N_432);
or U746 (N_746,N_220,N_110);
or U747 (N_747,N_405,N_314);
or U748 (N_748,N_42,N_393);
and U749 (N_749,N_449,N_368);
nor U750 (N_750,N_264,N_467);
nor U751 (N_751,N_148,N_201);
nor U752 (N_752,N_206,N_193);
nor U753 (N_753,N_272,N_135);
nand U754 (N_754,N_304,N_108);
or U755 (N_755,N_388,N_375);
nand U756 (N_756,N_129,N_44);
and U757 (N_757,N_48,N_222);
or U758 (N_758,N_56,N_494);
xor U759 (N_759,N_147,N_101);
and U760 (N_760,N_489,N_347);
or U761 (N_761,N_391,N_130);
nand U762 (N_762,N_264,N_293);
and U763 (N_763,N_227,N_85);
or U764 (N_764,N_233,N_411);
nor U765 (N_765,N_169,N_421);
nand U766 (N_766,N_42,N_61);
or U767 (N_767,N_483,N_421);
or U768 (N_768,N_378,N_374);
nor U769 (N_769,N_301,N_93);
nor U770 (N_770,N_336,N_98);
or U771 (N_771,N_429,N_418);
nor U772 (N_772,N_480,N_417);
nand U773 (N_773,N_168,N_299);
and U774 (N_774,N_167,N_422);
and U775 (N_775,N_214,N_92);
and U776 (N_776,N_241,N_247);
nor U777 (N_777,N_119,N_371);
nor U778 (N_778,N_390,N_97);
and U779 (N_779,N_288,N_300);
nor U780 (N_780,N_400,N_274);
and U781 (N_781,N_151,N_253);
or U782 (N_782,N_394,N_304);
and U783 (N_783,N_482,N_319);
or U784 (N_784,N_496,N_212);
or U785 (N_785,N_299,N_377);
nor U786 (N_786,N_126,N_55);
nand U787 (N_787,N_229,N_405);
nand U788 (N_788,N_427,N_423);
and U789 (N_789,N_217,N_346);
xor U790 (N_790,N_150,N_153);
and U791 (N_791,N_187,N_419);
and U792 (N_792,N_287,N_197);
and U793 (N_793,N_33,N_19);
nor U794 (N_794,N_259,N_220);
nor U795 (N_795,N_72,N_305);
nand U796 (N_796,N_336,N_44);
xor U797 (N_797,N_226,N_453);
and U798 (N_798,N_65,N_247);
and U799 (N_799,N_125,N_297);
and U800 (N_800,N_208,N_334);
nand U801 (N_801,N_268,N_192);
nand U802 (N_802,N_204,N_17);
nor U803 (N_803,N_324,N_343);
and U804 (N_804,N_351,N_15);
nor U805 (N_805,N_142,N_295);
and U806 (N_806,N_136,N_4);
nor U807 (N_807,N_175,N_1);
nand U808 (N_808,N_183,N_21);
and U809 (N_809,N_75,N_223);
or U810 (N_810,N_50,N_341);
nand U811 (N_811,N_202,N_345);
and U812 (N_812,N_311,N_406);
or U813 (N_813,N_485,N_69);
xnor U814 (N_814,N_272,N_13);
nor U815 (N_815,N_60,N_408);
or U816 (N_816,N_224,N_106);
nand U817 (N_817,N_474,N_432);
and U818 (N_818,N_328,N_87);
and U819 (N_819,N_147,N_452);
nor U820 (N_820,N_471,N_360);
and U821 (N_821,N_211,N_483);
and U822 (N_822,N_339,N_391);
nor U823 (N_823,N_169,N_136);
or U824 (N_824,N_343,N_192);
xor U825 (N_825,N_118,N_21);
and U826 (N_826,N_399,N_476);
nor U827 (N_827,N_40,N_55);
or U828 (N_828,N_339,N_350);
nand U829 (N_829,N_2,N_386);
or U830 (N_830,N_177,N_222);
nor U831 (N_831,N_63,N_247);
and U832 (N_832,N_261,N_432);
nand U833 (N_833,N_64,N_466);
or U834 (N_834,N_283,N_327);
nand U835 (N_835,N_492,N_389);
and U836 (N_836,N_289,N_58);
nor U837 (N_837,N_113,N_89);
or U838 (N_838,N_119,N_64);
xnor U839 (N_839,N_348,N_74);
nand U840 (N_840,N_22,N_469);
or U841 (N_841,N_125,N_280);
nor U842 (N_842,N_497,N_329);
nor U843 (N_843,N_147,N_244);
and U844 (N_844,N_187,N_184);
and U845 (N_845,N_4,N_325);
nor U846 (N_846,N_235,N_499);
or U847 (N_847,N_482,N_348);
nor U848 (N_848,N_298,N_418);
and U849 (N_849,N_91,N_383);
nand U850 (N_850,N_242,N_181);
and U851 (N_851,N_235,N_209);
or U852 (N_852,N_352,N_277);
nor U853 (N_853,N_58,N_188);
nand U854 (N_854,N_228,N_171);
and U855 (N_855,N_259,N_486);
and U856 (N_856,N_67,N_162);
or U857 (N_857,N_364,N_453);
nand U858 (N_858,N_32,N_221);
or U859 (N_859,N_338,N_88);
nand U860 (N_860,N_8,N_263);
nor U861 (N_861,N_340,N_30);
nor U862 (N_862,N_110,N_355);
and U863 (N_863,N_198,N_462);
or U864 (N_864,N_416,N_394);
nand U865 (N_865,N_268,N_400);
nand U866 (N_866,N_477,N_423);
nor U867 (N_867,N_250,N_39);
nand U868 (N_868,N_15,N_453);
nand U869 (N_869,N_203,N_51);
or U870 (N_870,N_77,N_187);
and U871 (N_871,N_453,N_21);
and U872 (N_872,N_455,N_248);
and U873 (N_873,N_251,N_382);
nand U874 (N_874,N_458,N_251);
or U875 (N_875,N_22,N_12);
nor U876 (N_876,N_381,N_476);
nor U877 (N_877,N_101,N_26);
and U878 (N_878,N_133,N_293);
nor U879 (N_879,N_78,N_260);
or U880 (N_880,N_20,N_303);
or U881 (N_881,N_51,N_266);
and U882 (N_882,N_183,N_171);
nand U883 (N_883,N_388,N_238);
or U884 (N_884,N_283,N_224);
or U885 (N_885,N_92,N_31);
nor U886 (N_886,N_409,N_287);
and U887 (N_887,N_221,N_319);
or U888 (N_888,N_291,N_166);
or U889 (N_889,N_301,N_375);
nor U890 (N_890,N_304,N_193);
nand U891 (N_891,N_5,N_68);
or U892 (N_892,N_232,N_11);
and U893 (N_893,N_192,N_455);
nor U894 (N_894,N_351,N_242);
nand U895 (N_895,N_51,N_108);
or U896 (N_896,N_273,N_446);
nor U897 (N_897,N_211,N_123);
and U898 (N_898,N_261,N_333);
and U899 (N_899,N_317,N_201);
and U900 (N_900,N_262,N_345);
xor U901 (N_901,N_241,N_274);
and U902 (N_902,N_332,N_74);
xor U903 (N_903,N_80,N_450);
or U904 (N_904,N_151,N_363);
and U905 (N_905,N_246,N_303);
and U906 (N_906,N_496,N_353);
nand U907 (N_907,N_316,N_283);
nor U908 (N_908,N_177,N_54);
nor U909 (N_909,N_441,N_89);
nand U910 (N_910,N_184,N_387);
nor U911 (N_911,N_306,N_448);
nand U912 (N_912,N_146,N_357);
or U913 (N_913,N_74,N_301);
xnor U914 (N_914,N_406,N_288);
or U915 (N_915,N_478,N_207);
nand U916 (N_916,N_54,N_357);
and U917 (N_917,N_40,N_369);
and U918 (N_918,N_40,N_225);
nand U919 (N_919,N_148,N_18);
or U920 (N_920,N_399,N_219);
nand U921 (N_921,N_164,N_4);
or U922 (N_922,N_300,N_480);
nor U923 (N_923,N_34,N_79);
nand U924 (N_924,N_497,N_381);
nand U925 (N_925,N_483,N_455);
nand U926 (N_926,N_141,N_488);
nand U927 (N_927,N_405,N_227);
or U928 (N_928,N_267,N_364);
nor U929 (N_929,N_26,N_243);
nand U930 (N_930,N_398,N_40);
or U931 (N_931,N_151,N_86);
and U932 (N_932,N_432,N_498);
nand U933 (N_933,N_108,N_258);
and U934 (N_934,N_408,N_58);
and U935 (N_935,N_435,N_80);
or U936 (N_936,N_404,N_415);
nor U937 (N_937,N_310,N_161);
or U938 (N_938,N_228,N_336);
or U939 (N_939,N_380,N_115);
nor U940 (N_940,N_22,N_234);
and U941 (N_941,N_393,N_457);
nand U942 (N_942,N_377,N_354);
nand U943 (N_943,N_182,N_317);
nand U944 (N_944,N_148,N_461);
nor U945 (N_945,N_346,N_310);
or U946 (N_946,N_187,N_103);
nor U947 (N_947,N_405,N_248);
and U948 (N_948,N_163,N_405);
nor U949 (N_949,N_253,N_333);
nand U950 (N_950,N_61,N_236);
nor U951 (N_951,N_269,N_18);
nand U952 (N_952,N_122,N_171);
nand U953 (N_953,N_436,N_91);
xnor U954 (N_954,N_193,N_226);
nor U955 (N_955,N_0,N_146);
and U956 (N_956,N_355,N_429);
nor U957 (N_957,N_384,N_367);
or U958 (N_958,N_89,N_486);
nor U959 (N_959,N_497,N_229);
nand U960 (N_960,N_367,N_266);
and U961 (N_961,N_198,N_309);
and U962 (N_962,N_328,N_194);
nor U963 (N_963,N_460,N_372);
nand U964 (N_964,N_191,N_281);
or U965 (N_965,N_344,N_144);
and U966 (N_966,N_34,N_338);
or U967 (N_967,N_451,N_465);
nor U968 (N_968,N_243,N_287);
or U969 (N_969,N_313,N_338);
nor U970 (N_970,N_5,N_158);
nand U971 (N_971,N_211,N_456);
or U972 (N_972,N_52,N_344);
or U973 (N_973,N_356,N_358);
nand U974 (N_974,N_417,N_499);
nand U975 (N_975,N_205,N_389);
nor U976 (N_976,N_20,N_279);
and U977 (N_977,N_107,N_349);
xnor U978 (N_978,N_494,N_457);
or U979 (N_979,N_207,N_346);
nand U980 (N_980,N_409,N_284);
nand U981 (N_981,N_358,N_300);
nand U982 (N_982,N_438,N_382);
and U983 (N_983,N_137,N_431);
nor U984 (N_984,N_138,N_314);
nor U985 (N_985,N_73,N_214);
nand U986 (N_986,N_216,N_474);
and U987 (N_987,N_354,N_90);
nor U988 (N_988,N_257,N_140);
and U989 (N_989,N_186,N_84);
and U990 (N_990,N_466,N_423);
nor U991 (N_991,N_41,N_116);
and U992 (N_992,N_470,N_139);
or U993 (N_993,N_314,N_216);
or U994 (N_994,N_235,N_148);
nand U995 (N_995,N_25,N_422);
or U996 (N_996,N_440,N_423);
or U997 (N_997,N_72,N_345);
nand U998 (N_998,N_329,N_468);
or U999 (N_999,N_318,N_478);
or U1000 (N_1000,N_870,N_900);
xnor U1001 (N_1001,N_626,N_763);
or U1002 (N_1002,N_618,N_876);
and U1003 (N_1003,N_556,N_836);
nor U1004 (N_1004,N_770,N_982);
or U1005 (N_1005,N_885,N_949);
and U1006 (N_1006,N_925,N_608);
and U1007 (N_1007,N_506,N_514);
nand U1008 (N_1008,N_839,N_599);
or U1009 (N_1009,N_808,N_968);
and U1010 (N_1010,N_892,N_877);
or U1011 (N_1011,N_894,N_541);
nor U1012 (N_1012,N_585,N_979);
and U1013 (N_1013,N_572,N_891);
or U1014 (N_1014,N_960,N_825);
nor U1015 (N_1015,N_622,N_881);
or U1016 (N_1016,N_577,N_997);
nand U1017 (N_1017,N_644,N_629);
and U1018 (N_1018,N_587,N_905);
or U1019 (N_1019,N_628,N_729);
or U1020 (N_1020,N_956,N_929);
nand U1021 (N_1021,N_961,N_927);
nor U1022 (N_1022,N_803,N_831);
nor U1023 (N_1023,N_589,N_606);
nand U1024 (N_1024,N_651,N_978);
or U1025 (N_1025,N_700,N_914);
or U1026 (N_1026,N_748,N_757);
nand U1027 (N_1027,N_665,N_650);
nor U1028 (N_1028,N_911,N_601);
nand U1029 (N_1029,N_709,N_687);
or U1030 (N_1030,N_612,N_584);
and U1031 (N_1031,N_965,N_641);
or U1032 (N_1032,N_555,N_815);
nand U1033 (N_1033,N_805,N_516);
nand U1034 (N_1034,N_916,N_718);
or U1035 (N_1035,N_594,N_691);
and U1036 (N_1036,N_731,N_926);
or U1037 (N_1037,N_851,N_521);
and U1038 (N_1038,N_844,N_546);
and U1039 (N_1039,N_645,N_795);
and U1040 (N_1040,N_526,N_602);
and U1041 (N_1041,N_898,N_674);
and U1042 (N_1042,N_764,N_551);
and U1043 (N_1043,N_828,N_820);
nor U1044 (N_1044,N_980,N_970);
nor U1045 (N_1045,N_532,N_504);
or U1046 (N_1046,N_793,N_663);
or U1047 (N_1047,N_574,N_837);
and U1048 (N_1048,N_936,N_821);
and U1049 (N_1049,N_642,N_661);
or U1050 (N_1050,N_706,N_550);
nor U1051 (N_1051,N_710,N_524);
or U1052 (N_1052,N_890,N_517);
nand U1053 (N_1053,N_684,N_683);
nand U1054 (N_1054,N_995,N_775);
and U1055 (N_1055,N_809,N_562);
nand U1056 (N_1056,N_946,N_848);
nand U1057 (N_1057,N_845,N_909);
and U1058 (N_1058,N_860,N_826);
or U1059 (N_1059,N_801,N_669);
and U1060 (N_1060,N_648,N_915);
nor U1061 (N_1061,N_662,N_954);
or U1062 (N_1062,N_944,N_868);
and U1063 (N_1063,N_694,N_703);
nor U1064 (N_1064,N_973,N_611);
nor U1065 (N_1065,N_981,N_552);
and U1066 (N_1066,N_505,N_678);
or U1067 (N_1067,N_908,N_668);
and U1068 (N_1068,N_922,N_639);
and U1069 (N_1069,N_571,N_969);
and U1070 (N_1070,N_653,N_971);
and U1071 (N_1071,N_972,N_704);
nand U1072 (N_1072,N_769,N_623);
or U1073 (N_1073,N_903,N_658);
nand U1074 (N_1074,N_660,N_986);
and U1075 (N_1075,N_761,N_525);
nor U1076 (N_1076,N_696,N_531);
nand U1077 (N_1077,N_701,N_707);
nand U1078 (N_1078,N_543,N_605);
nor U1079 (N_1079,N_588,N_907);
nor U1080 (N_1080,N_666,N_615);
and U1081 (N_1081,N_721,N_698);
or U1082 (N_1082,N_967,N_874);
nand U1083 (N_1083,N_865,N_501);
nand U1084 (N_1084,N_640,N_590);
nor U1085 (N_1085,N_859,N_542);
or U1086 (N_1086,N_869,N_933);
nand U1087 (N_1087,N_893,N_811);
nand U1088 (N_1088,N_744,N_964);
and U1089 (N_1089,N_609,N_654);
xor U1090 (N_1090,N_784,N_554);
or U1091 (N_1091,N_561,N_785);
nor U1092 (N_1092,N_579,N_742);
nor U1093 (N_1093,N_850,N_724);
nor U1094 (N_1094,N_994,N_682);
nor U1095 (N_1095,N_823,N_923);
and U1096 (N_1096,N_540,N_766);
or U1097 (N_1097,N_722,N_686);
and U1098 (N_1098,N_739,N_948);
or U1099 (N_1099,N_617,N_988);
or U1100 (N_1100,N_557,N_685);
nand U1101 (N_1101,N_732,N_798);
and U1102 (N_1102,N_671,N_632);
nor U1103 (N_1103,N_591,N_670);
nand U1104 (N_1104,N_902,N_595);
or U1105 (N_1105,N_963,N_884);
and U1106 (N_1106,N_509,N_690);
nor U1107 (N_1107,N_921,N_520);
or U1108 (N_1108,N_790,N_560);
or U1109 (N_1109,N_657,N_987);
nor U1110 (N_1110,N_582,N_693);
or U1111 (N_1111,N_538,N_941);
nand U1112 (N_1112,N_810,N_777);
nand U1113 (N_1113,N_912,N_985);
and U1114 (N_1114,N_723,N_887);
nor U1115 (N_1115,N_992,N_652);
and U1116 (N_1116,N_547,N_773);
or U1117 (N_1117,N_635,N_888);
nor U1118 (N_1118,N_816,N_958);
nand U1119 (N_1119,N_673,N_719);
or U1120 (N_1120,N_889,N_990);
or U1121 (N_1121,N_867,N_791);
nand U1122 (N_1122,N_563,N_737);
nor U1123 (N_1123,N_814,N_834);
or U1124 (N_1124,N_975,N_920);
and U1125 (N_1125,N_897,N_537);
nand U1126 (N_1126,N_679,N_846);
and U1127 (N_1127,N_756,N_910);
nand U1128 (N_1128,N_559,N_849);
or U1129 (N_1129,N_842,N_507);
nand U1130 (N_1130,N_730,N_533);
and U1131 (N_1131,N_812,N_676);
nand U1132 (N_1132,N_829,N_558);
nand U1133 (N_1133,N_774,N_976);
or U1134 (N_1134,N_983,N_932);
and U1135 (N_1135,N_545,N_959);
nor U1136 (N_1136,N_720,N_529);
or U1137 (N_1137,N_530,N_861);
nor U1138 (N_1138,N_621,N_699);
nor U1139 (N_1139,N_786,N_503);
nor U1140 (N_1140,N_797,N_536);
nor U1141 (N_1141,N_535,N_755);
nor U1142 (N_1142,N_638,N_962);
nand U1143 (N_1143,N_800,N_508);
nor U1144 (N_1144,N_855,N_938);
and U1145 (N_1145,N_767,N_840);
or U1146 (N_1146,N_620,N_752);
nand U1147 (N_1147,N_802,N_548);
or U1148 (N_1148,N_583,N_586);
or U1149 (N_1149,N_573,N_689);
or U1150 (N_1150,N_813,N_581);
nand U1151 (N_1151,N_955,N_511);
xor U1152 (N_1152,N_883,N_899);
nand U1153 (N_1153,N_760,N_569);
nor U1154 (N_1154,N_570,N_649);
and U1155 (N_1155,N_634,N_523);
nand U1156 (N_1156,N_534,N_715);
or U1157 (N_1157,N_789,N_780);
or U1158 (N_1158,N_950,N_672);
nor U1159 (N_1159,N_853,N_952);
or U1160 (N_1160,N_843,N_762);
nand U1161 (N_1161,N_940,N_782);
nand U1162 (N_1162,N_847,N_643);
and U1163 (N_1163,N_600,N_625);
or U1164 (N_1164,N_768,N_953);
nand U1165 (N_1165,N_928,N_688);
nor U1166 (N_1166,N_734,N_799);
or U1167 (N_1167,N_913,N_937);
nor U1168 (N_1168,N_779,N_794);
and U1169 (N_1169,N_746,N_675);
or U1170 (N_1170,N_667,N_714);
nor U1171 (N_1171,N_781,N_637);
nand U1172 (N_1172,N_984,N_872);
nor U1173 (N_1173,N_616,N_917);
or U1174 (N_1174,N_646,N_738);
nor U1175 (N_1175,N_568,N_610);
and U1176 (N_1176,N_864,N_624);
or U1177 (N_1177,N_655,N_603);
nand U1178 (N_1178,N_627,N_743);
or U1179 (N_1179,N_631,N_878);
nand U1180 (N_1180,N_996,N_566);
nor U1181 (N_1181,N_822,N_515);
nor U1182 (N_1182,N_510,N_765);
nor U1183 (N_1183,N_575,N_862);
and U1184 (N_1184,N_677,N_827);
or U1185 (N_1185,N_792,N_711);
nor U1186 (N_1186,N_957,N_614);
nand U1187 (N_1187,N_747,N_713);
and U1188 (N_1188,N_919,N_549);
and U1189 (N_1189,N_716,N_807);
nand U1190 (N_1190,N_783,N_680);
nand U1191 (N_1191,N_522,N_873);
and U1192 (N_1192,N_998,N_796);
nand U1193 (N_1193,N_871,N_527);
or U1194 (N_1194,N_564,N_727);
and U1195 (N_1195,N_934,N_702);
or U1196 (N_1196,N_513,N_945);
nor U1197 (N_1197,N_596,N_924);
nor U1198 (N_1198,N_630,N_906);
nor U1199 (N_1199,N_567,N_857);
or U1200 (N_1200,N_966,N_604);
or U1201 (N_1201,N_977,N_771);
nor U1202 (N_1202,N_712,N_758);
and U1203 (N_1203,N_951,N_772);
or U1204 (N_1204,N_863,N_659);
nand U1205 (N_1205,N_901,N_695);
nand U1206 (N_1206,N_776,N_544);
or U1207 (N_1207,N_824,N_750);
and U1208 (N_1208,N_692,N_880);
or U1209 (N_1209,N_512,N_735);
nand U1210 (N_1210,N_751,N_882);
nor U1211 (N_1211,N_597,N_759);
nor U1212 (N_1212,N_835,N_947);
or U1213 (N_1213,N_858,N_754);
nand U1214 (N_1214,N_939,N_619);
or U1215 (N_1215,N_833,N_841);
or U1216 (N_1216,N_999,N_519);
and U1217 (N_1217,N_832,N_817);
nor U1218 (N_1218,N_886,N_942);
nand U1219 (N_1219,N_580,N_681);
or U1220 (N_1220,N_741,N_819);
nor U1221 (N_1221,N_728,N_788);
nand U1222 (N_1222,N_787,N_806);
and U1223 (N_1223,N_656,N_930);
or U1224 (N_1224,N_664,N_725);
or U1225 (N_1225,N_854,N_993);
nor U1226 (N_1226,N_852,N_593);
nand U1227 (N_1227,N_935,N_745);
or U1228 (N_1228,N_705,N_518);
or U1229 (N_1229,N_895,N_804);
or U1230 (N_1230,N_607,N_502);
and U1231 (N_1231,N_989,N_753);
or U1232 (N_1232,N_553,N_636);
or U1233 (N_1233,N_647,N_717);
or U1234 (N_1234,N_991,N_598);
nor U1235 (N_1235,N_578,N_500);
nor U1236 (N_1236,N_749,N_879);
nor U1237 (N_1237,N_736,N_778);
and U1238 (N_1238,N_565,N_613);
and U1239 (N_1239,N_866,N_528);
or U1240 (N_1240,N_918,N_896);
nand U1241 (N_1241,N_592,N_726);
or U1242 (N_1242,N_539,N_697);
or U1243 (N_1243,N_818,N_838);
and U1244 (N_1244,N_830,N_904);
or U1245 (N_1245,N_943,N_733);
nor U1246 (N_1246,N_708,N_875);
xnor U1247 (N_1247,N_931,N_974);
nor U1248 (N_1248,N_740,N_856);
or U1249 (N_1249,N_576,N_633);
nor U1250 (N_1250,N_853,N_854);
or U1251 (N_1251,N_515,N_891);
nor U1252 (N_1252,N_814,N_636);
nand U1253 (N_1253,N_834,N_900);
and U1254 (N_1254,N_700,N_634);
or U1255 (N_1255,N_908,N_724);
nor U1256 (N_1256,N_639,N_753);
and U1257 (N_1257,N_777,N_553);
and U1258 (N_1258,N_600,N_695);
nor U1259 (N_1259,N_858,N_692);
xnor U1260 (N_1260,N_660,N_691);
and U1261 (N_1261,N_969,N_974);
nand U1262 (N_1262,N_867,N_744);
nand U1263 (N_1263,N_754,N_965);
or U1264 (N_1264,N_785,N_554);
or U1265 (N_1265,N_895,N_983);
nor U1266 (N_1266,N_815,N_683);
nand U1267 (N_1267,N_684,N_963);
nand U1268 (N_1268,N_895,N_794);
nor U1269 (N_1269,N_762,N_860);
nand U1270 (N_1270,N_935,N_882);
or U1271 (N_1271,N_515,N_853);
and U1272 (N_1272,N_666,N_710);
and U1273 (N_1273,N_700,N_680);
and U1274 (N_1274,N_706,N_700);
or U1275 (N_1275,N_999,N_587);
nor U1276 (N_1276,N_893,N_503);
and U1277 (N_1277,N_904,N_861);
nand U1278 (N_1278,N_623,N_747);
and U1279 (N_1279,N_650,N_689);
or U1280 (N_1280,N_884,N_983);
nor U1281 (N_1281,N_949,N_583);
or U1282 (N_1282,N_959,N_640);
and U1283 (N_1283,N_744,N_897);
or U1284 (N_1284,N_503,N_750);
nand U1285 (N_1285,N_622,N_815);
or U1286 (N_1286,N_536,N_587);
or U1287 (N_1287,N_811,N_998);
and U1288 (N_1288,N_784,N_576);
nand U1289 (N_1289,N_681,N_527);
and U1290 (N_1290,N_611,N_560);
nand U1291 (N_1291,N_623,N_695);
nand U1292 (N_1292,N_953,N_658);
nor U1293 (N_1293,N_840,N_900);
nand U1294 (N_1294,N_729,N_987);
nand U1295 (N_1295,N_963,N_692);
xor U1296 (N_1296,N_838,N_767);
or U1297 (N_1297,N_637,N_794);
and U1298 (N_1298,N_770,N_522);
and U1299 (N_1299,N_702,N_849);
nor U1300 (N_1300,N_613,N_582);
nand U1301 (N_1301,N_913,N_689);
nand U1302 (N_1302,N_503,N_832);
or U1303 (N_1303,N_814,N_968);
nand U1304 (N_1304,N_884,N_641);
nor U1305 (N_1305,N_543,N_555);
nor U1306 (N_1306,N_878,N_628);
and U1307 (N_1307,N_986,N_858);
nand U1308 (N_1308,N_769,N_727);
nand U1309 (N_1309,N_768,N_624);
or U1310 (N_1310,N_775,N_819);
nor U1311 (N_1311,N_746,N_520);
nor U1312 (N_1312,N_561,N_648);
or U1313 (N_1313,N_643,N_864);
nand U1314 (N_1314,N_881,N_688);
or U1315 (N_1315,N_964,N_691);
or U1316 (N_1316,N_700,N_554);
and U1317 (N_1317,N_698,N_542);
xnor U1318 (N_1318,N_875,N_765);
or U1319 (N_1319,N_975,N_950);
and U1320 (N_1320,N_503,N_908);
nor U1321 (N_1321,N_951,N_849);
and U1322 (N_1322,N_879,N_812);
or U1323 (N_1323,N_530,N_826);
or U1324 (N_1324,N_906,N_876);
nor U1325 (N_1325,N_687,N_678);
or U1326 (N_1326,N_827,N_580);
xnor U1327 (N_1327,N_709,N_625);
nor U1328 (N_1328,N_532,N_832);
and U1329 (N_1329,N_596,N_737);
or U1330 (N_1330,N_984,N_922);
nand U1331 (N_1331,N_614,N_959);
nor U1332 (N_1332,N_627,N_816);
and U1333 (N_1333,N_522,N_785);
nor U1334 (N_1334,N_947,N_744);
nor U1335 (N_1335,N_809,N_764);
nand U1336 (N_1336,N_582,N_785);
or U1337 (N_1337,N_728,N_786);
nor U1338 (N_1338,N_857,N_502);
nand U1339 (N_1339,N_808,N_597);
or U1340 (N_1340,N_626,N_943);
or U1341 (N_1341,N_715,N_958);
nand U1342 (N_1342,N_955,N_507);
and U1343 (N_1343,N_750,N_968);
nand U1344 (N_1344,N_892,N_712);
nor U1345 (N_1345,N_893,N_954);
or U1346 (N_1346,N_636,N_748);
and U1347 (N_1347,N_833,N_907);
nand U1348 (N_1348,N_939,N_923);
nor U1349 (N_1349,N_997,N_777);
nor U1350 (N_1350,N_801,N_760);
and U1351 (N_1351,N_687,N_764);
and U1352 (N_1352,N_604,N_669);
or U1353 (N_1353,N_528,N_920);
nand U1354 (N_1354,N_996,N_937);
and U1355 (N_1355,N_800,N_997);
nand U1356 (N_1356,N_971,N_766);
nor U1357 (N_1357,N_524,N_822);
nor U1358 (N_1358,N_701,N_975);
nand U1359 (N_1359,N_908,N_833);
nand U1360 (N_1360,N_515,N_901);
and U1361 (N_1361,N_941,N_837);
nand U1362 (N_1362,N_811,N_654);
nor U1363 (N_1363,N_675,N_838);
and U1364 (N_1364,N_961,N_674);
and U1365 (N_1365,N_904,N_604);
and U1366 (N_1366,N_831,N_953);
and U1367 (N_1367,N_737,N_992);
or U1368 (N_1368,N_698,N_550);
or U1369 (N_1369,N_532,N_776);
and U1370 (N_1370,N_995,N_895);
nand U1371 (N_1371,N_866,N_647);
and U1372 (N_1372,N_873,N_600);
nor U1373 (N_1373,N_921,N_580);
and U1374 (N_1374,N_778,N_781);
nor U1375 (N_1375,N_919,N_838);
nor U1376 (N_1376,N_628,N_639);
xnor U1377 (N_1377,N_768,N_868);
nor U1378 (N_1378,N_909,N_597);
and U1379 (N_1379,N_641,N_755);
nor U1380 (N_1380,N_532,N_698);
nand U1381 (N_1381,N_960,N_911);
or U1382 (N_1382,N_629,N_758);
nor U1383 (N_1383,N_530,N_692);
nand U1384 (N_1384,N_631,N_568);
nor U1385 (N_1385,N_852,N_502);
or U1386 (N_1386,N_625,N_988);
nand U1387 (N_1387,N_545,N_765);
or U1388 (N_1388,N_756,N_787);
xor U1389 (N_1389,N_835,N_553);
and U1390 (N_1390,N_793,N_778);
nor U1391 (N_1391,N_991,N_751);
and U1392 (N_1392,N_928,N_601);
nand U1393 (N_1393,N_701,N_657);
and U1394 (N_1394,N_802,N_694);
or U1395 (N_1395,N_622,N_718);
or U1396 (N_1396,N_753,N_555);
or U1397 (N_1397,N_530,N_986);
nor U1398 (N_1398,N_856,N_684);
or U1399 (N_1399,N_661,N_546);
or U1400 (N_1400,N_739,N_726);
nand U1401 (N_1401,N_568,N_857);
or U1402 (N_1402,N_575,N_536);
xor U1403 (N_1403,N_872,N_504);
or U1404 (N_1404,N_647,N_624);
nand U1405 (N_1405,N_649,N_954);
and U1406 (N_1406,N_997,N_532);
or U1407 (N_1407,N_733,N_521);
or U1408 (N_1408,N_847,N_764);
nor U1409 (N_1409,N_841,N_816);
nor U1410 (N_1410,N_719,N_865);
nor U1411 (N_1411,N_510,N_891);
nand U1412 (N_1412,N_777,N_656);
nor U1413 (N_1413,N_880,N_570);
or U1414 (N_1414,N_974,N_987);
nand U1415 (N_1415,N_724,N_972);
nand U1416 (N_1416,N_992,N_809);
and U1417 (N_1417,N_691,N_951);
nor U1418 (N_1418,N_504,N_991);
or U1419 (N_1419,N_857,N_672);
nor U1420 (N_1420,N_570,N_970);
nor U1421 (N_1421,N_603,N_505);
or U1422 (N_1422,N_863,N_783);
and U1423 (N_1423,N_674,N_598);
nor U1424 (N_1424,N_578,N_529);
nor U1425 (N_1425,N_707,N_552);
and U1426 (N_1426,N_574,N_892);
nor U1427 (N_1427,N_927,N_781);
nor U1428 (N_1428,N_913,N_971);
and U1429 (N_1429,N_728,N_734);
nand U1430 (N_1430,N_787,N_576);
nand U1431 (N_1431,N_579,N_500);
and U1432 (N_1432,N_918,N_703);
nand U1433 (N_1433,N_834,N_691);
nand U1434 (N_1434,N_742,N_997);
nand U1435 (N_1435,N_999,N_892);
or U1436 (N_1436,N_579,N_816);
nor U1437 (N_1437,N_694,N_898);
and U1438 (N_1438,N_745,N_988);
or U1439 (N_1439,N_606,N_851);
and U1440 (N_1440,N_851,N_791);
nor U1441 (N_1441,N_735,N_501);
nand U1442 (N_1442,N_685,N_657);
nand U1443 (N_1443,N_954,N_845);
nor U1444 (N_1444,N_789,N_529);
and U1445 (N_1445,N_895,N_846);
or U1446 (N_1446,N_537,N_922);
nand U1447 (N_1447,N_962,N_744);
nand U1448 (N_1448,N_543,N_923);
nor U1449 (N_1449,N_895,N_670);
or U1450 (N_1450,N_664,N_791);
or U1451 (N_1451,N_522,N_724);
nor U1452 (N_1452,N_775,N_776);
nor U1453 (N_1453,N_532,N_775);
or U1454 (N_1454,N_629,N_538);
nor U1455 (N_1455,N_933,N_881);
or U1456 (N_1456,N_698,N_942);
nand U1457 (N_1457,N_952,N_616);
nand U1458 (N_1458,N_830,N_510);
nor U1459 (N_1459,N_639,N_743);
or U1460 (N_1460,N_541,N_712);
and U1461 (N_1461,N_880,N_534);
nor U1462 (N_1462,N_529,N_832);
or U1463 (N_1463,N_846,N_962);
nand U1464 (N_1464,N_999,N_962);
nor U1465 (N_1465,N_963,N_519);
nor U1466 (N_1466,N_791,N_972);
nor U1467 (N_1467,N_530,N_645);
or U1468 (N_1468,N_799,N_948);
and U1469 (N_1469,N_788,N_993);
nand U1470 (N_1470,N_716,N_929);
and U1471 (N_1471,N_606,N_727);
nor U1472 (N_1472,N_595,N_553);
nor U1473 (N_1473,N_618,N_623);
or U1474 (N_1474,N_644,N_627);
or U1475 (N_1475,N_534,N_664);
nor U1476 (N_1476,N_732,N_862);
nand U1477 (N_1477,N_938,N_829);
or U1478 (N_1478,N_905,N_615);
and U1479 (N_1479,N_556,N_664);
xor U1480 (N_1480,N_841,N_533);
or U1481 (N_1481,N_691,N_947);
nand U1482 (N_1482,N_896,N_669);
and U1483 (N_1483,N_675,N_688);
nand U1484 (N_1484,N_729,N_860);
or U1485 (N_1485,N_734,N_837);
and U1486 (N_1486,N_583,N_521);
nand U1487 (N_1487,N_866,N_641);
or U1488 (N_1488,N_745,N_548);
nand U1489 (N_1489,N_767,N_856);
nor U1490 (N_1490,N_555,N_647);
and U1491 (N_1491,N_687,N_534);
and U1492 (N_1492,N_829,N_547);
nand U1493 (N_1493,N_586,N_959);
or U1494 (N_1494,N_617,N_537);
nand U1495 (N_1495,N_734,N_593);
or U1496 (N_1496,N_502,N_608);
and U1497 (N_1497,N_513,N_970);
nor U1498 (N_1498,N_872,N_759);
nor U1499 (N_1499,N_933,N_872);
nand U1500 (N_1500,N_1422,N_1462);
and U1501 (N_1501,N_1398,N_1088);
nand U1502 (N_1502,N_1059,N_1317);
or U1503 (N_1503,N_1382,N_1034);
nor U1504 (N_1504,N_1303,N_1170);
nor U1505 (N_1505,N_1139,N_1058);
and U1506 (N_1506,N_1135,N_1356);
nor U1507 (N_1507,N_1030,N_1477);
or U1508 (N_1508,N_1402,N_1005);
or U1509 (N_1509,N_1429,N_1183);
nand U1510 (N_1510,N_1033,N_1383);
or U1511 (N_1511,N_1066,N_1369);
and U1512 (N_1512,N_1167,N_1182);
nor U1513 (N_1513,N_1067,N_1334);
or U1514 (N_1514,N_1400,N_1372);
nand U1515 (N_1515,N_1096,N_1045);
nor U1516 (N_1516,N_1436,N_1404);
xnor U1517 (N_1517,N_1322,N_1163);
and U1518 (N_1518,N_1439,N_1407);
and U1519 (N_1519,N_1038,N_1287);
nor U1520 (N_1520,N_1017,N_1179);
nor U1521 (N_1521,N_1390,N_1242);
and U1522 (N_1522,N_1112,N_1450);
nor U1523 (N_1523,N_1110,N_1325);
and U1524 (N_1524,N_1251,N_1387);
nor U1525 (N_1525,N_1070,N_1246);
or U1526 (N_1526,N_1190,N_1457);
and U1527 (N_1527,N_1233,N_1037);
nand U1528 (N_1528,N_1078,N_1226);
nor U1529 (N_1529,N_1272,N_1494);
or U1530 (N_1530,N_1275,N_1492);
nand U1531 (N_1531,N_1090,N_1172);
nor U1532 (N_1532,N_1244,N_1248);
xor U1533 (N_1533,N_1164,N_1136);
or U1534 (N_1534,N_1147,N_1257);
or U1535 (N_1535,N_1211,N_1262);
nand U1536 (N_1536,N_1227,N_1294);
nand U1537 (N_1537,N_1203,N_1150);
nor U1538 (N_1538,N_1447,N_1384);
nand U1539 (N_1539,N_1185,N_1329);
and U1540 (N_1540,N_1451,N_1015);
and U1541 (N_1541,N_1003,N_1336);
and U1542 (N_1542,N_1491,N_1249);
and U1543 (N_1543,N_1016,N_1188);
or U1544 (N_1544,N_1344,N_1271);
and U1545 (N_1545,N_1231,N_1121);
and U1546 (N_1546,N_1419,N_1061);
and U1547 (N_1547,N_1196,N_1499);
nor U1548 (N_1548,N_1055,N_1254);
nand U1549 (N_1549,N_1452,N_1187);
and U1550 (N_1550,N_1392,N_1471);
nor U1551 (N_1551,N_1143,N_1308);
nand U1552 (N_1552,N_1414,N_1213);
and U1553 (N_1553,N_1026,N_1331);
and U1554 (N_1554,N_1201,N_1069);
nor U1555 (N_1555,N_1006,N_1218);
and U1556 (N_1556,N_1458,N_1286);
or U1557 (N_1557,N_1305,N_1367);
nor U1558 (N_1558,N_1184,N_1460);
xor U1559 (N_1559,N_1497,N_1145);
nand U1560 (N_1560,N_1191,N_1431);
nor U1561 (N_1561,N_1235,N_1194);
and U1562 (N_1562,N_1442,N_1337);
nor U1563 (N_1563,N_1154,N_1092);
nor U1564 (N_1564,N_1039,N_1330);
nor U1565 (N_1565,N_1130,N_1314);
or U1566 (N_1566,N_1470,N_1459);
nand U1567 (N_1567,N_1274,N_1104);
and U1568 (N_1568,N_1118,N_1009);
and U1569 (N_1569,N_1373,N_1386);
or U1570 (N_1570,N_1079,N_1239);
nand U1571 (N_1571,N_1115,N_1036);
nand U1572 (N_1572,N_1119,N_1173);
or U1573 (N_1573,N_1432,N_1498);
and U1574 (N_1574,N_1427,N_1266);
and U1575 (N_1575,N_1077,N_1290);
nand U1576 (N_1576,N_1466,N_1264);
or U1577 (N_1577,N_1029,N_1347);
nor U1578 (N_1578,N_1332,N_1171);
nor U1579 (N_1579,N_1043,N_1405);
or U1580 (N_1580,N_1062,N_1278);
and U1581 (N_1581,N_1221,N_1023);
nand U1582 (N_1582,N_1002,N_1052);
and U1583 (N_1583,N_1065,N_1165);
or U1584 (N_1584,N_1178,N_1391);
nor U1585 (N_1585,N_1376,N_1444);
or U1586 (N_1586,N_1351,N_1401);
nand U1587 (N_1587,N_1484,N_1157);
or U1588 (N_1588,N_1035,N_1028);
nand U1589 (N_1589,N_1428,N_1388);
and U1590 (N_1590,N_1081,N_1333);
or U1591 (N_1591,N_1189,N_1199);
nand U1592 (N_1592,N_1364,N_1206);
nor U1593 (N_1593,N_1479,N_1197);
xnor U1594 (N_1594,N_1365,N_1472);
nor U1595 (N_1595,N_1007,N_1141);
and U1596 (N_1596,N_1350,N_1378);
and U1597 (N_1597,N_1421,N_1265);
or U1598 (N_1598,N_1004,N_1267);
or U1599 (N_1599,N_1232,N_1486);
or U1600 (N_1600,N_1108,N_1072);
nor U1601 (N_1601,N_1149,N_1126);
and U1602 (N_1602,N_1449,N_1053);
or U1603 (N_1603,N_1087,N_1225);
nor U1604 (N_1604,N_1409,N_1389);
and U1605 (N_1605,N_1027,N_1056);
nor U1606 (N_1606,N_1301,N_1291);
and U1607 (N_1607,N_1379,N_1202);
nand U1608 (N_1608,N_1480,N_1073);
and U1609 (N_1609,N_1151,N_1464);
or U1610 (N_1610,N_1313,N_1021);
and U1611 (N_1611,N_1487,N_1395);
and U1612 (N_1612,N_1293,N_1277);
nand U1613 (N_1613,N_1496,N_1396);
or U1614 (N_1614,N_1476,N_1403);
or U1615 (N_1615,N_1381,N_1416);
and U1616 (N_1616,N_1175,N_1474);
and U1617 (N_1617,N_1495,N_1234);
and U1618 (N_1618,N_1100,N_1455);
and U1619 (N_1619,N_1148,N_1013);
nand U1620 (N_1620,N_1411,N_1155);
nand U1621 (N_1621,N_1423,N_1327);
nand U1622 (N_1622,N_1425,N_1068);
or U1623 (N_1623,N_1210,N_1114);
and U1624 (N_1624,N_1144,N_1306);
xor U1625 (N_1625,N_1268,N_1054);
or U1626 (N_1626,N_1128,N_1298);
nand U1627 (N_1627,N_1362,N_1352);
or U1628 (N_1628,N_1319,N_1214);
or U1629 (N_1629,N_1340,N_1270);
or U1630 (N_1630,N_1103,N_1074);
nand U1631 (N_1631,N_1415,N_1397);
nor U1632 (N_1632,N_1263,N_1208);
or U1633 (N_1633,N_1140,N_1348);
nor U1634 (N_1634,N_1134,N_1010);
nand U1635 (N_1635,N_1138,N_1323);
nand U1636 (N_1636,N_1261,N_1040);
or U1637 (N_1637,N_1209,N_1368);
xnor U1638 (N_1638,N_1309,N_1292);
and U1639 (N_1639,N_1160,N_1106);
nor U1640 (N_1640,N_1111,N_1342);
nor U1641 (N_1641,N_1241,N_1282);
and U1642 (N_1642,N_1085,N_1426);
nor U1643 (N_1643,N_1156,N_1176);
nor U1644 (N_1644,N_1080,N_1064);
xor U1645 (N_1645,N_1253,N_1424);
and U1646 (N_1646,N_1247,N_1363);
nor U1647 (N_1647,N_1252,N_1394);
nand U1648 (N_1648,N_1014,N_1276);
nor U1649 (N_1649,N_1255,N_1285);
or U1650 (N_1650,N_1137,N_1366);
nor U1651 (N_1651,N_1412,N_1359);
or U1652 (N_1652,N_1297,N_1049);
nand U1653 (N_1653,N_1453,N_1230);
or U1654 (N_1654,N_1012,N_1380);
or U1655 (N_1655,N_1228,N_1483);
nor U1656 (N_1656,N_1102,N_1299);
or U1657 (N_1657,N_1169,N_1441);
nor U1658 (N_1658,N_1360,N_1204);
xnor U1659 (N_1659,N_1469,N_1098);
and U1660 (N_1660,N_1042,N_1454);
nand U1661 (N_1661,N_1326,N_1166);
or U1662 (N_1662,N_1236,N_1355);
nand U1663 (N_1663,N_1418,N_1001);
or U1664 (N_1664,N_1320,N_1312);
and U1665 (N_1665,N_1060,N_1237);
or U1666 (N_1666,N_1446,N_1307);
nand U1667 (N_1667,N_1229,N_1180);
nor U1668 (N_1668,N_1093,N_1024);
nand U1669 (N_1669,N_1046,N_1349);
and U1670 (N_1670,N_1456,N_1113);
and U1671 (N_1671,N_1280,N_1374);
or U1672 (N_1672,N_1105,N_1063);
or U1673 (N_1673,N_1127,N_1243);
or U1674 (N_1674,N_1025,N_1047);
nand U1675 (N_1675,N_1430,N_1475);
nand U1676 (N_1676,N_1273,N_1324);
and U1677 (N_1677,N_1082,N_1399);
nand U1678 (N_1678,N_1361,N_1050);
and U1679 (N_1679,N_1107,N_1259);
xnor U1680 (N_1680,N_1289,N_1129);
and U1681 (N_1681,N_1200,N_1022);
nand U1682 (N_1682,N_1339,N_1142);
nand U1683 (N_1683,N_1094,N_1192);
nor U1684 (N_1684,N_1433,N_1000);
nand U1685 (N_1685,N_1260,N_1057);
nand U1686 (N_1686,N_1296,N_1153);
nor U1687 (N_1687,N_1420,N_1304);
nand U1688 (N_1688,N_1133,N_1250);
or U1689 (N_1689,N_1406,N_1269);
and U1690 (N_1690,N_1099,N_1410);
nor U1691 (N_1691,N_1120,N_1256);
nand U1692 (N_1692,N_1161,N_1467);
or U1693 (N_1693,N_1375,N_1101);
and U1694 (N_1694,N_1358,N_1125);
and U1695 (N_1695,N_1168,N_1343);
and U1696 (N_1696,N_1315,N_1437);
or U1697 (N_1697,N_1089,N_1489);
or U1698 (N_1698,N_1220,N_1493);
nor U1699 (N_1699,N_1044,N_1481);
nand U1700 (N_1700,N_1076,N_1473);
or U1701 (N_1701,N_1482,N_1109);
nand U1702 (N_1702,N_1300,N_1051);
or U1703 (N_1703,N_1198,N_1222);
nor U1704 (N_1704,N_1091,N_1478);
nand U1705 (N_1705,N_1131,N_1146);
and U1706 (N_1706,N_1440,N_1488);
nor U1707 (N_1707,N_1435,N_1310);
nor U1708 (N_1708,N_1321,N_1020);
and U1709 (N_1709,N_1357,N_1097);
or U1710 (N_1710,N_1186,N_1215);
nor U1711 (N_1711,N_1095,N_1193);
xnor U1712 (N_1712,N_1284,N_1032);
and U1713 (N_1713,N_1370,N_1338);
nor U1714 (N_1714,N_1302,N_1341);
or U1715 (N_1715,N_1345,N_1018);
or U1716 (N_1716,N_1354,N_1385);
and U1717 (N_1717,N_1443,N_1434);
nor U1718 (N_1718,N_1377,N_1031);
and U1719 (N_1719,N_1393,N_1205);
or U1720 (N_1720,N_1245,N_1195);
or U1721 (N_1721,N_1288,N_1448);
nand U1722 (N_1722,N_1238,N_1353);
nand U1723 (N_1723,N_1152,N_1159);
nor U1724 (N_1724,N_1117,N_1124);
or U1725 (N_1725,N_1413,N_1048);
or U1726 (N_1726,N_1041,N_1212);
or U1727 (N_1727,N_1019,N_1158);
nand U1728 (N_1728,N_1207,N_1465);
and U1729 (N_1729,N_1219,N_1328);
and U1730 (N_1730,N_1279,N_1318);
nand U1731 (N_1731,N_1240,N_1011);
and U1732 (N_1732,N_1223,N_1316);
nor U1733 (N_1733,N_1461,N_1075);
or U1734 (N_1734,N_1084,N_1490);
nor U1735 (N_1735,N_1408,N_1217);
or U1736 (N_1736,N_1468,N_1281);
and U1737 (N_1737,N_1335,N_1162);
xor U1738 (N_1738,N_1438,N_1071);
or U1739 (N_1739,N_1083,N_1224);
and U1740 (N_1740,N_1008,N_1485);
nor U1741 (N_1741,N_1463,N_1258);
and U1742 (N_1742,N_1216,N_1174);
and U1743 (N_1743,N_1283,N_1181);
nor U1744 (N_1744,N_1445,N_1417);
nor U1745 (N_1745,N_1086,N_1122);
or U1746 (N_1746,N_1371,N_1116);
xnor U1747 (N_1747,N_1346,N_1177);
or U1748 (N_1748,N_1132,N_1311);
or U1749 (N_1749,N_1123,N_1295);
nand U1750 (N_1750,N_1394,N_1452);
or U1751 (N_1751,N_1340,N_1158);
nand U1752 (N_1752,N_1221,N_1405);
nand U1753 (N_1753,N_1486,N_1265);
or U1754 (N_1754,N_1174,N_1069);
nand U1755 (N_1755,N_1101,N_1052);
nor U1756 (N_1756,N_1207,N_1036);
or U1757 (N_1757,N_1284,N_1090);
nor U1758 (N_1758,N_1461,N_1258);
nor U1759 (N_1759,N_1217,N_1278);
or U1760 (N_1760,N_1066,N_1247);
or U1761 (N_1761,N_1480,N_1125);
nand U1762 (N_1762,N_1110,N_1245);
nor U1763 (N_1763,N_1309,N_1250);
or U1764 (N_1764,N_1454,N_1270);
xor U1765 (N_1765,N_1209,N_1131);
nor U1766 (N_1766,N_1350,N_1331);
or U1767 (N_1767,N_1252,N_1325);
or U1768 (N_1768,N_1096,N_1326);
nor U1769 (N_1769,N_1315,N_1366);
and U1770 (N_1770,N_1200,N_1348);
nand U1771 (N_1771,N_1117,N_1140);
and U1772 (N_1772,N_1471,N_1447);
or U1773 (N_1773,N_1281,N_1091);
or U1774 (N_1774,N_1062,N_1001);
nor U1775 (N_1775,N_1272,N_1328);
or U1776 (N_1776,N_1383,N_1175);
nor U1777 (N_1777,N_1153,N_1043);
and U1778 (N_1778,N_1044,N_1027);
or U1779 (N_1779,N_1079,N_1255);
and U1780 (N_1780,N_1043,N_1093);
nor U1781 (N_1781,N_1212,N_1321);
and U1782 (N_1782,N_1376,N_1349);
nor U1783 (N_1783,N_1039,N_1137);
and U1784 (N_1784,N_1076,N_1341);
or U1785 (N_1785,N_1325,N_1246);
and U1786 (N_1786,N_1175,N_1019);
nor U1787 (N_1787,N_1186,N_1101);
or U1788 (N_1788,N_1095,N_1285);
nand U1789 (N_1789,N_1358,N_1088);
nor U1790 (N_1790,N_1443,N_1051);
nand U1791 (N_1791,N_1338,N_1447);
or U1792 (N_1792,N_1394,N_1445);
nor U1793 (N_1793,N_1152,N_1118);
and U1794 (N_1794,N_1142,N_1316);
and U1795 (N_1795,N_1220,N_1303);
and U1796 (N_1796,N_1363,N_1322);
nand U1797 (N_1797,N_1310,N_1110);
nand U1798 (N_1798,N_1353,N_1395);
nor U1799 (N_1799,N_1381,N_1099);
and U1800 (N_1800,N_1034,N_1120);
and U1801 (N_1801,N_1495,N_1046);
and U1802 (N_1802,N_1094,N_1477);
and U1803 (N_1803,N_1462,N_1324);
or U1804 (N_1804,N_1399,N_1385);
nor U1805 (N_1805,N_1017,N_1280);
nand U1806 (N_1806,N_1115,N_1394);
and U1807 (N_1807,N_1274,N_1132);
nor U1808 (N_1808,N_1147,N_1126);
nor U1809 (N_1809,N_1332,N_1044);
or U1810 (N_1810,N_1222,N_1189);
nand U1811 (N_1811,N_1186,N_1230);
nor U1812 (N_1812,N_1363,N_1113);
or U1813 (N_1813,N_1236,N_1411);
or U1814 (N_1814,N_1020,N_1077);
nand U1815 (N_1815,N_1452,N_1310);
or U1816 (N_1816,N_1207,N_1458);
nand U1817 (N_1817,N_1031,N_1447);
or U1818 (N_1818,N_1210,N_1001);
nand U1819 (N_1819,N_1292,N_1228);
nor U1820 (N_1820,N_1075,N_1216);
nor U1821 (N_1821,N_1270,N_1212);
or U1822 (N_1822,N_1370,N_1058);
and U1823 (N_1823,N_1365,N_1299);
or U1824 (N_1824,N_1470,N_1071);
nand U1825 (N_1825,N_1174,N_1086);
nor U1826 (N_1826,N_1041,N_1152);
nor U1827 (N_1827,N_1029,N_1111);
and U1828 (N_1828,N_1078,N_1496);
or U1829 (N_1829,N_1119,N_1104);
and U1830 (N_1830,N_1190,N_1127);
nor U1831 (N_1831,N_1455,N_1180);
or U1832 (N_1832,N_1376,N_1302);
or U1833 (N_1833,N_1101,N_1292);
nand U1834 (N_1834,N_1387,N_1273);
and U1835 (N_1835,N_1140,N_1434);
nor U1836 (N_1836,N_1128,N_1293);
or U1837 (N_1837,N_1027,N_1337);
nor U1838 (N_1838,N_1088,N_1154);
and U1839 (N_1839,N_1340,N_1021);
nand U1840 (N_1840,N_1495,N_1344);
xnor U1841 (N_1841,N_1127,N_1139);
or U1842 (N_1842,N_1489,N_1447);
nand U1843 (N_1843,N_1444,N_1188);
nor U1844 (N_1844,N_1074,N_1409);
nor U1845 (N_1845,N_1196,N_1486);
and U1846 (N_1846,N_1499,N_1364);
or U1847 (N_1847,N_1389,N_1453);
nor U1848 (N_1848,N_1265,N_1068);
nand U1849 (N_1849,N_1223,N_1110);
nor U1850 (N_1850,N_1377,N_1408);
nor U1851 (N_1851,N_1226,N_1359);
and U1852 (N_1852,N_1380,N_1181);
and U1853 (N_1853,N_1229,N_1221);
and U1854 (N_1854,N_1227,N_1461);
or U1855 (N_1855,N_1053,N_1125);
nor U1856 (N_1856,N_1061,N_1009);
or U1857 (N_1857,N_1351,N_1488);
or U1858 (N_1858,N_1413,N_1448);
or U1859 (N_1859,N_1353,N_1025);
nand U1860 (N_1860,N_1450,N_1486);
nor U1861 (N_1861,N_1165,N_1344);
xnor U1862 (N_1862,N_1186,N_1053);
and U1863 (N_1863,N_1155,N_1485);
nand U1864 (N_1864,N_1265,N_1222);
nor U1865 (N_1865,N_1378,N_1056);
nor U1866 (N_1866,N_1315,N_1206);
nor U1867 (N_1867,N_1220,N_1240);
nand U1868 (N_1868,N_1184,N_1267);
or U1869 (N_1869,N_1465,N_1213);
nor U1870 (N_1870,N_1309,N_1116);
nand U1871 (N_1871,N_1470,N_1387);
and U1872 (N_1872,N_1408,N_1498);
or U1873 (N_1873,N_1147,N_1245);
nand U1874 (N_1874,N_1130,N_1023);
nand U1875 (N_1875,N_1336,N_1184);
nand U1876 (N_1876,N_1187,N_1252);
or U1877 (N_1877,N_1425,N_1079);
nor U1878 (N_1878,N_1067,N_1088);
or U1879 (N_1879,N_1176,N_1384);
nor U1880 (N_1880,N_1112,N_1062);
nor U1881 (N_1881,N_1040,N_1252);
nand U1882 (N_1882,N_1013,N_1164);
or U1883 (N_1883,N_1023,N_1208);
xor U1884 (N_1884,N_1125,N_1294);
nor U1885 (N_1885,N_1449,N_1156);
nor U1886 (N_1886,N_1093,N_1415);
and U1887 (N_1887,N_1057,N_1024);
and U1888 (N_1888,N_1306,N_1486);
or U1889 (N_1889,N_1012,N_1184);
nand U1890 (N_1890,N_1356,N_1123);
nor U1891 (N_1891,N_1362,N_1140);
nor U1892 (N_1892,N_1156,N_1414);
xnor U1893 (N_1893,N_1175,N_1088);
or U1894 (N_1894,N_1328,N_1139);
nor U1895 (N_1895,N_1229,N_1350);
nor U1896 (N_1896,N_1249,N_1271);
nor U1897 (N_1897,N_1432,N_1027);
and U1898 (N_1898,N_1240,N_1144);
nand U1899 (N_1899,N_1345,N_1136);
or U1900 (N_1900,N_1497,N_1122);
xor U1901 (N_1901,N_1431,N_1016);
nor U1902 (N_1902,N_1151,N_1033);
and U1903 (N_1903,N_1247,N_1268);
nor U1904 (N_1904,N_1007,N_1483);
nand U1905 (N_1905,N_1407,N_1069);
nand U1906 (N_1906,N_1291,N_1292);
nand U1907 (N_1907,N_1201,N_1448);
nor U1908 (N_1908,N_1302,N_1078);
or U1909 (N_1909,N_1493,N_1399);
nand U1910 (N_1910,N_1373,N_1486);
and U1911 (N_1911,N_1485,N_1295);
and U1912 (N_1912,N_1251,N_1271);
or U1913 (N_1913,N_1494,N_1474);
nor U1914 (N_1914,N_1110,N_1156);
nand U1915 (N_1915,N_1055,N_1394);
xor U1916 (N_1916,N_1235,N_1011);
xnor U1917 (N_1917,N_1180,N_1197);
and U1918 (N_1918,N_1007,N_1282);
nor U1919 (N_1919,N_1027,N_1263);
nor U1920 (N_1920,N_1194,N_1046);
nor U1921 (N_1921,N_1425,N_1376);
or U1922 (N_1922,N_1227,N_1213);
and U1923 (N_1923,N_1288,N_1032);
nand U1924 (N_1924,N_1023,N_1030);
and U1925 (N_1925,N_1287,N_1367);
nor U1926 (N_1926,N_1268,N_1197);
or U1927 (N_1927,N_1377,N_1393);
nand U1928 (N_1928,N_1105,N_1310);
nor U1929 (N_1929,N_1075,N_1128);
nand U1930 (N_1930,N_1105,N_1338);
and U1931 (N_1931,N_1393,N_1358);
and U1932 (N_1932,N_1388,N_1092);
nand U1933 (N_1933,N_1300,N_1254);
xnor U1934 (N_1934,N_1099,N_1159);
nand U1935 (N_1935,N_1046,N_1280);
nand U1936 (N_1936,N_1051,N_1456);
nor U1937 (N_1937,N_1014,N_1325);
and U1938 (N_1938,N_1060,N_1021);
nand U1939 (N_1939,N_1265,N_1246);
or U1940 (N_1940,N_1371,N_1283);
nor U1941 (N_1941,N_1051,N_1220);
and U1942 (N_1942,N_1210,N_1002);
and U1943 (N_1943,N_1478,N_1211);
or U1944 (N_1944,N_1406,N_1284);
nand U1945 (N_1945,N_1262,N_1384);
nand U1946 (N_1946,N_1295,N_1362);
and U1947 (N_1947,N_1307,N_1279);
or U1948 (N_1948,N_1124,N_1350);
or U1949 (N_1949,N_1314,N_1416);
nand U1950 (N_1950,N_1114,N_1291);
and U1951 (N_1951,N_1032,N_1177);
and U1952 (N_1952,N_1398,N_1476);
xnor U1953 (N_1953,N_1034,N_1032);
or U1954 (N_1954,N_1030,N_1311);
or U1955 (N_1955,N_1079,N_1006);
nand U1956 (N_1956,N_1059,N_1045);
nand U1957 (N_1957,N_1492,N_1395);
and U1958 (N_1958,N_1335,N_1374);
nor U1959 (N_1959,N_1221,N_1456);
nand U1960 (N_1960,N_1007,N_1168);
nor U1961 (N_1961,N_1135,N_1499);
nor U1962 (N_1962,N_1277,N_1003);
and U1963 (N_1963,N_1267,N_1122);
nand U1964 (N_1964,N_1485,N_1373);
nand U1965 (N_1965,N_1261,N_1197);
or U1966 (N_1966,N_1041,N_1497);
and U1967 (N_1967,N_1464,N_1238);
nand U1968 (N_1968,N_1131,N_1161);
nor U1969 (N_1969,N_1472,N_1248);
nor U1970 (N_1970,N_1048,N_1460);
nor U1971 (N_1971,N_1096,N_1026);
or U1972 (N_1972,N_1220,N_1115);
nand U1973 (N_1973,N_1119,N_1404);
xnor U1974 (N_1974,N_1001,N_1381);
or U1975 (N_1975,N_1116,N_1263);
nor U1976 (N_1976,N_1184,N_1153);
or U1977 (N_1977,N_1129,N_1017);
nand U1978 (N_1978,N_1334,N_1038);
or U1979 (N_1979,N_1198,N_1165);
or U1980 (N_1980,N_1399,N_1325);
and U1981 (N_1981,N_1020,N_1147);
or U1982 (N_1982,N_1378,N_1108);
or U1983 (N_1983,N_1421,N_1317);
nand U1984 (N_1984,N_1438,N_1492);
and U1985 (N_1985,N_1188,N_1202);
or U1986 (N_1986,N_1121,N_1486);
nor U1987 (N_1987,N_1034,N_1310);
nor U1988 (N_1988,N_1118,N_1261);
or U1989 (N_1989,N_1135,N_1433);
or U1990 (N_1990,N_1030,N_1105);
or U1991 (N_1991,N_1092,N_1275);
and U1992 (N_1992,N_1228,N_1474);
or U1993 (N_1993,N_1441,N_1490);
nor U1994 (N_1994,N_1359,N_1445);
or U1995 (N_1995,N_1270,N_1245);
or U1996 (N_1996,N_1427,N_1073);
or U1997 (N_1997,N_1453,N_1034);
xor U1998 (N_1998,N_1493,N_1122);
nand U1999 (N_1999,N_1208,N_1120);
or U2000 (N_2000,N_1802,N_1864);
and U2001 (N_2001,N_1774,N_1665);
xor U2002 (N_2002,N_1571,N_1626);
nand U2003 (N_2003,N_1737,N_1575);
nor U2004 (N_2004,N_1557,N_1916);
xnor U2005 (N_2005,N_1506,N_1963);
and U2006 (N_2006,N_1943,N_1886);
nand U2007 (N_2007,N_1788,N_1949);
and U2008 (N_2008,N_1736,N_1545);
or U2009 (N_2009,N_1647,N_1507);
nor U2010 (N_2010,N_1751,N_1784);
nor U2011 (N_2011,N_1925,N_1778);
or U2012 (N_2012,N_1746,N_1681);
and U2013 (N_2013,N_1556,N_1903);
nor U2014 (N_2014,N_1710,N_1898);
nand U2015 (N_2015,N_1542,N_1798);
or U2016 (N_2016,N_1599,N_1603);
nor U2017 (N_2017,N_1514,N_1550);
nor U2018 (N_2018,N_1581,N_1801);
nor U2019 (N_2019,N_1752,N_1857);
and U2020 (N_2020,N_1919,N_1837);
nor U2021 (N_2021,N_1513,N_1867);
nor U2022 (N_2022,N_1560,N_1779);
or U2023 (N_2023,N_1823,N_1555);
or U2024 (N_2024,N_1716,N_1725);
or U2025 (N_2025,N_1985,N_1667);
and U2026 (N_2026,N_1965,N_1954);
nand U2027 (N_2027,N_1720,N_1889);
nand U2028 (N_2028,N_1905,N_1794);
nand U2029 (N_2029,N_1793,N_1882);
and U2030 (N_2030,N_1564,N_1825);
or U2031 (N_2031,N_1861,N_1990);
nand U2032 (N_2032,N_1782,N_1643);
nand U2033 (N_2033,N_1610,N_1912);
or U2034 (N_2034,N_1628,N_1944);
nand U2035 (N_2035,N_1713,N_1785);
nor U2036 (N_2036,N_1754,N_1934);
or U2037 (N_2037,N_1644,N_1553);
nand U2038 (N_2038,N_1589,N_1894);
nand U2039 (N_2039,N_1924,N_1881);
or U2040 (N_2040,N_1639,N_1698);
nand U2041 (N_2041,N_1563,N_1900);
and U2042 (N_2042,N_1756,N_1906);
nor U2043 (N_2043,N_1762,N_1691);
or U2044 (N_2044,N_1776,N_1760);
or U2045 (N_2045,N_1680,N_1645);
or U2046 (N_2046,N_1629,N_1917);
and U2047 (N_2047,N_1868,N_1614);
nand U2048 (N_2048,N_1574,N_1789);
nor U2049 (N_2049,N_1841,N_1638);
nand U2050 (N_2050,N_1862,N_1849);
and U2051 (N_2051,N_1674,N_1950);
or U2052 (N_2052,N_1997,N_1694);
or U2053 (N_2053,N_1512,N_1528);
xnor U2054 (N_2054,N_1933,N_1792);
or U2055 (N_2055,N_1980,N_1959);
and U2056 (N_2056,N_1878,N_1601);
or U2057 (N_2057,N_1559,N_1761);
or U2058 (N_2058,N_1937,N_1783);
nand U2059 (N_2059,N_1981,N_1987);
nor U2060 (N_2060,N_1809,N_1717);
nor U2061 (N_2061,N_1598,N_1953);
xor U2062 (N_2062,N_1757,N_1800);
or U2063 (N_2063,N_1653,N_1973);
or U2064 (N_2064,N_1524,N_1755);
nor U2065 (N_2065,N_1986,N_1781);
nor U2066 (N_2066,N_1676,N_1873);
nor U2067 (N_2067,N_1901,N_1697);
nand U2068 (N_2068,N_1657,N_1613);
or U2069 (N_2069,N_1687,N_1768);
nor U2070 (N_2070,N_1734,N_1650);
or U2071 (N_2071,N_1729,N_1991);
nand U2072 (N_2072,N_1835,N_1731);
nand U2073 (N_2073,N_1578,N_1688);
nand U2074 (N_2074,N_1926,N_1711);
and U2075 (N_2075,N_1723,N_1714);
nand U2076 (N_2076,N_1604,N_1646);
nand U2077 (N_2077,N_1743,N_1870);
nand U2078 (N_2078,N_1602,N_1952);
nor U2079 (N_2079,N_1904,N_1791);
nand U2080 (N_2080,N_1846,N_1840);
or U2081 (N_2081,N_1938,N_1732);
and U2082 (N_2082,N_1652,N_1527);
and U2083 (N_2083,N_1592,N_1709);
or U2084 (N_2084,N_1551,N_1648);
nand U2085 (N_2085,N_1741,N_1693);
or U2086 (N_2086,N_1617,N_1682);
or U2087 (N_2087,N_1967,N_1576);
or U2088 (N_2088,N_1523,N_1582);
nand U2089 (N_2089,N_1964,N_1655);
or U2090 (N_2090,N_1941,N_1955);
and U2091 (N_2091,N_1505,N_1567);
or U2092 (N_2092,N_1615,N_1662);
nor U2093 (N_2093,N_1910,N_1600);
nor U2094 (N_2094,N_1561,N_1642);
nand U2095 (N_2095,N_1974,N_1594);
nor U2096 (N_2096,N_1871,N_1875);
nor U2097 (N_2097,N_1773,N_1994);
nand U2098 (N_2098,N_1689,N_1738);
or U2099 (N_2099,N_1702,N_1529);
and U2100 (N_2100,N_1942,N_1771);
or U2101 (N_2101,N_1570,N_1921);
nor U2102 (N_2102,N_1803,N_1817);
nand U2103 (N_2103,N_1516,N_1855);
nor U2104 (N_2104,N_1962,N_1992);
nor U2105 (N_2105,N_1543,N_1908);
and U2106 (N_2106,N_1821,N_1532);
and U2107 (N_2107,N_1659,N_1863);
nor U2108 (N_2108,N_1632,N_1651);
or U2109 (N_2109,N_1805,N_1956);
or U2110 (N_2110,N_1663,N_1748);
nor U2111 (N_2111,N_1673,N_1923);
and U2112 (N_2112,N_1876,N_1562);
and U2113 (N_2113,N_1945,N_1995);
nand U2114 (N_2114,N_1568,N_1565);
and U2115 (N_2115,N_1931,N_1830);
or U2116 (N_2116,N_1728,N_1775);
nor U2117 (N_2117,N_1669,N_1631);
nor U2118 (N_2118,N_1984,N_1971);
nand U2119 (N_2119,N_1726,N_1538);
nor U2120 (N_2120,N_1854,N_1847);
nand U2121 (N_2121,N_1597,N_1544);
nand U2122 (N_2122,N_1972,N_1699);
or U2123 (N_2123,N_1636,N_1929);
nand U2124 (N_2124,N_1939,N_1704);
nand U2125 (N_2125,N_1504,N_1998);
nor U2126 (N_2126,N_1832,N_1612);
or U2127 (N_2127,N_1895,N_1838);
or U2128 (N_2128,N_1558,N_1874);
nand U2129 (N_2129,N_1843,N_1885);
nor U2130 (N_2130,N_1811,N_1915);
or U2131 (N_2131,N_1546,N_1526);
nand U2132 (N_2132,N_1552,N_1660);
nor U2133 (N_2133,N_1946,N_1742);
or U2134 (N_2134,N_1625,N_1958);
nand U2135 (N_2135,N_1880,N_1796);
xnor U2136 (N_2136,N_1727,N_1595);
nor U2137 (N_2137,N_1521,N_1596);
nor U2138 (N_2138,N_1797,N_1979);
nor U2139 (N_2139,N_1786,N_1914);
and U2140 (N_2140,N_1573,N_1707);
or U2141 (N_2141,N_1858,N_1848);
or U2142 (N_2142,N_1820,N_1606);
nand U2143 (N_2143,N_1899,N_1583);
nand U2144 (N_2144,N_1718,N_1739);
and U2145 (N_2145,N_1591,N_1547);
nand U2146 (N_2146,N_1509,N_1672);
nor U2147 (N_2147,N_1675,N_1866);
nor U2148 (N_2148,N_1759,N_1819);
nand U2149 (N_2149,N_1807,N_1519);
nor U2150 (N_2150,N_1508,N_1763);
nor U2151 (N_2151,N_1684,N_1670);
nor U2152 (N_2152,N_1608,N_1501);
or U2153 (N_2153,N_1982,N_1750);
nor U2154 (N_2154,N_1988,N_1593);
nand U2155 (N_2155,N_1622,N_1940);
and U2156 (N_2156,N_1585,N_1500);
nor U2157 (N_2157,N_1948,N_1587);
nor U2158 (N_2158,N_1812,N_1968);
nand U2159 (N_2159,N_1664,N_1765);
nor U2160 (N_2160,N_1865,N_1749);
and U2161 (N_2161,N_1810,N_1892);
nor U2162 (N_2162,N_1896,N_1656);
and U2163 (N_2163,N_1911,N_1996);
xor U2164 (N_2164,N_1511,N_1836);
or U2165 (N_2165,N_1586,N_1531);
or U2166 (N_2166,N_1851,N_1619);
or U2167 (N_2167,N_1719,N_1588);
and U2168 (N_2168,N_1683,N_1666);
nand U2169 (N_2169,N_1554,N_1533);
xor U2170 (N_2170,N_1883,N_1927);
and U2171 (N_2171,N_1745,N_1951);
nand U2172 (N_2172,N_1961,N_1834);
and U2173 (N_2173,N_1620,N_1517);
or U2174 (N_2174,N_1829,N_1549);
or U2175 (N_2175,N_1671,N_1658);
nor U2176 (N_2176,N_1913,N_1520);
nor U2177 (N_2177,N_1999,N_1540);
xor U2178 (N_2178,N_1695,N_1884);
or U2179 (N_2179,N_1686,N_1537);
or U2180 (N_2180,N_1887,N_1787);
or U2181 (N_2181,N_1534,N_1701);
nand U2182 (N_2182,N_1891,N_1569);
and U2183 (N_2183,N_1641,N_1983);
nor U2184 (N_2184,N_1877,N_1806);
xor U2185 (N_2185,N_1654,N_1907);
or U2186 (N_2186,N_1541,N_1932);
nand U2187 (N_2187,N_1502,N_1777);
nor U2188 (N_2188,N_1957,N_1535);
and U2189 (N_2189,N_1808,N_1989);
and U2190 (N_2190,N_1795,N_1634);
and U2191 (N_2191,N_1715,N_1577);
or U2192 (N_2192,N_1692,N_1518);
or U2193 (N_2193,N_1930,N_1758);
nand U2194 (N_2194,N_1767,N_1966);
nor U2195 (N_2195,N_1975,N_1548);
and U2196 (N_2196,N_1890,N_1678);
nand U2197 (N_2197,N_1539,N_1850);
and U2198 (N_2198,N_1839,N_1920);
nor U2199 (N_2199,N_1580,N_1708);
nand U2200 (N_2200,N_1833,N_1824);
nand U2201 (N_2201,N_1813,N_1814);
and U2202 (N_2202,N_1928,N_1633);
nand U2203 (N_2203,N_1515,N_1902);
and U2204 (N_2204,N_1844,N_1605);
nand U2205 (N_2205,N_1978,N_1584);
nand U2206 (N_2206,N_1909,N_1690);
or U2207 (N_2207,N_1769,N_1872);
and U2208 (N_2208,N_1503,N_1572);
and U2209 (N_2209,N_1827,N_1856);
nor U2210 (N_2210,N_1730,N_1816);
nor U2211 (N_2211,N_1828,N_1918);
or U2212 (N_2212,N_1790,N_1799);
nand U2213 (N_2213,N_1936,N_1935);
nor U2214 (N_2214,N_1640,N_1818);
nor U2215 (N_2215,N_1826,N_1609);
nor U2216 (N_2216,N_1530,N_1772);
or U2217 (N_2217,N_1627,N_1740);
nor U2218 (N_2218,N_1522,N_1611);
nor U2219 (N_2219,N_1616,N_1635);
and U2220 (N_2220,N_1747,N_1770);
or U2221 (N_2221,N_1621,N_1637);
or U2222 (N_2222,N_1510,N_1859);
and U2223 (N_2223,N_1744,N_1618);
nor U2224 (N_2224,N_1976,N_1735);
nor U2225 (N_2225,N_1815,N_1893);
or U2226 (N_2226,N_1525,N_1753);
nor U2227 (N_2227,N_1721,N_1852);
or U2228 (N_2228,N_1842,N_1685);
nor U2229 (N_2229,N_1977,N_1970);
or U2230 (N_2230,N_1649,N_1993);
nor U2231 (N_2231,N_1706,N_1853);
and U2232 (N_2232,N_1579,N_1624);
nor U2233 (N_2233,N_1764,N_1879);
xor U2234 (N_2234,N_1679,N_1566);
nor U2235 (N_2235,N_1888,N_1960);
or U2236 (N_2236,N_1668,N_1831);
nand U2237 (N_2237,N_1677,N_1804);
and U2238 (N_2238,N_1700,N_1630);
or U2239 (N_2239,N_1703,N_1623);
or U2240 (N_2240,N_1922,N_1780);
and U2241 (N_2241,N_1860,N_1969);
nor U2242 (N_2242,N_1822,N_1766);
or U2243 (N_2243,N_1590,N_1712);
or U2244 (N_2244,N_1845,N_1705);
and U2245 (N_2245,N_1722,N_1536);
or U2246 (N_2246,N_1897,N_1947);
and U2247 (N_2247,N_1661,N_1724);
or U2248 (N_2248,N_1607,N_1869);
and U2249 (N_2249,N_1733,N_1696);
or U2250 (N_2250,N_1934,N_1693);
nor U2251 (N_2251,N_1876,N_1611);
nand U2252 (N_2252,N_1830,N_1982);
nand U2253 (N_2253,N_1669,N_1791);
nand U2254 (N_2254,N_1562,N_1846);
and U2255 (N_2255,N_1771,N_1635);
or U2256 (N_2256,N_1687,N_1533);
nor U2257 (N_2257,N_1501,N_1536);
and U2258 (N_2258,N_1502,N_1641);
nand U2259 (N_2259,N_1949,N_1593);
nor U2260 (N_2260,N_1629,N_1963);
and U2261 (N_2261,N_1775,N_1617);
nor U2262 (N_2262,N_1825,N_1738);
nand U2263 (N_2263,N_1547,N_1777);
nor U2264 (N_2264,N_1934,N_1774);
nand U2265 (N_2265,N_1767,N_1926);
or U2266 (N_2266,N_1890,N_1832);
nor U2267 (N_2267,N_1675,N_1692);
xor U2268 (N_2268,N_1676,N_1707);
and U2269 (N_2269,N_1564,N_1710);
and U2270 (N_2270,N_1556,N_1896);
and U2271 (N_2271,N_1792,N_1630);
and U2272 (N_2272,N_1511,N_1601);
and U2273 (N_2273,N_1913,N_1548);
nand U2274 (N_2274,N_1617,N_1846);
and U2275 (N_2275,N_1513,N_1922);
nand U2276 (N_2276,N_1607,N_1851);
or U2277 (N_2277,N_1935,N_1861);
nand U2278 (N_2278,N_1581,N_1961);
nor U2279 (N_2279,N_1626,N_1838);
and U2280 (N_2280,N_1597,N_1981);
and U2281 (N_2281,N_1954,N_1677);
nor U2282 (N_2282,N_1907,N_1890);
nor U2283 (N_2283,N_1972,N_1765);
nand U2284 (N_2284,N_1874,N_1603);
nand U2285 (N_2285,N_1754,N_1504);
or U2286 (N_2286,N_1561,N_1692);
or U2287 (N_2287,N_1506,N_1955);
nand U2288 (N_2288,N_1650,N_1788);
nand U2289 (N_2289,N_1815,N_1776);
nor U2290 (N_2290,N_1966,N_1522);
nor U2291 (N_2291,N_1943,N_1652);
or U2292 (N_2292,N_1865,N_1897);
or U2293 (N_2293,N_1777,N_1601);
or U2294 (N_2294,N_1883,N_1664);
nand U2295 (N_2295,N_1816,N_1616);
nand U2296 (N_2296,N_1887,N_1637);
or U2297 (N_2297,N_1742,N_1975);
nor U2298 (N_2298,N_1794,N_1500);
nor U2299 (N_2299,N_1756,N_1992);
or U2300 (N_2300,N_1994,N_1785);
and U2301 (N_2301,N_1785,N_1526);
nor U2302 (N_2302,N_1703,N_1699);
or U2303 (N_2303,N_1694,N_1857);
and U2304 (N_2304,N_1745,N_1678);
or U2305 (N_2305,N_1862,N_1656);
nor U2306 (N_2306,N_1501,N_1663);
or U2307 (N_2307,N_1994,N_1749);
or U2308 (N_2308,N_1508,N_1597);
or U2309 (N_2309,N_1976,N_1612);
and U2310 (N_2310,N_1617,N_1821);
nor U2311 (N_2311,N_1530,N_1653);
nand U2312 (N_2312,N_1730,N_1796);
or U2313 (N_2313,N_1969,N_1919);
and U2314 (N_2314,N_1846,N_1943);
and U2315 (N_2315,N_1701,N_1945);
or U2316 (N_2316,N_1743,N_1971);
nand U2317 (N_2317,N_1773,N_1714);
nor U2318 (N_2318,N_1985,N_1977);
and U2319 (N_2319,N_1663,N_1691);
or U2320 (N_2320,N_1565,N_1955);
and U2321 (N_2321,N_1675,N_1820);
and U2322 (N_2322,N_1908,N_1993);
nand U2323 (N_2323,N_1666,N_1999);
or U2324 (N_2324,N_1931,N_1894);
or U2325 (N_2325,N_1608,N_1973);
or U2326 (N_2326,N_1899,N_1917);
or U2327 (N_2327,N_1722,N_1660);
nor U2328 (N_2328,N_1896,N_1694);
or U2329 (N_2329,N_1745,N_1756);
or U2330 (N_2330,N_1501,N_1975);
nand U2331 (N_2331,N_1564,N_1647);
nor U2332 (N_2332,N_1531,N_1917);
and U2333 (N_2333,N_1616,N_1550);
nand U2334 (N_2334,N_1713,N_1545);
nand U2335 (N_2335,N_1875,N_1553);
nor U2336 (N_2336,N_1962,N_1923);
nand U2337 (N_2337,N_1587,N_1711);
nand U2338 (N_2338,N_1519,N_1640);
nand U2339 (N_2339,N_1539,N_1779);
or U2340 (N_2340,N_1789,N_1918);
and U2341 (N_2341,N_1789,N_1867);
or U2342 (N_2342,N_1835,N_1628);
nor U2343 (N_2343,N_1839,N_1637);
nand U2344 (N_2344,N_1669,N_1841);
and U2345 (N_2345,N_1740,N_1917);
and U2346 (N_2346,N_1547,N_1687);
nand U2347 (N_2347,N_1566,N_1538);
or U2348 (N_2348,N_1918,N_1601);
or U2349 (N_2349,N_1704,N_1722);
and U2350 (N_2350,N_1958,N_1817);
nand U2351 (N_2351,N_1511,N_1937);
nand U2352 (N_2352,N_1713,N_1575);
or U2353 (N_2353,N_1617,N_1899);
and U2354 (N_2354,N_1987,N_1651);
nand U2355 (N_2355,N_1674,N_1980);
and U2356 (N_2356,N_1900,N_1513);
and U2357 (N_2357,N_1756,N_1583);
or U2358 (N_2358,N_1901,N_1808);
and U2359 (N_2359,N_1903,N_1747);
nand U2360 (N_2360,N_1727,N_1954);
and U2361 (N_2361,N_1546,N_1816);
nor U2362 (N_2362,N_1926,N_1999);
nand U2363 (N_2363,N_1994,N_1860);
and U2364 (N_2364,N_1643,N_1548);
nor U2365 (N_2365,N_1753,N_1727);
or U2366 (N_2366,N_1528,N_1896);
and U2367 (N_2367,N_1597,N_1657);
nand U2368 (N_2368,N_1844,N_1994);
and U2369 (N_2369,N_1566,N_1874);
nor U2370 (N_2370,N_1877,N_1755);
nand U2371 (N_2371,N_1530,N_1860);
or U2372 (N_2372,N_1668,N_1579);
or U2373 (N_2373,N_1818,N_1853);
or U2374 (N_2374,N_1608,N_1510);
or U2375 (N_2375,N_1588,N_1700);
nor U2376 (N_2376,N_1950,N_1743);
or U2377 (N_2377,N_1699,N_1725);
nand U2378 (N_2378,N_1665,N_1808);
and U2379 (N_2379,N_1838,N_1888);
nor U2380 (N_2380,N_1895,N_1582);
nor U2381 (N_2381,N_1689,N_1598);
xnor U2382 (N_2382,N_1777,N_1676);
and U2383 (N_2383,N_1649,N_1629);
and U2384 (N_2384,N_1516,N_1554);
nor U2385 (N_2385,N_1701,N_1540);
nand U2386 (N_2386,N_1963,N_1518);
or U2387 (N_2387,N_1859,N_1927);
and U2388 (N_2388,N_1694,N_1529);
nand U2389 (N_2389,N_1604,N_1580);
nor U2390 (N_2390,N_1713,N_1555);
or U2391 (N_2391,N_1534,N_1590);
or U2392 (N_2392,N_1782,N_1628);
or U2393 (N_2393,N_1734,N_1513);
nor U2394 (N_2394,N_1734,N_1626);
nor U2395 (N_2395,N_1976,N_1977);
nor U2396 (N_2396,N_1702,N_1897);
xor U2397 (N_2397,N_1554,N_1913);
nor U2398 (N_2398,N_1644,N_1609);
or U2399 (N_2399,N_1887,N_1960);
nand U2400 (N_2400,N_1788,N_1569);
nor U2401 (N_2401,N_1765,N_1788);
nand U2402 (N_2402,N_1908,N_1642);
nor U2403 (N_2403,N_1906,N_1861);
nor U2404 (N_2404,N_1840,N_1627);
or U2405 (N_2405,N_1825,N_1965);
nand U2406 (N_2406,N_1825,N_1671);
nand U2407 (N_2407,N_1524,N_1965);
and U2408 (N_2408,N_1684,N_1950);
nand U2409 (N_2409,N_1925,N_1856);
nand U2410 (N_2410,N_1874,N_1792);
and U2411 (N_2411,N_1845,N_1821);
and U2412 (N_2412,N_1976,N_1573);
and U2413 (N_2413,N_1553,N_1904);
or U2414 (N_2414,N_1809,N_1774);
and U2415 (N_2415,N_1959,N_1977);
nor U2416 (N_2416,N_1868,N_1696);
nor U2417 (N_2417,N_1663,N_1758);
or U2418 (N_2418,N_1996,N_1573);
or U2419 (N_2419,N_1966,N_1691);
or U2420 (N_2420,N_1655,N_1829);
or U2421 (N_2421,N_1603,N_1742);
nor U2422 (N_2422,N_1965,N_1898);
nor U2423 (N_2423,N_1698,N_1593);
or U2424 (N_2424,N_1980,N_1871);
or U2425 (N_2425,N_1720,N_1630);
nor U2426 (N_2426,N_1906,N_1645);
nand U2427 (N_2427,N_1603,N_1735);
nand U2428 (N_2428,N_1588,N_1907);
or U2429 (N_2429,N_1891,N_1521);
or U2430 (N_2430,N_1607,N_1780);
nor U2431 (N_2431,N_1974,N_1605);
nand U2432 (N_2432,N_1541,N_1563);
nand U2433 (N_2433,N_1833,N_1815);
nand U2434 (N_2434,N_1795,N_1681);
and U2435 (N_2435,N_1652,N_1900);
nand U2436 (N_2436,N_1883,N_1660);
and U2437 (N_2437,N_1708,N_1884);
nor U2438 (N_2438,N_1826,N_1578);
nand U2439 (N_2439,N_1663,N_1909);
or U2440 (N_2440,N_1767,N_1657);
or U2441 (N_2441,N_1906,N_1847);
and U2442 (N_2442,N_1982,N_1951);
and U2443 (N_2443,N_1524,N_1523);
or U2444 (N_2444,N_1612,N_1682);
nand U2445 (N_2445,N_1549,N_1556);
nand U2446 (N_2446,N_1732,N_1935);
nand U2447 (N_2447,N_1870,N_1758);
nor U2448 (N_2448,N_1586,N_1603);
nor U2449 (N_2449,N_1535,N_1611);
and U2450 (N_2450,N_1963,N_1665);
nand U2451 (N_2451,N_1782,N_1766);
and U2452 (N_2452,N_1579,N_1933);
and U2453 (N_2453,N_1653,N_1638);
nand U2454 (N_2454,N_1821,N_1691);
or U2455 (N_2455,N_1526,N_1551);
or U2456 (N_2456,N_1537,N_1983);
nor U2457 (N_2457,N_1652,N_1956);
nor U2458 (N_2458,N_1578,N_1836);
nand U2459 (N_2459,N_1735,N_1801);
nand U2460 (N_2460,N_1819,N_1604);
nor U2461 (N_2461,N_1674,N_1941);
and U2462 (N_2462,N_1932,N_1766);
nor U2463 (N_2463,N_1986,N_1663);
nor U2464 (N_2464,N_1571,N_1703);
and U2465 (N_2465,N_1988,N_1817);
or U2466 (N_2466,N_1706,N_1515);
and U2467 (N_2467,N_1994,N_1869);
nand U2468 (N_2468,N_1636,N_1815);
nand U2469 (N_2469,N_1888,N_1638);
or U2470 (N_2470,N_1605,N_1828);
and U2471 (N_2471,N_1769,N_1932);
or U2472 (N_2472,N_1921,N_1753);
nand U2473 (N_2473,N_1648,N_1755);
or U2474 (N_2474,N_1588,N_1735);
nand U2475 (N_2475,N_1635,N_1567);
or U2476 (N_2476,N_1799,N_1842);
or U2477 (N_2477,N_1527,N_1896);
or U2478 (N_2478,N_1660,N_1863);
and U2479 (N_2479,N_1952,N_1806);
nor U2480 (N_2480,N_1914,N_1845);
or U2481 (N_2481,N_1887,N_1750);
or U2482 (N_2482,N_1683,N_1543);
and U2483 (N_2483,N_1765,N_1775);
nor U2484 (N_2484,N_1873,N_1944);
or U2485 (N_2485,N_1824,N_1902);
nor U2486 (N_2486,N_1802,N_1584);
nand U2487 (N_2487,N_1661,N_1557);
or U2488 (N_2488,N_1559,N_1635);
or U2489 (N_2489,N_1860,N_1991);
and U2490 (N_2490,N_1850,N_1603);
nand U2491 (N_2491,N_1971,N_1604);
nor U2492 (N_2492,N_1508,N_1537);
or U2493 (N_2493,N_1638,N_1854);
nor U2494 (N_2494,N_1711,N_1659);
nand U2495 (N_2495,N_1670,N_1647);
and U2496 (N_2496,N_1753,N_1943);
and U2497 (N_2497,N_1829,N_1764);
nand U2498 (N_2498,N_1999,N_1648);
nor U2499 (N_2499,N_1558,N_1660);
nand U2500 (N_2500,N_2416,N_2106);
or U2501 (N_2501,N_2198,N_2456);
nor U2502 (N_2502,N_2023,N_2495);
nand U2503 (N_2503,N_2381,N_2287);
nand U2504 (N_2504,N_2107,N_2441);
and U2505 (N_2505,N_2015,N_2183);
or U2506 (N_2506,N_2174,N_2068);
or U2507 (N_2507,N_2387,N_2135);
or U2508 (N_2508,N_2476,N_2278);
nand U2509 (N_2509,N_2342,N_2446);
or U2510 (N_2510,N_2409,N_2449);
or U2511 (N_2511,N_2271,N_2269);
xnor U2512 (N_2512,N_2181,N_2266);
or U2513 (N_2513,N_2199,N_2100);
nand U2514 (N_2514,N_2038,N_2352);
nor U2515 (N_2515,N_2338,N_2263);
nand U2516 (N_2516,N_2036,N_2248);
nand U2517 (N_2517,N_2472,N_2072);
nand U2518 (N_2518,N_2480,N_2176);
or U2519 (N_2519,N_2325,N_2267);
or U2520 (N_2520,N_2259,N_2244);
or U2521 (N_2521,N_2185,N_2273);
xor U2522 (N_2522,N_2048,N_2317);
and U2523 (N_2523,N_2327,N_2356);
nor U2524 (N_2524,N_2272,N_2345);
and U2525 (N_2525,N_2066,N_2047);
nor U2526 (N_2526,N_2464,N_2247);
or U2527 (N_2527,N_2497,N_2055);
nor U2528 (N_2528,N_2237,N_2331);
nor U2529 (N_2529,N_2217,N_2291);
nand U2530 (N_2530,N_2286,N_2056);
nor U2531 (N_2531,N_2258,N_2438);
or U2532 (N_2532,N_2080,N_2367);
nor U2533 (N_2533,N_2488,N_2492);
or U2534 (N_2534,N_2444,N_2348);
nand U2535 (N_2535,N_2193,N_2284);
or U2536 (N_2536,N_2301,N_2486);
and U2537 (N_2537,N_2122,N_2282);
nand U2538 (N_2538,N_2389,N_2393);
or U2539 (N_2539,N_2123,N_2324);
or U2540 (N_2540,N_2159,N_2336);
nand U2541 (N_2541,N_2167,N_2128);
or U2542 (N_2542,N_2470,N_2017);
nor U2543 (N_2543,N_2354,N_2116);
or U2544 (N_2544,N_2083,N_2070);
nor U2545 (N_2545,N_2414,N_2455);
and U2546 (N_2546,N_2388,N_2028);
and U2547 (N_2547,N_2355,N_2081);
nor U2548 (N_2548,N_2090,N_2188);
and U2549 (N_2549,N_2344,N_2140);
or U2550 (N_2550,N_2264,N_2009);
nor U2551 (N_2551,N_2417,N_2133);
nand U2552 (N_2552,N_2316,N_2157);
and U2553 (N_2553,N_2137,N_2408);
or U2554 (N_2554,N_2311,N_2323);
or U2555 (N_2555,N_2042,N_2429);
and U2556 (N_2556,N_2005,N_2152);
or U2557 (N_2557,N_2415,N_2380);
nor U2558 (N_2558,N_2182,N_2216);
or U2559 (N_2559,N_2213,N_2277);
nand U2560 (N_2560,N_2363,N_2347);
and U2561 (N_2561,N_2466,N_2379);
and U2562 (N_2562,N_2397,N_2018);
or U2563 (N_2563,N_2184,N_2255);
nor U2564 (N_2564,N_2093,N_2427);
nand U2565 (N_2565,N_2453,N_2377);
or U2566 (N_2566,N_2307,N_2224);
and U2567 (N_2567,N_2296,N_2173);
nor U2568 (N_2568,N_2297,N_2111);
or U2569 (N_2569,N_2205,N_2396);
and U2570 (N_2570,N_2462,N_2463);
nor U2571 (N_2571,N_2221,N_2447);
and U2572 (N_2572,N_2285,N_2095);
and U2573 (N_2573,N_2346,N_2067);
nand U2574 (N_2574,N_2499,N_2156);
nand U2575 (N_2575,N_2308,N_2238);
and U2576 (N_2576,N_2321,N_2003);
or U2577 (N_2577,N_2059,N_2141);
or U2578 (N_2578,N_2457,N_2276);
and U2579 (N_2579,N_2050,N_2434);
or U2580 (N_2580,N_2143,N_2027);
and U2581 (N_2581,N_2451,N_2092);
nand U2582 (N_2582,N_2359,N_2085);
and U2583 (N_2583,N_2436,N_2306);
nand U2584 (N_2584,N_2114,N_2404);
nor U2585 (N_2585,N_2175,N_2362);
or U2586 (N_2586,N_2021,N_2121);
nor U2587 (N_2587,N_2011,N_2353);
and U2588 (N_2588,N_2340,N_2177);
or U2589 (N_2589,N_2274,N_2283);
nor U2590 (N_2590,N_2394,N_2033);
xnor U2591 (N_2591,N_2040,N_2169);
and U2592 (N_2592,N_2076,N_2110);
and U2593 (N_2593,N_2386,N_2171);
and U2594 (N_2594,N_2091,N_2089);
nor U2595 (N_2595,N_2010,N_2209);
nor U2596 (N_2596,N_2374,N_2298);
or U2597 (N_2597,N_2256,N_2117);
and U2598 (N_2598,N_2391,N_2052);
nor U2599 (N_2599,N_2315,N_2459);
or U2600 (N_2600,N_2086,N_2150);
nor U2601 (N_2601,N_2222,N_2134);
and U2602 (N_2602,N_2211,N_2236);
or U2603 (N_2603,N_2468,N_2037);
or U2604 (N_2604,N_2382,N_2422);
nor U2605 (N_2605,N_2000,N_2318);
or U2606 (N_2606,N_2025,N_2371);
nor U2607 (N_2607,N_2373,N_2477);
or U2608 (N_2608,N_2178,N_2138);
nand U2609 (N_2609,N_2293,N_2249);
nor U2610 (N_2610,N_2234,N_2425);
nor U2611 (N_2611,N_2461,N_2360);
nor U2612 (N_2612,N_2370,N_2158);
and U2613 (N_2613,N_2419,N_2219);
nor U2614 (N_2614,N_2019,N_2044);
and U2615 (N_2615,N_2192,N_2328);
nor U2616 (N_2616,N_2078,N_2399);
nor U2617 (N_2617,N_2479,N_2041);
xor U2618 (N_2618,N_2022,N_2473);
nand U2619 (N_2619,N_2426,N_2024);
nand U2620 (N_2620,N_2058,N_2246);
or U2621 (N_2621,N_2270,N_2074);
nor U2622 (N_2622,N_2223,N_2302);
nand U2623 (N_2623,N_2491,N_2229);
and U2624 (N_2624,N_2043,N_2368);
or U2625 (N_2625,N_2337,N_2197);
nand U2626 (N_2626,N_2132,N_2482);
or U2627 (N_2627,N_2309,N_2148);
nand U2628 (N_2628,N_2465,N_2295);
and U2629 (N_2629,N_2170,N_2413);
or U2630 (N_2630,N_2032,N_2478);
and U2631 (N_2631,N_2443,N_2400);
or U2632 (N_2632,N_2220,N_2190);
nor U2633 (N_2633,N_2361,N_2189);
nor U2634 (N_2634,N_2435,N_2314);
and U2635 (N_2635,N_2253,N_2226);
and U2636 (N_2636,N_2030,N_2496);
nand U2637 (N_2637,N_2231,N_2075);
and U2638 (N_2638,N_2180,N_2099);
nor U2639 (N_2639,N_2265,N_2228);
nand U2640 (N_2640,N_2279,N_2142);
and U2641 (N_2641,N_2412,N_2305);
and U2642 (N_2642,N_2402,N_2262);
or U2643 (N_2643,N_2421,N_2162);
nand U2644 (N_2644,N_2243,N_2418);
or U2645 (N_2645,N_2304,N_2233);
nand U2646 (N_2646,N_2250,N_2281);
nand U2647 (N_2647,N_2332,N_2372);
nor U2648 (N_2648,N_2016,N_2094);
or U2649 (N_2649,N_2241,N_2484);
nand U2650 (N_2650,N_2119,N_2115);
and U2651 (N_2651,N_2407,N_2212);
or U2652 (N_2652,N_2490,N_2452);
or U2653 (N_2653,N_2326,N_2280);
nor U2654 (N_2654,N_2062,N_2218);
nand U2655 (N_2655,N_2358,N_2410);
or U2656 (N_2656,N_2031,N_2063);
nor U2657 (N_2657,N_2144,N_2139);
or U2658 (N_2658,N_2108,N_2312);
or U2659 (N_2659,N_2384,N_2494);
and U2660 (N_2660,N_2214,N_2039);
or U2661 (N_2661,N_2104,N_2469);
and U2662 (N_2662,N_2460,N_2349);
and U2663 (N_2663,N_2411,N_2471);
nand U2664 (N_2664,N_2483,N_2498);
or U2665 (N_2665,N_2124,N_2034);
and U2666 (N_2666,N_2096,N_2423);
nand U2667 (N_2667,N_2392,N_2433);
nor U2668 (N_2668,N_2450,N_2061);
nor U2669 (N_2669,N_2369,N_2232);
nand U2670 (N_2670,N_2474,N_2118);
or U2671 (N_2671,N_2242,N_2378);
or U2672 (N_2672,N_2487,N_2299);
and U2673 (N_2673,N_2130,N_2254);
nor U2674 (N_2674,N_2060,N_2489);
and U2675 (N_2675,N_2261,N_2365);
nand U2676 (N_2676,N_2163,N_2292);
nor U2677 (N_2677,N_2245,N_2196);
or U2678 (N_2678,N_2268,N_2168);
and U2679 (N_2679,N_2161,N_2065);
and U2680 (N_2680,N_2204,N_2129);
or U2681 (N_2681,N_2004,N_2069);
nor U2682 (N_2682,N_2333,N_2339);
and U2683 (N_2683,N_2026,N_2225);
or U2684 (N_2684,N_2126,N_2475);
or U2685 (N_2685,N_2405,N_2227);
or U2686 (N_2686,N_2442,N_2105);
nand U2687 (N_2687,N_2406,N_2343);
or U2688 (N_2688,N_2252,N_2079);
nand U2689 (N_2689,N_2330,N_2160);
nor U2690 (N_2690,N_2002,N_2147);
and U2691 (N_2691,N_2029,N_2458);
xnor U2692 (N_2692,N_2350,N_2322);
or U2693 (N_2693,N_2401,N_2294);
and U2694 (N_2694,N_2432,N_2206);
nor U2695 (N_2695,N_2172,N_2437);
or U2696 (N_2696,N_2049,N_2208);
and U2697 (N_2697,N_2154,N_2390);
or U2698 (N_2698,N_2057,N_2125);
xor U2699 (N_2699,N_2319,N_2187);
and U2700 (N_2700,N_2230,N_2467);
nand U2701 (N_2701,N_2006,N_2166);
nor U2702 (N_2702,N_2289,N_2403);
and U2703 (N_2703,N_2375,N_2376);
and U2704 (N_2704,N_2014,N_2149);
or U2705 (N_2705,N_2300,N_2257);
nor U2706 (N_2706,N_2202,N_2383);
nor U2707 (N_2707,N_2303,N_2077);
nand U2708 (N_2708,N_2310,N_2430);
or U2709 (N_2709,N_2053,N_2153);
nand U2710 (N_2710,N_2357,N_2194);
and U2711 (N_2711,N_2440,N_2251);
nor U2712 (N_2712,N_2290,N_2087);
and U2713 (N_2713,N_2103,N_2054);
or U2714 (N_2714,N_2385,N_2448);
nor U2715 (N_2715,N_2165,N_2102);
and U2716 (N_2716,N_2275,N_2082);
nand U2717 (N_2717,N_2191,N_2203);
nand U2718 (N_2718,N_2200,N_2136);
xor U2719 (N_2719,N_2097,N_2329);
xnor U2720 (N_2720,N_2064,N_2364);
or U2721 (N_2721,N_2179,N_2098);
and U2722 (N_2722,N_2366,N_2109);
nor U2723 (N_2723,N_2424,N_2112);
xnor U2724 (N_2724,N_2260,N_2239);
nand U2725 (N_2725,N_2215,N_2335);
and U2726 (N_2726,N_2395,N_2051);
xnor U2727 (N_2727,N_2012,N_2240);
nor U2728 (N_2728,N_2164,N_2320);
nor U2729 (N_2729,N_2398,N_2207);
nand U2730 (N_2730,N_2146,N_2445);
nand U2731 (N_2731,N_2454,N_2313);
or U2732 (N_2732,N_2235,N_2113);
and U2733 (N_2733,N_2151,N_2334);
or U2734 (N_2734,N_2013,N_2431);
and U2735 (N_2735,N_2101,N_2428);
nor U2736 (N_2736,N_2493,N_2439);
nand U2737 (N_2737,N_2155,N_2351);
nor U2738 (N_2738,N_2420,N_2195);
nand U2739 (N_2739,N_2288,N_2481);
or U2740 (N_2740,N_2088,N_2120);
nor U2741 (N_2741,N_2045,N_2210);
nor U2742 (N_2742,N_2020,N_2084);
or U2743 (N_2743,N_2341,N_2007);
or U2744 (N_2744,N_2073,N_2001);
and U2745 (N_2745,N_2127,N_2046);
nor U2746 (N_2746,N_2201,N_2071);
or U2747 (N_2747,N_2145,N_2485);
or U2748 (N_2748,N_2186,N_2035);
nand U2749 (N_2749,N_2131,N_2008);
xnor U2750 (N_2750,N_2397,N_2057);
or U2751 (N_2751,N_2432,N_2250);
nand U2752 (N_2752,N_2393,N_2476);
nor U2753 (N_2753,N_2177,N_2145);
nand U2754 (N_2754,N_2443,N_2046);
and U2755 (N_2755,N_2008,N_2097);
nand U2756 (N_2756,N_2212,N_2327);
nor U2757 (N_2757,N_2031,N_2454);
nor U2758 (N_2758,N_2481,N_2024);
nor U2759 (N_2759,N_2132,N_2407);
and U2760 (N_2760,N_2105,N_2015);
or U2761 (N_2761,N_2260,N_2222);
nand U2762 (N_2762,N_2037,N_2080);
or U2763 (N_2763,N_2313,N_2258);
and U2764 (N_2764,N_2336,N_2327);
nor U2765 (N_2765,N_2104,N_2289);
nand U2766 (N_2766,N_2099,N_2151);
and U2767 (N_2767,N_2005,N_2410);
nand U2768 (N_2768,N_2156,N_2472);
nor U2769 (N_2769,N_2118,N_2399);
nor U2770 (N_2770,N_2355,N_2366);
and U2771 (N_2771,N_2058,N_2111);
or U2772 (N_2772,N_2018,N_2406);
nor U2773 (N_2773,N_2046,N_2320);
nor U2774 (N_2774,N_2086,N_2239);
or U2775 (N_2775,N_2023,N_2244);
and U2776 (N_2776,N_2270,N_2312);
and U2777 (N_2777,N_2204,N_2147);
nand U2778 (N_2778,N_2040,N_2367);
nand U2779 (N_2779,N_2144,N_2209);
nor U2780 (N_2780,N_2084,N_2014);
and U2781 (N_2781,N_2434,N_2149);
or U2782 (N_2782,N_2425,N_2486);
and U2783 (N_2783,N_2436,N_2141);
and U2784 (N_2784,N_2425,N_2136);
and U2785 (N_2785,N_2440,N_2493);
and U2786 (N_2786,N_2375,N_2017);
nand U2787 (N_2787,N_2439,N_2443);
and U2788 (N_2788,N_2298,N_2479);
nor U2789 (N_2789,N_2367,N_2391);
and U2790 (N_2790,N_2009,N_2388);
and U2791 (N_2791,N_2461,N_2377);
and U2792 (N_2792,N_2475,N_2010);
nor U2793 (N_2793,N_2144,N_2373);
or U2794 (N_2794,N_2042,N_2373);
nor U2795 (N_2795,N_2159,N_2158);
or U2796 (N_2796,N_2095,N_2351);
nor U2797 (N_2797,N_2096,N_2337);
or U2798 (N_2798,N_2119,N_2350);
or U2799 (N_2799,N_2043,N_2457);
nand U2800 (N_2800,N_2099,N_2360);
and U2801 (N_2801,N_2238,N_2404);
or U2802 (N_2802,N_2364,N_2349);
nor U2803 (N_2803,N_2422,N_2339);
nor U2804 (N_2804,N_2168,N_2018);
nand U2805 (N_2805,N_2198,N_2261);
or U2806 (N_2806,N_2332,N_2192);
and U2807 (N_2807,N_2485,N_2304);
nand U2808 (N_2808,N_2130,N_2230);
nor U2809 (N_2809,N_2464,N_2087);
or U2810 (N_2810,N_2087,N_2472);
nor U2811 (N_2811,N_2391,N_2301);
nor U2812 (N_2812,N_2138,N_2249);
and U2813 (N_2813,N_2123,N_2034);
nand U2814 (N_2814,N_2067,N_2066);
nor U2815 (N_2815,N_2087,N_2306);
nor U2816 (N_2816,N_2215,N_2019);
nor U2817 (N_2817,N_2349,N_2169);
and U2818 (N_2818,N_2228,N_2275);
nand U2819 (N_2819,N_2428,N_2436);
nor U2820 (N_2820,N_2448,N_2007);
and U2821 (N_2821,N_2065,N_2334);
nand U2822 (N_2822,N_2355,N_2402);
and U2823 (N_2823,N_2247,N_2006);
or U2824 (N_2824,N_2136,N_2145);
and U2825 (N_2825,N_2190,N_2060);
and U2826 (N_2826,N_2368,N_2074);
nor U2827 (N_2827,N_2303,N_2193);
nor U2828 (N_2828,N_2432,N_2067);
nor U2829 (N_2829,N_2498,N_2378);
or U2830 (N_2830,N_2089,N_2338);
nor U2831 (N_2831,N_2151,N_2258);
and U2832 (N_2832,N_2005,N_2498);
or U2833 (N_2833,N_2159,N_2319);
nor U2834 (N_2834,N_2046,N_2345);
or U2835 (N_2835,N_2367,N_2303);
xnor U2836 (N_2836,N_2005,N_2413);
and U2837 (N_2837,N_2353,N_2359);
or U2838 (N_2838,N_2141,N_2065);
and U2839 (N_2839,N_2045,N_2294);
or U2840 (N_2840,N_2040,N_2198);
nand U2841 (N_2841,N_2459,N_2414);
nand U2842 (N_2842,N_2289,N_2336);
or U2843 (N_2843,N_2193,N_2409);
and U2844 (N_2844,N_2456,N_2432);
nand U2845 (N_2845,N_2174,N_2233);
nand U2846 (N_2846,N_2135,N_2009);
or U2847 (N_2847,N_2282,N_2343);
nand U2848 (N_2848,N_2062,N_2192);
or U2849 (N_2849,N_2019,N_2221);
and U2850 (N_2850,N_2096,N_2065);
nor U2851 (N_2851,N_2058,N_2169);
and U2852 (N_2852,N_2205,N_2099);
and U2853 (N_2853,N_2297,N_2463);
and U2854 (N_2854,N_2014,N_2235);
or U2855 (N_2855,N_2100,N_2438);
nor U2856 (N_2856,N_2497,N_2365);
or U2857 (N_2857,N_2429,N_2161);
nand U2858 (N_2858,N_2481,N_2377);
and U2859 (N_2859,N_2026,N_2256);
nand U2860 (N_2860,N_2154,N_2050);
or U2861 (N_2861,N_2296,N_2190);
nand U2862 (N_2862,N_2056,N_2493);
nand U2863 (N_2863,N_2158,N_2161);
nand U2864 (N_2864,N_2130,N_2463);
and U2865 (N_2865,N_2003,N_2317);
nand U2866 (N_2866,N_2412,N_2064);
or U2867 (N_2867,N_2395,N_2307);
xor U2868 (N_2868,N_2074,N_2023);
nand U2869 (N_2869,N_2493,N_2497);
nor U2870 (N_2870,N_2372,N_2305);
and U2871 (N_2871,N_2372,N_2145);
nand U2872 (N_2872,N_2279,N_2016);
and U2873 (N_2873,N_2187,N_2099);
or U2874 (N_2874,N_2003,N_2131);
nand U2875 (N_2875,N_2405,N_2280);
and U2876 (N_2876,N_2474,N_2050);
nand U2877 (N_2877,N_2116,N_2490);
nand U2878 (N_2878,N_2357,N_2183);
nor U2879 (N_2879,N_2162,N_2101);
xnor U2880 (N_2880,N_2152,N_2130);
and U2881 (N_2881,N_2277,N_2090);
nor U2882 (N_2882,N_2194,N_2262);
and U2883 (N_2883,N_2381,N_2315);
or U2884 (N_2884,N_2290,N_2448);
or U2885 (N_2885,N_2492,N_2293);
nand U2886 (N_2886,N_2243,N_2321);
nand U2887 (N_2887,N_2116,N_2447);
or U2888 (N_2888,N_2207,N_2486);
and U2889 (N_2889,N_2217,N_2272);
and U2890 (N_2890,N_2164,N_2318);
or U2891 (N_2891,N_2313,N_2342);
and U2892 (N_2892,N_2471,N_2397);
and U2893 (N_2893,N_2128,N_2231);
nor U2894 (N_2894,N_2364,N_2449);
nor U2895 (N_2895,N_2119,N_2246);
or U2896 (N_2896,N_2161,N_2437);
nor U2897 (N_2897,N_2151,N_2177);
nor U2898 (N_2898,N_2480,N_2237);
or U2899 (N_2899,N_2327,N_2124);
and U2900 (N_2900,N_2102,N_2027);
nand U2901 (N_2901,N_2437,N_2366);
or U2902 (N_2902,N_2090,N_2401);
or U2903 (N_2903,N_2159,N_2117);
or U2904 (N_2904,N_2445,N_2197);
nor U2905 (N_2905,N_2481,N_2321);
and U2906 (N_2906,N_2019,N_2107);
and U2907 (N_2907,N_2436,N_2310);
nand U2908 (N_2908,N_2222,N_2005);
or U2909 (N_2909,N_2021,N_2380);
nand U2910 (N_2910,N_2320,N_2324);
nand U2911 (N_2911,N_2321,N_2341);
and U2912 (N_2912,N_2022,N_2310);
or U2913 (N_2913,N_2052,N_2246);
nand U2914 (N_2914,N_2131,N_2296);
nand U2915 (N_2915,N_2444,N_2341);
or U2916 (N_2916,N_2474,N_2438);
nand U2917 (N_2917,N_2254,N_2211);
nand U2918 (N_2918,N_2305,N_2127);
nor U2919 (N_2919,N_2110,N_2344);
nor U2920 (N_2920,N_2431,N_2017);
and U2921 (N_2921,N_2264,N_2224);
nor U2922 (N_2922,N_2132,N_2387);
nor U2923 (N_2923,N_2348,N_2003);
nor U2924 (N_2924,N_2313,N_2480);
and U2925 (N_2925,N_2227,N_2231);
and U2926 (N_2926,N_2255,N_2118);
and U2927 (N_2927,N_2327,N_2026);
nand U2928 (N_2928,N_2479,N_2188);
nor U2929 (N_2929,N_2467,N_2020);
and U2930 (N_2930,N_2389,N_2063);
nor U2931 (N_2931,N_2195,N_2364);
or U2932 (N_2932,N_2102,N_2337);
and U2933 (N_2933,N_2190,N_2151);
or U2934 (N_2934,N_2256,N_2317);
and U2935 (N_2935,N_2167,N_2268);
nand U2936 (N_2936,N_2194,N_2479);
and U2937 (N_2937,N_2321,N_2261);
nand U2938 (N_2938,N_2340,N_2403);
nor U2939 (N_2939,N_2257,N_2007);
nor U2940 (N_2940,N_2180,N_2148);
and U2941 (N_2941,N_2003,N_2475);
nor U2942 (N_2942,N_2037,N_2202);
or U2943 (N_2943,N_2261,N_2230);
and U2944 (N_2944,N_2312,N_2401);
nor U2945 (N_2945,N_2108,N_2321);
nand U2946 (N_2946,N_2187,N_2205);
and U2947 (N_2947,N_2396,N_2340);
or U2948 (N_2948,N_2443,N_2215);
nand U2949 (N_2949,N_2466,N_2269);
nand U2950 (N_2950,N_2114,N_2489);
or U2951 (N_2951,N_2171,N_2122);
nor U2952 (N_2952,N_2227,N_2212);
nand U2953 (N_2953,N_2146,N_2086);
nand U2954 (N_2954,N_2033,N_2066);
nand U2955 (N_2955,N_2370,N_2137);
nand U2956 (N_2956,N_2449,N_2426);
nor U2957 (N_2957,N_2402,N_2254);
or U2958 (N_2958,N_2242,N_2182);
and U2959 (N_2959,N_2124,N_2258);
nand U2960 (N_2960,N_2200,N_2364);
nor U2961 (N_2961,N_2314,N_2488);
nand U2962 (N_2962,N_2286,N_2300);
nor U2963 (N_2963,N_2377,N_2434);
nor U2964 (N_2964,N_2090,N_2497);
nand U2965 (N_2965,N_2392,N_2299);
and U2966 (N_2966,N_2249,N_2145);
nor U2967 (N_2967,N_2173,N_2037);
nand U2968 (N_2968,N_2386,N_2419);
or U2969 (N_2969,N_2321,N_2137);
nand U2970 (N_2970,N_2077,N_2482);
or U2971 (N_2971,N_2080,N_2103);
or U2972 (N_2972,N_2003,N_2205);
xnor U2973 (N_2973,N_2396,N_2329);
and U2974 (N_2974,N_2118,N_2371);
and U2975 (N_2975,N_2068,N_2223);
nand U2976 (N_2976,N_2304,N_2182);
and U2977 (N_2977,N_2153,N_2058);
or U2978 (N_2978,N_2303,N_2072);
nor U2979 (N_2979,N_2175,N_2443);
nor U2980 (N_2980,N_2177,N_2465);
or U2981 (N_2981,N_2281,N_2266);
and U2982 (N_2982,N_2414,N_2072);
or U2983 (N_2983,N_2256,N_2093);
and U2984 (N_2984,N_2213,N_2101);
nor U2985 (N_2985,N_2487,N_2006);
nor U2986 (N_2986,N_2063,N_2284);
nand U2987 (N_2987,N_2484,N_2082);
and U2988 (N_2988,N_2475,N_2085);
and U2989 (N_2989,N_2232,N_2336);
nand U2990 (N_2990,N_2247,N_2278);
nand U2991 (N_2991,N_2205,N_2170);
or U2992 (N_2992,N_2417,N_2238);
or U2993 (N_2993,N_2327,N_2194);
nand U2994 (N_2994,N_2049,N_2204);
or U2995 (N_2995,N_2395,N_2193);
nand U2996 (N_2996,N_2135,N_2258);
and U2997 (N_2997,N_2122,N_2186);
nor U2998 (N_2998,N_2298,N_2301);
or U2999 (N_2999,N_2361,N_2260);
xnor U3000 (N_3000,N_2683,N_2898);
nand U3001 (N_3001,N_2784,N_2518);
nand U3002 (N_3002,N_2821,N_2843);
nand U3003 (N_3003,N_2527,N_2867);
and U3004 (N_3004,N_2830,N_2576);
and U3005 (N_3005,N_2675,N_2988);
and U3006 (N_3006,N_2953,N_2610);
and U3007 (N_3007,N_2749,N_2906);
nand U3008 (N_3008,N_2738,N_2616);
or U3009 (N_3009,N_2710,N_2605);
or U3010 (N_3010,N_2724,N_2607);
or U3011 (N_3011,N_2554,N_2584);
and U3012 (N_3012,N_2513,N_2684);
and U3013 (N_3013,N_2729,N_2912);
nor U3014 (N_3014,N_2545,N_2794);
or U3015 (N_3015,N_2977,N_2868);
or U3016 (N_3016,N_2841,N_2742);
xor U3017 (N_3017,N_2721,N_2848);
and U3018 (N_3018,N_2884,N_2952);
nor U3019 (N_3019,N_2526,N_2731);
nand U3020 (N_3020,N_2842,N_2668);
or U3021 (N_3021,N_2549,N_2599);
nand U3022 (N_3022,N_2832,N_2822);
or U3023 (N_3023,N_2660,N_2533);
xor U3024 (N_3024,N_2747,N_2803);
and U3025 (N_3025,N_2946,N_2578);
nor U3026 (N_3026,N_2502,N_2878);
and U3027 (N_3027,N_2851,N_2839);
and U3028 (N_3028,N_2990,N_2500);
xor U3029 (N_3029,N_2857,N_2630);
and U3030 (N_3030,N_2809,N_2974);
or U3031 (N_3031,N_2662,N_2873);
nand U3032 (N_3032,N_2507,N_2654);
and U3033 (N_3033,N_2633,N_2824);
and U3034 (N_3034,N_2792,N_2618);
or U3035 (N_3035,N_2591,N_2590);
nand U3036 (N_3036,N_2674,N_2901);
nand U3037 (N_3037,N_2511,N_2850);
nor U3038 (N_3038,N_2913,N_2699);
and U3039 (N_3039,N_2734,N_2954);
nor U3040 (N_3040,N_2967,N_2916);
or U3041 (N_3041,N_2761,N_2657);
and U3042 (N_3042,N_2572,N_2997);
nor U3043 (N_3043,N_2845,N_2951);
nand U3044 (N_3044,N_2801,N_2891);
nand U3045 (N_3045,N_2930,N_2777);
or U3046 (N_3046,N_2628,N_2669);
nor U3047 (N_3047,N_2592,N_2750);
nor U3048 (N_3048,N_2785,N_2556);
and U3049 (N_3049,N_2661,N_2716);
and U3050 (N_3050,N_2732,N_2984);
nor U3051 (N_3051,N_2865,N_2604);
and U3052 (N_3052,N_2560,N_2987);
nand U3053 (N_3053,N_2547,N_2910);
nand U3054 (N_3054,N_2640,N_2852);
and U3055 (N_3055,N_2920,N_2757);
nor U3056 (N_3056,N_2712,N_2664);
nand U3057 (N_3057,N_2542,N_2594);
nor U3058 (N_3058,N_2564,N_2980);
nand U3059 (N_3059,N_2638,N_2575);
or U3060 (N_3060,N_2688,N_2771);
nor U3061 (N_3061,N_2506,N_2923);
nor U3062 (N_3062,N_2811,N_2790);
and U3063 (N_3063,N_2581,N_2634);
nand U3064 (N_3064,N_2553,N_2505);
or U3065 (N_3065,N_2515,N_2743);
and U3066 (N_3066,N_2753,N_2765);
and U3067 (N_3067,N_2966,N_2939);
or U3068 (N_3068,N_2601,N_2780);
or U3069 (N_3069,N_2998,N_2979);
xnor U3070 (N_3070,N_2817,N_2921);
and U3071 (N_3071,N_2562,N_2567);
and U3072 (N_3072,N_2972,N_2709);
or U3073 (N_3073,N_2836,N_2593);
nand U3074 (N_3074,N_2600,N_2512);
nand U3075 (N_3075,N_2529,N_2665);
xnor U3076 (N_3076,N_2825,N_2748);
nor U3077 (N_3077,N_2714,N_2508);
xnor U3078 (N_3078,N_2645,N_2537);
and U3079 (N_3079,N_2963,N_2565);
or U3080 (N_3080,N_2797,N_2677);
or U3081 (N_3081,N_2585,N_2917);
and U3082 (N_3082,N_2528,N_2615);
and U3083 (N_3083,N_2571,N_2658);
nor U3084 (N_3084,N_2597,N_2608);
nor U3085 (N_3085,N_2681,N_2978);
or U3086 (N_3086,N_2775,N_2713);
and U3087 (N_3087,N_2697,N_2859);
and U3088 (N_3088,N_2702,N_2929);
nor U3089 (N_3089,N_2989,N_2727);
or U3090 (N_3090,N_2762,N_2619);
and U3091 (N_3091,N_2760,N_2768);
nor U3092 (N_3092,N_2504,N_2999);
or U3093 (N_3093,N_2625,N_2517);
xor U3094 (N_3094,N_2530,N_2589);
nor U3095 (N_3095,N_2807,N_2755);
or U3096 (N_3096,N_2788,N_2623);
nand U3097 (N_3097,N_2812,N_2828);
nand U3098 (N_3098,N_2569,N_2687);
and U3099 (N_3099,N_2516,N_2892);
or U3100 (N_3100,N_2737,N_2538);
or U3101 (N_3101,N_2543,N_2719);
and U3102 (N_3102,N_2741,N_2586);
nand U3103 (N_3103,N_2981,N_2705);
xnor U3104 (N_3104,N_2875,N_2849);
and U3105 (N_3105,N_2961,N_2620);
nand U3106 (N_3106,N_2992,N_2795);
nand U3107 (N_3107,N_2514,N_2725);
nand U3108 (N_3108,N_2501,N_2776);
nand U3109 (N_3109,N_2635,N_2982);
nor U3110 (N_3110,N_2736,N_2927);
or U3111 (N_3111,N_2573,N_2626);
xor U3112 (N_3112,N_2864,N_2899);
and U3113 (N_3113,N_2744,N_2991);
and U3114 (N_3114,N_2770,N_2805);
or U3115 (N_3115,N_2889,N_2840);
or U3116 (N_3116,N_2940,N_2643);
and U3117 (N_3117,N_2903,N_2766);
nand U3118 (N_3118,N_2679,N_2596);
or U3119 (N_3119,N_2522,N_2796);
nor U3120 (N_3120,N_2598,N_2986);
nor U3121 (N_3121,N_2896,N_2994);
and U3122 (N_3122,N_2632,N_2609);
nand U3123 (N_3123,N_2968,N_2673);
or U3124 (N_3124,N_2872,N_2701);
and U3125 (N_3125,N_2694,N_2931);
xor U3126 (N_3126,N_2534,N_2723);
xnor U3127 (N_3127,N_2847,N_2950);
nand U3128 (N_3128,N_2810,N_2698);
nand U3129 (N_3129,N_2955,N_2733);
nand U3130 (N_3130,N_2676,N_2804);
nor U3131 (N_3131,N_2960,N_2639);
nand U3132 (N_3132,N_2861,N_2523);
nor U3133 (N_3133,N_2612,N_2708);
nand U3134 (N_3134,N_2745,N_2659);
nand U3135 (N_3135,N_2696,N_2902);
or U3136 (N_3136,N_2846,N_2831);
nand U3137 (N_3137,N_2787,N_2503);
nand U3138 (N_3138,N_2546,N_2863);
nand U3139 (N_3139,N_2566,N_2764);
and U3140 (N_3140,N_2800,N_2880);
and U3141 (N_3141,N_2704,N_2740);
or U3142 (N_3142,N_2877,N_2943);
or U3143 (N_3143,N_2922,N_2686);
nand U3144 (N_3144,N_2924,N_2641);
nor U3145 (N_3145,N_2651,N_2689);
and U3146 (N_3146,N_2541,N_2650);
nand U3147 (N_3147,N_2624,N_2959);
and U3148 (N_3148,N_2838,N_2579);
nor U3149 (N_3149,N_2636,N_2582);
nand U3150 (N_3150,N_2779,N_2844);
nand U3151 (N_3151,N_2962,N_2948);
or U3152 (N_3152,N_2897,N_2682);
nor U3153 (N_3153,N_2786,N_2672);
or U3154 (N_3154,N_2621,N_2938);
or U3155 (N_3155,N_2976,N_2835);
nor U3156 (N_3156,N_2879,N_2933);
or U3157 (N_3157,N_2778,N_2767);
nand U3158 (N_3158,N_2678,N_2829);
xor U3159 (N_3159,N_2793,N_2520);
or U3160 (N_3160,N_2552,N_2629);
nand U3161 (N_3161,N_2642,N_2914);
nand U3162 (N_3162,N_2570,N_2550);
nand U3163 (N_3163,N_2918,N_2854);
and U3164 (N_3164,N_2937,N_2957);
nor U3165 (N_3165,N_2870,N_2670);
and U3166 (N_3166,N_2646,N_2647);
and U3167 (N_3167,N_2965,N_2985);
nor U3168 (N_3168,N_2539,N_2752);
and U3169 (N_3169,N_2671,N_2819);
nor U3170 (N_3170,N_2690,N_2874);
and U3171 (N_3171,N_2995,N_2971);
xor U3172 (N_3172,N_2614,N_2622);
xor U3173 (N_3173,N_2525,N_2881);
nor U3174 (N_3174,N_2703,N_2858);
nand U3175 (N_3175,N_2885,N_2653);
nor U3176 (N_3176,N_2789,N_2866);
nand U3177 (N_3177,N_2956,N_2557);
nor U3178 (N_3178,N_2602,N_2758);
nand U3179 (N_3179,N_2540,N_2706);
nor U3180 (N_3180,N_2555,N_2637);
and U3181 (N_3181,N_2535,N_2548);
nand U3182 (N_3182,N_2739,N_2815);
nor U3183 (N_3183,N_2893,N_2595);
and U3184 (N_3184,N_2826,N_2886);
nor U3185 (N_3185,N_2656,N_2944);
nor U3186 (N_3186,N_2782,N_2876);
and U3187 (N_3187,N_2970,N_2856);
or U3188 (N_3188,N_2559,N_2587);
or U3189 (N_3189,N_2941,N_2648);
or U3190 (N_3190,N_2531,N_2655);
or U3191 (N_3191,N_2746,N_2945);
nor U3192 (N_3192,N_2915,N_2773);
or U3193 (N_3193,N_2769,N_2717);
and U3194 (N_3194,N_2942,N_2853);
and U3195 (N_3195,N_2958,N_2908);
nand U3196 (N_3196,N_2666,N_2900);
nand U3197 (N_3197,N_2925,N_2715);
or U3198 (N_3198,N_2759,N_2818);
nand U3199 (N_3199,N_2802,N_2855);
nor U3200 (N_3200,N_2799,N_2993);
or U3201 (N_3201,N_2580,N_2973);
and U3202 (N_3202,N_2860,N_2894);
nor U3203 (N_3203,N_2882,N_2983);
nand U3204 (N_3204,N_2911,N_2895);
nor U3205 (N_3205,N_2862,N_2551);
or U3206 (N_3206,N_2606,N_2627);
nor U3207 (N_3207,N_2693,N_2791);
or U3208 (N_3208,N_2772,N_2631);
xnor U3209 (N_3209,N_2837,N_2718);
nand U3210 (N_3210,N_2700,N_2722);
nand U3211 (N_3211,N_2577,N_2919);
nor U3212 (N_3212,N_2563,N_2820);
and U3213 (N_3213,N_2996,N_2935);
and U3214 (N_3214,N_2558,N_2603);
nor U3215 (N_3215,N_2969,N_2975);
nor U3216 (N_3216,N_2536,N_2947);
and U3217 (N_3217,N_2588,N_2680);
nand U3218 (N_3218,N_2926,N_2888);
nor U3219 (N_3219,N_2905,N_2833);
nand U3220 (N_3220,N_2932,N_2806);
xnor U3221 (N_3221,N_2936,N_2735);
nand U3222 (N_3222,N_2907,N_2928);
nor U3223 (N_3223,N_2568,N_2519);
or U3224 (N_3224,N_2964,N_2685);
nand U3225 (N_3225,N_2695,N_2692);
or U3226 (N_3226,N_2827,N_2871);
nand U3227 (N_3227,N_2613,N_2756);
nor U3228 (N_3228,N_2720,N_2532);
nor U3229 (N_3229,N_2561,N_2883);
and U3230 (N_3230,N_2904,N_2774);
nor U3231 (N_3231,N_2798,N_2707);
nand U3232 (N_3232,N_2611,N_2617);
nor U3233 (N_3233,N_2649,N_2663);
nand U3234 (N_3234,N_2816,N_2751);
nor U3235 (N_3235,N_2763,N_2887);
nand U3236 (N_3236,N_2667,N_2574);
and U3237 (N_3237,N_2644,N_2813);
nor U3238 (N_3238,N_2652,N_2808);
and U3239 (N_3239,N_2730,N_2909);
nand U3240 (N_3240,N_2583,N_2711);
nand U3241 (N_3241,N_2934,N_2521);
nor U3242 (N_3242,N_2869,N_2691);
and U3243 (N_3243,N_2890,N_2726);
or U3244 (N_3244,N_2509,N_2510);
and U3245 (N_3245,N_2949,N_2754);
nor U3246 (N_3246,N_2814,N_2781);
nand U3247 (N_3247,N_2728,N_2544);
nand U3248 (N_3248,N_2823,N_2524);
or U3249 (N_3249,N_2834,N_2783);
or U3250 (N_3250,N_2858,N_2611);
and U3251 (N_3251,N_2701,N_2696);
or U3252 (N_3252,N_2641,N_2872);
or U3253 (N_3253,N_2909,N_2787);
and U3254 (N_3254,N_2739,N_2717);
or U3255 (N_3255,N_2777,N_2839);
nand U3256 (N_3256,N_2728,N_2974);
and U3257 (N_3257,N_2684,N_2783);
and U3258 (N_3258,N_2550,N_2557);
or U3259 (N_3259,N_2574,N_2958);
nand U3260 (N_3260,N_2569,N_2826);
or U3261 (N_3261,N_2509,N_2753);
xnor U3262 (N_3262,N_2837,N_2731);
nor U3263 (N_3263,N_2725,N_2701);
nand U3264 (N_3264,N_2905,N_2681);
and U3265 (N_3265,N_2739,N_2772);
or U3266 (N_3266,N_2572,N_2763);
nor U3267 (N_3267,N_2827,N_2694);
nand U3268 (N_3268,N_2693,N_2884);
or U3269 (N_3269,N_2545,N_2892);
nand U3270 (N_3270,N_2539,N_2918);
nor U3271 (N_3271,N_2963,N_2626);
and U3272 (N_3272,N_2842,N_2736);
or U3273 (N_3273,N_2879,N_2941);
or U3274 (N_3274,N_2549,N_2880);
nor U3275 (N_3275,N_2732,N_2606);
or U3276 (N_3276,N_2969,N_2747);
and U3277 (N_3277,N_2707,N_2965);
or U3278 (N_3278,N_2984,N_2540);
nor U3279 (N_3279,N_2776,N_2805);
nand U3280 (N_3280,N_2755,N_2951);
nand U3281 (N_3281,N_2555,N_2678);
and U3282 (N_3282,N_2980,N_2598);
nand U3283 (N_3283,N_2802,N_2879);
nor U3284 (N_3284,N_2552,N_2911);
nor U3285 (N_3285,N_2565,N_2682);
nor U3286 (N_3286,N_2782,N_2594);
nor U3287 (N_3287,N_2960,N_2743);
nor U3288 (N_3288,N_2883,N_2905);
nand U3289 (N_3289,N_2530,N_2703);
xnor U3290 (N_3290,N_2770,N_2801);
nor U3291 (N_3291,N_2735,N_2717);
or U3292 (N_3292,N_2982,N_2622);
or U3293 (N_3293,N_2875,N_2652);
or U3294 (N_3294,N_2814,N_2842);
nor U3295 (N_3295,N_2779,N_2900);
nor U3296 (N_3296,N_2583,N_2681);
and U3297 (N_3297,N_2531,N_2786);
nor U3298 (N_3298,N_2772,N_2902);
xor U3299 (N_3299,N_2783,N_2673);
or U3300 (N_3300,N_2663,N_2652);
nand U3301 (N_3301,N_2816,N_2966);
or U3302 (N_3302,N_2712,N_2908);
or U3303 (N_3303,N_2951,N_2652);
nor U3304 (N_3304,N_2863,N_2571);
nor U3305 (N_3305,N_2793,N_2984);
nor U3306 (N_3306,N_2944,N_2823);
nand U3307 (N_3307,N_2881,N_2915);
nor U3308 (N_3308,N_2937,N_2871);
xnor U3309 (N_3309,N_2963,N_2538);
nand U3310 (N_3310,N_2793,N_2753);
and U3311 (N_3311,N_2626,N_2874);
and U3312 (N_3312,N_2628,N_2989);
or U3313 (N_3313,N_2788,N_2664);
nor U3314 (N_3314,N_2514,N_2708);
or U3315 (N_3315,N_2888,N_2688);
and U3316 (N_3316,N_2958,N_2891);
and U3317 (N_3317,N_2537,N_2664);
or U3318 (N_3318,N_2507,N_2632);
and U3319 (N_3319,N_2734,N_2793);
or U3320 (N_3320,N_2655,N_2523);
nand U3321 (N_3321,N_2590,N_2688);
or U3322 (N_3322,N_2511,N_2642);
nor U3323 (N_3323,N_2696,N_2946);
nor U3324 (N_3324,N_2590,N_2724);
nand U3325 (N_3325,N_2532,N_2799);
xnor U3326 (N_3326,N_2963,N_2740);
and U3327 (N_3327,N_2933,N_2644);
nor U3328 (N_3328,N_2941,N_2724);
and U3329 (N_3329,N_2711,N_2721);
nand U3330 (N_3330,N_2824,N_2570);
xor U3331 (N_3331,N_2622,N_2854);
and U3332 (N_3332,N_2722,N_2601);
nand U3333 (N_3333,N_2595,N_2921);
nor U3334 (N_3334,N_2742,N_2544);
nor U3335 (N_3335,N_2649,N_2744);
nand U3336 (N_3336,N_2666,N_2734);
nand U3337 (N_3337,N_2707,N_2739);
nand U3338 (N_3338,N_2527,N_2706);
nand U3339 (N_3339,N_2702,N_2769);
nor U3340 (N_3340,N_2706,N_2654);
or U3341 (N_3341,N_2718,N_2919);
or U3342 (N_3342,N_2654,N_2933);
and U3343 (N_3343,N_2522,N_2817);
nor U3344 (N_3344,N_2801,N_2874);
or U3345 (N_3345,N_2622,N_2607);
and U3346 (N_3346,N_2842,N_2520);
and U3347 (N_3347,N_2980,N_2691);
or U3348 (N_3348,N_2701,N_2643);
and U3349 (N_3349,N_2787,N_2680);
nor U3350 (N_3350,N_2663,N_2525);
and U3351 (N_3351,N_2592,N_2722);
and U3352 (N_3352,N_2601,N_2996);
nor U3353 (N_3353,N_2694,N_2606);
and U3354 (N_3354,N_2654,N_2736);
xor U3355 (N_3355,N_2677,N_2822);
and U3356 (N_3356,N_2597,N_2978);
and U3357 (N_3357,N_2684,N_2784);
and U3358 (N_3358,N_2586,N_2816);
nand U3359 (N_3359,N_2672,N_2630);
nand U3360 (N_3360,N_2797,N_2719);
nor U3361 (N_3361,N_2662,N_2974);
and U3362 (N_3362,N_2701,N_2968);
and U3363 (N_3363,N_2745,N_2827);
and U3364 (N_3364,N_2648,N_2949);
nand U3365 (N_3365,N_2641,N_2916);
and U3366 (N_3366,N_2525,N_2747);
or U3367 (N_3367,N_2562,N_2999);
or U3368 (N_3368,N_2932,N_2893);
nand U3369 (N_3369,N_2729,N_2833);
xor U3370 (N_3370,N_2869,N_2896);
or U3371 (N_3371,N_2529,N_2738);
nand U3372 (N_3372,N_2520,N_2690);
and U3373 (N_3373,N_2568,N_2929);
and U3374 (N_3374,N_2925,N_2868);
or U3375 (N_3375,N_2862,N_2514);
nand U3376 (N_3376,N_2658,N_2635);
and U3377 (N_3377,N_2557,N_2513);
nand U3378 (N_3378,N_2805,N_2605);
or U3379 (N_3379,N_2733,N_2679);
nand U3380 (N_3380,N_2950,N_2944);
or U3381 (N_3381,N_2934,N_2576);
nor U3382 (N_3382,N_2579,N_2972);
nand U3383 (N_3383,N_2949,N_2729);
nand U3384 (N_3384,N_2826,N_2787);
and U3385 (N_3385,N_2861,N_2822);
nand U3386 (N_3386,N_2781,N_2532);
and U3387 (N_3387,N_2675,N_2777);
and U3388 (N_3388,N_2663,N_2621);
or U3389 (N_3389,N_2846,N_2512);
or U3390 (N_3390,N_2918,N_2771);
nand U3391 (N_3391,N_2587,N_2512);
or U3392 (N_3392,N_2758,N_2612);
or U3393 (N_3393,N_2897,N_2875);
nand U3394 (N_3394,N_2893,N_2886);
nand U3395 (N_3395,N_2620,N_2925);
nand U3396 (N_3396,N_2728,N_2980);
or U3397 (N_3397,N_2962,N_2604);
nor U3398 (N_3398,N_2789,N_2545);
or U3399 (N_3399,N_2757,N_2689);
nor U3400 (N_3400,N_2604,N_2708);
nor U3401 (N_3401,N_2914,N_2507);
nor U3402 (N_3402,N_2954,N_2584);
or U3403 (N_3403,N_2547,N_2536);
nand U3404 (N_3404,N_2810,N_2725);
or U3405 (N_3405,N_2960,N_2545);
xor U3406 (N_3406,N_2658,N_2851);
xor U3407 (N_3407,N_2771,N_2642);
nor U3408 (N_3408,N_2658,N_2552);
nor U3409 (N_3409,N_2827,N_2540);
or U3410 (N_3410,N_2713,N_2764);
nor U3411 (N_3411,N_2648,N_2897);
or U3412 (N_3412,N_2659,N_2933);
and U3413 (N_3413,N_2898,N_2990);
and U3414 (N_3414,N_2915,N_2741);
and U3415 (N_3415,N_2907,N_2884);
nor U3416 (N_3416,N_2666,N_2866);
or U3417 (N_3417,N_2673,N_2615);
or U3418 (N_3418,N_2994,N_2718);
or U3419 (N_3419,N_2874,N_2514);
nor U3420 (N_3420,N_2990,N_2872);
or U3421 (N_3421,N_2738,N_2990);
and U3422 (N_3422,N_2789,N_2647);
and U3423 (N_3423,N_2981,N_2665);
nand U3424 (N_3424,N_2872,N_2632);
or U3425 (N_3425,N_2780,N_2925);
and U3426 (N_3426,N_2739,N_2708);
or U3427 (N_3427,N_2792,N_2690);
nand U3428 (N_3428,N_2863,N_2507);
nand U3429 (N_3429,N_2889,N_2536);
nor U3430 (N_3430,N_2807,N_2980);
and U3431 (N_3431,N_2546,N_2656);
nand U3432 (N_3432,N_2846,N_2543);
nand U3433 (N_3433,N_2620,N_2943);
or U3434 (N_3434,N_2913,N_2837);
nor U3435 (N_3435,N_2919,N_2814);
nor U3436 (N_3436,N_2546,N_2652);
and U3437 (N_3437,N_2552,N_2631);
nand U3438 (N_3438,N_2796,N_2904);
or U3439 (N_3439,N_2514,N_2607);
nor U3440 (N_3440,N_2846,N_2871);
and U3441 (N_3441,N_2556,N_2742);
nand U3442 (N_3442,N_2926,N_2874);
or U3443 (N_3443,N_2577,N_2590);
or U3444 (N_3444,N_2586,N_2647);
nor U3445 (N_3445,N_2792,N_2652);
nor U3446 (N_3446,N_2576,N_2607);
xor U3447 (N_3447,N_2849,N_2895);
or U3448 (N_3448,N_2809,N_2638);
or U3449 (N_3449,N_2759,N_2674);
nor U3450 (N_3450,N_2787,N_2533);
and U3451 (N_3451,N_2654,N_2513);
nor U3452 (N_3452,N_2716,N_2734);
nand U3453 (N_3453,N_2793,N_2719);
and U3454 (N_3454,N_2568,N_2686);
or U3455 (N_3455,N_2728,N_2768);
nand U3456 (N_3456,N_2849,N_2584);
nand U3457 (N_3457,N_2846,N_2663);
and U3458 (N_3458,N_2521,N_2681);
or U3459 (N_3459,N_2921,N_2827);
nor U3460 (N_3460,N_2521,N_2690);
or U3461 (N_3461,N_2590,N_2715);
and U3462 (N_3462,N_2578,N_2770);
and U3463 (N_3463,N_2955,N_2554);
nand U3464 (N_3464,N_2896,N_2623);
and U3465 (N_3465,N_2522,N_2747);
and U3466 (N_3466,N_2649,N_2839);
and U3467 (N_3467,N_2897,N_2975);
and U3468 (N_3468,N_2644,N_2908);
nor U3469 (N_3469,N_2617,N_2839);
nor U3470 (N_3470,N_2865,N_2940);
or U3471 (N_3471,N_2698,N_2849);
nor U3472 (N_3472,N_2662,N_2944);
nor U3473 (N_3473,N_2612,N_2522);
nand U3474 (N_3474,N_2825,N_2804);
nor U3475 (N_3475,N_2968,N_2659);
nand U3476 (N_3476,N_2613,N_2778);
nor U3477 (N_3477,N_2874,N_2927);
nand U3478 (N_3478,N_2705,N_2953);
nor U3479 (N_3479,N_2651,N_2780);
nor U3480 (N_3480,N_2602,N_2899);
nor U3481 (N_3481,N_2740,N_2874);
xnor U3482 (N_3482,N_2507,N_2801);
and U3483 (N_3483,N_2562,N_2861);
nor U3484 (N_3484,N_2510,N_2677);
and U3485 (N_3485,N_2974,N_2623);
nor U3486 (N_3486,N_2758,N_2849);
nand U3487 (N_3487,N_2529,N_2991);
or U3488 (N_3488,N_2932,N_2656);
nor U3489 (N_3489,N_2895,N_2957);
or U3490 (N_3490,N_2671,N_2553);
nor U3491 (N_3491,N_2514,N_2631);
nor U3492 (N_3492,N_2771,N_2821);
and U3493 (N_3493,N_2523,N_2604);
nor U3494 (N_3494,N_2898,N_2770);
and U3495 (N_3495,N_2601,N_2825);
or U3496 (N_3496,N_2831,N_2724);
nor U3497 (N_3497,N_2793,N_2522);
or U3498 (N_3498,N_2761,N_2925);
and U3499 (N_3499,N_2534,N_2845);
nor U3500 (N_3500,N_3111,N_3001);
nand U3501 (N_3501,N_3430,N_3158);
xor U3502 (N_3502,N_3302,N_3141);
and U3503 (N_3503,N_3088,N_3192);
nand U3504 (N_3504,N_3054,N_3032);
and U3505 (N_3505,N_3243,N_3062);
and U3506 (N_3506,N_3320,N_3377);
or U3507 (N_3507,N_3431,N_3157);
and U3508 (N_3508,N_3250,N_3145);
and U3509 (N_3509,N_3021,N_3403);
nand U3510 (N_3510,N_3372,N_3266);
nor U3511 (N_3511,N_3394,N_3240);
nand U3512 (N_3512,N_3360,N_3438);
or U3513 (N_3513,N_3080,N_3354);
nor U3514 (N_3514,N_3335,N_3125);
and U3515 (N_3515,N_3100,N_3009);
or U3516 (N_3516,N_3436,N_3131);
nand U3517 (N_3517,N_3330,N_3391);
or U3518 (N_3518,N_3288,N_3139);
nand U3519 (N_3519,N_3077,N_3228);
or U3520 (N_3520,N_3204,N_3257);
nand U3521 (N_3521,N_3282,N_3388);
and U3522 (N_3522,N_3310,N_3115);
and U3523 (N_3523,N_3448,N_3027);
nor U3524 (N_3524,N_3406,N_3223);
nand U3525 (N_3525,N_3346,N_3016);
nand U3526 (N_3526,N_3437,N_3311);
nand U3527 (N_3527,N_3269,N_3252);
or U3528 (N_3528,N_3461,N_3319);
nand U3529 (N_3529,N_3083,N_3334);
nand U3530 (N_3530,N_3270,N_3482);
nand U3531 (N_3531,N_3143,N_3091);
nor U3532 (N_3532,N_3118,N_3036);
and U3533 (N_3533,N_3155,N_3127);
nor U3534 (N_3534,N_3312,N_3201);
nand U3535 (N_3535,N_3366,N_3273);
nand U3536 (N_3536,N_3457,N_3162);
nand U3537 (N_3537,N_3220,N_3480);
nor U3538 (N_3538,N_3276,N_3426);
nand U3539 (N_3539,N_3134,N_3408);
nor U3540 (N_3540,N_3196,N_3284);
nand U3541 (N_3541,N_3447,N_3468);
nor U3542 (N_3542,N_3290,N_3488);
and U3543 (N_3543,N_3393,N_3254);
nor U3544 (N_3544,N_3443,N_3364);
and U3545 (N_3545,N_3385,N_3031);
nor U3546 (N_3546,N_3093,N_3460);
and U3547 (N_3547,N_3025,N_3184);
nand U3548 (N_3548,N_3211,N_3170);
nor U3549 (N_3549,N_3244,N_3253);
and U3550 (N_3550,N_3389,N_3456);
xor U3551 (N_3551,N_3344,N_3082);
xor U3552 (N_3552,N_3275,N_3453);
nand U3553 (N_3553,N_3322,N_3487);
nand U3554 (N_3554,N_3168,N_3029);
nor U3555 (N_3555,N_3313,N_3180);
nor U3556 (N_3556,N_3493,N_3351);
or U3557 (N_3557,N_3237,N_3151);
xor U3558 (N_3558,N_3300,N_3173);
and U3559 (N_3559,N_3022,N_3202);
nand U3560 (N_3560,N_3245,N_3114);
nand U3561 (N_3561,N_3217,N_3070);
or U3562 (N_3562,N_3489,N_3316);
and U3563 (N_3563,N_3410,N_3090);
nor U3564 (N_3564,N_3038,N_3048);
nand U3565 (N_3565,N_3246,N_3017);
and U3566 (N_3566,N_3342,N_3081);
nand U3567 (N_3567,N_3265,N_3117);
nor U3568 (N_3568,N_3105,N_3400);
nor U3569 (N_3569,N_3104,N_3185);
nor U3570 (N_3570,N_3293,N_3248);
nand U3571 (N_3571,N_3323,N_3378);
nor U3572 (N_3572,N_3361,N_3309);
nand U3573 (N_3573,N_3485,N_3238);
nor U3574 (N_3574,N_3119,N_3386);
and U3575 (N_3575,N_3398,N_3049);
and U3576 (N_3576,N_3150,N_3107);
or U3577 (N_3577,N_3010,N_3263);
nor U3578 (N_3578,N_3186,N_3262);
nor U3579 (N_3579,N_3109,N_3007);
nor U3580 (N_3580,N_3033,N_3073);
or U3581 (N_3581,N_3006,N_3218);
nand U3582 (N_3582,N_3225,N_3110);
nand U3583 (N_3583,N_3333,N_3494);
and U3584 (N_3584,N_3165,N_3210);
and U3585 (N_3585,N_3056,N_3481);
or U3586 (N_3586,N_3242,N_3195);
nor U3587 (N_3587,N_3348,N_3096);
or U3588 (N_3588,N_3241,N_3325);
and U3589 (N_3589,N_3261,N_3176);
and U3590 (N_3590,N_3414,N_3187);
nand U3591 (N_3591,N_3296,N_3317);
nand U3592 (N_3592,N_3412,N_3120);
and U3593 (N_3593,N_3129,N_3422);
nand U3594 (N_3594,N_3340,N_3402);
and U3595 (N_3595,N_3439,N_3286);
xor U3596 (N_3596,N_3067,N_3023);
or U3597 (N_3597,N_3321,N_3053);
nand U3598 (N_3598,N_3078,N_3037);
and U3599 (N_3599,N_3205,N_3281);
and U3600 (N_3600,N_3208,N_3128);
nor U3601 (N_3601,N_3459,N_3075);
nor U3602 (N_3602,N_3287,N_3188);
or U3603 (N_3603,N_3214,N_3369);
nand U3604 (N_3604,N_3024,N_3163);
and U3605 (N_3605,N_3365,N_3490);
and U3606 (N_3606,N_3015,N_3452);
nor U3607 (N_3607,N_3458,N_3209);
nor U3608 (N_3608,N_3471,N_3301);
and U3609 (N_3609,N_3464,N_3148);
nand U3610 (N_3610,N_3079,N_3387);
or U3611 (N_3611,N_3427,N_3147);
or U3612 (N_3612,N_3271,N_3052);
and U3613 (N_3613,N_3356,N_3433);
or U3614 (N_3614,N_3251,N_3071);
or U3615 (N_3615,N_3446,N_3318);
nor U3616 (N_3616,N_3470,N_3442);
nand U3617 (N_3617,N_3200,N_3449);
nand U3618 (N_3618,N_3428,N_3484);
and U3619 (N_3619,N_3383,N_3046);
nor U3620 (N_3620,N_3297,N_3455);
or U3621 (N_3621,N_3472,N_3370);
nor U3622 (N_3622,N_3206,N_3051);
xor U3623 (N_3623,N_3429,N_3355);
or U3624 (N_3624,N_3182,N_3374);
nand U3625 (N_3625,N_3064,N_3035);
or U3626 (N_3626,N_3095,N_3183);
and U3627 (N_3627,N_3123,N_3435);
or U3628 (N_3628,N_3172,N_3230);
nand U3629 (N_3629,N_3216,N_3102);
nor U3630 (N_3630,N_3327,N_3441);
and U3631 (N_3631,N_3434,N_3474);
nor U3632 (N_3632,N_3255,N_3349);
and U3633 (N_3633,N_3154,N_3042);
or U3634 (N_3634,N_3454,N_3171);
and U3635 (N_3635,N_3280,N_3231);
and U3636 (N_3636,N_3417,N_3368);
nor U3637 (N_3637,N_3373,N_3068);
or U3638 (N_3638,N_3404,N_3332);
or U3639 (N_3639,N_3138,N_3126);
nor U3640 (N_3640,N_3203,N_3416);
and U3641 (N_3641,N_3283,N_3363);
and U3642 (N_3642,N_3178,N_3177);
nor U3643 (N_3643,N_3175,N_3226);
or U3644 (N_3644,N_3142,N_3432);
nor U3645 (N_3645,N_3166,N_3299);
nor U3646 (N_3646,N_3491,N_3020);
nor U3647 (N_3647,N_3411,N_3199);
or U3648 (N_3648,N_3390,N_3087);
and U3649 (N_3649,N_3121,N_3133);
nor U3650 (N_3650,N_3419,N_3486);
and U3651 (N_3651,N_3045,N_3181);
or U3652 (N_3652,N_3063,N_3278);
and U3653 (N_3653,N_3292,N_3477);
or U3654 (N_3654,N_3074,N_3329);
xnor U3655 (N_3655,N_3149,N_3190);
nand U3656 (N_3656,N_3084,N_3294);
or U3657 (N_3657,N_3445,N_3161);
nand U3658 (N_3658,N_3350,N_3314);
nand U3659 (N_3659,N_3272,N_3153);
nor U3660 (N_3660,N_3169,N_3267);
nand U3661 (N_3661,N_3089,N_3112);
and U3662 (N_3662,N_3338,N_3232);
and U3663 (N_3663,N_3189,N_3086);
nand U3664 (N_3664,N_3308,N_3498);
and U3665 (N_3665,N_3003,N_3331);
nor U3666 (N_3666,N_3291,N_3397);
nand U3667 (N_3667,N_3156,N_3274);
or U3668 (N_3668,N_3337,N_3124);
or U3669 (N_3669,N_3092,N_3066);
nand U3670 (N_3670,N_3315,N_3179);
nand U3671 (N_3671,N_3152,N_3106);
or U3672 (N_3672,N_3420,N_3357);
or U3673 (N_3673,N_3072,N_3164);
or U3674 (N_3674,N_3116,N_3463);
and U3675 (N_3675,N_3144,N_3167);
xor U3676 (N_3676,N_3306,N_3011);
or U3677 (N_3677,N_3496,N_3019);
and U3678 (N_3678,N_3047,N_3399);
or U3679 (N_3679,N_3159,N_3444);
nor U3680 (N_3680,N_3057,N_3098);
and U3681 (N_3681,N_3101,N_3130);
nor U3682 (N_3682,N_3339,N_3371);
nand U3683 (N_3683,N_3065,N_3012);
nand U3684 (N_3684,N_3197,N_3040);
nor U3685 (N_3685,N_3499,N_3008);
and U3686 (N_3686,N_3212,N_3303);
nor U3687 (N_3687,N_3085,N_3352);
nor U3688 (N_3688,N_3440,N_3094);
nand U3689 (N_3689,N_3324,N_3384);
nand U3690 (N_3690,N_3039,N_3043);
and U3691 (N_3691,N_3140,N_3425);
nand U3692 (N_3692,N_3466,N_3343);
and U3693 (N_3693,N_3375,N_3041);
nor U3694 (N_3694,N_3227,N_3061);
and U3695 (N_3695,N_3215,N_3413);
and U3696 (N_3696,N_3328,N_3268);
and U3697 (N_3697,N_3396,N_3059);
and U3698 (N_3698,N_3376,N_3401);
and U3699 (N_3699,N_3213,N_3259);
and U3700 (N_3700,N_3279,N_3362);
nand U3701 (N_3701,N_3260,N_3450);
or U3702 (N_3702,N_3013,N_3002);
nand U3703 (N_3703,N_3160,N_3113);
nor U3704 (N_3704,N_3285,N_3359);
and U3705 (N_3705,N_3018,N_3030);
and U3706 (N_3706,N_3239,N_3277);
nor U3707 (N_3707,N_3194,N_3392);
nand U3708 (N_3708,N_3380,N_3326);
nand U3709 (N_3709,N_3307,N_3465);
nand U3710 (N_3710,N_3219,N_3367);
or U3711 (N_3711,N_3418,N_3395);
and U3712 (N_3712,N_3264,N_3233);
and U3713 (N_3713,N_3050,N_3108);
nor U3714 (N_3714,N_3132,N_3497);
nand U3715 (N_3715,N_3235,N_3295);
and U3716 (N_3716,N_3415,N_3193);
nor U3717 (N_3717,N_3221,N_3000);
xor U3718 (N_3718,N_3146,N_3492);
nand U3719 (N_3719,N_3467,N_3097);
and U3720 (N_3720,N_3345,N_3451);
and U3721 (N_3721,N_3407,N_3207);
nand U3722 (N_3722,N_3224,N_3341);
or U3723 (N_3723,N_3473,N_3256);
nand U3724 (N_3724,N_3236,N_3103);
nor U3725 (N_3725,N_3249,N_3469);
nor U3726 (N_3726,N_3135,N_3191);
or U3727 (N_3727,N_3174,N_3034);
or U3728 (N_3728,N_3136,N_3382);
nor U3729 (N_3729,N_3304,N_3005);
nand U3730 (N_3730,N_3222,N_3409);
and U3731 (N_3731,N_3423,N_3379);
nand U3732 (N_3732,N_3058,N_3495);
nor U3733 (N_3733,N_3358,N_3122);
nor U3734 (N_3734,N_3421,N_3044);
nand U3735 (N_3735,N_3198,N_3247);
nor U3736 (N_3736,N_3353,N_3405);
nor U3737 (N_3737,N_3137,N_3055);
nand U3738 (N_3738,N_3234,N_3462);
nand U3739 (N_3739,N_3289,N_3076);
and U3740 (N_3740,N_3026,N_3424);
nand U3741 (N_3741,N_3475,N_3028);
or U3742 (N_3742,N_3483,N_3478);
or U3743 (N_3743,N_3347,N_3476);
nand U3744 (N_3744,N_3336,N_3381);
nand U3745 (N_3745,N_3014,N_3069);
or U3746 (N_3746,N_3004,N_3298);
nand U3747 (N_3747,N_3060,N_3305);
or U3748 (N_3748,N_3229,N_3479);
or U3749 (N_3749,N_3258,N_3099);
xor U3750 (N_3750,N_3267,N_3075);
nor U3751 (N_3751,N_3104,N_3296);
nand U3752 (N_3752,N_3175,N_3264);
nor U3753 (N_3753,N_3296,N_3251);
nand U3754 (N_3754,N_3431,N_3034);
and U3755 (N_3755,N_3160,N_3392);
nand U3756 (N_3756,N_3422,N_3352);
xor U3757 (N_3757,N_3362,N_3273);
nand U3758 (N_3758,N_3341,N_3228);
nand U3759 (N_3759,N_3088,N_3352);
nor U3760 (N_3760,N_3177,N_3135);
and U3761 (N_3761,N_3038,N_3179);
nor U3762 (N_3762,N_3284,N_3000);
nand U3763 (N_3763,N_3328,N_3018);
nor U3764 (N_3764,N_3350,N_3483);
nor U3765 (N_3765,N_3130,N_3368);
or U3766 (N_3766,N_3470,N_3407);
or U3767 (N_3767,N_3043,N_3014);
nand U3768 (N_3768,N_3189,N_3412);
or U3769 (N_3769,N_3084,N_3271);
nand U3770 (N_3770,N_3195,N_3260);
nand U3771 (N_3771,N_3097,N_3389);
nor U3772 (N_3772,N_3435,N_3015);
or U3773 (N_3773,N_3069,N_3022);
or U3774 (N_3774,N_3132,N_3220);
and U3775 (N_3775,N_3380,N_3140);
or U3776 (N_3776,N_3297,N_3131);
and U3777 (N_3777,N_3310,N_3378);
nor U3778 (N_3778,N_3194,N_3445);
nand U3779 (N_3779,N_3186,N_3356);
or U3780 (N_3780,N_3205,N_3284);
or U3781 (N_3781,N_3394,N_3142);
or U3782 (N_3782,N_3123,N_3099);
or U3783 (N_3783,N_3481,N_3471);
nor U3784 (N_3784,N_3085,N_3137);
or U3785 (N_3785,N_3308,N_3111);
and U3786 (N_3786,N_3323,N_3250);
nor U3787 (N_3787,N_3254,N_3075);
and U3788 (N_3788,N_3355,N_3005);
nand U3789 (N_3789,N_3265,N_3125);
xnor U3790 (N_3790,N_3191,N_3289);
nor U3791 (N_3791,N_3130,N_3473);
or U3792 (N_3792,N_3118,N_3359);
nor U3793 (N_3793,N_3035,N_3043);
nor U3794 (N_3794,N_3280,N_3202);
and U3795 (N_3795,N_3222,N_3187);
nor U3796 (N_3796,N_3145,N_3388);
and U3797 (N_3797,N_3427,N_3162);
nand U3798 (N_3798,N_3022,N_3271);
or U3799 (N_3799,N_3405,N_3310);
or U3800 (N_3800,N_3321,N_3078);
nor U3801 (N_3801,N_3024,N_3066);
nand U3802 (N_3802,N_3326,N_3288);
nand U3803 (N_3803,N_3327,N_3198);
nand U3804 (N_3804,N_3101,N_3429);
nand U3805 (N_3805,N_3045,N_3073);
nand U3806 (N_3806,N_3139,N_3064);
nand U3807 (N_3807,N_3178,N_3181);
or U3808 (N_3808,N_3231,N_3085);
and U3809 (N_3809,N_3016,N_3159);
nand U3810 (N_3810,N_3449,N_3323);
and U3811 (N_3811,N_3228,N_3458);
nor U3812 (N_3812,N_3041,N_3482);
or U3813 (N_3813,N_3110,N_3127);
nand U3814 (N_3814,N_3324,N_3351);
and U3815 (N_3815,N_3253,N_3095);
and U3816 (N_3816,N_3043,N_3102);
nor U3817 (N_3817,N_3263,N_3289);
and U3818 (N_3818,N_3213,N_3091);
and U3819 (N_3819,N_3450,N_3196);
or U3820 (N_3820,N_3068,N_3005);
nand U3821 (N_3821,N_3495,N_3153);
nand U3822 (N_3822,N_3409,N_3384);
nand U3823 (N_3823,N_3082,N_3143);
or U3824 (N_3824,N_3194,N_3030);
and U3825 (N_3825,N_3097,N_3275);
or U3826 (N_3826,N_3430,N_3198);
and U3827 (N_3827,N_3142,N_3446);
and U3828 (N_3828,N_3372,N_3034);
nor U3829 (N_3829,N_3404,N_3414);
and U3830 (N_3830,N_3165,N_3006);
nand U3831 (N_3831,N_3105,N_3464);
nor U3832 (N_3832,N_3087,N_3248);
or U3833 (N_3833,N_3474,N_3292);
or U3834 (N_3834,N_3046,N_3434);
xor U3835 (N_3835,N_3420,N_3013);
nand U3836 (N_3836,N_3000,N_3492);
or U3837 (N_3837,N_3498,N_3175);
or U3838 (N_3838,N_3346,N_3450);
or U3839 (N_3839,N_3063,N_3451);
or U3840 (N_3840,N_3038,N_3087);
nor U3841 (N_3841,N_3385,N_3432);
nand U3842 (N_3842,N_3025,N_3124);
and U3843 (N_3843,N_3424,N_3110);
nand U3844 (N_3844,N_3119,N_3295);
xor U3845 (N_3845,N_3216,N_3359);
nor U3846 (N_3846,N_3454,N_3388);
nor U3847 (N_3847,N_3075,N_3125);
and U3848 (N_3848,N_3346,N_3004);
or U3849 (N_3849,N_3004,N_3390);
nand U3850 (N_3850,N_3450,N_3343);
nor U3851 (N_3851,N_3021,N_3080);
nor U3852 (N_3852,N_3444,N_3095);
and U3853 (N_3853,N_3119,N_3470);
or U3854 (N_3854,N_3217,N_3345);
and U3855 (N_3855,N_3281,N_3006);
nand U3856 (N_3856,N_3406,N_3229);
nand U3857 (N_3857,N_3227,N_3041);
or U3858 (N_3858,N_3230,N_3229);
and U3859 (N_3859,N_3101,N_3113);
nand U3860 (N_3860,N_3373,N_3317);
nand U3861 (N_3861,N_3403,N_3122);
or U3862 (N_3862,N_3401,N_3302);
xnor U3863 (N_3863,N_3159,N_3465);
or U3864 (N_3864,N_3413,N_3104);
or U3865 (N_3865,N_3393,N_3262);
and U3866 (N_3866,N_3292,N_3190);
and U3867 (N_3867,N_3210,N_3434);
and U3868 (N_3868,N_3452,N_3311);
nor U3869 (N_3869,N_3037,N_3327);
and U3870 (N_3870,N_3199,N_3154);
or U3871 (N_3871,N_3423,N_3421);
and U3872 (N_3872,N_3225,N_3459);
and U3873 (N_3873,N_3482,N_3060);
nor U3874 (N_3874,N_3073,N_3272);
nor U3875 (N_3875,N_3031,N_3122);
or U3876 (N_3876,N_3172,N_3000);
and U3877 (N_3877,N_3263,N_3032);
and U3878 (N_3878,N_3349,N_3218);
and U3879 (N_3879,N_3085,N_3183);
nor U3880 (N_3880,N_3487,N_3374);
and U3881 (N_3881,N_3014,N_3397);
nand U3882 (N_3882,N_3284,N_3069);
and U3883 (N_3883,N_3374,N_3206);
and U3884 (N_3884,N_3022,N_3354);
and U3885 (N_3885,N_3416,N_3161);
and U3886 (N_3886,N_3068,N_3325);
nand U3887 (N_3887,N_3423,N_3454);
nor U3888 (N_3888,N_3281,N_3438);
or U3889 (N_3889,N_3406,N_3161);
nor U3890 (N_3890,N_3400,N_3439);
or U3891 (N_3891,N_3269,N_3353);
xor U3892 (N_3892,N_3160,N_3043);
or U3893 (N_3893,N_3429,N_3214);
nor U3894 (N_3894,N_3484,N_3319);
or U3895 (N_3895,N_3441,N_3452);
and U3896 (N_3896,N_3498,N_3144);
nor U3897 (N_3897,N_3369,N_3365);
and U3898 (N_3898,N_3022,N_3218);
nand U3899 (N_3899,N_3289,N_3000);
and U3900 (N_3900,N_3330,N_3380);
xor U3901 (N_3901,N_3451,N_3318);
nor U3902 (N_3902,N_3298,N_3287);
or U3903 (N_3903,N_3475,N_3231);
or U3904 (N_3904,N_3438,N_3483);
nor U3905 (N_3905,N_3273,N_3377);
nand U3906 (N_3906,N_3326,N_3165);
nor U3907 (N_3907,N_3000,N_3401);
nor U3908 (N_3908,N_3315,N_3394);
xor U3909 (N_3909,N_3095,N_3273);
and U3910 (N_3910,N_3322,N_3348);
and U3911 (N_3911,N_3046,N_3483);
nor U3912 (N_3912,N_3481,N_3417);
and U3913 (N_3913,N_3211,N_3251);
or U3914 (N_3914,N_3072,N_3039);
nand U3915 (N_3915,N_3274,N_3150);
nor U3916 (N_3916,N_3292,N_3492);
xor U3917 (N_3917,N_3237,N_3080);
nand U3918 (N_3918,N_3264,N_3090);
nor U3919 (N_3919,N_3213,N_3360);
and U3920 (N_3920,N_3341,N_3130);
nor U3921 (N_3921,N_3393,N_3444);
nand U3922 (N_3922,N_3375,N_3228);
nor U3923 (N_3923,N_3065,N_3465);
and U3924 (N_3924,N_3156,N_3054);
or U3925 (N_3925,N_3176,N_3029);
nor U3926 (N_3926,N_3244,N_3481);
nand U3927 (N_3927,N_3313,N_3001);
or U3928 (N_3928,N_3121,N_3131);
and U3929 (N_3929,N_3002,N_3331);
nor U3930 (N_3930,N_3444,N_3018);
and U3931 (N_3931,N_3469,N_3165);
and U3932 (N_3932,N_3260,N_3018);
nand U3933 (N_3933,N_3242,N_3324);
and U3934 (N_3934,N_3168,N_3081);
nand U3935 (N_3935,N_3245,N_3004);
and U3936 (N_3936,N_3224,N_3144);
and U3937 (N_3937,N_3158,N_3067);
nor U3938 (N_3938,N_3376,N_3221);
and U3939 (N_3939,N_3232,N_3351);
and U3940 (N_3940,N_3415,N_3480);
or U3941 (N_3941,N_3228,N_3282);
nand U3942 (N_3942,N_3000,N_3301);
nor U3943 (N_3943,N_3353,N_3291);
and U3944 (N_3944,N_3365,N_3436);
or U3945 (N_3945,N_3100,N_3332);
nand U3946 (N_3946,N_3140,N_3189);
nor U3947 (N_3947,N_3308,N_3184);
nor U3948 (N_3948,N_3280,N_3371);
nor U3949 (N_3949,N_3186,N_3318);
nand U3950 (N_3950,N_3325,N_3342);
nand U3951 (N_3951,N_3338,N_3083);
and U3952 (N_3952,N_3086,N_3169);
nand U3953 (N_3953,N_3022,N_3002);
or U3954 (N_3954,N_3459,N_3081);
or U3955 (N_3955,N_3475,N_3165);
and U3956 (N_3956,N_3162,N_3420);
and U3957 (N_3957,N_3161,N_3381);
and U3958 (N_3958,N_3192,N_3195);
and U3959 (N_3959,N_3285,N_3453);
or U3960 (N_3960,N_3327,N_3018);
nand U3961 (N_3961,N_3460,N_3244);
nor U3962 (N_3962,N_3443,N_3388);
nand U3963 (N_3963,N_3099,N_3291);
nor U3964 (N_3964,N_3447,N_3439);
nor U3965 (N_3965,N_3272,N_3388);
nand U3966 (N_3966,N_3313,N_3489);
and U3967 (N_3967,N_3080,N_3125);
xnor U3968 (N_3968,N_3271,N_3381);
and U3969 (N_3969,N_3040,N_3265);
nor U3970 (N_3970,N_3406,N_3213);
or U3971 (N_3971,N_3315,N_3476);
nand U3972 (N_3972,N_3465,N_3064);
and U3973 (N_3973,N_3148,N_3193);
nand U3974 (N_3974,N_3320,N_3447);
or U3975 (N_3975,N_3426,N_3187);
or U3976 (N_3976,N_3048,N_3355);
and U3977 (N_3977,N_3121,N_3107);
or U3978 (N_3978,N_3342,N_3489);
xor U3979 (N_3979,N_3478,N_3273);
nor U3980 (N_3980,N_3299,N_3188);
or U3981 (N_3981,N_3244,N_3091);
or U3982 (N_3982,N_3183,N_3344);
and U3983 (N_3983,N_3391,N_3050);
nor U3984 (N_3984,N_3223,N_3193);
and U3985 (N_3985,N_3354,N_3467);
nand U3986 (N_3986,N_3499,N_3407);
nor U3987 (N_3987,N_3470,N_3374);
and U3988 (N_3988,N_3481,N_3055);
and U3989 (N_3989,N_3212,N_3470);
nand U3990 (N_3990,N_3092,N_3324);
and U3991 (N_3991,N_3212,N_3421);
nor U3992 (N_3992,N_3315,N_3297);
or U3993 (N_3993,N_3436,N_3097);
and U3994 (N_3994,N_3066,N_3112);
nand U3995 (N_3995,N_3371,N_3402);
nand U3996 (N_3996,N_3220,N_3456);
or U3997 (N_3997,N_3187,N_3348);
nor U3998 (N_3998,N_3218,N_3047);
nor U3999 (N_3999,N_3116,N_3231);
or U4000 (N_4000,N_3883,N_3542);
and U4001 (N_4001,N_3573,N_3811);
nor U4002 (N_4002,N_3941,N_3868);
nand U4003 (N_4003,N_3981,N_3676);
nand U4004 (N_4004,N_3846,N_3614);
or U4005 (N_4005,N_3949,N_3528);
nor U4006 (N_4006,N_3774,N_3964);
nor U4007 (N_4007,N_3596,N_3936);
nand U4008 (N_4008,N_3983,N_3572);
and U4009 (N_4009,N_3689,N_3996);
nand U4010 (N_4010,N_3782,N_3744);
nand U4011 (N_4011,N_3968,N_3533);
or U4012 (N_4012,N_3587,N_3647);
and U4013 (N_4013,N_3957,N_3526);
nand U4014 (N_4014,N_3829,N_3884);
nand U4015 (N_4015,N_3805,N_3831);
and U4016 (N_4016,N_3904,N_3856);
nand U4017 (N_4017,N_3928,N_3939);
nand U4018 (N_4018,N_3807,N_3621);
nand U4019 (N_4019,N_3615,N_3631);
nand U4020 (N_4020,N_3530,N_3986);
or U4021 (N_4021,N_3612,N_3879);
nor U4022 (N_4022,N_3806,N_3732);
nand U4023 (N_4023,N_3854,N_3804);
nand U4024 (N_4024,N_3842,N_3687);
nor U4025 (N_4025,N_3875,N_3849);
nor U4026 (N_4026,N_3626,N_3857);
or U4027 (N_4027,N_3843,N_3963);
or U4028 (N_4028,N_3755,N_3855);
nand U4029 (N_4029,N_3720,N_3509);
or U4030 (N_4030,N_3808,N_3645);
or U4031 (N_4031,N_3965,N_3922);
or U4032 (N_4032,N_3903,N_3802);
nand U4033 (N_4033,N_3771,N_3895);
nand U4034 (N_4034,N_3999,N_3640);
nor U4035 (N_4035,N_3628,N_3836);
nor U4036 (N_4036,N_3770,N_3582);
or U4037 (N_4037,N_3564,N_3945);
nand U4038 (N_4038,N_3905,N_3906);
nand U4039 (N_4039,N_3588,N_3861);
and U4040 (N_4040,N_3951,N_3694);
nand U4041 (N_4041,N_3544,N_3798);
and U4042 (N_4042,N_3644,N_3518);
nand U4043 (N_4043,N_3577,N_3757);
nand U4044 (N_4044,N_3671,N_3508);
nor U4045 (N_4045,N_3664,N_3723);
nand U4046 (N_4046,N_3944,N_3899);
nand U4047 (N_4047,N_3625,N_3736);
nand U4048 (N_4048,N_3975,N_3791);
and U4049 (N_4049,N_3651,N_3701);
nor U4050 (N_4050,N_3595,N_3622);
nor U4051 (N_4051,N_3926,N_3923);
nor U4052 (N_4052,N_3746,N_3649);
and U4053 (N_4053,N_3876,N_3624);
and U4054 (N_4054,N_3616,N_3589);
and U4055 (N_4055,N_3734,N_3885);
nand U4056 (N_4056,N_3768,N_3979);
and U4057 (N_4057,N_3580,N_3684);
nor U4058 (N_4058,N_3873,N_3900);
nand U4059 (N_4059,N_3597,N_3910);
and U4060 (N_4060,N_3716,N_3972);
and U4061 (N_4061,N_3514,N_3692);
nor U4062 (N_4062,N_3602,N_3813);
and U4063 (N_4063,N_3792,N_3947);
or U4064 (N_4064,N_3515,N_3554);
and U4065 (N_4065,N_3666,N_3618);
or U4066 (N_4066,N_3713,N_3810);
or U4067 (N_4067,N_3718,N_3599);
and U4068 (N_4068,N_3823,N_3998);
nor U4069 (N_4069,N_3966,N_3838);
or U4070 (N_4070,N_3632,N_3889);
nor U4071 (N_4071,N_3605,N_3866);
and U4072 (N_4072,N_3652,N_3667);
or U4073 (N_4073,N_3893,N_3953);
or U4074 (N_4074,N_3933,N_3613);
nor U4075 (N_4075,N_3752,N_3794);
nor U4076 (N_4076,N_3887,N_3783);
nand U4077 (N_4077,N_3541,N_3686);
nand U4078 (N_4078,N_3555,N_3727);
nor U4079 (N_4079,N_3679,N_3677);
and U4080 (N_4080,N_3575,N_3784);
nand U4081 (N_4081,N_3545,N_3547);
and U4082 (N_4082,N_3704,N_3673);
nand U4083 (N_4083,N_3971,N_3609);
nand U4084 (N_4084,N_3961,N_3568);
or U4085 (N_4085,N_3516,N_3705);
xor U4086 (N_4086,N_3984,N_3658);
nor U4087 (N_4087,N_3988,N_3674);
and U4088 (N_4088,N_3506,N_3559);
or U4089 (N_4089,N_3741,N_3912);
nand U4090 (N_4090,N_3598,N_3916);
or U4091 (N_4091,N_3995,N_3583);
or U4092 (N_4092,N_3991,N_3987);
and U4093 (N_4093,N_3865,N_3517);
and U4094 (N_4094,N_3604,N_3918);
or U4095 (N_4095,N_3501,N_3639);
nand U4096 (N_4096,N_3584,N_3691);
and U4097 (N_4097,N_3814,N_3540);
nor U4098 (N_4098,N_3698,N_3512);
or U4099 (N_4099,N_3897,N_3919);
or U4100 (N_4100,N_3769,N_3997);
nand U4101 (N_4101,N_3858,N_3924);
nor U4102 (N_4102,N_3730,N_3778);
nand U4103 (N_4103,N_3825,N_3859);
and U4104 (N_4104,N_3860,N_3608);
and U4105 (N_4105,N_3969,N_3753);
nand U4106 (N_4106,N_3513,N_3648);
nand U4107 (N_4107,N_3661,N_3830);
and U4108 (N_4108,N_3617,N_3525);
nand U4109 (N_4109,N_3759,N_3634);
nor U4110 (N_4110,N_3646,N_3816);
xor U4111 (N_4111,N_3940,N_3956);
or U4112 (N_4112,N_3735,N_3777);
and U4113 (N_4113,N_3915,N_3817);
and U4114 (N_4114,N_3740,N_3657);
nand U4115 (N_4115,N_3750,N_3524);
nor U4116 (N_4116,N_3781,N_3950);
nand U4117 (N_4117,N_3994,N_3815);
or U4118 (N_4118,N_3581,N_3837);
nor U4119 (N_4119,N_3891,N_3980);
or U4120 (N_4120,N_3603,N_3901);
and U4121 (N_4121,N_3502,N_3785);
or U4122 (N_4122,N_3764,N_3717);
and U4123 (N_4123,N_3952,N_3948);
or U4124 (N_4124,N_3894,N_3650);
or U4125 (N_4125,N_3557,N_3749);
nor U4126 (N_4126,N_3930,N_3641);
nor U4127 (N_4127,N_3714,N_3914);
and U4128 (N_4128,N_3707,N_3574);
nand U4129 (N_4129,N_3793,N_3549);
or U4130 (N_4130,N_3722,N_3586);
nand U4131 (N_4131,N_3668,N_3982);
nand U4132 (N_4132,N_3729,N_3503);
nand U4133 (N_4133,N_3934,N_3611);
or U4134 (N_4134,N_3537,N_3719);
nand U4135 (N_4135,N_3678,N_3977);
nor U4136 (N_4136,N_3571,N_3620);
and U4137 (N_4137,N_3702,N_3619);
or U4138 (N_4138,N_3786,N_3754);
nand U4139 (N_4139,N_3760,N_3710);
nor U4140 (N_4140,N_3536,N_3826);
nand U4141 (N_4141,N_3959,N_3960);
xor U4142 (N_4142,N_3693,N_3630);
or U4143 (N_4143,N_3908,N_3505);
and U4144 (N_4144,N_3696,N_3902);
or U4145 (N_4145,N_3762,N_3763);
nor U4146 (N_4146,N_3553,N_3844);
or U4147 (N_4147,N_3896,N_3772);
nand U4148 (N_4148,N_3569,N_3742);
and U4149 (N_4149,N_3690,N_3728);
and U4150 (N_4150,N_3898,N_3931);
nor U4151 (N_4151,N_3872,N_3504);
or U4152 (N_4152,N_3978,N_3765);
and U4153 (N_4153,N_3847,N_3797);
xnor U4154 (N_4154,N_3637,N_3954);
nor U4155 (N_4155,N_3882,N_3565);
nand U4156 (N_4156,N_3921,N_3993);
nor U4157 (N_4157,N_3510,N_3758);
and U4158 (N_4158,N_3820,N_3539);
nor U4159 (N_4159,N_3800,N_3532);
nor U4160 (N_4160,N_3890,N_3682);
nand U4161 (N_4161,N_3824,N_3976);
nand U4162 (N_4162,N_3747,N_3695);
nand U4163 (N_4163,N_3579,N_3534);
or U4164 (N_4164,N_3552,N_3548);
nand U4165 (N_4165,N_3932,N_3967);
nor U4166 (N_4166,N_3725,N_3703);
nor U4167 (N_4167,N_3828,N_3685);
nand U4168 (N_4168,N_3775,N_3946);
or U4169 (N_4169,N_3610,N_3590);
nand U4170 (N_4170,N_3839,N_3853);
nor U4171 (N_4171,N_3567,N_3809);
or U4172 (N_4172,N_3958,N_3561);
nand U4173 (N_4173,N_3560,N_3527);
or U4174 (N_4174,N_3990,N_3925);
xor U4175 (N_4175,N_3818,N_3594);
or U4176 (N_4176,N_3803,N_3636);
nand U4177 (N_4177,N_3745,N_3606);
nor U4178 (N_4178,N_3662,N_3985);
and U4179 (N_4179,N_3845,N_3708);
nor U4180 (N_4180,N_3989,N_3507);
nand U4181 (N_4181,N_3938,N_3788);
or U4182 (N_4182,N_3670,N_3672);
nand U4183 (N_4183,N_3973,N_3869);
xor U4184 (N_4184,N_3653,N_3550);
xnor U4185 (N_4185,N_3731,N_3779);
or U4186 (N_4186,N_3819,N_3748);
nand U4187 (N_4187,N_3766,N_3911);
nor U4188 (N_4188,N_3867,N_3688);
and U4189 (N_4189,N_3715,N_3870);
nand U4190 (N_4190,N_3737,N_3665);
and U4191 (N_4191,N_3700,N_3607);
nand U4192 (N_4192,N_3712,N_3871);
and U4193 (N_4193,N_3909,N_3827);
nand U4194 (N_4194,N_3751,N_3551);
and U4195 (N_4195,N_3521,N_3638);
nor U4196 (N_4196,N_3822,N_3576);
nand U4197 (N_4197,N_3711,N_3937);
or U4198 (N_4198,N_3529,N_3880);
nand U4199 (N_4199,N_3558,N_3511);
and U4200 (N_4200,N_3790,N_3538);
and U4201 (N_4201,N_3962,N_3593);
or U4202 (N_4202,N_3546,N_3724);
nand U4203 (N_4203,N_3833,N_3929);
xor U4204 (N_4204,N_3739,N_3500);
or U4205 (N_4205,N_3835,N_3773);
nand U4206 (N_4206,N_3578,N_3892);
and U4207 (N_4207,N_3681,N_3834);
and U4208 (N_4208,N_3848,N_3850);
nor U4209 (N_4209,N_3680,N_3776);
or U4210 (N_4210,N_3683,N_3821);
nand U4211 (N_4211,N_3974,N_3520);
or U4212 (N_4212,N_3881,N_3699);
and U4213 (N_4213,N_3955,N_3733);
nand U4214 (N_4214,N_3851,N_3863);
nor U4215 (N_4215,N_3756,N_3907);
and U4216 (N_4216,N_3864,N_3697);
and U4217 (N_4217,N_3927,N_3642);
nand U4218 (N_4218,N_3543,N_3886);
and U4219 (N_4219,N_3852,N_3706);
nand U4220 (N_4220,N_3629,N_3942);
nor U4221 (N_4221,N_3627,N_3888);
and U4222 (N_4222,N_3877,N_3709);
nand U4223 (N_4223,N_3663,N_3660);
and U4224 (N_4224,N_3799,N_3654);
and U4225 (N_4225,N_3920,N_3669);
or U4226 (N_4226,N_3787,N_3878);
or U4227 (N_4227,N_3935,N_3801);
nand U4228 (N_4228,N_3767,N_3743);
or U4229 (N_4229,N_3585,N_3633);
nand U4230 (N_4230,N_3563,N_3795);
or U4231 (N_4231,N_3812,N_3570);
and U4232 (N_4232,N_3556,N_3531);
nand U4233 (N_4233,N_3600,N_3643);
or U4234 (N_4234,N_3874,N_3601);
nor U4235 (N_4235,N_3659,N_3591);
and U4236 (N_4236,N_3635,N_3780);
or U4237 (N_4237,N_3841,N_3726);
nand U4238 (N_4238,N_3943,N_3562);
nand U4239 (N_4239,N_3522,N_3535);
or U4240 (N_4240,N_3523,N_3992);
and U4241 (N_4241,N_3623,N_3917);
or U4242 (N_4242,N_3721,N_3796);
or U4243 (N_4243,N_3913,N_3655);
nor U4244 (N_4244,N_3675,N_3832);
nand U4245 (N_4245,N_3970,N_3840);
or U4246 (N_4246,N_3656,N_3761);
nor U4247 (N_4247,N_3789,N_3592);
and U4248 (N_4248,N_3862,N_3738);
or U4249 (N_4249,N_3519,N_3566);
nand U4250 (N_4250,N_3746,N_3765);
nor U4251 (N_4251,N_3757,N_3653);
nor U4252 (N_4252,N_3742,N_3909);
nor U4253 (N_4253,N_3600,N_3969);
and U4254 (N_4254,N_3657,N_3647);
nand U4255 (N_4255,N_3785,N_3912);
and U4256 (N_4256,N_3753,N_3751);
xnor U4257 (N_4257,N_3983,N_3818);
nor U4258 (N_4258,N_3765,N_3603);
nor U4259 (N_4259,N_3823,N_3830);
and U4260 (N_4260,N_3889,N_3947);
and U4261 (N_4261,N_3616,N_3693);
nor U4262 (N_4262,N_3667,N_3502);
and U4263 (N_4263,N_3592,N_3580);
nand U4264 (N_4264,N_3579,N_3751);
and U4265 (N_4265,N_3935,N_3899);
and U4266 (N_4266,N_3616,N_3741);
nor U4267 (N_4267,N_3719,N_3573);
nand U4268 (N_4268,N_3970,N_3716);
or U4269 (N_4269,N_3537,N_3627);
nor U4270 (N_4270,N_3701,N_3592);
or U4271 (N_4271,N_3705,N_3951);
nor U4272 (N_4272,N_3638,N_3916);
nor U4273 (N_4273,N_3641,N_3682);
nor U4274 (N_4274,N_3834,N_3886);
and U4275 (N_4275,N_3939,N_3616);
nand U4276 (N_4276,N_3747,N_3639);
and U4277 (N_4277,N_3874,N_3891);
or U4278 (N_4278,N_3745,N_3536);
nand U4279 (N_4279,N_3656,N_3653);
or U4280 (N_4280,N_3522,N_3917);
and U4281 (N_4281,N_3518,N_3885);
nor U4282 (N_4282,N_3621,N_3509);
nor U4283 (N_4283,N_3971,N_3568);
and U4284 (N_4284,N_3713,N_3678);
xor U4285 (N_4285,N_3576,N_3778);
or U4286 (N_4286,N_3529,N_3717);
or U4287 (N_4287,N_3945,N_3541);
nand U4288 (N_4288,N_3927,N_3512);
nor U4289 (N_4289,N_3536,N_3578);
nor U4290 (N_4290,N_3574,N_3732);
nand U4291 (N_4291,N_3791,N_3776);
nor U4292 (N_4292,N_3781,N_3619);
and U4293 (N_4293,N_3926,N_3528);
and U4294 (N_4294,N_3637,N_3588);
or U4295 (N_4295,N_3885,N_3599);
nand U4296 (N_4296,N_3629,N_3957);
or U4297 (N_4297,N_3994,N_3998);
and U4298 (N_4298,N_3519,N_3768);
or U4299 (N_4299,N_3596,N_3844);
nor U4300 (N_4300,N_3797,N_3891);
nor U4301 (N_4301,N_3910,N_3651);
nand U4302 (N_4302,N_3839,N_3780);
nor U4303 (N_4303,N_3829,N_3967);
nor U4304 (N_4304,N_3527,N_3870);
and U4305 (N_4305,N_3653,N_3501);
nand U4306 (N_4306,N_3787,N_3979);
and U4307 (N_4307,N_3751,N_3552);
or U4308 (N_4308,N_3663,N_3827);
nor U4309 (N_4309,N_3549,N_3622);
and U4310 (N_4310,N_3944,N_3525);
nand U4311 (N_4311,N_3573,N_3825);
and U4312 (N_4312,N_3757,N_3976);
nand U4313 (N_4313,N_3901,N_3759);
or U4314 (N_4314,N_3720,N_3734);
nand U4315 (N_4315,N_3946,N_3914);
nor U4316 (N_4316,N_3995,N_3906);
nand U4317 (N_4317,N_3690,N_3503);
nor U4318 (N_4318,N_3953,N_3920);
nand U4319 (N_4319,N_3662,N_3774);
or U4320 (N_4320,N_3852,N_3977);
nor U4321 (N_4321,N_3611,N_3546);
nand U4322 (N_4322,N_3514,N_3776);
and U4323 (N_4323,N_3957,N_3604);
and U4324 (N_4324,N_3567,N_3759);
nand U4325 (N_4325,N_3678,N_3827);
nand U4326 (N_4326,N_3692,N_3547);
nand U4327 (N_4327,N_3704,N_3509);
nor U4328 (N_4328,N_3716,N_3961);
and U4329 (N_4329,N_3562,N_3560);
nor U4330 (N_4330,N_3738,N_3968);
or U4331 (N_4331,N_3757,N_3560);
and U4332 (N_4332,N_3939,N_3993);
nand U4333 (N_4333,N_3647,N_3844);
nor U4334 (N_4334,N_3859,N_3694);
and U4335 (N_4335,N_3597,N_3616);
or U4336 (N_4336,N_3623,N_3984);
nand U4337 (N_4337,N_3726,N_3652);
and U4338 (N_4338,N_3630,N_3842);
or U4339 (N_4339,N_3567,N_3743);
and U4340 (N_4340,N_3547,N_3894);
nor U4341 (N_4341,N_3651,N_3897);
nor U4342 (N_4342,N_3566,N_3974);
nand U4343 (N_4343,N_3590,N_3621);
and U4344 (N_4344,N_3614,N_3576);
nand U4345 (N_4345,N_3872,N_3686);
or U4346 (N_4346,N_3666,N_3913);
and U4347 (N_4347,N_3752,N_3637);
nand U4348 (N_4348,N_3539,N_3519);
nand U4349 (N_4349,N_3522,N_3971);
nor U4350 (N_4350,N_3859,N_3707);
or U4351 (N_4351,N_3855,N_3910);
and U4352 (N_4352,N_3853,N_3611);
nor U4353 (N_4353,N_3935,N_3642);
nor U4354 (N_4354,N_3679,N_3765);
or U4355 (N_4355,N_3991,N_3533);
nand U4356 (N_4356,N_3657,N_3971);
nand U4357 (N_4357,N_3602,N_3805);
or U4358 (N_4358,N_3596,N_3508);
nand U4359 (N_4359,N_3714,N_3727);
or U4360 (N_4360,N_3806,N_3804);
nor U4361 (N_4361,N_3764,N_3809);
and U4362 (N_4362,N_3510,N_3817);
and U4363 (N_4363,N_3627,N_3953);
nor U4364 (N_4364,N_3870,N_3958);
nor U4365 (N_4365,N_3506,N_3600);
nand U4366 (N_4366,N_3671,N_3542);
or U4367 (N_4367,N_3587,N_3550);
or U4368 (N_4368,N_3666,N_3722);
xnor U4369 (N_4369,N_3594,N_3872);
nor U4370 (N_4370,N_3929,N_3604);
nand U4371 (N_4371,N_3833,N_3626);
nor U4372 (N_4372,N_3653,N_3942);
and U4373 (N_4373,N_3873,N_3649);
nor U4374 (N_4374,N_3868,N_3758);
and U4375 (N_4375,N_3502,N_3529);
or U4376 (N_4376,N_3617,N_3688);
or U4377 (N_4377,N_3787,N_3895);
or U4378 (N_4378,N_3981,N_3663);
or U4379 (N_4379,N_3711,N_3660);
and U4380 (N_4380,N_3544,N_3989);
and U4381 (N_4381,N_3556,N_3701);
nand U4382 (N_4382,N_3580,N_3972);
nor U4383 (N_4383,N_3587,N_3878);
nand U4384 (N_4384,N_3800,N_3758);
and U4385 (N_4385,N_3609,N_3795);
nand U4386 (N_4386,N_3564,N_3850);
or U4387 (N_4387,N_3757,N_3872);
nor U4388 (N_4388,N_3978,N_3755);
nor U4389 (N_4389,N_3881,N_3852);
nor U4390 (N_4390,N_3606,N_3880);
nor U4391 (N_4391,N_3729,N_3836);
or U4392 (N_4392,N_3808,N_3535);
and U4393 (N_4393,N_3675,N_3792);
nand U4394 (N_4394,N_3759,N_3540);
nor U4395 (N_4395,N_3552,N_3750);
or U4396 (N_4396,N_3870,N_3938);
or U4397 (N_4397,N_3645,N_3802);
nand U4398 (N_4398,N_3719,N_3855);
and U4399 (N_4399,N_3675,N_3990);
nand U4400 (N_4400,N_3553,N_3816);
nand U4401 (N_4401,N_3744,N_3680);
nand U4402 (N_4402,N_3542,N_3942);
and U4403 (N_4403,N_3935,N_3921);
nand U4404 (N_4404,N_3647,N_3875);
nand U4405 (N_4405,N_3524,N_3707);
nor U4406 (N_4406,N_3949,N_3628);
or U4407 (N_4407,N_3733,N_3601);
and U4408 (N_4408,N_3850,N_3513);
or U4409 (N_4409,N_3853,N_3692);
nor U4410 (N_4410,N_3828,N_3827);
and U4411 (N_4411,N_3721,N_3916);
and U4412 (N_4412,N_3928,N_3881);
nand U4413 (N_4413,N_3714,N_3539);
nor U4414 (N_4414,N_3912,N_3517);
and U4415 (N_4415,N_3509,N_3794);
nand U4416 (N_4416,N_3702,N_3738);
and U4417 (N_4417,N_3515,N_3729);
and U4418 (N_4418,N_3500,N_3691);
nand U4419 (N_4419,N_3978,N_3712);
or U4420 (N_4420,N_3628,N_3824);
and U4421 (N_4421,N_3677,N_3957);
or U4422 (N_4422,N_3642,N_3993);
or U4423 (N_4423,N_3573,N_3736);
nand U4424 (N_4424,N_3570,N_3918);
or U4425 (N_4425,N_3921,N_3715);
or U4426 (N_4426,N_3955,N_3598);
and U4427 (N_4427,N_3594,N_3611);
nand U4428 (N_4428,N_3972,N_3552);
and U4429 (N_4429,N_3738,N_3582);
nand U4430 (N_4430,N_3756,N_3769);
and U4431 (N_4431,N_3992,N_3822);
and U4432 (N_4432,N_3528,N_3698);
and U4433 (N_4433,N_3709,N_3544);
nor U4434 (N_4434,N_3522,N_3685);
or U4435 (N_4435,N_3517,N_3821);
nor U4436 (N_4436,N_3905,N_3816);
nor U4437 (N_4437,N_3534,N_3547);
or U4438 (N_4438,N_3749,N_3720);
nand U4439 (N_4439,N_3904,N_3566);
nor U4440 (N_4440,N_3512,N_3803);
nor U4441 (N_4441,N_3817,N_3934);
xnor U4442 (N_4442,N_3762,N_3520);
and U4443 (N_4443,N_3713,N_3703);
nor U4444 (N_4444,N_3938,N_3514);
nand U4445 (N_4445,N_3547,N_3660);
nand U4446 (N_4446,N_3706,N_3584);
or U4447 (N_4447,N_3602,N_3851);
and U4448 (N_4448,N_3545,N_3537);
or U4449 (N_4449,N_3799,N_3942);
or U4450 (N_4450,N_3560,N_3659);
and U4451 (N_4451,N_3577,N_3804);
nand U4452 (N_4452,N_3778,N_3737);
nor U4453 (N_4453,N_3515,N_3995);
nor U4454 (N_4454,N_3782,N_3965);
and U4455 (N_4455,N_3866,N_3739);
nor U4456 (N_4456,N_3984,N_3993);
nor U4457 (N_4457,N_3540,N_3647);
nand U4458 (N_4458,N_3882,N_3577);
nand U4459 (N_4459,N_3508,N_3661);
nand U4460 (N_4460,N_3529,N_3735);
nor U4461 (N_4461,N_3656,N_3618);
nor U4462 (N_4462,N_3992,N_3732);
or U4463 (N_4463,N_3549,N_3783);
or U4464 (N_4464,N_3503,N_3937);
or U4465 (N_4465,N_3505,N_3939);
and U4466 (N_4466,N_3694,N_3920);
nor U4467 (N_4467,N_3958,N_3898);
and U4468 (N_4468,N_3931,N_3946);
nand U4469 (N_4469,N_3905,N_3711);
and U4470 (N_4470,N_3864,N_3616);
or U4471 (N_4471,N_3706,N_3898);
and U4472 (N_4472,N_3591,N_3551);
or U4473 (N_4473,N_3936,N_3840);
and U4474 (N_4474,N_3984,N_3644);
or U4475 (N_4475,N_3965,N_3831);
and U4476 (N_4476,N_3574,N_3593);
and U4477 (N_4477,N_3989,N_3972);
nand U4478 (N_4478,N_3904,N_3850);
nand U4479 (N_4479,N_3533,N_3710);
nand U4480 (N_4480,N_3952,N_3507);
nor U4481 (N_4481,N_3883,N_3650);
nor U4482 (N_4482,N_3726,N_3879);
and U4483 (N_4483,N_3926,N_3619);
nand U4484 (N_4484,N_3930,N_3666);
nand U4485 (N_4485,N_3608,N_3596);
or U4486 (N_4486,N_3871,N_3673);
nand U4487 (N_4487,N_3600,N_3795);
nor U4488 (N_4488,N_3849,N_3869);
and U4489 (N_4489,N_3613,N_3537);
or U4490 (N_4490,N_3768,N_3559);
nand U4491 (N_4491,N_3821,N_3504);
and U4492 (N_4492,N_3909,N_3691);
and U4493 (N_4493,N_3913,N_3738);
nand U4494 (N_4494,N_3586,N_3813);
nand U4495 (N_4495,N_3721,N_3794);
xnor U4496 (N_4496,N_3537,N_3707);
nor U4497 (N_4497,N_3893,N_3695);
or U4498 (N_4498,N_3718,N_3949);
and U4499 (N_4499,N_3621,N_3919);
and U4500 (N_4500,N_4308,N_4231);
nand U4501 (N_4501,N_4462,N_4410);
or U4502 (N_4502,N_4419,N_4254);
or U4503 (N_4503,N_4348,N_4489);
or U4504 (N_4504,N_4443,N_4343);
nor U4505 (N_4505,N_4272,N_4420);
nor U4506 (N_4506,N_4166,N_4131);
nand U4507 (N_4507,N_4279,N_4426);
nand U4508 (N_4508,N_4468,N_4390);
nor U4509 (N_4509,N_4003,N_4371);
nor U4510 (N_4510,N_4025,N_4028);
xnor U4511 (N_4511,N_4138,N_4071);
nand U4512 (N_4512,N_4212,N_4140);
or U4513 (N_4513,N_4347,N_4320);
nor U4514 (N_4514,N_4268,N_4185);
nor U4515 (N_4515,N_4394,N_4305);
xnor U4516 (N_4516,N_4139,N_4043);
and U4517 (N_4517,N_4041,N_4039);
nand U4518 (N_4518,N_4341,N_4016);
and U4519 (N_4519,N_4022,N_4467);
nand U4520 (N_4520,N_4366,N_4129);
and U4521 (N_4521,N_4407,N_4454);
and U4522 (N_4522,N_4321,N_4284);
and U4523 (N_4523,N_4157,N_4178);
and U4524 (N_4524,N_4481,N_4463);
and U4525 (N_4525,N_4309,N_4474);
and U4526 (N_4526,N_4108,N_4170);
or U4527 (N_4527,N_4069,N_4063);
nand U4528 (N_4528,N_4261,N_4336);
nor U4529 (N_4529,N_4109,N_4154);
or U4530 (N_4530,N_4058,N_4115);
nand U4531 (N_4531,N_4496,N_4062);
nand U4532 (N_4532,N_4297,N_4223);
nand U4533 (N_4533,N_4213,N_4285);
xnor U4534 (N_4534,N_4357,N_4358);
nand U4535 (N_4535,N_4018,N_4097);
or U4536 (N_4536,N_4056,N_4262);
or U4537 (N_4537,N_4110,N_4265);
and U4538 (N_4538,N_4064,N_4125);
and U4539 (N_4539,N_4456,N_4252);
and U4540 (N_4540,N_4447,N_4165);
and U4541 (N_4541,N_4246,N_4104);
nand U4542 (N_4542,N_4092,N_4255);
or U4543 (N_4543,N_4106,N_4217);
nand U4544 (N_4544,N_4449,N_4082);
or U4545 (N_4545,N_4179,N_4114);
nand U4546 (N_4546,N_4382,N_4205);
nor U4547 (N_4547,N_4403,N_4368);
xor U4548 (N_4548,N_4460,N_4107);
xnor U4549 (N_4549,N_4180,N_4015);
or U4550 (N_4550,N_4423,N_4073);
nand U4551 (N_4551,N_4220,N_4075);
or U4552 (N_4552,N_4037,N_4375);
nand U4553 (N_4553,N_4381,N_4036);
nand U4554 (N_4554,N_4136,N_4488);
nand U4555 (N_4555,N_4406,N_4388);
and U4556 (N_4556,N_4155,N_4159);
or U4557 (N_4557,N_4392,N_4156);
or U4558 (N_4558,N_4291,N_4427);
or U4559 (N_4559,N_4337,N_4006);
nor U4560 (N_4560,N_4280,N_4144);
or U4561 (N_4561,N_4293,N_4070);
and U4562 (N_4562,N_4163,N_4451);
nor U4563 (N_4563,N_4226,N_4486);
nor U4564 (N_4564,N_4356,N_4049);
nor U4565 (N_4565,N_4493,N_4266);
and U4566 (N_4566,N_4495,N_4300);
and U4567 (N_4567,N_4401,N_4499);
nand U4568 (N_4568,N_4278,N_4283);
and U4569 (N_4569,N_4301,N_4079);
and U4570 (N_4570,N_4353,N_4333);
and U4571 (N_4571,N_4076,N_4210);
and U4572 (N_4572,N_4424,N_4100);
nor U4573 (N_4573,N_4415,N_4004);
nand U4574 (N_4574,N_4450,N_4497);
and U4575 (N_4575,N_4033,N_4169);
nand U4576 (N_4576,N_4096,N_4351);
nor U4577 (N_4577,N_4304,N_4490);
nor U4578 (N_4578,N_4314,N_4000);
nor U4579 (N_4579,N_4142,N_4409);
or U4580 (N_4580,N_4483,N_4149);
and U4581 (N_4581,N_4471,N_4350);
or U4582 (N_4582,N_4319,N_4440);
nor U4583 (N_4583,N_4445,N_4273);
nand U4584 (N_4584,N_4235,N_4020);
or U4585 (N_4585,N_4077,N_4380);
nand U4586 (N_4586,N_4362,N_4355);
nor U4587 (N_4587,N_4292,N_4001);
and U4588 (N_4588,N_4202,N_4168);
nand U4589 (N_4589,N_4122,N_4247);
and U4590 (N_4590,N_4167,N_4444);
nor U4591 (N_4591,N_4418,N_4377);
nand U4592 (N_4592,N_4085,N_4386);
nor U4593 (N_4593,N_4051,N_4074);
nand U4594 (N_4594,N_4188,N_4479);
nor U4595 (N_4595,N_4325,N_4295);
nand U4596 (N_4596,N_4038,N_4439);
or U4597 (N_4597,N_4208,N_4172);
nor U4598 (N_4598,N_4431,N_4236);
xnor U4599 (N_4599,N_4365,N_4339);
and U4600 (N_4600,N_4067,N_4099);
nor U4601 (N_4601,N_4199,N_4050);
and U4602 (N_4602,N_4316,N_4225);
nor U4603 (N_4603,N_4430,N_4143);
or U4604 (N_4604,N_4412,N_4322);
or U4605 (N_4605,N_4492,N_4118);
nor U4606 (N_4606,N_4303,N_4219);
and U4607 (N_4607,N_4413,N_4414);
or U4608 (N_4608,N_4132,N_4234);
nand U4609 (N_4609,N_4434,N_4194);
and U4610 (N_4610,N_4196,N_4453);
and U4611 (N_4611,N_4089,N_4171);
or U4612 (N_4612,N_4152,N_4281);
nor U4613 (N_4613,N_4014,N_4200);
or U4614 (N_4614,N_4083,N_4206);
or U4615 (N_4615,N_4428,N_4233);
nor U4616 (N_4616,N_4105,N_4398);
or U4617 (N_4617,N_4080,N_4387);
nand U4618 (N_4618,N_4019,N_4193);
nor U4619 (N_4619,N_4465,N_4094);
and U4620 (N_4620,N_4175,N_4340);
and U4621 (N_4621,N_4310,N_4189);
or U4622 (N_4622,N_4209,N_4017);
and U4623 (N_4623,N_4197,N_4057);
nand U4624 (N_4624,N_4035,N_4250);
or U4625 (N_4625,N_4068,N_4251);
or U4626 (N_4626,N_4191,N_4151);
nand U4627 (N_4627,N_4240,N_4120);
or U4628 (N_4628,N_4186,N_4317);
or U4629 (N_4629,N_4065,N_4203);
nor U4630 (N_4630,N_4446,N_4150);
or U4631 (N_4631,N_4369,N_4072);
nand U4632 (N_4632,N_4329,N_4248);
or U4633 (N_4633,N_4135,N_4258);
or U4634 (N_4634,N_4269,N_4026);
or U4635 (N_4635,N_4103,N_4346);
nor U4636 (N_4636,N_4482,N_4306);
nand U4637 (N_4637,N_4148,N_4081);
and U4638 (N_4638,N_4095,N_4271);
or U4639 (N_4639,N_4374,N_4393);
and U4640 (N_4640,N_4345,N_4121);
nand U4641 (N_4641,N_4048,N_4024);
and U4642 (N_4642,N_4147,N_4086);
and U4643 (N_4643,N_4184,N_4181);
and U4644 (N_4644,N_4034,N_4298);
and U4645 (N_4645,N_4290,N_4249);
nor U4646 (N_4646,N_4124,N_4128);
or U4647 (N_4647,N_4422,N_4243);
or U4648 (N_4648,N_4494,N_4241);
nand U4649 (N_4649,N_4245,N_4123);
nor U4650 (N_4650,N_4127,N_4327);
and U4651 (N_4651,N_4146,N_4111);
and U4652 (N_4652,N_4432,N_4360);
and U4653 (N_4653,N_4173,N_4055);
nor U4654 (N_4654,N_4417,N_4260);
nor U4655 (N_4655,N_4384,N_4416);
nand U4656 (N_4656,N_4002,N_4311);
nand U4657 (N_4657,N_4441,N_4257);
or U4658 (N_4658,N_4045,N_4376);
xor U4659 (N_4659,N_4389,N_4397);
xor U4660 (N_4660,N_4359,N_4400);
and U4661 (N_4661,N_4455,N_4112);
and U4662 (N_4662,N_4078,N_4029);
and U4663 (N_4663,N_4373,N_4484);
nor U4664 (N_4664,N_4183,N_4237);
nor U4665 (N_4665,N_4402,N_4378);
nand U4666 (N_4666,N_4330,N_4141);
and U4667 (N_4667,N_4385,N_4093);
nor U4668 (N_4668,N_4054,N_4338);
or U4669 (N_4669,N_4023,N_4021);
nand U4670 (N_4670,N_4161,N_4469);
or U4671 (N_4671,N_4195,N_4204);
or U4672 (N_4672,N_4405,N_4383);
nor U4673 (N_4673,N_4164,N_4046);
nor U4674 (N_4674,N_4399,N_4008);
nor U4675 (N_4675,N_4174,N_4349);
nand U4676 (N_4676,N_4344,N_4032);
and U4677 (N_4677,N_4287,N_4053);
and U4678 (N_4678,N_4084,N_4228);
nand U4679 (N_4679,N_4176,N_4372);
or U4680 (N_4680,N_4192,N_4498);
nand U4681 (N_4681,N_4294,N_4088);
nor U4682 (N_4682,N_4211,N_4429);
nor U4683 (N_4683,N_4059,N_4060);
and U4684 (N_4684,N_4364,N_4130);
nand U4685 (N_4685,N_4354,N_4207);
and U4686 (N_4686,N_4090,N_4040);
and U4687 (N_4687,N_4425,N_4464);
nor U4688 (N_4688,N_4277,N_4491);
xnor U4689 (N_4689,N_4324,N_4027);
nor U4690 (N_4690,N_4012,N_4145);
and U4691 (N_4691,N_4201,N_4153);
nor U4692 (N_4692,N_4487,N_4315);
nand U4693 (N_4693,N_4408,N_4274);
nor U4694 (N_4694,N_4473,N_4031);
or U4695 (N_4695,N_4232,N_4326);
nor U4696 (N_4696,N_4052,N_4323);
nor U4697 (N_4697,N_4335,N_4087);
and U4698 (N_4698,N_4459,N_4448);
or U4699 (N_4699,N_4244,N_4263);
and U4700 (N_4700,N_4442,N_4466);
nand U4701 (N_4701,N_4238,N_4119);
nor U4702 (N_4702,N_4276,N_4066);
or U4703 (N_4703,N_4370,N_4352);
or U4704 (N_4704,N_4182,N_4475);
nand U4705 (N_4705,N_4190,N_4224);
and U4706 (N_4706,N_4332,N_4411);
nand U4707 (N_4707,N_4458,N_4379);
nand U4708 (N_4708,N_4457,N_4478);
xor U4709 (N_4709,N_4229,N_4286);
nand U4710 (N_4710,N_4101,N_4328);
and U4711 (N_4711,N_4296,N_4342);
or U4712 (N_4712,N_4331,N_4299);
nor U4713 (N_4713,N_4162,N_4396);
or U4714 (N_4714,N_4098,N_4134);
nor U4715 (N_4715,N_4361,N_4334);
and U4716 (N_4716,N_4476,N_4230);
nand U4717 (N_4717,N_4367,N_4198);
and U4718 (N_4718,N_4264,N_4282);
and U4719 (N_4719,N_4275,N_4007);
nor U4720 (N_4720,N_4116,N_4126);
nor U4721 (N_4721,N_4470,N_4435);
and U4722 (N_4722,N_4160,N_4061);
xnor U4723 (N_4723,N_4437,N_4158);
nor U4724 (N_4724,N_4461,N_4404);
nand U4725 (N_4725,N_4009,N_4363);
or U4726 (N_4726,N_4117,N_4477);
or U4727 (N_4727,N_4013,N_4480);
or U4728 (N_4728,N_4102,N_4288);
nand U4729 (N_4729,N_4239,N_4289);
and U4730 (N_4730,N_4438,N_4221);
nand U4731 (N_4731,N_4177,N_4307);
nor U4732 (N_4732,N_4133,N_4242);
nand U4733 (N_4733,N_4472,N_4214);
and U4734 (N_4734,N_4030,N_4421);
nand U4735 (N_4735,N_4137,N_4042);
nor U4736 (N_4736,N_4259,N_4391);
and U4737 (N_4737,N_4227,N_4485);
nand U4738 (N_4738,N_4253,N_4005);
and U4739 (N_4739,N_4318,N_4270);
nor U4740 (N_4740,N_4011,N_4436);
nor U4741 (N_4741,N_4313,N_4010);
nand U4742 (N_4742,N_4187,N_4222);
and U4743 (N_4743,N_4216,N_4113);
nand U4744 (N_4744,N_4312,N_4091);
or U4745 (N_4745,N_4302,N_4256);
and U4746 (N_4746,N_4218,N_4433);
nand U4747 (N_4747,N_4267,N_4395);
nand U4748 (N_4748,N_4452,N_4215);
nand U4749 (N_4749,N_4047,N_4044);
or U4750 (N_4750,N_4048,N_4063);
nor U4751 (N_4751,N_4182,N_4105);
nor U4752 (N_4752,N_4310,N_4165);
or U4753 (N_4753,N_4050,N_4123);
or U4754 (N_4754,N_4337,N_4206);
nand U4755 (N_4755,N_4339,N_4069);
nand U4756 (N_4756,N_4040,N_4483);
nand U4757 (N_4757,N_4088,N_4243);
and U4758 (N_4758,N_4429,N_4358);
or U4759 (N_4759,N_4147,N_4053);
or U4760 (N_4760,N_4107,N_4194);
or U4761 (N_4761,N_4394,N_4323);
nor U4762 (N_4762,N_4119,N_4249);
and U4763 (N_4763,N_4205,N_4066);
nand U4764 (N_4764,N_4190,N_4026);
and U4765 (N_4765,N_4419,N_4313);
or U4766 (N_4766,N_4298,N_4329);
and U4767 (N_4767,N_4050,N_4462);
nor U4768 (N_4768,N_4387,N_4420);
nor U4769 (N_4769,N_4244,N_4421);
nand U4770 (N_4770,N_4286,N_4331);
or U4771 (N_4771,N_4476,N_4416);
and U4772 (N_4772,N_4297,N_4368);
or U4773 (N_4773,N_4222,N_4485);
nand U4774 (N_4774,N_4059,N_4043);
or U4775 (N_4775,N_4021,N_4319);
and U4776 (N_4776,N_4117,N_4006);
or U4777 (N_4777,N_4221,N_4218);
and U4778 (N_4778,N_4216,N_4367);
nand U4779 (N_4779,N_4334,N_4215);
nor U4780 (N_4780,N_4129,N_4361);
nor U4781 (N_4781,N_4186,N_4022);
or U4782 (N_4782,N_4191,N_4454);
and U4783 (N_4783,N_4349,N_4263);
nand U4784 (N_4784,N_4006,N_4292);
or U4785 (N_4785,N_4196,N_4060);
nor U4786 (N_4786,N_4308,N_4460);
nand U4787 (N_4787,N_4220,N_4056);
or U4788 (N_4788,N_4185,N_4476);
or U4789 (N_4789,N_4202,N_4498);
and U4790 (N_4790,N_4219,N_4360);
nand U4791 (N_4791,N_4428,N_4172);
nor U4792 (N_4792,N_4460,N_4497);
and U4793 (N_4793,N_4283,N_4277);
or U4794 (N_4794,N_4165,N_4368);
nand U4795 (N_4795,N_4021,N_4449);
or U4796 (N_4796,N_4055,N_4431);
nor U4797 (N_4797,N_4447,N_4069);
or U4798 (N_4798,N_4439,N_4405);
and U4799 (N_4799,N_4064,N_4230);
or U4800 (N_4800,N_4008,N_4064);
nor U4801 (N_4801,N_4289,N_4361);
nor U4802 (N_4802,N_4218,N_4148);
nor U4803 (N_4803,N_4332,N_4067);
or U4804 (N_4804,N_4302,N_4421);
xor U4805 (N_4805,N_4494,N_4056);
and U4806 (N_4806,N_4463,N_4174);
and U4807 (N_4807,N_4292,N_4232);
nand U4808 (N_4808,N_4350,N_4198);
and U4809 (N_4809,N_4493,N_4223);
and U4810 (N_4810,N_4049,N_4292);
nor U4811 (N_4811,N_4422,N_4038);
nand U4812 (N_4812,N_4125,N_4007);
nor U4813 (N_4813,N_4372,N_4207);
or U4814 (N_4814,N_4132,N_4099);
and U4815 (N_4815,N_4356,N_4121);
nand U4816 (N_4816,N_4106,N_4303);
and U4817 (N_4817,N_4445,N_4023);
and U4818 (N_4818,N_4112,N_4272);
and U4819 (N_4819,N_4145,N_4202);
nand U4820 (N_4820,N_4468,N_4317);
and U4821 (N_4821,N_4135,N_4236);
or U4822 (N_4822,N_4015,N_4236);
or U4823 (N_4823,N_4310,N_4384);
or U4824 (N_4824,N_4007,N_4255);
nor U4825 (N_4825,N_4065,N_4152);
nor U4826 (N_4826,N_4493,N_4125);
or U4827 (N_4827,N_4357,N_4149);
nand U4828 (N_4828,N_4246,N_4296);
or U4829 (N_4829,N_4011,N_4332);
and U4830 (N_4830,N_4245,N_4099);
and U4831 (N_4831,N_4406,N_4139);
nor U4832 (N_4832,N_4371,N_4384);
and U4833 (N_4833,N_4040,N_4431);
nand U4834 (N_4834,N_4422,N_4418);
or U4835 (N_4835,N_4264,N_4142);
or U4836 (N_4836,N_4026,N_4005);
and U4837 (N_4837,N_4112,N_4498);
nand U4838 (N_4838,N_4300,N_4188);
or U4839 (N_4839,N_4035,N_4115);
or U4840 (N_4840,N_4472,N_4051);
or U4841 (N_4841,N_4061,N_4252);
nand U4842 (N_4842,N_4185,N_4044);
nand U4843 (N_4843,N_4312,N_4342);
or U4844 (N_4844,N_4114,N_4063);
and U4845 (N_4845,N_4152,N_4349);
xor U4846 (N_4846,N_4398,N_4193);
and U4847 (N_4847,N_4350,N_4223);
or U4848 (N_4848,N_4031,N_4043);
nor U4849 (N_4849,N_4275,N_4233);
and U4850 (N_4850,N_4382,N_4017);
nand U4851 (N_4851,N_4058,N_4298);
and U4852 (N_4852,N_4082,N_4381);
and U4853 (N_4853,N_4361,N_4405);
nor U4854 (N_4854,N_4187,N_4263);
nor U4855 (N_4855,N_4282,N_4124);
or U4856 (N_4856,N_4329,N_4172);
nor U4857 (N_4857,N_4160,N_4496);
or U4858 (N_4858,N_4316,N_4300);
or U4859 (N_4859,N_4202,N_4420);
nor U4860 (N_4860,N_4285,N_4132);
nand U4861 (N_4861,N_4412,N_4131);
or U4862 (N_4862,N_4263,N_4005);
nand U4863 (N_4863,N_4342,N_4346);
or U4864 (N_4864,N_4347,N_4472);
nand U4865 (N_4865,N_4206,N_4413);
and U4866 (N_4866,N_4244,N_4214);
or U4867 (N_4867,N_4383,N_4431);
and U4868 (N_4868,N_4120,N_4396);
or U4869 (N_4869,N_4478,N_4238);
nand U4870 (N_4870,N_4278,N_4470);
nor U4871 (N_4871,N_4199,N_4258);
and U4872 (N_4872,N_4173,N_4387);
and U4873 (N_4873,N_4428,N_4306);
and U4874 (N_4874,N_4423,N_4149);
or U4875 (N_4875,N_4085,N_4070);
nand U4876 (N_4876,N_4316,N_4126);
nand U4877 (N_4877,N_4135,N_4481);
nand U4878 (N_4878,N_4287,N_4191);
nor U4879 (N_4879,N_4248,N_4105);
nand U4880 (N_4880,N_4498,N_4334);
xor U4881 (N_4881,N_4190,N_4398);
or U4882 (N_4882,N_4025,N_4488);
nand U4883 (N_4883,N_4300,N_4359);
and U4884 (N_4884,N_4410,N_4312);
or U4885 (N_4885,N_4427,N_4368);
nor U4886 (N_4886,N_4392,N_4329);
nand U4887 (N_4887,N_4040,N_4180);
nand U4888 (N_4888,N_4437,N_4317);
nand U4889 (N_4889,N_4164,N_4319);
or U4890 (N_4890,N_4194,N_4378);
or U4891 (N_4891,N_4227,N_4478);
or U4892 (N_4892,N_4057,N_4165);
nor U4893 (N_4893,N_4126,N_4247);
nand U4894 (N_4894,N_4065,N_4069);
nor U4895 (N_4895,N_4066,N_4235);
or U4896 (N_4896,N_4411,N_4139);
nor U4897 (N_4897,N_4095,N_4315);
and U4898 (N_4898,N_4013,N_4206);
or U4899 (N_4899,N_4241,N_4239);
or U4900 (N_4900,N_4164,N_4082);
and U4901 (N_4901,N_4008,N_4046);
nand U4902 (N_4902,N_4307,N_4012);
or U4903 (N_4903,N_4324,N_4265);
nand U4904 (N_4904,N_4099,N_4181);
and U4905 (N_4905,N_4074,N_4493);
and U4906 (N_4906,N_4422,N_4145);
and U4907 (N_4907,N_4005,N_4366);
and U4908 (N_4908,N_4402,N_4252);
nor U4909 (N_4909,N_4412,N_4369);
and U4910 (N_4910,N_4112,N_4278);
and U4911 (N_4911,N_4381,N_4452);
nor U4912 (N_4912,N_4023,N_4169);
nand U4913 (N_4913,N_4379,N_4250);
and U4914 (N_4914,N_4296,N_4187);
nor U4915 (N_4915,N_4137,N_4093);
or U4916 (N_4916,N_4263,N_4134);
and U4917 (N_4917,N_4290,N_4027);
nand U4918 (N_4918,N_4440,N_4404);
xor U4919 (N_4919,N_4061,N_4382);
nand U4920 (N_4920,N_4016,N_4220);
or U4921 (N_4921,N_4201,N_4307);
nor U4922 (N_4922,N_4420,N_4291);
nor U4923 (N_4923,N_4187,N_4071);
or U4924 (N_4924,N_4015,N_4182);
nand U4925 (N_4925,N_4048,N_4098);
nor U4926 (N_4926,N_4285,N_4296);
nor U4927 (N_4927,N_4199,N_4274);
or U4928 (N_4928,N_4243,N_4076);
nand U4929 (N_4929,N_4226,N_4478);
nand U4930 (N_4930,N_4348,N_4262);
xor U4931 (N_4931,N_4228,N_4041);
and U4932 (N_4932,N_4264,N_4155);
or U4933 (N_4933,N_4319,N_4083);
or U4934 (N_4934,N_4437,N_4037);
nand U4935 (N_4935,N_4319,N_4165);
nor U4936 (N_4936,N_4168,N_4197);
or U4937 (N_4937,N_4295,N_4212);
nand U4938 (N_4938,N_4200,N_4424);
and U4939 (N_4939,N_4404,N_4432);
and U4940 (N_4940,N_4036,N_4378);
or U4941 (N_4941,N_4243,N_4366);
or U4942 (N_4942,N_4465,N_4123);
or U4943 (N_4943,N_4456,N_4059);
or U4944 (N_4944,N_4213,N_4021);
nor U4945 (N_4945,N_4237,N_4428);
and U4946 (N_4946,N_4484,N_4192);
xnor U4947 (N_4947,N_4096,N_4072);
nor U4948 (N_4948,N_4067,N_4170);
nand U4949 (N_4949,N_4025,N_4151);
nand U4950 (N_4950,N_4281,N_4053);
nor U4951 (N_4951,N_4063,N_4268);
and U4952 (N_4952,N_4144,N_4169);
and U4953 (N_4953,N_4042,N_4116);
or U4954 (N_4954,N_4046,N_4343);
or U4955 (N_4955,N_4273,N_4489);
or U4956 (N_4956,N_4339,N_4471);
and U4957 (N_4957,N_4449,N_4482);
or U4958 (N_4958,N_4256,N_4412);
and U4959 (N_4959,N_4211,N_4266);
and U4960 (N_4960,N_4340,N_4387);
or U4961 (N_4961,N_4102,N_4088);
or U4962 (N_4962,N_4220,N_4232);
or U4963 (N_4963,N_4327,N_4328);
nor U4964 (N_4964,N_4088,N_4201);
and U4965 (N_4965,N_4406,N_4116);
nor U4966 (N_4966,N_4345,N_4339);
and U4967 (N_4967,N_4401,N_4094);
nor U4968 (N_4968,N_4342,N_4308);
or U4969 (N_4969,N_4085,N_4406);
or U4970 (N_4970,N_4010,N_4137);
nand U4971 (N_4971,N_4086,N_4156);
nor U4972 (N_4972,N_4002,N_4390);
and U4973 (N_4973,N_4498,N_4492);
or U4974 (N_4974,N_4101,N_4431);
nor U4975 (N_4975,N_4303,N_4035);
nor U4976 (N_4976,N_4160,N_4019);
nor U4977 (N_4977,N_4421,N_4094);
and U4978 (N_4978,N_4310,N_4386);
nor U4979 (N_4979,N_4214,N_4491);
nand U4980 (N_4980,N_4020,N_4101);
or U4981 (N_4981,N_4211,N_4282);
nor U4982 (N_4982,N_4290,N_4337);
or U4983 (N_4983,N_4480,N_4290);
and U4984 (N_4984,N_4193,N_4344);
nand U4985 (N_4985,N_4054,N_4374);
nor U4986 (N_4986,N_4079,N_4001);
nor U4987 (N_4987,N_4183,N_4174);
or U4988 (N_4988,N_4015,N_4316);
and U4989 (N_4989,N_4040,N_4031);
or U4990 (N_4990,N_4085,N_4191);
or U4991 (N_4991,N_4175,N_4216);
nor U4992 (N_4992,N_4485,N_4476);
nand U4993 (N_4993,N_4409,N_4201);
or U4994 (N_4994,N_4157,N_4324);
nand U4995 (N_4995,N_4315,N_4326);
nor U4996 (N_4996,N_4080,N_4146);
nor U4997 (N_4997,N_4001,N_4350);
or U4998 (N_4998,N_4423,N_4063);
and U4999 (N_4999,N_4165,N_4135);
nand UO_0 (O_0,N_4892,N_4860);
nand UO_1 (O_1,N_4603,N_4730);
nand UO_2 (O_2,N_4593,N_4885);
and UO_3 (O_3,N_4504,N_4675);
nand UO_4 (O_4,N_4941,N_4822);
and UO_5 (O_5,N_4738,N_4797);
or UO_6 (O_6,N_4563,N_4930);
nor UO_7 (O_7,N_4680,N_4894);
and UO_8 (O_8,N_4685,N_4615);
or UO_9 (O_9,N_4670,N_4819);
or UO_10 (O_10,N_4678,N_4577);
and UO_11 (O_11,N_4608,N_4722);
nor UO_12 (O_12,N_4996,N_4572);
nand UO_13 (O_13,N_4693,N_4828);
or UO_14 (O_14,N_4728,N_4858);
or UO_15 (O_15,N_4729,N_4787);
or UO_16 (O_16,N_4855,N_4599);
and UO_17 (O_17,N_4672,N_4947);
or UO_18 (O_18,N_4959,N_4699);
and UO_19 (O_19,N_4545,N_4781);
and UO_20 (O_20,N_4803,N_4743);
nand UO_21 (O_21,N_4674,N_4869);
or UO_22 (O_22,N_4798,N_4557);
nand UO_23 (O_23,N_4978,N_4689);
or UO_24 (O_24,N_4814,N_4840);
and UO_25 (O_25,N_4914,N_4757);
nor UO_26 (O_26,N_4835,N_4758);
nor UO_27 (O_27,N_4724,N_4910);
nand UO_28 (O_28,N_4922,N_4886);
and UO_29 (O_29,N_4592,N_4986);
and UO_30 (O_30,N_4641,N_4660);
or UO_31 (O_31,N_4772,N_4801);
nor UO_32 (O_32,N_4839,N_4673);
or UO_33 (O_33,N_4715,N_4813);
nand UO_34 (O_34,N_4541,N_4834);
nand UO_35 (O_35,N_4774,N_4569);
nand UO_36 (O_36,N_4513,N_4568);
or UO_37 (O_37,N_4850,N_4980);
and UO_38 (O_38,N_4697,N_4826);
and UO_39 (O_39,N_4921,N_4979);
nand UO_40 (O_40,N_4887,N_4558);
nand UO_41 (O_41,N_4765,N_4923);
and UO_42 (O_42,N_4856,N_4879);
or UO_43 (O_43,N_4842,N_4529);
nand UO_44 (O_44,N_4695,N_4939);
nor UO_45 (O_45,N_4851,N_4708);
nor UO_46 (O_46,N_4588,N_4793);
and UO_47 (O_47,N_4824,N_4548);
or UO_48 (O_48,N_4610,N_4741);
nand UO_49 (O_49,N_4812,N_4877);
nand UO_50 (O_50,N_4852,N_4817);
nand UO_51 (O_51,N_4517,N_4586);
nor UO_52 (O_52,N_4811,N_4882);
or UO_53 (O_53,N_4790,N_4677);
or UO_54 (O_54,N_4861,N_4655);
nor UO_55 (O_55,N_4833,N_4507);
and UO_56 (O_56,N_4760,N_4888);
nor UO_57 (O_57,N_4521,N_4849);
nand UO_58 (O_58,N_4759,N_4536);
nand UO_59 (O_59,N_4827,N_4512);
nor UO_60 (O_60,N_4532,N_4909);
and UO_61 (O_61,N_4755,N_4717);
nand UO_62 (O_62,N_4648,N_4580);
nor UO_63 (O_63,N_4546,N_4795);
nor UO_64 (O_64,N_4962,N_4775);
or UO_65 (O_65,N_4684,N_4666);
and UO_66 (O_66,N_4725,N_4987);
nand UO_67 (O_67,N_4989,N_4613);
and UO_68 (O_68,N_4727,N_4919);
or UO_69 (O_69,N_4515,N_4720);
and UO_70 (O_70,N_4714,N_4686);
nor UO_71 (O_71,N_4734,N_4762);
or UO_72 (O_72,N_4590,N_4881);
nor UO_73 (O_73,N_4898,N_4969);
or UO_74 (O_74,N_4607,N_4912);
or UO_75 (O_75,N_4671,N_4531);
and UO_76 (O_76,N_4573,N_4505);
and UO_77 (O_77,N_4927,N_4631);
nand UO_78 (O_78,N_4705,N_4584);
and UO_79 (O_79,N_4838,N_4668);
nand UO_80 (O_80,N_4846,N_4810);
nand UO_81 (O_81,N_4773,N_4944);
and UO_82 (O_82,N_4973,N_4691);
and UO_83 (O_83,N_4506,N_4538);
and UO_84 (O_84,N_4514,N_4763);
nand UO_85 (O_85,N_4650,N_4816);
and UO_86 (O_86,N_4931,N_4832);
and UO_87 (O_87,N_4552,N_4634);
nor UO_88 (O_88,N_4736,N_4562);
xor UO_89 (O_89,N_4530,N_4777);
and UO_90 (O_90,N_4591,N_4518);
nand UO_91 (O_91,N_4988,N_4718);
or UO_92 (O_92,N_4690,N_4875);
and UO_93 (O_93,N_4768,N_4957);
nor UO_94 (O_94,N_4873,N_4761);
or UO_95 (O_95,N_4564,N_4742);
nor UO_96 (O_96,N_4915,N_4924);
nor UO_97 (O_97,N_4534,N_4965);
nor UO_98 (O_98,N_4786,N_4503);
or UO_99 (O_99,N_4789,N_4874);
or UO_100 (O_100,N_4891,N_4982);
nor UO_101 (O_101,N_4556,N_4770);
or UO_102 (O_102,N_4866,N_4616);
nand UO_103 (O_103,N_4731,N_4703);
nor UO_104 (O_104,N_4566,N_4639);
or UO_105 (O_105,N_4792,N_4997);
nand UO_106 (O_106,N_4600,N_4948);
nand UO_107 (O_107,N_4527,N_4756);
nor UO_108 (O_108,N_4553,N_4779);
and UO_109 (O_109,N_4776,N_4745);
xor UO_110 (O_110,N_4565,N_4544);
nor UO_111 (O_111,N_4589,N_4806);
and UO_112 (O_112,N_4519,N_4716);
nand UO_113 (O_113,N_4665,N_4872);
nor UO_114 (O_114,N_4526,N_4999);
or UO_115 (O_115,N_4904,N_4637);
and UO_116 (O_116,N_4954,N_4604);
nor UO_117 (O_117,N_4669,N_4896);
nor UO_118 (O_118,N_4707,N_4913);
nor UO_119 (O_119,N_4878,N_4901);
and UO_120 (O_120,N_4642,N_4946);
or UO_121 (O_121,N_4619,N_4895);
and UO_122 (O_122,N_4953,N_4547);
and UO_123 (O_123,N_4737,N_4949);
and UO_124 (O_124,N_4870,N_4719);
or UO_125 (O_125,N_4581,N_4543);
nor UO_126 (O_126,N_4994,N_4733);
or UO_127 (O_127,N_4884,N_4653);
or UO_128 (O_128,N_4929,N_4501);
xnor UO_129 (O_129,N_4542,N_4845);
nand UO_130 (O_130,N_4934,N_4754);
or UO_131 (O_131,N_4995,N_4985);
nor UO_132 (O_132,N_4511,N_4682);
nand UO_133 (O_133,N_4570,N_4907);
nor UO_134 (O_134,N_4862,N_4975);
or UO_135 (O_135,N_4847,N_4751);
or UO_136 (O_136,N_4778,N_4611);
and UO_137 (O_137,N_4902,N_4630);
nor UO_138 (O_138,N_4906,N_4749);
xor UO_139 (O_139,N_4576,N_4926);
or UO_140 (O_140,N_4594,N_4694);
and UO_141 (O_141,N_4918,N_4702);
nor UO_142 (O_142,N_4876,N_4711);
nand UO_143 (O_143,N_4522,N_4952);
and UO_144 (O_144,N_4647,N_4739);
or UO_145 (O_145,N_4917,N_4807);
or UO_146 (O_146,N_4706,N_4785);
nor UO_147 (O_147,N_4533,N_4900);
nand UO_148 (O_148,N_4516,N_4945);
nand UO_149 (O_149,N_4618,N_4747);
and UO_150 (O_150,N_4823,N_4614);
or UO_151 (O_151,N_4574,N_4897);
and UO_152 (O_152,N_4925,N_4808);
xor UO_153 (O_153,N_4667,N_4632);
and UO_154 (O_154,N_4649,N_4723);
xor UO_155 (O_155,N_4967,N_4943);
nor UO_156 (O_156,N_4899,N_4679);
nor UO_157 (O_157,N_4571,N_4645);
nor UO_158 (O_158,N_4753,N_4783);
nor UO_159 (O_159,N_4990,N_4796);
nor UO_160 (O_160,N_4601,N_4799);
nand UO_161 (O_161,N_4889,N_4830);
nand UO_162 (O_162,N_4968,N_4628);
xnor UO_163 (O_163,N_4585,N_4550);
and UO_164 (O_164,N_4579,N_4502);
and UO_165 (O_165,N_4712,N_4865);
nor UO_166 (O_166,N_4829,N_4942);
nor UO_167 (O_167,N_4750,N_4843);
or UO_168 (O_168,N_4582,N_4976);
nand UO_169 (O_169,N_4520,N_4800);
and UO_170 (O_170,N_4890,N_4936);
and UO_171 (O_171,N_4549,N_4864);
or UO_172 (O_172,N_4597,N_4971);
nor UO_173 (O_173,N_4651,N_4932);
or UO_174 (O_174,N_4525,N_4744);
nor UO_175 (O_175,N_4509,N_4868);
and UO_176 (O_176,N_4908,N_4788);
nor UO_177 (O_177,N_4626,N_4794);
xor UO_178 (O_178,N_4983,N_4821);
and UO_179 (O_179,N_4940,N_4629);
or UO_180 (O_180,N_4937,N_4960);
or UO_181 (O_181,N_4784,N_4804);
nor UO_182 (O_182,N_4955,N_4848);
nand UO_183 (O_183,N_4539,N_4578);
nor UO_184 (O_184,N_4559,N_4998);
nor UO_185 (O_185,N_4583,N_4735);
or UO_186 (O_186,N_4625,N_4598);
or UO_187 (O_187,N_4646,N_4853);
and UO_188 (O_188,N_4740,N_4698);
nand UO_189 (O_189,N_4508,N_4688);
or UO_190 (O_190,N_4620,N_4748);
and UO_191 (O_191,N_4713,N_4654);
and UO_192 (O_192,N_4606,N_4836);
nor UO_193 (O_193,N_4791,N_4841);
nand UO_194 (O_194,N_4818,N_4658);
nor UO_195 (O_195,N_4867,N_4766);
nand UO_196 (O_196,N_4681,N_4732);
or UO_197 (O_197,N_4704,N_4863);
or UO_198 (O_198,N_4709,N_4602);
or UO_199 (O_199,N_4524,N_4561);
nand UO_200 (O_200,N_4981,N_4809);
nor UO_201 (O_201,N_4664,N_4991);
or UO_202 (O_202,N_4933,N_4974);
nor UO_203 (O_203,N_4780,N_4659);
nor UO_204 (O_204,N_4764,N_4961);
nand UO_205 (O_205,N_4871,N_4644);
or UO_206 (O_206,N_4710,N_4609);
and UO_207 (O_207,N_4595,N_4964);
nor UO_208 (O_208,N_4657,N_4640);
and UO_209 (O_209,N_4956,N_4963);
or UO_210 (O_210,N_4950,N_4831);
nand UO_211 (O_211,N_4893,N_4771);
nor UO_212 (O_212,N_4883,N_4938);
and UO_213 (O_213,N_4555,N_4928);
or UO_214 (O_214,N_4920,N_4551);
nand UO_215 (O_215,N_4605,N_4854);
or UO_216 (O_216,N_4916,N_4769);
or UO_217 (O_217,N_4635,N_4903);
nand UO_218 (O_218,N_4746,N_4623);
or UO_219 (O_219,N_4540,N_4627);
and UO_220 (O_220,N_4567,N_4596);
nor UO_221 (O_221,N_4656,N_4621);
nand UO_222 (O_222,N_4683,N_4970);
and UO_223 (O_223,N_4805,N_4844);
nand UO_224 (O_224,N_4837,N_4638);
or UO_225 (O_225,N_4624,N_4663);
and UO_226 (O_226,N_4701,N_4984);
and UO_227 (O_227,N_4935,N_4700);
or UO_228 (O_228,N_4951,N_4972);
nor UO_229 (O_229,N_4911,N_4687);
or UO_230 (O_230,N_4652,N_4528);
nor UO_231 (O_231,N_4575,N_4802);
nand UO_232 (O_232,N_4752,N_4622);
nand UO_233 (O_233,N_4782,N_4993);
or UO_234 (O_234,N_4857,N_4633);
or UO_235 (O_235,N_4696,N_4587);
nand UO_236 (O_236,N_4820,N_4560);
nand UO_237 (O_237,N_4815,N_4636);
nor UO_238 (O_238,N_4966,N_4617);
nand UO_239 (O_239,N_4535,N_4767);
or UO_240 (O_240,N_4977,N_4661);
nand UO_241 (O_241,N_4523,N_4676);
and UO_242 (O_242,N_4859,N_4500);
nand UO_243 (O_243,N_4662,N_4554);
nor UO_244 (O_244,N_4905,N_4692);
or UO_245 (O_245,N_4992,N_4721);
nor UO_246 (O_246,N_4825,N_4958);
nand UO_247 (O_247,N_4510,N_4612);
and UO_248 (O_248,N_4880,N_4726);
or UO_249 (O_249,N_4643,N_4537);
or UO_250 (O_250,N_4919,N_4847);
nand UO_251 (O_251,N_4767,N_4519);
or UO_252 (O_252,N_4798,N_4610);
and UO_253 (O_253,N_4656,N_4549);
nand UO_254 (O_254,N_4731,N_4854);
nand UO_255 (O_255,N_4534,N_4976);
nand UO_256 (O_256,N_4768,N_4653);
or UO_257 (O_257,N_4996,N_4718);
or UO_258 (O_258,N_4526,N_4667);
and UO_259 (O_259,N_4793,N_4723);
nand UO_260 (O_260,N_4512,N_4688);
nor UO_261 (O_261,N_4852,N_4743);
or UO_262 (O_262,N_4654,N_4740);
and UO_263 (O_263,N_4667,N_4708);
or UO_264 (O_264,N_4918,N_4837);
or UO_265 (O_265,N_4858,N_4761);
nor UO_266 (O_266,N_4762,N_4733);
nor UO_267 (O_267,N_4960,N_4756);
and UO_268 (O_268,N_4870,N_4704);
and UO_269 (O_269,N_4913,N_4910);
nor UO_270 (O_270,N_4953,N_4724);
or UO_271 (O_271,N_4962,N_4974);
nor UO_272 (O_272,N_4709,N_4566);
nand UO_273 (O_273,N_4834,N_4699);
or UO_274 (O_274,N_4820,N_4798);
nand UO_275 (O_275,N_4718,N_4744);
nor UO_276 (O_276,N_4617,N_4561);
nor UO_277 (O_277,N_4959,N_4509);
nor UO_278 (O_278,N_4673,N_4830);
and UO_279 (O_279,N_4507,N_4881);
nor UO_280 (O_280,N_4977,N_4935);
nand UO_281 (O_281,N_4832,N_4740);
and UO_282 (O_282,N_4506,N_4999);
or UO_283 (O_283,N_4995,N_4573);
or UO_284 (O_284,N_4520,N_4572);
and UO_285 (O_285,N_4519,N_4976);
or UO_286 (O_286,N_4621,N_4974);
xor UO_287 (O_287,N_4583,N_4868);
and UO_288 (O_288,N_4569,N_4843);
or UO_289 (O_289,N_4916,N_4639);
nand UO_290 (O_290,N_4979,N_4657);
nand UO_291 (O_291,N_4501,N_4893);
xnor UO_292 (O_292,N_4816,N_4596);
and UO_293 (O_293,N_4543,N_4937);
nand UO_294 (O_294,N_4593,N_4630);
and UO_295 (O_295,N_4943,N_4807);
nor UO_296 (O_296,N_4973,N_4611);
nor UO_297 (O_297,N_4668,N_4573);
and UO_298 (O_298,N_4934,N_4867);
nor UO_299 (O_299,N_4608,N_4688);
and UO_300 (O_300,N_4581,N_4672);
or UO_301 (O_301,N_4658,N_4737);
nor UO_302 (O_302,N_4681,N_4535);
and UO_303 (O_303,N_4600,N_4938);
nand UO_304 (O_304,N_4827,N_4580);
nand UO_305 (O_305,N_4997,N_4633);
or UO_306 (O_306,N_4689,N_4950);
or UO_307 (O_307,N_4663,N_4543);
or UO_308 (O_308,N_4831,N_4806);
nor UO_309 (O_309,N_4951,N_4814);
or UO_310 (O_310,N_4616,N_4830);
nor UO_311 (O_311,N_4588,N_4769);
nor UO_312 (O_312,N_4925,N_4672);
and UO_313 (O_313,N_4642,N_4658);
nand UO_314 (O_314,N_4761,N_4870);
and UO_315 (O_315,N_4672,N_4792);
and UO_316 (O_316,N_4901,N_4569);
nor UO_317 (O_317,N_4585,N_4844);
nor UO_318 (O_318,N_4964,N_4739);
nand UO_319 (O_319,N_4677,N_4927);
or UO_320 (O_320,N_4671,N_4771);
and UO_321 (O_321,N_4658,N_4742);
nand UO_322 (O_322,N_4706,N_4573);
nor UO_323 (O_323,N_4727,N_4833);
nor UO_324 (O_324,N_4562,N_4529);
and UO_325 (O_325,N_4727,N_4584);
nor UO_326 (O_326,N_4833,N_4789);
nand UO_327 (O_327,N_4511,N_4547);
or UO_328 (O_328,N_4970,N_4868);
and UO_329 (O_329,N_4746,N_4978);
nand UO_330 (O_330,N_4612,N_4795);
nor UO_331 (O_331,N_4737,N_4909);
and UO_332 (O_332,N_4968,N_4932);
or UO_333 (O_333,N_4647,N_4523);
nor UO_334 (O_334,N_4560,N_4605);
nor UO_335 (O_335,N_4838,N_4761);
or UO_336 (O_336,N_4581,N_4580);
nor UO_337 (O_337,N_4861,N_4719);
nand UO_338 (O_338,N_4703,N_4747);
or UO_339 (O_339,N_4593,N_4856);
nand UO_340 (O_340,N_4527,N_4907);
and UO_341 (O_341,N_4589,N_4768);
and UO_342 (O_342,N_4781,N_4621);
or UO_343 (O_343,N_4966,N_4534);
or UO_344 (O_344,N_4851,N_4894);
nand UO_345 (O_345,N_4550,N_4539);
nand UO_346 (O_346,N_4934,N_4548);
nand UO_347 (O_347,N_4798,N_4857);
nand UO_348 (O_348,N_4664,N_4768);
nor UO_349 (O_349,N_4746,N_4836);
and UO_350 (O_350,N_4549,N_4607);
nor UO_351 (O_351,N_4925,N_4759);
and UO_352 (O_352,N_4931,N_4683);
and UO_353 (O_353,N_4948,N_4526);
nor UO_354 (O_354,N_4596,N_4531);
or UO_355 (O_355,N_4669,N_4544);
or UO_356 (O_356,N_4882,N_4641);
xor UO_357 (O_357,N_4917,N_4752);
or UO_358 (O_358,N_4978,N_4775);
xnor UO_359 (O_359,N_4699,N_4747);
or UO_360 (O_360,N_4720,N_4529);
and UO_361 (O_361,N_4725,N_4788);
nor UO_362 (O_362,N_4714,N_4514);
and UO_363 (O_363,N_4996,N_4599);
xor UO_364 (O_364,N_4995,N_4702);
and UO_365 (O_365,N_4850,N_4851);
and UO_366 (O_366,N_4606,N_4847);
or UO_367 (O_367,N_4859,N_4592);
nand UO_368 (O_368,N_4502,N_4711);
or UO_369 (O_369,N_4765,N_4796);
and UO_370 (O_370,N_4771,N_4764);
and UO_371 (O_371,N_4937,N_4570);
nor UO_372 (O_372,N_4510,N_4941);
nand UO_373 (O_373,N_4917,N_4857);
or UO_374 (O_374,N_4701,N_4576);
nor UO_375 (O_375,N_4512,N_4873);
nand UO_376 (O_376,N_4692,N_4530);
nor UO_377 (O_377,N_4569,N_4880);
nor UO_378 (O_378,N_4639,N_4719);
and UO_379 (O_379,N_4786,N_4779);
nand UO_380 (O_380,N_4591,N_4863);
and UO_381 (O_381,N_4982,N_4871);
nor UO_382 (O_382,N_4571,N_4657);
and UO_383 (O_383,N_4907,N_4868);
or UO_384 (O_384,N_4893,N_4658);
or UO_385 (O_385,N_4773,N_4601);
nor UO_386 (O_386,N_4699,N_4582);
or UO_387 (O_387,N_4500,N_4745);
and UO_388 (O_388,N_4633,N_4963);
xor UO_389 (O_389,N_4644,N_4710);
and UO_390 (O_390,N_4540,N_4848);
and UO_391 (O_391,N_4929,N_4755);
nor UO_392 (O_392,N_4931,N_4905);
nand UO_393 (O_393,N_4931,N_4771);
nor UO_394 (O_394,N_4815,N_4932);
nand UO_395 (O_395,N_4982,N_4537);
nand UO_396 (O_396,N_4991,N_4533);
or UO_397 (O_397,N_4799,N_4506);
nor UO_398 (O_398,N_4898,N_4821);
or UO_399 (O_399,N_4671,N_4942);
and UO_400 (O_400,N_4813,N_4570);
and UO_401 (O_401,N_4818,N_4919);
xor UO_402 (O_402,N_4789,N_4958);
nor UO_403 (O_403,N_4567,N_4800);
and UO_404 (O_404,N_4947,N_4896);
or UO_405 (O_405,N_4683,N_4514);
or UO_406 (O_406,N_4865,N_4693);
nand UO_407 (O_407,N_4870,N_4722);
nand UO_408 (O_408,N_4513,N_4886);
nand UO_409 (O_409,N_4647,N_4798);
nor UO_410 (O_410,N_4621,N_4561);
nand UO_411 (O_411,N_4860,N_4703);
and UO_412 (O_412,N_4684,N_4571);
nand UO_413 (O_413,N_4592,N_4667);
or UO_414 (O_414,N_4977,N_4822);
or UO_415 (O_415,N_4846,N_4818);
nor UO_416 (O_416,N_4600,N_4815);
nand UO_417 (O_417,N_4867,N_4663);
and UO_418 (O_418,N_4659,N_4808);
nand UO_419 (O_419,N_4602,N_4604);
or UO_420 (O_420,N_4950,N_4912);
and UO_421 (O_421,N_4600,N_4864);
nand UO_422 (O_422,N_4512,N_4851);
nor UO_423 (O_423,N_4553,N_4552);
nor UO_424 (O_424,N_4672,N_4864);
nand UO_425 (O_425,N_4970,N_4781);
nand UO_426 (O_426,N_4757,N_4982);
nor UO_427 (O_427,N_4626,N_4891);
nand UO_428 (O_428,N_4523,N_4934);
xnor UO_429 (O_429,N_4825,N_4507);
nand UO_430 (O_430,N_4517,N_4606);
and UO_431 (O_431,N_4840,N_4569);
nand UO_432 (O_432,N_4663,N_4854);
or UO_433 (O_433,N_4701,N_4980);
and UO_434 (O_434,N_4999,N_4548);
and UO_435 (O_435,N_4958,N_4884);
or UO_436 (O_436,N_4713,N_4875);
nand UO_437 (O_437,N_4958,N_4721);
and UO_438 (O_438,N_4658,N_4950);
nand UO_439 (O_439,N_4876,N_4602);
nand UO_440 (O_440,N_4834,N_4943);
nand UO_441 (O_441,N_4524,N_4644);
and UO_442 (O_442,N_4751,N_4864);
or UO_443 (O_443,N_4537,N_4704);
or UO_444 (O_444,N_4890,N_4597);
or UO_445 (O_445,N_4908,N_4644);
nor UO_446 (O_446,N_4530,N_4895);
nor UO_447 (O_447,N_4936,N_4648);
nand UO_448 (O_448,N_4747,N_4644);
and UO_449 (O_449,N_4958,N_4800);
and UO_450 (O_450,N_4987,N_4834);
or UO_451 (O_451,N_4883,N_4673);
nor UO_452 (O_452,N_4664,N_4920);
or UO_453 (O_453,N_4643,N_4718);
xnor UO_454 (O_454,N_4712,N_4734);
nand UO_455 (O_455,N_4771,N_4938);
nand UO_456 (O_456,N_4554,N_4846);
and UO_457 (O_457,N_4641,N_4535);
nand UO_458 (O_458,N_4685,N_4776);
nand UO_459 (O_459,N_4651,N_4735);
and UO_460 (O_460,N_4975,N_4940);
or UO_461 (O_461,N_4851,N_4550);
nor UO_462 (O_462,N_4986,N_4706);
xnor UO_463 (O_463,N_4968,N_4874);
xnor UO_464 (O_464,N_4652,N_4625);
nor UO_465 (O_465,N_4803,N_4549);
nand UO_466 (O_466,N_4508,N_4592);
nand UO_467 (O_467,N_4511,N_4895);
nand UO_468 (O_468,N_4819,N_4928);
nor UO_469 (O_469,N_4627,N_4653);
nand UO_470 (O_470,N_4890,N_4966);
nand UO_471 (O_471,N_4970,N_4778);
nor UO_472 (O_472,N_4978,N_4550);
and UO_473 (O_473,N_4754,N_4597);
nor UO_474 (O_474,N_4694,N_4689);
and UO_475 (O_475,N_4500,N_4994);
nand UO_476 (O_476,N_4531,N_4982);
nand UO_477 (O_477,N_4768,N_4619);
or UO_478 (O_478,N_4517,N_4669);
or UO_479 (O_479,N_4679,N_4693);
nand UO_480 (O_480,N_4607,N_4586);
and UO_481 (O_481,N_4993,N_4851);
nor UO_482 (O_482,N_4524,N_4761);
nand UO_483 (O_483,N_4901,N_4968);
nand UO_484 (O_484,N_4872,N_4537);
or UO_485 (O_485,N_4862,N_4574);
nand UO_486 (O_486,N_4793,N_4902);
and UO_487 (O_487,N_4772,N_4806);
nand UO_488 (O_488,N_4875,N_4857);
nor UO_489 (O_489,N_4830,N_4842);
nand UO_490 (O_490,N_4598,N_4594);
nor UO_491 (O_491,N_4776,N_4902);
nand UO_492 (O_492,N_4716,N_4988);
and UO_493 (O_493,N_4996,N_4855);
or UO_494 (O_494,N_4807,N_4513);
nand UO_495 (O_495,N_4500,N_4533);
nor UO_496 (O_496,N_4704,N_4554);
and UO_497 (O_497,N_4642,N_4552);
nor UO_498 (O_498,N_4660,N_4605);
nand UO_499 (O_499,N_4892,N_4638);
nor UO_500 (O_500,N_4876,N_4505);
or UO_501 (O_501,N_4657,N_4974);
nand UO_502 (O_502,N_4894,N_4865);
or UO_503 (O_503,N_4640,N_4923);
and UO_504 (O_504,N_4522,N_4515);
nor UO_505 (O_505,N_4546,N_4602);
nor UO_506 (O_506,N_4563,N_4533);
nand UO_507 (O_507,N_4607,N_4555);
or UO_508 (O_508,N_4725,N_4723);
nor UO_509 (O_509,N_4557,N_4661);
nor UO_510 (O_510,N_4856,N_4964);
or UO_511 (O_511,N_4907,N_4551);
nor UO_512 (O_512,N_4762,N_4893);
and UO_513 (O_513,N_4733,N_4713);
nand UO_514 (O_514,N_4730,N_4754);
nor UO_515 (O_515,N_4973,N_4672);
nor UO_516 (O_516,N_4841,N_4546);
xor UO_517 (O_517,N_4522,N_4555);
nor UO_518 (O_518,N_4649,N_4714);
nand UO_519 (O_519,N_4897,N_4586);
nand UO_520 (O_520,N_4606,N_4607);
nand UO_521 (O_521,N_4610,N_4559);
and UO_522 (O_522,N_4888,N_4613);
nand UO_523 (O_523,N_4984,N_4953);
nand UO_524 (O_524,N_4876,N_4945);
and UO_525 (O_525,N_4637,N_4542);
nor UO_526 (O_526,N_4962,N_4743);
nand UO_527 (O_527,N_4679,N_4892);
nor UO_528 (O_528,N_4501,N_4800);
and UO_529 (O_529,N_4996,N_4567);
or UO_530 (O_530,N_4922,N_4854);
or UO_531 (O_531,N_4527,N_4601);
nand UO_532 (O_532,N_4708,N_4934);
and UO_533 (O_533,N_4706,N_4664);
or UO_534 (O_534,N_4559,N_4841);
and UO_535 (O_535,N_4510,N_4750);
nand UO_536 (O_536,N_4738,N_4886);
nand UO_537 (O_537,N_4668,N_4705);
nand UO_538 (O_538,N_4979,N_4872);
xor UO_539 (O_539,N_4779,N_4574);
or UO_540 (O_540,N_4513,N_4609);
nor UO_541 (O_541,N_4769,N_4743);
and UO_542 (O_542,N_4856,N_4812);
xor UO_543 (O_543,N_4763,N_4557);
nor UO_544 (O_544,N_4999,N_4646);
or UO_545 (O_545,N_4959,N_4643);
or UO_546 (O_546,N_4810,N_4917);
and UO_547 (O_547,N_4690,N_4896);
or UO_548 (O_548,N_4871,N_4613);
xnor UO_549 (O_549,N_4594,N_4828);
nand UO_550 (O_550,N_4893,N_4727);
and UO_551 (O_551,N_4795,N_4564);
nor UO_552 (O_552,N_4984,N_4897);
and UO_553 (O_553,N_4877,N_4780);
and UO_554 (O_554,N_4699,N_4725);
nand UO_555 (O_555,N_4601,N_4666);
nor UO_556 (O_556,N_4972,N_4601);
and UO_557 (O_557,N_4790,N_4997);
or UO_558 (O_558,N_4805,N_4975);
nor UO_559 (O_559,N_4617,N_4680);
nand UO_560 (O_560,N_4577,N_4797);
nor UO_561 (O_561,N_4683,N_4879);
or UO_562 (O_562,N_4613,N_4511);
nor UO_563 (O_563,N_4858,N_4884);
nand UO_564 (O_564,N_4574,N_4981);
or UO_565 (O_565,N_4923,N_4877);
or UO_566 (O_566,N_4864,N_4838);
nor UO_567 (O_567,N_4933,N_4747);
and UO_568 (O_568,N_4556,N_4979);
nor UO_569 (O_569,N_4646,N_4847);
nor UO_570 (O_570,N_4898,N_4924);
or UO_571 (O_571,N_4565,N_4827);
nor UO_572 (O_572,N_4709,N_4584);
nand UO_573 (O_573,N_4826,N_4560);
nand UO_574 (O_574,N_4653,N_4776);
nor UO_575 (O_575,N_4659,N_4791);
nor UO_576 (O_576,N_4894,N_4693);
and UO_577 (O_577,N_4628,N_4923);
nor UO_578 (O_578,N_4777,N_4872);
nand UO_579 (O_579,N_4550,N_4943);
nand UO_580 (O_580,N_4542,N_4572);
nand UO_581 (O_581,N_4828,N_4612);
or UO_582 (O_582,N_4823,N_4865);
and UO_583 (O_583,N_4909,N_4543);
nor UO_584 (O_584,N_4526,N_4511);
nor UO_585 (O_585,N_4995,N_4831);
nor UO_586 (O_586,N_4968,N_4580);
or UO_587 (O_587,N_4511,N_4729);
nor UO_588 (O_588,N_4556,N_4811);
nor UO_589 (O_589,N_4862,N_4988);
nand UO_590 (O_590,N_4987,N_4606);
or UO_591 (O_591,N_4906,N_4878);
xnor UO_592 (O_592,N_4855,N_4578);
or UO_593 (O_593,N_4623,N_4981);
and UO_594 (O_594,N_4526,N_4665);
or UO_595 (O_595,N_4524,N_4663);
and UO_596 (O_596,N_4545,N_4619);
xor UO_597 (O_597,N_4539,N_4942);
nand UO_598 (O_598,N_4948,N_4660);
and UO_599 (O_599,N_4915,N_4613);
or UO_600 (O_600,N_4537,N_4558);
nor UO_601 (O_601,N_4912,N_4854);
nand UO_602 (O_602,N_4808,N_4568);
nor UO_603 (O_603,N_4540,N_4604);
nand UO_604 (O_604,N_4511,N_4541);
and UO_605 (O_605,N_4887,N_4503);
or UO_606 (O_606,N_4945,N_4965);
xnor UO_607 (O_607,N_4772,N_4737);
nand UO_608 (O_608,N_4940,N_4884);
nor UO_609 (O_609,N_4751,N_4555);
nand UO_610 (O_610,N_4594,N_4712);
or UO_611 (O_611,N_4975,N_4620);
and UO_612 (O_612,N_4831,N_4952);
or UO_613 (O_613,N_4661,N_4733);
and UO_614 (O_614,N_4856,N_4679);
nand UO_615 (O_615,N_4599,N_4973);
nand UO_616 (O_616,N_4647,N_4951);
nor UO_617 (O_617,N_4783,N_4825);
nand UO_618 (O_618,N_4989,N_4878);
nand UO_619 (O_619,N_4830,N_4634);
and UO_620 (O_620,N_4546,N_4783);
xnor UO_621 (O_621,N_4525,N_4796);
or UO_622 (O_622,N_4899,N_4983);
xnor UO_623 (O_623,N_4892,N_4606);
nor UO_624 (O_624,N_4989,N_4542);
and UO_625 (O_625,N_4833,N_4591);
or UO_626 (O_626,N_4923,N_4598);
nand UO_627 (O_627,N_4839,N_4606);
and UO_628 (O_628,N_4642,N_4781);
and UO_629 (O_629,N_4604,N_4655);
and UO_630 (O_630,N_4681,N_4776);
nor UO_631 (O_631,N_4542,N_4926);
nand UO_632 (O_632,N_4714,N_4532);
nand UO_633 (O_633,N_4825,N_4692);
and UO_634 (O_634,N_4703,N_4891);
and UO_635 (O_635,N_4919,N_4596);
or UO_636 (O_636,N_4954,N_4926);
nor UO_637 (O_637,N_4593,N_4760);
and UO_638 (O_638,N_4897,N_4594);
and UO_639 (O_639,N_4635,N_4890);
or UO_640 (O_640,N_4787,N_4976);
and UO_641 (O_641,N_4534,N_4933);
or UO_642 (O_642,N_4635,N_4660);
xnor UO_643 (O_643,N_4973,N_4631);
or UO_644 (O_644,N_4690,N_4564);
or UO_645 (O_645,N_4811,N_4730);
nand UO_646 (O_646,N_4633,N_4992);
nor UO_647 (O_647,N_4894,N_4904);
xnor UO_648 (O_648,N_4508,N_4721);
or UO_649 (O_649,N_4675,N_4752);
or UO_650 (O_650,N_4790,N_4513);
or UO_651 (O_651,N_4967,N_4540);
nand UO_652 (O_652,N_4897,N_4612);
and UO_653 (O_653,N_4992,N_4773);
nand UO_654 (O_654,N_4534,N_4887);
nand UO_655 (O_655,N_4775,N_4854);
nand UO_656 (O_656,N_4575,N_4883);
or UO_657 (O_657,N_4583,N_4925);
nand UO_658 (O_658,N_4765,N_4703);
nand UO_659 (O_659,N_4716,N_4846);
nand UO_660 (O_660,N_4563,N_4663);
nand UO_661 (O_661,N_4626,N_4758);
nor UO_662 (O_662,N_4894,N_4928);
nor UO_663 (O_663,N_4921,N_4699);
nand UO_664 (O_664,N_4558,N_4749);
or UO_665 (O_665,N_4712,N_4693);
nand UO_666 (O_666,N_4539,N_4697);
nand UO_667 (O_667,N_4909,N_4879);
xnor UO_668 (O_668,N_4513,N_4659);
or UO_669 (O_669,N_4885,N_4529);
nor UO_670 (O_670,N_4724,N_4872);
or UO_671 (O_671,N_4930,N_4874);
nand UO_672 (O_672,N_4945,N_4784);
or UO_673 (O_673,N_4677,N_4862);
and UO_674 (O_674,N_4946,N_4745);
nand UO_675 (O_675,N_4774,N_4647);
nor UO_676 (O_676,N_4886,N_4911);
nand UO_677 (O_677,N_4685,N_4884);
or UO_678 (O_678,N_4693,N_4624);
and UO_679 (O_679,N_4691,N_4762);
or UO_680 (O_680,N_4899,N_4904);
and UO_681 (O_681,N_4897,N_4947);
or UO_682 (O_682,N_4608,N_4872);
and UO_683 (O_683,N_4562,N_4723);
or UO_684 (O_684,N_4961,N_4802);
or UO_685 (O_685,N_4810,N_4710);
nor UO_686 (O_686,N_4950,N_4703);
xor UO_687 (O_687,N_4969,N_4704);
and UO_688 (O_688,N_4999,N_4676);
or UO_689 (O_689,N_4904,N_4728);
and UO_690 (O_690,N_4880,N_4714);
nand UO_691 (O_691,N_4685,N_4690);
and UO_692 (O_692,N_4924,N_4788);
or UO_693 (O_693,N_4768,N_4640);
nor UO_694 (O_694,N_4611,N_4541);
nor UO_695 (O_695,N_4761,N_4839);
nand UO_696 (O_696,N_4828,N_4742);
and UO_697 (O_697,N_4959,N_4809);
and UO_698 (O_698,N_4941,N_4670);
or UO_699 (O_699,N_4502,N_4653);
nand UO_700 (O_700,N_4857,N_4945);
nand UO_701 (O_701,N_4769,N_4609);
or UO_702 (O_702,N_4534,N_4814);
nor UO_703 (O_703,N_4823,N_4555);
or UO_704 (O_704,N_4866,N_4603);
nand UO_705 (O_705,N_4848,N_4976);
nor UO_706 (O_706,N_4892,N_4915);
nor UO_707 (O_707,N_4810,N_4877);
nand UO_708 (O_708,N_4809,N_4568);
or UO_709 (O_709,N_4919,N_4710);
or UO_710 (O_710,N_4630,N_4579);
and UO_711 (O_711,N_4757,N_4600);
nor UO_712 (O_712,N_4814,N_4514);
and UO_713 (O_713,N_4941,N_4825);
nand UO_714 (O_714,N_4963,N_4897);
and UO_715 (O_715,N_4608,N_4975);
or UO_716 (O_716,N_4634,N_4910);
and UO_717 (O_717,N_4738,N_4506);
or UO_718 (O_718,N_4633,N_4661);
nand UO_719 (O_719,N_4816,N_4531);
nor UO_720 (O_720,N_4669,N_4683);
nor UO_721 (O_721,N_4621,N_4855);
nand UO_722 (O_722,N_4998,N_4704);
nand UO_723 (O_723,N_4711,N_4729);
or UO_724 (O_724,N_4956,N_4868);
and UO_725 (O_725,N_4728,N_4613);
nand UO_726 (O_726,N_4775,N_4774);
nand UO_727 (O_727,N_4611,N_4688);
xor UO_728 (O_728,N_4836,N_4961);
or UO_729 (O_729,N_4620,N_4576);
xnor UO_730 (O_730,N_4970,N_4875);
nand UO_731 (O_731,N_4682,N_4599);
nand UO_732 (O_732,N_4676,N_4746);
or UO_733 (O_733,N_4635,N_4564);
nor UO_734 (O_734,N_4704,N_4764);
nor UO_735 (O_735,N_4923,N_4772);
nand UO_736 (O_736,N_4936,N_4523);
nor UO_737 (O_737,N_4805,N_4803);
and UO_738 (O_738,N_4808,N_4816);
and UO_739 (O_739,N_4899,N_4750);
or UO_740 (O_740,N_4866,N_4688);
nor UO_741 (O_741,N_4788,N_4854);
or UO_742 (O_742,N_4610,N_4666);
and UO_743 (O_743,N_4797,N_4630);
and UO_744 (O_744,N_4856,N_4617);
or UO_745 (O_745,N_4568,N_4724);
nand UO_746 (O_746,N_4841,N_4735);
or UO_747 (O_747,N_4586,N_4762);
nor UO_748 (O_748,N_4577,N_4885);
nor UO_749 (O_749,N_4735,N_4979);
and UO_750 (O_750,N_4975,N_4546);
nor UO_751 (O_751,N_4785,N_4810);
or UO_752 (O_752,N_4913,N_4708);
or UO_753 (O_753,N_4721,N_4768);
or UO_754 (O_754,N_4883,N_4674);
or UO_755 (O_755,N_4827,N_4575);
or UO_756 (O_756,N_4509,N_4910);
nor UO_757 (O_757,N_4777,N_4959);
or UO_758 (O_758,N_4956,N_4653);
or UO_759 (O_759,N_4560,N_4981);
and UO_760 (O_760,N_4997,N_4878);
nand UO_761 (O_761,N_4926,N_4560);
xnor UO_762 (O_762,N_4523,N_4869);
nand UO_763 (O_763,N_4726,N_4650);
and UO_764 (O_764,N_4645,N_4813);
and UO_765 (O_765,N_4890,N_4841);
nand UO_766 (O_766,N_4584,N_4605);
nor UO_767 (O_767,N_4584,N_4920);
or UO_768 (O_768,N_4904,N_4507);
or UO_769 (O_769,N_4690,N_4582);
or UO_770 (O_770,N_4774,N_4759);
nor UO_771 (O_771,N_4584,N_4870);
nand UO_772 (O_772,N_4878,N_4628);
and UO_773 (O_773,N_4669,N_4723);
nand UO_774 (O_774,N_4619,N_4681);
xor UO_775 (O_775,N_4935,N_4843);
or UO_776 (O_776,N_4697,N_4810);
nor UO_777 (O_777,N_4987,N_4899);
nor UO_778 (O_778,N_4682,N_4704);
nor UO_779 (O_779,N_4837,N_4764);
and UO_780 (O_780,N_4863,N_4737);
or UO_781 (O_781,N_4552,N_4786);
and UO_782 (O_782,N_4850,N_4511);
nor UO_783 (O_783,N_4642,N_4513);
nand UO_784 (O_784,N_4795,N_4577);
nor UO_785 (O_785,N_4788,N_4824);
nor UO_786 (O_786,N_4591,N_4640);
nand UO_787 (O_787,N_4797,N_4775);
nand UO_788 (O_788,N_4600,N_4878);
or UO_789 (O_789,N_4856,N_4880);
nand UO_790 (O_790,N_4552,N_4811);
nor UO_791 (O_791,N_4694,N_4803);
or UO_792 (O_792,N_4778,N_4536);
and UO_793 (O_793,N_4898,N_4949);
nor UO_794 (O_794,N_4675,N_4714);
nor UO_795 (O_795,N_4705,N_4656);
or UO_796 (O_796,N_4694,N_4755);
nand UO_797 (O_797,N_4733,N_4627);
nor UO_798 (O_798,N_4765,N_4883);
nor UO_799 (O_799,N_4661,N_4745);
nor UO_800 (O_800,N_4585,N_4975);
nor UO_801 (O_801,N_4904,N_4618);
nor UO_802 (O_802,N_4885,N_4788);
nand UO_803 (O_803,N_4603,N_4608);
xor UO_804 (O_804,N_4926,N_4806);
and UO_805 (O_805,N_4502,N_4567);
nor UO_806 (O_806,N_4885,N_4740);
nor UO_807 (O_807,N_4562,N_4533);
and UO_808 (O_808,N_4785,N_4959);
or UO_809 (O_809,N_4903,N_4825);
and UO_810 (O_810,N_4594,N_4560);
nor UO_811 (O_811,N_4777,N_4565);
nand UO_812 (O_812,N_4584,N_4857);
nor UO_813 (O_813,N_4817,N_4718);
or UO_814 (O_814,N_4721,N_4775);
nor UO_815 (O_815,N_4605,N_4507);
and UO_816 (O_816,N_4942,N_4627);
or UO_817 (O_817,N_4955,N_4899);
nand UO_818 (O_818,N_4711,N_4640);
and UO_819 (O_819,N_4626,N_4592);
and UO_820 (O_820,N_4762,N_4610);
or UO_821 (O_821,N_4906,N_4764);
and UO_822 (O_822,N_4940,N_4830);
nand UO_823 (O_823,N_4694,N_4669);
or UO_824 (O_824,N_4681,N_4912);
nor UO_825 (O_825,N_4846,N_4829);
and UO_826 (O_826,N_4669,N_4554);
and UO_827 (O_827,N_4893,N_4703);
nor UO_828 (O_828,N_4634,N_4932);
nand UO_829 (O_829,N_4781,N_4720);
nand UO_830 (O_830,N_4528,N_4866);
or UO_831 (O_831,N_4542,N_4976);
nand UO_832 (O_832,N_4954,N_4529);
and UO_833 (O_833,N_4776,N_4511);
and UO_834 (O_834,N_4779,N_4784);
and UO_835 (O_835,N_4900,N_4579);
nor UO_836 (O_836,N_4867,N_4937);
or UO_837 (O_837,N_4525,N_4711);
and UO_838 (O_838,N_4541,N_4978);
or UO_839 (O_839,N_4872,N_4571);
nor UO_840 (O_840,N_4583,N_4750);
and UO_841 (O_841,N_4783,N_4992);
nand UO_842 (O_842,N_4708,N_4590);
nor UO_843 (O_843,N_4820,N_4797);
nor UO_844 (O_844,N_4918,N_4566);
and UO_845 (O_845,N_4578,N_4683);
nor UO_846 (O_846,N_4882,N_4994);
and UO_847 (O_847,N_4918,N_4754);
and UO_848 (O_848,N_4632,N_4672);
nor UO_849 (O_849,N_4954,N_4788);
and UO_850 (O_850,N_4581,N_4808);
or UO_851 (O_851,N_4857,N_4677);
and UO_852 (O_852,N_4566,N_4592);
nor UO_853 (O_853,N_4828,N_4913);
nor UO_854 (O_854,N_4960,N_4760);
or UO_855 (O_855,N_4808,N_4725);
or UO_856 (O_856,N_4844,N_4998);
or UO_857 (O_857,N_4738,N_4993);
nand UO_858 (O_858,N_4817,N_4654);
nor UO_859 (O_859,N_4992,N_4972);
nor UO_860 (O_860,N_4887,N_4697);
and UO_861 (O_861,N_4554,N_4802);
nor UO_862 (O_862,N_4551,N_4957);
or UO_863 (O_863,N_4763,N_4926);
and UO_864 (O_864,N_4951,N_4755);
nor UO_865 (O_865,N_4901,N_4894);
nand UO_866 (O_866,N_4883,N_4994);
and UO_867 (O_867,N_4907,N_4563);
and UO_868 (O_868,N_4903,N_4654);
and UO_869 (O_869,N_4561,N_4546);
and UO_870 (O_870,N_4990,N_4550);
or UO_871 (O_871,N_4706,N_4655);
or UO_872 (O_872,N_4536,N_4548);
or UO_873 (O_873,N_4643,N_4878);
and UO_874 (O_874,N_4870,N_4626);
and UO_875 (O_875,N_4940,N_4608);
nand UO_876 (O_876,N_4740,N_4782);
nor UO_877 (O_877,N_4724,N_4669);
nor UO_878 (O_878,N_4666,N_4812);
or UO_879 (O_879,N_4582,N_4854);
nand UO_880 (O_880,N_4954,N_4972);
and UO_881 (O_881,N_4529,N_4537);
or UO_882 (O_882,N_4688,N_4800);
nand UO_883 (O_883,N_4523,N_4568);
nand UO_884 (O_884,N_4739,N_4885);
and UO_885 (O_885,N_4649,N_4932);
and UO_886 (O_886,N_4914,N_4745);
or UO_887 (O_887,N_4682,N_4917);
nor UO_888 (O_888,N_4937,N_4707);
nand UO_889 (O_889,N_4749,N_4894);
and UO_890 (O_890,N_4706,N_4804);
and UO_891 (O_891,N_4769,N_4654);
or UO_892 (O_892,N_4738,N_4908);
nand UO_893 (O_893,N_4774,N_4922);
or UO_894 (O_894,N_4512,N_4994);
and UO_895 (O_895,N_4604,N_4803);
nor UO_896 (O_896,N_4751,N_4706);
and UO_897 (O_897,N_4997,N_4546);
nor UO_898 (O_898,N_4881,N_4518);
nor UO_899 (O_899,N_4877,N_4512);
and UO_900 (O_900,N_4821,N_4923);
or UO_901 (O_901,N_4582,N_4569);
or UO_902 (O_902,N_4730,N_4785);
and UO_903 (O_903,N_4532,N_4702);
nand UO_904 (O_904,N_4527,N_4875);
nand UO_905 (O_905,N_4796,N_4767);
and UO_906 (O_906,N_4546,N_4628);
and UO_907 (O_907,N_4880,N_4504);
nor UO_908 (O_908,N_4522,N_4948);
or UO_909 (O_909,N_4577,N_4956);
or UO_910 (O_910,N_4683,N_4672);
nand UO_911 (O_911,N_4740,N_4874);
nand UO_912 (O_912,N_4598,N_4773);
or UO_913 (O_913,N_4564,N_4925);
nor UO_914 (O_914,N_4729,N_4641);
xor UO_915 (O_915,N_4521,N_4999);
and UO_916 (O_916,N_4537,N_4695);
xor UO_917 (O_917,N_4752,N_4645);
nand UO_918 (O_918,N_4707,N_4756);
or UO_919 (O_919,N_4819,N_4509);
and UO_920 (O_920,N_4825,N_4682);
nor UO_921 (O_921,N_4517,N_4919);
or UO_922 (O_922,N_4909,N_4948);
nand UO_923 (O_923,N_4820,N_4835);
and UO_924 (O_924,N_4611,N_4982);
nor UO_925 (O_925,N_4573,N_4924);
nor UO_926 (O_926,N_4903,N_4902);
or UO_927 (O_927,N_4553,N_4821);
or UO_928 (O_928,N_4511,N_4845);
or UO_929 (O_929,N_4732,N_4743);
and UO_930 (O_930,N_4738,N_4592);
or UO_931 (O_931,N_4853,N_4582);
or UO_932 (O_932,N_4620,N_4862);
nand UO_933 (O_933,N_4906,N_4962);
and UO_934 (O_934,N_4666,N_4576);
nor UO_935 (O_935,N_4652,N_4894);
nor UO_936 (O_936,N_4932,N_4848);
nand UO_937 (O_937,N_4864,N_4742);
or UO_938 (O_938,N_4549,N_4965);
or UO_939 (O_939,N_4519,N_4612);
nor UO_940 (O_940,N_4934,N_4617);
nand UO_941 (O_941,N_4661,N_4501);
nand UO_942 (O_942,N_4776,N_4637);
or UO_943 (O_943,N_4921,N_4955);
nor UO_944 (O_944,N_4610,N_4620);
or UO_945 (O_945,N_4893,N_4995);
nand UO_946 (O_946,N_4690,N_4535);
nand UO_947 (O_947,N_4779,N_4974);
xnor UO_948 (O_948,N_4732,N_4712);
or UO_949 (O_949,N_4897,N_4609);
and UO_950 (O_950,N_4629,N_4588);
or UO_951 (O_951,N_4909,N_4601);
and UO_952 (O_952,N_4954,N_4810);
and UO_953 (O_953,N_4625,N_4939);
nor UO_954 (O_954,N_4934,N_4833);
nand UO_955 (O_955,N_4867,N_4782);
and UO_956 (O_956,N_4643,N_4857);
or UO_957 (O_957,N_4715,N_4691);
or UO_958 (O_958,N_4706,N_4941);
nor UO_959 (O_959,N_4999,N_4670);
nor UO_960 (O_960,N_4587,N_4892);
nand UO_961 (O_961,N_4929,N_4662);
nor UO_962 (O_962,N_4912,N_4943);
or UO_963 (O_963,N_4831,N_4571);
or UO_964 (O_964,N_4522,N_4847);
or UO_965 (O_965,N_4791,N_4682);
or UO_966 (O_966,N_4892,N_4651);
or UO_967 (O_967,N_4609,N_4822);
nand UO_968 (O_968,N_4587,N_4662);
nor UO_969 (O_969,N_4802,N_4843);
nor UO_970 (O_970,N_4927,N_4732);
and UO_971 (O_971,N_4648,N_4767);
nor UO_972 (O_972,N_4664,N_4726);
and UO_973 (O_973,N_4905,N_4585);
nand UO_974 (O_974,N_4687,N_4736);
or UO_975 (O_975,N_4958,N_4976);
and UO_976 (O_976,N_4893,N_4500);
nand UO_977 (O_977,N_4888,N_4636);
nor UO_978 (O_978,N_4896,N_4734);
xor UO_979 (O_979,N_4610,N_4586);
or UO_980 (O_980,N_4580,N_4517);
and UO_981 (O_981,N_4856,N_4536);
xor UO_982 (O_982,N_4648,N_4918);
xnor UO_983 (O_983,N_4992,N_4669);
and UO_984 (O_984,N_4938,N_4925);
and UO_985 (O_985,N_4897,N_4852);
and UO_986 (O_986,N_4830,N_4559);
or UO_987 (O_987,N_4617,N_4590);
xnor UO_988 (O_988,N_4882,N_4782);
and UO_989 (O_989,N_4521,N_4519);
or UO_990 (O_990,N_4717,N_4909);
or UO_991 (O_991,N_4902,N_4504);
and UO_992 (O_992,N_4930,N_4523);
nand UO_993 (O_993,N_4873,N_4892);
nor UO_994 (O_994,N_4555,N_4532);
nand UO_995 (O_995,N_4630,N_4629);
or UO_996 (O_996,N_4591,N_4585);
nor UO_997 (O_997,N_4926,N_4620);
and UO_998 (O_998,N_4966,N_4709);
and UO_999 (O_999,N_4564,N_4812);
endmodule