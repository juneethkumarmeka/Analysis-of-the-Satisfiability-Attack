module basic_500_3000_500_15_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_438,In_278);
and U1 (N_1,In_200,In_364);
or U2 (N_2,In_426,In_37);
and U3 (N_3,In_7,In_411);
nand U4 (N_4,In_400,In_223);
or U5 (N_5,In_1,In_15);
nor U6 (N_6,In_422,In_106);
nor U7 (N_7,In_417,In_67);
nand U8 (N_8,In_43,In_347);
nand U9 (N_9,In_160,In_336);
and U10 (N_10,In_194,In_314);
nor U11 (N_11,In_195,In_392);
xnor U12 (N_12,In_159,In_430);
nor U13 (N_13,In_482,In_253);
nor U14 (N_14,In_76,In_330);
xor U15 (N_15,In_36,In_313);
nor U16 (N_16,In_45,In_345);
nor U17 (N_17,In_465,In_468);
and U18 (N_18,In_369,In_265);
and U19 (N_19,In_326,In_229);
nor U20 (N_20,In_157,In_351);
nor U21 (N_21,In_379,In_332);
nor U22 (N_22,In_376,In_499);
or U23 (N_23,In_286,In_473);
and U24 (N_24,In_252,In_335);
or U25 (N_25,In_377,In_448);
and U26 (N_26,In_375,In_139);
or U27 (N_27,In_466,In_264);
nor U28 (N_28,In_105,In_18);
nor U29 (N_29,In_40,In_96);
nand U30 (N_30,In_236,In_151);
and U31 (N_31,In_249,In_290);
and U32 (N_32,In_387,In_74);
nand U33 (N_33,In_109,In_235);
nand U34 (N_34,In_220,In_32);
nor U35 (N_35,In_414,In_359);
nor U36 (N_36,In_239,In_172);
and U37 (N_37,In_383,In_108);
nand U38 (N_38,In_193,In_85);
nand U39 (N_39,In_184,In_386);
or U40 (N_40,In_101,In_120);
nand U41 (N_41,In_207,In_24);
nand U42 (N_42,In_479,In_55);
and U43 (N_43,In_111,In_115);
and U44 (N_44,In_363,In_140);
nand U45 (N_45,In_215,In_384);
or U46 (N_46,In_51,In_256);
or U47 (N_47,In_353,In_149);
or U48 (N_48,In_315,In_135);
nor U49 (N_49,In_487,In_268);
nor U50 (N_50,In_457,In_308);
or U51 (N_51,In_324,In_127);
nor U52 (N_52,In_154,In_14);
nand U53 (N_53,In_8,In_441);
nor U54 (N_54,In_431,In_209);
or U55 (N_55,In_196,In_243);
xor U56 (N_56,In_344,In_167);
nor U57 (N_57,In_453,In_77);
or U58 (N_58,In_83,In_445);
nor U59 (N_59,In_251,In_285);
and U60 (N_60,In_263,In_131);
nand U61 (N_61,In_19,In_233);
nand U62 (N_62,In_30,In_355);
nand U63 (N_63,In_170,In_2);
nand U64 (N_64,In_318,In_93);
and U65 (N_65,In_44,In_132);
nand U66 (N_66,In_173,In_10);
nor U67 (N_67,In_238,In_272);
or U68 (N_68,In_449,In_283);
or U69 (N_69,In_291,In_87);
and U70 (N_70,In_31,In_186);
and U71 (N_71,In_33,In_153);
and U72 (N_72,In_124,In_425);
xor U73 (N_73,In_381,In_248);
nor U74 (N_74,In_306,In_419);
or U75 (N_75,In_46,In_57);
and U76 (N_76,In_434,In_491);
nor U77 (N_77,In_295,In_292);
nand U78 (N_78,In_446,In_79);
nand U79 (N_79,In_126,In_257);
nand U80 (N_80,In_394,In_179);
or U81 (N_81,In_224,In_316);
nand U82 (N_82,In_452,In_174);
nor U83 (N_83,In_432,In_294);
nand U84 (N_84,In_475,In_152);
and U85 (N_85,In_439,In_338);
nor U86 (N_86,In_389,In_218);
or U87 (N_87,In_423,In_302);
nand U88 (N_88,In_322,In_150);
or U89 (N_89,In_429,In_420);
or U90 (N_90,In_192,In_496);
and U91 (N_91,In_6,In_370);
nor U92 (N_92,In_399,In_407);
and U93 (N_93,In_130,In_143);
nand U94 (N_94,In_16,In_25);
xor U95 (N_95,In_462,In_89);
or U96 (N_96,In_365,In_418);
or U97 (N_97,In_175,In_99);
nand U98 (N_98,In_279,In_360);
nor U99 (N_99,In_169,In_176);
nand U100 (N_100,In_357,In_110);
nand U101 (N_101,In_262,In_97);
nor U102 (N_102,In_346,In_191);
nand U103 (N_103,In_447,In_444);
and U104 (N_104,In_199,In_297);
nand U105 (N_105,In_421,In_82);
nand U106 (N_106,In_497,In_320);
and U107 (N_107,In_492,In_61);
nor U108 (N_108,In_408,In_480);
nand U109 (N_109,In_107,In_323);
nor U110 (N_110,In_352,In_488);
nor U111 (N_111,In_467,In_266);
nand U112 (N_112,In_12,In_78);
and U113 (N_113,In_328,In_133);
nor U114 (N_114,In_197,In_329);
nor U115 (N_115,In_495,In_189);
nor U116 (N_116,In_354,In_39);
or U117 (N_117,In_455,In_208);
nand U118 (N_118,In_41,In_202);
and U119 (N_119,In_185,In_433);
nand U120 (N_120,In_403,In_361);
or U121 (N_121,In_141,In_288);
nor U122 (N_122,In_312,In_289);
nand U123 (N_123,In_62,In_410);
nor U124 (N_124,In_60,In_216);
nand U125 (N_125,In_22,In_222);
nand U126 (N_126,In_374,In_21);
or U127 (N_127,In_86,In_398);
and U128 (N_128,In_118,In_246);
nor U129 (N_129,In_481,In_284);
or U130 (N_130,In_68,In_64);
and U131 (N_131,In_260,In_282);
and U132 (N_132,In_443,In_413);
nor U133 (N_133,In_119,In_472);
or U134 (N_134,In_300,In_80);
or U135 (N_135,In_305,In_307);
nand U136 (N_136,In_158,In_134);
nor U137 (N_137,In_146,In_56);
nor U138 (N_138,In_415,In_340);
nor U139 (N_139,In_214,In_227);
nor U140 (N_140,In_450,In_47);
or U141 (N_141,In_245,In_95);
nand U142 (N_142,In_104,In_221);
xnor U143 (N_143,In_485,In_319);
nand U144 (N_144,In_123,In_180);
nor U145 (N_145,In_397,In_366);
and U146 (N_146,In_116,In_117);
and U147 (N_147,In_5,In_406);
or U148 (N_148,In_136,In_50);
nor U149 (N_149,In_404,In_163);
nor U150 (N_150,In_331,In_91);
and U151 (N_151,In_287,In_201);
or U152 (N_152,In_372,In_81);
nand U153 (N_153,In_38,In_402);
nand U154 (N_154,In_145,In_327);
nor U155 (N_155,In_90,In_490);
nand U156 (N_156,In_231,In_293);
nand U157 (N_157,In_210,In_321);
nor U158 (N_158,In_20,In_471);
nand U159 (N_159,In_65,In_476);
or U160 (N_160,In_17,In_122);
or U161 (N_161,In_9,In_275);
and U162 (N_162,In_416,In_52);
nor U163 (N_163,In_382,In_232);
or U164 (N_164,In_54,In_178);
and U165 (N_165,In_226,In_137);
nor U166 (N_166,In_470,In_486);
nand U167 (N_167,In_269,In_325);
or U168 (N_168,In_212,In_343);
or U169 (N_169,In_211,In_190);
or U170 (N_170,In_464,In_396);
nor U171 (N_171,In_92,In_254);
nor U172 (N_172,In_166,In_401);
and U173 (N_173,In_277,In_128);
nand U174 (N_174,In_59,In_53);
and U175 (N_175,In_26,In_469);
and U176 (N_176,In_230,In_459);
and U177 (N_177,In_0,In_270);
and U178 (N_178,In_255,In_484);
nand U179 (N_179,In_409,In_342);
and U180 (N_180,In_390,In_155);
or U181 (N_181,In_349,In_205);
nor U182 (N_182,In_388,In_165);
and U183 (N_183,In_156,In_427);
or U184 (N_184,In_113,In_296);
or U185 (N_185,In_225,In_273);
xnor U186 (N_186,In_267,In_436);
nor U187 (N_187,In_378,In_494);
or U188 (N_188,In_49,In_168);
nand U189 (N_189,In_34,In_247);
nor U190 (N_190,In_242,In_63);
nor U191 (N_191,In_188,In_4);
nor U192 (N_192,In_395,In_13);
nand U193 (N_193,In_348,In_42);
and U194 (N_194,In_187,In_271);
nor U195 (N_195,In_385,In_456);
nor U196 (N_196,In_73,In_27);
and U197 (N_197,In_198,In_206);
and U198 (N_198,In_98,In_380);
nand U199 (N_199,In_48,In_303);
and U200 (N_200,N_185,In_234);
nand U201 (N_201,N_197,N_71);
or U202 (N_202,N_146,N_129);
nand U203 (N_203,In_317,N_128);
nand U204 (N_204,In_237,N_103);
or U205 (N_205,N_144,N_79);
nor U206 (N_206,N_32,In_281);
nor U207 (N_207,N_198,N_11);
nor U208 (N_208,In_451,N_125);
nor U209 (N_209,N_59,In_483);
nand U210 (N_210,N_21,N_132);
nor U211 (N_211,N_161,In_35);
or U212 (N_212,N_50,In_371);
or U213 (N_213,N_72,In_181);
and U214 (N_214,N_199,N_26);
and U215 (N_215,In_478,In_489);
or U216 (N_216,In_28,N_149);
or U217 (N_217,In_121,In_298);
nand U218 (N_218,In_177,In_463);
or U219 (N_219,N_151,N_81);
nand U220 (N_220,N_135,N_189);
nand U221 (N_221,In_240,N_173);
nand U222 (N_222,N_51,N_119);
nand U223 (N_223,N_184,In_3);
and U224 (N_224,N_3,N_101);
nor U225 (N_225,N_140,N_171);
or U226 (N_226,In_213,In_337);
or U227 (N_227,N_16,In_183);
or U228 (N_228,In_368,In_498);
nand U229 (N_229,N_166,In_162);
nand U230 (N_230,In_280,N_22);
nand U231 (N_231,N_83,In_142);
or U232 (N_232,N_45,N_66);
and U233 (N_233,In_428,N_40);
nand U234 (N_234,N_5,In_276);
nand U235 (N_235,N_195,N_82);
or U236 (N_236,N_186,N_70);
or U237 (N_237,N_164,N_158);
and U238 (N_238,N_13,In_258);
nand U239 (N_239,In_309,N_124);
and U240 (N_240,N_87,N_8);
nand U241 (N_241,N_46,N_133);
and U242 (N_242,N_93,N_56);
or U243 (N_243,N_139,N_183);
or U244 (N_244,N_172,N_115);
and U245 (N_245,N_194,N_112);
or U246 (N_246,In_440,In_412);
and U247 (N_247,N_169,In_144);
nor U248 (N_248,In_102,In_474);
or U249 (N_249,N_36,N_58);
nor U250 (N_250,N_117,In_460);
and U251 (N_251,N_9,N_145);
xor U252 (N_252,N_108,N_134);
and U253 (N_253,In_333,N_123);
xnor U254 (N_254,In_261,N_35);
and U255 (N_255,N_90,N_6);
nor U256 (N_256,N_19,N_181);
xor U257 (N_257,In_58,N_76);
nand U258 (N_258,In_148,In_138);
xnor U259 (N_259,N_127,In_66);
nor U260 (N_260,N_29,In_391);
or U261 (N_261,N_191,N_153);
nand U262 (N_262,N_23,N_49);
nand U263 (N_263,N_96,N_24);
nand U264 (N_264,N_157,N_20);
nor U265 (N_265,In_29,N_187);
and U266 (N_266,N_34,N_10);
and U267 (N_267,N_137,N_105);
nor U268 (N_268,In_164,In_112);
nor U269 (N_269,N_28,N_114);
and U270 (N_270,In_219,N_156);
nand U271 (N_271,In_103,In_350);
and U272 (N_272,N_111,In_69);
xnor U273 (N_273,N_27,N_95);
xnor U274 (N_274,In_23,N_12);
and U275 (N_275,N_179,N_41);
xor U276 (N_276,In_393,N_38);
nor U277 (N_277,In_250,N_106);
xnor U278 (N_278,In_100,In_125);
and U279 (N_279,N_86,N_92);
or U280 (N_280,In_454,N_69);
xnor U281 (N_281,N_188,N_73);
nand U282 (N_282,N_162,N_2);
or U283 (N_283,In_129,In_334);
nand U284 (N_284,N_136,In_217);
nor U285 (N_285,N_53,N_64);
and U286 (N_286,N_170,N_65);
and U287 (N_287,N_174,N_61);
nand U288 (N_288,In_367,N_68);
and U289 (N_289,In_311,N_1);
nor U290 (N_290,N_44,N_54);
xor U291 (N_291,In_299,N_178);
and U292 (N_292,N_177,In_339);
nand U293 (N_293,N_42,In_274);
or U294 (N_294,In_114,N_180);
xor U295 (N_295,N_160,In_88);
xnor U296 (N_296,N_60,N_154);
or U297 (N_297,In_461,N_107);
or U298 (N_298,N_110,N_182);
or U299 (N_299,N_47,In_84);
nor U300 (N_300,In_458,N_91);
nand U301 (N_301,In_11,N_39);
nor U302 (N_302,N_15,N_80);
nor U303 (N_303,N_138,In_147);
nand U304 (N_304,In_70,N_147);
nand U305 (N_305,N_7,N_100);
nor U306 (N_306,In_424,N_165);
and U307 (N_307,N_104,In_405);
nand U308 (N_308,N_4,N_102);
and U309 (N_309,In_442,In_171);
nor U310 (N_310,N_196,In_182);
nand U311 (N_311,N_152,N_159);
and U312 (N_312,N_57,N_131);
or U313 (N_313,N_176,In_71);
nor U314 (N_314,N_175,N_30);
nor U315 (N_315,In_310,N_67);
xnor U316 (N_316,N_190,In_244);
nor U317 (N_317,N_109,In_477);
nand U318 (N_318,N_98,In_362);
nand U319 (N_319,In_358,N_97);
nor U320 (N_320,In_435,In_204);
nor U321 (N_321,N_167,N_118);
nand U322 (N_322,N_121,N_78);
or U323 (N_323,N_163,N_113);
or U324 (N_324,N_17,N_74);
nand U325 (N_325,In_94,N_75);
nor U326 (N_326,In_72,N_48);
and U327 (N_327,In_304,In_341);
nand U328 (N_328,In_75,N_148);
nor U329 (N_329,N_168,In_259);
xor U330 (N_330,N_142,N_88);
nor U331 (N_331,N_62,N_77);
nand U332 (N_332,N_99,N_143);
nor U333 (N_333,N_37,N_85);
or U334 (N_334,In_437,N_25);
or U335 (N_335,In_228,N_130);
and U336 (N_336,N_43,N_116);
nand U337 (N_337,N_18,N_126);
or U338 (N_338,N_14,N_52);
and U339 (N_339,N_0,N_193);
nor U340 (N_340,In_301,N_55);
and U341 (N_341,In_203,N_89);
or U342 (N_342,N_94,N_122);
and U343 (N_343,N_150,N_120);
and U344 (N_344,In_241,In_356);
and U345 (N_345,N_141,N_33);
and U346 (N_346,In_493,N_192);
nor U347 (N_347,N_84,In_373);
and U348 (N_348,N_31,N_63);
or U349 (N_349,N_155,In_161);
nand U350 (N_350,N_152,N_108);
nor U351 (N_351,In_393,N_56);
nor U352 (N_352,In_463,N_199);
or U353 (N_353,N_149,In_358);
and U354 (N_354,N_56,N_191);
or U355 (N_355,N_194,In_11);
nor U356 (N_356,N_181,N_6);
nand U357 (N_357,In_171,N_167);
nand U358 (N_358,In_144,N_93);
nand U359 (N_359,N_47,N_88);
nor U360 (N_360,In_88,N_149);
xor U361 (N_361,In_442,N_11);
and U362 (N_362,N_83,In_311);
nor U363 (N_363,N_64,In_310);
nand U364 (N_364,In_219,N_171);
nor U365 (N_365,In_204,N_195);
and U366 (N_366,N_99,In_451);
and U367 (N_367,N_37,N_34);
and U368 (N_368,N_168,In_261);
nand U369 (N_369,N_181,In_442);
nor U370 (N_370,N_20,N_71);
and U371 (N_371,In_161,N_60);
nor U372 (N_372,In_112,N_134);
nand U373 (N_373,In_478,N_129);
and U374 (N_374,In_405,N_114);
or U375 (N_375,In_391,In_280);
nand U376 (N_376,N_157,N_60);
nand U377 (N_377,N_60,In_164);
nand U378 (N_378,N_92,N_171);
nand U379 (N_379,N_138,N_123);
nor U380 (N_380,N_183,N_102);
nand U381 (N_381,In_317,N_173);
nand U382 (N_382,N_143,N_189);
and U383 (N_383,N_114,N_38);
and U384 (N_384,In_228,N_181);
and U385 (N_385,In_28,N_72);
and U386 (N_386,N_130,In_244);
or U387 (N_387,In_362,In_259);
nand U388 (N_388,N_194,N_7);
nor U389 (N_389,In_483,In_204);
and U390 (N_390,N_73,N_32);
or U391 (N_391,In_58,N_110);
and U392 (N_392,N_72,N_95);
or U393 (N_393,In_144,N_36);
nor U394 (N_394,N_181,N_197);
or U395 (N_395,N_125,N_132);
or U396 (N_396,N_13,N_159);
nor U397 (N_397,N_105,N_109);
and U398 (N_398,In_317,N_99);
xor U399 (N_399,In_103,In_435);
or U400 (N_400,N_364,N_218);
nor U401 (N_401,N_349,N_363);
or U402 (N_402,N_241,N_390);
nand U403 (N_403,N_226,N_329);
or U404 (N_404,N_348,N_286);
and U405 (N_405,N_288,N_382);
nand U406 (N_406,N_359,N_303);
nor U407 (N_407,N_287,N_207);
nor U408 (N_408,N_362,N_396);
or U409 (N_409,N_267,N_335);
and U410 (N_410,N_262,N_320);
or U411 (N_411,N_245,N_238);
or U412 (N_412,N_330,N_203);
and U413 (N_413,N_264,N_334);
nand U414 (N_414,N_270,N_361);
and U415 (N_415,N_388,N_315);
nor U416 (N_416,N_391,N_277);
nand U417 (N_417,N_380,N_229);
and U418 (N_418,N_208,N_310);
nor U419 (N_419,N_338,N_222);
or U420 (N_420,N_231,N_296);
and U421 (N_421,N_344,N_216);
nand U422 (N_422,N_341,N_283);
nor U423 (N_423,N_394,N_299);
nand U424 (N_424,N_379,N_302);
and U425 (N_425,N_221,N_251);
or U426 (N_426,N_351,N_263);
or U427 (N_427,N_342,N_383);
or U428 (N_428,N_331,N_276);
nor U429 (N_429,N_300,N_274);
nor U430 (N_430,N_386,N_212);
or U431 (N_431,N_244,N_206);
and U432 (N_432,N_255,N_378);
nor U433 (N_433,N_311,N_210);
or U434 (N_434,N_202,N_314);
nand U435 (N_435,N_318,N_399);
and U436 (N_436,N_317,N_301);
nor U437 (N_437,N_393,N_304);
and U438 (N_438,N_224,N_260);
and U439 (N_439,N_230,N_384);
or U440 (N_440,N_392,N_339);
and U441 (N_441,N_326,N_272);
nor U442 (N_442,N_239,N_345);
and U443 (N_443,N_259,N_346);
and U444 (N_444,N_305,N_282);
nor U445 (N_445,N_225,N_316);
and U446 (N_446,N_324,N_281);
and U447 (N_447,N_232,N_217);
and U448 (N_448,N_257,N_371);
nor U449 (N_449,N_297,N_369);
and U450 (N_450,N_271,N_356);
nand U451 (N_451,N_347,N_366);
and U452 (N_452,N_375,N_385);
and U453 (N_453,N_309,N_332);
and U454 (N_454,N_358,N_248);
or U455 (N_455,N_295,N_340);
and U456 (N_456,N_389,N_343);
nor U457 (N_457,N_360,N_327);
or U458 (N_458,N_201,N_292);
xor U459 (N_459,N_254,N_242);
nor U460 (N_460,N_307,N_228);
and U461 (N_461,N_294,N_219);
and U462 (N_462,N_275,N_265);
nand U463 (N_463,N_377,N_354);
or U464 (N_464,N_337,N_372);
nand U465 (N_465,N_289,N_205);
nor U466 (N_466,N_323,N_365);
nand U467 (N_467,N_352,N_290);
nor U468 (N_468,N_235,N_322);
or U469 (N_469,N_278,N_285);
nor U470 (N_470,N_333,N_373);
or U471 (N_471,N_336,N_353);
nand U472 (N_472,N_215,N_227);
nor U473 (N_473,N_236,N_268);
or U474 (N_474,N_398,N_211);
or U475 (N_475,N_233,N_397);
and U476 (N_476,N_204,N_243);
nand U477 (N_477,N_279,N_367);
nor U478 (N_478,N_240,N_298);
nor U479 (N_479,N_284,N_247);
or U480 (N_480,N_223,N_256);
and U481 (N_481,N_328,N_293);
and U482 (N_482,N_266,N_355);
and U483 (N_483,N_200,N_319);
and U484 (N_484,N_246,N_370);
or U485 (N_485,N_252,N_209);
nand U486 (N_486,N_249,N_306);
and U487 (N_487,N_253,N_291);
and U488 (N_488,N_261,N_273);
nand U489 (N_489,N_308,N_220);
and U490 (N_490,N_213,N_234);
or U491 (N_491,N_214,N_269);
and U492 (N_492,N_387,N_258);
nand U493 (N_493,N_374,N_280);
or U494 (N_494,N_325,N_312);
or U495 (N_495,N_350,N_381);
nand U496 (N_496,N_368,N_395);
and U497 (N_497,N_357,N_250);
nor U498 (N_498,N_313,N_237);
nand U499 (N_499,N_321,N_376);
and U500 (N_500,N_324,N_289);
nand U501 (N_501,N_238,N_202);
nor U502 (N_502,N_277,N_290);
and U503 (N_503,N_330,N_318);
nor U504 (N_504,N_329,N_265);
and U505 (N_505,N_315,N_360);
xnor U506 (N_506,N_364,N_201);
nand U507 (N_507,N_216,N_255);
nor U508 (N_508,N_304,N_313);
nor U509 (N_509,N_338,N_220);
or U510 (N_510,N_317,N_335);
nor U511 (N_511,N_278,N_208);
nor U512 (N_512,N_262,N_379);
and U513 (N_513,N_343,N_329);
or U514 (N_514,N_357,N_256);
nand U515 (N_515,N_278,N_273);
or U516 (N_516,N_238,N_206);
nor U517 (N_517,N_351,N_238);
or U518 (N_518,N_359,N_380);
nor U519 (N_519,N_218,N_387);
nand U520 (N_520,N_217,N_398);
nand U521 (N_521,N_222,N_263);
or U522 (N_522,N_364,N_238);
nor U523 (N_523,N_239,N_371);
nor U524 (N_524,N_287,N_338);
or U525 (N_525,N_286,N_218);
and U526 (N_526,N_288,N_268);
or U527 (N_527,N_281,N_222);
and U528 (N_528,N_351,N_214);
or U529 (N_529,N_350,N_210);
and U530 (N_530,N_300,N_361);
nor U531 (N_531,N_272,N_200);
nand U532 (N_532,N_318,N_218);
and U533 (N_533,N_237,N_238);
and U534 (N_534,N_246,N_228);
xor U535 (N_535,N_207,N_367);
nor U536 (N_536,N_292,N_272);
or U537 (N_537,N_238,N_273);
nand U538 (N_538,N_207,N_380);
nor U539 (N_539,N_283,N_301);
nor U540 (N_540,N_389,N_234);
or U541 (N_541,N_364,N_284);
nor U542 (N_542,N_341,N_251);
and U543 (N_543,N_278,N_396);
nand U544 (N_544,N_288,N_337);
or U545 (N_545,N_200,N_353);
and U546 (N_546,N_304,N_255);
and U547 (N_547,N_313,N_383);
nand U548 (N_548,N_388,N_242);
nand U549 (N_549,N_398,N_359);
or U550 (N_550,N_331,N_375);
nand U551 (N_551,N_327,N_303);
and U552 (N_552,N_377,N_262);
and U553 (N_553,N_268,N_377);
nor U554 (N_554,N_340,N_200);
and U555 (N_555,N_374,N_376);
nor U556 (N_556,N_320,N_347);
or U557 (N_557,N_346,N_251);
and U558 (N_558,N_374,N_270);
nor U559 (N_559,N_236,N_271);
nand U560 (N_560,N_269,N_346);
nor U561 (N_561,N_328,N_332);
nor U562 (N_562,N_266,N_299);
and U563 (N_563,N_211,N_345);
or U564 (N_564,N_387,N_244);
and U565 (N_565,N_374,N_253);
nor U566 (N_566,N_320,N_230);
nor U567 (N_567,N_214,N_381);
nor U568 (N_568,N_334,N_203);
and U569 (N_569,N_245,N_394);
nand U570 (N_570,N_275,N_389);
nor U571 (N_571,N_229,N_253);
or U572 (N_572,N_318,N_275);
nor U573 (N_573,N_305,N_236);
or U574 (N_574,N_227,N_301);
or U575 (N_575,N_306,N_304);
or U576 (N_576,N_385,N_365);
or U577 (N_577,N_395,N_201);
nand U578 (N_578,N_315,N_243);
nor U579 (N_579,N_355,N_370);
nor U580 (N_580,N_308,N_299);
and U581 (N_581,N_212,N_333);
and U582 (N_582,N_298,N_279);
or U583 (N_583,N_391,N_238);
nor U584 (N_584,N_251,N_276);
nand U585 (N_585,N_289,N_252);
or U586 (N_586,N_253,N_389);
and U587 (N_587,N_219,N_269);
nor U588 (N_588,N_240,N_247);
nand U589 (N_589,N_351,N_203);
nand U590 (N_590,N_246,N_358);
nand U591 (N_591,N_283,N_381);
or U592 (N_592,N_213,N_201);
nor U593 (N_593,N_218,N_371);
nor U594 (N_594,N_338,N_200);
and U595 (N_595,N_377,N_382);
or U596 (N_596,N_248,N_285);
nand U597 (N_597,N_363,N_274);
and U598 (N_598,N_257,N_367);
nor U599 (N_599,N_397,N_218);
or U600 (N_600,N_533,N_484);
or U601 (N_601,N_436,N_514);
and U602 (N_602,N_580,N_463);
and U603 (N_603,N_487,N_465);
nand U604 (N_604,N_479,N_500);
and U605 (N_605,N_432,N_468);
nor U606 (N_606,N_518,N_460);
nand U607 (N_607,N_483,N_585);
and U608 (N_608,N_488,N_525);
or U609 (N_609,N_534,N_467);
and U610 (N_610,N_446,N_564);
nand U611 (N_611,N_576,N_473);
or U612 (N_612,N_437,N_400);
nor U613 (N_613,N_438,N_428);
or U614 (N_614,N_563,N_586);
nor U615 (N_615,N_521,N_471);
nor U616 (N_616,N_526,N_490);
nand U617 (N_617,N_413,N_548);
nand U618 (N_618,N_502,N_451);
or U619 (N_619,N_540,N_424);
or U620 (N_620,N_419,N_551);
nand U621 (N_621,N_578,N_594);
nor U622 (N_622,N_567,N_477);
nor U623 (N_623,N_452,N_401);
nand U624 (N_624,N_486,N_539);
nand U625 (N_625,N_530,N_415);
or U626 (N_626,N_547,N_542);
nand U627 (N_627,N_423,N_513);
or U628 (N_628,N_412,N_427);
nand U629 (N_629,N_455,N_565);
and U630 (N_630,N_442,N_449);
nand U631 (N_631,N_430,N_404);
and U632 (N_632,N_566,N_497);
and U633 (N_633,N_596,N_407);
or U634 (N_634,N_470,N_405);
or U635 (N_635,N_402,N_506);
and U636 (N_636,N_549,N_543);
nor U637 (N_637,N_433,N_426);
and U638 (N_638,N_571,N_541);
and U639 (N_639,N_410,N_509);
nand U640 (N_640,N_453,N_511);
and U641 (N_641,N_589,N_418);
or U642 (N_642,N_577,N_527);
or U643 (N_643,N_510,N_579);
nor U644 (N_644,N_573,N_590);
nand U645 (N_645,N_560,N_458);
nand U646 (N_646,N_457,N_441);
nand U647 (N_647,N_522,N_422);
xor U648 (N_648,N_599,N_425);
nand U649 (N_649,N_538,N_535);
nand U650 (N_650,N_469,N_492);
and U651 (N_651,N_501,N_411);
nand U652 (N_652,N_443,N_498);
nor U653 (N_653,N_505,N_550);
or U654 (N_654,N_508,N_447);
or U655 (N_655,N_588,N_545);
nor U656 (N_656,N_557,N_528);
nand U657 (N_657,N_466,N_481);
nor U658 (N_658,N_429,N_461);
nand U659 (N_659,N_558,N_403);
nand U660 (N_660,N_524,N_459);
or U661 (N_661,N_570,N_523);
and U662 (N_662,N_507,N_478);
nor U663 (N_663,N_552,N_431);
nor U664 (N_664,N_475,N_489);
nor U665 (N_665,N_417,N_499);
nand U666 (N_666,N_450,N_517);
and U667 (N_667,N_435,N_476);
nand U668 (N_668,N_598,N_536);
or U669 (N_669,N_503,N_519);
and U670 (N_670,N_406,N_515);
nor U671 (N_671,N_480,N_587);
nor U672 (N_672,N_472,N_583);
and U673 (N_673,N_554,N_474);
xor U674 (N_674,N_531,N_584);
nand U675 (N_675,N_482,N_553);
or U676 (N_676,N_462,N_444);
nor U677 (N_677,N_597,N_555);
xnor U678 (N_678,N_537,N_496);
nor U679 (N_679,N_494,N_409);
nand U680 (N_680,N_414,N_562);
or U681 (N_681,N_581,N_592);
and U682 (N_682,N_493,N_559);
or U683 (N_683,N_591,N_572);
and U684 (N_684,N_456,N_561);
and U685 (N_685,N_464,N_582);
nor U686 (N_686,N_546,N_512);
or U687 (N_687,N_421,N_485);
nand U688 (N_688,N_568,N_556);
or U689 (N_689,N_495,N_593);
nor U690 (N_690,N_575,N_491);
nand U691 (N_691,N_532,N_445);
nor U692 (N_692,N_544,N_440);
or U693 (N_693,N_595,N_504);
nand U694 (N_694,N_516,N_448);
nand U695 (N_695,N_420,N_408);
nor U696 (N_696,N_434,N_416);
nand U697 (N_697,N_454,N_574);
or U698 (N_698,N_529,N_439);
nor U699 (N_699,N_520,N_569);
xnor U700 (N_700,N_406,N_526);
or U701 (N_701,N_430,N_460);
and U702 (N_702,N_518,N_486);
xnor U703 (N_703,N_467,N_577);
nor U704 (N_704,N_464,N_468);
nor U705 (N_705,N_497,N_541);
nand U706 (N_706,N_453,N_593);
nor U707 (N_707,N_459,N_485);
nor U708 (N_708,N_569,N_459);
nand U709 (N_709,N_457,N_546);
nand U710 (N_710,N_550,N_547);
nor U711 (N_711,N_458,N_478);
and U712 (N_712,N_599,N_415);
nor U713 (N_713,N_403,N_438);
or U714 (N_714,N_503,N_445);
nor U715 (N_715,N_450,N_424);
nor U716 (N_716,N_528,N_400);
nor U717 (N_717,N_438,N_599);
nor U718 (N_718,N_403,N_493);
and U719 (N_719,N_548,N_426);
nand U720 (N_720,N_473,N_579);
or U721 (N_721,N_401,N_562);
and U722 (N_722,N_559,N_429);
nand U723 (N_723,N_505,N_588);
nor U724 (N_724,N_441,N_403);
or U725 (N_725,N_508,N_477);
nor U726 (N_726,N_557,N_582);
or U727 (N_727,N_546,N_550);
or U728 (N_728,N_499,N_508);
and U729 (N_729,N_527,N_452);
nor U730 (N_730,N_499,N_415);
nor U731 (N_731,N_500,N_402);
nor U732 (N_732,N_406,N_598);
and U733 (N_733,N_588,N_594);
nor U734 (N_734,N_441,N_524);
nand U735 (N_735,N_440,N_568);
and U736 (N_736,N_415,N_446);
nor U737 (N_737,N_572,N_589);
or U738 (N_738,N_582,N_598);
or U739 (N_739,N_530,N_519);
or U740 (N_740,N_462,N_536);
and U741 (N_741,N_411,N_400);
or U742 (N_742,N_554,N_419);
nand U743 (N_743,N_439,N_588);
and U744 (N_744,N_597,N_593);
or U745 (N_745,N_570,N_482);
and U746 (N_746,N_578,N_412);
or U747 (N_747,N_452,N_559);
nor U748 (N_748,N_559,N_512);
or U749 (N_749,N_453,N_581);
nand U750 (N_750,N_498,N_591);
nand U751 (N_751,N_501,N_479);
and U752 (N_752,N_548,N_404);
nor U753 (N_753,N_470,N_453);
nor U754 (N_754,N_420,N_460);
or U755 (N_755,N_504,N_473);
nand U756 (N_756,N_599,N_463);
nor U757 (N_757,N_461,N_596);
or U758 (N_758,N_425,N_433);
nand U759 (N_759,N_537,N_596);
nand U760 (N_760,N_423,N_494);
or U761 (N_761,N_433,N_578);
nand U762 (N_762,N_417,N_531);
nand U763 (N_763,N_403,N_440);
or U764 (N_764,N_565,N_513);
and U765 (N_765,N_559,N_510);
nor U766 (N_766,N_457,N_440);
nor U767 (N_767,N_445,N_431);
nand U768 (N_768,N_484,N_562);
and U769 (N_769,N_419,N_548);
and U770 (N_770,N_501,N_504);
and U771 (N_771,N_507,N_548);
nand U772 (N_772,N_537,N_563);
nor U773 (N_773,N_491,N_409);
nor U774 (N_774,N_539,N_437);
or U775 (N_775,N_590,N_435);
nand U776 (N_776,N_481,N_485);
and U777 (N_777,N_539,N_585);
and U778 (N_778,N_434,N_575);
or U779 (N_779,N_520,N_415);
and U780 (N_780,N_478,N_455);
nand U781 (N_781,N_550,N_585);
and U782 (N_782,N_595,N_458);
and U783 (N_783,N_436,N_446);
nor U784 (N_784,N_548,N_599);
nand U785 (N_785,N_487,N_483);
nor U786 (N_786,N_461,N_575);
nor U787 (N_787,N_539,N_495);
nand U788 (N_788,N_560,N_436);
or U789 (N_789,N_432,N_530);
or U790 (N_790,N_584,N_493);
nand U791 (N_791,N_432,N_556);
nor U792 (N_792,N_525,N_453);
and U793 (N_793,N_404,N_449);
nor U794 (N_794,N_472,N_577);
nand U795 (N_795,N_491,N_570);
or U796 (N_796,N_465,N_453);
or U797 (N_797,N_461,N_534);
or U798 (N_798,N_516,N_420);
nor U799 (N_799,N_437,N_499);
nor U800 (N_800,N_742,N_785);
nor U801 (N_801,N_701,N_646);
nand U802 (N_802,N_657,N_601);
nor U803 (N_803,N_789,N_730);
nand U804 (N_804,N_723,N_645);
xnor U805 (N_805,N_665,N_712);
or U806 (N_806,N_647,N_672);
nand U807 (N_807,N_690,N_615);
nand U808 (N_808,N_744,N_724);
nor U809 (N_809,N_697,N_791);
nand U810 (N_810,N_614,N_639);
or U811 (N_811,N_671,N_698);
or U812 (N_812,N_654,N_727);
or U813 (N_813,N_661,N_768);
nor U814 (N_814,N_670,N_644);
nor U815 (N_815,N_777,N_632);
or U816 (N_816,N_638,N_634);
and U817 (N_817,N_626,N_737);
or U818 (N_818,N_685,N_678);
nor U819 (N_819,N_694,N_709);
or U820 (N_820,N_771,N_649);
or U821 (N_821,N_676,N_655);
nor U822 (N_822,N_703,N_790);
nor U823 (N_823,N_714,N_659);
and U824 (N_824,N_782,N_793);
nand U825 (N_825,N_754,N_682);
and U826 (N_826,N_795,N_721);
and U827 (N_827,N_758,N_648);
nor U828 (N_828,N_766,N_767);
or U829 (N_829,N_708,N_731);
xnor U830 (N_830,N_786,N_713);
and U831 (N_831,N_666,N_692);
nand U832 (N_832,N_700,N_711);
nand U833 (N_833,N_618,N_761);
and U834 (N_834,N_728,N_624);
nand U835 (N_835,N_629,N_696);
and U836 (N_836,N_740,N_600);
or U837 (N_837,N_612,N_738);
and U838 (N_838,N_608,N_720);
nand U839 (N_839,N_695,N_680);
and U840 (N_840,N_707,N_686);
xor U841 (N_841,N_610,N_733);
nor U842 (N_842,N_797,N_735);
or U843 (N_843,N_622,N_617);
nor U844 (N_844,N_764,N_725);
and U845 (N_845,N_788,N_656);
and U846 (N_846,N_718,N_674);
nand U847 (N_847,N_663,N_779);
and U848 (N_848,N_691,N_778);
nor U849 (N_849,N_631,N_775);
and U850 (N_850,N_687,N_660);
nor U851 (N_851,N_602,N_621);
or U852 (N_852,N_623,N_605);
nand U853 (N_853,N_751,N_799);
and U854 (N_854,N_794,N_736);
or U855 (N_855,N_673,N_772);
nor U856 (N_856,N_668,N_706);
and U857 (N_857,N_755,N_759);
or U858 (N_858,N_726,N_625);
nor U859 (N_859,N_653,N_773);
or U860 (N_860,N_604,N_717);
or U861 (N_861,N_677,N_710);
nor U862 (N_862,N_783,N_620);
or U863 (N_863,N_732,N_636);
and U864 (N_864,N_715,N_650);
and U865 (N_865,N_628,N_763);
nand U866 (N_866,N_641,N_633);
or U867 (N_867,N_750,N_781);
or U868 (N_868,N_667,N_719);
nand U869 (N_869,N_705,N_637);
and U870 (N_870,N_679,N_640);
or U871 (N_871,N_609,N_787);
nor U872 (N_872,N_741,N_684);
or U873 (N_873,N_769,N_643);
nor U874 (N_874,N_642,N_683);
nor U875 (N_875,N_681,N_753);
nand U876 (N_876,N_748,N_765);
and U877 (N_877,N_747,N_664);
nand U878 (N_878,N_630,N_774);
or U879 (N_879,N_746,N_603);
and U880 (N_880,N_780,N_792);
nor U881 (N_881,N_743,N_757);
or U882 (N_882,N_651,N_611);
and U883 (N_883,N_762,N_688);
nor U884 (N_884,N_749,N_669);
or U885 (N_885,N_675,N_798);
or U886 (N_886,N_739,N_613);
nand U887 (N_887,N_776,N_729);
or U888 (N_888,N_607,N_770);
and U889 (N_889,N_652,N_635);
and U890 (N_890,N_796,N_716);
and U891 (N_891,N_756,N_722);
and U892 (N_892,N_662,N_689);
and U893 (N_893,N_702,N_760);
nor U894 (N_894,N_704,N_606);
nand U895 (N_895,N_734,N_627);
nand U896 (N_896,N_616,N_784);
or U897 (N_897,N_699,N_619);
or U898 (N_898,N_693,N_745);
and U899 (N_899,N_658,N_752);
xor U900 (N_900,N_755,N_752);
xnor U901 (N_901,N_772,N_712);
and U902 (N_902,N_680,N_734);
or U903 (N_903,N_627,N_780);
nor U904 (N_904,N_784,N_753);
and U905 (N_905,N_650,N_698);
nand U906 (N_906,N_722,N_690);
nor U907 (N_907,N_700,N_607);
and U908 (N_908,N_725,N_799);
nand U909 (N_909,N_601,N_730);
or U910 (N_910,N_661,N_666);
nand U911 (N_911,N_671,N_727);
and U912 (N_912,N_643,N_742);
or U913 (N_913,N_663,N_645);
nor U914 (N_914,N_795,N_739);
and U915 (N_915,N_607,N_610);
nor U916 (N_916,N_617,N_755);
or U917 (N_917,N_707,N_625);
nand U918 (N_918,N_606,N_696);
or U919 (N_919,N_747,N_658);
or U920 (N_920,N_773,N_600);
and U921 (N_921,N_632,N_676);
nand U922 (N_922,N_621,N_659);
and U923 (N_923,N_639,N_628);
nand U924 (N_924,N_673,N_768);
nand U925 (N_925,N_679,N_777);
nor U926 (N_926,N_781,N_744);
and U927 (N_927,N_666,N_626);
nor U928 (N_928,N_703,N_728);
or U929 (N_929,N_697,N_638);
nor U930 (N_930,N_756,N_604);
nand U931 (N_931,N_708,N_758);
or U932 (N_932,N_777,N_641);
nand U933 (N_933,N_716,N_612);
and U934 (N_934,N_763,N_632);
nor U935 (N_935,N_787,N_737);
nor U936 (N_936,N_786,N_602);
and U937 (N_937,N_610,N_655);
nand U938 (N_938,N_637,N_662);
and U939 (N_939,N_636,N_737);
and U940 (N_940,N_670,N_672);
or U941 (N_941,N_619,N_762);
and U942 (N_942,N_675,N_757);
or U943 (N_943,N_635,N_672);
or U944 (N_944,N_693,N_645);
and U945 (N_945,N_769,N_757);
nor U946 (N_946,N_652,N_778);
nor U947 (N_947,N_661,N_781);
or U948 (N_948,N_623,N_784);
nand U949 (N_949,N_631,N_607);
nor U950 (N_950,N_660,N_772);
nand U951 (N_951,N_722,N_656);
nor U952 (N_952,N_693,N_721);
nor U953 (N_953,N_622,N_609);
nand U954 (N_954,N_777,N_624);
and U955 (N_955,N_642,N_616);
or U956 (N_956,N_682,N_783);
nand U957 (N_957,N_710,N_688);
or U958 (N_958,N_713,N_698);
and U959 (N_959,N_758,N_761);
nand U960 (N_960,N_622,N_671);
nand U961 (N_961,N_789,N_746);
or U962 (N_962,N_721,N_681);
nand U963 (N_963,N_742,N_786);
or U964 (N_964,N_640,N_677);
and U965 (N_965,N_742,N_677);
and U966 (N_966,N_726,N_703);
or U967 (N_967,N_708,N_736);
or U968 (N_968,N_714,N_736);
nand U969 (N_969,N_636,N_683);
xnor U970 (N_970,N_642,N_757);
nand U971 (N_971,N_675,N_700);
and U972 (N_972,N_703,N_734);
or U973 (N_973,N_789,N_671);
or U974 (N_974,N_743,N_747);
and U975 (N_975,N_680,N_773);
or U976 (N_976,N_714,N_723);
nand U977 (N_977,N_609,N_702);
xnor U978 (N_978,N_768,N_737);
nor U979 (N_979,N_701,N_630);
nand U980 (N_980,N_642,N_778);
nand U981 (N_981,N_764,N_667);
nand U982 (N_982,N_668,N_633);
and U983 (N_983,N_669,N_686);
nand U984 (N_984,N_704,N_738);
or U985 (N_985,N_782,N_731);
and U986 (N_986,N_770,N_772);
nor U987 (N_987,N_616,N_718);
nand U988 (N_988,N_744,N_644);
or U989 (N_989,N_685,N_756);
nor U990 (N_990,N_662,N_619);
nand U991 (N_991,N_652,N_617);
and U992 (N_992,N_707,N_775);
or U993 (N_993,N_750,N_735);
and U994 (N_994,N_700,N_638);
nor U995 (N_995,N_629,N_725);
or U996 (N_996,N_778,N_722);
and U997 (N_997,N_649,N_674);
and U998 (N_998,N_690,N_675);
or U999 (N_999,N_739,N_774);
or U1000 (N_1000,N_871,N_997);
and U1001 (N_1001,N_942,N_807);
and U1002 (N_1002,N_994,N_901);
xnor U1003 (N_1003,N_861,N_813);
xor U1004 (N_1004,N_889,N_808);
or U1005 (N_1005,N_816,N_951);
and U1006 (N_1006,N_828,N_998);
nor U1007 (N_1007,N_982,N_983);
nand U1008 (N_1008,N_842,N_934);
nor U1009 (N_1009,N_995,N_905);
nor U1010 (N_1010,N_872,N_919);
or U1011 (N_1011,N_963,N_866);
or U1012 (N_1012,N_948,N_988);
and U1013 (N_1013,N_917,N_814);
or U1014 (N_1014,N_804,N_823);
and U1015 (N_1015,N_967,N_897);
nor U1016 (N_1016,N_817,N_910);
nand U1017 (N_1017,N_930,N_892);
nand U1018 (N_1018,N_932,N_939);
nor U1019 (N_1019,N_959,N_941);
nand U1020 (N_1020,N_975,N_940);
xor U1021 (N_1021,N_853,N_971);
nand U1022 (N_1022,N_890,N_943);
nand U1023 (N_1023,N_906,N_949);
nand U1024 (N_1024,N_887,N_805);
or U1025 (N_1025,N_830,N_916);
nand U1026 (N_1026,N_819,N_836);
nand U1027 (N_1027,N_914,N_978);
and U1028 (N_1028,N_874,N_815);
or U1029 (N_1029,N_829,N_857);
or U1030 (N_1030,N_809,N_841);
nand U1031 (N_1031,N_926,N_843);
or U1032 (N_1032,N_960,N_894);
nand U1033 (N_1033,N_947,N_979);
and U1034 (N_1034,N_863,N_945);
and U1035 (N_1035,N_803,N_875);
nand U1036 (N_1036,N_908,N_925);
nand U1037 (N_1037,N_800,N_810);
nand U1038 (N_1038,N_964,N_981);
nor U1039 (N_1039,N_920,N_922);
nor U1040 (N_1040,N_877,N_990);
or U1041 (N_1041,N_969,N_895);
nor U1042 (N_1042,N_958,N_848);
nor U1043 (N_1043,N_952,N_965);
nor U1044 (N_1044,N_953,N_844);
or U1045 (N_1045,N_986,N_899);
nor U1046 (N_1046,N_893,N_806);
nand U1047 (N_1047,N_931,N_865);
nand U1048 (N_1048,N_936,N_824);
and U1049 (N_1049,N_938,N_812);
or U1050 (N_1050,N_858,N_878);
nor U1051 (N_1051,N_825,N_838);
nand U1052 (N_1052,N_869,N_900);
or U1053 (N_1053,N_933,N_846);
or U1054 (N_1054,N_904,N_885);
and U1055 (N_1055,N_854,N_884);
or U1056 (N_1056,N_826,N_849);
or U1057 (N_1057,N_903,N_859);
nand U1058 (N_1058,N_862,N_973);
or U1059 (N_1059,N_851,N_977);
nand U1060 (N_1060,N_970,N_937);
and U1061 (N_1061,N_818,N_852);
or U1062 (N_1062,N_870,N_912);
nor U1063 (N_1063,N_944,N_840);
or U1064 (N_1064,N_911,N_927);
or U1065 (N_1065,N_909,N_837);
or U1066 (N_1066,N_820,N_915);
nand U1067 (N_1067,N_886,N_860);
or U1068 (N_1068,N_864,N_928);
or U1069 (N_1069,N_991,N_923);
nand U1070 (N_1070,N_883,N_822);
or U1071 (N_1071,N_989,N_856);
or U1072 (N_1072,N_888,N_831);
nor U1073 (N_1073,N_972,N_929);
and U1074 (N_1074,N_879,N_881);
or U1075 (N_1075,N_855,N_946);
and U1076 (N_1076,N_913,N_873);
xnor U1077 (N_1077,N_966,N_834);
nor U1078 (N_1078,N_876,N_867);
or U1079 (N_1079,N_801,N_868);
and U1080 (N_1080,N_999,N_850);
nand U1081 (N_1081,N_847,N_821);
and U1082 (N_1082,N_835,N_902);
and U1083 (N_1083,N_957,N_980);
nor U1084 (N_1084,N_962,N_811);
and U1085 (N_1085,N_992,N_845);
or U1086 (N_1086,N_896,N_918);
nor U1087 (N_1087,N_880,N_985);
nand U1088 (N_1088,N_907,N_987);
and U1089 (N_1089,N_935,N_921);
nor U1090 (N_1090,N_956,N_955);
nand U1091 (N_1091,N_976,N_832);
or U1092 (N_1092,N_891,N_898);
nor U1093 (N_1093,N_827,N_833);
nor U1094 (N_1094,N_954,N_984);
or U1095 (N_1095,N_839,N_802);
nand U1096 (N_1096,N_974,N_882);
nand U1097 (N_1097,N_924,N_961);
nand U1098 (N_1098,N_968,N_950);
or U1099 (N_1099,N_993,N_996);
and U1100 (N_1100,N_985,N_805);
or U1101 (N_1101,N_922,N_804);
nand U1102 (N_1102,N_948,N_846);
and U1103 (N_1103,N_886,N_997);
and U1104 (N_1104,N_978,N_822);
and U1105 (N_1105,N_863,N_970);
and U1106 (N_1106,N_976,N_815);
nand U1107 (N_1107,N_831,N_936);
nand U1108 (N_1108,N_897,N_800);
nand U1109 (N_1109,N_864,N_850);
nand U1110 (N_1110,N_818,N_809);
nand U1111 (N_1111,N_992,N_996);
or U1112 (N_1112,N_942,N_954);
or U1113 (N_1113,N_881,N_889);
nand U1114 (N_1114,N_931,N_851);
or U1115 (N_1115,N_809,N_907);
or U1116 (N_1116,N_817,N_848);
or U1117 (N_1117,N_881,N_890);
or U1118 (N_1118,N_826,N_981);
and U1119 (N_1119,N_987,N_802);
nand U1120 (N_1120,N_957,N_913);
nand U1121 (N_1121,N_851,N_994);
and U1122 (N_1122,N_893,N_903);
and U1123 (N_1123,N_844,N_827);
xnor U1124 (N_1124,N_867,N_886);
nand U1125 (N_1125,N_813,N_845);
or U1126 (N_1126,N_863,N_802);
nand U1127 (N_1127,N_863,N_867);
or U1128 (N_1128,N_864,N_888);
nor U1129 (N_1129,N_954,N_844);
and U1130 (N_1130,N_938,N_874);
nor U1131 (N_1131,N_972,N_800);
or U1132 (N_1132,N_916,N_839);
and U1133 (N_1133,N_854,N_952);
and U1134 (N_1134,N_941,N_948);
nand U1135 (N_1135,N_840,N_880);
xor U1136 (N_1136,N_947,N_927);
or U1137 (N_1137,N_895,N_842);
or U1138 (N_1138,N_908,N_924);
nand U1139 (N_1139,N_896,N_877);
or U1140 (N_1140,N_822,N_966);
nor U1141 (N_1141,N_851,N_949);
nand U1142 (N_1142,N_938,N_885);
nand U1143 (N_1143,N_834,N_859);
nand U1144 (N_1144,N_986,N_957);
and U1145 (N_1145,N_802,N_943);
nor U1146 (N_1146,N_923,N_899);
or U1147 (N_1147,N_927,N_969);
or U1148 (N_1148,N_970,N_945);
nor U1149 (N_1149,N_974,N_819);
or U1150 (N_1150,N_955,N_803);
and U1151 (N_1151,N_964,N_903);
or U1152 (N_1152,N_812,N_883);
nor U1153 (N_1153,N_869,N_862);
nor U1154 (N_1154,N_837,N_880);
or U1155 (N_1155,N_878,N_900);
nor U1156 (N_1156,N_821,N_997);
and U1157 (N_1157,N_920,N_930);
nor U1158 (N_1158,N_865,N_926);
xor U1159 (N_1159,N_999,N_961);
or U1160 (N_1160,N_987,N_939);
or U1161 (N_1161,N_960,N_889);
nor U1162 (N_1162,N_859,N_809);
nand U1163 (N_1163,N_902,N_970);
nor U1164 (N_1164,N_896,N_843);
and U1165 (N_1165,N_950,N_831);
and U1166 (N_1166,N_821,N_834);
nor U1167 (N_1167,N_963,N_973);
or U1168 (N_1168,N_996,N_930);
or U1169 (N_1169,N_806,N_908);
xnor U1170 (N_1170,N_846,N_868);
and U1171 (N_1171,N_926,N_930);
nor U1172 (N_1172,N_929,N_852);
or U1173 (N_1173,N_840,N_951);
nor U1174 (N_1174,N_905,N_922);
nand U1175 (N_1175,N_918,N_872);
nor U1176 (N_1176,N_819,N_821);
nor U1177 (N_1177,N_967,N_922);
and U1178 (N_1178,N_959,N_808);
nor U1179 (N_1179,N_858,N_907);
or U1180 (N_1180,N_893,N_883);
and U1181 (N_1181,N_852,N_840);
nand U1182 (N_1182,N_983,N_990);
nor U1183 (N_1183,N_882,N_856);
nand U1184 (N_1184,N_892,N_981);
xor U1185 (N_1185,N_828,N_801);
nor U1186 (N_1186,N_987,N_949);
nand U1187 (N_1187,N_801,N_962);
or U1188 (N_1188,N_885,N_871);
or U1189 (N_1189,N_950,N_930);
nand U1190 (N_1190,N_834,N_857);
and U1191 (N_1191,N_851,N_892);
or U1192 (N_1192,N_977,N_926);
nand U1193 (N_1193,N_915,N_923);
or U1194 (N_1194,N_968,N_897);
or U1195 (N_1195,N_912,N_923);
and U1196 (N_1196,N_829,N_813);
and U1197 (N_1197,N_956,N_808);
and U1198 (N_1198,N_836,N_864);
nand U1199 (N_1199,N_971,N_935);
nand U1200 (N_1200,N_1091,N_1142);
nand U1201 (N_1201,N_1051,N_1013);
or U1202 (N_1202,N_1009,N_1116);
and U1203 (N_1203,N_1169,N_1043);
and U1204 (N_1204,N_1149,N_1045);
nor U1205 (N_1205,N_1153,N_1016);
nand U1206 (N_1206,N_1165,N_1038);
or U1207 (N_1207,N_1133,N_1088);
xor U1208 (N_1208,N_1176,N_1046);
and U1209 (N_1209,N_1121,N_1030);
nand U1210 (N_1210,N_1053,N_1063);
and U1211 (N_1211,N_1190,N_1044);
nand U1212 (N_1212,N_1001,N_1035);
xnor U1213 (N_1213,N_1093,N_1011);
nand U1214 (N_1214,N_1168,N_1156);
xor U1215 (N_1215,N_1171,N_1104);
nor U1216 (N_1216,N_1005,N_1058);
nor U1217 (N_1217,N_1074,N_1070);
nand U1218 (N_1218,N_1055,N_1184);
and U1219 (N_1219,N_1188,N_1081);
nand U1220 (N_1220,N_1015,N_1049);
nor U1221 (N_1221,N_1021,N_1075);
or U1222 (N_1222,N_1034,N_1130);
nor U1223 (N_1223,N_1199,N_1109);
or U1224 (N_1224,N_1019,N_1177);
xor U1225 (N_1225,N_1164,N_1112);
nor U1226 (N_1226,N_1098,N_1192);
and U1227 (N_1227,N_1159,N_1064);
nand U1228 (N_1228,N_1067,N_1024);
and U1229 (N_1229,N_1111,N_1071);
and U1230 (N_1230,N_1061,N_1079);
nor U1231 (N_1231,N_1148,N_1134);
nor U1232 (N_1232,N_1196,N_1185);
nand U1233 (N_1233,N_1180,N_1131);
nor U1234 (N_1234,N_1060,N_1135);
or U1235 (N_1235,N_1107,N_1124);
nand U1236 (N_1236,N_1052,N_1047);
nor U1237 (N_1237,N_1189,N_1191);
and U1238 (N_1238,N_1096,N_1139);
nand U1239 (N_1239,N_1007,N_1150);
nor U1240 (N_1240,N_1087,N_1160);
or U1241 (N_1241,N_1161,N_1042);
nand U1242 (N_1242,N_1078,N_1017);
and U1243 (N_1243,N_1039,N_1028);
or U1244 (N_1244,N_1105,N_1186);
or U1245 (N_1245,N_1167,N_1158);
and U1246 (N_1246,N_1118,N_1122);
nor U1247 (N_1247,N_1166,N_1033);
nand U1248 (N_1248,N_1173,N_1018);
or U1249 (N_1249,N_1100,N_1140);
nand U1250 (N_1250,N_1006,N_1179);
and U1251 (N_1251,N_1069,N_1012);
nand U1252 (N_1252,N_1084,N_1141);
nor U1253 (N_1253,N_1066,N_1023);
nor U1254 (N_1254,N_1117,N_1114);
nand U1255 (N_1255,N_1125,N_1086);
nor U1256 (N_1256,N_1092,N_1065);
and U1257 (N_1257,N_1126,N_1050);
or U1258 (N_1258,N_1103,N_1123);
xnor U1259 (N_1259,N_1073,N_1082);
nand U1260 (N_1260,N_1041,N_1032);
xor U1261 (N_1261,N_1110,N_1094);
or U1262 (N_1262,N_1068,N_1095);
or U1263 (N_1263,N_1193,N_1002);
xor U1264 (N_1264,N_1195,N_1090);
nor U1265 (N_1265,N_1197,N_1027);
and U1266 (N_1266,N_1025,N_1144);
and U1267 (N_1267,N_1108,N_1182);
nand U1268 (N_1268,N_1020,N_1054);
nand U1269 (N_1269,N_1022,N_1194);
nor U1270 (N_1270,N_1057,N_1031);
nor U1271 (N_1271,N_1136,N_1101);
and U1272 (N_1272,N_1099,N_1026);
nor U1273 (N_1273,N_1062,N_1138);
nor U1274 (N_1274,N_1040,N_1056);
nor U1275 (N_1275,N_1172,N_1076);
nand U1276 (N_1276,N_1119,N_1102);
nand U1277 (N_1277,N_1154,N_1128);
or U1278 (N_1278,N_1151,N_1077);
nor U1279 (N_1279,N_1163,N_1113);
nor U1280 (N_1280,N_1187,N_1162);
nand U1281 (N_1281,N_1036,N_1059);
nor U1282 (N_1282,N_1175,N_1029);
nor U1283 (N_1283,N_1198,N_1129);
nor U1284 (N_1284,N_1120,N_1147);
nor U1285 (N_1285,N_1000,N_1127);
nand U1286 (N_1286,N_1170,N_1003);
or U1287 (N_1287,N_1072,N_1106);
or U1288 (N_1288,N_1083,N_1146);
nand U1289 (N_1289,N_1155,N_1174);
and U1290 (N_1290,N_1080,N_1014);
or U1291 (N_1291,N_1157,N_1085);
or U1292 (N_1292,N_1115,N_1137);
nor U1293 (N_1293,N_1183,N_1132);
nand U1294 (N_1294,N_1010,N_1152);
xnor U1295 (N_1295,N_1008,N_1097);
nand U1296 (N_1296,N_1089,N_1143);
or U1297 (N_1297,N_1178,N_1181);
nor U1298 (N_1298,N_1145,N_1004);
or U1299 (N_1299,N_1037,N_1048);
nand U1300 (N_1300,N_1143,N_1174);
and U1301 (N_1301,N_1021,N_1197);
nor U1302 (N_1302,N_1179,N_1019);
nand U1303 (N_1303,N_1064,N_1140);
nor U1304 (N_1304,N_1126,N_1183);
nand U1305 (N_1305,N_1198,N_1023);
or U1306 (N_1306,N_1013,N_1135);
nand U1307 (N_1307,N_1114,N_1034);
and U1308 (N_1308,N_1140,N_1004);
or U1309 (N_1309,N_1047,N_1034);
and U1310 (N_1310,N_1172,N_1074);
nand U1311 (N_1311,N_1059,N_1018);
or U1312 (N_1312,N_1185,N_1153);
and U1313 (N_1313,N_1193,N_1059);
or U1314 (N_1314,N_1115,N_1131);
nand U1315 (N_1315,N_1089,N_1003);
or U1316 (N_1316,N_1027,N_1083);
and U1317 (N_1317,N_1024,N_1057);
or U1318 (N_1318,N_1057,N_1198);
nor U1319 (N_1319,N_1139,N_1037);
nor U1320 (N_1320,N_1132,N_1002);
nor U1321 (N_1321,N_1028,N_1162);
and U1322 (N_1322,N_1116,N_1199);
and U1323 (N_1323,N_1130,N_1102);
nand U1324 (N_1324,N_1146,N_1141);
nand U1325 (N_1325,N_1041,N_1138);
or U1326 (N_1326,N_1117,N_1182);
xnor U1327 (N_1327,N_1085,N_1127);
and U1328 (N_1328,N_1174,N_1060);
xor U1329 (N_1329,N_1099,N_1069);
and U1330 (N_1330,N_1079,N_1087);
and U1331 (N_1331,N_1181,N_1092);
or U1332 (N_1332,N_1064,N_1122);
and U1333 (N_1333,N_1051,N_1075);
and U1334 (N_1334,N_1125,N_1123);
nor U1335 (N_1335,N_1101,N_1056);
or U1336 (N_1336,N_1183,N_1192);
nor U1337 (N_1337,N_1168,N_1157);
and U1338 (N_1338,N_1189,N_1175);
or U1339 (N_1339,N_1000,N_1141);
nand U1340 (N_1340,N_1081,N_1101);
nor U1341 (N_1341,N_1089,N_1046);
nor U1342 (N_1342,N_1143,N_1117);
nand U1343 (N_1343,N_1018,N_1144);
xnor U1344 (N_1344,N_1169,N_1165);
or U1345 (N_1345,N_1058,N_1156);
or U1346 (N_1346,N_1061,N_1180);
and U1347 (N_1347,N_1026,N_1116);
or U1348 (N_1348,N_1088,N_1158);
or U1349 (N_1349,N_1091,N_1174);
or U1350 (N_1350,N_1008,N_1186);
nand U1351 (N_1351,N_1070,N_1183);
nand U1352 (N_1352,N_1091,N_1071);
or U1353 (N_1353,N_1120,N_1080);
and U1354 (N_1354,N_1138,N_1092);
nand U1355 (N_1355,N_1161,N_1009);
and U1356 (N_1356,N_1076,N_1158);
nand U1357 (N_1357,N_1152,N_1137);
and U1358 (N_1358,N_1197,N_1091);
or U1359 (N_1359,N_1084,N_1153);
nor U1360 (N_1360,N_1100,N_1005);
nand U1361 (N_1361,N_1034,N_1019);
xor U1362 (N_1362,N_1030,N_1154);
or U1363 (N_1363,N_1193,N_1178);
nor U1364 (N_1364,N_1034,N_1057);
and U1365 (N_1365,N_1039,N_1166);
and U1366 (N_1366,N_1024,N_1046);
or U1367 (N_1367,N_1107,N_1021);
nor U1368 (N_1368,N_1078,N_1029);
nor U1369 (N_1369,N_1189,N_1018);
and U1370 (N_1370,N_1029,N_1063);
and U1371 (N_1371,N_1145,N_1106);
or U1372 (N_1372,N_1030,N_1182);
and U1373 (N_1373,N_1138,N_1184);
nor U1374 (N_1374,N_1127,N_1105);
and U1375 (N_1375,N_1042,N_1011);
and U1376 (N_1376,N_1151,N_1034);
nor U1377 (N_1377,N_1084,N_1119);
nor U1378 (N_1378,N_1169,N_1109);
nor U1379 (N_1379,N_1067,N_1018);
xnor U1380 (N_1380,N_1147,N_1031);
and U1381 (N_1381,N_1115,N_1067);
and U1382 (N_1382,N_1051,N_1138);
nand U1383 (N_1383,N_1092,N_1158);
nor U1384 (N_1384,N_1021,N_1161);
nand U1385 (N_1385,N_1173,N_1147);
nor U1386 (N_1386,N_1183,N_1082);
nand U1387 (N_1387,N_1101,N_1068);
and U1388 (N_1388,N_1198,N_1096);
nor U1389 (N_1389,N_1001,N_1122);
nor U1390 (N_1390,N_1061,N_1073);
nor U1391 (N_1391,N_1189,N_1176);
nand U1392 (N_1392,N_1064,N_1196);
nand U1393 (N_1393,N_1154,N_1185);
nand U1394 (N_1394,N_1112,N_1116);
and U1395 (N_1395,N_1106,N_1096);
nand U1396 (N_1396,N_1087,N_1012);
and U1397 (N_1397,N_1169,N_1148);
and U1398 (N_1398,N_1002,N_1175);
nor U1399 (N_1399,N_1102,N_1121);
nor U1400 (N_1400,N_1238,N_1375);
and U1401 (N_1401,N_1202,N_1330);
nand U1402 (N_1402,N_1343,N_1248);
and U1403 (N_1403,N_1292,N_1203);
nor U1404 (N_1404,N_1295,N_1313);
nor U1405 (N_1405,N_1241,N_1372);
nor U1406 (N_1406,N_1322,N_1383);
nand U1407 (N_1407,N_1337,N_1321);
nor U1408 (N_1408,N_1293,N_1351);
or U1409 (N_1409,N_1266,N_1365);
nor U1410 (N_1410,N_1256,N_1288);
xnor U1411 (N_1411,N_1396,N_1304);
nor U1412 (N_1412,N_1283,N_1220);
or U1413 (N_1413,N_1234,N_1356);
and U1414 (N_1414,N_1331,N_1391);
nand U1415 (N_1415,N_1252,N_1328);
nor U1416 (N_1416,N_1346,N_1291);
and U1417 (N_1417,N_1214,N_1382);
or U1418 (N_1418,N_1260,N_1355);
and U1419 (N_1419,N_1385,N_1341);
nand U1420 (N_1420,N_1389,N_1222);
and U1421 (N_1421,N_1251,N_1349);
nor U1422 (N_1422,N_1231,N_1243);
or U1423 (N_1423,N_1395,N_1239);
nor U1424 (N_1424,N_1399,N_1212);
nand U1425 (N_1425,N_1297,N_1338);
nand U1426 (N_1426,N_1388,N_1277);
xnor U1427 (N_1427,N_1370,N_1289);
nor U1428 (N_1428,N_1264,N_1254);
nor U1429 (N_1429,N_1270,N_1242);
or U1430 (N_1430,N_1369,N_1285);
nand U1431 (N_1431,N_1280,N_1250);
or U1432 (N_1432,N_1275,N_1324);
xnor U1433 (N_1433,N_1235,N_1310);
nand U1434 (N_1434,N_1286,N_1317);
nor U1435 (N_1435,N_1348,N_1249);
nand U1436 (N_1436,N_1281,N_1368);
nand U1437 (N_1437,N_1378,N_1269);
nor U1438 (N_1438,N_1230,N_1255);
xnor U1439 (N_1439,N_1263,N_1287);
nand U1440 (N_1440,N_1237,N_1229);
and U1441 (N_1441,N_1332,N_1279);
and U1442 (N_1442,N_1367,N_1381);
and U1443 (N_1443,N_1278,N_1205);
or U1444 (N_1444,N_1392,N_1209);
or U1445 (N_1445,N_1300,N_1232);
or U1446 (N_1446,N_1312,N_1350);
nand U1447 (N_1447,N_1345,N_1262);
and U1448 (N_1448,N_1236,N_1299);
or U1449 (N_1449,N_1276,N_1353);
and U1450 (N_1450,N_1366,N_1354);
nand U1451 (N_1451,N_1327,N_1342);
nand U1452 (N_1452,N_1397,N_1224);
nand U1453 (N_1453,N_1273,N_1318);
or U1454 (N_1454,N_1240,N_1233);
and U1455 (N_1455,N_1210,N_1225);
and U1456 (N_1456,N_1207,N_1267);
and U1457 (N_1457,N_1221,N_1290);
nor U1458 (N_1458,N_1352,N_1258);
xor U1459 (N_1459,N_1364,N_1272);
nor U1460 (N_1460,N_1259,N_1393);
and U1461 (N_1461,N_1315,N_1371);
nand U1462 (N_1462,N_1308,N_1340);
nand U1463 (N_1463,N_1336,N_1306);
and U1464 (N_1464,N_1326,N_1215);
or U1465 (N_1465,N_1363,N_1329);
and U1466 (N_1466,N_1339,N_1211);
and U1467 (N_1467,N_1380,N_1379);
or U1468 (N_1468,N_1325,N_1374);
or U1469 (N_1469,N_1386,N_1314);
nand U1470 (N_1470,N_1303,N_1216);
and U1471 (N_1471,N_1390,N_1257);
or U1472 (N_1472,N_1357,N_1245);
nor U1473 (N_1473,N_1323,N_1309);
nor U1474 (N_1474,N_1347,N_1261);
or U1475 (N_1475,N_1228,N_1274);
nand U1476 (N_1476,N_1227,N_1282);
nand U1477 (N_1477,N_1398,N_1246);
nor U1478 (N_1478,N_1384,N_1359);
nand U1479 (N_1479,N_1284,N_1387);
xnor U1480 (N_1480,N_1361,N_1294);
nand U1481 (N_1481,N_1296,N_1394);
and U1482 (N_1482,N_1223,N_1244);
and U1483 (N_1483,N_1358,N_1206);
or U1484 (N_1484,N_1302,N_1362);
or U1485 (N_1485,N_1301,N_1219);
nand U1486 (N_1486,N_1333,N_1200);
nor U1487 (N_1487,N_1217,N_1268);
nor U1488 (N_1488,N_1298,N_1204);
nor U1489 (N_1489,N_1344,N_1335);
and U1490 (N_1490,N_1201,N_1311);
xnor U1491 (N_1491,N_1271,N_1213);
nand U1492 (N_1492,N_1208,N_1218);
nand U1493 (N_1493,N_1307,N_1373);
nand U1494 (N_1494,N_1334,N_1377);
and U1495 (N_1495,N_1265,N_1316);
or U1496 (N_1496,N_1376,N_1253);
nor U1497 (N_1497,N_1305,N_1319);
nor U1498 (N_1498,N_1247,N_1360);
nor U1499 (N_1499,N_1320,N_1226);
nor U1500 (N_1500,N_1360,N_1214);
nand U1501 (N_1501,N_1345,N_1351);
or U1502 (N_1502,N_1229,N_1316);
and U1503 (N_1503,N_1386,N_1266);
nor U1504 (N_1504,N_1354,N_1353);
nor U1505 (N_1505,N_1254,N_1207);
or U1506 (N_1506,N_1386,N_1385);
or U1507 (N_1507,N_1202,N_1203);
xor U1508 (N_1508,N_1261,N_1262);
nor U1509 (N_1509,N_1293,N_1223);
nor U1510 (N_1510,N_1349,N_1240);
or U1511 (N_1511,N_1254,N_1302);
and U1512 (N_1512,N_1214,N_1294);
and U1513 (N_1513,N_1240,N_1253);
or U1514 (N_1514,N_1319,N_1223);
nor U1515 (N_1515,N_1310,N_1331);
and U1516 (N_1516,N_1379,N_1216);
or U1517 (N_1517,N_1289,N_1368);
or U1518 (N_1518,N_1257,N_1332);
nand U1519 (N_1519,N_1381,N_1264);
or U1520 (N_1520,N_1355,N_1300);
nor U1521 (N_1521,N_1358,N_1242);
nand U1522 (N_1522,N_1329,N_1210);
nor U1523 (N_1523,N_1252,N_1324);
and U1524 (N_1524,N_1217,N_1227);
nand U1525 (N_1525,N_1309,N_1317);
nor U1526 (N_1526,N_1233,N_1280);
and U1527 (N_1527,N_1251,N_1270);
or U1528 (N_1528,N_1202,N_1363);
nand U1529 (N_1529,N_1334,N_1273);
or U1530 (N_1530,N_1287,N_1240);
nand U1531 (N_1531,N_1316,N_1354);
and U1532 (N_1532,N_1246,N_1282);
xnor U1533 (N_1533,N_1357,N_1206);
nand U1534 (N_1534,N_1387,N_1301);
nand U1535 (N_1535,N_1219,N_1261);
nand U1536 (N_1536,N_1251,N_1357);
and U1537 (N_1537,N_1293,N_1330);
nor U1538 (N_1538,N_1321,N_1360);
and U1539 (N_1539,N_1282,N_1294);
and U1540 (N_1540,N_1217,N_1322);
nand U1541 (N_1541,N_1260,N_1367);
and U1542 (N_1542,N_1312,N_1238);
or U1543 (N_1543,N_1383,N_1291);
nor U1544 (N_1544,N_1355,N_1357);
nand U1545 (N_1545,N_1361,N_1355);
and U1546 (N_1546,N_1236,N_1391);
or U1547 (N_1547,N_1367,N_1224);
and U1548 (N_1548,N_1284,N_1287);
or U1549 (N_1549,N_1322,N_1315);
or U1550 (N_1550,N_1385,N_1351);
and U1551 (N_1551,N_1221,N_1363);
or U1552 (N_1552,N_1374,N_1221);
nor U1553 (N_1553,N_1262,N_1342);
xnor U1554 (N_1554,N_1282,N_1363);
nand U1555 (N_1555,N_1287,N_1388);
or U1556 (N_1556,N_1269,N_1262);
xnor U1557 (N_1557,N_1397,N_1271);
nor U1558 (N_1558,N_1307,N_1257);
nand U1559 (N_1559,N_1317,N_1354);
or U1560 (N_1560,N_1268,N_1334);
and U1561 (N_1561,N_1306,N_1391);
nand U1562 (N_1562,N_1304,N_1359);
or U1563 (N_1563,N_1222,N_1312);
nand U1564 (N_1564,N_1373,N_1313);
and U1565 (N_1565,N_1319,N_1337);
and U1566 (N_1566,N_1331,N_1293);
nand U1567 (N_1567,N_1220,N_1258);
or U1568 (N_1568,N_1273,N_1251);
and U1569 (N_1569,N_1394,N_1289);
nand U1570 (N_1570,N_1244,N_1286);
nor U1571 (N_1571,N_1246,N_1342);
or U1572 (N_1572,N_1206,N_1257);
xnor U1573 (N_1573,N_1314,N_1200);
or U1574 (N_1574,N_1224,N_1207);
nand U1575 (N_1575,N_1294,N_1337);
nand U1576 (N_1576,N_1393,N_1323);
nor U1577 (N_1577,N_1230,N_1384);
and U1578 (N_1578,N_1273,N_1366);
nor U1579 (N_1579,N_1303,N_1282);
nand U1580 (N_1580,N_1397,N_1392);
nor U1581 (N_1581,N_1286,N_1283);
nand U1582 (N_1582,N_1357,N_1200);
and U1583 (N_1583,N_1231,N_1378);
or U1584 (N_1584,N_1396,N_1307);
and U1585 (N_1585,N_1356,N_1289);
nand U1586 (N_1586,N_1219,N_1300);
nand U1587 (N_1587,N_1315,N_1289);
and U1588 (N_1588,N_1393,N_1394);
and U1589 (N_1589,N_1396,N_1224);
nand U1590 (N_1590,N_1371,N_1272);
xor U1591 (N_1591,N_1267,N_1378);
or U1592 (N_1592,N_1371,N_1245);
nor U1593 (N_1593,N_1369,N_1333);
or U1594 (N_1594,N_1374,N_1314);
nand U1595 (N_1595,N_1366,N_1397);
nor U1596 (N_1596,N_1250,N_1218);
nor U1597 (N_1597,N_1293,N_1270);
and U1598 (N_1598,N_1351,N_1360);
or U1599 (N_1599,N_1244,N_1218);
or U1600 (N_1600,N_1582,N_1487);
and U1601 (N_1601,N_1496,N_1428);
or U1602 (N_1602,N_1546,N_1598);
or U1603 (N_1603,N_1436,N_1540);
nor U1604 (N_1604,N_1505,N_1574);
nor U1605 (N_1605,N_1541,N_1431);
and U1606 (N_1606,N_1458,N_1473);
or U1607 (N_1607,N_1561,N_1575);
nor U1608 (N_1608,N_1430,N_1572);
and U1609 (N_1609,N_1414,N_1420);
and U1610 (N_1610,N_1450,N_1417);
or U1611 (N_1611,N_1587,N_1583);
nand U1612 (N_1612,N_1599,N_1509);
or U1613 (N_1613,N_1443,N_1565);
and U1614 (N_1614,N_1454,N_1516);
nor U1615 (N_1615,N_1491,N_1567);
and U1616 (N_1616,N_1478,N_1493);
nand U1617 (N_1617,N_1468,N_1477);
and U1618 (N_1618,N_1498,N_1576);
or U1619 (N_1619,N_1453,N_1515);
nor U1620 (N_1620,N_1560,N_1568);
nand U1621 (N_1621,N_1497,N_1494);
nor U1622 (N_1622,N_1472,N_1533);
and U1623 (N_1623,N_1595,N_1554);
nand U1624 (N_1624,N_1528,N_1558);
nand U1625 (N_1625,N_1525,N_1448);
nand U1626 (N_1626,N_1427,N_1482);
nand U1627 (N_1627,N_1407,N_1523);
nand U1628 (N_1628,N_1594,N_1511);
nand U1629 (N_1629,N_1530,N_1542);
nand U1630 (N_1630,N_1463,N_1518);
nor U1631 (N_1631,N_1578,N_1492);
and U1632 (N_1632,N_1481,N_1597);
and U1633 (N_1633,N_1429,N_1421);
nor U1634 (N_1634,N_1466,N_1504);
and U1635 (N_1635,N_1566,N_1461);
and U1636 (N_1636,N_1571,N_1513);
nand U1637 (N_1637,N_1545,N_1527);
or U1638 (N_1638,N_1418,N_1562);
or U1639 (N_1639,N_1474,N_1438);
nand U1640 (N_1640,N_1520,N_1410);
nor U1641 (N_1641,N_1586,N_1537);
or U1642 (N_1642,N_1544,N_1532);
and U1643 (N_1643,N_1547,N_1507);
nor U1644 (N_1644,N_1512,N_1593);
nand U1645 (N_1645,N_1579,N_1549);
and U1646 (N_1646,N_1510,N_1415);
nand U1647 (N_1647,N_1551,N_1488);
nand U1648 (N_1648,N_1423,N_1591);
nand U1649 (N_1649,N_1441,N_1413);
and U1650 (N_1650,N_1573,N_1419);
nand U1651 (N_1651,N_1535,N_1529);
nor U1652 (N_1652,N_1548,N_1440);
or U1653 (N_1653,N_1403,N_1452);
or U1654 (N_1654,N_1500,N_1451);
and U1655 (N_1655,N_1499,N_1552);
or U1656 (N_1656,N_1464,N_1449);
xnor U1657 (N_1657,N_1405,N_1506);
nor U1658 (N_1658,N_1495,N_1580);
and U1659 (N_1659,N_1485,N_1435);
nand U1660 (N_1660,N_1471,N_1408);
nand U1661 (N_1661,N_1483,N_1534);
nand U1662 (N_1662,N_1588,N_1457);
nand U1663 (N_1663,N_1446,N_1445);
or U1664 (N_1664,N_1589,N_1592);
or U1665 (N_1665,N_1432,N_1536);
and U1666 (N_1666,N_1412,N_1437);
and U1667 (N_1667,N_1460,N_1459);
nand U1668 (N_1668,N_1411,N_1503);
nand U1669 (N_1669,N_1401,N_1508);
nand U1670 (N_1670,N_1563,N_1590);
and U1671 (N_1671,N_1426,N_1559);
nor U1672 (N_1672,N_1462,N_1486);
nand U1673 (N_1673,N_1434,N_1501);
nand U1674 (N_1674,N_1425,N_1400);
nand U1675 (N_1675,N_1455,N_1479);
nand U1676 (N_1676,N_1553,N_1465);
xnor U1677 (N_1677,N_1584,N_1475);
or U1678 (N_1678,N_1539,N_1480);
or U1679 (N_1679,N_1402,N_1524);
nor U1680 (N_1680,N_1422,N_1521);
and U1681 (N_1681,N_1433,N_1538);
nand U1682 (N_1682,N_1404,N_1556);
or U1683 (N_1683,N_1519,N_1447);
and U1684 (N_1684,N_1557,N_1531);
or U1685 (N_1685,N_1543,N_1489);
nand U1686 (N_1686,N_1550,N_1469);
nor U1687 (N_1687,N_1424,N_1502);
or U1688 (N_1688,N_1476,N_1596);
or U1689 (N_1689,N_1416,N_1442);
nand U1690 (N_1690,N_1409,N_1581);
nor U1691 (N_1691,N_1526,N_1514);
nand U1692 (N_1692,N_1467,N_1484);
or U1693 (N_1693,N_1490,N_1522);
nand U1694 (N_1694,N_1439,N_1570);
nor U1695 (N_1695,N_1517,N_1470);
xor U1696 (N_1696,N_1577,N_1555);
or U1697 (N_1697,N_1406,N_1585);
nor U1698 (N_1698,N_1564,N_1569);
nand U1699 (N_1699,N_1456,N_1444);
or U1700 (N_1700,N_1529,N_1478);
nand U1701 (N_1701,N_1589,N_1584);
nand U1702 (N_1702,N_1585,N_1557);
nor U1703 (N_1703,N_1594,N_1473);
or U1704 (N_1704,N_1421,N_1458);
nand U1705 (N_1705,N_1544,N_1535);
xor U1706 (N_1706,N_1493,N_1445);
or U1707 (N_1707,N_1431,N_1587);
or U1708 (N_1708,N_1439,N_1583);
nor U1709 (N_1709,N_1536,N_1555);
nand U1710 (N_1710,N_1498,N_1483);
or U1711 (N_1711,N_1512,N_1525);
nor U1712 (N_1712,N_1455,N_1489);
nand U1713 (N_1713,N_1409,N_1512);
or U1714 (N_1714,N_1491,N_1407);
nand U1715 (N_1715,N_1508,N_1480);
and U1716 (N_1716,N_1407,N_1582);
and U1717 (N_1717,N_1534,N_1570);
nand U1718 (N_1718,N_1418,N_1405);
nor U1719 (N_1719,N_1552,N_1563);
and U1720 (N_1720,N_1524,N_1492);
and U1721 (N_1721,N_1514,N_1597);
or U1722 (N_1722,N_1403,N_1546);
and U1723 (N_1723,N_1468,N_1455);
nor U1724 (N_1724,N_1579,N_1458);
nor U1725 (N_1725,N_1528,N_1409);
or U1726 (N_1726,N_1540,N_1558);
nand U1727 (N_1727,N_1553,N_1524);
or U1728 (N_1728,N_1570,N_1499);
nor U1729 (N_1729,N_1570,N_1483);
xnor U1730 (N_1730,N_1456,N_1405);
and U1731 (N_1731,N_1583,N_1585);
and U1732 (N_1732,N_1406,N_1407);
nand U1733 (N_1733,N_1564,N_1521);
nand U1734 (N_1734,N_1434,N_1516);
and U1735 (N_1735,N_1443,N_1559);
nand U1736 (N_1736,N_1509,N_1448);
or U1737 (N_1737,N_1478,N_1448);
or U1738 (N_1738,N_1543,N_1555);
nor U1739 (N_1739,N_1455,N_1472);
nor U1740 (N_1740,N_1597,N_1592);
nor U1741 (N_1741,N_1474,N_1486);
and U1742 (N_1742,N_1514,N_1437);
nand U1743 (N_1743,N_1544,N_1519);
or U1744 (N_1744,N_1424,N_1418);
or U1745 (N_1745,N_1449,N_1570);
or U1746 (N_1746,N_1552,N_1525);
nor U1747 (N_1747,N_1416,N_1530);
nand U1748 (N_1748,N_1488,N_1592);
nor U1749 (N_1749,N_1544,N_1524);
nand U1750 (N_1750,N_1455,N_1575);
and U1751 (N_1751,N_1443,N_1510);
nor U1752 (N_1752,N_1437,N_1489);
nand U1753 (N_1753,N_1568,N_1451);
or U1754 (N_1754,N_1486,N_1502);
and U1755 (N_1755,N_1508,N_1499);
nor U1756 (N_1756,N_1452,N_1542);
and U1757 (N_1757,N_1598,N_1539);
or U1758 (N_1758,N_1468,N_1404);
nand U1759 (N_1759,N_1484,N_1411);
and U1760 (N_1760,N_1407,N_1497);
nor U1761 (N_1761,N_1512,N_1480);
nor U1762 (N_1762,N_1541,N_1509);
nand U1763 (N_1763,N_1419,N_1579);
nand U1764 (N_1764,N_1516,N_1407);
nor U1765 (N_1765,N_1596,N_1495);
or U1766 (N_1766,N_1467,N_1547);
or U1767 (N_1767,N_1593,N_1463);
xor U1768 (N_1768,N_1483,N_1460);
and U1769 (N_1769,N_1536,N_1469);
nand U1770 (N_1770,N_1419,N_1431);
nand U1771 (N_1771,N_1452,N_1431);
and U1772 (N_1772,N_1437,N_1562);
or U1773 (N_1773,N_1482,N_1433);
or U1774 (N_1774,N_1507,N_1402);
nor U1775 (N_1775,N_1571,N_1496);
and U1776 (N_1776,N_1513,N_1546);
nor U1777 (N_1777,N_1581,N_1445);
and U1778 (N_1778,N_1537,N_1552);
and U1779 (N_1779,N_1599,N_1426);
nor U1780 (N_1780,N_1480,N_1450);
nor U1781 (N_1781,N_1503,N_1536);
and U1782 (N_1782,N_1572,N_1530);
nor U1783 (N_1783,N_1447,N_1458);
nand U1784 (N_1784,N_1448,N_1575);
and U1785 (N_1785,N_1595,N_1443);
nand U1786 (N_1786,N_1528,N_1435);
nand U1787 (N_1787,N_1529,N_1470);
nand U1788 (N_1788,N_1546,N_1578);
nor U1789 (N_1789,N_1413,N_1529);
or U1790 (N_1790,N_1513,N_1548);
nor U1791 (N_1791,N_1428,N_1422);
nand U1792 (N_1792,N_1591,N_1532);
or U1793 (N_1793,N_1403,N_1565);
and U1794 (N_1794,N_1545,N_1478);
and U1795 (N_1795,N_1455,N_1430);
nand U1796 (N_1796,N_1509,N_1434);
and U1797 (N_1797,N_1410,N_1504);
and U1798 (N_1798,N_1441,N_1427);
nor U1799 (N_1799,N_1413,N_1516);
or U1800 (N_1800,N_1798,N_1615);
or U1801 (N_1801,N_1737,N_1725);
nor U1802 (N_1802,N_1670,N_1696);
and U1803 (N_1803,N_1671,N_1713);
and U1804 (N_1804,N_1754,N_1767);
nor U1805 (N_1805,N_1699,N_1739);
nor U1806 (N_1806,N_1619,N_1632);
and U1807 (N_1807,N_1637,N_1784);
and U1808 (N_1808,N_1766,N_1789);
and U1809 (N_1809,N_1674,N_1622);
nor U1810 (N_1810,N_1773,N_1662);
nor U1811 (N_1811,N_1608,N_1609);
xnor U1812 (N_1812,N_1748,N_1745);
and U1813 (N_1813,N_1704,N_1779);
xnor U1814 (N_1814,N_1669,N_1783);
and U1815 (N_1815,N_1738,N_1661);
nor U1816 (N_1816,N_1647,N_1648);
and U1817 (N_1817,N_1723,N_1709);
xor U1818 (N_1818,N_1657,N_1697);
nor U1819 (N_1819,N_1603,N_1781);
or U1820 (N_1820,N_1715,N_1797);
nand U1821 (N_1821,N_1763,N_1734);
and U1822 (N_1822,N_1787,N_1654);
nand U1823 (N_1823,N_1719,N_1721);
or U1824 (N_1824,N_1782,N_1668);
nor U1825 (N_1825,N_1790,N_1614);
and U1826 (N_1826,N_1651,N_1616);
nor U1827 (N_1827,N_1610,N_1761);
nor U1828 (N_1828,N_1605,N_1703);
and U1829 (N_1829,N_1730,N_1753);
and U1830 (N_1830,N_1683,N_1618);
nand U1831 (N_1831,N_1684,N_1688);
nor U1832 (N_1832,N_1646,N_1634);
nand U1833 (N_1833,N_1746,N_1791);
nor U1834 (N_1834,N_1695,N_1762);
nor U1835 (N_1835,N_1677,N_1707);
nor U1836 (N_1836,N_1621,N_1720);
nand U1837 (N_1837,N_1617,N_1726);
or U1838 (N_1838,N_1642,N_1606);
and U1839 (N_1839,N_1757,N_1649);
or U1840 (N_1840,N_1752,N_1686);
or U1841 (N_1841,N_1626,N_1679);
nand U1842 (N_1842,N_1771,N_1724);
or U1843 (N_1843,N_1629,N_1628);
and U1844 (N_1844,N_1728,N_1612);
or U1845 (N_1845,N_1635,N_1625);
nand U1846 (N_1846,N_1700,N_1630);
nor U1847 (N_1847,N_1690,N_1794);
or U1848 (N_1848,N_1799,N_1764);
nand U1849 (N_1849,N_1639,N_1792);
and U1850 (N_1850,N_1682,N_1653);
or U1851 (N_1851,N_1636,N_1710);
nand U1852 (N_1852,N_1772,N_1750);
or U1853 (N_1853,N_1643,N_1613);
and U1854 (N_1854,N_1698,N_1667);
xnor U1855 (N_1855,N_1600,N_1604);
and U1856 (N_1856,N_1623,N_1760);
and U1857 (N_1857,N_1638,N_1685);
nand U1858 (N_1858,N_1693,N_1733);
and U1859 (N_1859,N_1602,N_1687);
or U1860 (N_1860,N_1691,N_1756);
or U1861 (N_1861,N_1735,N_1749);
nand U1862 (N_1862,N_1644,N_1718);
xnor U1863 (N_1863,N_1722,N_1640);
nor U1864 (N_1864,N_1742,N_1743);
nor U1865 (N_1865,N_1770,N_1717);
and U1866 (N_1866,N_1633,N_1776);
nand U1867 (N_1867,N_1607,N_1705);
nand U1868 (N_1868,N_1786,N_1675);
nor U1869 (N_1869,N_1740,N_1780);
nor U1870 (N_1870,N_1673,N_1601);
and U1871 (N_1871,N_1681,N_1795);
xnor U1872 (N_1872,N_1775,N_1706);
or U1873 (N_1873,N_1708,N_1663);
or U1874 (N_1874,N_1774,N_1777);
nor U1875 (N_1875,N_1731,N_1714);
and U1876 (N_1876,N_1736,N_1631);
nand U1877 (N_1877,N_1650,N_1678);
nor U1878 (N_1878,N_1694,N_1676);
nor U1879 (N_1879,N_1744,N_1701);
or U1880 (N_1880,N_1716,N_1732);
and U1881 (N_1881,N_1658,N_1692);
or U1882 (N_1882,N_1680,N_1665);
and U1883 (N_1883,N_1727,N_1712);
and U1884 (N_1884,N_1611,N_1796);
or U1885 (N_1885,N_1672,N_1769);
nand U1886 (N_1886,N_1793,N_1778);
nand U1887 (N_1887,N_1759,N_1758);
nor U1888 (N_1888,N_1702,N_1627);
or U1889 (N_1889,N_1755,N_1641);
nand U1890 (N_1890,N_1741,N_1645);
or U1891 (N_1891,N_1666,N_1664);
or U1892 (N_1892,N_1659,N_1655);
and U1893 (N_1893,N_1768,N_1689);
or U1894 (N_1894,N_1751,N_1711);
nor U1895 (N_1895,N_1620,N_1788);
nor U1896 (N_1896,N_1765,N_1785);
nor U1897 (N_1897,N_1624,N_1656);
and U1898 (N_1898,N_1660,N_1729);
xor U1899 (N_1899,N_1652,N_1747);
or U1900 (N_1900,N_1613,N_1672);
nor U1901 (N_1901,N_1619,N_1664);
and U1902 (N_1902,N_1603,N_1710);
nor U1903 (N_1903,N_1609,N_1788);
nand U1904 (N_1904,N_1633,N_1609);
nor U1905 (N_1905,N_1799,N_1686);
or U1906 (N_1906,N_1754,N_1696);
or U1907 (N_1907,N_1775,N_1793);
nand U1908 (N_1908,N_1756,N_1609);
nor U1909 (N_1909,N_1702,N_1643);
nor U1910 (N_1910,N_1609,N_1739);
or U1911 (N_1911,N_1776,N_1725);
nand U1912 (N_1912,N_1688,N_1689);
and U1913 (N_1913,N_1776,N_1639);
nor U1914 (N_1914,N_1618,N_1785);
and U1915 (N_1915,N_1684,N_1672);
nand U1916 (N_1916,N_1661,N_1665);
and U1917 (N_1917,N_1742,N_1784);
or U1918 (N_1918,N_1695,N_1621);
nor U1919 (N_1919,N_1670,N_1732);
nor U1920 (N_1920,N_1726,N_1626);
xor U1921 (N_1921,N_1641,N_1745);
nand U1922 (N_1922,N_1726,N_1650);
nand U1923 (N_1923,N_1651,N_1683);
nand U1924 (N_1924,N_1683,N_1789);
nand U1925 (N_1925,N_1692,N_1605);
nor U1926 (N_1926,N_1794,N_1798);
and U1927 (N_1927,N_1610,N_1743);
and U1928 (N_1928,N_1789,N_1613);
or U1929 (N_1929,N_1714,N_1674);
nand U1930 (N_1930,N_1626,N_1611);
nor U1931 (N_1931,N_1636,N_1613);
or U1932 (N_1932,N_1693,N_1600);
nor U1933 (N_1933,N_1742,N_1702);
and U1934 (N_1934,N_1622,N_1708);
nand U1935 (N_1935,N_1642,N_1672);
nor U1936 (N_1936,N_1679,N_1611);
and U1937 (N_1937,N_1785,N_1743);
or U1938 (N_1938,N_1673,N_1645);
or U1939 (N_1939,N_1676,N_1657);
nand U1940 (N_1940,N_1618,N_1716);
or U1941 (N_1941,N_1697,N_1622);
nor U1942 (N_1942,N_1629,N_1620);
nor U1943 (N_1943,N_1739,N_1632);
nor U1944 (N_1944,N_1737,N_1772);
or U1945 (N_1945,N_1663,N_1680);
nor U1946 (N_1946,N_1633,N_1751);
nor U1947 (N_1947,N_1749,N_1700);
and U1948 (N_1948,N_1649,N_1666);
nand U1949 (N_1949,N_1753,N_1720);
nor U1950 (N_1950,N_1757,N_1681);
nor U1951 (N_1951,N_1601,N_1631);
or U1952 (N_1952,N_1757,N_1720);
and U1953 (N_1953,N_1675,N_1757);
or U1954 (N_1954,N_1752,N_1693);
and U1955 (N_1955,N_1641,N_1771);
or U1956 (N_1956,N_1627,N_1741);
nand U1957 (N_1957,N_1640,N_1788);
nand U1958 (N_1958,N_1728,N_1602);
or U1959 (N_1959,N_1784,N_1756);
and U1960 (N_1960,N_1735,N_1715);
and U1961 (N_1961,N_1691,N_1787);
and U1962 (N_1962,N_1711,N_1677);
nor U1963 (N_1963,N_1732,N_1672);
nand U1964 (N_1964,N_1604,N_1786);
and U1965 (N_1965,N_1606,N_1640);
nor U1966 (N_1966,N_1623,N_1734);
and U1967 (N_1967,N_1615,N_1783);
nor U1968 (N_1968,N_1699,N_1786);
xnor U1969 (N_1969,N_1612,N_1711);
and U1970 (N_1970,N_1619,N_1742);
nor U1971 (N_1971,N_1769,N_1737);
or U1972 (N_1972,N_1722,N_1780);
nor U1973 (N_1973,N_1633,N_1793);
nand U1974 (N_1974,N_1793,N_1784);
or U1975 (N_1975,N_1729,N_1741);
and U1976 (N_1976,N_1605,N_1728);
xnor U1977 (N_1977,N_1749,N_1654);
and U1978 (N_1978,N_1670,N_1791);
and U1979 (N_1979,N_1682,N_1685);
nor U1980 (N_1980,N_1768,N_1610);
or U1981 (N_1981,N_1720,N_1611);
nand U1982 (N_1982,N_1789,N_1773);
nand U1983 (N_1983,N_1668,N_1622);
or U1984 (N_1984,N_1616,N_1786);
nor U1985 (N_1985,N_1634,N_1665);
and U1986 (N_1986,N_1751,N_1674);
xor U1987 (N_1987,N_1785,N_1761);
and U1988 (N_1988,N_1781,N_1720);
nand U1989 (N_1989,N_1798,N_1758);
nor U1990 (N_1990,N_1767,N_1704);
nor U1991 (N_1991,N_1786,N_1609);
nand U1992 (N_1992,N_1780,N_1648);
or U1993 (N_1993,N_1725,N_1706);
nand U1994 (N_1994,N_1741,N_1646);
and U1995 (N_1995,N_1751,N_1612);
nand U1996 (N_1996,N_1763,N_1608);
or U1997 (N_1997,N_1612,N_1688);
or U1998 (N_1998,N_1682,N_1708);
nand U1999 (N_1999,N_1691,N_1631);
nor U2000 (N_2000,N_1806,N_1903);
nand U2001 (N_2001,N_1846,N_1937);
nor U2002 (N_2002,N_1867,N_1948);
xor U2003 (N_2003,N_1821,N_1823);
nand U2004 (N_2004,N_1935,N_1832);
or U2005 (N_2005,N_1887,N_1839);
and U2006 (N_2006,N_1920,N_1801);
nand U2007 (N_2007,N_1904,N_1871);
or U2008 (N_2008,N_1908,N_1844);
nor U2009 (N_2009,N_1959,N_1919);
nor U2010 (N_2010,N_1983,N_1838);
and U2011 (N_2011,N_1944,N_1829);
and U2012 (N_2012,N_1893,N_1899);
nand U2013 (N_2013,N_1863,N_1927);
nor U2014 (N_2014,N_1909,N_1986);
or U2015 (N_2015,N_1860,N_1825);
nor U2016 (N_2016,N_1856,N_1964);
or U2017 (N_2017,N_1884,N_1984);
or U2018 (N_2018,N_1818,N_1954);
nor U2019 (N_2019,N_1942,N_1892);
nor U2020 (N_2020,N_1872,N_1814);
nand U2021 (N_2021,N_1947,N_1805);
nand U2022 (N_2022,N_1896,N_1941);
or U2023 (N_2023,N_1866,N_1882);
or U2024 (N_2024,N_1848,N_1924);
or U2025 (N_2025,N_1962,N_1878);
nand U2026 (N_2026,N_1979,N_1841);
nor U2027 (N_2027,N_1881,N_1971);
nor U2028 (N_2028,N_1906,N_1833);
and U2029 (N_2029,N_1850,N_1934);
or U2030 (N_2030,N_1836,N_1880);
nor U2031 (N_2031,N_1890,N_1802);
nand U2032 (N_2032,N_1912,N_1928);
and U2033 (N_2033,N_1968,N_1803);
or U2034 (N_2034,N_1943,N_1950);
nor U2035 (N_2035,N_1857,N_1945);
nand U2036 (N_2036,N_1988,N_1898);
and U2037 (N_2037,N_1868,N_1967);
nand U2038 (N_2038,N_1949,N_1834);
nand U2039 (N_2039,N_1917,N_1812);
nand U2040 (N_2040,N_1862,N_1966);
xnor U2041 (N_2041,N_1996,N_1901);
or U2042 (N_2042,N_1972,N_1817);
or U2043 (N_2043,N_1933,N_1930);
xor U2044 (N_2044,N_1990,N_1888);
and U2045 (N_2045,N_1830,N_1816);
nor U2046 (N_2046,N_1873,N_1815);
nor U2047 (N_2047,N_1865,N_1940);
and U2048 (N_2048,N_1932,N_1993);
or U2049 (N_2049,N_1910,N_1975);
nor U2050 (N_2050,N_1902,N_1831);
nor U2051 (N_2051,N_1999,N_1938);
nand U2052 (N_2052,N_1822,N_1922);
or U2053 (N_2053,N_1809,N_1891);
nand U2054 (N_2054,N_1936,N_1987);
xor U2055 (N_2055,N_1824,N_1911);
or U2056 (N_2056,N_1808,N_1913);
nor U2057 (N_2057,N_1982,N_1907);
and U2058 (N_2058,N_1965,N_1960);
xnor U2059 (N_2059,N_1842,N_1875);
or U2060 (N_2060,N_1951,N_1870);
nor U2061 (N_2061,N_1998,N_1952);
nor U2062 (N_2062,N_1918,N_1883);
nand U2063 (N_2063,N_1991,N_1837);
or U2064 (N_2064,N_1953,N_1864);
or U2065 (N_2065,N_1970,N_1992);
or U2066 (N_2066,N_1939,N_1874);
or U2067 (N_2067,N_1956,N_1851);
nand U2068 (N_2068,N_1859,N_1820);
or U2069 (N_2069,N_1855,N_1914);
and U2070 (N_2070,N_1895,N_1826);
nand U2071 (N_2071,N_1957,N_1819);
nand U2072 (N_2072,N_1858,N_1969);
or U2073 (N_2073,N_1807,N_1900);
nor U2074 (N_2074,N_1977,N_1886);
nand U2075 (N_2075,N_1925,N_1827);
or U2076 (N_2076,N_1915,N_1879);
nor U2077 (N_2077,N_1813,N_1843);
and U2078 (N_2078,N_1978,N_1997);
or U2079 (N_2079,N_1853,N_1955);
or U2080 (N_2080,N_1985,N_1994);
and U2081 (N_2081,N_1961,N_1921);
or U2082 (N_2082,N_1800,N_1811);
nand U2083 (N_2083,N_1981,N_1926);
or U2084 (N_2084,N_1854,N_1889);
nor U2085 (N_2085,N_1973,N_1958);
or U2086 (N_2086,N_1946,N_1894);
or U2087 (N_2087,N_1852,N_1995);
nand U2088 (N_2088,N_1897,N_1931);
nor U2089 (N_2089,N_1849,N_1989);
nor U2090 (N_2090,N_1804,N_1876);
nor U2091 (N_2091,N_1916,N_1828);
or U2092 (N_2092,N_1929,N_1923);
and U2093 (N_2093,N_1877,N_1810);
or U2094 (N_2094,N_1905,N_1835);
nor U2095 (N_2095,N_1963,N_1974);
xnor U2096 (N_2096,N_1840,N_1869);
nor U2097 (N_2097,N_1976,N_1845);
nand U2098 (N_2098,N_1885,N_1847);
nand U2099 (N_2099,N_1980,N_1861);
nand U2100 (N_2100,N_1958,N_1863);
or U2101 (N_2101,N_1908,N_1953);
nor U2102 (N_2102,N_1920,N_1966);
or U2103 (N_2103,N_1898,N_1897);
nand U2104 (N_2104,N_1803,N_1919);
and U2105 (N_2105,N_1928,N_1803);
and U2106 (N_2106,N_1807,N_1947);
and U2107 (N_2107,N_1832,N_1838);
or U2108 (N_2108,N_1899,N_1939);
nand U2109 (N_2109,N_1811,N_1951);
and U2110 (N_2110,N_1851,N_1888);
nand U2111 (N_2111,N_1909,N_1833);
or U2112 (N_2112,N_1848,N_1946);
nor U2113 (N_2113,N_1994,N_1900);
nand U2114 (N_2114,N_1967,N_1802);
and U2115 (N_2115,N_1952,N_1823);
and U2116 (N_2116,N_1985,N_1895);
or U2117 (N_2117,N_1978,N_1850);
and U2118 (N_2118,N_1818,N_1920);
and U2119 (N_2119,N_1925,N_1886);
and U2120 (N_2120,N_1821,N_1819);
and U2121 (N_2121,N_1809,N_1917);
or U2122 (N_2122,N_1914,N_1987);
and U2123 (N_2123,N_1852,N_1927);
nor U2124 (N_2124,N_1865,N_1855);
nor U2125 (N_2125,N_1984,N_1922);
xor U2126 (N_2126,N_1918,N_1825);
nand U2127 (N_2127,N_1913,N_1897);
nand U2128 (N_2128,N_1842,N_1936);
and U2129 (N_2129,N_1829,N_1995);
or U2130 (N_2130,N_1916,N_1969);
and U2131 (N_2131,N_1964,N_1880);
or U2132 (N_2132,N_1895,N_1842);
nor U2133 (N_2133,N_1952,N_1872);
nor U2134 (N_2134,N_1865,N_1803);
or U2135 (N_2135,N_1825,N_1958);
nand U2136 (N_2136,N_1886,N_1814);
or U2137 (N_2137,N_1890,N_1875);
nor U2138 (N_2138,N_1905,N_1903);
nor U2139 (N_2139,N_1863,N_1815);
nand U2140 (N_2140,N_1952,N_1942);
and U2141 (N_2141,N_1819,N_1841);
or U2142 (N_2142,N_1985,N_1820);
and U2143 (N_2143,N_1967,N_1935);
and U2144 (N_2144,N_1978,N_1827);
nand U2145 (N_2145,N_1839,N_1994);
nand U2146 (N_2146,N_1943,N_1932);
nand U2147 (N_2147,N_1973,N_1908);
and U2148 (N_2148,N_1924,N_1907);
nor U2149 (N_2149,N_1812,N_1868);
or U2150 (N_2150,N_1856,N_1897);
nand U2151 (N_2151,N_1881,N_1878);
nand U2152 (N_2152,N_1984,N_1874);
nor U2153 (N_2153,N_1820,N_1969);
or U2154 (N_2154,N_1811,N_1819);
nor U2155 (N_2155,N_1978,N_1938);
nor U2156 (N_2156,N_1854,N_1880);
nor U2157 (N_2157,N_1971,N_1801);
nand U2158 (N_2158,N_1805,N_1937);
nand U2159 (N_2159,N_1838,N_1833);
nand U2160 (N_2160,N_1915,N_1854);
and U2161 (N_2161,N_1898,N_1849);
nand U2162 (N_2162,N_1886,N_1937);
or U2163 (N_2163,N_1996,N_1848);
and U2164 (N_2164,N_1912,N_1983);
or U2165 (N_2165,N_1831,N_1910);
nor U2166 (N_2166,N_1976,N_1980);
nand U2167 (N_2167,N_1929,N_1800);
or U2168 (N_2168,N_1827,N_1814);
or U2169 (N_2169,N_1831,N_1898);
nand U2170 (N_2170,N_1800,N_1829);
nor U2171 (N_2171,N_1840,N_1958);
nand U2172 (N_2172,N_1838,N_1879);
nor U2173 (N_2173,N_1824,N_1913);
nand U2174 (N_2174,N_1844,N_1994);
and U2175 (N_2175,N_1993,N_1926);
or U2176 (N_2176,N_1813,N_1920);
or U2177 (N_2177,N_1918,N_1878);
and U2178 (N_2178,N_1985,N_1802);
and U2179 (N_2179,N_1884,N_1843);
nand U2180 (N_2180,N_1851,N_1998);
nor U2181 (N_2181,N_1956,N_1843);
nand U2182 (N_2182,N_1998,N_1843);
or U2183 (N_2183,N_1846,N_1874);
xnor U2184 (N_2184,N_1869,N_1924);
nand U2185 (N_2185,N_1899,N_1873);
and U2186 (N_2186,N_1999,N_1966);
nand U2187 (N_2187,N_1920,N_1906);
nor U2188 (N_2188,N_1960,N_1920);
xor U2189 (N_2189,N_1870,N_1973);
or U2190 (N_2190,N_1870,N_1900);
and U2191 (N_2191,N_1922,N_1973);
or U2192 (N_2192,N_1826,N_1921);
nand U2193 (N_2193,N_1907,N_1888);
nor U2194 (N_2194,N_1907,N_1908);
and U2195 (N_2195,N_1953,N_1911);
nor U2196 (N_2196,N_1999,N_1862);
and U2197 (N_2197,N_1876,N_1987);
or U2198 (N_2198,N_1961,N_1937);
and U2199 (N_2199,N_1989,N_1862);
or U2200 (N_2200,N_2025,N_2167);
nor U2201 (N_2201,N_2075,N_2145);
nor U2202 (N_2202,N_2160,N_2034);
nor U2203 (N_2203,N_2115,N_2000);
and U2204 (N_2204,N_2006,N_2012);
nand U2205 (N_2205,N_2141,N_2114);
and U2206 (N_2206,N_2125,N_2051);
and U2207 (N_2207,N_2013,N_2149);
and U2208 (N_2208,N_2066,N_2181);
or U2209 (N_2209,N_2178,N_2162);
nor U2210 (N_2210,N_2107,N_2113);
and U2211 (N_2211,N_2117,N_2148);
or U2212 (N_2212,N_2039,N_2171);
nor U2213 (N_2213,N_2062,N_2129);
or U2214 (N_2214,N_2147,N_2169);
nand U2215 (N_2215,N_2187,N_2031);
nor U2216 (N_2216,N_2104,N_2170);
or U2217 (N_2217,N_2055,N_2180);
nand U2218 (N_2218,N_2046,N_2021);
nor U2219 (N_2219,N_2077,N_2019);
nor U2220 (N_2220,N_2023,N_2166);
or U2221 (N_2221,N_2049,N_2068);
nor U2222 (N_2222,N_2111,N_2057);
and U2223 (N_2223,N_2079,N_2142);
or U2224 (N_2224,N_2179,N_2128);
nor U2225 (N_2225,N_2159,N_2199);
or U2226 (N_2226,N_2008,N_2082);
nor U2227 (N_2227,N_2018,N_2030);
nand U2228 (N_2228,N_2097,N_2016);
nand U2229 (N_2229,N_2014,N_2092);
nand U2230 (N_2230,N_2106,N_2120);
or U2231 (N_2231,N_2132,N_2157);
nand U2232 (N_2232,N_2146,N_2080);
or U2233 (N_2233,N_2083,N_2088);
nor U2234 (N_2234,N_2011,N_2053);
nor U2235 (N_2235,N_2151,N_2101);
nand U2236 (N_2236,N_2121,N_2193);
and U2237 (N_2237,N_2076,N_2067);
nor U2238 (N_2238,N_2081,N_2110);
and U2239 (N_2239,N_2005,N_2070);
xnor U2240 (N_2240,N_2186,N_2029);
and U2241 (N_2241,N_2112,N_2060);
nand U2242 (N_2242,N_2143,N_2084);
or U2243 (N_2243,N_2048,N_2040);
or U2244 (N_2244,N_2096,N_2135);
or U2245 (N_2245,N_2189,N_2036);
nor U2246 (N_2246,N_2172,N_2054);
and U2247 (N_2247,N_2109,N_2131);
nand U2248 (N_2248,N_2024,N_2022);
nor U2249 (N_2249,N_2196,N_2122);
or U2250 (N_2250,N_2150,N_2140);
nand U2251 (N_2251,N_2123,N_2116);
or U2252 (N_2252,N_2017,N_2126);
nand U2253 (N_2253,N_2105,N_2183);
or U2254 (N_2254,N_2056,N_2165);
or U2255 (N_2255,N_2042,N_2063);
and U2256 (N_2256,N_2194,N_2087);
or U2257 (N_2257,N_2156,N_2064);
or U2258 (N_2258,N_2119,N_2007);
and U2259 (N_2259,N_2099,N_2168);
xnor U2260 (N_2260,N_2103,N_2093);
or U2261 (N_2261,N_2153,N_2020);
and U2262 (N_2262,N_2137,N_2139);
nor U2263 (N_2263,N_2094,N_2033);
or U2264 (N_2264,N_2004,N_2163);
nand U2265 (N_2265,N_2136,N_2001);
and U2266 (N_2266,N_2061,N_2124);
or U2267 (N_2267,N_2118,N_2144);
nor U2268 (N_2268,N_2102,N_2032);
xnor U2269 (N_2269,N_2047,N_2191);
and U2270 (N_2270,N_2050,N_2002);
and U2271 (N_2271,N_2072,N_2195);
or U2272 (N_2272,N_2100,N_2134);
or U2273 (N_2273,N_2065,N_2044);
or U2274 (N_2274,N_2027,N_2108);
nand U2275 (N_2275,N_2197,N_2089);
xor U2276 (N_2276,N_2161,N_2130);
or U2277 (N_2277,N_2133,N_2177);
or U2278 (N_2278,N_2154,N_2015);
and U2279 (N_2279,N_2090,N_2164);
nor U2280 (N_2280,N_2173,N_2184);
and U2281 (N_2281,N_2028,N_2127);
and U2282 (N_2282,N_2185,N_2071);
nor U2283 (N_2283,N_2188,N_2069);
and U2284 (N_2284,N_2035,N_2138);
and U2285 (N_2285,N_2192,N_2045);
and U2286 (N_2286,N_2058,N_2038);
nand U2287 (N_2287,N_2198,N_2052);
nor U2288 (N_2288,N_2182,N_2091);
and U2289 (N_2289,N_2174,N_2074);
and U2290 (N_2290,N_2086,N_2152);
nor U2291 (N_2291,N_2190,N_2010);
nor U2292 (N_2292,N_2158,N_2085);
or U2293 (N_2293,N_2041,N_2043);
nand U2294 (N_2294,N_2078,N_2003);
nand U2295 (N_2295,N_2176,N_2009);
or U2296 (N_2296,N_2098,N_2175);
and U2297 (N_2297,N_2026,N_2059);
and U2298 (N_2298,N_2037,N_2155);
and U2299 (N_2299,N_2095,N_2073);
nor U2300 (N_2300,N_2147,N_2030);
or U2301 (N_2301,N_2138,N_2102);
and U2302 (N_2302,N_2000,N_2054);
nand U2303 (N_2303,N_2176,N_2059);
nor U2304 (N_2304,N_2153,N_2031);
nand U2305 (N_2305,N_2149,N_2048);
or U2306 (N_2306,N_2194,N_2157);
or U2307 (N_2307,N_2133,N_2008);
nor U2308 (N_2308,N_2095,N_2196);
or U2309 (N_2309,N_2109,N_2108);
nor U2310 (N_2310,N_2181,N_2033);
nand U2311 (N_2311,N_2056,N_2135);
nand U2312 (N_2312,N_2121,N_2153);
and U2313 (N_2313,N_2066,N_2043);
nor U2314 (N_2314,N_2126,N_2107);
nor U2315 (N_2315,N_2065,N_2174);
nor U2316 (N_2316,N_2110,N_2140);
or U2317 (N_2317,N_2097,N_2199);
or U2318 (N_2318,N_2078,N_2096);
nand U2319 (N_2319,N_2050,N_2001);
or U2320 (N_2320,N_2170,N_2052);
nand U2321 (N_2321,N_2097,N_2141);
nor U2322 (N_2322,N_2058,N_2055);
or U2323 (N_2323,N_2059,N_2143);
and U2324 (N_2324,N_2142,N_2164);
and U2325 (N_2325,N_2088,N_2095);
or U2326 (N_2326,N_2193,N_2040);
nand U2327 (N_2327,N_2097,N_2126);
and U2328 (N_2328,N_2199,N_2031);
nor U2329 (N_2329,N_2027,N_2034);
nor U2330 (N_2330,N_2132,N_2146);
nand U2331 (N_2331,N_2011,N_2197);
or U2332 (N_2332,N_2121,N_2016);
nand U2333 (N_2333,N_2191,N_2071);
and U2334 (N_2334,N_2031,N_2198);
nor U2335 (N_2335,N_2168,N_2106);
nor U2336 (N_2336,N_2014,N_2097);
and U2337 (N_2337,N_2067,N_2044);
and U2338 (N_2338,N_2173,N_2032);
or U2339 (N_2339,N_2109,N_2119);
or U2340 (N_2340,N_2137,N_2004);
nand U2341 (N_2341,N_2103,N_2153);
and U2342 (N_2342,N_2148,N_2021);
or U2343 (N_2343,N_2022,N_2078);
xnor U2344 (N_2344,N_2062,N_2029);
xor U2345 (N_2345,N_2160,N_2148);
nand U2346 (N_2346,N_2128,N_2199);
nor U2347 (N_2347,N_2148,N_2095);
and U2348 (N_2348,N_2006,N_2162);
and U2349 (N_2349,N_2118,N_2081);
or U2350 (N_2350,N_2091,N_2068);
nand U2351 (N_2351,N_2104,N_2013);
and U2352 (N_2352,N_2160,N_2017);
nand U2353 (N_2353,N_2023,N_2055);
and U2354 (N_2354,N_2099,N_2151);
nand U2355 (N_2355,N_2188,N_2130);
and U2356 (N_2356,N_2132,N_2052);
and U2357 (N_2357,N_2049,N_2007);
or U2358 (N_2358,N_2176,N_2154);
or U2359 (N_2359,N_2165,N_2199);
or U2360 (N_2360,N_2060,N_2039);
nand U2361 (N_2361,N_2176,N_2036);
nor U2362 (N_2362,N_2127,N_2009);
and U2363 (N_2363,N_2115,N_2061);
nand U2364 (N_2364,N_2001,N_2165);
and U2365 (N_2365,N_2012,N_2103);
nor U2366 (N_2366,N_2009,N_2194);
nor U2367 (N_2367,N_2080,N_2075);
or U2368 (N_2368,N_2112,N_2164);
nand U2369 (N_2369,N_2161,N_2074);
and U2370 (N_2370,N_2033,N_2169);
nand U2371 (N_2371,N_2008,N_2093);
nor U2372 (N_2372,N_2028,N_2042);
nor U2373 (N_2373,N_2165,N_2173);
nor U2374 (N_2374,N_2176,N_2174);
or U2375 (N_2375,N_2028,N_2167);
nand U2376 (N_2376,N_2144,N_2127);
or U2377 (N_2377,N_2122,N_2112);
nand U2378 (N_2378,N_2050,N_2178);
nor U2379 (N_2379,N_2011,N_2128);
nand U2380 (N_2380,N_2141,N_2060);
and U2381 (N_2381,N_2094,N_2130);
or U2382 (N_2382,N_2011,N_2106);
nand U2383 (N_2383,N_2194,N_2183);
or U2384 (N_2384,N_2140,N_2042);
and U2385 (N_2385,N_2036,N_2132);
nand U2386 (N_2386,N_2070,N_2157);
nor U2387 (N_2387,N_2040,N_2116);
nand U2388 (N_2388,N_2001,N_2115);
or U2389 (N_2389,N_2026,N_2057);
nor U2390 (N_2390,N_2148,N_2059);
nor U2391 (N_2391,N_2015,N_2003);
nand U2392 (N_2392,N_2041,N_2089);
or U2393 (N_2393,N_2109,N_2181);
nand U2394 (N_2394,N_2010,N_2029);
nor U2395 (N_2395,N_2184,N_2190);
or U2396 (N_2396,N_2035,N_2199);
or U2397 (N_2397,N_2028,N_2183);
nor U2398 (N_2398,N_2106,N_2179);
nor U2399 (N_2399,N_2007,N_2101);
or U2400 (N_2400,N_2395,N_2351);
nand U2401 (N_2401,N_2271,N_2341);
nand U2402 (N_2402,N_2280,N_2363);
and U2403 (N_2403,N_2301,N_2339);
nor U2404 (N_2404,N_2379,N_2333);
and U2405 (N_2405,N_2359,N_2305);
and U2406 (N_2406,N_2371,N_2294);
and U2407 (N_2407,N_2335,N_2377);
and U2408 (N_2408,N_2259,N_2376);
nand U2409 (N_2409,N_2212,N_2211);
and U2410 (N_2410,N_2257,N_2355);
or U2411 (N_2411,N_2242,N_2399);
nand U2412 (N_2412,N_2261,N_2295);
nand U2413 (N_2413,N_2243,N_2283);
nand U2414 (N_2414,N_2297,N_2336);
and U2415 (N_2415,N_2380,N_2249);
or U2416 (N_2416,N_2235,N_2375);
nand U2417 (N_2417,N_2238,N_2344);
or U2418 (N_2418,N_2269,N_2389);
or U2419 (N_2419,N_2313,N_2292);
nand U2420 (N_2420,N_2362,N_2205);
xnor U2421 (N_2421,N_2265,N_2390);
nand U2422 (N_2422,N_2207,N_2391);
nand U2423 (N_2423,N_2353,N_2231);
and U2424 (N_2424,N_2378,N_2307);
nand U2425 (N_2425,N_2366,N_2346);
nand U2426 (N_2426,N_2310,N_2356);
xor U2427 (N_2427,N_2274,N_2219);
nand U2428 (N_2428,N_2228,N_2288);
nand U2429 (N_2429,N_2327,N_2369);
or U2430 (N_2430,N_2203,N_2309);
nor U2431 (N_2431,N_2251,N_2202);
or U2432 (N_2432,N_2276,N_2392);
nor U2433 (N_2433,N_2232,N_2230);
nand U2434 (N_2434,N_2221,N_2284);
or U2435 (N_2435,N_2299,N_2239);
nor U2436 (N_2436,N_2210,N_2298);
or U2437 (N_2437,N_2314,N_2322);
nor U2438 (N_2438,N_2350,N_2222);
nand U2439 (N_2439,N_2384,N_2291);
and U2440 (N_2440,N_2244,N_2328);
or U2441 (N_2441,N_2370,N_2319);
or U2442 (N_2442,N_2394,N_2357);
nand U2443 (N_2443,N_2208,N_2387);
or U2444 (N_2444,N_2343,N_2381);
and U2445 (N_2445,N_2247,N_2348);
xnor U2446 (N_2446,N_2223,N_2303);
nand U2447 (N_2447,N_2216,N_2386);
nor U2448 (N_2448,N_2285,N_2396);
nand U2449 (N_2449,N_2293,N_2260);
nand U2450 (N_2450,N_2287,N_2226);
or U2451 (N_2451,N_2360,N_2334);
nand U2452 (N_2452,N_2349,N_2254);
or U2453 (N_2453,N_2241,N_2318);
nor U2454 (N_2454,N_2236,N_2325);
and U2455 (N_2455,N_2258,N_2218);
and U2456 (N_2456,N_2250,N_2372);
nor U2457 (N_2457,N_2281,N_2255);
and U2458 (N_2458,N_2213,N_2367);
or U2459 (N_2459,N_2321,N_2234);
nand U2460 (N_2460,N_2383,N_2365);
nand U2461 (N_2461,N_2275,N_2253);
and U2462 (N_2462,N_2224,N_2340);
and U2463 (N_2463,N_2245,N_2374);
or U2464 (N_2464,N_2308,N_2272);
xor U2465 (N_2465,N_2278,N_2316);
nor U2466 (N_2466,N_2315,N_2296);
or U2467 (N_2467,N_2329,N_2342);
or U2468 (N_2468,N_2277,N_2323);
and U2469 (N_2469,N_2302,N_2273);
nand U2470 (N_2470,N_2206,N_2338);
or U2471 (N_2471,N_2364,N_2358);
nand U2472 (N_2472,N_2252,N_2267);
and U2473 (N_2473,N_2268,N_2289);
and U2474 (N_2474,N_2217,N_2270);
nor U2475 (N_2475,N_2320,N_2337);
xor U2476 (N_2476,N_2347,N_2200);
and U2477 (N_2477,N_2304,N_2240);
nor U2478 (N_2478,N_2306,N_2330);
or U2479 (N_2479,N_2282,N_2332);
and U2480 (N_2480,N_2388,N_2246);
nand U2481 (N_2481,N_2215,N_2227);
nand U2482 (N_2482,N_2324,N_2266);
nor U2483 (N_2483,N_2352,N_2311);
nand U2484 (N_2484,N_2279,N_2256);
nor U2485 (N_2485,N_2361,N_2317);
nor U2486 (N_2486,N_2373,N_2385);
or U2487 (N_2487,N_2326,N_2398);
nand U2488 (N_2488,N_2262,N_2368);
nor U2489 (N_2489,N_2204,N_2220);
nand U2490 (N_2490,N_2331,N_2237);
or U2491 (N_2491,N_2393,N_2201);
or U2492 (N_2492,N_2248,N_2263);
or U2493 (N_2493,N_2354,N_2300);
nor U2494 (N_2494,N_2286,N_2264);
nand U2495 (N_2495,N_2382,N_2209);
nand U2496 (N_2496,N_2225,N_2233);
and U2497 (N_2497,N_2229,N_2214);
or U2498 (N_2498,N_2397,N_2312);
nand U2499 (N_2499,N_2290,N_2345);
nor U2500 (N_2500,N_2279,N_2272);
and U2501 (N_2501,N_2274,N_2289);
nor U2502 (N_2502,N_2253,N_2374);
xnor U2503 (N_2503,N_2320,N_2350);
nor U2504 (N_2504,N_2265,N_2343);
nand U2505 (N_2505,N_2391,N_2216);
and U2506 (N_2506,N_2236,N_2254);
nand U2507 (N_2507,N_2348,N_2362);
nand U2508 (N_2508,N_2361,N_2352);
nor U2509 (N_2509,N_2352,N_2393);
nor U2510 (N_2510,N_2221,N_2211);
nand U2511 (N_2511,N_2246,N_2357);
and U2512 (N_2512,N_2256,N_2232);
xor U2513 (N_2513,N_2376,N_2229);
and U2514 (N_2514,N_2271,N_2303);
or U2515 (N_2515,N_2338,N_2214);
and U2516 (N_2516,N_2281,N_2380);
or U2517 (N_2517,N_2397,N_2206);
nand U2518 (N_2518,N_2230,N_2234);
and U2519 (N_2519,N_2286,N_2293);
nor U2520 (N_2520,N_2259,N_2258);
nand U2521 (N_2521,N_2340,N_2351);
and U2522 (N_2522,N_2371,N_2325);
and U2523 (N_2523,N_2230,N_2362);
nor U2524 (N_2524,N_2228,N_2347);
and U2525 (N_2525,N_2321,N_2203);
or U2526 (N_2526,N_2247,N_2363);
nor U2527 (N_2527,N_2294,N_2380);
and U2528 (N_2528,N_2214,N_2235);
or U2529 (N_2529,N_2323,N_2397);
or U2530 (N_2530,N_2380,N_2312);
nand U2531 (N_2531,N_2371,N_2224);
nor U2532 (N_2532,N_2331,N_2371);
and U2533 (N_2533,N_2295,N_2349);
nor U2534 (N_2534,N_2338,N_2245);
nor U2535 (N_2535,N_2365,N_2227);
nand U2536 (N_2536,N_2248,N_2300);
and U2537 (N_2537,N_2256,N_2245);
nor U2538 (N_2538,N_2249,N_2376);
and U2539 (N_2539,N_2286,N_2239);
or U2540 (N_2540,N_2323,N_2262);
or U2541 (N_2541,N_2391,N_2206);
or U2542 (N_2542,N_2205,N_2252);
nand U2543 (N_2543,N_2274,N_2301);
or U2544 (N_2544,N_2348,N_2384);
nand U2545 (N_2545,N_2211,N_2329);
and U2546 (N_2546,N_2358,N_2235);
nand U2547 (N_2547,N_2244,N_2229);
and U2548 (N_2548,N_2229,N_2374);
or U2549 (N_2549,N_2285,N_2302);
nor U2550 (N_2550,N_2288,N_2330);
nand U2551 (N_2551,N_2372,N_2297);
nor U2552 (N_2552,N_2203,N_2269);
nor U2553 (N_2553,N_2334,N_2309);
nor U2554 (N_2554,N_2246,N_2229);
and U2555 (N_2555,N_2205,N_2243);
nor U2556 (N_2556,N_2252,N_2297);
and U2557 (N_2557,N_2299,N_2272);
nand U2558 (N_2558,N_2398,N_2302);
xnor U2559 (N_2559,N_2229,N_2320);
or U2560 (N_2560,N_2286,N_2276);
or U2561 (N_2561,N_2376,N_2216);
and U2562 (N_2562,N_2396,N_2391);
and U2563 (N_2563,N_2377,N_2395);
nand U2564 (N_2564,N_2389,N_2390);
or U2565 (N_2565,N_2389,N_2316);
and U2566 (N_2566,N_2372,N_2365);
or U2567 (N_2567,N_2227,N_2330);
nor U2568 (N_2568,N_2251,N_2263);
nand U2569 (N_2569,N_2311,N_2236);
nor U2570 (N_2570,N_2221,N_2355);
nor U2571 (N_2571,N_2267,N_2245);
nand U2572 (N_2572,N_2390,N_2220);
and U2573 (N_2573,N_2320,N_2334);
nor U2574 (N_2574,N_2215,N_2264);
nand U2575 (N_2575,N_2344,N_2231);
nor U2576 (N_2576,N_2283,N_2230);
nand U2577 (N_2577,N_2300,N_2290);
and U2578 (N_2578,N_2283,N_2284);
nand U2579 (N_2579,N_2240,N_2361);
and U2580 (N_2580,N_2216,N_2383);
nor U2581 (N_2581,N_2329,N_2233);
nor U2582 (N_2582,N_2317,N_2276);
nor U2583 (N_2583,N_2346,N_2228);
or U2584 (N_2584,N_2375,N_2224);
and U2585 (N_2585,N_2234,N_2292);
and U2586 (N_2586,N_2340,N_2398);
and U2587 (N_2587,N_2215,N_2380);
nor U2588 (N_2588,N_2357,N_2286);
nand U2589 (N_2589,N_2311,N_2230);
and U2590 (N_2590,N_2383,N_2346);
or U2591 (N_2591,N_2261,N_2283);
xor U2592 (N_2592,N_2335,N_2312);
nor U2593 (N_2593,N_2365,N_2266);
or U2594 (N_2594,N_2225,N_2329);
or U2595 (N_2595,N_2360,N_2251);
and U2596 (N_2596,N_2365,N_2213);
nand U2597 (N_2597,N_2393,N_2328);
or U2598 (N_2598,N_2221,N_2318);
nand U2599 (N_2599,N_2382,N_2345);
or U2600 (N_2600,N_2402,N_2448);
nor U2601 (N_2601,N_2449,N_2518);
or U2602 (N_2602,N_2418,N_2435);
nand U2603 (N_2603,N_2598,N_2471);
or U2604 (N_2604,N_2547,N_2454);
and U2605 (N_2605,N_2401,N_2420);
nand U2606 (N_2606,N_2446,N_2429);
nand U2607 (N_2607,N_2512,N_2575);
nor U2608 (N_2608,N_2493,N_2408);
nor U2609 (N_2609,N_2470,N_2593);
nor U2610 (N_2610,N_2467,N_2428);
nand U2611 (N_2611,N_2578,N_2568);
nand U2612 (N_2612,N_2499,N_2464);
and U2613 (N_2613,N_2555,N_2431);
and U2614 (N_2614,N_2447,N_2466);
and U2615 (N_2615,N_2452,N_2495);
or U2616 (N_2616,N_2583,N_2477);
xor U2617 (N_2617,N_2417,N_2425);
and U2618 (N_2618,N_2554,N_2438);
and U2619 (N_2619,N_2460,N_2521);
or U2620 (N_2620,N_2528,N_2421);
or U2621 (N_2621,N_2469,N_2517);
or U2622 (N_2622,N_2462,N_2461);
nand U2623 (N_2623,N_2474,N_2523);
nand U2624 (N_2624,N_2492,N_2529);
nand U2625 (N_2625,N_2441,N_2596);
or U2626 (N_2626,N_2488,N_2584);
or U2627 (N_2627,N_2473,N_2497);
nor U2628 (N_2628,N_2451,N_2487);
nor U2629 (N_2629,N_2409,N_2534);
nor U2630 (N_2630,N_2545,N_2567);
and U2631 (N_2631,N_2522,N_2405);
and U2632 (N_2632,N_2480,N_2573);
nor U2633 (N_2633,N_2513,N_2566);
and U2634 (N_2634,N_2579,N_2450);
nor U2635 (N_2635,N_2414,N_2501);
nand U2636 (N_2636,N_2430,N_2535);
or U2637 (N_2637,N_2542,N_2515);
nand U2638 (N_2638,N_2476,N_2509);
and U2639 (N_2639,N_2538,N_2577);
xnor U2640 (N_2640,N_2455,N_2550);
and U2641 (N_2641,N_2486,N_2597);
nand U2642 (N_2642,N_2591,N_2525);
and U2643 (N_2643,N_2472,N_2416);
nor U2644 (N_2644,N_2475,N_2500);
nand U2645 (N_2645,N_2502,N_2503);
or U2646 (N_2646,N_2558,N_2582);
xor U2647 (N_2647,N_2404,N_2444);
nor U2648 (N_2648,N_2571,N_2531);
nand U2649 (N_2649,N_2433,N_2560);
or U2650 (N_2650,N_2457,N_2490);
xor U2651 (N_2651,N_2561,N_2539);
and U2652 (N_2652,N_2599,N_2595);
nor U2653 (N_2653,N_2533,N_2496);
nand U2654 (N_2654,N_2443,N_2419);
or U2655 (N_2655,N_2413,N_2516);
nand U2656 (N_2656,N_2442,N_2526);
nand U2657 (N_2657,N_2507,N_2543);
and U2658 (N_2658,N_2572,N_2463);
and U2659 (N_2659,N_2432,N_2489);
nor U2660 (N_2660,N_2423,N_2506);
nor U2661 (N_2661,N_2562,N_2415);
and U2662 (N_2662,N_2586,N_2559);
nor U2663 (N_2663,N_2505,N_2569);
xor U2664 (N_2664,N_2594,N_2580);
and U2665 (N_2665,N_2589,N_2479);
nand U2666 (N_2666,N_2403,N_2422);
or U2667 (N_2667,N_2494,N_2574);
nor U2668 (N_2668,N_2514,N_2581);
and U2669 (N_2669,N_2536,N_2453);
nand U2670 (N_2670,N_2465,N_2427);
nor U2671 (N_2671,N_2590,N_2524);
nor U2672 (N_2672,N_2548,N_2437);
nand U2673 (N_2673,N_2556,N_2410);
nand U2674 (N_2674,N_2532,N_2519);
nand U2675 (N_2675,N_2468,N_2540);
nor U2676 (N_2676,N_2483,N_2587);
nor U2677 (N_2677,N_2412,N_2439);
nand U2678 (N_2678,N_2553,N_2588);
or U2679 (N_2679,N_2498,N_2434);
nand U2680 (N_2680,N_2481,N_2440);
or U2681 (N_2681,N_2510,N_2557);
nand U2682 (N_2682,N_2458,N_2576);
nand U2683 (N_2683,N_2406,N_2478);
nand U2684 (N_2684,N_2407,N_2445);
nand U2685 (N_2685,N_2459,N_2563);
or U2686 (N_2686,N_2541,N_2546);
or U2687 (N_2687,N_2411,N_2436);
or U2688 (N_2688,N_2564,N_2504);
nand U2689 (N_2689,N_2585,N_2549);
nand U2690 (N_2690,N_2511,N_2530);
and U2691 (N_2691,N_2544,N_2552);
nor U2692 (N_2692,N_2570,N_2400);
nor U2693 (N_2693,N_2482,N_2565);
nor U2694 (N_2694,N_2551,N_2426);
or U2695 (N_2695,N_2456,N_2491);
nor U2696 (N_2696,N_2592,N_2520);
nor U2697 (N_2697,N_2537,N_2485);
nor U2698 (N_2698,N_2527,N_2508);
nor U2699 (N_2699,N_2424,N_2484);
nor U2700 (N_2700,N_2485,N_2461);
nand U2701 (N_2701,N_2439,N_2542);
nand U2702 (N_2702,N_2420,N_2574);
and U2703 (N_2703,N_2583,N_2520);
and U2704 (N_2704,N_2527,N_2524);
nand U2705 (N_2705,N_2426,N_2545);
or U2706 (N_2706,N_2585,N_2542);
nor U2707 (N_2707,N_2444,N_2439);
or U2708 (N_2708,N_2444,N_2592);
and U2709 (N_2709,N_2476,N_2559);
and U2710 (N_2710,N_2474,N_2491);
and U2711 (N_2711,N_2567,N_2522);
and U2712 (N_2712,N_2519,N_2514);
nor U2713 (N_2713,N_2432,N_2540);
or U2714 (N_2714,N_2466,N_2589);
and U2715 (N_2715,N_2544,N_2557);
nor U2716 (N_2716,N_2429,N_2557);
and U2717 (N_2717,N_2566,N_2414);
nor U2718 (N_2718,N_2500,N_2487);
or U2719 (N_2719,N_2498,N_2501);
nor U2720 (N_2720,N_2541,N_2523);
or U2721 (N_2721,N_2459,N_2481);
nand U2722 (N_2722,N_2550,N_2457);
nand U2723 (N_2723,N_2446,N_2412);
and U2724 (N_2724,N_2519,N_2570);
and U2725 (N_2725,N_2575,N_2546);
nand U2726 (N_2726,N_2424,N_2411);
nand U2727 (N_2727,N_2591,N_2401);
nor U2728 (N_2728,N_2547,N_2439);
nand U2729 (N_2729,N_2531,N_2427);
nand U2730 (N_2730,N_2561,N_2596);
or U2731 (N_2731,N_2551,N_2526);
nand U2732 (N_2732,N_2480,N_2442);
nand U2733 (N_2733,N_2482,N_2575);
xnor U2734 (N_2734,N_2598,N_2556);
nand U2735 (N_2735,N_2493,N_2400);
and U2736 (N_2736,N_2574,N_2596);
and U2737 (N_2737,N_2453,N_2482);
and U2738 (N_2738,N_2403,N_2555);
nand U2739 (N_2739,N_2575,N_2496);
xor U2740 (N_2740,N_2589,N_2512);
nor U2741 (N_2741,N_2599,N_2422);
or U2742 (N_2742,N_2544,N_2426);
and U2743 (N_2743,N_2587,N_2564);
nor U2744 (N_2744,N_2436,N_2474);
nand U2745 (N_2745,N_2427,N_2440);
nand U2746 (N_2746,N_2500,N_2511);
and U2747 (N_2747,N_2581,N_2462);
nor U2748 (N_2748,N_2542,N_2560);
or U2749 (N_2749,N_2446,N_2400);
or U2750 (N_2750,N_2526,N_2465);
nor U2751 (N_2751,N_2566,N_2461);
and U2752 (N_2752,N_2441,N_2566);
nor U2753 (N_2753,N_2464,N_2586);
nand U2754 (N_2754,N_2500,N_2441);
nor U2755 (N_2755,N_2509,N_2472);
nor U2756 (N_2756,N_2473,N_2441);
and U2757 (N_2757,N_2429,N_2464);
and U2758 (N_2758,N_2490,N_2431);
nor U2759 (N_2759,N_2461,N_2580);
nand U2760 (N_2760,N_2541,N_2591);
and U2761 (N_2761,N_2439,N_2436);
nand U2762 (N_2762,N_2593,N_2472);
nor U2763 (N_2763,N_2421,N_2459);
or U2764 (N_2764,N_2474,N_2482);
nor U2765 (N_2765,N_2439,N_2401);
nand U2766 (N_2766,N_2595,N_2524);
or U2767 (N_2767,N_2422,N_2472);
or U2768 (N_2768,N_2428,N_2463);
nor U2769 (N_2769,N_2560,N_2486);
and U2770 (N_2770,N_2593,N_2483);
nor U2771 (N_2771,N_2580,N_2582);
or U2772 (N_2772,N_2559,N_2457);
and U2773 (N_2773,N_2447,N_2537);
nor U2774 (N_2774,N_2543,N_2552);
and U2775 (N_2775,N_2459,N_2489);
and U2776 (N_2776,N_2561,N_2598);
or U2777 (N_2777,N_2594,N_2560);
nand U2778 (N_2778,N_2402,N_2481);
nand U2779 (N_2779,N_2581,N_2481);
and U2780 (N_2780,N_2588,N_2474);
nand U2781 (N_2781,N_2453,N_2548);
or U2782 (N_2782,N_2595,N_2489);
and U2783 (N_2783,N_2486,N_2459);
xnor U2784 (N_2784,N_2597,N_2446);
nand U2785 (N_2785,N_2524,N_2583);
nor U2786 (N_2786,N_2429,N_2511);
and U2787 (N_2787,N_2542,N_2568);
nor U2788 (N_2788,N_2526,N_2496);
or U2789 (N_2789,N_2554,N_2538);
nor U2790 (N_2790,N_2556,N_2403);
or U2791 (N_2791,N_2529,N_2519);
or U2792 (N_2792,N_2428,N_2585);
nand U2793 (N_2793,N_2522,N_2539);
and U2794 (N_2794,N_2456,N_2496);
nor U2795 (N_2795,N_2496,N_2406);
and U2796 (N_2796,N_2505,N_2555);
and U2797 (N_2797,N_2428,N_2509);
nor U2798 (N_2798,N_2491,N_2564);
and U2799 (N_2799,N_2477,N_2486);
nor U2800 (N_2800,N_2641,N_2654);
and U2801 (N_2801,N_2704,N_2645);
nand U2802 (N_2802,N_2670,N_2703);
and U2803 (N_2803,N_2618,N_2620);
nor U2804 (N_2804,N_2776,N_2615);
and U2805 (N_2805,N_2621,N_2724);
or U2806 (N_2806,N_2757,N_2610);
and U2807 (N_2807,N_2632,N_2760);
and U2808 (N_2808,N_2788,N_2752);
or U2809 (N_2809,N_2790,N_2695);
nand U2810 (N_2810,N_2700,N_2715);
and U2811 (N_2811,N_2678,N_2701);
nor U2812 (N_2812,N_2606,N_2635);
nand U2813 (N_2813,N_2722,N_2791);
nand U2814 (N_2814,N_2794,N_2667);
nand U2815 (N_2815,N_2633,N_2736);
nand U2816 (N_2816,N_2718,N_2772);
and U2817 (N_2817,N_2717,N_2764);
or U2818 (N_2818,N_2696,N_2751);
nand U2819 (N_2819,N_2622,N_2676);
nor U2820 (N_2820,N_2723,N_2769);
nand U2821 (N_2821,N_2627,N_2775);
nand U2822 (N_2822,N_2681,N_2677);
and U2823 (N_2823,N_2680,N_2787);
or U2824 (N_2824,N_2694,N_2662);
xor U2825 (N_2825,N_2755,N_2767);
and U2826 (N_2826,N_2626,N_2738);
nand U2827 (N_2827,N_2664,N_2669);
nand U2828 (N_2828,N_2653,N_2684);
nor U2829 (N_2829,N_2719,N_2728);
or U2830 (N_2830,N_2640,N_2793);
or U2831 (N_2831,N_2781,N_2631);
and U2832 (N_2832,N_2666,N_2609);
xnor U2833 (N_2833,N_2657,N_2605);
nor U2834 (N_2834,N_2686,N_2756);
and U2835 (N_2835,N_2766,N_2705);
or U2836 (N_2836,N_2792,N_2659);
nor U2837 (N_2837,N_2786,N_2629);
nor U2838 (N_2838,N_2762,N_2691);
nor U2839 (N_2839,N_2727,N_2785);
and U2840 (N_2840,N_2789,N_2779);
nand U2841 (N_2841,N_2730,N_2647);
nand U2842 (N_2842,N_2726,N_2674);
and U2843 (N_2843,N_2748,N_2797);
and U2844 (N_2844,N_2683,N_2668);
and U2845 (N_2845,N_2697,N_2690);
and U2846 (N_2846,N_2783,N_2709);
nand U2847 (N_2847,N_2780,N_2759);
nor U2848 (N_2848,N_2619,N_2650);
and U2849 (N_2849,N_2624,N_2744);
nand U2850 (N_2850,N_2644,N_2600);
or U2851 (N_2851,N_2665,N_2737);
nand U2852 (N_2852,N_2685,N_2692);
nand U2853 (N_2853,N_2660,N_2702);
nor U2854 (N_2854,N_2689,N_2673);
nor U2855 (N_2855,N_2616,N_2698);
and U2856 (N_2856,N_2774,N_2603);
nor U2857 (N_2857,N_2617,N_2763);
or U2858 (N_2858,N_2799,N_2754);
or U2859 (N_2859,N_2639,N_2636);
and U2860 (N_2860,N_2712,N_2604);
and U2861 (N_2861,N_2743,N_2648);
nor U2862 (N_2862,N_2651,N_2740);
nand U2863 (N_2863,N_2777,N_2601);
nor U2864 (N_2864,N_2658,N_2773);
nand U2865 (N_2865,N_2771,N_2634);
or U2866 (N_2866,N_2699,N_2638);
nor U2867 (N_2867,N_2642,N_2746);
nand U2868 (N_2868,N_2649,N_2679);
nand U2869 (N_2869,N_2725,N_2770);
and U2870 (N_2870,N_2623,N_2735);
nor U2871 (N_2871,N_2671,N_2782);
nand U2872 (N_2872,N_2646,N_2784);
nand U2873 (N_2873,N_2706,N_2687);
or U2874 (N_2874,N_2675,N_2655);
or U2875 (N_2875,N_2768,N_2613);
or U2876 (N_2876,N_2795,N_2682);
or U2877 (N_2877,N_2672,N_2652);
or U2878 (N_2878,N_2628,N_2753);
nand U2879 (N_2879,N_2796,N_2749);
or U2880 (N_2880,N_2625,N_2612);
nand U2881 (N_2881,N_2731,N_2602);
nor U2882 (N_2882,N_2630,N_2721);
xnor U2883 (N_2883,N_2661,N_2729);
or U2884 (N_2884,N_2741,N_2614);
nand U2885 (N_2885,N_2607,N_2693);
nand U2886 (N_2886,N_2608,N_2643);
and U2887 (N_2887,N_2714,N_2758);
nand U2888 (N_2888,N_2739,N_2710);
nor U2889 (N_2889,N_2663,N_2745);
and U2890 (N_2890,N_2713,N_2747);
nand U2891 (N_2891,N_2637,N_2656);
nor U2892 (N_2892,N_2720,N_2716);
and U2893 (N_2893,N_2742,N_2798);
and U2894 (N_2894,N_2688,N_2765);
and U2895 (N_2895,N_2611,N_2734);
nand U2896 (N_2896,N_2732,N_2711);
nor U2897 (N_2897,N_2733,N_2778);
nor U2898 (N_2898,N_2761,N_2750);
and U2899 (N_2899,N_2707,N_2708);
nand U2900 (N_2900,N_2693,N_2766);
and U2901 (N_2901,N_2791,N_2666);
and U2902 (N_2902,N_2764,N_2785);
nor U2903 (N_2903,N_2662,N_2707);
nand U2904 (N_2904,N_2616,N_2658);
nand U2905 (N_2905,N_2717,N_2735);
or U2906 (N_2906,N_2758,N_2622);
and U2907 (N_2907,N_2605,N_2752);
or U2908 (N_2908,N_2606,N_2647);
nor U2909 (N_2909,N_2769,N_2795);
nand U2910 (N_2910,N_2685,N_2748);
nor U2911 (N_2911,N_2635,N_2662);
nand U2912 (N_2912,N_2707,N_2612);
or U2913 (N_2913,N_2765,N_2714);
nor U2914 (N_2914,N_2766,N_2729);
and U2915 (N_2915,N_2791,N_2772);
and U2916 (N_2916,N_2653,N_2619);
nor U2917 (N_2917,N_2756,N_2674);
or U2918 (N_2918,N_2779,N_2701);
or U2919 (N_2919,N_2683,N_2650);
nand U2920 (N_2920,N_2696,N_2694);
and U2921 (N_2921,N_2773,N_2767);
or U2922 (N_2922,N_2663,N_2743);
and U2923 (N_2923,N_2796,N_2713);
or U2924 (N_2924,N_2655,N_2717);
nor U2925 (N_2925,N_2787,N_2748);
nand U2926 (N_2926,N_2695,N_2652);
or U2927 (N_2927,N_2695,N_2615);
nor U2928 (N_2928,N_2777,N_2621);
nor U2929 (N_2929,N_2737,N_2713);
nor U2930 (N_2930,N_2796,N_2784);
or U2931 (N_2931,N_2605,N_2645);
and U2932 (N_2932,N_2721,N_2752);
nor U2933 (N_2933,N_2668,N_2734);
or U2934 (N_2934,N_2673,N_2632);
xnor U2935 (N_2935,N_2782,N_2606);
or U2936 (N_2936,N_2662,N_2759);
nand U2937 (N_2937,N_2669,N_2732);
xor U2938 (N_2938,N_2636,N_2612);
nor U2939 (N_2939,N_2776,N_2738);
and U2940 (N_2940,N_2725,N_2722);
nor U2941 (N_2941,N_2795,N_2775);
or U2942 (N_2942,N_2753,N_2617);
or U2943 (N_2943,N_2608,N_2731);
nand U2944 (N_2944,N_2782,N_2614);
nor U2945 (N_2945,N_2615,N_2740);
nand U2946 (N_2946,N_2612,N_2683);
nor U2947 (N_2947,N_2697,N_2631);
or U2948 (N_2948,N_2705,N_2775);
nor U2949 (N_2949,N_2794,N_2790);
or U2950 (N_2950,N_2708,N_2610);
or U2951 (N_2951,N_2688,N_2624);
nand U2952 (N_2952,N_2725,N_2792);
or U2953 (N_2953,N_2683,N_2739);
or U2954 (N_2954,N_2658,N_2637);
nand U2955 (N_2955,N_2623,N_2777);
and U2956 (N_2956,N_2696,N_2739);
nor U2957 (N_2957,N_2766,N_2646);
nand U2958 (N_2958,N_2694,N_2607);
nor U2959 (N_2959,N_2671,N_2775);
or U2960 (N_2960,N_2662,N_2649);
nand U2961 (N_2961,N_2761,N_2753);
and U2962 (N_2962,N_2783,N_2732);
or U2963 (N_2963,N_2668,N_2793);
or U2964 (N_2964,N_2695,N_2770);
or U2965 (N_2965,N_2765,N_2770);
or U2966 (N_2966,N_2646,N_2731);
nand U2967 (N_2967,N_2605,N_2677);
nor U2968 (N_2968,N_2799,N_2737);
and U2969 (N_2969,N_2712,N_2676);
nand U2970 (N_2970,N_2771,N_2670);
nor U2971 (N_2971,N_2726,N_2734);
or U2972 (N_2972,N_2663,N_2750);
nor U2973 (N_2973,N_2763,N_2651);
nor U2974 (N_2974,N_2662,N_2633);
and U2975 (N_2975,N_2647,N_2712);
nor U2976 (N_2976,N_2799,N_2740);
xnor U2977 (N_2977,N_2775,N_2711);
or U2978 (N_2978,N_2726,N_2713);
or U2979 (N_2979,N_2719,N_2737);
nor U2980 (N_2980,N_2743,N_2767);
and U2981 (N_2981,N_2791,N_2717);
nand U2982 (N_2982,N_2723,N_2765);
or U2983 (N_2983,N_2752,N_2778);
and U2984 (N_2984,N_2747,N_2739);
nor U2985 (N_2985,N_2729,N_2693);
nor U2986 (N_2986,N_2731,N_2708);
and U2987 (N_2987,N_2675,N_2769);
and U2988 (N_2988,N_2689,N_2755);
nor U2989 (N_2989,N_2716,N_2660);
and U2990 (N_2990,N_2747,N_2638);
nand U2991 (N_2991,N_2643,N_2774);
nor U2992 (N_2992,N_2704,N_2613);
nor U2993 (N_2993,N_2673,N_2653);
nand U2994 (N_2994,N_2634,N_2678);
nor U2995 (N_2995,N_2778,N_2754);
nor U2996 (N_2996,N_2754,N_2711);
and U2997 (N_2997,N_2706,N_2711);
nor U2998 (N_2998,N_2673,N_2734);
and U2999 (N_2999,N_2703,N_2662);
nand UO_0 (O_0,N_2995,N_2805);
nor UO_1 (O_1,N_2918,N_2831);
or UO_2 (O_2,N_2802,N_2987);
and UO_3 (O_3,N_2904,N_2975);
or UO_4 (O_4,N_2920,N_2957);
nor UO_5 (O_5,N_2858,N_2908);
nand UO_6 (O_6,N_2958,N_2828);
and UO_7 (O_7,N_2868,N_2985);
and UO_8 (O_8,N_2809,N_2980);
nor UO_9 (O_9,N_2999,N_2994);
or UO_10 (O_10,N_2942,N_2861);
nor UO_11 (O_11,N_2887,N_2978);
and UO_12 (O_12,N_2924,N_2945);
xnor UO_13 (O_13,N_2849,N_2899);
and UO_14 (O_14,N_2955,N_2867);
and UO_15 (O_15,N_2962,N_2922);
and UO_16 (O_16,N_2934,N_2921);
nor UO_17 (O_17,N_2923,N_2984);
and UO_18 (O_18,N_2927,N_2818);
nor UO_19 (O_19,N_2990,N_2916);
nand UO_20 (O_20,N_2824,N_2979);
nand UO_21 (O_21,N_2996,N_2825);
and UO_22 (O_22,N_2911,N_2977);
and UO_23 (O_23,N_2829,N_2865);
or UO_24 (O_24,N_2917,N_2915);
xor UO_25 (O_25,N_2866,N_2813);
nor UO_26 (O_26,N_2953,N_2823);
nand UO_27 (O_27,N_2933,N_2885);
or UO_28 (O_28,N_2998,N_2848);
nand UO_29 (O_29,N_2811,N_2935);
nand UO_30 (O_30,N_2870,N_2983);
and UO_31 (O_31,N_2949,N_2986);
and UO_32 (O_32,N_2929,N_2896);
or UO_33 (O_33,N_2940,N_2952);
nand UO_34 (O_34,N_2863,N_2902);
and UO_35 (O_35,N_2954,N_2956);
or UO_36 (O_36,N_2857,N_2821);
nor UO_37 (O_37,N_2807,N_2835);
nand UO_38 (O_38,N_2841,N_2910);
or UO_39 (O_39,N_2886,N_2888);
and UO_40 (O_40,N_2842,N_2951);
or UO_41 (O_41,N_2972,N_2897);
and UO_42 (O_42,N_2822,N_2851);
nand UO_43 (O_43,N_2879,N_2932);
nor UO_44 (O_44,N_2838,N_2905);
and UO_45 (O_45,N_2854,N_2968);
nand UO_46 (O_46,N_2846,N_2875);
nor UO_47 (O_47,N_2872,N_2852);
and UO_48 (O_48,N_2836,N_2860);
nand UO_49 (O_49,N_2890,N_2815);
nand UO_50 (O_50,N_2859,N_2943);
and UO_51 (O_51,N_2901,N_2817);
nand UO_52 (O_52,N_2873,N_2830);
or UO_53 (O_53,N_2981,N_2840);
nor UO_54 (O_54,N_2844,N_2970);
and UO_55 (O_55,N_2993,N_2938);
or UO_56 (O_56,N_2876,N_2903);
xor UO_57 (O_57,N_2883,N_2966);
nor UO_58 (O_58,N_2941,N_2937);
and UO_59 (O_59,N_2950,N_2961);
nor UO_60 (O_60,N_2832,N_2810);
and UO_61 (O_61,N_2967,N_2856);
nor UO_62 (O_62,N_2965,N_2837);
and UO_63 (O_63,N_2827,N_2880);
and UO_64 (O_64,N_2892,N_2936);
nand UO_65 (O_65,N_2882,N_2812);
and UO_66 (O_66,N_2845,N_2847);
and UO_67 (O_67,N_2874,N_2826);
nor UO_68 (O_68,N_2804,N_2900);
or UO_69 (O_69,N_2928,N_2948);
nand UO_70 (O_70,N_2925,N_2862);
nor UO_71 (O_71,N_2895,N_2871);
and UO_72 (O_72,N_2839,N_2833);
nor UO_73 (O_73,N_2930,N_2906);
and UO_74 (O_74,N_2960,N_2806);
nand UO_75 (O_75,N_2808,N_2814);
and UO_76 (O_76,N_2878,N_2801);
nand UO_77 (O_77,N_2800,N_2819);
nand UO_78 (O_78,N_2969,N_2894);
nand UO_79 (O_79,N_2881,N_2988);
nand UO_80 (O_80,N_2869,N_2947);
nor UO_81 (O_81,N_2914,N_2919);
nand UO_82 (O_82,N_2971,N_2982);
and UO_83 (O_83,N_2891,N_2959);
nor UO_84 (O_84,N_2991,N_2974);
or UO_85 (O_85,N_2926,N_2843);
nand UO_86 (O_86,N_2893,N_2884);
nand UO_87 (O_87,N_2964,N_2909);
nand UO_88 (O_88,N_2976,N_2992);
nand UO_89 (O_89,N_2939,N_2834);
and UO_90 (O_90,N_2946,N_2944);
nand UO_91 (O_91,N_2997,N_2853);
and UO_92 (O_92,N_2889,N_2803);
nand UO_93 (O_93,N_2877,N_2855);
or UO_94 (O_94,N_2816,N_2989);
and UO_95 (O_95,N_2913,N_2850);
nand UO_96 (O_96,N_2907,N_2820);
and UO_97 (O_97,N_2898,N_2963);
nor UO_98 (O_98,N_2864,N_2973);
and UO_99 (O_99,N_2931,N_2912);
or UO_100 (O_100,N_2849,N_2999);
nand UO_101 (O_101,N_2830,N_2986);
and UO_102 (O_102,N_2991,N_2866);
nor UO_103 (O_103,N_2999,N_2820);
nand UO_104 (O_104,N_2889,N_2863);
nor UO_105 (O_105,N_2868,N_2917);
nor UO_106 (O_106,N_2925,N_2844);
nand UO_107 (O_107,N_2874,N_2891);
nand UO_108 (O_108,N_2987,N_2821);
nand UO_109 (O_109,N_2831,N_2808);
nand UO_110 (O_110,N_2987,N_2997);
and UO_111 (O_111,N_2995,N_2807);
nand UO_112 (O_112,N_2815,N_2928);
and UO_113 (O_113,N_2829,N_2816);
nand UO_114 (O_114,N_2824,N_2813);
nor UO_115 (O_115,N_2840,N_2910);
nor UO_116 (O_116,N_2992,N_2956);
and UO_117 (O_117,N_2890,N_2969);
or UO_118 (O_118,N_2857,N_2907);
nor UO_119 (O_119,N_2914,N_2857);
nor UO_120 (O_120,N_2804,N_2936);
and UO_121 (O_121,N_2982,N_2966);
or UO_122 (O_122,N_2935,N_2952);
and UO_123 (O_123,N_2861,N_2903);
nor UO_124 (O_124,N_2947,N_2845);
and UO_125 (O_125,N_2941,N_2913);
and UO_126 (O_126,N_2933,N_2881);
nor UO_127 (O_127,N_2811,N_2857);
or UO_128 (O_128,N_2972,N_2954);
or UO_129 (O_129,N_2961,N_2888);
nand UO_130 (O_130,N_2912,N_2986);
and UO_131 (O_131,N_2830,N_2884);
or UO_132 (O_132,N_2835,N_2885);
nor UO_133 (O_133,N_2806,N_2883);
or UO_134 (O_134,N_2840,N_2894);
nand UO_135 (O_135,N_2876,N_2964);
and UO_136 (O_136,N_2932,N_2956);
nor UO_137 (O_137,N_2934,N_2949);
nand UO_138 (O_138,N_2901,N_2873);
or UO_139 (O_139,N_2993,N_2859);
nand UO_140 (O_140,N_2943,N_2911);
and UO_141 (O_141,N_2818,N_2877);
or UO_142 (O_142,N_2920,N_2914);
or UO_143 (O_143,N_2857,N_2961);
nor UO_144 (O_144,N_2925,N_2851);
nand UO_145 (O_145,N_2832,N_2954);
or UO_146 (O_146,N_2920,N_2901);
nand UO_147 (O_147,N_2961,N_2942);
and UO_148 (O_148,N_2864,N_2984);
nor UO_149 (O_149,N_2883,N_2997);
or UO_150 (O_150,N_2879,N_2916);
nand UO_151 (O_151,N_2965,N_2940);
or UO_152 (O_152,N_2830,N_2856);
nand UO_153 (O_153,N_2821,N_2977);
and UO_154 (O_154,N_2894,N_2944);
and UO_155 (O_155,N_2849,N_2894);
nor UO_156 (O_156,N_2923,N_2958);
nor UO_157 (O_157,N_2998,N_2941);
nor UO_158 (O_158,N_2986,N_2988);
or UO_159 (O_159,N_2991,N_2802);
nand UO_160 (O_160,N_2803,N_2823);
and UO_161 (O_161,N_2958,N_2954);
nor UO_162 (O_162,N_2884,N_2853);
and UO_163 (O_163,N_2942,N_2906);
xnor UO_164 (O_164,N_2950,N_2828);
nor UO_165 (O_165,N_2909,N_2938);
nor UO_166 (O_166,N_2847,N_2808);
and UO_167 (O_167,N_2876,N_2946);
or UO_168 (O_168,N_2921,N_2994);
nor UO_169 (O_169,N_2854,N_2904);
or UO_170 (O_170,N_2989,N_2874);
nand UO_171 (O_171,N_2873,N_2975);
or UO_172 (O_172,N_2826,N_2986);
and UO_173 (O_173,N_2954,N_2910);
nor UO_174 (O_174,N_2897,N_2986);
or UO_175 (O_175,N_2951,N_2981);
or UO_176 (O_176,N_2933,N_2832);
nor UO_177 (O_177,N_2853,N_2950);
and UO_178 (O_178,N_2857,N_2927);
nand UO_179 (O_179,N_2844,N_2917);
and UO_180 (O_180,N_2978,N_2846);
nand UO_181 (O_181,N_2994,N_2954);
nand UO_182 (O_182,N_2877,N_2971);
nor UO_183 (O_183,N_2907,N_2867);
nand UO_184 (O_184,N_2940,N_2869);
and UO_185 (O_185,N_2811,N_2816);
nor UO_186 (O_186,N_2905,N_2901);
nand UO_187 (O_187,N_2924,N_2944);
and UO_188 (O_188,N_2913,N_2961);
and UO_189 (O_189,N_2994,N_2975);
and UO_190 (O_190,N_2971,N_2825);
nor UO_191 (O_191,N_2868,N_2961);
nand UO_192 (O_192,N_2982,N_2858);
and UO_193 (O_193,N_2859,N_2964);
nand UO_194 (O_194,N_2800,N_2918);
and UO_195 (O_195,N_2853,N_2819);
or UO_196 (O_196,N_2860,N_2964);
or UO_197 (O_197,N_2848,N_2827);
and UO_198 (O_198,N_2967,N_2875);
or UO_199 (O_199,N_2993,N_2951);
nand UO_200 (O_200,N_2899,N_2822);
nand UO_201 (O_201,N_2984,N_2837);
nor UO_202 (O_202,N_2853,N_2877);
or UO_203 (O_203,N_2985,N_2962);
and UO_204 (O_204,N_2993,N_2910);
nand UO_205 (O_205,N_2985,N_2931);
nand UO_206 (O_206,N_2835,N_2902);
and UO_207 (O_207,N_2998,N_2984);
nor UO_208 (O_208,N_2901,N_2889);
or UO_209 (O_209,N_2860,N_2845);
nor UO_210 (O_210,N_2911,N_2927);
nand UO_211 (O_211,N_2912,N_2992);
nor UO_212 (O_212,N_2816,N_2805);
or UO_213 (O_213,N_2997,N_2921);
xnor UO_214 (O_214,N_2920,N_2894);
nand UO_215 (O_215,N_2905,N_2886);
and UO_216 (O_216,N_2993,N_2909);
nor UO_217 (O_217,N_2922,N_2809);
nor UO_218 (O_218,N_2877,N_2881);
and UO_219 (O_219,N_2921,N_2989);
or UO_220 (O_220,N_2966,N_2809);
nand UO_221 (O_221,N_2979,N_2960);
nor UO_222 (O_222,N_2989,N_2920);
nand UO_223 (O_223,N_2813,N_2890);
and UO_224 (O_224,N_2883,N_2840);
or UO_225 (O_225,N_2844,N_2900);
and UO_226 (O_226,N_2922,N_2878);
nand UO_227 (O_227,N_2883,N_2977);
nor UO_228 (O_228,N_2924,N_2962);
and UO_229 (O_229,N_2932,N_2851);
and UO_230 (O_230,N_2887,N_2881);
or UO_231 (O_231,N_2929,N_2940);
and UO_232 (O_232,N_2940,N_2937);
or UO_233 (O_233,N_2846,N_2821);
or UO_234 (O_234,N_2882,N_2933);
and UO_235 (O_235,N_2837,N_2855);
or UO_236 (O_236,N_2859,N_2920);
nand UO_237 (O_237,N_2822,N_2890);
nand UO_238 (O_238,N_2887,N_2993);
nand UO_239 (O_239,N_2833,N_2842);
or UO_240 (O_240,N_2913,N_2806);
or UO_241 (O_241,N_2859,N_2834);
nor UO_242 (O_242,N_2902,N_2932);
xnor UO_243 (O_243,N_2834,N_2836);
xnor UO_244 (O_244,N_2849,N_2942);
nor UO_245 (O_245,N_2982,N_2854);
nor UO_246 (O_246,N_2989,N_2990);
and UO_247 (O_247,N_2803,N_2893);
nor UO_248 (O_248,N_2991,N_2819);
nand UO_249 (O_249,N_2821,N_2926);
and UO_250 (O_250,N_2891,N_2857);
or UO_251 (O_251,N_2900,N_2828);
and UO_252 (O_252,N_2892,N_2845);
nor UO_253 (O_253,N_2850,N_2820);
or UO_254 (O_254,N_2917,N_2910);
nand UO_255 (O_255,N_2967,N_2817);
and UO_256 (O_256,N_2945,N_2868);
nand UO_257 (O_257,N_2833,N_2975);
nor UO_258 (O_258,N_2968,N_2929);
or UO_259 (O_259,N_2999,N_2916);
or UO_260 (O_260,N_2805,N_2864);
nand UO_261 (O_261,N_2994,N_2806);
and UO_262 (O_262,N_2979,N_2935);
and UO_263 (O_263,N_2839,N_2954);
nor UO_264 (O_264,N_2861,N_2830);
or UO_265 (O_265,N_2873,N_2816);
and UO_266 (O_266,N_2896,N_2856);
or UO_267 (O_267,N_2896,N_2804);
nor UO_268 (O_268,N_2926,N_2875);
and UO_269 (O_269,N_2988,N_2987);
nor UO_270 (O_270,N_2864,N_2840);
and UO_271 (O_271,N_2868,N_2829);
or UO_272 (O_272,N_2863,N_2961);
or UO_273 (O_273,N_2861,N_2922);
nand UO_274 (O_274,N_2851,N_2985);
nand UO_275 (O_275,N_2921,N_2885);
and UO_276 (O_276,N_2820,N_2838);
and UO_277 (O_277,N_2879,N_2974);
nor UO_278 (O_278,N_2806,N_2958);
xnor UO_279 (O_279,N_2987,N_2878);
or UO_280 (O_280,N_2979,N_2889);
nand UO_281 (O_281,N_2851,N_2903);
nor UO_282 (O_282,N_2954,N_2976);
and UO_283 (O_283,N_2926,N_2831);
and UO_284 (O_284,N_2948,N_2834);
or UO_285 (O_285,N_2917,N_2817);
and UO_286 (O_286,N_2880,N_2817);
and UO_287 (O_287,N_2996,N_2936);
or UO_288 (O_288,N_2828,N_2917);
nor UO_289 (O_289,N_2961,N_2890);
or UO_290 (O_290,N_2840,N_2857);
nor UO_291 (O_291,N_2894,N_2911);
and UO_292 (O_292,N_2942,N_2933);
and UO_293 (O_293,N_2953,N_2960);
nand UO_294 (O_294,N_2839,N_2840);
and UO_295 (O_295,N_2953,N_2864);
xor UO_296 (O_296,N_2982,N_2979);
and UO_297 (O_297,N_2867,N_2944);
nand UO_298 (O_298,N_2923,N_2834);
nand UO_299 (O_299,N_2821,N_2916);
nor UO_300 (O_300,N_2966,N_2970);
nor UO_301 (O_301,N_2849,N_2976);
or UO_302 (O_302,N_2936,N_2954);
or UO_303 (O_303,N_2949,N_2821);
and UO_304 (O_304,N_2844,N_2954);
and UO_305 (O_305,N_2878,N_2963);
nand UO_306 (O_306,N_2948,N_2878);
and UO_307 (O_307,N_2944,N_2866);
or UO_308 (O_308,N_2924,N_2932);
or UO_309 (O_309,N_2933,N_2883);
nor UO_310 (O_310,N_2948,N_2815);
xor UO_311 (O_311,N_2959,N_2800);
or UO_312 (O_312,N_2898,N_2815);
and UO_313 (O_313,N_2892,N_2853);
and UO_314 (O_314,N_2848,N_2907);
or UO_315 (O_315,N_2987,N_2897);
or UO_316 (O_316,N_2910,N_2919);
and UO_317 (O_317,N_2845,N_2846);
nor UO_318 (O_318,N_2902,N_2983);
and UO_319 (O_319,N_2873,N_2870);
or UO_320 (O_320,N_2849,N_2992);
nor UO_321 (O_321,N_2996,N_2935);
and UO_322 (O_322,N_2919,N_2876);
or UO_323 (O_323,N_2896,N_2949);
nor UO_324 (O_324,N_2861,N_2824);
or UO_325 (O_325,N_2893,N_2812);
nand UO_326 (O_326,N_2867,N_2823);
nor UO_327 (O_327,N_2979,N_2902);
nand UO_328 (O_328,N_2849,N_2858);
and UO_329 (O_329,N_2862,N_2965);
and UO_330 (O_330,N_2949,N_2857);
or UO_331 (O_331,N_2813,N_2861);
nor UO_332 (O_332,N_2873,N_2890);
or UO_333 (O_333,N_2878,N_2938);
nand UO_334 (O_334,N_2845,N_2865);
nor UO_335 (O_335,N_2944,N_2855);
or UO_336 (O_336,N_2845,N_2823);
or UO_337 (O_337,N_2931,N_2915);
and UO_338 (O_338,N_2903,N_2899);
or UO_339 (O_339,N_2988,N_2939);
and UO_340 (O_340,N_2931,N_2845);
or UO_341 (O_341,N_2871,N_2910);
nand UO_342 (O_342,N_2980,N_2993);
and UO_343 (O_343,N_2853,N_2824);
and UO_344 (O_344,N_2879,N_2810);
nor UO_345 (O_345,N_2830,N_2807);
and UO_346 (O_346,N_2953,N_2965);
nand UO_347 (O_347,N_2958,N_2900);
nor UO_348 (O_348,N_2870,N_2956);
xor UO_349 (O_349,N_2905,N_2851);
or UO_350 (O_350,N_2819,N_2922);
nand UO_351 (O_351,N_2940,N_2927);
and UO_352 (O_352,N_2817,N_2977);
nand UO_353 (O_353,N_2878,N_2872);
nor UO_354 (O_354,N_2972,N_2833);
nor UO_355 (O_355,N_2971,N_2808);
nand UO_356 (O_356,N_2825,N_2909);
nor UO_357 (O_357,N_2913,N_2940);
or UO_358 (O_358,N_2897,N_2956);
nand UO_359 (O_359,N_2883,N_2853);
nor UO_360 (O_360,N_2923,N_2955);
and UO_361 (O_361,N_2817,N_2841);
nand UO_362 (O_362,N_2875,N_2825);
nand UO_363 (O_363,N_2940,N_2951);
or UO_364 (O_364,N_2984,N_2808);
nor UO_365 (O_365,N_2908,N_2879);
or UO_366 (O_366,N_2952,N_2921);
or UO_367 (O_367,N_2927,N_2977);
or UO_368 (O_368,N_2827,N_2812);
or UO_369 (O_369,N_2907,N_2854);
nor UO_370 (O_370,N_2982,N_2994);
or UO_371 (O_371,N_2825,N_2931);
and UO_372 (O_372,N_2853,N_2800);
nor UO_373 (O_373,N_2900,N_2871);
or UO_374 (O_374,N_2839,N_2927);
or UO_375 (O_375,N_2927,N_2908);
or UO_376 (O_376,N_2809,N_2931);
nand UO_377 (O_377,N_2871,N_2889);
and UO_378 (O_378,N_2923,N_2840);
and UO_379 (O_379,N_2949,N_2985);
and UO_380 (O_380,N_2888,N_2825);
or UO_381 (O_381,N_2940,N_2839);
and UO_382 (O_382,N_2804,N_2818);
or UO_383 (O_383,N_2966,N_2983);
nor UO_384 (O_384,N_2930,N_2849);
and UO_385 (O_385,N_2887,N_2990);
and UO_386 (O_386,N_2807,N_2819);
and UO_387 (O_387,N_2974,N_2876);
nand UO_388 (O_388,N_2978,N_2944);
nor UO_389 (O_389,N_2822,N_2913);
nor UO_390 (O_390,N_2823,N_2898);
and UO_391 (O_391,N_2833,N_2816);
nand UO_392 (O_392,N_2985,N_2810);
nor UO_393 (O_393,N_2902,N_2847);
or UO_394 (O_394,N_2859,N_2900);
nand UO_395 (O_395,N_2953,N_2955);
nor UO_396 (O_396,N_2983,N_2815);
and UO_397 (O_397,N_2904,N_2886);
nand UO_398 (O_398,N_2875,N_2889);
or UO_399 (O_399,N_2955,N_2914);
nand UO_400 (O_400,N_2951,N_2861);
or UO_401 (O_401,N_2852,N_2882);
or UO_402 (O_402,N_2923,N_2873);
xnor UO_403 (O_403,N_2817,N_2882);
nand UO_404 (O_404,N_2963,N_2841);
and UO_405 (O_405,N_2912,N_2981);
nor UO_406 (O_406,N_2951,N_2964);
nand UO_407 (O_407,N_2811,N_2840);
nor UO_408 (O_408,N_2949,N_2872);
or UO_409 (O_409,N_2875,N_2886);
and UO_410 (O_410,N_2983,N_2900);
nand UO_411 (O_411,N_2812,N_2938);
or UO_412 (O_412,N_2833,N_2911);
xor UO_413 (O_413,N_2902,N_2908);
nand UO_414 (O_414,N_2992,N_2968);
nor UO_415 (O_415,N_2941,N_2930);
or UO_416 (O_416,N_2935,N_2987);
nand UO_417 (O_417,N_2914,N_2816);
or UO_418 (O_418,N_2849,N_2831);
or UO_419 (O_419,N_2828,N_2830);
nand UO_420 (O_420,N_2974,N_2936);
nor UO_421 (O_421,N_2917,N_2808);
nor UO_422 (O_422,N_2937,N_2976);
nand UO_423 (O_423,N_2961,N_2870);
or UO_424 (O_424,N_2952,N_2892);
nand UO_425 (O_425,N_2801,N_2886);
and UO_426 (O_426,N_2910,N_2979);
nor UO_427 (O_427,N_2944,N_2969);
nand UO_428 (O_428,N_2801,N_2852);
nor UO_429 (O_429,N_2944,N_2868);
and UO_430 (O_430,N_2938,N_2917);
and UO_431 (O_431,N_2877,N_2897);
and UO_432 (O_432,N_2932,N_2986);
xnor UO_433 (O_433,N_2981,N_2936);
nand UO_434 (O_434,N_2899,N_2971);
nand UO_435 (O_435,N_2880,N_2940);
nor UO_436 (O_436,N_2945,N_2972);
nor UO_437 (O_437,N_2832,N_2857);
nand UO_438 (O_438,N_2915,N_2908);
or UO_439 (O_439,N_2805,N_2947);
nor UO_440 (O_440,N_2913,N_2938);
and UO_441 (O_441,N_2812,N_2873);
and UO_442 (O_442,N_2969,N_2922);
nand UO_443 (O_443,N_2914,N_2917);
nand UO_444 (O_444,N_2928,N_2983);
nor UO_445 (O_445,N_2991,N_2907);
and UO_446 (O_446,N_2832,N_2969);
nand UO_447 (O_447,N_2903,N_2887);
nand UO_448 (O_448,N_2825,N_2919);
nor UO_449 (O_449,N_2807,N_2964);
or UO_450 (O_450,N_2866,N_2858);
nor UO_451 (O_451,N_2979,N_2883);
and UO_452 (O_452,N_2801,N_2803);
and UO_453 (O_453,N_2879,N_2985);
and UO_454 (O_454,N_2814,N_2969);
nor UO_455 (O_455,N_2909,N_2984);
nand UO_456 (O_456,N_2938,N_2886);
or UO_457 (O_457,N_2880,N_2809);
or UO_458 (O_458,N_2830,N_2903);
xor UO_459 (O_459,N_2918,N_2829);
and UO_460 (O_460,N_2820,N_2944);
or UO_461 (O_461,N_2965,N_2971);
nor UO_462 (O_462,N_2824,N_2908);
nand UO_463 (O_463,N_2956,N_2835);
nand UO_464 (O_464,N_2925,N_2984);
nand UO_465 (O_465,N_2836,N_2800);
nand UO_466 (O_466,N_2814,N_2826);
nand UO_467 (O_467,N_2962,N_2927);
and UO_468 (O_468,N_2927,N_2806);
or UO_469 (O_469,N_2850,N_2947);
or UO_470 (O_470,N_2853,N_2990);
or UO_471 (O_471,N_2830,N_2976);
nand UO_472 (O_472,N_2934,N_2857);
nor UO_473 (O_473,N_2819,N_2971);
nand UO_474 (O_474,N_2886,N_2808);
nor UO_475 (O_475,N_2896,N_2987);
and UO_476 (O_476,N_2894,N_2845);
nand UO_477 (O_477,N_2919,N_2814);
and UO_478 (O_478,N_2823,N_2965);
nand UO_479 (O_479,N_2992,N_2854);
nor UO_480 (O_480,N_2975,N_2867);
nor UO_481 (O_481,N_2832,N_2992);
or UO_482 (O_482,N_2953,N_2928);
nand UO_483 (O_483,N_2959,N_2857);
or UO_484 (O_484,N_2863,N_2972);
nor UO_485 (O_485,N_2803,N_2963);
xnor UO_486 (O_486,N_2900,N_2839);
nor UO_487 (O_487,N_2831,N_2992);
or UO_488 (O_488,N_2893,N_2994);
nand UO_489 (O_489,N_2929,N_2860);
or UO_490 (O_490,N_2836,N_2866);
nor UO_491 (O_491,N_2888,N_2880);
or UO_492 (O_492,N_2921,N_2801);
and UO_493 (O_493,N_2993,N_2835);
or UO_494 (O_494,N_2841,N_2801);
or UO_495 (O_495,N_2986,N_2968);
nand UO_496 (O_496,N_2863,N_2869);
nor UO_497 (O_497,N_2863,N_2947);
and UO_498 (O_498,N_2803,N_2845);
nand UO_499 (O_499,N_2853,N_2821);
endmodule