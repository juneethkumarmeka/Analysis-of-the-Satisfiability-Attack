module basic_500_3000_500_15_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_339,In_347);
nand U1 (N_1,In_160,In_389);
nor U2 (N_2,In_401,In_155);
and U3 (N_3,In_144,In_212);
or U4 (N_4,In_345,In_124);
or U5 (N_5,In_56,In_327);
nand U6 (N_6,In_117,In_430);
and U7 (N_7,In_78,In_385);
nor U8 (N_8,In_73,In_461);
or U9 (N_9,In_485,In_261);
nor U10 (N_10,In_397,In_265);
and U11 (N_11,In_6,In_443);
and U12 (N_12,In_184,In_278);
xnor U13 (N_13,In_448,In_340);
nand U14 (N_14,In_442,In_412);
nor U15 (N_15,In_491,In_264);
or U16 (N_16,In_380,In_497);
or U17 (N_17,In_115,In_426);
nand U18 (N_18,In_0,In_89);
nor U19 (N_19,In_378,In_427);
nand U20 (N_20,In_473,In_197);
and U21 (N_21,In_464,In_23);
nor U22 (N_22,In_239,In_13);
and U23 (N_23,In_478,In_210);
and U24 (N_24,In_268,In_422);
or U25 (N_25,In_163,In_175);
and U26 (N_26,In_365,In_384);
or U27 (N_27,In_146,In_61);
and U28 (N_28,In_468,In_475);
nor U29 (N_29,In_208,In_387);
nand U30 (N_30,In_279,In_52);
nand U31 (N_31,In_315,In_31);
nand U32 (N_32,In_43,In_157);
nor U33 (N_33,In_220,In_330);
and U34 (N_34,In_323,In_394);
nor U35 (N_35,In_60,In_313);
nor U36 (N_36,In_293,In_272);
nor U37 (N_37,In_12,In_71);
nand U38 (N_38,In_351,In_181);
nand U39 (N_39,In_375,In_454);
or U40 (N_40,In_236,In_27);
nand U41 (N_41,In_198,In_98);
nor U42 (N_42,In_74,In_428);
and U43 (N_43,In_64,In_70);
nor U44 (N_44,In_492,In_67);
xnor U45 (N_45,In_472,In_241);
nor U46 (N_46,In_455,In_34);
or U47 (N_47,In_259,In_128);
and U48 (N_48,In_438,In_221);
or U49 (N_49,In_307,In_270);
nor U50 (N_50,In_29,In_263);
and U51 (N_51,In_53,In_18);
nor U52 (N_52,In_479,In_217);
nor U53 (N_53,In_229,In_228);
nor U54 (N_54,In_143,In_247);
or U55 (N_55,In_425,In_266);
and U56 (N_56,In_164,In_90);
nand U57 (N_57,In_242,In_3);
or U58 (N_58,In_363,In_314);
nor U59 (N_59,In_85,In_233);
and U60 (N_60,In_255,In_100);
nand U61 (N_61,In_230,In_133);
nand U62 (N_62,In_459,In_406);
nor U63 (N_63,In_77,In_226);
nand U64 (N_64,In_306,In_321);
xnor U65 (N_65,In_285,In_420);
nor U66 (N_66,In_59,In_84);
xor U67 (N_67,In_48,In_349);
and U68 (N_68,In_431,In_134);
nor U69 (N_69,In_203,In_361);
nand U70 (N_70,In_209,In_395);
nand U71 (N_71,In_246,In_130);
or U72 (N_72,In_477,In_445);
or U73 (N_73,In_119,In_167);
and U74 (N_74,In_196,In_334);
nand U75 (N_75,In_471,In_114);
and U76 (N_76,In_486,In_251);
or U77 (N_77,In_487,In_419);
nor U78 (N_78,In_372,In_222);
nand U79 (N_79,In_45,In_493);
nor U80 (N_80,In_244,In_123);
and U81 (N_81,In_125,In_170);
nor U82 (N_82,In_106,In_42);
or U83 (N_83,In_151,In_317);
and U84 (N_84,In_149,In_450);
nor U85 (N_85,In_153,In_168);
and U86 (N_86,In_194,In_109);
or U87 (N_87,In_411,In_207);
or U88 (N_88,In_54,In_413);
nor U89 (N_89,In_316,In_324);
nor U90 (N_90,In_267,In_352);
nor U91 (N_91,In_201,In_7);
or U92 (N_92,In_470,In_105);
nand U93 (N_93,In_116,In_416);
or U94 (N_94,In_190,In_68);
nand U95 (N_95,In_399,In_171);
nor U96 (N_96,In_325,In_386);
nand U97 (N_97,In_495,In_137);
and U98 (N_98,In_252,In_158);
xnor U99 (N_99,In_274,In_187);
and U100 (N_100,In_258,In_102);
and U101 (N_101,In_288,In_338);
and U102 (N_102,In_50,In_333);
or U103 (N_103,In_211,In_367);
and U104 (N_104,In_331,In_140);
nand U105 (N_105,In_318,In_441);
or U106 (N_106,In_499,In_482);
or U107 (N_107,In_152,In_358);
nor U108 (N_108,In_498,In_199);
and U109 (N_109,In_302,In_421);
nand U110 (N_110,In_447,In_218);
nor U111 (N_111,In_120,In_118);
and U112 (N_112,In_15,In_185);
nand U113 (N_113,In_465,In_11);
or U114 (N_114,In_180,In_249);
nor U115 (N_115,In_296,In_300);
nand U116 (N_116,In_176,In_235);
or U117 (N_117,In_126,In_357);
xnor U118 (N_118,In_245,In_72);
or U119 (N_119,In_277,In_28);
and U120 (N_120,In_99,In_166);
nor U121 (N_121,In_282,In_16);
or U122 (N_122,In_418,In_22);
nand U123 (N_123,In_446,In_295);
nand U124 (N_124,In_474,In_122);
and U125 (N_125,In_273,In_253);
xor U126 (N_126,In_14,In_169);
nand U127 (N_127,In_355,In_494);
xor U128 (N_128,In_80,In_369);
nand U129 (N_129,In_206,In_410);
xnor U130 (N_130,In_88,In_192);
nor U131 (N_131,In_139,In_41);
xor U132 (N_132,In_329,In_256);
or U133 (N_133,In_257,In_488);
or U134 (N_134,In_141,In_213);
nor U135 (N_135,In_32,In_103);
or U136 (N_136,In_284,In_310);
and U137 (N_137,In_359,In_110);
nor U138 (N_138,In_405,In_240);
and U139 (N_139,In_275,In_66);
or U140 (N_140,In_215,In_309);
nand U141 (N_141,In_86,In_286);
nand U142 (N_142,In_336,In_271);
nor U143 (N_143,In_423,In_371);
xnor U144 (N_144,In_483,In_453);
nor U145 (N_145,In_38,In_335);
nor U146 (N_146,In_381,In_379);
or U147 (N_147,In_107,In_280);
nand U148 (N_148,In_342,In_104);
or U149 (N_149,In_154,In_466);
nand U150 (N_150,In_82,In_414);
nand U151 (N_151,In_200,In_129);
nand U152 (N_152,In_276,In_290);
nand U153 (N_153,In_436,In_35);
nor U154 (N_154,In_2,In_311);
and U155 (N_155,In_58,In_219);
xnor U156 (N_156,In_9,In_204);
or U157 (N_157,In_223,In_353);
nand U158 (N_158,In_248,In_402);
and U159 (N_159,In_434,In_186);
and U160 (N_160,In_156,In_127);
nor U161 (N_161,In_65,In_409);
nor U162 (N_162,In_388,In_289);
nor U163 (N_163,In_173,In_283);
and U164 (N_164,In_408,In_36);
xor U165 (N_165,In_243,In_93);
and U166 (N_166,In_326,In_303);
nand U167 (N_167,In_193,In_97);
and U168 (N_168,In_188,In_94);
or U169 (N_169,In_496,In_404);
and U170 (N_170,In_292,In_96);
nor U171 (N_171,In_112,In_396);
and U172 (N_172,In_299,In_10);
nor U173 (N_173,In_269,In_69);
nor U174 (N_174,In_17,In_392);
xnor U175 (N_175,In_332,In_490);
or U176 (N_176,In_113,In_121);
and U177 (N_177,In_469,In_452);
or U178 (N_178,In_376,In_362);
nor U179 (N_179,In_234,In_480);
and U180 (N_180,In_294,In_75);
and U181 (N_181,In_145,In_354);
or U182 (N_182,In_44,In_189);
nand U183 (N_183,In_195,In_4);
nand U184 (N_184,In_214,In_225);
xnor U185 (N_185,In_159,In_26);
or U186 (N_186,In_20,In_301);
or U187 (N_187,In_460,In_417);
nor U188 (N_188,In_91,In_463);
nor U189 (N_189,In_319,In_174);
or U190 (N_190,In_135,In_328);
nor U191 (N_191,In_202,In_224);
and U192 (N_192,In_254,In_320);
nand U193 (N_193,In_343,In_462);
and U194 (N_194,In_432,In_348);
or U195 (N_195,In_391,In_341);
and U196 (N_196,In_393,In_232);
or U197 (N_197,In_178,In_312);
and U198 (N_198,In_37,In_429);
nor U199 (N_199,In_46,In_5);
and U200 (N_200,N_117,N_16);
nand U201 (N_201,N_74,In_131);
nor U202 (N_202,N_50,In_57);
nand U203 (N_203,In_400,In_298);
or U204 (N_204,N_44,N_132);
nand U205 (N_205,In_449,N_109);
or U206 (N_206,In_183,N_49);
nor U207 (N_207,N_147,In_435);
or U208 (N_208,In_19,N_181);
and U209 (N_209,N_70,N_29);
and U210 (N_210,N_173,In_238);
and U211 (N_211,In_382,In_407);
and U212 (N_212,In_356,N_164);
and U213 (N_213,N_183,In_142);
nand U214 (N_214,N_121,N_103);
or U215 (N_215,N_76,N_37);
nand U216 (N_216,In_49,N_139);
nand U217 (N_217,N_38,N_150);
nand U218 (N_218,N_25,In_262);
or U219 (N_219,N_174,N_54);
nor U220 (N_220,N_130,N_72);
nor U221 (N_221,N_186,N_171);
nand U222 (N_222,N_57,N_56);
nor U223 (N_223,In_87,N_39);
and U224 (N_224,N_69,In_62);
nand U225 (N_225,N_125,In_177);
or U226 (N_226,N_152,N_13);
or U227 (N_227,In_231,N_196);
or U228 (N_228,In_161,N_133);
nand U229 (N_229,In_383,In_370);
nand U230 (N_230,N_89,N_3);
nor U231 (N_231,N_94,N_167);
nor U232 (N_232,N_120,In_147);
nor U233 (N_233,N_51,N_151);
or U234 (N_234,N_2,N_82);
nor U235 (N_235,In_39,N_184);
and U236 (N_236,In_291,N_27);
or U237 (N_237,N_159,In_237);
and U238 (N_238,N_185,In_366);
and U239 (N_239,N_144,In_21);
and U240 (N_240,In_360,In_456);
nor U241 (N_241,In_1,In_95);
nor U242 (N_242,N_135,N_178);
nor U243 (N_243,N_46,N_116);
and U244 (N_244,N_84,N_63);
nand U245 (N_245,N_138,N_58);
and U246 (N_246,In_484,N_55);
nor U247 (N_247,N_137,N_21);
and U248 (N_248,In_368,In_81);
nand U249 (N_249,In_403,N_47);
nor U250 (N_250,N_195,In_458);
nand U251 (N_251,In_55,In_305);
nand U252 (N_252,N_110,N_5);
nand U253 (N_253,N_68,N_60);
or U254 (N_254,N_119,N_192);
and U255 (N_255,N_154,In_51);
and U256 (N_256,N_0,N_65);
or U257 (N_257,N_124,N_160);
nor U258 (N_258,In_467,N_31);
nor U259 (N_259,In_179,N_112);
nand U260 (N_260,N_93,In_433);
and U261 (N_261,N_157,N_42);
and U262 (N_262,In_439,N_129);
nand U263 (N_263,In_287,In_364);
and U264 (N_264,N_170,N_26);
nand U265 (N_265,N_142,N_100);
nor U266 (N_266,N_156,In_440);
or U267 (N_267,In_136,N_41);
and U268 (N_268,N_126,N_180);
xnor U269 (N_269,N_87,N_97);
and U270 (N_270,N_88,In_322);
or U271 (N_271,In_182,In_451);
nor U272 (N_272,N_104,N_95);
nand U273 (N_273,In_79,In_8);
and U274 (N_274,N_6,N_23);
nand U275 (N_275,N_66,N_198);
nand U276 (N_276,In_172,In_250);
nor U277 (N_277,N_153,N_80);
xnor U278 (N_278,In_476,N_77);
nand U279 (N_279,In_191,N_14);
nor U280 (N_280,N_115,In_165);
and U281 (N_281,N_179,N_158);
nand U282 (N_282,N_197,N_32);
nand U283 (N_283,N_122,N_92);
nand U284 (N_284,In_24,In_281);
or U285 (N_285,In_25,N_34);
nor U286 (N_286,N_146,In_63);
and U287 (N_287,N_99,N_148);
nor U288 (N_288,In_350,N_165);
nand U289 (N_289,N_24,N_98);
and U290 (N_290,In_216,N_59);
or U291 (N_291,N_83,In_260);
nand U292 (N_292,In_489,N_162);
xor U293 (N_293,N_64,N_71);
or U294 (N_294,In_390,In_92);
nor U295 (N_295,N_176,In_132);
nor U296 (N_296,N_175,In_437);
nand U297 (N_297,N_182,N_101);
xnor U298 (N_298,N_168,N_194);
nor U299 (N_299,N_78,N_189);
and U300 (N_300,In_308,N_199);
nand U301 (N_301,N_166,In_47);
nor U302 (N_302,N_188,In_415);
and U303 (N_303,N_85,In_108);
nand U304 (N_304,In_297,In_76);
and U305 (N_305,N_191,N_33);
nor U306 (N_306,N_163,N_161);
nor U307 (N_307,N_17,N_140);
nor U308 (N_308,N_79,N_19);
nor U309 (N_309,N_86,N_73);
nand U310 (N_310,N_118,N_18);
and U311 (N_311,In_162,N_40);
nor U312 (N_312,In_33,N_1);
and U313 (N_313,N_114,N_190);
xnor U314 (N_314,In_227,N_193);
nand U315 (N_315,In_373,N_187);
and U316 (N_316,N_149,N_62);
nand U317 (N_317,N_30,In_344);
xor U318 (N_318,N_127,N_4);
nor U319 (N_319,N_7,N_134);
and U320 (N_320,N_52,In_101);
or U321 (N_321,N_107,In_83);
or U322 (N_322,N_22,In_148);
nand U323 (N_323,In_30,N_90);
and U324 (N_324,In_205,N_136);
xnor U325 (N_325,N_61,N_9);
or U326 (N_326,N_35,In_398);
or U327 (N_327,N_177,In_304);
and U328 (N_328,N_169,N_91);
nor U329 (N_329,N_102,N_141);
or U330 (N_330,N_131,N_20);
or U331 (N_331,In_346,In_481);
and U332 (N_332,In_337,In_424);
or U333 (N_333,N_48,N_45);
or U334 (N_334,In_111,N_81);
nor U335 (N_335,N_67,N_12);
nor U336 (N_336,In_138,N_123);
nor U337 (N_337,N_10,N_106);
xor U338 (N_338,N_113,N_8);
and U339 (N_339,N_155,In_377);
and U340 (N_340,N_143,N_145);
nand U341 (N_341,N_128,N_15);
nand U342 (N_342,N_96,In_40);
nor U343 (N_343,N_105,N_11);
and U344 (N_344,In_444,N_36);
nand U345 (N_345,N_111,In_150);
or U346 (N_346,N_53,In_457);
or U347 (N_347,N_43,N_108);
xor U348 (N_348,N_172,N_28);
nor U349 (N_349,N_75,In_374);
nor U350 (N_350,In_451,In_87);
nor U351 (N_351,N_69,N_79);
and U352 (N_352,In_366,N_7);
and U353 (N_353,N_186,N_8);
nand U354 (N_354,In_451,N_11);
nand U355 (N_355,In_437,In_382);
and U356 (N_356,In_132,N_48);
nor U357 (N_357,N_154,N_35);
and U358 (N_358,N_149,N_7);
and U359 (N_359,N_174,N_33);
nor U360 (N_360,N_158,N_102);
or U361 (N_361,N_0,In_360);
xnor U362 (N_362,In_476,N_132);
nor U363 (N_363,N_20,In_262);
or U364 (N_364,In_92,In_360);
or U365 (N_365,In_373,N_12);
or U366 (N_366,N_13,N_105);
xor U367 (N_367,N_115,In_33);
or U368 (N_368,In_250,N_7);
or U369 (N_369,In_19,In_403);
and U370 (N_370,N_195,N_157);
nand U371 (N_371,N_29,N_159);
or U372 (N_372,N_40,N_10);
or U373 (N_373,In_403,N_19);
or U374 (N_374,N_72,N_33);
and U375 (N_375,N_161,In_444);
xnor U376 (N_376,N_2,N_39);
or U377 (N_377,N_100,N_140);
or U378 (N_378,In_95,In_360);
or U379 (N_379,N_44,N_178);
or U380 (N_380,N_45,In_62);
or U381 (N_381,N_80,N_72);
nand U382 (N_382,In_322,N_150);
nor U383 (N_383,N_167,N_49);
nor U384 (N_384,N_135,N_2);
or U385 (N_385,N_168,N_91);
nand U386 (N_386,N_26,In_250);
xor U387 (N_387,In_92,N_53);
nand U388 (N_388,N_118,In_30);
and U389 (N_389,N_52,N_36);
and U390 (N_390,N_180,In_138);
and U391 (N_391,N_148,N_16);
nand U392 (N_392,N_196,In_83);
nand U393 (N_393,N_184,In_366);
or U394 (N_394,In_439,N_134);
nand U395 (N_395,N_173,N_35);
nor U396 (N_396,N_30,In_238);
nor U397 (N_397,N_63,N_27);
nor U398 (N_398,N_2,In_132);
nand U399 (N_399,In_398,In_182);
or U400 (N_400,N_319,N_226);
and U401 (N_401,N_353,N_372);
nand U402 (N_402,N_206,N_259);
or U403 (N_403,N_279,N_282);
nand U404 (N_404,N_313,N_263);
nand U405 (N_405,N_257,N_365);
or U406 (N_406,N_342,N_285);
nand U407 (N_407,N_309,N_204);
or U408 (N_408,N_237,N_258);
nand U409 (N_409,N_231,N_228);
or U410 (N_410,N_356,N_205);
or U411 (N_411,N_223,N_300);
and U412 (N_412,N_273,N_201);
and U413 (N_413,N_280,N_227);
and U414 (N_414,N_245,N_334);
and U415 (N_415,N_325,N_304);
or U416 (N_416,N_330,N_307);
nand U417 (N_417,N_338,N_397);
or U418 (N_418,N_302,N_351);
xor U419 (N_419,N_200,N_386);
or U420 (N_420,N_346,N_367);
nor U421 (N_421,N_390,N_350);
and U422 (N_422,N_392,N_221);
nor U423 (N_423,N_389,N_260);
and U424 (N_424,N_222,N_375);
nor U425 (N_425,N_332,N_361);
nor U426 (N_426,N_362,N_208);
nor U427 (N_427,N_381,N_305);
nor U428 (N_428,N_219,N_378);
or U429 (N_429,N_229,N_250);
xnor U430 (N_430,N_268,N_318);
and U431 (N_431,N_331,N_267);
nand U432 (N_432,N_252,N_294);
nor U433 (N_433,N_395,N_271);
nand U434 (N_434,N_391,N_202);
and U435 (N_435,N_303,N_370);
nand U436 (N_436,N_239,N_248);
nand U437 (N_437,N_276,N_398);
nor U438 (N_438,N_242,N_308);
nor U439 (N_439,N_306,N_393);
nand U440 (N_440,N_380,N_217);
or U441 (N_441,N_256,N_265);
and U442 (N_442,N_310,N_246);
nor U443 (N_443,N_377,N_211);
or U444 (N_444,N_321,N_327);
and U445 (N_445,N_274,N_388);
xnor U446 (N_446,N_295,N_328);
nand U447 (N_447,N_266,N_255);
and U448 (N_448,N_337,N_272);
nor U449 (N_449,N_329,N_207);
or U450 (N_450,N_360,N_230);
nor U451 (N_451,N_251,N_264);
and U452 (N_452,N_317,N_335);
nand U453 (N_453,N_296,N_323);
and U454 (N_454,N_312,N_281);
nor U455 (N_455,N_314,N_209);
nor U456 (N_456,N_366,N_254);
or U457 (N_457,N_363,N_345);
nor U458 (N_458,N_286,N_326);
nor U459 (N_459,N_284,N_355);
nor U460 (N_460,N_347,N_243);
nor U461 (N_461,N_357,N_224);
nor U462 (N_462,N_374,N_288);
and U463 (N_463,N_235,N_341);
xor U464 (N_464,N_244,N_299);
and U465 (N_465,N_315,N_262);
and U466 (N_466,N_379,N_348);
nand U467 (N_467,N_311,N_247);
nand U468 (N_468,N_384,N_210);
and U469 (N_469,N_316,N_234);
and U470 (N_470,N_240,N_213);
and U471 (N_471,N_373,N_336);
or U472 (N_472,N_343,N_333);
and U473 (N_473,N_289,N_369);
or U474 (N_474,N_249,N_324);
and U475 (N_475,N_352,N_269);
nor U476 (N_476,N_292,N_368);
nand U477 (N_477,N_349,N_290);
nor U478 (N_478,N_322,N_241);
nand U479 (N_479,N_385,N_253);
or U480 (N_480,N_358,N_382);
or U481 (N_481,N_301,N_359);
nand U482 (N_482,N_399,N_320);
and U483 (N_483,N_236,N_215);
nand U484 (N_484,N_291,N_396);
xor U485 (N_485,N_216,N_277);
xor U486 (N_486,N_283,N_278);
nand U487 (N_487,N_344,N_218);
and U488 (N_488,N_212,N_275);
nand U489 (N_489,N_238,N_214);
or U490 (N_490,N_297,N_203);
xor U491 (N_491,N_354,N_340);
nand U492 (N_492,N_232,N_293);
xnor U493 (N_493,N_383,N_287);
xnor U494 (N_494,N_339,N_376);
and U495 (N_495,N_371,N_225);
or U496 (N_496,N_261,N_394);
nor U497 (N_497,N_387,N_270);
or U498 (N_498,N_364,N_233);
and U499 (N_499,N_220,N_298);
nand U500 (N_500,N_329,N_333);
nor U501 (N_501,N_225,N_379);
or U502 (N_502,N_358,N_252);
or U503 (N_503,N_242,N_377);
or U504 (N_504,N_224,N_275);
and U505 (N_505,N_332,N_313);
and U506 (N_506,N_270,N_233);
nand U507 (N_507,N_353,N_326);
and U508 (N_508,N_269,N_234);
nand U509 (N_509,N_269,N_377);
nor U510 (N_510,N_282,N_383);
nor U511 (N_511,N_301,N_381);
xor U512 (N_512,N_254,N_297);
or U513 (N_513,N_349,N_386);
xnor U514 (N_514,N_292,N_226);
or U515 (N_515,N_367,N_306);
and U516 (N_516,N_341,N_288);
nor U517 (N_517,N_345,N_383);
xor U518 (N_518,N_251,N_316);
nor U519 (N_519,N_383,N_289);
or U520 (N_520,N_252,N_360);
and U521 (N_521,N_242,N_226);
and U522 (N_522,N_331,N_396);
nor U523 (N_523,N_392,N_253);
or U524 (N_524,N_315,N_357);
nand U525 (N_525,N_329,N_212);
or U526 (N_526,N_218,N_203);
nor U527 (N_527,N_341,N_397);
nor U528 (N_528,N_357,N_351);
or U529 (N_529,N_308,N_390);
or U530 (N_530,N_357,N_279);
or U531 (N_531,N_255,N_233);
or U532 (N_532,N_243,N_391);
and U533 (N_533,N_382,N_329);
nand U534 (N_534,N_207,N_246);
and U535 (N_535,N_295,N_263);
and U536 (N_536,N_336,N_355);
nor U537 (N_537,N_381,N_206);
nor U538 (N_538,N_393,N_339);
nor U539 (N_539,N_382,N_222);
or U540 (N_540,N_226,N_328);
nand U541 (N_541,N_216,N_372);
or U542 (N_542,N_335,N_290);
and U543 (N_543,N_279,N_220);
nand U544 (N_544,N_333,N_394);
or U545 (N_545,N_382,N_345);
and U546 (N_546,N_370,N_230);
nand U547 (N_547,N_265,N_396);
nand U548 (N_548,N_251,N_224);
and U549 (N_549,N_379,N_347);
nand U550 (N_550,N_355,N_395);
nand U551 (N_551,N_332,N_394);
nor U552 (N_552,N_352,N_369);
or U553 (N_553,N_356,N_239);
nor U554 (N_554,N_245,N_362);
nor U555 (N_555,N_309,N_222);
nand U556 (N_556,N_380,N_224);
nor U557 (N_557,N_214,N_347);
or U558 (N_558,N_330,N_343);
or U559 (N_559,N_373,N_340);
nor U560 (N_560,N_379,N_262);
nand U561 (N_561,N_375,N_396);
nand U562 (N_562,N_333,N_309);
and U563 (N_563,N_292,N_210);
or U564 (N_564,N_386,N_355);
or U565 (N_565,N_200,N_389);
xor U566 (N_566,N_257,N_260);
and U567 (N_567,N_297,N_260);
nor U568 (N_568,N_283,N_228);
and U569 (N_569,N_292,N_246);
or U570 (N_570,N_208,N_236);
xnor U571 (N_571,N_247,N_331);
or U572 (N_572,N_200,N_339);
or U573 (N_573,N_297,N_277);
or U574 (N_574,N_242,N_200);
nor U575 (N_575,N_234,N_218);
nor U576 (N_576,N_316,N_360);
or U577 (N_577,N_307,N_279);
or U578 (N_578,N_375,N_340);
xnor U579 (N_579,N_311,N_367);
and U580 (N_580,N_244,N_293);
nor U581 (N_581,N_334,N_338);
or U582 (N_582,N_222,N_294);
or U583 (N_583,N_312,N_243);
nor U584 (N_584,N_337,N_308);
nand U585 (N_585,N_269,N_341);
nor U586 (N_586,N_348,N_292);
and U587 (N_587,N_339,N_305);
nor U588 (N_588,N_361,N_281);
nand U589 (N_589,N_293,N_276);
and U590 (N_590,N_273,N_216);
xnor U591 (N_591,N_370,N_382);
xnor U592 (N_592,N_284,N_202);
nor U593 (N_593,N_360,N_314);
nor U594 (N_594,N_363,N_226);
nand U595 (N_595,N_347,N_349);
nand U596 (N_596,N_274,N_203);
or U597 (N_597,N_230,N_300);
nor U598 (N_598,N_288,N_347);
and U599 (N_599,N_213,N_378);
xor U600 (N_600,N_517,N_491);
and U601 (N_601,N_480,N_419);
and U602 (N_602,N_416,N_420);
and U603 (N_603,N_503,N_466);
or U604 (N_604,N_552,N_469);
nor U605 (N_605,N_559,N_405);
or U606 (N_606,N_428,N_429);
nor U607 (N_607,N_477,N_565);
and U608 (N_608,N_571,N_496);
and U609 (N_609,N_561,N_533);
nor U610 (N_610,N_510,N_485);
nand U611 (N_611,N_529,N_579);
or U612 (N_612,N_439,N_442);
nor U613 (N_613,N_551,N_520);
or U614 (N_614,N_583,N_468);
or U615 (N_615,N_563,N_575);
nand U616 (N_616,N_505,N_572);
or U617 (N_617,N_523,N_495);
and U618 (N_618,N_435,N_471);
and U619 (N_619,N_599,N_576);
or U620 (N_620,N_417,N_438);
or U621 (N_621,N_446,N_534);
or U622 (N_622,N_511,N_537);
and U623 (N_623,N_545,N_421);
xnor U624 (N_624,N_492,N_444);
nand U625 (N_625,N_504,N_456);
and U626 (N_626,N_443,N_432);
nand U627 (N_627,N_506,N_573);
or U628 (N_628,N_598,N_596);
and U629 (N_629,N_459,N_554);
or U630 (N_630,N_487,N_555);
and U631 (N_631,N_549,N_461);
nand U632 (N_632,N_586,N_441);
nand U633 (N_633,N_585,N_525);
nor U634 (N_634,N_502,N_424);
nor U635 (N_635,N_472,N_515);
nor U636 (N_636,N_445,N_406);
nand U637 (N_637,N_595,N_548);
or U638 (N_638,N_513,N_589);
or U639 (N_639,N_474,N_423);
nand U640 (N_640,N_518,N_475);
xnor U641 (N_641,N_526,N_498);
nor U642 (N_642,N_581,N_574);
nor U643 (N_643,N_490,N_514);
xnor U644 (N_644,N_591,N_546);
or U645 (N_645,N_519,N_497);
or U646 (N_646,N_566,N_426);
or U647 (N_647,N_412,N_409);
nand U648 (N_648,N_584,N_407);
nand U649 (N_649,N_507,N_422);
and U650 (N_650,N_413,N_531);
nand U651 (N_651,N_535,N_478);
or U652 (N_652,N_536,N_587);
nor U653 (N_653,N_500,N_430);
and U654 (N_654,N_541,N_401);
nand U655 (N_655,N_452,N_489);
nor U656 (N_656,N_481,N_564);
or U657 (N_657,N_493,N_524);
xor U658 (N_658,N_528,N_449);
or U659 (N_659,N_470,N_437);
nand U660 (N_660,N_508,N_450);
nand U661 (N_661,N_453,N_580);
nor U662 (N_662,N_562,N_404);
or U663 (N_663,N_547,N_482);
or U664 (N_664,N_462,N_544);
or U665 (N_665,N_557,N_542);
nor U666 (N_666,N_532,N_556);
nor U667 (N_667,N_577,N_484);
and U668 (N_668,N_558,N_418);
nor U669 (N_669,N_494,N_464);
nand U670 (N_670,N_458,N_516);
and U671 (N_671,N_440,N_451);
and U672 (N_672,N_486,N_415);
nand U673 (N_673,N_593,N_434);
nor U674 (N_674,N_427,N_578);
or U675 (N_675,N_588,N_411);
or U676 (N_676,N_448,N_543);
or U677 (N_677,N_463,N_560);
and U678 (N_678,N_447,N_460);
nand U679 (N_679,N_570,N_592);
nand U680 (N_680,N_509,N_467);
and U681 (N_681,N_569,N_455);
and U682 (N_682,N_410,N_590);
or U683 (N_683,N_499,N_567);
and U684 (N_684,N_476,N_454);
or U685 (N_685,N_521,N_425);
and U686 (N_686,N_479,N_527);
or U687 (N_687,N_550,N_522);
or U688 (N_688,N_433,N_400);
nand U689 (N_689,N_539,N_582);
nor U690 (N_690,N_431,N_553);
nand U691 (N_691,N_473,N_538);
xor U692 (N_692,N_457,N_512);
or U693 (N_693,N_501,N_465);
or U694 (N_694,N_568,N_414);
xnor U695 (N_695,N_408,N_402);
xnor U696 (N_696,N_530,N_488);
or U697 (N_697,N_436,N_597);
and U698 (N_698,N_540,N_594);
and U699 (N_699,N_483,N_403);
nor U700 (N_700,N_594,N_539);
nand U701 (N_701,N_480,N_443);
nand U702 (N_702,N_451,N_522);
or U703 (N_703,N_462,N_568);
nand U704 (N_704,N_431,N_415);
nor U705 (N_705,N_510,N_548);
or U706 (N_706,N_468,N_476);
nand U707 (N_707,N_594,N_479);
nand U708 (N_708,N_409,N_423);
nand U709 (N_709,N_433,N_569);
or U710 (N_710,N_483,N_525);
nand U711 (N_711,N_491,N_512);
or U712 (N_712,N_538,N_503);
nand U713 (N_713,N_533,N_572);
nor U714 (N_714,N_475,N_575);
nand U715 (N_715,N_554,N_467);
and U716 (N_716,N_539,N_435);
nor U717 (N_717,N_410,N_503);
nor U718 (N_718,N_535,N_450);
and U719 (N_719,N_436,N_408);
nand U720 (N_720,N_594,N_549);
or U721 (N_721,N_473,N_403);
or U722 (N_722,N_574,N_595);
nand U723 (N_723,N_572,N_574);
nand U724 (N_724,N_484,N_492);
nor U725 (N_725,N_573,N_428);
nor U726 (N_726,N_536,N_433);
or U727 (N_727,N_464,N_491);
nand U728 (N_728,N_520,N_435);
nor U729 (N_729,N_503,N_579);
and U730 (N_730,N_575,N_495);
or U731 (N_731,N_542,N_548);
and U732 (N_732,N_519,N_554);
nand U733 (N_733,N_446,N_516);
nand U734 (N_734,N_400,N_426);
nor U735 (N_735,N_509,N_533);
or U736 (N_736,N_535,N_479);
nor U737 (N_737,N_452,N_440);
or U738 (N_738,N_476,N_542);
nor U739 (N_739,N_533,N_579);
nor U740 (N_740,N_513,N_539);
or U741 (N_741,N_474,N_421);
and U742 (N_742,N_546,N_421);
or U743 (N_743,N_574,N_435);
nand U744 (N_744,N_417,N_420);
or U745 (N_745,N_459,N_406);
nor U746 (N_746,N_451,N_507);
or U747 (N_747,N_444,N_485);
nand U748 (N_748,N_525,N_534);
and U749 (N_749,N_438,N_510);
nor U750 (N_750,N_458,N_447);
nor U751 (N_751,N_438,N_437);
or U752 (N_752,N_565,N_450);
nor U753 (N_753,N_571,N_478);
or U754 (N_754,N_523,N_533);
xor U755 (N_755,N_510,N_582);
nor U756 (N_756,N_507,N_466);
nor U757 (N_757,N_579,N_520);
or U758 (N_758,N_488,N_468);
nand U759 (N_759,N_490,N_462);
nor U760 (N_760,N_493,N_569);
nand U761 (N_761,N_562,N_402);
or U762 (N_762,N_435,N_467);
xor U763 (N_763,N_541,N_411);
nand U764 (N_764,N_432,N_507);
and U765 (N_765,N_519,N_482);
and U766 (N_766,N_533,N_422);
or U767 (N_767,N_425,N_529);
xor U768 (N_768,N_461,N_440);
nand U769 (N_769,N_426,N_440);
and U770 (N_770,N_523,N_491);
or U771 (N_771,N_501,N_581);
and U772 (N_772,N_445,N_590);
or U773 (N_773,N_556,N_550);
and U774 (N_774,N_463,N_404);
nor U775 (N_775,N_500,N_442);
nor U776 (N_776,N_480,N_524);
xnor U777 (N_777,N_509,N_429);
nor U778 (N_778,N_512,N_549);
and U779 (N_779,N_581,N_520);
nand U780 (N_780,N_510,N_594);
or U781 (N_781,N_411,N_472);
nor U782 (N_782,N_458,N_489);
and U783 (N_783,N_407,N_442);
or U784 (N_784,N_514,N_572);
nor U785 (N_785,N_402,N_531);
and U786 (N_786,N_516,N_515);
nor U787 (N_787,N_465,N_454);
or U788 (N_788,N_576,N_561);
and U789 (N_789,N_572,N_455);
or U790 (N_790,N_501,N_476);
nor U791 (N_791,N_571,N_436);
nand U792 (N_792,N_463,N_442);
or U793 (N_793,N_420,N_487);
nor U794 (N_794,N_557,N_421);
xnor U795 (N_795,N_564,N_580);
or U796 (N_796,N_453,N_594);
and U797 (N_797,N_582,N_450);
or U798 (N_798,N_550,N_412);
or U799 (N_799,N_567,N_463);
or U800 (N_800,N_751,N_617);
xor U801 (N_801,N_671,N_660);
and U802 (N_802,N_661,N_600);
or U803 (N_803,N_710,N_695);
nand U804 (N_804,N_722,N_648);
nor U805 (N_805,N_713,N_606);
and U806 (N_806,N_662,N_707);
nand U807 (N_807,N_618,N_604);
or U808 (N_808,N_761,N_746);
nand U809 (N_809,N_686,N_740);
and U810 (N_810,N_764,N_634);
and U811 (N_811,N_691,N_765);
or U812 (N_812,N_784,N_715);
nand U813 (N_813,N_635,N_666);
and U814 (N_814,N_673,N_745);
nor U815 (N_815,N_766,N_655);
xnor U816 (N_816,N_629,N_681);
and U817 (N_817,N_682,N_690);
nor U818 (N_818,N_756,N_781);
and U819 (N_819,N_731,N_744);
xor U820 (N_820,N_789,N_783);
nand U821 (N_821,N_643,N_770);
and U822 (N_822,N_718,N_675);
or U823 (N_823,N_752,N_650);
and U824 (N_824,N_753,N_657);
or U825 (N_825,N_620,N_637);
nor U826 (N_826,N_772,N_610);
nand U827 (N_827,N_743,N_747);
nor U828 (N_828,N_679,N_796);
and U829 (N_829,N_645,N_795);
nor U830 (N_830,N_644,N_797);
or U831 (N_831,N_669,N_667);
nand U832 (N_832,N_725,N_785);
nand U833 (N_833,N_654,N_638);
or U834 (N_834,N_670,N_723);
nand U835 (N_835,N_627,N_658);
or U836 (N_836,N_632,N_708);
and U837 (N_837,N_641,N_750);
and U838 (N_838,N_714,N_623);
xnor U839 (N_839,N_721,N_678);
xnor U840 (N_840,N_768,N_732);
and U841 (N_841,N_738,N_697);
nor U842 (N_842,N_613,N_776);
nor U843 (N_843,N_664,N_735);
nand U844 (N_844,N_733,N_779);
nor U845 (N_845,N_711,N_626);
nand U846 (N_846,N_622,N_612);
nand U847 (N_847,N_742,N_668);
nand U848 (N_848,N_615,N_773);
nand U849 (N_849,N_692,N_705);
and U850 (N_850,N_663,N_737);
nand U851 (N_851,N_696,N_603);
and U852 (N_852,N_728,N_704);
xnor U853 (N_853,N_611,N_726);
nor U854 (N_854,N_672,N_724);
nand U855 (N_855,N_774,N_631);
xor U856 (N_856,N_685,N_799);
and U857 (N_857,N_702,N_736);
xnor U858 (N_858,N_621,N_601);
and U859 (N_859,N_763,N_607);
nand U860 (N_860,N_748,N_793);
or U861 (N_861,N_769,N_755);
nand U862 (N_862,N_777,N_758);
or U863 (N_863,N_616,N_619);
xnor U864 (N_864,N_754,N_786);
nand U865 (N_865,N_741,N_649);
nand U866 (N_866,N_720,N_739);
nand U867 (N_867,N_633,N_780);
and U868 (N_868,N_647,N_646);
nand U869 (N_869,N_734,N_767);
or U870 (N_870,N_703,N_614);
or U871 (N_871,N_656,N_782);
xor U872 (N_872,N_602,N_677);
or U873 (N_873,N_749,N_693);
or U874 (N_874,N_642,N_636);
nor U875 (N_875,N_630,N_791);
or U876 (N_876,N_730,N_694);
or U877 (N_877,N_688,N_771);
xnor U878 (N_878,N_798,N_700);
or U879 (N_879,N_628,N_699);
nand U880 (N_880,N_717,N_760);
or U881 (N_881,N_729,N_790);
nand U882 (N_882,N_609,N_625);
xor U883 (N_883,N_698,N_687);
nor U884 (N_884,N_762,N_709);
nor U885 (N_885,N_680,N_757);
or U886 (N_886,N_775,N_674);
and U887 (N_887,N_639,N_716);
nor U888 (N_888,N_792,N_653);
or U889 (N_889,N_778,N_706);
nor U890 (N_890,N_787,N_640);
or U891 (N_891,N_759,N_684);
nand U892 (N_892,N_624,N_605);
nor U893 (N_893,N_659,N_719);
and U894 (N_894,N_727,N_652);
and U895 (N_895,N_651,N_794);
nand U896 (N_896,N_689,N_712);
nand U897 (N_897,N_683,N_665);
nor U898 (N_898,N_608,N_788);
or U899 (N_899,N_676,N_701);
nand U900 (N_900,N_675,N_702);
or U901 (N_901,N_742,N_616);
and U902 (N_902,N_606,N_639);
xor U903 (N_903,N_793,N_746);
and U904 (N_904,N_674,N_647);
nand U905 (N_905,N_747,N_631);
or U906 (N_906,N_690,N_639);
and U907 (N_907,N_766,N_711);
nand U908 (N_908,N_616,N_615);
and U909 (N_909,N_633,N_656);
nor U910 (N_910,N_750,N_711);
and U911 (N_911,N_780,N_654);
nand U912 (N_912,N_693,N_625);
or U913 (N_913,N_738,N_768);
nand U914 (N_914,N_685,N_751);
nor U915 (N_915,N_725,N_749);
nand U916 (N_916,N_617,N_640);
and U917 (N_917,N_714,N_703);
xnor U918 (N_918,N_677,N_795);
nor U919 (N_919,N_657,N_602);
xnor U920 (N_920,N_699,N_718);
nand U921 (N_921,N_735,N_663);
nand U922 (N_922,N_681,N_758);
nor U923 (N_923,N_719,N_611);
or U924 (N_924,N_729,N_764);
nor U925 (N_925,N_695,N_730);
nor U926 (N_926,N_638,N_699);
nand U927 (N_927,N_644,N_653);
or U928 (N_928,N_642,N_612);
nor U929 (N_929,N_731,N_630);
and U930 (N_930,N_792,N_741);
nor U931 (N_931,N_666,N_795);
and U932 (N_932,N_725,N_750);
nor U933 (N_933,N_661,N_676);
xnor U934 (N_934,N_676,N_796);
and U935 (N_935,N_732,N_606);
xnor U936 (N_936,N_784,N_738);
nor U937 (N_937,N_703,N_729);
and U938 (N_938,N_705,N_719);
nand U939 (N_939,N_739,N_745);
xnor U940 (N_940,N_661,N_606);
xnor U941 (N_941,N_663,N_747);
nor U942 (N_942,N_747,N_783);
nor U943 (N_943,N_711,N_761);
xnor U944 (N_944,N_738,N_638);
nand U945 (N_945,N_702,N_745);
or U946 (N_946,N_795,N_626);
or U947 (N_947,N_605,N_634);
nand U948 (N_948,N_658,N_623);
or U949 (N_949,N_639,N_685);
nor U950 (N_950,N_706,N_711);
nand U951 (N_951,N_741,N_779);
nand U952 (N_952,N_781,N_761);
and U953 (N_953,N_660,N_715);
nand U954 (N_954,N_769,N_731);
xnor U955 (N_955,N_692,N_674);
xnor U956 (N_956,N_603,N_784);
nand U957 (N_957,N_679,N_741);
and U958 (N_958,N_633,N_629);
xor U959 (N_959,N_635,N_615);
and U960 (N_960,N_719,N_734);
or U961 (N_961,N_704,N_622);
nand U962 (N_962,N_684,N_757);
and U963 (N_963,N_672,N_744);
or U964 (N_964,N_692,N_715);
nand U965 (N_965,N_784,N_653);
or U966 (N_966,N_613,N_646);
and U967 (N_967,N_785,N_792);
nand U968 (N_968,N_614,N_779);
nor U969 (N_969,N_679,N_706);
nor U970 (N_970,N_754,N_675);
nand U971 (N_971,N_765,N_702);
nor U972 (N_972,N_729,N_697);
and U973 (N_973,N_663,N_787);
and U974 (N_974,N_781,N_779);
and U975 (N_975,N_681,N_767);
or U976 (N_976,N_707,N_708);
nand U977 (N_977,N_613,N_667);
or U978 (N_978,N_681,N_733);
nor U979 (N_979,N_759,N_726);
and U980 (N_980,N_776,N_630);
nand U981 (N_981,N_787,N_723);
or U982 (N_982,N_748,N_720);
nor U983 (N_983,N_746,N_628);
and U984 (N_984,N_730,N_645);
xnor U985 (N_985,N_786,N_784);
or U986 (N_986,N_696,N_605);
nor U987 (N_987,N_628,N_772);
or U988 (N_988,N_700,N_661);
and U989 (N_989,N_676,N_624);
or U990 (N_990,N_700,N_744);
xnor U991 (N_991,N_782,N_732);
nand U992 (N_992,N_789,N_714);
nor U993 (N_993,N_601,N_787);
and U994 (N_994,N_603,N_642);
nand U995 (N_995,N_743,N_680);
nand U996 (N_996,N_634,N_712);
or U997 (N_997,N_719,N_741);
nor U998 (N_998,N_649,N_635);
nor U999 (N_999,N_788,N_618);
or U1000 (N_1000,N_958,N_853);
xnor U1001 (N_1001,N_992,N_960);
nor U1002 (N_1002,N_940,N_865);
or U1003 (N_1003,N_860,N_896);
nor U1004 (N_1004,N_912,N_815);
and U1005 (N_1005,N_955,N_988);
or U1006 (N_1006,N_805,N_876);
nor U1007 (N_1007,N_903,N_938);
or U1008 (N_1008,N_852,N_904);
nor U1009 (N_1009,N_870,N_901);
nand U1010 (N_1010,N_924,N_926);
nand U1011 (N_1011,N_922,N_907);
nand U1012 (N_1012,N_919,N_878);
nor U1013 (N_1013,N_918,N_961);
or U1014 (N_1014,N_933,N_847);
and U1015 (N_1015,N_845,N_839);
nor U1016 (N_1016,N_964,N_818);
xnor U1017 (N_1017,N_905,N_858);
and U1018 (N_1018,N_850,N_902);
xor U1019 (N_1019,N_952,N_813);
or U1020 (N_1020,N_976,N_833);
nand U1021 (N_1021,N_829,N_925);
and U1022 (N_1022,N_939,N_898);
nor U1023 (N_1023,N_928,N_911);
nand U1024 (N_1024,N_894,N_801);
nor U1025 (N_1025,N_825,N_835);
nand U1026 (N_1026,N_900,N_956);
and U1027 (N_1027,N_985,N_866);
nor U1028 (N_1028,N_927,N_814);
nand U1029 (N_1029,N_859,N_944);
nand U1030 (N_1030,N_856,N_855);
xor U1031 (N_1031,N_830,N_950);
or U1032 (N_1032,N_920,N_991);
nand U1033 (N_1033,N_846,N_824);
nand U1034 (N_1034,N_862,N_973);
and U1035 (N_1035,N_972,N_947);
or U1036 (N_1036,N_989,N_854);
or U1037 (N_1037,N_808,N_891);
and U1038 (N_1038,N_978,N_826);
or U1039 (N_1039,N_931,N_867);
or U1040 (N_1040,N_809,N_934);
nor U1041 (N_1041,N_914,N_953);
or U1042 (N_1042,N_948,N_857);
and U1043 (N_1043,N_999,N_916);
xnor U1044 (N_1044,N_910,N_849);
or U1045 (N_1045,N_966,N_974);
nor U1046 (N_1046,N_946,N_868);
or U1047 (N_1047,N_828,N_877);
nor U1048 (N_1048,N_832,N_893);
nor U1049 (N_1049,N_831,N_915);
and U1050 (N_1050,N_840,N_864);
and U1051 (N_1051,N_863,N_842);
nor U1052 (N_1052,N_951,N_921);
or U1053 (N_1053,N_879,N_967);
nand U1054 (N_1054,N_886,N_871);
and U1055 (N_1055,N_890,N_937);
nand U1056 (N_1056,N_816,N_923);
nor U1057 (N_1057,N_983,N_959);
nand U1058 (N_1058,N_990,N_980);
nor U1059 (N_1059,N_897,N_930);
xnor U1060 (N_1060,N_848,N_874);
or U1061 (N_1061,N_810,N_889);
or U1062 (N_1062,N_899,N_975);
nor U1063 (N_1063,N_872,N_941);
nand U1064 (N_1064,N_971,N_822);
or U1065 (N_1065,N_885,N_913);
and U1066 (N_1066,N_882,N_819);
xor U1067 (N_1067,N_895,N_800);
nand U1068 (N_1068,N_861,N_883);
nand U1069 (N_1069,N_851,N_837);
nand U1070 (N_1070,N_957,N_977);
nand U1071 (N_1071,N_892,N_984);
or U1072 (N_1072,N_881,N_875);
nand U1073 (N_1073,N_804,N_880);
nor U1074 (N_1074,N_935,N_827);
nand U1075 (N_1075,N_981,N_811);
and U1076 (N_1076,N_993,N_942);
and U1077 (N_1077,N_987,N_841);
or U1078 (N_1078,N_995,N_909);
nor U1079 (N_1079,N_954,N_962);
or U1080 (N_1080,N_807,N_997);
xor U1081 (N_1081,N_986,N_908);
or U1082 (N_1082,N_823,N_982);
xor U1083 (N_1083,N_906,N_844);
nand U1084 (N_1084,N_994,N_888);
and U1085 (N_1085,N_806,N_884);
and U1086 (N_1086,N_817,N_812);
nor U1087 (N_1087,N_873,N_945);
nor U1088 (N_1088,N_803,N_836);
and U1089 (N_1089,N_936,N_821);
nand U1090 (N_1090,N_887,N_949);
nor U1091 (N_1091,N_963,N_834);
nand U1092 (N_1092,N_820,N_996);
nand U1093 (N_1093,N_943,N_843);
nand U1094 (N_1094,N_917,N_969);
or U1095 (N_1095,N_979,N_869);
xor U1096 (N_1096,N_968,N_970);
and U1097 (N_1097,N_932,N_929);
nor U1098 (N_1098,N_802,N_838);
nor U1099 (N_1099,N_998,N_965);
nand U1100 (N_1100,N_854,N_990);
nand U1101 (N_1101,N_932,N_983);
nor U1102 (N_1102,N_884,N_915);
nor U1103 (N_1103,N_958,N_893);
or U1104 (N_1104,N_963,N_927);
and U1105 (N_1105,N_995,N_966);
nand U1106 (N_1106,N_888,N_975);
nor U1107 (N_1107,N_805,N_960);
and U1108 (N_1108,N_939,N_964);
nor U1109 (N_1109,N_814,N_970);
or U1110 (N_1110,N_840,N_959);
nand U1111 (N_1111,N_906,N_950);
xor U1112 (N_1112,N_834,N_850);
nor U1113 (N_1113,N_938,N_842);
nand U1114 (N_1114,N_913,N_841);
nand U1115 (N_1115,N_849,N_936);
nand U1116 (N_1116,N_811,N_990);
nor U1117 (N_1117,N_931,N_823);
xor U1118 (N_1118,N_818,N_960);
nor U1119 (N_1119,N_877,N_847);
nand U1120 (N_1120,N_808,N_961);
and U1121 (N_1121,N_814,N_834);
nor U1122 (N_1122,N_800,N_924);
and U1123 (N_1123,N_940,N_954);
xnor U1124 (N_1124,N_915,N_955);
or U1125 (N_1125,N_953,N_949);
nor U1126 (N_1126,N_981,N_804);
nor U1127 (N_1127,N_836,N_860);
nand U1128 (N_1128,N_825,N_846);
or U1129 (N_1129,N_945,N_875);
and U1130 (N_1130,N_843,N_842);
or U1131 (N_1131,N_802,N_928);
or U1132 (N_1132,N_857,N_903);
nand U1133 (N_1133,N_972,N_915);
nor U1134 (N_1134,N_847,N_972);
nand U1135 (N_1135,N_969,N_970);
xor U1136 (N_1136,N_911,N_932);
nor U1137 (N_1137,N_849,N_901);
xnor U1138 (N_1138,N_883,N_943);
and U1139 (N_1139,N_912,N_906);
and U1140 (N_1140,N_906,N_897);
or U1141 (N_1141,N_925,N_888);
nand U1142 (N_1142,N_893,N_800);
or U1143 (N_1143,N_965,N_882);
nor U1144 (N_1144,N_914,N_885);
nor U1145 (N_1145,N_974,N_997);
and U1146 (N_1146,N_978,N_955);
and U1147 (N_1147,N_980,N_952);
and U1148 (N_1148,N_844,N_884);
or U1149 (N_1149,N_825,N_954);
or U1150 (N_1150,N_929,N_967);
nand U1151 (N_1151,N_997,N_836);
nor U1152 (N_1152,N_917,N_822);
nand U1153 (N_1153,N_932,N_874);
xor U1154 (N_1154,N_936,N_954);
or U1155 (N_1155,N_953,N_975);
nor U1156 (N_1156,N_938,N_822);
nand U1157 (N_1157,N_918,N_805);
nor U1158 (N_1158,N_956,N_809);
nand U1159 (N_1159,N_867,N_833);
or U1160 (N_1160,N_970,N_995);
nand U1161 (N_1161,N_913,N_810);
and U1162 (N_1162,N_843,N_986);
xnor U1163 (N_1163,N_812,N_931);
nand U1164 (N_1164,N_899,N_919);
or U1165 (N_1165,N_988,N_852);
nor U1166 (N_1166,N_886,N_990);
nor U1167 (N_1167,N_827,N_860);
and U1168 (N_1168,N_953,N_933);
or U1169 (N_1169,N_936,N_900);
and U1170 (N_1170,N_947,N_953);
nand U1171 (N_1171,N_904,N_987);
nand U1172 (N_1172,N_812,N_916);
or U1173 (N_1173,N_820,N_978);
or U1174 (N_1174,N_991,N_966);
xnor U1175 (N_1175,N_876,N_859);
and U1176 (N_1176,N_809,N_815);
and U1177 (N_1177,N_862,N_841);
nand U1178 (N_1178,N_855,N_833);
or U1179 (N_1179,N_861,N_999);
nor U1180 (N_1180,N_983,N_878);
or U1181 (N_1181,N_962,N_849);
nor U1182 (N_1182,N_901,N_883);
nor U1183 (N_1183,N_812,N_962);
nand U1184 (N_1184,N_953,N_970);
and U1185 (N_1185,N_855,N_937);
or U1186 (N_1186,N_859,N_884);
nor U1187 (N_1187,N_974,N_898);
or U1188 (N_1188,N_891,N_908);
nand U1189 (N_1189,N_985,N_903);
nand U1190 (N_1190,N_802,N_861);
or U1191 (N_1191,N_995,N_831);
nand U1192 (N_1192,N_920,N_936);
nand U1193 (N_1193,N_822,N_803);
nand U1194 (N_1194,N_956,N_879);
and U1195 (N_1195,N_991,N_883);
nor U1196 (N_1196,N_835,N_860);
or U1197 (N_1197,N_886,N_873);
and U1198 (N_1198,N_880,N_836);
nand U1199 (N_1199,N_938,N_904);
nand U1200 (N_1200,N_1108,N_1060);
nor U1201 (N_1201,N_1094,N_1149);
nor U1202 (N_1202,N_1146,N_1188);
nand U1203 (N_1203,N_1107,N_1101);
or U1204 (N_1204,N_1098,N_1004);
nand U1205 (N_1205,N_1158,N_1033);
nor U1206 (N_1206,N_1115,N_1062);
and U1207 (N_1207,N_1071,N_1134);
nand U1208 (N_1208,N_1017,N_1087);
and U1209 (N_1209,N_1056,N_1170);
or U1210 (N_1210,N_1190,N_1061);
xnor U1211 (N_1211,N_1121,N_1184);
nand U1212 (N_1212,N_1041,N_1103);
or U1213 (N_1213,N_1072,N_1112);
nor U1214 (N_1214,N_1145,N_1142);
and U1215 (N_1215,N_1049,N_1076);
nor U1216 (N_1216,N_1074,N_1147);
and U1217 (N_1217,N_1157,N_1109);
and U1218 (N_1218,N_1036,N_1032);
and U1219 (N_1219,N_1128,N_1009);
or U1220 (N_1220,N_1152,N_1097);
nor U1221 (N_1221,N_1106,N_1192);
and U1222 (N_1222,N_1092,N_1090);
and U1223 (N_1223,N_1059,N_1169);
and U1224 (N_1224,N_1113,N_1163);
nand U1225 (N_1225,N_1085,N_1166);
or U1226 (N_1226,N_1150,N_1114);
or U1227 (N_1227,N_1104,N_1068);
or U1228 (N_1228,N_1116,N_1037);
nand U1229 (N_1229,N_1148,N_1105);
nand U1230 (N_1230,N_1013,N_1005);
nand U1231 (N_1231,N_1155,N_1167);
xor U1232 (N_1232,N_1038,N_1132);
nand U1233 (N_1233,N_1057,N_1137);
nor U1234 (N_1234,N_1077,N_1133);
and U1235 (N_1235,N_1124,N_1173);
and U1236 (N_1236,N_1075,N_1069);
nor U1237 (N_1237,N_1018,N_1034);
or U1238 (N_1238,N_1043,N_1144);
nand U1239 (N_1239,N_1143,N_1099);
nand U1240 (N_1240,N_1138,N_1182);
nand U1241 (N_1241,N_1047,N_1045);
or U1242 (N_1242,N_1187,N_1016);
nor U1243 (N_1243,N_1174,N_1080);
or U1244 (N_1244,N_1102,N_1179);
and U1245 (N_1245,N_1064,N_1010);
nor U1246 (N_1246,N_1088,N_1198);
and U1247 (N_1247,N_1089,N_1176);
nor U1248 (N_1248,N_1154,N_1086);
or U1249 (N_1249,N_1185,N_1175);
and U1250 (N_1250,N_1058,N_1055);
or U1251 (N_1251,N_1189,N_1141);
nor U1252 (N_1252,N_1079,N_1139);
xnor U1253 (N_1253,N_1140,N_1096);
or U1254 (N_1254,N_1180,N_1070);
nor U1255 (N_1255,N_1196,N_1127);
xor U1256 (N_1256,N_1000,N_1122);
xnor U1257 (N_1257,N_1181,N_1031);
nand U1258 (N_1258,N_1199,N_1073);
or U1259 (N_1259,N_1091,N_1156);
and U1260 (N_1260,N_1164,N_1026);
or U1261 (N_1261,N_1151,N_1153);
and U1262 (N_1262,N_1118,N_1131);
nor U1263 (N_1263,N_1135,N_1191);
or U1264 (N_1264,N_1160,N_1052);
xnor U1265 (N_1265,N_1012,N_1020);
nand U1266 (N_1266,N_1029,N_1039);
nand U1267 (N_1267,N_1129,N_1123);
or U1268 (N_1268,N_1007,N_1044);
or U1269 (N_1269,N_1053,N_1014);
or U1270 (N_1270,N_1195,N_1008);
nand U1271 (N_1271,N_1083,N_1050);
nand U1272 (N_1272,N_1065,N_1126);
nand U1273 (N_1273,N_1183,N_1111);
and U1274 (N_1274,N_1125,N_1117);
xor U1275 (N_1275,N_1119,N_1081);
xor U1276 (N_1276,N_1165,N_1023);
and U1277 (N_1277,N_1161,N_1002);
nor U1278 (N_1278,N_1051,N_1120);
and U1279 (N_1279,N_1178,N_1110);
nor U1280 (N_1280,N_1006,N_1027);
or U1281 (N_1281,N_1063,N_1162);
nor U1282 (N_1282,N_1024,N_1003);
or U1283 (N_1283,N_1054,N_1040);
or U1284 (N_1284,N_1130,N_1193);
and U1285 (N_1285,N_1030,N_1177);
xor U1286 (N_1286,N_1028,N_1011);
nand U1287 (N_1287,N_1035,N_1159);
and U1288 (N_1288,N_1001,N_1042);
or U1289 (N_1289,N_1021,N_1048);
and U1290 (N_1290,N_1136,N_1046);
or U1291 (N_1291,N_1025,N_1186);
nor U1292 (N_1292,N_1084,N_1095);
nor U1293 (N_1293,N_1067,N_1015);
or U1294 (N_1294,N_1093,N_1066);
nand U1295 (N_1295,N_1022,N_1197);
and U1296 (N_1296,N_1078,N_1082);
nand U1297 (N_1297,N_1019,N_1172);
nor U1298 (N_1298,N_1168,N_1194);
and U1299 (N_1299,N_1171,N_1100);
nand U1300 (N_1300,N_1005,N_1139);
nand U1301 (N_1301,N_1194,N_1000);
and U1302 (N_1302,N_1187,N_1188);
nand U1303 (N_1303,N_1028,N_1014);
and U1304 (N_1304,N_1093,N_1005);
and U1305 (N_1305,N_1085,N_1094);
nor U1306 (N_1306,N_1163,N_1012);
or U1307 (N_1307,N_1024,N_1186);
or U1308 (N_1308,N_1090,N_1061);
and U1309 (N_1309,N_1138,N_1086);
and U1310 (N_1310,N_1075,N_1157);
nor U1311 (N_1311,N_1169,N_1167);
nand U1312 (N_1312,N_1081,N_1001);
or U1313 (N_1313,N_1041,N_1016);
nor U1314 (N_1314,N_1186,N_1126);
nand U1315 (N_1315,N_1066,N_1004);
xnor U1316 (N_1316,N_1027,N_1192);
nor U1317 (N_1317,N_1183,N_1008);
nor U1318 (N_1318,N_1147,N_1015);
and U1319 (N_1319,N_1178,N_1085);
and U1320 (N_1320,N_1135,N_1114);
or U1321 (N_1321,N_1055,N_1195);
or U1322 (N_1322,N_1101,N_1002);
xnor U1323 (N_1323,N_1114,N_1053);
xnor U1324 (N_1324,N_1108,N_1132);
and U1325 (N_1325,N_1048,N_1057);
or U1326 (N_1326,N_1003,N_1159);
nor U1327 (N_1327,N_1117,N_1112);
or U1328 (N_1328,N_1119,N_1025);
nor U1329 (N_1329,N_1034,N_1138);
xor U1330 (N_1330,N_1104,N_1158);
or U1331 (N_1331,N_1008,N_1022);
nor U1332 (N_1332,N_1191,N_1027);
xor U1333 (N_1333,N_1070,N_1035);
nand U1334 (N_1334,N_1146,N_1055);
or U1335 (N_1335,N_1077,N_1162);
nand U1336 (N_1336,N_1185,N_1027);
nor U1337 (N_1337,N_1090,N_1112);
xnor U1338 (N_1338,N_1110,N_1108);
or U1339 (N_1339,N_1177,N_1106);
and U1340 (N_1340,N_1111,N_1188);
and U1341 (N_1341,N_1187,N_1080);
and U1342 (N_1342,N_1096,N_1156);
nand U1343 (N_1343,N_1127,N_1100);
or U1344 (N_1344,N_1037,N_1100);
nand U1345 (N_1345,N_1085,N_1023);
and U1346 (N_1346,N_1010,N_1050);
nand U1347 (N_1347,N_1082,N_1115);
and U1348 (N_1348,N_1001,N_1103);
and U1349 (N_1349,N_1174,N_1112);
nand U1350 (N_1350,N_1189,N_1171);
nand U1351 (N_1351,N_1045,N_1063);
nand U1352 (N_1352,N_1174,N_1036);
or U1353 (N_1353,N_1065,N_1181);
xor U1354 (N_1354,N_1140,N_1084);
nor U1355 (N_1355,N_1025,N_1154);
and U1356 (N_1356,N_1154,N_1096);
and U1357 (N_1357,N_1061,N_1079);
nand U1358 (N_1358,N_1139,N_1076);
nor U1359 (N_1359,N_1180,N_1102);
and U1360 (N_1360,N_1019,N_1096);
nor U1361 (N_1361,N_1159,N_1192);
and U1362 (N_1362,N_1043,N_1182);
and U1363 (N_1363,N_1008,N_1094);
nand U1364 (N_1364,N_1145,N_1165);
and U1365 (N_1365,N_1186,N_1097);
nor U1366 (N_1366,N_1121,N_1145);
or U1367 (N_1367,N_1000,N_1159);
nand U1368 (N_1368,N_1021,N_1029);
nand U1369 (N_1369,N_1106,N_1112);
and U1370 (N_1370,N_1195,N_1182);
or U1371 (N_1371,N_1055,N_1051);
and U1372 (N_1372,N_1004,N_1193);
or U1373 (N_1373,N_1164,N_1166);
and U1374 (N_1374,N_1009,N_1095);
or U1375 (N_1375,N_1042,N_1194);
nand U1376 (N_1376,N_1014,N_1103);
xnor U1377 (N_1377,N_1156,N_1059);
nand U1378 (N_1378,N_1097,N_1148);
xnor U1379 (N_1379,N_1108,N_1071);
nor U1380 (N_1380,N_1043,N_1154);
or U1381 (N_1381,N_1103,N_1081);
and U1382 (N_1382,N_1092,N_1075);
nor U1383 (N_1383,N_1067,N_1004);
nor U1384 (N_1384,N_1198,N_1117);
nor U1385 (N_1385,N_1098,N_1138);
nand U1386 (N_1386,N_1019,N_1188);
or U1387 (N_1387,N_1007,N_1047);
or U1388 (N_1388,N_1001,N_1031);
nor U1389 (N_1389,N_1119,N_1166);
or U1390 (N_1390,N_1133,N_1007);
nand U1391 (N_1391,N_1121,N_1062);
nor U1392 (N_1392,N_1105,N_1085);
nand U1393 (N_1393,N_1181,N_1122);
or U1394 (N_1394,N_1043,N_1173);
nand U1395 (N_1395,N_1001,N_1010);
and U1396 (N_1396,N_1002,N_1153);
nor U1397 (N_1397,N_1135,N_1082);
or U1398 (N_1398,N_1086,N_1097);
nor U1399 (N_1399,N_1148,N_1132);
and U1400 (N_1400,N_1261,N_1370);
or U1401 (N_1401,N_1234,N_1221);
xnor U1402 (N_1402,N_1229,N_1225);
or U1403 (N_1403,N_1232,N_1351);
or U1404 (N_1404,N_1364,N_1222);
nand U1405 (N_1405,N_1201,N_1392);
nor U1406 (N_1406,N_1327,N_1286);
and U1407 (N_1407,N_1335,N_1242);
xnor U1408 (N_1408,N_1316,N_1211);
or U1409 (N_1409,N_1203,N_1281);
nand U1410 (N_1410,N_1332,N_1302);
nand U1411 (N_1411,N_1226,N_1352);
and U1412 (N_1412,N_1340,N_1207);
or U1413 (N_1413,N_1200,N_1236);
xnor U1414 (N_1414,N_1257,N_1385);
nor U1415 (N_1415,N_1377,N_1224);
xor U1416 (N_1416,N_1235,N_1363);
nor U1417 (N_1417,N_1326,N_1284);
nor U1418 (N_1418,N_1294,N_1379);
nor U1419 (N_1419,N_1338,N_1274);
or U1420 (N_1420,N_1240,N_1321);
or U1421 (N_1421,N_1271,N_1208);
nor U1422 (N_1422,N_1277,N_1381);
nand U1423 (N_1423,N_1398,N_1218);
nor U1424 (N_1424,N_1368,N_1213);
nand U1425 (N_1425,N_1394,N_1375);
nand U1426 (N_1426,N_1355,N_1388);
xor U1427 (N_1427,N_1339,N_1250);
or U1428 (N_1428,N_1353,N_1228);
and U1429 (N_1429,N_1241,N_1373);
nor U1430 (N_1430,N_1356,N_1290);
nand U1431 (N_1431,N_1246,N_1389);
nor U1432 (N_1432,N_1296,N_1273);
nor U1433 (N_1433,N_1251,N_1387);
or U1434 (N_1434,N_1386,N_1308);
nand U1435 (N_1435,N_1249,N_1255);
and U1436 (N_1436,N_1244,N_1365);
and U1437 (N_1437,N_1342,N_1292);
nand U1438 (N_1438,N_1265,N_1333);
nor U1439 (N_1439,N_1260,N_1305);
nor U1440 (N_1440,N_1272,N_1285);
nand U1441 (N_1441,N_1336,N_1259);
or U1442 (N_1442,N_1227,N_1346);
xnor U1443 (N_1443,N_1315,N_1372);
or U1444 (N_1444,N_1202,N_1393);
or U1445 (N_1445,N_1238,N_1350);
xnor U1446 (N_1446,N_1380,N_1237);
nor U1447 (N_1447,N_1312,N_1279);
nand U1448 (N_1448,N_1288,N_1348);
or U1449 (N_1449,N_1344,N_1289);
nor U1450 (N_1450,N_1280,N_1362);
and U1451 (N_1451,N_1253,N_1390);
or U1452 (N_1452,N_1345,N_1205);
and U1453 (N_1453,N_1267,N_1295);
or U1454 (N_1454,N_1310,N_1206);
or U1455 (N_1455,N_1299,N_1269);
nand U1456 (N_1456,N_1215,N_1395);
xnor U1457 (N_1457,N_1314,N_1256);
and U1458 (N_1458,N_1204,N_1254);
or U1459 (N_1459,N_1297,N_1374);
nand U1460 (N_1460,N_1298,N_1307);
nand U1461 (N_1461,N_1396,N_1317);
or U1462 (N_1462,N_1301,N_1270);
or U1463 (N_1463,N_1230,N_1268);
nor U1464 (N_1464,N_1247,N_1354);
nor U1465 (N_1465,N_1369,N_1347);
and U1466 (N_1466,N_1209,N_1233);
and U1467 (N_1467,N_1366,N_1319);
nor U1468 (N_1468,N_1275,N_1282);
nand U1469 (N_1469,N_1266,N_1283);
and U1470 (N_1470,N_1287,N_1349);
xor U1471 (N_1471,N_1384,N_1360);
or U1472 (N_1472,N_1318,N_1313);
nand U1473 (N_1473,N_1276,N_1239);
nor U1474 (N_1474,N_1243,N_1262);
nor U1475 (N_1475,N_1311,N_1293);
nand U1476 (N_1476,N_1359,N_1331);
nor U1477 (N_1477,N_1391,N_1357);
xor U1478 (N_1478,N_1328,N_1343);
nor U1479 (N_1479,N_1397,N_1371);
or U1480 (N_1480,N_1337,N_1214);
and U1481 (N_1481,N_1300,N_1216);
xnor U1482 (N_1482,N_1382,N_1220);
nor U1483 (N_1483,N_1264,N_1219);
nand U1484 (N_1484,N_1330,N_1263);
nor U1485 (N_1485,N_1258,N_1245);
nor U1486 (N_1486,N_1323,N_1217);
or U1487 (N_1487,N_1320,N_1231);
or U1488 (N_1488,N_1252,N_1383);
and U1489 (N_1489,N_1309,N_1291);
and U1490 (N_1490,N_1329,N_1306);
nor U1491 (N_1491,N_1324,N_1358);
nand U1492 (N_1492,N_1367,N_1212);
nor U1493 (N_1493,N_1248,N_1341);
nand U1494 (N_1494,N_1322,N_1223);
xnor U1495 (N_1495,N_1325,N_1361);
nand U1496 (N_1496,N_1376,N_1303);
nor U1497 (N_1497,N_1304,N_1399);
nor U1498 (N_1498,N_1278,N_1378);
nor U1499 (N_1499,N_1334,N_1210);
nand U1500 (N_1500,N_1268,N_1214);
or U1501 (N_1501,N_1299,N_1227);
or U1502 (N_1502,N_1356,N_1372);
xnor U1503 (N_1503,N_1279,N_1244);
and U1504 (N_1504,N_1234,N_1300);
or U1505 (N_1505,N_1232,N_1345);
nand U1506 (N_1506,N_1212,N_1298);
nand U1507 (N_1507,N_1283,N_1377);
nor U1508 (N_1508,N_1342,N_1375);
nor U1509 (N_1509,N_1296,N_1201);
nand U1510 (N_1510,N_1394,N_1312);
and U1511 (N_1511,N_1240,N_1367);
nor U1512 (N_1512,N_1258,N_1247);
xnor U1513 (N_1513,N_1375,N_1340);
and U1514 (N_1514,N_1348,N_1231);
xor U1515 (N_1515,N_1334,N_1360);
or U1516 (N_1516,N_1292,N_1369);
xnor U1517 (N_1517,N_1214,N_1263);
and U1518 (N_1518,N_1270,N_1378);
nand U1519 (N_1519,N_1340,N_1344);
nor U1520 (N_1520,N_1342,N_1321);
nor U1521 (N_1521,N_1388,N_1329);
nand U1522 (N_1522,N_1370,N_1336);
and U1523 (N_1523,N_1206,N_1240);
nor U1524 (N_1524,N_1350,N_1364);
nand U1525 (N_1525,N_1299,N_1265);
nand U1526 (N_1526,N_1211,N_1286);
or U1527 (N_1527,N_1295,N_1283);
nand U1528 (N_1528,N_1223,N_1266);
or U1529 (N_1529,N_1305,N_1327);
nand U1530 (N_1530,N_1243,N_1211);
nand U1531 (N_1531,N_1266,N_1389);
nor U1532 (N_1532,N_1389,N_1302);
nand U1533 (N_1533,N_1317,N_1253);
nor U1534 (N_1534,N_1242,N_1217);
or U1535 (N_1535,N_1258,N_1204);
nor U1536 (N_1536,N_1275,N_1265);
nand U1537 (N_1537,N_1288,N_1290);
nor U1538 (N_1538,N_1265,N_1217);
nand U1539 (N_1539,N_1303,N_1342);
xor U1540 (N_1540,N_1205,N_1369);
nor U1541 (N_1541,N_1220,N_1222);
and U1542 (N_1542,N_1382,N_1366);
or U1543 (N_1543,N_1216,N_1325);
nor U1544 (N_1544,N_1299,N_1258);
and U1545 (N_1545,N_1399,N_1212);
xor U1546 (N_1546,N_1217,N_1384);
nand U1547 (N_1547,N_1252,N_1372);
and U1548 (N_1548,N_1355,N_1335);
and U1549 (N_1549,N_1393,N_1218);
nor U1550 (N_1550,N_1387,N_1304);
nor U1551 (N_1551,N_1313,N_1315);
and U1552 (N_1552,N_1398,N_1239);
nor U1553 (N_1553,N_1320,N_1249);
and U1554 (N_1554,N_1249,N_1289);
and U1555 (N_1555,N_1203,N_1265);
nand U1556 (N_1556,N_1397,N_1201);
xor U1557 (N_1557,N_1312,N_1223);
nor U1558 (N_1558,N_1214,N_1373);
nand U1559 (N_1559,N_1375,N_1356);
xor U1560 (N_1560,N_1274,N_1207);
xor U1561 (N_1561,N_1373,N_1323);
nand U1562 (N_1562,N_1304,N_1274);
or U1563 (N_1563,N_1260,N_1274);
nor U1564 (N_1564,N_1252,N_1231);
or U1565 (N_1565,N_1201,N_1360);
nor U1566 (N_1566,N_1267,N_1224);
nand U1567 (N_1567,N_1253,N_1201);
nor U1568 (N_1568,N_1283,N_1357);
nand U1569 (N_1569,N_1379,N_1305);
nor U1570 (N_1570,N_1361,N_1333);
or U1571 (N_1571,N_1392,N_1216);
nand U1572 (N_1572,N_1317,N_1254);
or U1573 (N_1573,N_1389,N_1254);
and U1574 (N_1574,N_1219,N_1203);
and U1575 (N_1575,N_1264,N_1345);
nand U1576 (N_1576,N_1213,N_1369);
or U1577 (N_1577,N_1390,N_1319);
and U1578 (N_1578,N_1324,N_1263);
and U1579 (N_1579,N_1240,N_1228);
and U1580 (N_1580,N_1281,N_1248);
nand U1581 (N_1581,N_1388,N_1235);
and U1582 (N_1582,N_1341,N_1226);
nand U1583 (N_1583,N_1252,N_1205);
or U1584 (N_1584,N_1216,N_1246);
nand U1585 (N_1585,N_1285,N_1349);
or U1586 (N_1586,N_1363,N_1288);
nand U1587 (N_1587,N_1321,N_1314);
or U1588 (N_1588,N_1203,N_1205);
and U1589 (N_1589,N_1326,N_1384);
nor U1590 (N_1590,N_1346,N_1208);
or U1591 (N_1591,N_1319,N_1396);
xor U1592 (N_1592,N_1309,N_1387);
or U1593 (N_1593,N_1352,N_1278);
nor U1594 (N_1594,N_1389,N_1315);
and U1595 (N_1595,N_1377,N_1227);
and U1596 (N_1596,N_1372,N_1321);
nor U1597 (N_1597,N_1211,N_1235);
or U1598 (N_1598,N_1240,N_1227);
or U1599 (N_1599,N_1358,N_1292);
xor U1600 (N_1600,N_1402,N_1475);
and U1601 (N_1601,N_1472,N_1491);
or U1602 (N_1602,N_1572,N_1576);
or U1603 (N_1603,N_1528,N_1400);
xor U1604 (N_1604,N_1485,N_1506);
and U1605 (N_1605,N_1539,N_1466);
nand U1606 (N_1606,N_1465,N_1579);
or U1607 (N_1607,N_1574,N_1544);
and U1608 (N_1608,N_1449,N_1422);
or U1609 (N_1609,N_1518,N_1487);
nor U1610 (N_1610,N_1540,N_1451);
nand U1611 (N_1611,N_1412,N_1421);
nor U1612 (N_1612,N_1547,N_1503);
and U1613 (N_1613,N_1563,N_1500);
nor U1614 (N_1614,N_1599,N_1470);
and U1615 (N_1615,N_1512,N_1498);
nor U1616 (N_1616,N_1440,N_1510);
and U1617 (N_1617,N_1502,N_1418);
or U1618 (N_1618,N_1549,N_1509);
or U1619 (N_1619,N_1586,N_1480);
or U1620 (N_1620,N_1526,N_1478);
or U1621 (N_1621,N_1474,N_1513);
or U1622 (N_1622,N_1520,N_1592);
or U1623 (N_1623,N_1531,N_1501);
nand U1624 (N_1624,N_1476,N_1593);
nor U1625 (N_1625,N_1555,N_1468);
nand U1626 (N_1626,N_1427,N_1588);
xnor U1627 (N_1627,N_1435,N_1447);
nand U1628 (N_1628,N_1587,N_1515);
or U1629 (N_1629,N_1523,N_1553);
nand U1630 (N_1630,N_1573,N_1493);
or U1631 (N_1631,N_1413,N_1444);
nand U1632 (N_1632,N_1446,N_1471);
nand U1633 (N_1633,N_1445,N_1458);
or U1634 (N_1634,N_1537,N_1557);
nor U1635 (N_1635,N_1562,N_1483);
or U1636 (N_1636,N_1516,N_1519);
nand U1637 (N_1637,N_1495,N_1589);
nor U1638 (N_1638,N_1431,N_1454);
or U1639 (N_1639,N_1443,N_1424);
or U1640 (N_1640,N_1558,N_1482);
and U1641 (N_1641,N_1541,N_1556);
xnor U1642 (N_1642,N_1423,N_1492);
nand U1643 (N_1643,N_1591,N_1479);
nor U1644 (N_1644,N_1517,N_1542);
and U1645 (N_1645,N_1401,N_1559);
nor U1646 (N_1646,N_1404,N_1565);
xor U1647 (N_1647,N_1533,N_1434);
nor U1648 (N_1648,N_1550,N_1554);
nor U1649 (N_1649,N_1429,N_1484);
nand U1650 (N_1650,N_1580,N_1594);
nand U1651 (N_1651,N_1408,N_1436);
or U1652 (N_1652,N_1551,N_1567);
and U1653 (N_1653,N_1499,N_1419);
and U1654 (N_1654,N_1425,N_1530);
and U1655 (N_1655,N_1564,N_1420);
nor U1656 (N_1656,N_1438,N_1538);
nor U1657 (N_1657,N_1463,N_1439);
nand U1658 (N_1658,N_1457,N_1546);
or U1659 (N_1659,N_1494,N_1504);
nor U1660 (N_1660,N_1426,N_1453);
nand U1661 (N_1661,N_1409,N_1570);
or U1662 (N_1662,N_1583,N_1585);
and U1663 (N_1663,N_1543,N_1441);
or U1664 (N_1664,N_1473,N_1469);
nor U1665 (N_1665,N_1522,N_1464);
nor U1666 (N_1666,N_1561,N_1584);
nor U1667 (N_1667,N_1407,N_1581);
nor U1668 (N_1668,N_1486,N_1417);
nand U1669 (N_1669,N_1406,N_1496);
nor U1670 (N_1670,N_1416,N_1582);
or U1671 (N_1671,N_1452,N_1535);
xnor U1672 (N_1672,N_1505,N_1497);
nand U1673 (N_1673,N_1430,N_1460);
and U1674 (N_1674,N_1511,N_1536);
nand U1675 (N_1675,N_1433,N_1590);
nor U1676 (N_1676,N_1477,N_1577);
nand U1677 (N_1677,N_1552,N_1450);
or U1678 (N_1678,N_1405,N_1595);
or U1679 (N_1679,N_1410,N_1403);
nor U1680 (N_1680,N_1432,N_1428);
and U1681 (N_1681,N_1575,N_1507);
and U1682 (N_1682,N_1521,N_1448);
and U1683 (N_1683,N_1437,N_1545);
and U1684 (N_1684,N_1459,N_1442);
nand U1685 (N_1685,N_1560,N_1596);
xor U1686 (N_1686,N_1481,N_1566);
and U1687 (N_1687,N_1490,N_1597);
nand U1688 (N_1688,N_1527,N_1514);
and U1689 (N_1689,N_1524,N_1598);
nor U1690 (N_1690,N_1414,N_1489);
nand U1691 (N_1691,N_1456,N_1534);
nand U1692 (N_1692,N_1411,N_1455);
nor U1693 (N_1693,N_1462,N_1461);
and U1694 (N_1694,N_1568,N_1467);
xnor U1695 (N_1695,N_1529,N_1488);
xor U1696 (N_1696,N_1525,N_1532);
xor U1697 (N_1697,N_1508,N_1571);
and U1698 (N_1698,N_1578,N_1415);
and U1699 (N_1699,N_1548,N_1569);
and U1700 (N_1700,N_1548,N_1438);
nand U1701 (N_1701,N_1406,N_1466);
or U1702 (N_1702,N_1441,N_1570);
nand U1703 (N_1703,N_1426,N_1492);
and U1704 (N_1704,N_1478,N_1540);
xnor U1705 (N_1705,N_1494,N_1539);
nand U1706 (N_1706,N_1563,N_1424);
and U1707 (N_1707,N_1563,N_1505);
nand U1708 (N_1708,N_1490,N_1580);
and U1709 (N_1709,N_1572,N_1565);
or U1710 (N_1710,N_1530,N_1462);
or U1711 (N_1711,N_1509,N_1596);
nor U1712 (N_1712,N_1438,N_1587);
and U1713 (N_1713,N_1574,N_1581);
and U1714 (N_1714,N_1558,N_1471);
nand U1715 (N_1715,N_1467,N_1534);
nor U1716 (N_1716,N_1484,N_1487);
or U1717 (N_1717,N_1464,N_1599);
xnor U1718 (N_1718,N_1463,N_1546);
and U1719 (N_1719,N_1516,N_1402);
xor U1720 (N_1720,N_1544,N_1594);
xor U1721 (N_1721,N_1419,N_1535);
nand U1722 (N_1722,N_1433,N_1475);
or U1723 (N_1723,N_1449,N_1487);
and U1724 (N_1724,N_1409,N_1574);
and U1725 (N_1725,N_1483,N_1413);
nand U1726 (N_1726,N_1532,N_1595);
and U1727 (N_1727,N_1569,N_1419);
xnor U1728 (N_1728,N_1581,N_1512);
nand U1729 (N_1729,N_1586,N_1433);
nand U1730 (N_1730,N_1502,N_1478);
and U1731 (N_1731,N_1565,N_1402);
or U1732 (N_1732,N_1417,N_1427);
nand U1733 (N_1733,N_1403,N_1478);
nor U1734 (N_1734,N_1431,N_1586);
or U1735 (N_1735,N_1577,N_1488);
or U1736 (N_1736,N_1516,N_1542);
nor U1737 (N_1737,N_1490,N_1457);
or U1738 (N_1738,N_1523,N_1458);
nand U1739 (N_1739,N_1441,N_1497);
nor U1740 (N_1740,N_1563,N_1550);
nand U1741 (N_1741,N_1585,N_1560);
and U1742 (N_1742,N_1576,N_1591);
and U1743 (N_1743,N_1421,N_1423);
or U1744 (N_1744,N_1520,N_1435);
and U1745 (N_1745,N_1458,N_1408);
and U1746 (N_1746,N_1515,N_1577);
nor U1747 (N_1747,N_1440,N_1431);
or U1748 (N_1748,N_1488,N_1519);
nand U1749 (N_1749,N_1531,N_1565);
nor U1750 (N_1750,N_1519,N_1413);
and U1751 (N_1751,N_1542,N_1515);
and U1752 (N_1752,N_1594,N_1415);
or U1753 (N_1753,N_1471,N_1429);
nand U1754 (N_1754,N_1558,N_1402);
or U1755 (N_1755,N_1469,N_1572);
nor U1756 (N_1756,N_1564,N_1447);
or U1757 (N_1757,N_1491,N_1452);
nor U1758 (N_1758,N_1504,N_1577);
or U1759 (N_1759,N_1450,N_1480);
and U1760 (N_1760,N_1473,N_1491);
nor U1761 (N_1761,N_1548,N_1533);
nor U1762 (N_1762,N_1530,N_1493);
nand U1763 (N_1763,N_1590,N_1557);
nor U1764 (N_1764,N_1407,N_1592);
nand U1765 (N_1765,N_1410,N_1568);
and U1766 (N_1766,N_1586,N_1424);
or U1767 (N_1767,N_1480,N_1420);
nor U1768 (N_1768,N_1428,N_1430);
or U1769 (N_1769,N_1466,N_1423);
nor U1770 (N_1770,N_1497,N_1405);
and U1771 (N_1771,N_1511,N_1400);
nor U1772 (N_1772,N_1574,N_1439);
xnor U1773 (N_1773,N_1505,N_1579);
and U1774 (N_1774,N_1569,N_1475);
or U1775 (N_1775,N_1444,N_1460);
and U1776 (N_1776,N_1533,N_1403);
nor U1777 (N_1777,N_1439,N_1598);
or U1778 (N_1778,N_1505,N_1465);
nor U1779 (N_1779,N_1424,N_1580);
nor U1780 (N_1780,N_1496,N_1536);
nor U1781 (N_1781,N_1501,N_1556);
and U1782 (N_1782,N_1498,N_1456);
nor U1783 (N_1783,N_1438,N_1509);
nand U1784 (N_1784,N_1445,N_1491);
or U1785 (N_1785,N_1485,N_1582);
and U1786 (N_1786,N_1414,N_1443);
nor U1787 (N_1787,N_1596,N_1583);
xnor U1788 (N_1788,N_1563,N_1569);
and U1789 (N_1789,N_1482,N_1517);
and U1790 (N_1790,N_1487,N_1413);
or U1791 (N_1791,N_1487,N_1573);
nand U1792 (N_1792,N_1558,N_1439);
and U1793 (N_1793,N_1472,N_1495);
nor U1794 (N_1794,N_1559,N_1418);
or U1795 (N_1795,N_1579,N_1412);
or U1796 (N_1796,N_1571,N_1498);
xnor U1797 (N_1797,N_1488,N_1417);
or U1798 (N_1798,N_1430,N_1527);
and U1799 (N_1799,N_1581,N_1551);
and U1800 (N_1800,N_1717,N_1790);
nor U1801 (N_1801,N_1765,N_1629);
xnor U1802 (N_1802,N_1628,N_1627);
and U1803 (N_1803,N_1793,N_1640);
nand U1804 (N_1804,N_1773,N_1604);
or U1805 (N_1805,N_1723,N_1700);
or U1806 (N_1806,N_1608,N_1733);
or U1807 (N_1807,N_1797,N_1669);
nand U1808 (N_1808,N_1743,N_1637);
nor U1809 (N_1809,N_1636,N_1737);
or U1810 (N_1810,N_1692,N_1704);
nand U1811 (N_1811,N_1634,N_1788);
nor U1812 (N_1812,N_1691,N_1665);
and U1813 (N_1813,N_1658,N_1660);
nor U1814 (N_1814,N_1698,N_1772);
nand U1815 (N_1815,N_1792,N_1719);
xnor U1816 (N_1816,N_1656,N_1798);
xor U1817 (N_1817,N_1767,N_1646);
and U1818 (N_1818,N_1664,N_1683);
and U1819 (N_1819,N_1643,N_1710);
nor U1820 (N_1820,N_1757,N_1707);
nor U1821 (N_1821,N_1653,N_1701);
nand U1822 (N_1822,N_1620,N_1672);
xnor U1823 (N_1823,N_1779,N_1739);
nor U1824 (N_1824,N_1766,N_1674);
nor U1825 (N_1825,N_1769,N_1736);
xor U1826 (N_1826,N_1601,N_1771);
xor U1827 (N_1827,N_1730,N_1624);
nor U1828 (N_1828,N_1789,N_1652);
xor U1829 (N_1829,N_1610,N_1679);
and U1830 (N_1830,N_1649,N_1682);
nand U1831 (N_1831,N_1748,N_1661);
nand U1832 (N_1832,N_1638,N_1676);
nor U1833 (N_1833,N_1740,N_1746);
nor U1834 (N_1834,N_1785,N_1729);
and U1835 (N_1835,N_1671,N_1651);
or U1836 (N_1836,N_1712,N_1630);
or U1837 (N_1837,N_1684,N_1603);
and U1838 (N_1838,N_1632,N_1670);
nand U1839 (N_1839,N_1696,N_1657);
xnor U1840 (N_1840,N_1768,N_1741);
or U1841 (N_1841,N_1609,N_1745);
nand U1842 (N_1842,N_1605,N_1787);
or U1843 (N_1843,N_1613,N_1764);
xor U1844 (N_1844,N_1686,N_1612);
xnor U1845 (N_1845,N_1781,N_1715);
nor U1846 (N_1846,N_1731,N_1666);
and U1847 (N_1847,N_1780,N_1687);
and U1848 (N_1848,N_1648,N_1783);
nand U1849 (N_1849,N_1786,N_1694);
nand U1850 (N_1850,N_1626,N_1749);
or U1851 (N_1851,N_1633,N_1776);
nor U1852 (N_1852,N_1728,N_1617);
and U1853 (N_1853,N_1727,N_1706);
nor U1854 (N_1854,N_1752,N_1755);
or U1855 (N_1855,N_1751,N_1725);
xnor U1856 (N_1856,N_1711,N_1759);
nor U1857 (N_1857,N_1796,N_1675);
nor U1858 (N_1858,N_1635,N_1690);
xor U1859 (N_1859,N_1744,N_1721);
and U1860 (N_1860,N_1763,N_1654);
and U1861 (N_1861,N_1750,N_1703);
or U1862 (N_1862,N_1747,N_1623);
or U1863 (N_1863,N_1602,N_1774);
nor U1864 (N_1864,N_1735,N_1647);
nor U1865 (N_1865,N_1784,N_1724);
nor U1866 (N_1866,N_1695,N_1732);
nor U1867 (N_1867,N_1775,N_1689);
nand U1868 (N_1868,N_1734,N_1615);
and U1869 (N_1869,N_1693,N_1625);
nor U1870 (N_1870,N_1645,N_1708);
or U1871 (N_1871,N_1718,N_1697);
or U1872 (N_1872,N_1662,N_1667);
xor U1873 (N_1873,N_1713,N_1606);
and U1874 (N_1874,N_1681,N_1619);
or U1875 (N_1875,N_1795,N_1644);
xnor U1876 (N_1876,N_1611,N_1709);
or U1877 (N_1877,N_1770,N_1756);
nand U1878 (N_1878,N_1663,N_1621);
or U1879 (N_1879,N_1726,N_1673);
or U1880 (N_1880,N_1762,N_1761);
and U1881 (N_1881,N_1631,N_1722);
nor U1882 (N_1882,N_1641,N_1720);
and U1883 (N_1883,N_1782,N_1618);
nand U1884 (N_1884,N_1668,N_1607);
xor U1885 (N_1885,N_1714,N_1680);
nand U1886 (N_1886,N_1753,N_1754);
or U1887 (N_1887,N_1742,N_1614);
nor U1888 (N_1888,N_1622,N_1738);
nand U1889 (N_1889,N_1677,N_1642);
or U1890 (N_1890,N_1705,N_1760);
or U1891 (N_1891,N_1699,N_1794);
nand U1892 (N_1892,N_1702,N_1616);
nor U1893 (N_1893,N_1685,N_1600);
or U1894 (N_1894,N_1639,N_1650);
nor U1895 (N_1895,N_1791,N_1778);
nor U1896 (N_1896,N_1659,N_1678);
or U1897 (N_1897,N_1716,N_1688);
nand U1898 (N_1898,N_1655,N_1777);
or U1899 (N_1899,N_1799,N_1758);
nand U1900 (N_1900,N_1658,N_1690);
nand U1901 (N_1901,N_1761,N_1622);
nor U1902 (N_1902,N_1619,N_1724);
and U1903 (N_1903,N_1795,N_1625);
nand U1904 (N_1904,N_1775,N_1738);
and U1905 (N_1905,N_1680,N_1661);
nor U1906 (N_1906,N_1625,N_1618);
or U1907 (N_1907,N_1762,N_1642);
nor U1908 (N_1908,N_1622,N_1606);
nand U1909 (N_1909,N_1707,N_1697);
and U1910 (N_1910,N_1690,N_1734);
and U1911 (N_1911,N_1752,N_1787);
xnor U1912 (N_1912,N_1661,N_1633);
nand U1913 (N_1913,N_1762,N_1649);
nor U1914 (N_1914,N_1662,N_1612);
nor U1915 (N_1915,N_1622,N_1644);
or U1916 (N_1916,N_1636,N_1703);
or U1917 (N_1917,N_1761,N_1707);
nand U1918 (N_1918,N_1673,N_1759);
and U1919 (N_1919,N_1680,N_1631);
xnor U1920 (N_1920,N_1771,N_1654);
nand U1921 (N_1921,N_1656,N_1601);
or U1922 (N_1922,N_1644,N_1651);
nand U1923 (N_1923,N_1616,N_1667);
nor U1924 (N_1924,N_1627,N_1722);
nand U1925 (N_1925,N_1627,N_1675);
and U1926 (N_1926,N_1688,N_1778);
nand U1927 (N_1927,N_1644,N_1635);
and U1928 (N_1928,N_1678,N_1706);
and U1929 (N_1929,N_1639,N_1741);
and U1930 (N_1930,N_1709,N_1765);
nand U1931 (N_1931,N_1689,N_1603);
nor U1932 (N_1932,N_1740,N_1672);
nand U1933 (N_1933,N_1678,N_1600);
nor U1934 (N_1934,N_1771,N_1625);
nor U1935 (N_1935,N_1655,N_1727);
or U1936 (N_1936,N_1648,N_1771);
nand U1937 (N_1937,N_1793,N_1770);
nor U1938 (N_1938,N_1619,N_1685);
nand U1939 (N_1939,N_1674,N_1750);
nor U1940 (N_1940,N_1609,N_1692);
and U1941 (N_1941,N_1724,N_1606);
and U1942 (N_1942,N_1673,N_1668);
nor U1943 (N_1943,N_1685,N_1672);
nand U1944 (N_1944,N_1782,N_1690);
nand U1945 (N_1945,N_1726,N_1680);
nor U1946 (N_1946,N_1696,N_1751);
xor U1947 (N_1947,N_1782,N_1791);
and U1948 (N_1948,N_1623,N_1657);
nand U1949 (N_1949,N_1646,N_1698);
nor U1950 (N_1950,N_1767,N_1743);
nand U1951 (N_1951,N_1785,N_1606);
nor U1952 (N_1952,N_1629,N_1730);
or U1953 (N_1953,N_1677,N_1766);
or U1954 (N_1954,N_1625,N_1615);
and U1955 (N_1955,N_1744,N_1785);
and U1956 (N_1956,N_1687,N_1608);
and U1957 (N_1957,N_1743,N_1780);
or U1958 (N_1958,N_1608,N_1752);
xnor U1959 (N_1959,N_1657,N_1685);
nand U1960 (N_1960,N_1713,N_1654);
and U1961 (N_1961,N_1794,N_1677);
xnor U1962 (N_1962,N_1626,N_1667);
and U1963 (N_1963,N_1654,N_1720);
nor U1964 (N_1964,N_1711,N_1716);
nor U1965 (N_1965,N_1632,N_1751);
or U1966 (N_1966,N_1649,N_1709);
xnor U1967 (N_1967,N_1706,N_1786);
and U1968 (N_1968,N_1794,N_1766);
nor U1969 (N_1969,N_1630,N_1746);
nand U1970 (N_1970,N_1621,N_1729);
nand U1971 (N_1971,N_1778,N_1755);
or U1972 (N_1972,N_1701,N_1687);
nand U1973 (N_1973,N_1642,N_1615);
nor U1974 (N_1974,N_1792,N_1669);
nand U1975 (N_1975,N_1655,N_1615);
or U1976 (N_1976,N_1777,N_1705);
nor U1977 (N_1977,N_1658,N_1764);
nor U1978 (N_1978,N_1734,N_1640);
or U1979 (N_1979,N_1693,N_1762);
nand U1980 (N_1980,N_1721,N_1627);
nor U1981 (N_1981,N_1626,N_1628);
nand U1982 (N_1982,N_1606,N_1748);
or U1983 (N_1983,N_1736,N_1724);
nor U1984 (N_1984,N_1748,N_1702);
nand U1985 (N_1985,N_1667,N_1635);
or U1986 (N_1986,N_1720,N_1736);
nor U1987 (N_1987,N_1605,N_1708);
or U1988 (N_1988,N_1668,N_1791);
nand U1989 (N_1989,N_1715,N_1639);
nor U1990 (N_1990,N_1756,N_1600);
and U1991 (N_1991,N_1711,N_1792);
or U1992 (N_1992,N_1612,N_1704);
nor U1993 (N_1993,N_1683,N_1794);
nand U1994 (N_1994,N_1660,N_1760);
xor U1995 (N_1995,N_1747,N_1792);
and U1996 (N_1996,N_1668,N_1705);
nor U1997 (N_1997,N_1726,N_1712);
nor U1998 (N_1998,N_1719,N_1671);
xnor U1999 (N_1999,N_1709,N_1767);
or U2000 (N_2000,N_1888,N_1958);
or U2001 (N_2001,N_1815,N_1806);
xnor U2002 (N_2002,N_1994,N_1939);
or U2003 (N_2003,N_1930,N_1973);
and U2004 (N_2004,N_1975,N_1972);
or U2005 (N_2005,N_1970,N_1848);
nor U2006 (N_2006,N_1867,N_1827);
nand U2007 (N_2007,N_1976,N_1928);
and U2008 (N_2008,N_1863,N_1948);
xor U2009 (N_2009,N_1938,N_1922);
nor U2010 (N_2010,N_1864,N_1807);
or U2011 (N_2011,N_1907,N_1802);
nor U2012 (N_2012,N_1974,N_1904);
or U2013 (N_2013,N_1838,N_1847);
nor U2014 (N_2014,N_1971,N_1991);
nor U2015 (N_2015,N_1893,N_1966);
and U2016 (N_2016,N_1917,N_1881);
or U2017 (N_2017,N_1821,N_1862);
nor U2018 (N_2018,N_1990,N_1896);
nor U2019 (N_2019,N_1836,N_1925);
xnor U2020 (N_2020,N_1978,N_1825);
and U2021 (N_2021,N_1983,N_1801);
and U2022 (N_2022,N_1870,N_1872);
xnor U2023 (N_2023,N_1897,N_1859);
and U2024 (N_2024,N_1871,N_1852);
or U2025 (N_2025,N_1915,N_1850);
nor U2026 (N_2026,N_1944,N_1811);
nand U2027 (N_2027,N_1865,N_1860);
or U2028 (N_2028,N_1887,N_1936);
or U2029 (N_2029,N_1968,N_1960);
xor U2030 (N_2030,N_1844,N_1895);
nor U2031 (N_2031,N_1842,N_1841);
xnor U2032 (N_2032,N_1984,N_1998);
nor U2033 (N_2033,N_1942,N_1935);
and U2034 (N_2034,N_1967,N_1992);
nand U2035 (N_2035,N_1800,N_1927);
nor U2036 (N_2036,N_1892,N_1828);
nor U2037 (N_2037,N_1817,N_1949);
nand U2038 (N_2038,N_1876,N_1996);
nand U2039 (N_2039,N_1995,N_1977);
and U2040 (N_2040,N_1875,N_1901);
and U2041 (N_2041,N_1882,N_1869);
xor U2042 (N_2042,N_1814,N_1880);
or U2043 (N_2043,N_1985,N_1906);
and U2044 (N_2044,N_1955,N_1986);
nor U2045 (N_2045,N_1854,N_1809);
nor U2046 (N_2046,N_1961,N_1829);
or U2047 (N_2047,N_1931,N_1954);
nor U2048 (N_2048,N_1858,N_1988);
xor U2049 (N_2049,N_1804,N_1840);
nand U2050 (N_2050,N_1835,N_1959);
xnor U2051 (N_2051,N_1839,N_1818);
and U2052 (N_2052,N_1879,N_1868);
nand U2053 (N_2053,N_1826,N_1919);
nor U2054 (N_2054,N_1980,N_1909);
or U2055 (N_2055,N_1889,N_1857);
and U2056 (N_2056,N_1932,N_1830);
or U2057 (N_2057,N_1957,N_1831);
and U2058 (N_2058,N_1979,N_1834);
nand U2059 (N_2059,N_1902,N_1987);
nand U2060 (N_2060,N_1941,N_1845);
and U2061 (N_2061,N_1920,N_1837);
nor U2062 (N_2062,N_1946,N_1926);
and U2063 (N_2063,N_1823,N_1912);
and U2064 (N_2064,N_1886,N_1894);
xnor U2065 (N_2065,N_1861,N_1933);
and U2066 (N_2066,N_1810,N_1833);
or U2067 (N_2067,N_1947,N_1934);
or U2068 (N_2068,N_1885,N_1808);
or U2069 (N_2069,N_1940,N_1964);
nor U2070 (N_2070,N_1819,N_1999);
nand U2071 (N_2071,N_1898,N_1853);
xor U2072 (N_2072,N_1822,N_1877);
or U2073 (N_2073,N_1911,N_1929);
nor U2074 (N_2074,N_1951,N_1908);
nor U2075 (N_2075,N_1913,N_1916);
and U2076 (N_2076,N_1803,N_1846);
and U2077 (N_2077,N_1855,N_1963);
nand U2078 (N_2078,N_1891,N_1981);
nor U2079 (N_2079,N_1899,N_1965);
xor U2080 (N_2080,N_1878,N_1923);
nor U2081 (N_2081,N_1824,N_1997);
nand U2082 (N_2082,N_1952,N_1937);
or U2083 (N_2083,N_1805,N_1945);
or U2084 (N_2084,N_1890,N_1812);
nor U2085 (N_2085,N_1900,N_1832);
xor U2086 (N_2086,N_1956,N_1813);
nand U2087 (N_2087,N_1918,N_1903);
nand U2088 (N_2088,N_1905,N_1953);
and U2089 (N_2089,N_1884,N_1989);
nor U2090 (N_2090,N_1943,N_1849);
nor U2091 (N_2091,N_1914,N_1921);
or U2092 (N_2092,N_1820,N_1969);
and U2093 (N_2093,N_1816,N_1962);
nor U2094 (N_2094,N_1866,N_1924);
nand U2095 (N_2095,N_1950,N_1982);
or U2096 (N_2096,N_1843,N_1856);
or U2097 (N_2097,N_1874,N_1993);
and U2098 (N_2098,N_1910,N_1851);
nor U2099 (N_2099,N_1883,N_1873);
or U2100 (N_2100,N_1882,N_1831);
nor U2101 (N_2101,N_1832,N_1841);
and U2102 (N_2102,N_1921,N_1837);
nand U2103 (N_2103,N_1949,N_1900);
nor U2104 (N_2104,N_1953,N_1944);
or U2105 (N_2105,N_1925,N_1991);
and U2106 (N_2106,N_1839,N_1938);
xor U2107 (N_2107,N_1909,N_1989);
and U2108 (N_2108,N_1976,N_1989);
or U2109 (N_2109,N_1810,N_1996);
nand U2110 (N_2110,N_1905,N_1874);
nand U2111 (N_2111,N_1862,N_1963);
or U2112 (N_2112,N_1995,N_1896);
nand U2113 (N_2113,N_1872,N_1981);
or U2114 (N_2114,N_1882,N_1824);
nor U2115 (N_2115,N_1860,N_1858);
nor U2116 (N_2116,N_1890,N_1928);
nand U2117 (N_2117,N_1947,N_1820);
and U2118 (N_2118,N_1960,N_1861);
and U2119 (N_2119,N_1883,N_1931);
xnor U2120 (N_2120,N_1824,N_1884);
or U2121 (N_2121,N_1972,N_1860);
or U2122 (N_2122,N_1908,N_1978);
xor U2123 (N_2123,N_1869,N_1816);
xor U2124 (N_2124,N_1872,N_1899);
nor U2125 (N_2125,N_1861,N_1954);
nand U2126 (N_2126,N_1908,N_1817);
or U2127 (N_2127,N_1852,N_1809);
or U2128 (N_2128,N_1804,N_1957);
xnor U2129 (N_2129,N_1996,N_1873);
and U2130 (N_2130,N_1947,N_1823);
nand U2131 (N_2131,N_1947,N_1957);
and U2132 (N_2132,N_1865,N_1974);
nor U2133 (N_2133,N_1827,N_1938);
nor U2134 (N_2134,N_1911,N_1921);
nand U2135 (N_2135,N_1936,N_1819);
nor U2136 (N_2136,N_1859,N_1972);
and U2137 (N_2137,N_1982,N_1885);
xor U2138 (N_2138,N_1963,N_1952);
or U2139 (N_2139,N_1808,N_1867);
and U2140 (N_2140,N_1895,N_1876);
xnor U2141 (N_2141,N_1836,N_1869);
nor U2142 (N_2142,N_1879,N_1836);
and U2143 (N_2143,N_1938,N_1913);
or U2144 (N_2144,N_1908,N_1874);
nand U2145 (N_2145,N_1814,N_1986);
or U2146 (N_2146,N_1969,N_1999);
or U2147 (N_2147,N_1964,N_1896);
and U2148 (N_2148,N_1854,N_1973);
xor U2149 (N_2149,N_1806,N_1945);
or U2150 (N_2150,N_1893,N_1974);
nor U2151 (N_2151,N_1848,N_1934);
nor U2152 (N_2152,N_1900,N_1920);
and U2153 (N_2153,N_1900,N_1956);
or U2154 (N_2154,N_1804,N_1980);
and U2155 (N_2155,N_1959,N_1952);
or U2156 (N_2156,N_1930,N_1825);
and U2157 (N_2157,N_1823,N_1885);
nand U2158 (N_2158,N_1908,N_1967);
or U2159 (N_2159,N_1843,N_1988);
or U2160 (N_2160,N_1954,N_1839);
nand U2161 (N_2161,N_1981,N_1989);
nand U2162 (N_2162,N_1970,N_1872);
or U2163 (N_2163,N_1987,N_1905);
nand U2164 (N_2164,N_1965,N_1936);
xnor U2165 (N_2165,N_1919,N_1968);
and U2166 (N_2166,N_1963,N_1883);
and U2167 (N_2167,N_1962,N_1920);
nand U2168 (N_2168,N_1866,N_1926);
nor U2169 (N_2169,N_1936,N_1996);
and U2170 (N_2170,N_1808,N_1980);
and U2171 (N_2171,N_1976,N_1812);
and U2172 (N_2172,N_1907,N_1997);
nor U2173 (N_2173,N_1810,N_1832);
nand U2174 (N_2174,N_1829,N_1802);
nand U2175 (N_2175,N_1873,N_1886);
or U2176 (N_2176,N_1908,N_1827);
and U2177 (N_2177,N_1835,N_1900);
or U2178 (N_2178,N_1945,N_1950);
nand U2179 (N_2179,N_1932,N_1964);
and U2180 (N_2180,N_1809,N_1965);
or U2181 (N_2181,N_1829,N_1800);
and U2182 (N_2182,N_1856,N_1929);
nand U2183 (N_2183,N_1961,N_1885);
nand U2184 (N_2184,N_1853,N_1854);
and U2185 (N_2185,N_1819,N_1829);
and U2186 (N_2186,N_1850,N_1881);
nor U2187 (N_2187,N_1986,N_1892);
nor U2188 (N_2188,N_1979,N_1959);
nor U2189 (N_2189,N_1820,N_1866);
nand U2190 (N_2190,N_1986,N_1872);
nand U2191 (N_2191,N_1809,N_1900);
or U2192 (N_2192,N_1973,N_1815);
and U2193 (N_2193,N_1854,N_1859);
and U2194 (N_2194,N_1905,N_1811);
nand U2195 (N_2195,N_1986,N_1807);
and U2196 (N_2196,N_1878,N_1807);
nor U2197 (N_2197,N_1983,N_1850);
nor U2198 (N_2198,N_1990,N_1828);
or U2199 (N_2199,N_1865,N_1945);
nand U2200 (N_2200,N_2072,N_2164);
xor U2201 (N_2201,N_2078,N_2048);
nor U2202 (N_2202,N_2087,N_2045);
nor U2203 (N_2203,N_2055,N_2168);
and U2204 (N_2204,N_2059,N_2190);
or U2205 (N_2205,N_2003,N_2046);
and U2206 (N_2206,N_2134,N_2157);
or U2207 (N_2207,N_2101,N_2060);
or U2208 (N_2208,N_2061,N_2135);
nor U2209 (N_2209,N_2155,N_2024);
and U2210 (N_2210,N_2035,N_2083);
nand U2211 (N_2211,N_2097,N_2093);
or U2212 (N_2212,N_2012,N_2033);
nor U2213 (N_2213,N_2032,N_2139);
or U2214 (N_2214,N_2016,N_2014);
and U2215 (N_2215,N_2129,N_2044);
and U2216 (N_2216,N_2007,N_2183);
nor U2217 (N_2217,N_2099,N_2165);
nand U2218 (N_2218,N_2138,N_2023);
and U2219 (N_2219,N_2119,N_2006);
and U2220 (N_2220,N_2043,N_2040);
nor U2221 (N_2221,N_2025,N_2075);
or U2222 (N_2222,N_2166,N_2154);
nand U2223 (N_2223,N_2151,N_2047);
or U2224 (N_2224,N_2123,N_2121);
nor U2225 (N_2225,N_2175,N_2037);
and U2226 (N_2226,N_2140,N_2100);
or U2227 (N_2227,N_2130,N_2098);
nor U2228 (N_2228,N_2053,N_2118);
nor U2229 (N_2229,N_2158,N_2126);
nor U2230 (N_2230,N_2052,N_2115);
xor U2231 (N_2231,N_2018,N_2107);
and U2232 (N_2232,N_2178,N_2149);
or U2233 (N_2233,N_2105,N_2112);
or U2234 (N_2234,N_2030,N_2195);
nand U2235 (N_2235,N_2022,N_2196);
nor U2236 (N_2236,N_2182,N_2077);
or U2237 (N_2237,N_2029,N_2017);
or U2238 (N_2238,N_2049,N_2056);
nor U2239 (N_2239,N_2148,N_2137);
and U2240 (N_2240,N_2125,N_2142);
nor U2241 (N_2241,N_2038,N_2079);
nand U2242 (N_2242,N_2054,N_2092);
nor U2243 (N_2243,N_2095,N_2062);
or U2244 (N_2244,N_2191,N_2069);
nor U2245 (N_2245,N_2192,N_2124);
and U2246 (N_2246,N_2180,N_2013);
nor U2247 (N_2247,N_2171,N_2132);
and U2248 (N_2248,N_2005,N_2074);
or U2249 (N_2249,N_2108,N_2004);
nand U2250 (N_2250,N_2187,N_2064);
nor U2251 (N_2251,N_2010,N_2146);
nand U2252 (N_2252,N_2184,N_2081);
nor U2253 (N_2253,N_2051,N_2021);
or U2254 (N_2254,N_2156,N_2039);
and U2255 (N_2255,N_2117,N_2167);
and U2256 (N_2256,N_2026,N_2084);
or U2257 (N_2257,N_2113,N_2088);
nor U2258 (N_2258,N_2152,N_2194);
nor U2259 (N_2259,N_2094,N_2160);
nor U2260 (N_2260,N_2034,N_2036);
xor U2261 (N_2261,N_2193,N_2080);
or U2262 (N_2262,N_2089,N_2147);
nand U2263 (N_2263,N_2104,N_2001);
nor U2264 (N_2264,N_2188,N_2066);
and U2265 (N_2265,N_2071,N_2106);
or U2266 (N_2266,N_2073,N_2199);
nand U2267 (N_2267,N_2179,N_2086);
and U2268 (N_2268,N_2082,N_2065);
nor U2269 (N_2269,N_2031,N_2145);
nor U2270 (N_2270,N_2186,N_2063);
nand U2271 (N_2271,N_2070,N_2103);
or U2272 (N_2272,N_2120,N_2085);
xor U2273 (N_2273,N_2028,N_2114);
nor U2274 (N_2274,N_2041,N_2111);
and U2275 (N_2275,N_2185,N_2068);
xor U2276 (N_2276,N_2096,N_2131);
or U2277 (N_2277,N_2122,N_2189);
and U2278 (N_2278,N_2136,N_2091);
nand U2279 (N_2279,N_2163,N_2162);
nor U2280 (N_2280,N_2002,N_2177);
nand U2281 (N_2281,N_2116,N_2027);
nor U2282 (N_2282,N_2173,N_2133);
nand U2283 (N_2283,N_2181,N_2019);
and U2284 (N_2284,N_2090,N_2159);
nand U2285 (N_2285,N_2058,N_2008);
nor U2286 (N_2286,N_2076,N_2153);
and U2287 (N_2287,N_2198,N_2197);
nand U2288 (N_2288,N_2011,N_2174);
and U2289 (N_2289,N_2102,N_2161);
and U2290 (N_2290,N_2000,N_2141);
xnor U2291 (N_2291,N_2067,N_2170);
nand U2292 (N_2292,N_2109,N_2172);
or U2293 (N_2293,N_2015,N_2042);
or U2294 (N_2294,N_2143,N_2050);
or U2295 (N_2295,N_2144,N_2110);
and U2296 (N_2296,N_2057,N_2020);
nor U2297 (N_2297,N_2128,N_2150);
and U2298 (N_2298,N_2169,N_2009);
nand U2299 (N_2299,N_2127,N_2176);
or U2300 (N_2300,N_2058,N_2137);
and U2301 (N_2301,N_2048,N_2081);
or U2302 (N_2302,N_2169,N_2187);
or U2303 (N_2303,N_2151,N_2049);
or U2304 (N_2304,N_2172,N_2043);
xor U2305 (N_2305,N_2118,N_2183);
or U2306 (N_2306,N_2014,N_2097);
nand U2307 (N_2307,N_2180,N_2083);
or U2308 (N_2308,N_2016,N_2105);
nand U2309 (N_2309,N_2002,N_2009);
or U2310 (N_2310,N_2095,N_2074);
or U2311 (N_2311,N_2020,N_2000);
and U2312 (N_2312,N_2119,N_2093);
nand U2313 (N_2313,N_2096,N_2042);
nor U2314 (N_2314,N_2184,N_2086);
and U2315 (N_2315,N_2084,N_2122);
or U2316 (N_2316,N_2040,N_2015);
nand U2317 (N_2317,N_2157,N_2080);
and U2318 (N_2318,N_2114,N_2078);
or U2319 (N_2319,N_2177,N_2171);
nor U2320 (N_2320,N_2153,N_2039);
or U2321 (N_2321,N_2096,N_2147);
or U2322 (N_2322,N_2151,N_2079);
and U2323 (N_2323,N_2008,N_2119);
nand U2324 (N_2324,N_2151,N_2137);
or U2325 (N_2325,N_2030,N_2138);
xor U2326 (N_2326,N_2067,N_2150);
and U2327 (N_2327,N_2117,N_2077);
and U2328 (N_2328,N_2040,N_2116);
or U2329 (N_2329,N_2189,N_2039);
nand U2330 (N_2330,N_2111,N_2156);
nor U2331 (N_2331,N_2076,N_2027);
and U2332 (N_2332,N_2164,N_2187);
nor U2333 (N_2333,N_2178,N_2193);
nor U2334 (N_2334,N_2138,N_2086);
xor U2335 (N_2335,N_2097,N_2178);
nor U2336 (N_2336,N_2066,N_2012);
nand U2337 (N_2337,N_2152,N_2089);
or U2338 (N_2338,N_2108,N_2185);
nand U2339 (N_2339,N_2129,N_2080);
xor U2340 (N_2340,N_2107,N_2051);
nor U2341 (N_2341,N_2177,N_2036);
or U2342 (N_2342,N_2110,N_2012);
or U2343 (N_2343,N_2152,N_2049);
nand U2344 (N_2344,N_2047,N_2087);
nand U2345 (N_2345,N_2086,N_2115);
and U2346 (N_2346,N_2094,N_2198);
and U2347 (N_2347,N_2134,N_2176);
nand U2348 (N_2348,N_2133,N_2050);
or U2349 (N_2349,N_2130,N_2165);
nor U2350 (N_2350,N_2154,N_2025);
nand U2351 (N_2351,N_2075,N_2003);
nor U2352 (N_2352,N_2161,N_2104);
nand U2353 (N_2353,N_2065,N_2161);
xnor U2354 (N_2354,N_2093,N_2179);
nand U2355 (N_2355,N_2083,N_2025);
xnor U2356 (N_2356,N_2177,N_2197);
xnor U2357 (N_2357,N_2162,N_2146);
and U2358 (N_2358,N_2150,N_2197);
nor U2359 (N_2359,N_2161,N_2019);
and U2360 (N_2360,N_2048,N_2199);
or U2361 (N_2361,N_2051,N_2140);
xor U2362 (N_2362,N_2141,N_2124);
nor U2363 (N_2363,N_2105,N_2117);
and U2364 (N_2364,N_2057,N_2041);
or U2365 (N_2365,N_2041,N_2141);
nand U2366 (N_2366,N_2152,N_2016);
nand U2367 (N_2367,N_2155,N_2005);
nor U2368 (N_2368,N_2081,N_2031);
nand U2369 (N_2369,N_2166,N_2059);
and U2370 (N_2370,N_2156,N_2069);
xor U2371 (N_2371,N_2037,N_2040);
nor U2372 (N_2372,N_2046,N_2189);
nor U2373 (N_2373,N_2182,N_2116);
nand U2374 (N_2374,N_2172,N_2091);
or U2375 (N_2375,N_2137,N_2192);
nand U2376 (N_2376,N_2116,N_2043);
nand U2377 (N_2377,N_2141,N_2177);
or U2378 (N_2378,N_2098,N_2131);
nor U2379 (N_2379,N_2185,N_2060);
and U2380 (N_2380,N_2108,N_2161);
xor U2381 (N_2381,N_2177,N_2040);
xnor U2382 (N_2382,N_2136,N_2172);
or U2383 (N_2383,N_2026,N_2024);
and U2384 (N_2384,N_2169,N_2129);
and U2385 (N_2385,N_2138,N_2085);
or U2386 (N_2386,N_2128,N_2156);
nor U2387 (N_2387,N_2023,N_2142);
and U2388 (N_2388,N_2144,N_2132);
nand U2389 (N_2389,N_2114,N_2071);
nand U2390 (N_2390,N_2021,N_2110);
nand U2391 (N_2391,N_2087,N_2145);
nand U2392 (N_2392,N_2107,N_2113);
or U2393 (N_2393,N_2132,N_2136);
or U2394 (N_2394,N_2130,N_2007);
and U2395 (N_2395,N_2030,N_2191);
nor U2396 (N_2396,N_2149,N_2167);
nand U2397 (N_2397,N_2198,N_2117);
nand U2398 (N_2398,N_2049,N_2053);
nor U2399 (N_2399,N_2105,N_2059);
nand U2400 (N_2400,N_2379,N_2249);
and U2401 (N_2401,N_2342,N_2390);
xor U2402 (N_2402,N_2202,N_2252);
nand U2403 (N_2403,N_2224,N_2303);
nand U2404 (N_2404,N_2346,N_2354);
or U2405 (N_2405,N_2326,N_2276);
xor U2406 (N_2406,N_2348,N_2353);
or U2407 (N_2407,N_2371,N_2318);
or U2408 (N_2408,N_2228,N_2360);
or U2409 (N_2409,N_2344,N_2349);
or U2410 (N_2410,N_2278,N_2361);
nor U2411 (N_2411,N_2381,N_2279);
nor U2412 (N_2412,N_2386,N_2334);
and U2413 (N_2413,N_2359,N_2241);
nand U2414 (N_2414,N_2367,N_2218);
xnor U2415 (N_2415,N_2294,N_2337);
and U2416 (N_2416,N_2319,N_2331);
nor U2417 (N_2417,N_2213,N_2216);
nor U2418 (N_2418,N_2247,N_2292);
nor U2419 (N_2419,N_2270,N_2350);
nand U2420 (N_2420,N_2338,N_2383);
or U2421 (N_2421,N_2320,N_2322);
xnor U2422 (N_2422,N_2255,N_2280);
nor U2423 (N_2423,N_2340,N_2323);
nand U2424 (N_2424,N_2201,N_2351);
and U2425 (N_2425,N_2356,N_2394);
xnor U2426 (N_2426,N_2261,N_2208);
nor U2427 (N_2427,N_2329,N_2358);
nand U2428 (N_2428,N_2253,N_2288);
or U2429 (N_2429,N_2328,N_2364);
nor U2430 (N_2430,N_2231,N_2388);
and U2431 (N_2431,N_2306,N_2372);
nand U2432 (N_2432,N_2374,N_2248);
or U2433 (N_2433,N_2312,N_2399);
nor U2434 (N_2434,N_2225,N_2263);
and U2435 (N_2435,N_2352,N_2309);
and U2436 (N_2436,N_2339,N_2244);
and U2437 (N_2437,N_2265,N_2389);
and U2438 (N_2438,N_2363,N_2254);
or U2439 (N_2439,N_2211,N_2365);
and U2440 (N_2440,N_2203,N_2223);
nand U2441 (N_2441,N_2215,N_2221);
nand U2442 (N_2442,N_2251,N_2264);
or U2443 (N_2443,N_2267,N_2219);
and U2444 (N_2444,N_2395,N_2283);
nand U2445 (N_2445,N_2384,N_2233);
or U2446 (N_2446,N_2281,N_2305);
or U2447 (N_2447,N_2355,N_2207);
and U2448 (N_2448,N_2277,N_2236);
and U2449 (N_2449,N_2327,N_2396);
xnor U2450 (N_2450,N_2273,N_2290);
nand U2451 (N_2451,N_2313,N_2333);
nand U2452 (N_2452,N_2378,N_2234);
xnor U2453 (N_2453,N_2245,N_2298);
or U2454 (N_2454,N_2256,N_2391);
and U2455 (N_2455,N_2382,N_2209);
nand U2456 (N_2456,N_2239,N_2226);
or U2457 (N_2457,N_2242,N_2250);
nor U2458 (N_2458,N_2302,N_2325);
and U2459 (N_2459,N_2398,N_2291);
or U2460 (N_2460,N_2299,N_2377);
or U2461 (N_2461,N_2336,N_2205);
nor U2462 (N_2462,N_2300,N_2343);
and U2463 (N_2463,N_2341,N_2200);
nand U2464 (N_2464,N_2235,N_2269);
nand U2465 (N_2465,N_2321,N_2227);
nor U2466 (N_2466,N_2232,N_2308);
xnor U2467 (N_2467,N_2284,N_2266);
nor U2468 (N_2468,N_2380,N_2316);
nor U2469 (N_2469,N_2373,N_2307);
nand U2470 (N_2470,N_2257,N_2237);
nor U2471 (N_2471,N_2315,N_2230);
or U2472 (N_2472,N_2397,N_2393);
or U2473 (N_2473,N_2330,N_2376);
nor U2474 (N_2474,N_2310,N_2220);
and U2475 (N_2475,N_2287,N_2275);
or U2476 (N_2476,N_2304,N_2296);
xnor U2477 (N_2477,N_2282,N_2272);
nor U2478 (N_2478,N_2262,N_2314);
nand U2479 (N_2479,N_2240,N_2259);
and U2480 (N_2480,N_2246,N_2229);
or U2481 (N_2481,N_2295,N_2274);
and U2482 (N_2482,N_2332,N_2210);
or U2483 (N_2483,N_2214,N_2238);
or U2484 (N_2484,N_2335,N_2293);
nor U2485 (N_2485,N_2345,N_2347);
or U2486 (N_2486,N_2222,N_2243);
or U2487 (N_2487,N_2286,N_2271);
or U2488 (N_2488,N_2357,N_2392);
or U2489 (N_2489,N_2370,N_2212);
and U2490 (N_2490,N_2260,N_2285);
and U2491 (N_2491,N_2375,N_2301);
and U2492 (N_2492,N_2362,N_2311);
nor U2493 (N_2493,N_2366,N_2258);
nor U2494 (N_2494,N_2217,N_2268);
nand U2495 (N_2495,N_2297,N_2368);
xnor U2496 (N_2496,N_2324,N_2385);
and U2497 (N_2497,N_2204,N_2369);
nor U2498 (N_2498,N_2317,N_2289);
or U2499 (N_2499,N_2387,N_2206);
and U2500 (N_2500,N_2256,N_2243);
and U2501 (N_2501,N_2240,N_2235);
nor U2502 (N_2502,N_2356,N_2214);
nor U2503 (N_2503,N_2226,N_2298);
nor U2504 (N_2504,N_2329,N_2328);
nand U2505 (N_2505,N_2335,N_2301);
or U2506 (N_2506,N_2248,N_2251);
xor U2507 (N_2507,N_2212,N_2247);
nor U2508 (N_2508,N_2376,N_2241);
and U2509 (N_2509,N_2334,N_2273);
nor U2510 (N_2510,N_2255,N_2337);
nand U2511 (N_2511,N_2286,N_2230);
or U2512 (N_2512,N_2338,N_2297);
nand U2513 (N_2513,N_2230,N_2225);
nand U2514 (N_2514,N_2300,N_2358);
or U2515 (N_2515,N_2348,N_2366);
and U2516 (N_2516,N_2237,N_2328);
and U2517 (N_2517,N_2261,N_2315);
or U2518 (N_2518,N_2339,N_2340);
nor U2519 (N_2519,N_2361,N_2240);
nand U2520 (N_2520,N_2381,N_2320);
nor U2521 (N_2521,N_2267,N_2361);
or U2522 (N_2522,N_2385,N_2299);
or U2523 (N_2523,N_2384,N_2364);
and U2524 (N_2524,N_2333,N_2212);
and U2525 (N_2525,N_2220,N_2382);
or U2526 (N_2526,N_2209,N_2393);
or U2527 (N_2527,N_2225,N_2376);
nand U2528 (N_2528,N_2212,N_2223);
or U2529 (N_2529,N_2233,N_2362);
nand U2530 (N_2530,N_2319,N_2340);
and U2531 (N_2531,N_2379,N_2377);
nand U2532 (N_2532,N_2270,N_2231);
and U2533 (N_2533,N_2319,N_2318);
nor U2534 (N_2534,N_2200,N_2330);
and U2535 (N_2535,N_2288,N_2380);
or U2536 (N_2536,N_2377,N_2338);
and U2537 (N_2537,N_2204,N_2357);
nor U2538 (N_2538,N_2333,N_2339);
or U2539 (N_2539,N_2212,N_2368);
or U2540 (N_2540,N_2223,N_2317);
and U2541 (N_2541,N_2303,N_2248);
nand U2542 (N_2542,N_2311,N_2276);
and U2543 (N_2543,N_2260,N_2366);
xor U2544 (N_2544,N_2348,N_2293);
nand U2545 (N_2545,N_2252,N_2249);
nand U2546 (N_2546,N_2362,N_2235);
nand U2547 (N_2547,N_2383,N_2369);
nor U2548 (N_2548,N_2242,N_2397);
nand U2549 (N_2549,N_2295,N_2324);
or U2550 (N_2550,N_2247,N_2233);
xor U2551 (N_2551,N_2365,N_2253);
and U2552 (N_2552,N_2396,N_2374);
nor U2553 (N_2553,N_2363,N_2339);
or U2554 (N_2554,N_2303,N_2384);
and U2555 (N_2555,N_2249,N_2260);
xnor U2556 (N_2556,N_2357,N_2274);
nand U2557 (N_2557,N_2282,N_2277);
nand U2558 (N_2558,N_2279,N_2281);
and U2559 (N_2559,N_2262,N_2343);
and U2560 (N_2560,N_2252,N_2268);
or U2561 (N_2561,N_2278,N_2280);
and U2562 (N_2562,N_2253,N_2370);
xnor U2563 (N_2563,N_2334,N_2323);
nor U2564 (N_2564,N_2286,N_2394);
or U2565 (N_2565,N_2216,N_2315);
and U2566 (N_2566,N_2294,N_2216);
xor U2567 (N_2567,N_2330,N_2363);
nor U2568 (N_2568,N_2290,N_2231);
nand U2569 (N_2569,N_2214,N_2300);
and U2570 (N_2570,N_2281,N_2367);
nand U2571 (N_2571,N_2297,N_2273);
nor U2572 (N_2572,N_2310,N_2363);
or U2573 (N_2573,N_2303,N_2337);
and U2574 (N_2574,N_2247,N_2224);
nor U2575 (N_2575,N_2276,N_2229);
nor U2576 (N_2576,N_2373,N_2388);
nor U2577 (N_2577,N_2238,N_2311);
xor U2578 (N_2578,N_2378,N_2398);
nand U2579 (N_2579,N_2335,N_2267);
nor U2580 (N_2580,N_2382,N_2369);
or U2581 (N_2581,N_2363,N_2271);
nor U2582 (N_2582,N_2307,N_2332);
or U2583 (N_2583,N_2314,N_2293);
or U2584 (N_2584,N_2213,N_2341);
and U2585 (N_2585,N_2304,N_2323);
nor U2586 (N_2586,N_2262,N_2395);
or U2587 (N_2587,N_2210,N_2364);
or U2588 (N_2588,N_2301,N_2222);
nand U2589 (N_2589,N_2214,N_2297);
nor U2590 (N_2590,N_2212,N_2350);
nor U2591 (N_2591,N_2329,N_2386);
or U2592 (N_2592,N_2213,N_2353);
or U2593 (N_2593,N_2335,N_2325);
nor U2594 (N_2594,N_2254,N_2289);
or U2595 (N_2595,N_2372,N_2381);
and U2596 (N_2596,N_2354,N_2221);
nand U2597 (N_2597,N_2362,N_2274);
nor U2598 (N_2598,N_2391,N_2228);
nand U2599 (N_2599,N_2289,N_2311);
nand U2600 (N_2600,N_2549,N_2500);
or U2601 (N_2601,N_2458,N_2497);
nor U2602 (N_2602,N_2423,N_2416);
nor U2603 (N_2603,N_2566,N_2495);
nand U2604 (N_2604,N_2578,N_2511);
or U2605 (N_2605,N_2457,N_2563);
or U2606 (N_2606,N_2502,N_2471);
nor U2607 (N_2607,N_2463,N_2545);
or U2608 (N_2608,N_2547,N_2521);
or U2609 (N_2609,N_2572,N_2482);
or U2610 (N_2610,N_2498,N_2470);
nand U2611 (N_2611,N_2591,N_2474);
or U2612 (N_2612,N_2577,N_2571);
xor U2613 (N_2613,N_2408,N_2592);
and U2614 (N_2614,N_2433,N_2524);
or U2615 (N_2615,N_2435,N_2558);
or U2616 (N_2616,N_2476,N_2442);
and U2617 (N_2617,N_2402,N_2503);
nand U2618 (N_2618,N_2553,N_2430);
nand U2619 (N_2619,N_2425,N_2538);
or U2620 (N_2620,N_2598,N_2445);
or U2621 (N_2621,N_2462,N_2515);
and U2622 (N_2622,N_2585,N_2443);
or U2623 (N_2623,N_2493,N_2528);
nand U2624 (N_2624,N_2459,N_2552);
and U2625 (N_2625,N_2599,N_2542);
nor U2626 (N_2626,N_2472,N_2436);
nand U2627 (N_2627,N_2478,N_2514);
nor U2628 (N_2628,N_2557,N_2569);
nand U2629 (N_2629,N_2450,N_2505);
or U2630 (N_2630,N_2589,N_2525);
and U2631 (N_2631,N_2492,N_2507);
nand U2632 (N_2632,N_2584,N_2449);
xnor U2633 (N_2633,N_2579,N_2551);
nand U2634 (N_2634,N_2526,N_2586);
or U2635 (N_2635,N_2484,N_2481);
and U2636 (N_2636,N_2483,N_2581);
and U2637 (N_2637,N_2494,N_2401);
or U2638 (N_2638,N_2570,N_2565);
nand U2639 (N_2639,N_2509,N_2460);
nor U2640 (N_2640,N_2439,N_2582);
and U2641 (N_2641,N_2455,N_2420);
and U2642 (N_2642,N_2466,N_2480);
nor U2643 (N_2643,N_2597,N_2554);
nand U2644 (N_2644,N_2588,N_2533);
nand U2645 (N_2645,N_2534,N_2537);
nor U2646 (N_2646,N_2539,N_2441);
or U2647 (N_2647,N_2501,N_2594);
nor U2648 (N_2648,N_2556,N_2574);
nor U2649 (N_2649,N_2590,N_2475);
nand U2650 (N_2650,N_2550,N_2488);
and U2651 (N_2651,N_2432,N_2535);
nor U2652 (N_2652,N_2527,N_2587);
nor U2653 (N_2653,N_2520,N_2448);
nand U2654 (N_2654,N_2409,N_2583);
or U2655 (N_2655,N_2499,N_2504);
or U2656 (N_2656,N_2548,N_2469);
nand U2657 (N_2657,N_2485,N_2529);
or U2658 (N_2658,N_2513,N_2519);
and U2659 (N_2659,N_2424,N_2446);
or U2660 (N_2660,N_2516,N_2560);
nor U2661 (N_2661,N_2422,N_2555);
or U2662 (N_2662,N_2438,N_2486);
or U2663 (N_2663,N_2400,N_2532);
xor U2664 (N_2664,N_2530,N_2540);
nand U2665 (N_2665,N_2543,N_2465);
or U2666 (N_2666,N_2419,N_2447);
and U2667 (N_2667,N_2580,N_2575);
xnor U2668 (N_2668,N_2406,N_2414);
nand U2669 (N_2669,N_2451,N_2421);
nand U2670 (N_2670,N_2541,N_2489);
nand U2671 (N_2671,N_2437,N_2576);
nand U2672 (N_2672,N_2567,N_2561);
and U2673 (N_2673,N_2407,N_2413);
nor U2674 (N_2674,N_2536,N_2454);
nand U2675 (N_2675,N_2440,N_2434);
nor U2676 (N_2676,N_2523,N_2559);
or U2677 (N_2677,N_2467,N_2428);
and U2678 (N_2678,N_2405,N_2477);
nand U2679 (N_2679,N_2453,N_2456);
and U2680 (N_2680,N_2411,N_2444);
and U2681 (N_2681,N_2418,N_2452);
and U2682 (N_2682,N_2487,N_2544);
or U2683 (N_2683,N_2490,N_2568);
or U2684 (N_2684,N_2415,N_2496);
xor U2685 (N_2685,N_2508,N_2417);
and U2686 (N_2686,N_2595,N_2512);
nand U2687 (N_2687,N_2573,N_2426);
nor U2688 (N_2688,N_2412,N_2593);
and U2689 (N_2689,N_2429,N_2427);
nand U2690 (N_2690,N_2562,N_2473);
or U2691 (N_2691,N_2518,N_2522);
nor U2692 (N_2692,N_2506,N_2403);
nand U2693 (N_2693,N_2531,N_2517);
nand U2694 (N_2694,N_2510,N_2461);
nor U2695 (N_2695,N_2564,N_2546);
nand U2696 (N_2696,N_2431,N_2479);
nand U2697 (N_2697,N_2491,N_2468);
or U2698 (N_2698,N_2596,N_2410);
and U2699 (N_2699,N_2404,N_2464);
xor U2700 (N_2700,N_2495,N_2545);
xnor U2701 (N_2701,N_2569,N_2550);
and U2702 (N_2702,N_2469,N_2513);
nand U2703 (N_2703,N_2558,N_2458);
or U2704 (N_2704,N_2526,N_2593);
or U2705 (N_2705,N_2549,N_2522);
and U2706 (N_2706,N_2451,N_2543);
nor U2707 (N_2707,N_2502,N_2551);
or U2708 (N_2708,N_2442,N_2432);
nor U2709 (N_2709,N_2523,N_2505);
nand U2710 (N_2710,N_2559,N_2461);
nand U2711 (N_2711,N_2436,N_2432);
nor U2712 (N_2712,N_2454,N_2492);
nand U2713 (N_2713,N_2416,N_2401);
or U2714 (N_2714,N_2548,N_2485);
nand U2715 (N_2715,N_2402,N_2492);
and U2716 (N_2716,N_2455,N_2421);
and U2717 (N_2717,N_2437,N_2435);
or U2718 (N_2718,N_2571,N_2449);
and U2719 (N_2719,N_2539,N_2511);
xnor U2720 (N_2720,N_2467,N_2505);
nor U2721 (N_2721,N_2417,N_2559);
xor U2722 (N_2722,N_2561,N_2431);
or U2723 (N_2723,N_2432,N_2514);
or U2724 (N_2724,N_2478,N_2577);
nand U2725 (N_2725,N_2527,N_2490);
or U2726 (N_2726,N_2599,N_2518);
nand U2727 (N_2727,N_2538,N_2586);
xor U2728 (N_2728,N_2447,N_2404);
or U2729 (N_2729,N_2496,N_2511);
nand U2730 (N_2730,N_2568,N_2574);
and U2731 (N_2731,N_2534,N_2586);
and U2732 (N_2732,N_2456,N_2552);
nor U2733 (N_2733,N_2555,N_2494);
nor U2734 (N_2734,N_2589,N_2566);
nand U2735 (N_2735,N_2554,N_2502);
nor U2736 (N_2736,N_2591,N_2464);
or U2737 (N_2737,N_2541,N_2598);
xnor U2738 (N_2738,N_2417,N_2488);
and U2739 (N_2739,N_2466,N_2524);
xor U2740 (N_2740,N_2596,N_2462);
nand U2741 (N_2741,N_2551,N_2414);
nand U2742 (N_2742,N_2440,N_2480);
xnor U2743 (N_2743,N_2419,N_2533);
and U2744 (N_2744,N_2423,N_2467);
nor U2745 (N_2745,N_2482,N_2546);
xnor U2746 (N_2746,N_2466,N_2586);
nor U2747 (N_2747,N_2523,N_2590);
nand U2748 (N_2748,N_2482,N_2402);
nor U2749 (N_2749,N_2532,N_2518);
and U2750 (N_2750,N_2442,N_2500);
and U2751 (N_2751,N_2405,N_2435);
and U2752 (N_2752,N_2597,N_2598);
or U2753 (N_2753,N_2498,N_2594);
nand U2754 (N_2754,N_2437,N_2409);
and U2755 (N_2755,N_2476,N_2404);
nor U2756 (N_2756,N_2522,N_2417);
and U2757 (N_2757,N_2456,N_2548);
or U2758 (N_2758,N_2531,N_2528);
nand U2759 (N_2759,N_2583,N_2552);
or U2760 (N_2760,N_2580,N_2588);
nand U2761 (N_2761,N_2467,N_2491);
nand U2762 (N_2762,N_2420,N_2457);
or U2763 (N_2763,N_2590,N_2500);
nand U2764 (N_2764,N_2591,N_2534);
nand U2765 (N_2765,N_2502,N_2575);
xor U2766 (N_2766,N_2576,N_2548);
nand U2767 (N_2767,N_2446,N_2531);
and U2768 (N_2768,N_2509,N_2429);
and U2769 (N_2769,N_2449,N_2445);
nor U2770 (N_2770,N_2436,N_2401);
xnor U2771 (N_2771,N_2454,N_2520);
and U2772 (N_2772,N_2587,N_2571);
xnor U2773 (N_2773,N_2487,N_2504);
or U2774 (N_2774,N_2599,N_2490);
nor U2775 (N_2775,N_2447,N_2401);
nand U2776 (N_2776,N_2575,N_2576);
or U2777 (N_2777,N_2444,N_2431);
nand U2778 (N_2778,N_2563,N_2455);
nor U2779 (N_2779,N_2529,N_2462);
or U2780 (N_2780,N_2534,N_2492);
nand U2781 (N_2781,N_2414,N_2478);
nor U2782 (N_2782,N_2498,N_2504);
or U2783 (N_2783,N_2585,N_2475);
nor U2784 (N_2784,N_2415,N_2411);
nor U2785 (N_2785,N_2436,N_2506);
or U2786 (N_2786,N_2422,N_2585);
or U2787 (N_2787,N_2551,N_2578);
nor U2788 (N_2788,N_2585,N_2489);
and U2789 (N_2789,N_2448,N_2430);
and U2790 (N_2790,N_2452,N_2514);
or U2791 (N_2791,N_2420,N_2431);
nor U2792 (N_2792,N_2536,N_2407);
nand U2793 (N_2793,N_2543,N_2558);
nor U2794 (N_2794,N_2590,N_2561);
nor U2795 (N_2795,N_2478,N_2456);
nor U2796 (N_2796,N_2453,N_2531);
or U2797 (N_2797,N_2452,N_2599);
or U2798 (N_2798,N_2509,N_2518);
nand U2799 (N_2799,N_2543,N_2566);
or U2800 (N_2800,N_2710,N_2755);
and U2801 (N_2801,N_2611,N_2768);
or U2802 (N_2802,N_2707,N_2797);
and U2803 (N_2803,N_2704,N_2667);
or U2804 (N_2804,N_2762,N_2673);
nand U2805 (N_2805,N_2692,N_2701);
nor U2806 (N_2806,N_2703,N_2770);
and U2807 (N_2807,N_2625,N_2614);
and U2808 (N_2808,N_2690,N_2641);
nand U2809 (N_2809,N_2757,N_2685);
and U2810 (N_2810,N_2785,N_2767);
and U2811 (N_2811,N_2706,N_2695);
nor U2812 (N_2812,N_2780,N_2786);
nand U2813 (N_2813,N_2605,N_2769);
or U2814 (N_2814,N_2604,N_2718);
nor U2815 (N_2815,N_2680,N_2663);
nor U2816 (N_2816,N_2603,N_2721);
nor U2817 (N_2817,N_2630,N_2631);
nand U2818 (N_2818,N_2615,N_2745);
nand U2819 (N_2819,N_2618,N_2645);
xnor U2820 (N_2820,N_2682,N_2664);
nor U2821 (N_2821,N_2602,N_2782);
nand U2822 (N_2822,N_2727,N_2709);
nor U2823 (N_2823,N_2705,N_2660);
or U2824 (N_2824,N_2699,N_2662);
and U2825 (N_2825,N_2672,N_2650);
and U2826 (N_2826,N_2734,N_2624);
and U2827 (N_2827,N_2732,N_2788);
or U2828 (N_2828,N_2717,N_2617);
nand U2829 (N_2829,N_2772,N_2616);
and U2830 (N_2830,N_2665,N_2669);
and U2831 (N_2831,N_2775,N_2713);
nor U2832 (N_2832,N_2653,N_2798);
and U2833 (N_2833,N_2750,N_2626);
xnor U2834 (N_2834,N_2647,N_2627);
nor U2835 (N_2835,N_2688,N_2670);
and U2836 (N_2836,N_2621,N_2729);
nand U2837 (N_2837,N_2787,N_2689);
and U2838 (N_2838,N_2691,N_2760);
and U2839 (N_2839,N_2679,N_2693);
nor U2840 (N_2840,N_2675,N_2684);
or U2841 (N_2841,N_2799,N_2697);
nand U2842 (N_2842,N_2678,N_2607);
and U2843 (N_2843,N_2714,N_2702);
and U2844 (N_2844,N_2640,N_2716);
nor U2845 (N_2845,N_2642,N_2742);
and U2846 (N_2846,N_2711,N_2676);
nor U2847 (N_2847,N_2759,N_2756);
and U2848 (N_2848,N_2600,N_2712);
or U2849 (N_2849,N_2737,N_2773);
or U2850 (N_2850,N_2781,N_2700);
nand U2851 (N_2851,N_2637,N_2698);
and U2852 (N_2852,N_2765,N_2741);
or U2853 (N_2853,N_2636,N_2620);
or U2854 (N_2854,N_2613,N_2779);
nand U2855 (N_2855,N_2736,N_2683);
or U2856 (N_2856,N_2666,N_2635);
xnor U2857 (N_2857,N_2654,N_2790);
nor U2858 (N_2858,N_2687,N_2612);
and U2859 (N_2859,N_2726,N_2795);
xor U2860 (N_2860,N_2789,N_2656);
or U2861 (N_2861,N_2784,N_2606);
and U2862 (N_2862,N_2661,N_2761);
nand U2863 (N_2863,N_2724,N_2766);
or U2864 (N_2864,N_2694,N_2719);
nand U2865 (N_2865,N_2651,N_2601);
xor U2866 (N_2866,N_2658,N_2791);
nor U2867 (N_2867,N_2735,N_2733);
and U2868 (N_2868,N_2752,N_2731);
nand U2869 (N_2869,N_2722,N_2659);
nor U2870 (N_2870,N_2623,N_2681);
xnor U2871 (N_2871,N_2793,N_2668);
nand U2872 (N_2872,N_2655,N_2629);
nand U2873 (N_2873,N_2748,N_2708);
and U2874 (N_2874,N_2744,N_2730);
and U2875 (N_2875,N_2634,N_2725);
or U2876 (N_2876,N_2646,N_2674);
nand U2877 (N_2877,N_2738,N_2764);
or U2878 (N_2878,N_2740,N_2622);
nand U2879 (N_2879,N_2608,N_2639);
and U2880 (N_2880,N_2783,N_2715);
nor U2881 (N_2881,N_2758,N_2794);
xnor U2882 (N_2882,N_2628,N_2657);
nor U2883 (N_2883,N_2644,N_2633);
and U2884 (N_2884,N_2638,N_2796);
xnor U2885 (N_2885,N_2746,N_2749);
nand U2886 (N_2886,N_2609,N_2753);
and U2887 (N_2887,N_2774,N_2739);
nor U2888 (N_2888,N_2619,N_2743);
nand U2889 (N_2889,N_2771,N_2728);
and U2890 (N_2890,N_2643,N_2792);
nand U2891 (N_2891,N_2632,N_2754);
xnor U2892 (N_2892,N_2723,N_2763);
nor U2893 (N_2893,N_2652,N_2778);
xor U2894 (N_2894,N_2777,N_2649);
and U2895 (N_2895,N_2686,N_2776);
and U2896 (N_2896,N_2610,N_2696);
nor U2897 (N_2897,N_2747,N_2671);
or U2898 (N_2898,N_2720,N_2751);
and U2899 (N_2899,N_2648,N_2677);
and U2900 (N_2900,N_2736,N_2771);
xor U2901 (N_2901,N_2684,N_2667);
and U2902 (N_2902,N_2633,N_2704);
nor U2903 (N_2903,N_2630,N_2677);
or U2904 (N_2904,N_2665,N_2744);
nor U2905 (N_2905,N_2786,N_2723);
nor U2906 (N_2906,N_2724,N_2799);
and U2907 (N_2907,N_2711,N_2612);
nand U2908 (N_2908,N_2606,N_2616);
or U2909 (N_2909,N_2602,N_2772);
and U2910 (N_2910,N_2691,N_2742);
xor U2911 (N_2911,N_2792,N_2639);
or U2912 (N_2912,N_2688,N_2781);
xor U2913 (N_2913,N_2714,N_2690);
and U2914 (N_2914,N_2753,N_2752);
or U2915 (N_2915,N_2683,N_2633);
nor U2916 (N_2916,N_2705,N_2777);
xor U2917 (N_2917,N_2693,N_2612);
nand U2918 (N_2918,N_2787,N_2749);
or U2919 (N_2919,N_2695,N_2616);
xor U2920 (N_2920,N_2680,N_2755);
or U2921 (N_2921,N_2724,N_2797);
nand U2922 (N_2922,N_2755,N_2661);
nor U2923 (N_2923,N_2796,N_2755);
and U2924 (N_2924,N_2779,N_2782);
xnor U2925 (N_2925,N_2665,N_2786);
nor U2926 (N_2926,N_2772,N_2727);
nand U2927 (N_2927,N_2691,N_2703);
or U2928 (N_2928,N_2708,N_2755);
nand U2929 (N_2929,N_2708,N_2689);
and U2930 (N_2930,N_2679,N_2603);
nand U2931 (N_2931,N_2703,N_2652);
nand U2932 (N_2932,N_2625,N_2773);
xnor U2933 (N_2933,N_2797,N_2757);
or U2934 (N_2934,N_2717,N_2723);
nand U2935 (N_2935,N_2636,N_2772);
nand U2936 (N_2936,N_2645,N_2776);
and U2937 (N_2937,N_2629,N_2676);
and U2938 (N_2938,N_2607,N_2769);
nor U2939 (N_2939,N_2734,N_2693);
nor U2940 (N_2940,N_2756,N_2760);
nor U2941 (N_2941,N_2665,N_2643);
or U2942 (N_2942,N_2723,N_2796);
xor U2943 (N_2943,N_2666,N_2798);
nor U2944 (N_2944,N_2768,N_2657);
or U2945 (N_2945,N_2736,N_2667);
or U2946 (N_2946,N_2694,N_2763);
or U2947 (N_2947,N_2654,N_2708);
nor U2948 (N_2948,N_2617,N_2624);
and U2949 (N_2949,N_2633,N_2640);
nand U2950 (N_2950,N_2636,N_2602);
nand U2951 (N_2951,N_2774,N_2636);
and U2952 (N_2952,N_2760,N_2604);
and U2953 (N_2953,N_2604,N_2660);
and U2954 (N_2954,N_2729,N_2696);
nor U2955 (N_2955,N_2622,N_2634);
nor U2956 (N_2956,N_2627,N_2707);
and U2957 (N_2957,N_2671,N_2678);
nor U2958 (N_2958,N_2796,N_2695);
nor U2959 (N_2959,N_2679,N_2789);
xnor U2960 (N_2960,N_2683,N_2665);
xnor U2961 (N_2961,N_2739,N_2756);
nor U2962 (N_2962,N_2641,N_2681);
xor U2963 (N_2963,N_2630,N_2765);
and U2964 (N_2964,N_2719,N_2607);
or U2965 (N_2965,N_2782,N_2681);
nor U2966 (N_2966,N_2704,N_2750);
nand U2967 (N_2967,N_2625,N_2709);
or U2968 (N_2968,N_2654,N_2784);
nor U2969 (N_2969,N_2743,N_2738);
nor U2970 (N_2970,N_2648,N_2678);
xor U2971 (N_2971,N_2720,N_2625);
nor U2972 (N_2972,N_2664,N_2661);
and U2973 (N_2973,N_2727,N_2620);
xor U2974 (N_2974,N_2790,N_2763);
and U2975 (N_2975,N_2673,N_2741);
and U2976 (N_2976,N_2601,N_2657);
and U2977 (N_2977,N_2776,N_2671);
or U2978 (N_2978,N_2668,N_2720);
and U2979 (N_2979,N_2692,N_2774);
nand U2980 (N_2980,N_2725,N_2718);
nand U2981 (N_2981,N_2752,N_2604);
or U2982 (N_2982,N_2790,N_2624);
xnor U2983 (N_2983,N_2689,N_2654);
xnor U2984 (N_2984,N_2755,N_2699);
nand U2985 (N_2985,N_2687,N_2748);
or U2986 (N_2986,N_2782,N_2770);
and U2987 (N_2987,N_2790,N_2631);
or U2988 (N_2988,N_2652,N_2617);
or U2989 (N_2989,N_2625,N_2688);
or U2990 (N_2990,N_2770,N_2606);
or U2991 (N_2991,N_2645,N_2792);
or U2992 (N_2992,N_2692,N_2685);
and U2993 (N_2993,N_2667,N_2671);
nand U2994 (N_2994,N_2614,N_2666);
nor U2995 (N_2995,N_2708,N_2601);
or U2996 (N_2996,N_2671,N_2712);
nor U2997 (N_2997,N_2681,N_2799);
nand U2998 (N_2998,N_2662,N_2762);
and U2999 (N_2999,N_2662,N_2634);
nand UO_0 (O_0,N_2916,N_2920);
and UO_1 (O_1,N_2886,N_2804);
nor UO_2 (O_2,N_2880,N_2825);
nor UO_3 (O_3,N_2841,N_2963);
xnor UO_4 (O_4,N_2848,N_2930);
or UO_5 (O_5,N_2887,N_2924);
or UO_6 (O_6,N_2818,N_2821);
or UO_7 (O_7,N_2948,N_2883);
and UO_8 (O_8,N_2875,N_2929);
nor UO_9 (O_9,N_2942,N_2871);
nor UO_10 (O_10,N_2838,N_2826);
and UO_11 (O_11,N_2890,N_2975);
or UO_12 (O_12,N_2867,N_2876);
and UO_13 (O_13,N_2809,N_2981);
nand UO_14 (O_14,N_2979,N_2943);
or UO_15 (O_15,N_2952,N_2895);
nand UO_16 (O_16,N_2878,N_2976);
nand UO_17 (O_17,N_2915,N_2800);
and UO_18 (O_18,N_2859,N_2803);
and UO_19 (O_19,N_2947,N_2937);
nor UO_20 (O_20,N_2901,N_2899);
and UO_21 (O_21,N_2870,N_2802);
or UO_22 (O_22,N_2862,N_2970);
and UO_23 (O_23,N_2957,N_2971);
and UO_24 (O_24,N_2819,N_2908);
nor UO_25 (O_25,N_2842,N_2810);
or UO_26 (O_26,N_2808,N_2989);
nand UO_27 (O_27,N_2852,N_2933);
and UO_28 (O_28,N_2868,N_2982);
nor UO_29 (O_29,N_2977,N_2974);
and UO_30 (O_30,N_2815,N_2836);
xnor UO_31 (O_31,N_2997,N_2950);
or UO_32 (O_32,N_2961,N_2900);
nand UO_33 (O_33,N_2839,N_2824);
or UO_34 (O_34,N_2837,N_2965);
nand UO_35 (O_35,N_2832,N_2991);
nand UO_36 (O_36,N_2850,N_2938);
or UO_37 (O_37,N_2892,N_2881);
or UO_38 (O_38,N_2993,N_2851);
or UO_39 (O_39,N_2806,N_2857);
and UO_40 (O_40,N_2820,N_2972);
nand UO_41 (O_41,N_2807,N_2918);
nor UO_42 (O_42,N_2829,N_2994);
or UO_43 (O_43,N_2902,N_2864);
nand UO_44 (O_44,N_2967,N_2903);
nor UO_45 (O_45,N_2854,N_2934);
nor UO_46 (O_46,N_2898,N_2905);
nor UO_47 (O_47,N_2823,N_2966);
xor UO_48 (O_48,N_2985,N_2874);
nor UO_49 (O_49,N_2834,N_2831);
nor UO_50 (O_50,N_2885,N_2987);
nor UO_51 (O_51,N_2984,N_2827);
nand UO_52 (O_52,N_2928,N_2865);
or UO_53 (O_53,N_2889,N_2995);
nand UO_54 (O_54,N_2983,N_2962);
xnor UO_55 (O_55,N_2830,N_2805);
nand UO_56 (O_56,N_2860,N_2907);
nand UO_57 (O_57,N_2855,N_2922);
and UO_58 (O_58,N_2990,N_2861);
or UO_59 (O_59,N_2906,N_2944);
nand UO_60 (O_60,N_2911,N_2949);
or UO_61 (O_61,N_2833,N_2847);
and UO_62 (O_62,N_2925,N_2873);
nor UO_63 (O_63,N_2960,N_2904);
or UO_64 (O_64,N_2939,N_2884);
nand UO_65 (O_65,N_2910,N_2986);
or UO_66 (O_66,N_2973,N_2882);
or UO_67 (O_67,N_2998,N_2816);
nor UO_68 (O_68,N_2914,N_2921);
and UO_69 (O_69,N_2877,N_2814);
nand UO_70 (O_70,N_2956,N_2945);
or UO_71 (O_71,N_2955,N_2988);
nand UO_72 (O_72,N_2931,N_2856);
nand UO_73 (O_73,N_2980,N_2872);
or UO_74 (O_74,N_2936,N_2888);
and UO_75 (O_75,N_2845,N_2849);
and UO_76 (O_76,N_2840,N_2959);
xor UO_77 (O_77,N_2968,N_2935);
nor UO_78 (O_78,N_2869,N_2893);
nor UO_79 (O_79,N_2894,N_2941);
nor UO_80 (O_80,N_2919,N_2996);
xnor UO_81 (O_81,N_2958,N_2858);
and UO_82 (O_82,N_2946,N_2917);
nor UO_83 (O_83,N_2927,N_2843);
or UO_84 (O_84,N_2896,N_2953);
nand UO_85 (O_85,N_2926,N_2822);
nand UO_86 (O_86,N_2964,N_2992);
xnor UO_87 (O_87,N_2912,N_2940);
xor UO_88 (O_88,N_2866,N_2913);
nor UO_89 (O_89,N_2853,N_2863);
nor UO_90 (O_90,N_2835,N_2954);
and UO_91 (O_91,N_2879,N_2999);
xor UO_92 (O_92,N_2817,N_2891);
or UO_93 (O_93,N_2828,N_2813);
or UO_94 (O_94,N_2909,N_2923);
or UO_95 (O_95,N_2951,N_2811);
or UO_96 (O_96,N_2897,N_2932);
or UO_97 (O_97,N_2844,N_2978);
or UO_98 (O_98,N_2801,N_2969);
nand UO_99 (O_99,N_2846,N_2812);
xor UO_100 (O_100,N_2952,N_2942);
nand UO_101 (O_101,N_2865,N_2932);
nor UO_102 (O_102,N_2902,N_2912);
nand UO_103 (O_103,N_2889,N_2861);
xnor UO_104 (O_104,N_2810,N_2992);
and UO_105 (O_105,N_2981,N_2909);
nor UO_106 (O_106,N_2836,N_2867);
nand UO_107 (O_107,N_2937,N_2868);
nand UO_108 (O_108,N_2992,N_2845);
nand UO_109 (O_109,N_2925,N_2894);
xor UO_110 (O_110,N_2995,N_2947);
nor UO_111 (O_111,N_2881,N_2995);
nand UO_112 (O_112,N_2948,N_2866);
xor UO_113 (O_113,N_2814,N_2888);
and UO_114 (O_114,N_2878,N_2861);
nor UO_115 (O_115,N_2936,N_2951);
or UO_116 (O_116,N_2932,N_2886);
and UO_117 (O_117,N_2976,N_2849);
or UO_118 (O_118,N_2936,N_2922);
nand UO_119 (O_119,N_2996,N_2902);
nand UO_120 (O_120,N_2929,N_2944);
or UO_121 (O_121,N_2963,N_2882);
and UO_122 (O_122,N_2975,N_2978);
and UO_123 (O_123,N_2854,N_2945);
nor UO_124 (O_124,N_2806,N_2988);
nor UO_125 (O_125,N_2928,N_2903);
nor UO_126 (O_126,N_2921,N_2992);
and UO_127 (O_127,N_2987,N_2829);
nor UO_128 (O_128,N_2971,N_2833);
and UO_129 (O_129,N_2942,N_2931);
nand UO_130 (O_130,N_2823,N_2815);
nor UO_131 (O_131,N_2818,N_2815);
xnor UO_132 (O_132,N_2852,N_2922);
or UO_133 (O_133,N_2822,N_2860);
nor UO_134 (O_134,N_2973,N_2918);
or UO_135 (O_135,N_2952,N_2820);
or UO_136 (O_136,N_2806,N_2918);
xor UO_137 (O_137,N_2880,N_2813);
and UO_138 (O_138,N_2961,N_2819);
and UO_139 (O_139,N_2837,N_2963);
nand UO_140 (O_140,N_2969,N_2813);
nand UO_141 (O_141,N_2811,N_2966);
nand UO_142 (O_142,N_2966,N_2914);
or UO_143 (O_143,N_2953,N_2809);
nand UO_144 (O_144,N_2864,N_2978);
and UO_145 (O_145,N_2834,N_2892);
nor UO_146 (O_146,N_2817,N_2979);
or UO_147 (O_147,N_2949,N_2843);
nand UO_148 (O_148,N_2873,N_2923);
nor UO_149 (O_149,N_2855,N_2864);
nand UO_150 (O_150,N_2867,N_2954);
and UO_151 (O_151,N_2827,N_2995);
nor UO_152 (O_152,N_2860,N_2881);
or UO_153 (O_153,N_2828,N_2904);
and UO_154 (O_154,N_2838,N_2996);
and UO_155 (O_155,N_2882,N_2807);
and UO_156 (O_156,N_2864,N_2819);
or UO_157 (O_157,N_2976,N_2824);
or UO_158 (O_158,N_2956,N_2870);
nand UO_159 (O_159,N_2988,N_2856);
or UO_160 (O_160,N_2936,N_2945);
nand UO_161 (O_161,N_2914,N_2857);
and UO_162 (O_162,N_2829,N_2957);
or UO_163 (O_163,N_2912,N_2850);
or UO_164 (O_164,N_2853,N_2905);
nor UO_165 (O_165,N_2947,N_2816);
and UO_166 (O_166,N_2859,N_2860);
nand UO_167 (O_167,N_2977,N_2928);
nand UO_168 (O_168,N_2845,N_2838);
and UO_169 (O_169,N_2897,N_2831);
and UO_170 (O_170,N_2846,N_2835);
and UO_171 (O_171,N_2976,N_2829);
or UO_172 (O_172,N_2976,N_2822);
nand UO_173 (O_173,N_2941,N_2850);
and UO_174 (O_174,N_2849,N_2939);
or UO_175 (O_175,N_2853,N_2948);
or UO_176 (O_176,N_2962,N_2807);
or UO_177 (O_177,N_2876,N_2978);
or UO_178 (O_178,N_2934,N_2814);
nand UO_179 (O_179,N_2921,N_2916);
or UO_180 (O_180,N_2812,N_2960);
and UO_181 (O_181,N_2899,N_2839);
and UO_182 (O_182,N_2855,N_2930);
or UO_183 (O_183,N_2971,N_2866);
nor UO_184 (O_184,N_2961,N_2929);
nor UO_185 (O_185,N_2947,N_2993);
nor UO_186 (O_186,N_2829,N_2836);
xor UO_187 (O_187,N_2846,N_2862);
nand UO_188 (O_188,N_2986,N_2990);
or UO_189 (O_189,N_2858,N_2845);
nor UO_190 (O_190,N_2944,N_2901);
and UO_191 (O_191,N_2935,N_2945);
xnor UO_192 (O_192,N_2904,N_2906);
and UO_193 (O_193,N_2930,N_2901);
xor UO_194 (O_194,N_2878,N_2882);
or UO_195 (O_195,N_2875,N_2818);
nor UO_196 (O_196,N_2832,N_2977);
or UO_197 (O_197,N_2854,N_2991);
and UO_198 (O_198,N_2870,N_2904);
or UO_199 (O_199,N_2914,N_2938);
or UO_200 (O_200,N_2976,N_2953);
xor UO_201 (O_201,N_2852,N_2816);
nor UO_202 (O_202,N_2868,N_2922);
nor UO_203 (O_203,N_2946,N_2957);
nand UO_204 (O_204,N_2883,N_2833);
nand UO_205 (O_205,N_2853,N_2929);
or UO_206 (O_206,N_2953,N_2925);
and UO_207 (O_207,N_2945,N_2963);
nand UO_208 (O_208,N_2869,N_2881);
or UO_209 (O_209,N_2898,N_2843);
or UO_210 (O_210,N_2821,N_2869);
nand UO_211 (O_211,N_2821,N_2985);
and UO_212 (O_212,N_2910,N_2812);
or UO_213 (O_213,N_2887,N_2986);
xnor UO_214 (O_214,N_2841,N_2885);
or UO_215 (O_215,N_2899,N_2907);
or UO_216 (O_216,N_2979,N_2813);
and UO_217 (O_217,N_2881,N_2986);
nand UO_218 (O_218,N_2847,N_2899);
and UO_219 (O_219,N_2974,N_2870);
or UO_220 (O_220,N_2952,N_2862);
and UO_221 (O_221,N_2801,N_2828);
nand UO_222 (O_222,N_2951,N_2850);
or UO_223 (O_223,N_2885,N_2935);
nand UO_224 (O_224,N_2948,N_2805);
nand UO_225 (O_225,N_2879,N_2911);
or UO_226 (O_226,N_2951,N_2827);
nand UO_227 (O_227,N_2871,N_2999);
or UO_228 (O_228,N_2822,N_2989);
nor UO_229 (O_229,N_2819,N_2890);
and UO_230 (O_230,N_2929,N_2870);
nor UO_231 (O_231,N_2816,N_2984);
and UO_232 (O_232,N_2955,N_2800);
and UO_233 (O_233,N_2856,N_2987);
xor UO_234 (O_234,N_2959,N_2829);
and UO_235 (O_235,N_2835,N_2865);
or UO_236 (O_236,N_2904,N_2929);
and UO_237 (O_237,N_2959,N_2972);
nand UO_238 (O_238,N_2967,N_2825);
xnor UO_239 (O_239,N_2848,N_2991);
nand UO_240 (O_240,N_2800,N_2808);
or UO_241 (O_241,N_2871,N_2979);
or UO_242 (O_242,N_2927,N_2946);
nor UO_243 (O_243,N_2878,N_2886);
and UO_244 (O_244,N_2805,N_2986);
nand UO_245 (O_245,N_2952,N_2999);
or UO_246 (O_246,N_2928,N_2972);
nor UO_247 (O_247,N_2856,N_2865);
nor UO_248 (O_248,N_2886,N_2855);
and UO_249 (O_249,N_2992,N_2955);
and UO_250 (O_250,N_2824,N_2903);
nand UO_251 (O_251,N_2894,N_2848);
xnor UO_252 (O_252,N_2936,N_2824);
xnor UO_253 (O_253,N_2936,N_2846);
or UO_254 (O_254,N_2810,N_2998);
nand UO_255 (O_255,N_2908,N_2904);
or UO_256 (O_256,N_2907,N_2867);
and UO_257 (O_257,N_2945,N_2928);
nand UO_258 (O_258,N_2870,N_2848);
and UO_259 (O_259,N_2813,N_2948);
xor UO_260 (O_260,N_2807,N_2891);
or UO_261 (O_261,N_2925,N_2901);
nor UO_262 (O_262,N_2976,N_2979);
nand UO_263 (O_263,N_2982,N_2836);
xor UO_264 (O_264,N_2897,N_2974);
or UO_265 (O_265,N_2884,N_2937);
and UO_266 (O_266,N_2938,N_2807);
and UO_267 (O_267,N_2898,N_2986);
nor UO_268 (O_268,N_2930,N_2814);
nor UO_269 (O_269,N_2960,N_2907);
nor UO_270 (O_270,N_2890,N_2984);
nor UO_271 (O_271,N_2831,N_2957);
nand UO_272 (O_272,N_2893,N_2824);
nor UO_273 (O_273,N_2900,N_2911);
nor UO_274 (O_274,N_2886,N_2895);
nor UO_275 (O_275,N_2931,N_2850);
nand UO_276 (O_276,N_2954,N_2930);
xnor UO_277 (O_277,N_2869,N_2997);
and UO_278 (O_278,N_2860,N_2931);
xnor UO_279 (O_279,N_2802,N_2883);
or UO_280 (O_280,N_2947,N_2812);
xor UO_281 (O_281,N_2952,N_2817);
nand UO_282 (O_282,N_2996,N_2968);
or UO_283 (O_283,N_2892,N_2837);
xor UO_284 (O_284,N_2898,N_2844);
or UO_285 (O_285,N_2913,N_2918);
and UO_286 (O_286,N_2806,N_2913);
nor UO_287 (O_287,N_2881,N_2858);
nor UO_288 (O_288,N_2909,N_2962);
nand UO_289 (O_289,N_2925,N_2829);
and UO_290 (O_290,N_2900,N_2953);
or UO_291 (O_291,N_2924,N_2909);
nor UO_292 (O_292,N_2933,N_2886);
or UO_293 (O_293,N_2823,N_2824);
and UO_294 (O_294,N_2866,N_2946);
or UO_295 (O_295,N_2897,N_2944);
xnor UO_296 (O_296,N_2952,N_2917);
xor UO_297 (O_297,N_2813,N_2863);
xnor UO_298 (O_298,N_2853,N_2928);
nand UO_299 (O_299,N_2946,N_2945);
or UO_300 (O_300,N_2845,N_2996);
nor UO_301 (O_301,N_2984,N_2808);
nor UO_302 (O_302,N_2810,N_2903);
and UO_303 (O_303,N_2889,N_2836);
nand UO_304 (O_304,N_2853,N_2849);
and UO_305 (O_305,N_2821,N_2847);
or UO_306 (O_306,N_2875,N_2864);
nand UO_307 (O_307,N_2841,N_2831);
nand UO_308 (O_308,N_2847,N_2870);
and UO_309 (O_309,N_2845,N_2944);
xnor UO_310 (O_310,N_2988,N_2864);
and UO_311 (O_311,N_2824,N_2950);
and UO_312 (O_312,N_2858,N_2943);
or UO_313 (O_313,N_2837,N_2946);
nor UO_314 (O_314,N_2840,N_2880);
or UO_315 (O_315,N_2992,N_2837);
nor UO_316 (O_316,N_2948,N_2855);
nand UO_317 (O_317,N_2906,N_2844);
and UO_318 (O_318,N_2998,N_2846);
nor UO_319 (O_319,N_2802,N_2962);
xor UO_320 (O_320,N_2819,N_2945);
nand UO_321 (O_321,N_2910,N_2805);
nor UO_322 (O_322,N_2955,N_2933);
or UO_323 (O_323,N_2879,N_2895);
nor UO_324 (O_324,N_2966,N_2804);
or UO_325 (O_325,N_2835,N_2820);
nor UO_326 (O_326,N_2926,N_2805);
or UO_327 (O_327,N_2945,N_2807);
nor UO_328 (O_328,N_2808,N_2985);
nand UO_329 (O_329,N_2845,N_2894);
and UO_330 (O_330,N_2945,N_2996);
or UO_331 (O_331,N_2942,N_2996);
nand UO_332 (O_332,N_2827,N_2821);
xor UO_333 (O_333,N_2852,N_2932);
xnor UO_334 (O_334,N_2865,N_2815);
nor UO_335 (O_335,N_2811,N_2989);
and UO_336 (O_336,N_2810,N_2839);
and UO_337 (O_337,N_2875,N_2950);
nor UO_338 (O_338,N_2942,N_2977);
nand UO_339 (O_339,N_2848,N_2927);
or UO_340 (O_340,N_2876,N_2814);
nor UO_341 (O_341,N_2986,N_2842);
nor UO_342 (O_342,N_2849,N_2840);
nand UO_343 (O_343,N_2818,N_2884);
or UO_344 (O_344,N_2973,N_2873);
or UO_345 (O_345,N_2990,N_2967);
and UO_346 (O_346,N_2923,N_2895);
and UO_347 (O_347,N_2896,N_2844);
nor UO_348 (O_348,N_2814,N_2965);
nor UO_349 (O_349,N_2969,N_2952);
xnor UO_350 (O_350,N_2840,N_2818);
and UO_351 (O_351,N_2817,N_2989);
xor UO_352 (O_352,N_2971,N_2949);
and UO_353 (O_353,N_2903,N_2933);
xor UO_354 (O_354,N_2898,N_2985);
or UO_355 (O_355,N_2813,N_2913);
or UO_356 (O_356,N_2892,N_2916);
and UO_357 (O_357,N_2918,N_2891);
nand UO_358 (O_358,N_2997,N_2828);
or UO_359 (O_359,N_2971,N_2983);
nand UO_360 (O_360,N_2883,N_2827);
nand UO_361 (O_361,N_2922,N_2847);
or UO_362 (O_362,N_2813,N_2837);
nor UO_363 (O_363,N_2933,N_2805);
or UO_364 (O_364,N_2800,N_2905);
nand UO_365 (O_365,N_2803,N_2811);
nand UO_366 (O_366,N_2808,N_2967);
nand UO_367 (O_367,N_2991,N_2923);
nor UO_368 (O_368,N_2988,N_2827);
nand UO_369 (O_369,N_2874,N_2840);
nand UO_370 (O_370,N_2937,N_2866);
xnor UO_371 (O_371,N_2815,N_2811);
nand UO_372 (O_372,N_2818,N_2812);
xor UO_373 (O_373,N_2983,N_2843);
xnor UO_374 (O_374,N_2984,N_2913);
nand UO_375 (O_375,N_2817,N_2815);
nand UO_376 (O_376,N_2882,N_2947);
nand UO_377 (O_377,N_2880,N_2908);
or UO_378 (O_378,N_2862,N_2997);
nand UO_379 (O_379,N_2910,N_2856);
and UO_380 (O_380,N_2918,N_2809);
nor UO_381 (O_381,N_2903,N_2948);
nor UO_382 (O_382,N_2934,N_2881);
and UO_383 (O_383,N_2969,N_2887);
and UO_384 (O_384,N_2879,N_2978);
or UO_385 (O_385,N_2948,N_2909);
xnor UO_386 (O_386,N_2967,N_2869);
nand UO_387 (O_387,N_2812,N_2948);
and UO_388 (O_388,N_2956,N_2896);
and UO_389 (O_389,N_2925,N_2859);
and UO_390 (O_390,N_2969,N_2964);
nand UO_391 (O_391,N_2832,N_2852);
nand UO_392 (O_392,N_2839,N_2993);
or UO_393 (O_393,N_2884,N_2833);
nand UO_394 (O_394,N_2882,N_2979);
nand UO_395 (O_395,N_2971,N_2895);
xor UO_396 (O_396,N_2928,N_2877);
nor UO_397 (O_397,N_2963,N_2807);
and UO_398 (O_398,N_2828,N_2851);
or UO_399 (O_399,N_2884,N_2932);
or UO_400 (O_400,N_2806,N_2991);
nand UO_401 (O_401,N_2855,N_2918);
nor UO_402 (O_402,N_2969,N_2942);
nor UO_403 (O_403,N_2916,N_2990);
and UO_404 (O_404,N_2975,N_2948);
nand UO_405 (O_405,N_2926,N_2901);
xnor UO_406 (O_406,N_2917,N_2833);
or UO_407 (O_407,N_2805,N_2970);
or UO_408 (O_408,N_2931,N_2950);
or UO_409 (O_409,N_2863,N_2906);
nand UO_410 (O_410,N_2918,N_2820);
and UO_411 (O_411,N_2958,N_2820);
nand UO_412 (O_412,N_2822,N_2947);
nor UO_413 (O_413,N_2833,N_2904);
nand UO_414 (O_414,N_2996,N_2872);
or UO_415 (O_415,N_2899,N_2842);
nor UO_416 (O_416,N_2943,N_2809);
and UO_417 (O_417,N_2964,N_2931);
and UO_418 (O_418,N_2848,N_2813);
or UO_419 (O_419,N_2945,N_2921);
and UO_420 (O_420,N_2857,N_2935);
nor UO_421 (O_421,N_2855,N_2981);
and UO_422 (O_422,N_2870,N_2912);
and UO_423 (O_423,N_2876,N_2906);
nand UO_424 (O_424,N_2970,N_2849);
nor UO_425 (O_425,N_2902,N_2919);
xnor UO_426 (O_426,N_2975,N_2865);
and UO_427 (O_427,N_2933,N_2932);
or UO_428 (O_428,N_2938,N_2803);
nor UO_429 (O_429,N_2805,N_2892);
xnor UO_430 (O_430,N_2974,N_2998);
nor UO_431 (O_431,N_2973,N_2938);
nor UO_432 (O_432,N_2889,N_2866);
nor UO_433 (O_433,N_2900,N_2993);
nand UO_434 (O_434,N_2992,N_2888);
or UO_435 (O_435,N_2953,N_2937);
xnor UO_436 (O_436,N_2861,N_2825);
and UO_437 (O_437,N_2823,N_2822);
or UO_438 (O_438,N_2970,N_2851);
and UO_439 (O_439,N_2893,N_2847);
nand UO_440 (O_440,N_2830,N_2948);
nor UO_441 (O_441,N_2903,N_2916);
or UO_442 (O_442,N_2939,N_2951);
nand UO_443 (O_443,N_2823,N_2957);
or UO_444 (O_444,N_2915,N_2911);
or UO_445 (O_445,N_2816,N_2969);
and UO_446 (O_446,N_2877,N_2866);
xnor UO_447 (O_447,N_2912,N_2982);
or UO_448 (O_448,N_2858,N_2856);
nor UO_449 (O_449,N_2995,N_2808);
nand UO_450 (O_450,N_2981,N_2801);
nor UO_451 (O_451,N_2919,N_2893);
nor UO_452 (O_452,N_2841,N_2905);
or UO_453 (O_453,N_2945,N_2867);
or UO_454 (O_454,N_2940,N_2992);
nand UO_455 (O_455,N_2998,N_2809);
and UO_456 (O_456,N_2804,N_2830);
nand UO_457 (O_457,N_2878,N_2888);
nor UO_458 (O_458,N_2963,N_2931);
and UO_459 (O_459,N_2893,N_2886);
and UO_460 (O_460,N_2958,N_2951);
and UO_461 (O_461,N_2900,N_2918);
or UO_462 (O_462,N_2822,N_2843);
and UO_463 (O_463,N_2884,N_2970);
or UO_464 (O_464,N_2850,N_2899);
xnor UO_465 (O_465,N_2830,N_2961);
nor UO_466 (O_466,N_2961,N_2902);
and UO_467 (O_467,N_2924,N_2809);
and UO_468 (O_468,N_2903,N_2800);
nor UO_469 (O_469,N_2856,N_2999);
or UO_470 (O_470,N_2926,N_2864);
and UO_471 (O_471,N_2885,N_2922);
or UO_472 (O_472,N_2905,N_2995);
or UO_473 (O_473,N_2897,N_2836);
nand UO_474 (O_474,N_2809,N_2801);
or UO_475 (O_475,N_2853,N_2886);
or UO_476 (O_476,N_2860,N_2925);
nand UO_477 (O_477,N_2964,N_2913);
and UO_478 (O_478,N_2879,N_2886);
nor UO_479 (O_479,N_2944,N_2960);
and UO_480 (O_480,N_2954,N_2855);
nand UO_481 (O_481,N_2942,N_2970);
nor UO_482 (O_482,N_2806,N_2962);
nor UO_483 (O_483,N_2925,N_2832);
nand UO_484 (O_484,N_2876,N_2909);
nor UO_485 (O_485,N_2934,N_2978);
and UO_486 (O_486,N_2811,N_2871);
and UO_487 (O_487,N_2873,N_2993);
xor UO_488 (O_488,N_2912,N_2864);
nand UO_489 (O_489,N_2827,N_2868);
nand UO_490 (O_490,N_2828,N_2887);
nand UO_491 (O_491,N_2919,N_2878);
nor UO_492 (O_492,N_2846,N_2916);
or UO_493 (O_493,N_2841,N_2986);
nand UO_494 (O_494,N_2936,N_2907);
nor UO_495 (O_495,N_2936,N_2811);
and UO_496 (O_496,N_2854,N_2926);
or UO_497 (O_497,N_2890,N_2864);
or UO_498 (O_498,N_2804,N_2906);
and UO_499 (O_499,N_2934,N_2816);
endmodule