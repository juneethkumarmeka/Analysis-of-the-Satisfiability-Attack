module basic_500_3000_500_3_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_454,In_492);
and U1 (N_1,In_154,In_251);
or U2 (N_2,In_243,In_128);
xnor U3 (N_3,In_194,In_377);
or U4 (N_4,In_350,In_408);
or U5 (N_5,In_294,In_139);
or U6 (N_6,In_233,In_435);
nand U7 (N_7,In_257,In_478);
nand U8 (N_8,In_415,In_145);
and U9 (N_9,In_115,In_4);
nand U10 (N_10,In_354,In_467);
and U11 (N_11,In_369,In_453);
nor U12 (N_12,In_353,In_303);
nor U13 (N_13,In_304,In_44);
xor U14 (N_14,In_308,In_281);
nor U15 (N_15,In_211,In_288);
and U16 (N_16,In_252,In_168);
nor U17 (N_17,In_360,In_3);
or U18 (N_18,In_229,In_12);
nand U19 (N_19,In_420,In_30);
xor U20 (N_20,In_23,In_10);
nand U21 (N_21,In_374,In_334);
or U22 (N_22,In_276,In_287);
and U23 (N_23,In_269,In_410);
xor U24 (N_24,In_56,In_385);
or U25 (N_25,In_275,In_62);
nand U26 (N_26,In_297,In_476);
or U27 (N_27,In_51,In_307);
xor U28 (N_28,In_480,In_31);
nand U29 (N_29,In_73,In_326);
nor U30 (N_30,In_47,In_365);
and U31 (N_31,In_298,In_392);
or U32 (N_32,In_80,In_263);
xor U33 (N_33,In_412,In_310);
nor U34 (N_34,In_177,In_498);
xor U35 (N_35,In_125,In_0);
nor U36 (N_36,In_235,In_173);
or U37 (N_37,In_126,In_349);
and U38 (N_38,In_259,In_7);
nand U39 (N_39,In_239,In_367);
nand U40 (N_40,In_25,In_40);
or U41 (N_41,In_371,In_38);
nor U42 (N_42,In_430,In_496);
or U43 (N_43,In_195,In_84);
xor U44 (N_44,In_19,In_336);
nor U45 (N_45,In_449,In_351);
and U46 (N_46,In_277,In_149);
and U47 (N_47,In_245,In_99);
nand U48 (N_48,In_335,In_213);
nand U49 (N_49,In_104,In_98);
or U50 (N_50,In_322,In_345);
and U51 (N_51,In_90,In_438);
nand U52 (N_52,In_300,In_387);
nor U53 (N_53,In_272,In_469);
or U54 (N_54,In_198,In_58);
nor U55 (N_55,In_89,In_83);
nand U56 (N_56,In_162,In_112);
and U57 (N_57,In_301,In_455);
and U58 (N_58,In_127,In_103);
nor U59 (N_59,In_376,In_53);
and U60 (N_60,In_343,In_161);
and U61 (N_61,In_232,In_241);
or U62 (N_62,In_65,In_129);
nor U63 (N_63,In_339,In_186);
nand U64 (N_64,In_486,In_429);
and U65 (N_65,In_144,In_366);
xor U66 (N_66,In_111,In_383);
or U67 (N_67,In_290,In_416);
nand U68 (N_68,In_156,In_167);
nor U69 (N_69,In_442,In_33);
or U70 (N_70,In_215,In_197);
nor U71 (N_71,In_78,In_372);
and U72 (N_72,In_400,In_95);
nand U73 (N_73,In_2,In_439);
nor U74 (N_74,In_222,In_337);
nand U75 (N_75,In_52,In_255);
and U76 (N_76,In_75,In_118);
nand U77 (N_77,In_176,In_234);
xor U78 (N_78,In_179,In_148);
and U79 (N_79,In_175,In_192);
and U80 (N_80,In_274,In_218);
xnor U81 (N_81,In_483,In_368);
nand U82 (N_82,In_42,In_158);
or U83 (N_83,In_169,In_36);
and U84 (N_84,In_137,In_85);
nor U85 (N_85,In_153,In_187);
or U86 (N_86,In_191,In_221);
nand U87 (N_87,In_100,In_352);
xor U88 (N_88,In_97,In_423);
nand U89 (N_89,In_379,In_163);
and U90 (N_90,In_384,In_133);
nand U91 (N_91,In_27,In_450);
xor U92 (N_92,In_338,In_39);
nor U93 (N_93,In_87,In_481);
or U94 (N_94,In_451,In_487);
or U95 (N_95,In_463,In_43);
and U96 (N_96,In_214,In_131);
nand U97 (N_97,In_50,In_160);
and U98 (N_98,In_204,In_182);
and U99 (N_99,In_15,In_254);
nor U100 (N_100,In_348,In_452);
nor U101 (N_101,In_74,In_475);
nand U102 (N_102,In_291,In_240);
xor U103 (N_103,In_93,In_421);
and U104 (N_104,In_292,In_230);
nor U105 (N_105,In_437,In_142);
nor U106 (N_106,In_1,In_344);
or U107 (N_107,In_262,In_200);
nand U108 (N_108,In_238,In_306);
nand U109 (N_109,In_431,In_157);
or U110 (N_110,In_271,In_361);
xnor U111 (N_111,In_325,In_35);
nor U112 (N_112,In_305,In_462);
nor U113 (N_113,In_426,In_121);
and U114 (N_114,In_331,In_69);
and U115 (N_115,In_286,In_120);
and U116 (N_116,In_249,In_67);
or U117 (N_117,In_296,In_72);
and U118 (N_118,In_18,In_318);
nand U119 (N_119,In_401,In_236);
or U120 (N_120,In_293,In_491);
and U121 (N_121,In_468,In_440);
nor U122 (N_122,In_405,In_356);
nor U123 (N_123,In_201,In_273);
and U124 (N_124,In_242,In_409);
nand U125 (N_125,In_268,In_364);
nand U126 (N_126,In_116,In_295);
nor U127 (N_127,In_22,In_330);
and U128 (N_128,In_311,In_494);
nand U129 (N_129,In_285,In_185);
nand U130 (N_130,In_5,In_282);
or U131 (N_131,In_323,In_267);
nor U132 (N_132,In_28,In_414);
xnor U133 (N_133,In_81,In_147);
nand U134 (N_134,In_382,In_122);
xor U135 (N_135,In_219,In_224);
or U136 (N_136,In_46,In_444);
nand U137 (N_137,In_474,In_477);
nand U138 (N_138,In_391,In_208);
nand U139 (N_139,In_457,In_495);
nand U140 (N_140,In_403,In_102);
and U141 (N_141,In_203,In_63);
nand U142 (N_142,In_394,In_212);
xor U143 (N_143,In_346,In_178);
or U144 (N_144,In_256,In_425);
or U145 (N_145,In_398,In_433);
nand U146 (N_146,In_375,In_270);
xnor U147 (N_147,In_280,In_166);
xnor U148 (N_148,In_370,In_159);
nand U149 (N_149,In_332,In_493);
nand U150 (N_150,In_109,In_210);
nor U151 (N_151,In_471,In_54);
nand U152 (N_152,In_217,In_59);
nor U153 (N_153,In_283,In_315);
nor U154 (N_154,In_94,In_473);
nor U155 (N_155,In_101,In_181);
and U156 (N_156,In_319,In_258);
or U157 (N_157,In_441,In_316);
or U158 (N_158,In_373,In_49);
or U159 (N_159,In_406,In_165);
or U160 (N_160,In_328,In_150);
and U161 (N_161,In_261,In_151);
nor U162 (N_162,In_207,In_199);
and U163 (N_163,In_13,In_180);
or U164 (N_164,In_289,In_60);
and U165 (N_165,In_279,In_174);
nand U166 (N_166,In_34,In_189);
or U167 (N_167,In_246,In_14);
xor U168 (N_168,In_313,In_223);
xor U169 (N_169,In_489,In_184);
xor U170 (N_170,In_340,In_458);
or U171 (N_171,In_11,In_193);
nor U172 (N_172,In_393,In_237);
and U173 (N_173,In_183,In_41);
or U174 (N_174,In_45,In_17);
or U175 (N_175,In_432,In_299);
nor U176 (N_176,In_357,In_260);
xnor U177 (N_177,In_446,In_29);
nand U178 (N_178,In_266,In_143);
and U179 (N_179,In_76,In_397);
or U180 (N_180,In_472,In_170);
nand U181 (N_181,In_264,In_381);
nand U182 (N_182,In_106,In_404);
and U183 (N_183,In_314,In_228);
nand U184 (N_184,In_427,In_284);
or U185 (N_185,In_8,In_302);
nor U186 (N_186,In_16,In_21);
nor U187 (N_187,In_390,In_466);
or U188 (N_188,In_77,In_464);
nand U189 (N_189,In_92,In_138);
nor U190 (N_190,In_359,In_231);
xnor U191 (N_191,In_309,In_113);
and U192 (N_192,In_134,In_119);
nor U193 (N_193,In_497,In_362);
and U194 (N_194,In_465,In_55);
or U195 (N_195,In_188,In_342);
nand U196 (N_196,In_399,In_171);
and U197 (N_197,In_26,In_490);
and U198 (N_198,In_135,In_424);
nand U199 (N_199,In_61,In_389);
nand U200 (N_200,In_155,In_378);
and U201 (N_201,In_205,In_460);
nor U202 (N_202,In_419,In_312);
nand U203 (N_203,In_244,In_220);
and U204 (N_204,In_459,In_448);
and U205 (N_205,In_411,In_88);
or U206 (N_206,In_417,In_402);
or U207 (N_207,In_434,In_68);
nand U208 (N_208,In_445,In_253);
and U209 (N_209,In_140,In_324);
nand U210 (N_210,In_443,In_422);
nand U211 (N_211,In_79,In_202);
and U212 (N_212,In_82,In_132);
nor U213 (N_213,In_57,In_436);
or U214 (N_214,In_114,In_248);
nand U215 (N_215,In_190,In_482);
nand U216 (N_216,In_456,In_70);
nor U217 (N_217,In_428,In_152);
or U218 (N_218,In_136,In_164);
and U219 (N_219,In_321,In_363);
nand U220 (N_220,In_278,In_407);
and U221 (N_221,In_447,In_48);
nand U222 (N_222,In_146,In_333);
xor U223 (N_223,In_485,In_6);
nand U224 (N_224,In_380,In_24);
xor U225 (N_225,In_206,In_250);
or U226 (N_226,In_358,In_227);
xnor U227 (N_227,In_327,In_386);
and U228 (N_228,In_124,In_172);
or U229 (N_229,In_225,In_32);
or U230 (N_230,In_317,In_395);
nor U231 (N_231,In_107,In_108);
and U232 (N_232,In_499,In_123);
and U233 (N_233,In_91,In_110);
nand U234 (N_234,In_141,In_265);
nand U235 (N_235,In_355,In_461);
or U236 (N_236,In_64,In_396);
and U237 (N_237,In_479,In_71);
and U238 (N_238,In_226,In_86);
xor U239 (N_239,In_105,In_20);
nor U240 (N_240,In_196,In_470);
or U241 (N_241,In_66,In_388);
and U242 (N_242,In_320,In_418);
and U243 (N_243,In_130,In_37);
and U244 (N_244,In_209,In_347);
and U245 (N_245,In_484,In_329);
and U246 (N_246,In_216,In_488);
nand U247 (N_247,In_413,In_9);
and U248 (N_248,In_96,In_117);
and U249 (N_249,In_247,In_341);
nor U250 (N_250,In_192,In_334);
or U251 (N_251,In_321,In_246);
xnor U252 (N_252,In_260,In_34);
and U253 (N_253,In_366,In_229);
or U254 (N_254,In_107,In_376);
nand U255 (N_255,In_210,In_185);
nor U256 (N_256,In_46,In_60);
nor U257 (N_257,In_457,In_151);
nand U258 (N_258,In_85,In_261);
nand U259 (N_259,In_87,In_152);
or U260 (N_260,In_182,In_200);
xor U261 (N_261,In_246,In_82);
or U262 (N_262,In_336,In_160);
xor U263 (N_263,In_486,In_337);
or U264 (N_264,In_458,In_152);
or U265 (N_265,In_230,In_61);
nor U266 (N_266,In_130,In_31);
nand U267 (N_267,In_260,In_27);
nor U268 (N_268,In_72,In_168);
nor U269 (N_269,In_389,In_145);
nor U270 (N_270,In_223,In_328);
nand U271 (N_271,In_241,In_366);
nand U272 (N_272,In_123,In_290);
nand U273 (N_273,In_426,In_218);
or U274 (N_274,In_494,In_137);
and U275 (N_275,In_75,In_434);
or U276 (N_276,In_246,In_12);
nand U277 (N_277,In_36,In_487);
or U278 (N_278,In_272,In_39);
or U279 (N_279,In_456,In_186);
or U280 (N_280,In_127,In_259);
and U281 (N_281,In_75,In_404);
nor U282 (N_282,In_350,In_378);
or U283 (N_283,In_81,In_465);
nand U284 (N_284,In_147,In_207);
nor U285 (N_285,In_371,In_63);
nor U286 (N_286,In_211,In_178);
nor U287 (N_287,In_310,In_357);
and U288 (N_288,In_163,In_181);
and U289 (N_289,In_179,In_7);
nor U290 (N_290,In_421,In_180);
and U291 (N_291,In_22,In_403);
and U292 (N_292,In_468,In_206);
nand U293 (N_293,In_474,In_329);
or U294 (N_294,In_22,In_203);
nand U295 (N_295,In_213,In_278);
or U296 (N_296,In_186,In_459);
and U297 (N_297,In_42,In_271);
nand U298 (N_298,In_157,In_381);
or U299 (N_299,In_61,In_287);
or U300 (N_300,In_496,In_171);
nor U301 (N_301,In_261,In_316);
and U302 (N_302,In_310,In_117);
xor U303 (N_303,In_261,In_122);
or U304 (N_304,In_355,In_460);
or U305 (N_305,In_406,In_482);
nor U306 (N_306,In_165,In_335);
xnor U307 (N_307,In_358,In_273);
and U308 (N_308,In_427,In_198);
nand U309 (N_309,In_466,In_116);
xnor U310 (N_310,In_81,In_38);
and U311 (N_311,In_219,In_157);
or U312 (N_312,In_23,In_280);
and U313 (N_313,In_195,In_191);
nor U314 (N_314,In_484,In_399);
xor U315 (N_315,In_238,In_175);
and U316 (N_316,In_33,In_395);
or U317 (N_317,In_462,In_336);
xor U318 (N_318,In_78,In_299);
xnor U319 (N_319,In_233,In_425);
or U320 (N_320,In_48,In_5);
and U321 (N_321,In_34,In_210);
nor U322 (N_322,In_161,In_386);
nand U323 (N_323,In_54,In_258);
nor U324 (N_324,In_380,In_304);
xor U325 (N_325,In_318,In_316);
nand U326 (N_326,In_137,In_422);
and U327 (N_327,In_154,In_151);
nor U328 (N_328,In_272,In_236);
or U329 (N_329,In_95,In_317);
or U330 (N_330,In_315,In_371);
nand U331 (N_331,In_459,In_306);
or U332 (N_332,In_413,In_143);
nor U333 (N_333,In_206,In_111);
xor U334 (N_334,In_352,In_61);
nor U335 (N_335,In_446,In_416);
xor U336 (N_336,In_286,In_96);
or U337 (N_337,In_127,In_134);
xnor U338 (N_338,In_208,In_448);
nand U339 (N_339,In_382,In_306);
nand U340 (N_340,In_61,In_450);
nand U341 (N_341,In_190,In_360);
and U342 (N_342,In_473,In_264);
or U343 (N_343,In_264,In_146);
nor U344 (N_344,In_143,In_280);
or U345 (N_345,In_246,In_263);
nand U346 (N_346,In_284,In_494);
xnor U347 (N_347,In_262,In_323);
or U348 (N_348,In_181,In_94);
nand U349 (N_349,In_146,In_68);
and U350 (N_350,In_122,In_117);
or U351 (N_351,In_463,In_310);
nor U352 (N_352,In_370,In_4);
or U353 (N_353,In_164,In_33);
xor U354 (N_354,In_235,In_392);
and U355 (N_355,In_386,In_242);
or U356 (N_356,In_299,In_20);
and U357 (N_357,In_236,In_233);
xor U358 (N_358,In_216,In_19);
xor U359 (N_359,In_137,In_327);
nand U360 (N_360,In_3,In_352);
and U361 (N_361,In_300,In_475);
nand U362 (N_362,In_127,In_8);
nand U363 (N_363,In_49,In_231);
xor U364 (N_364,In_52,In_379);
nand U365 (N_365,In_132,In_467);
nor U366 (N_366,In_203,In_91);
nor U367 (N_367,In_489,In_371);
nor U368 (N_368,In_101,In_254);
and U369 (N_369,In_410,In_45);
or U370 (N_370,In_131,In_413);
nor U371 (N_371,In_59,In_219);
or U372 (N_372,In_161,In_139);
nor U373 (N_373,In_161,In_381);
xnor U374 (N_374,In_265,In_401);
or U375 (N_375,In_291,In_7);
nor U376 (N_376,In_77,In_184);
and U377 (N_377,In_394,In_337);
nand U378 (N_378,In_23,In_1);
nand U379 (N_379,In_270,In_84);
and U380 (N_380,In_322,In_343);
nor U381 (N_381,In_369,In_4);
nand U382 (N_382,In_146,In_99);
nand U383 (N_383,In_309,In_258);
and U384 (N_384,In_365,In_422);
nand U385 (N_385,In_444,In_481);
or U386 (N_386,In_190,In_445);
nand U387 (N_387,In_235,In_399);
nand U388 (N_388,In_321,In_113);
nand U389 (N_389,In_274,In_488);
and U390 (N_390,In_358,In_181);
nor U391 (N_391,In_289,In_175);
nand U392 (N_392,In_421,In_92);
or U393 (N_393,In_83,In_218);
nor U394 (N_394,In_298,In_376);
or U395 (N_395,In_99,In_371);
or U396 (N_396,In_120,In_449);
nor U397 (N_397,In_56,In_316);
nand U398 (N_398,In_24,In_31);
or U399 (N_399,In_292,In_98);
nor U400 (N_400,In_29,In_275);
nand U401 (N_401,In_423,In_229);
nand U402 (N_402,In_76,In_159);
nor U403 (N_403,In_235,In_328);
nor U404 (N_404,In_448,In_340);
nand U405 (N_405,In_239,In_338);
nor U406 (N_406,In_455,In_268);
nand U407 (N_407,In_42,In_60);
or U408 (N_408,In_233,In_348);
and U409 (N_409,In_32,In_101);
xnor U410 (N_410,In_39,In_109);
nor U411 (N_411,In_294,In_490);
nand U412 (N_412,In_429,In_131);
nand U413 (N_413,In_490,In_4);
or U414 (N_414,In_98,In_497);
nor U415 (N_415,In_99,In_493);
nand U416 (N_416,In_57,In_375);
nand U417 (N_417,In_212,In_259);
and U418 (N_418,In_361,In_256);
nor U419 (N_419,In_189,In_408);
nand U420 (N_420,In_409,In_235);
and U421 (N_421,In_395,In_459);
or U422 (N_422,In_277,In_106);
and U423 (N_423,In_311,In_165);
nor U424 (N_424,In_317,In_434);
nand U425 (N_425,In_278,In_198);
nor U426 (N_426,In_116,In_385);
nor U427 (N_427,In_319,In_123);
nor U428 (N_428,In_217,In_454);
nor U429 (N_429,In_162,In_24);
nor U430 (N_430,In_140,In_371);
or U431 (N_431,In_125,In_308);
xor U432 (N_432,In_182,In_83);
nor U433 (N_433,In_470,In_249);
nor U434 (N_434,In_100,In_239);
nor U435 (N_435,In_273,In_345);
xor U436 (N_436,In_156,In_385);
or U437 (N_437,In_426,In_443);
nor U438 (N_438,In_307,In_230);
nor U439 (N_439,In_83,In_104);
or U440 (N_440,In_81,In_477);
or U441 (N_441,In_415,In_122);
and U442 (N_442,In_359,In_28);
nand U443 (N_443,In_315,In_417);
or U444 (N_444,In_81,In_372);
nand U445 (N_445,In_295,In_303);
and U446 (N_446,In_192,In_187);
or U447 (N_447,In_195,In_149);
nand U448 (N_448,In_328,In_290);
or U449 (N_449,In_377,In_190);
or U450 (N_450,In_257,In_217);
nand U451 (N_451,In_50,In_397);
nor U452 (N_452,In_12,In_131);
xor U453 (N_453,In_201,In_136);
nor U454 (N_454,In_437,In_53);
xnor U455 (N_455,In_87,In_494);
nor U456 (N_456,In_108,In_67);
xor U457 (N_457,In_62,In_493);
and U458 (N_458,In_466,In_483);
nand U459 (N_459,In_379,In_231);
or U460 (N_460,In_200,In_165);
nor U461 (N_461,In_369,In_234);
xor U462 (N_462,In_266,In_289);
or U463 (N_463,In_306,In_27);
nand U464 (N_464,In_432,In_307);
or U465 (N_465,In_32,In_14);
nand U466 (N_466,In_375,In_320);
or U467 (N_467,In_64,In_341);
or U468 (N_468,In_40,In_346);
nand U469 (N_469,In_484,In_177);
or U470 (N_470,In_476,In_77);
nand U471 (N_471,In_117,In_143);
or U472 (N_472,In_357,In_322);
nor U473 (N_473,In_67,In_496);
nor U474 (N_474,In_138,In_93);
nand U475 (N_475,In_181,In_488);
nand U476 (N_476,In_363,In_32);
nor U477 (N_477,In_128,In_223);
or U478 (N_478,In_53,In_348);
nand U479 (N_479,In_319,In_115);
nand U480 (N_480,In_461,In_71);
xnor U481 (N_481,In_374,In_18);
or U482 (N_482,In_488,In_320);
nand U483 (N_483,In_395,In_38);
or U484 (N_484,In_295,In_86);
nor U485 (N_485,In_212,In_336);
nor U486 (N_486,In_167,In_134);
nand U487 (N_487,In_242,In_413);
nor U488 (N_488,In_27,In_100);
or U489 (N_489,In_50,In_319);
nand U490 (N_490,In_305,In_495);
and U491 (N_491,In_315,In_179);
or U492 (N_492,In_183,In_139);
nor U493 (N_493,In_22,In_499);
and U494 (N_494,In_90,In_270);
xor U495 (N_495,In_299,In_280);
or U496 (N_496,In_151,In_323);
nand U497 (N_497,In_254,In_194);
and U498 (N_498,In_281,In_100);
and U499 (N_499,In_90,In_20);
nor U500 (N_500,In_249,In_79);
nor U501 (N_501,In_300,In_48);
and U502 (N_502,In_353,In_275);
nor U503 (N_503,In_414,In_104);
or U504 (N_504,In_309,In_99);
and U505 (N_505,In_144,In_421);
xor U506 (N_506,In_210,In_217);
and U507 (N_507,In_37,In_181);
nand U508 (N_508,In_306,In_318);
and U509 (N_509,In_283,In_80);
nor U510 (N_510,In_318,In_482);
or U511 (N_511,In_148,In_340);
and U512 (N_512,In_415,In_61);
nor U513 (N_513,In_131,In_419);
nand U514 (N_514,In_441,In_429);
nand U515 (N_515,In_25,In_119);
and U516 (N_516,In_422,In_249);
and U517 (N_517,In_194,In_478);
nor U518 (N_518,In_148,In_407);
and U519 (N_519,In_292,In_109);
or U520 (N_520,In_176,In_486);
or U521 (N_521,In_237,In_406);
xor U522 (N_522,In_133,In_74);
or U523 (N_523,In_182,In_328);
nand U524 (N_524,In_99,In_499);
nand U525 (N_525,In_365,In_300);
and U526 (N_526,In_109,In_368);
nor U527 (N_527,In_478,In_53);
nand U528 (N_528,In_199,In_161);
nor U529 (N_529,In_21,In_79);
and U530 (N_530,In_412,In_253);
and U531 (N_531,In_392,In_409);
nand U532 (N_532,In_74,In_55);
or U533 (N_533,In_398,In_428);
nor U534 (N_534,In_11,In_33);
nand U535 (N_535,In_462,In_30);
or U536 (N_536,In_396,In_401);
and U537 (N_537,In_268,In_243);
xnor U538 (N_538,In_234,In_168);
and U539 (N_539,In_181,In_36);
nor U540 (N_540,In_377,In_429);
or U541 (N_541,In_280,In_427);
or U542 (N_542,In_247,In_277);
or U543 (N_543,In_198,In_71);
nand U544 (N_544,In_256,In_490);
or U545 (N_545,In_380,In_449);
or U546 (N_546,In_348,In_237);
and U547 (N_547,In_107,In_54);
or U548 (N_548,In_343,In_414);
and U549 (N_549,In_62,In_96);
nand U550 (N_550,In_143,In_438);
xor U551 (N_551,In_308,In_411);
nor U552 (N_552,In_158,In_279);
and U553 (N_553,In_396,In_467);
or U554 (N_554,In_245,In_328);
xnor U555 (N_555,In_22,In_491);
and U556 (N_556,In_49,In_355);
nor U557 (N_557,In_77,In_297);
or U558 (N_558,In_258,In_494);
nor U559 (N_559,In_358,In_447);
nor U560 (N_560,In_269,In_95);
and U561 (N_561,In_439,In_195);
nor U562 (N_562,In_197,In_179);
and U563 (N_563,In_181,In_413);
nor U564 (N_564,In_319,In_384);
and U565 (N_565,In_439,In_383);
nand U566 (N_566,In_77,In_136);
nor U567 (N_567,In_424,In_390);
nand U568 (N_568,In_79,In_186);
nand U569 (N_569,In_298,In_439);
xor U570 (N_570,In_440,In_89);
or U571 (N_571,In_372,In_150);
nand U572 (N_572,In_481,In_345);
xnor U573 (N_573,In_253,In_233);
nor U574 (N_574,In_306,In_399);
or U575 (N_575,In_28,In_272);
nor U576 (N_576,In_384,In_132);
or U577 (N_577,In_465,In_32);
nand U578 (N_578,In_58,In_311);
and U579 (N_579,In_76,In_423);
or U580 (N_580,In_266,In_328);
and U581 (N_581,In_318,In_60);
nor U582 (N_582,In_466,In_342);
nand U583 (N_583,In_291,In_246);
nand U584 (N_584,In_162,In_168);
nor U585 (N_585,In_396,In_48);
nor U586 (N_586,In_366,In_314);
or U587 (N_587,In_409,In_196);
nand U588 (N_588,In_428,In_16);
nand U589 (N_589,In_437,In_271);
nor U590 (N_590,In_111,In_392);
nand U591 (N_591,In_214,In_243);
or U592 (N_592,In_291,In_266);
and U593 (N_593,In_201,In_156);
nor U594 (N_594,In_75,In_371);
and U595 (N_595,In_272,In_263);
and U596 (N_596,In_24,In_352);
or U597 (N_597,In_230,In_421);
and U598 (N_598,In_401,In_162);
nor U599 (N_599,In_297,In_293);
nor U600 (N_600,In_289,In_192);
nor U601 (N_601,In_409,In_161);
and U602 (N_602,In_45,In_1);
nor U603 (N_603,In_210,In_26);
nor U604 (N_604,In_425,In_390);
nor U605 (N_605,In_110,In_365);
nand U606 (N_606,In_406,In_124);
nand U607 (N_607,In_124,In_185);
nand U608 (N_608,In_143,In_393);
or U609 (N_609,In_29,In_244);
and U610 (N_610,In_27,In_438);
and U611 (N_611,In_240,In_446);
nor U612 (N_612,In_490,In_428);
nor U613 (N_613,In_194,In_21);
nor U614 (N_614,In_294,In_415);
and U615 (N_615,In_332,In_398);
nor U616 (N_616,In_354,In_191);
and U617 (N_617,In_496,In_207);
nor U618 (N_618,In_222,In_394);
and U619 (N_619,In_287,In_201);
nor U620 (N_620,In_165,In_22);
or U621 (N_621,In_10,In_441);
or U622 (N_622,In_328,In_126);
nor U623 (N_623,In_274,In_242);
nor U624 (N_624,In_20,In_68);
nand U625 (N_625,In_117,In_409);
nand U626 (N_626,In_122,In_344);
nor U627 (N_627,In_239,In_417);
nor U628 (N_628,In_130,In_279);
and U629 (N_629,In_286,In_236);
or U630 (N_630,In_27,In_7);
and U631 (N_631,In_21,In_366);
xnor U632 (N_632,In_469,In_244);
and U633 (N_633,In_354,In_382);
and U634 (N_634,In_240,In_253);
xnor U635 (N_635,In_338,In_7);
or U636 (N_636,In_434,In_350);
nor U637 (N_637,In_460,In_449);
xnor U638 (N_638,In_73,In_312);
and U639 (N_639,In_311,In_189);
nand U640 (N_640,In_350,In_110);
xor U641 (N_641,In_442,In_373);
nand U642 (N_642,In_466,In_91);
nand U643 (N_643,In_121,In_275);
xnor U644 (N_644,In_264,In_494);
nand U645 (N_645,In_404,In_171);
and U646 (N_646,In_448,In_96);
and U647 (N_647,In_491,In_66);
and U648 (N_648,In_112,In_321);
nand U649 (N_649,In_18,In_224);
nand U650 (N_650,In_369,In_80);
nor U651 (N_651,In_191,In_459);
and U652 (N_652,In_227,In_431);
nand U653 (N_653,In_280,In_204);
and U654 (N_654,In_313,In_260);
and U655 (N_655,In_87,In_256);
nor U656 (N_656,In_339,In_167);
nand U657 (N_657,In_392,In_80);
nand U658 (N_658,In_254,In_110);
nor U659 (N_659,In_79,In_55);
xor U660 (N_660,In_491,In_414);
and U661 (N_661,In_335,In_169);
or U662 (N_662,In_227,In_293);
nor U663 (N_663,In_287,In_378);
nor U664 (N_664,In_72,In_399);
or U665 (N_665,In_423,In_149);
nand U666 (N_666,In_162,In_141);
or U667 (N_667,In_455,In_155);
xor U668 (N_668,In_306,In_245);
nand U669 (N_669,In_285,In_238);
nor U670 (N_670,In_210,In_220);
nor U671 (N_671,In_151,In_10);
nand U672 (N_672,In_156,In_175);
nor U673 (N_673,In_103,In_141);
nand U674 (N_674,In_453,In_164);
or U675 (N_675,In_101,In_351);
nand U676 (N_676,In_283,In_157);
nand U677 (N_677,In_13,In_87);
nor U678 (N_678,In_290,In_468);
nor U679 (N_679,In_454,In_429);
nor U680 (N_680,In_69,In_287);
or U681 (N_681,In_327,In_38);
nor U682 (N_682,In_360,In_402);
nor U683 (N_683,In_122,In_265);
or U684 (N_684,In_473,In_208);
nand U685 (N_685,In_412,In_295);
nand U686 (N_686,In_253,In_205);
nor U687 (N_687,In_288,In_415);
or U688 (N_688,In_465,In_345);
nand U689 (N_689,In_8,In_102);
nand U690 (N_690,In_64,In_143);
xnor U691 (N_691,In_213,In_96);
or U692 (N_692,In_480,In_343);
nand U693 (N_693,In_115,In_77);
or U694 (N_694,In_11,In_212);
or U695 (N_695,In_456,In_60);
xnor U696 (N_696,In_198,In_193);
or U697 (N_697,In_238,In_288);
nand U698 (N_698,In_95,In_92);
or U699 (N_699,In_429,In_483);
nand U700 (N_700,In_309,In_42);
or U701 (N_701,In_341,In_408);
xnor U702 (N_702,In_166,In_466);
xor U703 (N_703,In_75,In_357);
nand U704 (N_704,In_321,In_362);
or U705 (N_705,In_90,In_203);
and U706 (N_706,In_129,In_66);
or U707 (N_707,In_356,In_434);
or U708 (N_708,In_85,In_240);
xnor U709 (N_709,In_90,In_399);
nand U710 (N_710,In_236,In_347);
nor U711 (N_711,In_199,In_91);
or U712 (N_712,In_97,In_401);
nand U713 (N_713,In_322,In_417);
nor U714 (N_714,In_134,In_122);
or U715 (N_715,In_391,In_68);
xnor U716 (N_716,In_208,In_394);
and U717 (N_717,In_458,In_270);
nor U718 (N_718,In_141,In_145);
or U719 (N_719,In_244,In_468);
and U720 (N_720,In_323,In_244);
nor U721 (N_721,In_486,In_38);
nor U722 (N_722,In_102,In_340);
nand U723 (N_723,In_72,In_25);
and U724 (N_724,In_458,In_312);
and U725 (N_725,In_43,In_437);
xor U726 (N_726,In_368,In_153);
nor U727 (N_727,In_365,In_167);
nor U728 (N_728,In_147,In_401);
and U729 (N_729,In_97,In_46);
and U730 (N_730,In_251,In_480);
or U731 (N_731,In_257,In_107);
or U732 (N_732,In_100,In_198);
nor U733 (N_733,In_447,In_214);
nor U734 (N_734,In_129,In_452);
and U735 (N_735,In_116,In_494);
xnor U736 (N_736,In_60,In_189);
or U737 (N_737,In_145,In_208);
or U738 (N_738,In_365,In_359);
and U739 (N_739,In_21,In_62);
nor U740 (N_740,In_391,In_124);
xnor U741 (N_741,In_359,In_213);
nor U742 (N_742,In_97,In_472);
xor U743 (N_743,In_436,In_80);
and U744 (N_744,In_373,In_162);
xor U745 (N_745,In_48,In_382);
and U746 (N_746,In_110,In_143);
nand U747 (N_747,In_44,In_26);
and U748 (N_748,In_90,In_392);
xor U749 (N_749,In_302,In_400);
or U750 (N_750,In_110,In_342);
or U751 (N_751,In_48,In_102);
or U752 (N_752,In_278,In_369);
or U753 (N_753,In_212,In_196);
nor U754 (N_754,In_370,In_105);
nor U755 (N_755,In_98,In_51);
and U756 (N_756,In_396,In_218);
nand U757 (N_757,In_441,In_162);
or U758 (N_758,In_298,In_20);
and U759 (N_759,In_397,In_121);
nor U760 (N_760,In_328,In_370);
nand U761 (N_761,In_496,In_122);
nand U762 (N_762,In_256,In_345);
nand U763 (N_763,In_354,In_408);
nand U764 (N_764,In_391,In_202);
nand U765 (N_765,In_284,In_210);
or U766 (N_766,In_26,In_432);
nand U767 (N_767,In_294,In_457);
and U768 (N_768,In_54,In_406);
or U769 (N_769,In_90,In_235);
nand U770 (N_770,In_499,In_490);
and U771 (N_771,In_464,In_416);
or U772 (N_772,In_422,In_184);
nand U773 (N_773,In_337,In_261);
and U774 (N_774,In_132,In_25);
nor U775 (N_775,In_240,In_357);
xnor U776 (N_776,In_60,In_201);
nor U777 (N_777,In_270,In_413);
and U778 (N_778,In_440,In_404);
or U779 (N_779,In_136,In_413);
nor U780 (N_780,In_244,In_90);
nand U781 (N_781,In_164,In_42);
or U782 (N_782,In_392,In_215);
and U783 (N_783,In_386,In_375);
and U784 (N_784,In_311,In_135);
and U785 (N_785,In_109,In_157);
nand U786 (N_786,In_22,In_35);
or U787 (N_787,In_325,In_150);
or U788 (N_788,In_224,In_242);
xnor U789 (N_789,In_489,In_370);
nand U790 (N_790,In_464,In_173);
and U791 (N_791,In_286,In_140);
nor U792 (N_792,In_417,In_2);
or U793 (N_793,In_403,In_18);
nand U794 (N_794,In_96,In_250);
and U795 (N_795,In_349,In_274);
nand U796 (N_796,In_184,In_173);
nand U797 (N_797,In_433,In_73);
or U798 (N_798,In_333,In_272);
and U799 (N_799,In_186,In_164);
nor U800 (N_800,In_400,In_147);
nand U801 (N_801,In_242,In_194);
and U802 (N_802,In_273,In_311);
and U803 (N_803,In_259,In_191);
or U804 (N_804,In_115,In_239);
nor U805 (N_805,In_253,In_485);
and U806 (N_806,In_441,In_22);
or U807 (N_807,In_413,In_219);
and U808 (N_808,In_70,In_234);
or U809 (N_809,In_68,In_194);
or U810 (N_810,In_447,In_18);
nor U811 (N_811,In_232,In_464);
and U812 (N_812,In_35,In_317);
or U813 (N_813,In_163,In_339);
nand U814 (N_814,In_461,In_277);
or U815 (N_815,In_121,In_128);
nor U816 (N_816,In_359,In_382);
or U817 (N_817,In_133,In_130);
nor U818 (N_818,In_297,In_217);
or U819 (N_819,In_257,In_230);
xnor U820 (N_820,In_275,In_392);
xnor U821 (N_821,In_177,In_494);
and U822 (N_822,In_245,In_138);
and U823 (N_823,In_274,In_161);
nand U824 (N_824,In_74,In_223);
nand U825 (N_825,In_207,In_201);
nor U826 (N_826,In_90,In_207);
nand U827 (N_827,In_146,In_29);
nor U828 (N_828,In_486,In_431);
or U829 (N_829,In_218,In_353);
nor U830 (N_830,In_319,In_70);
nor U831 (N_831,In_406,In_7);
nand U832 (N_832,In_250,In_325);
nor U833 (N_833,In_68,In_71);
or U834 (N_834,In_386,In_143);
and U835 (N_835,In_262,In_102);
or U836 (N_836,In_260,In_151);
or U837 (N_837,In_29,In_380);
or U838 (N_838,In_70,In_359);
and U839 (N_839,In_257,In_452);
and U840 (N_840,In_471,In_155);
nor U841 (N_841,In_270,In_179);
and U842 (N_842,In_296,In_249);
and U843 (N_843,In_211,In_169);
and U844 (N_844,In_155,In_460);
and U845 (N_845,In_223,In_414);
or U846 (N_846,In_313,In_200);
nor U847 (N_847,In_444,In_166);
nand U848 (N_848,In_458,In_364);
or U849 (N_849,In_36,In_175);
nand U850 (N_850,In_484,In_30);
and U851 (N_851,In_117,In_218);
nand U852 (N_852,In_290,In_422);
and U853 (N_853,In_419,In_149);
or U854 (N_854,In_97,In_200);
nand U855 (N_855,In_374,In_494);
or U856 (N_856,In_369,In_249);
xnor U857 (N_857,In_139,In_57);
or U858 (N_858,In_197,In_294);
nor U859 (N_859,In_129,In_472);
nor U860 (N_860,In_19,In_90);
and U861 (N_861,In_247,In_147);
and U862 (N_862,In_86,In_428);
nor U863 (N_863,In_337,In_365);
nor U864 (N_864,In_474,In_449);
nand U865 (N_865,In_88,In_10);
and U866 (N_866,In_459,In_178);
nor U867 (N_867,In_140,In_449);
nand U868 (N_868,In_90,In_3);
nand U869 (N_869,In_223,In_375);
and U870 (N_870,In_109,In_265);
and U871 (N_871,In_341,In_450);
nand U872 (N_872,In_239,In_246);
xor U873 (N_873,In_237,In_357);
xnor U874 (N_874,In_449,In_416);
or U875 (N_875,In_205,In_249);
or U876 (N_876,In_310,In_342);
nor U877 (N_877,In_436,In_342);
xnor U878 (N_878,In_383,In_457);
nor U879 (N_879,In_219,In_401);
nor U880 (N_880,In_156,In_54);
nand U881 (N_881,In_242,In_345);
nor U882 (N_882,In_249,In_374);
nor U883 (N_883,In_123,In_133);
or U884 (N_884,In_122,In_364);
nor U885 (N_885,In_483,In_14);
or U886 (N_886,In_358,In_431);
nand U887 (N_887,In_288,In_351);
nor U888 (N_888,In_300,In_11);
and U889 (N_889,In_267,In_135);
and U890 (N_890,In_27,In_213);
nor U891 (N_891,In_492,In_380);
and U892 (N_892,In_400,In_253);
and U893 (N_893,In_136,In_310);
or U894 (N_894,In_461,In_268);
nor U895 (N_895,In_470,In_7);
or U896 (N_896,In_214,In_245);
nor U897 (N_897,In_40,In_343);
nand U898 (N_898,In_137,In_304);
nand U899 (N_899,In_209,In_246);
or U900 (N_900,In_313,In_108);
nor U901 (N_901,In_11,In_247);
nand U902 (N_902,In_404,In_69);
and U903 (N_903,In_386,In_360);
and U904 (N_904,In_378,In_224);
nor U905 (N_905,In_167,In_210);
or U906 (N_906,In_375,In_131);
nor U907 (N_907,In_272,In_399);
nand U908 (N_908,In_467,In_21);
nor U909 (N_909,In_102,In_3);
or U910 (N_910,In_427,In_456);
and U911 (N_911,In_127,In_125);
nand U912 (N_912,In_203,In_370);
and U913 (N_913,In_33,In_465);
nand U914 (N_914,In_312,In_337);
nand U915 (N_915,In_384,In_62);
or U916 (N_916,In_161,In_492);
and U917 (N_917,In_117,In_212);
and U918 (N_918,In_470,In_286);
nand U919 (N_919,In_343,In_202);
nor U920 (N_920,In_242,In_344);
or U921 (N_921,In_1,In_483);
nand U922 (N_922,In_57,In_367);
or U923 (N_923,In_68,In_361);
and U924 (N_924,In_194,In_440);
and U925 (N_925,In_455,In_287);
and U926 (N_926,In_204,In_461);
nand U927 (N_927,In_93,In_20);
nand U928 (N_928,In_26,In_392);
nand U929 (N_929,In_313,In_116);
or U930 (N_930,In_40,In_179);
xnor U931 (N_931,In_319,In_425);
nor U932 (N_932,In_424,In_385);
nand U933 (N_933,In_171,In_444);
nand U934 (N_934,In_37,In_246);
and U935 (N_935,In_447,In_137);
nor U936 (N_936,In_125,In_286);
or U937 (N_937,In_134,In_173);
or U938 (N_938,In_272,In_105);
nor U939 (N_939,In_52,In_4);
or U940 (N_940,In_202,In_99);
and U941 (N_941,In_248,In_72);
nor U942 (N_942,In_135,In_489);
xnor U943 (N_943,In_358,In_297);
xnor U944 (N_944,In_12,In_211);
nor U945 (N_945,In_492,In_382);
and U946 (N_946,In_350,In_324);
nor U947 (N_947,In_34,In_342);
nor U948 (N_948,In_360,In_174);
and U949 (N_949,In_299,In_222);
xor U950 (N_950,In_20,In_261);
xnor U951 (N_951,In_172,In_151);
nor U952 (N_952,In_132,In_387);
and U953 (N_953,In_2,In_22);
or U954 (N_954,In_234,In_64);
nor U955 (N_955,In_216,In_97);
nand U956 (N_956,In_379,In_313);
or U957 (N_957,In_486,In_131);
nor U958 (N_958,In_241,In_324);
nor U959 (N_959,In_90,In_218);
and U960 (N_960,In_484,In_95);
and U961 (N_961,In_428,In_393);
nor U962 (N_962,In_85,In_293);
or U963 (N_963,In_66,In_464);
and U964 (N_964,In_431,In_69);
or U965 (N_965,In_372,In_209);
nor U966 (N_966,In_108,In_447);
and U967 (N_967,In_91,In_263);
nor U968 (N_968,In_36,In_17);
and U969 (N_969,In_436,In_229);
nor U970 (N_970,In_268,In_99);
or U971 (N_971,In_51,In_251);
and U972 (N_972,In_367,In_348);
xor U973 (N_973,In_450,In_427);
and U974 (N_974,In_217,In_49);
or U975 (N_975,In_247,In_170);
nor U976 (N_976,In_259,In_395);
nand U977 (N_977,In_474,In_321);
nor U978 (N_978,In_164,In_191);
xnor U979 (N_979,In_373,In_1);
nand U980 (N_980,In_135,In_317);
nand U981 (N_981,In_33,In_298);
nor U982 (N_982,In_167,In_253);
or U983 (N_983,In_88,In_448);
and U984 (N_984,In_40,In_156);
nand U985 (N_985,In_119,In_38);
and U986 (N_986,In_397,In_38);
nor U987 (N_987,In_480,In_422);
nand U988 (N_988,In_98,In_490);
or U989 (N_989,In_309,In_367);
nor U990 (N_990,In_261,In_239);
or U991 (N_991,In_379,In_111);
and U992 (N_992,In_413,In_127);
nand U993 (N_993,In_453,In_25);
nand U994 (N_994,In_78,In_205);
or U995 (N_995,In_279,In_94);
or U996 (N_996,In_212,In_325);
xnor U997 (N_997,In_21,In_377);
nor U998 (N_998,In_377,In_330);
and U999 (N_999,In_165,In_448);
nand U1000 (N_1000,N_741,N_233);
and U1001 (N_1001,N_414,N_579);
nand U1002 (N_1002,N_739,N_522);
xnor U1003 (N_1003,N_296,N_416);
nor U1004 (N_1004,N_891,N_870);
nor U1005 (N_1005,N_877,N_720);
nand U1006 (N_1006,N_230,N_694);
or U1007 (N_1007,N_583,N_271);
nand U1008 (N_1008,N_422,N_104);
nand U1009 (N_1009,N_18,N_688);
nor U1010 (N_1010,N_175,N_386);
nor U1011 (N_1011,N_991,N_406);
and U1012 (N_1012,N_237,N_508);
or U1013 (N_1013,N_184,N_982);
nand U1014 (N_1014,N_192,N_849);
nor U1015 (N_1015,N_675,N_353);
or U1016 (N_1016,N_277,N_150);
and U1017 (N_1017,N_248,N_68);
or U1018 (N_1018,N_232,N_904);
nor U1019 (N_1019,N_698,N_956);
or U1020 (N_1020,N_518,N_286);
and U1021 (N_1021,N_63,N_722);
nand U1022 (N_1022,N_993,N_341);
and U1023 (N_1023,N_844,N_28);
nor U1024 (N_1024,N_37,N_415);
or U1025 (N_1025,N_785,N_926);
or U1026 (N_1026,N_862,N_968);
or U1027 (N_1027,N_738,N_110);
and U1028 (N_1028,N_839,N_626);
or U1029 (N_1029,N_874,N_348);
or U1030 (N_1030,N_501,N_813);
nand U1031 (N_1031,N_859,N_268);
and U1032 (N_1032,N_140,N_704);
nand U1033 (N_1033,N_605,N_735);
nor U1034 (N_1034,N_354,N_371);
and U1035 (N_1035,N_683,N_533);
nand U1036 (N_1036,N_73,N_352);
nand U1037 (N_1037,N_99,N_447);
or U1038 (N_1038,N_6,N_56);
nor U1039 (N_1039,N_337,N_498);
or U1040 (N_1040,N_466,N_152);
xnor U1041 (N_1041,N_798,N_95);
nand U1042 (N_1042,N_200,N_419);
and U1043 (N_1043,N_223,N_322);
and U1044 (N_1044,N_360,N_196);
and U1045 (N_1045,N_850,N_912);
xnor U1046 (N_1046,N_823,N_506);
and U1047 (N_1047,N_436,N_94);
xnor U1048 (N_1048,N_914,N_726);
nand U1049 (N_1049,N_328,N_393);
nor U1050 (N_1050,N_437,N_604);
or U1051 (N_1051,N_892,N_784);
nor U1052 (N_1052,N_293,N_611);
and U1053 (N_1053,N_111,N_960);
nor U1054 (N_1054,N_176,N_668);
or U1055 (N_1055,N_343,N_682);
and U1056 (N_1056,N_32,N_998);
or U1057 (N_1057,N_616,N_287);
or U1058 (N_1058,N_433,N_78);
and U1059 (N_1059,N_34,N_539);
and U1060 (N_1060,N_356,N_247);
nor U1061 (N_1061,N_229,N_679);
nor U1062 (N_1062,N_880,N_902);
nand U1063 (N_1063,N_655,N_796);
or U1064 (N_1064,N_70,N_962);
and U1065 (N_1065,N_217,N_194);
nand U1066 (N_1066,N_922,N_561);
nor U1067 (N_1067,N_527,N_687);
xor U1068 (N_1068,N_878,N_555);
nor U1069 (N_1069,N_568,N_995);
or U1070 (N_1070,N_462,N_314);
or U1071 (N_1071,N_100,N_510);
and U1072 (N_1072,N_969,N_310);
nor U1073 (N_1073,N_239,N_146);
or U1074 (N_1074,N_2,N_967);
or U1075 (N_1075,N_731,N_358);
nor U1076 (N_1076,N_743,N_584);
nand U1077 (N_1077,N_214,N_820);
or U1078 (N_1078,N_893,N_985);
and U1079 (N_1079,N_629,N_715);
xnor U1080 (N_1080,N_622,N_390);
nor U1081 (N_1081,N_559,N_427);
nor U1082 (N_1082,N_806,N_123);
or U1083 (N_1083,N_75,N_252);
or U1084 (N_1084,N_674,N_1);
or U1085 (N_1085,N_85,N_791);
or U1086 (N_1086,N_428,N_977);
nor U1087 (N_1087,N_573,N_472);
and U1088 (N_1088,N_215,N_795);
nand U1089 (N_1089,N_621,N_281);
nor U1090 (N_1090,N_334,N_854);
xor U1091 (N_1091,N_261,N_940);
nor U1092 (N_1092,N_109,N_638);
and U1093 (N_1093,N_942,N_576);
and U1094 (N_1094,N_582,N_167);
or U1095 (N_1095,N_244,N_966);
nor U1096 (N_1096,N_402,N_202);
nor U1097 (N_1097,N_551,N_366);
nor U1098 (N_1098,N_524,N_478);
nor U1099 (N_1099,N_391,N_166);
nand U1100 (N_1100,N_340,N_157);
and U1101 (N_1101,N_41,N_950);
nand U1102 (N_1102,N_558,N_297);
nand U1103 (N_1103,N_550,N_786);
nand U1104 (N_1104,N_836,N_882);
or U1105 (N_1105,N_464,N_23);
or U1106 (N_1106,N_613,N_114);
or U1107 (N_1107,N_285,N_938);
and U1108 (N_1108,N_490,N_650);
and U1109 (N_1109,N_936,N_696);
xor U1110 (N_1110,N_44,N_553);
or U1111 (N_1111,N_178,N_772);
nand U1112 (N_1112,N_544,N_908);
nor U1113 (N_1113,N_807,N_295);
nor U1114 (N_1114,N_47,N_760);
and U1115 (N_1115,N_482,N_917);
or U1116 (N_1116,N_319,N_292);
or U1117 (N_1117,N_843,N_377);
and U1118 (N_1118,N_925,N_378);
or U1119 (N_1119,N_549,N_746);
nand U1120 (N_1120,N_141,N_987);
and U1121 (N_1121,N_153,N_879);
and U1122 (N_1122,N_845,N_900);
nor U1123 (N_1123,N_690,N_72);
and U1124 (N_1124,N_211,N_886);
and U1125 (N_1125,N_164,N_595);
or U1126 (N_1126,N_983,N_842);
or U1127 (N_1127,N_990,N_21);
nand U1128 (N_1128,N_923,N_523);
and U1129 (N_1129,N_106,N_329);
nor U1130 (N_1130,N_748,N_131);
or U1131 (N_1131,N_779,N_607);
or U1132 (N_1132,N_661,N_442);
or U1133 (N_1133,N_747,N_405);
and U1134 (N_1134,N_161,N_137);
xor U1135 (N_1135,N_564,N_221);
nand U1136 (N_1136,N_617,N_288);
or U1137 (N_1137,N_231,N_413);
nor U1138 (N_1138,N_569,N_663);
nand U1139 (N_1139,N_376,N_970);
nand U1140 (N_1140,N_440,N_275);
and U1141 (N_1141,N_774,N_491);
or U1142 (N_1142,N_973,N_809);
or U1143 (N_1143,N_636,N_17);
or U1144 (N_1144,N_226,N_480);
nand U1145 (N_1145,N_603,N_461);
or U1146 (N_1146,N_708,N_717);
nor U1147 (N_1147,N_189,N_812);
nand U1148 (N_1148,N_24,N_811);
or U1149 (N_1149,N_97,N_703);
nand U1150 (N_1150,N_554,N_545);
xor U1151 (N_1151,N_205,N_208);
and U1152 (N_1152,N_896,N_915);
or U1153 (N_1153,N_115,N_173);
and U1154 (N_1154,N_804,N_656);
and U1155 (N_1155,N_361,N_869);
and U1156 (N_1156,N_289,N_51);
or U1157 (N_1157,N_417,N_602);
nand U1158 (N_1158,N_61,N_160);
nand U1159 (N_1159,N_623,N_136);
nand U1160 (N_1160,N_372,N_635);
nand U1161 (N_1161,N_392,N_66);
and U1162 (N_1162,N_955,N_815);
and U1163 (N_1163,N_919,N_448);
xnor U1164 (N_1164,N_680,N_941);
nor U1165 (N_1165,N_62,N_35);
and U1166 (N_1166,N_643,N_625);
and U1167 (N_1167,N_557,N_238);
nand U1168 (N_1168,N_338,N_997);
nor U1169 (N_1169,N_734,N_280);
or U1170 (N_1170,N_409,N_716);
and U1171 (N_1171,N_504,N_875);
and U1172 (N_1172,N_156,N_646);
nand U1173 (N_1173,N_566,N_267);
nor U1174 (N_1174,N_630,N_283);
nand U1175 (N_1175,N_446,N_457);
nor U1176 (N_1176,N_677,N_924);
nand U1177 (N_1177,N_155,N_327);
nand U1178 (N_1178,N_592,N_505);
or U1179 (N_1179,N_108,N_119);
or U1180 (N_1180,N_455,N_712);
and U1181 (N_1181,N_702,N_978);
or U1182 (N_1182,N_79,N_395);
nand U1183 (N_1183,N_52,N_362);
nand U1184 (N_1184,N_305,N_188);
nor U1185 (N_1185,N_57,N_374);
and U1186 (N_1186,N_400,N_133);
and U1187 (N_1187,N_245,N_364);
and U1188 (N_1188,N_718,N_183);
nor U1189 (N_1189,N_947,N_441);
or U1190 (N_1190,N_777,N_837);
or U1191 (N_1191,N_606,N_769);
xnor U1192 (N_1192,N_793,N_468);
or U1193 (N_1193,N_383,N_531);
or U1194 (N_1194,N_686,N_313);
xor U1195 (N_1195,N_494,N_856);
nor U1196 (N_1196,N_979,N_794);
or U1197 (N_1197,N_540,N_996);
nand U1198 (N_1198,N_681,N_359);
nand U1199 (N_1199,N_596,N_719);
or U1200 (N_1200,N_113,N_81);
and U1201 (N_1201,N_42,N_972);
xor U1202 (N_1202,N_989,N_534);
nand U1203 (N_1203,N_253,N_312);
nor U1204 (N_1204,N_935,N_671);
or U1205 (N_1205,N_631,N_577);
or U1206 (N_1206,N_654,N_840);
nand U1207 (N_1207,N_380,N_43);
xnor U1208 (N_1208,N_496,N_833);
nand U1209 (N_1209,N_556,N_756);
nand U1210 (N_1210,N_740,N_162);
nor U1211 (N_1211,N_601,N_209);
and U1212 (N_1212,N_810,N_771);
nor U1213 (N_1213,N_235,N_357);
or U1214 (N_1214,N_615,N_13);
or U1215 (N_1215,N_701,N_775);
and U1216 (N_1216,N_116,N_570);
nand U1217 (N_1217,N_302,N_884);
and U1218 (N_1218,N_450,N_339);
nor U1219 (N_1219,N_259,N_787);
and U1220 (N_1220,N_742,N_600);
or U1221 (N_1221,N_346,N_29);
or U1222 (N_1222,N_254,N_883);
nor U1223 (N_1223,N_538,N_790);
and U1224 (N_1224,N_483,N_326);
nand U1225 (N_1225,N_332,N_665);
or U1226 (N_1226,N_282,N_828);
nand U1227 (N_1227,N_961,N_265);
or U1228 (N_1228,N_198,N_432);
nor U1229 (N_1229,N_379,N_789);
nor U1230 (N_1230,N_610,N_250);
or U1231 (N_1231,N_971,N_976);
and U1232 (N_1232,N_709,N_224);
or U1233 (N_1233,N_459,N_894);
xor U1234 (N_1234,N_20,N_516);
and U1235 (N_1235,N_49,N_486);
nand U1236 (N_1236,N_799,N_881);
nand U1237 (N_1237,N_632,N_475);
or U1238 (N_1238,N_86,N_946);
nand U1239 (N_1239,N_673,N_633);
or U1240 (N_1240,N_449,N_456);
nor U1241 (N_1241,N_721,N_39);
and U1242 (N_1242,N_788,N_365);
nor U1243 (N_1243,N_102,N_48);
and U1244 (N_1244,N_838,N_768);
nor U1245 (N_1245,N_382,N_445);
xnor U1246 (N_1246,N_389,N_325);
xor U1247 (N_1247,N_401,N_575);
and U1248 (N_1248,N_901,N_429);
or U1249 (N_1249,N_817,N_418);
nor U1250 (N_1250,N_725,N_255);
nand U1251 (N_1251,N_397,N_814);
or U1252 (N_1252,N_916,N_930);
xnor U1253 (N_1253,N_135,N_444);
nand U1254 (N_1254,N_857,N_780);
xnor U1255 (N_1255,N_163,N_762);
nor U1256 (N_1256,N_773,N_599);
nand U1257 (N_1257,N_170,N_492);
nand U1258 (N_1258,N_578,N_776);
nor U1259 (N_1259,N_168,N_808);
nand U1260 (N_1260,N_649,N_127);
or U1261 (N_1261,N_349,N_321);
nor U1262 (N_1262,N_71,N_994);
nand U1263 (N_1263,N_782,N_749);
or U1264 (N_1264,N_619,N_125);
nor U1265 (N_1265,N_481,N_565);
or U1266 (N_1266,N_846,N_803);
nand U1267 (N_1267,N_639,N_537);
and U1268 (N_1268,N_19,N_98);
nand U1269 (N_1269,N_80,N_819);
and U1270 (N_1270,N_130,N_699);
nor U1271 (N_1271,N_648,N_805);
or U1272 (N_1272,N_195,N_503);
nor U1273 (N_1273,N_301,N_608);
nor U1274 (N_1274,N_46,N_934);
nand U1275 (N_1275,N_107,N_944);
nor U1276 (N_1276,N_50,N_246);
nand U1277 (N_1277,N_647,N_954);
or U1278 (N_1278,N_937,N_399);
and U1279 (N_1279,N_580,N_560);
and U1280 (N_1280,N_197,N_887);
or U1281 (N_1281,N_3,N_324);
or U1282 (N_1282,N_974,N_404);
nand U1283 (N_1283,N_477,N_236);
nand U1284 (N_1284,N_451,N_586);
and U1285 (N_1285,N_112,N_588);
nand U1286 (N_1286,N_890,N_899);
or U1287 (N_1287,N_847,N_407);
nand U1288 (N_1288,N_350,N_543);
nor U1289 (N_1289,N_851,N_30);
and U1290 (N_1290,N_951,N_871);
nor U1291 (N_1291,N_792,N_678);
nor U1292 (N_1292,N_585,N_865);
nor U1293 (N_1293,N_889,N_278);
or U1294 (N_1294,N_965,N_500);
nor U1295 (N_1295,N_920,N_210);
or U1296 (N_1296,N_258,N_905);
xnor U1297 (N_1297,N_40,N_520);
or U1298 (N_1298,N_454,N_727);
nand U1299 (N_1299,N_315,N_467);
or U1300 (N_1300,N_535,N_958);
or U1301 (N_1301,N_122,N_530);
nor U1302 (N_1302,N_853,N_58);
nor U1303 (N_1303,N_485,N_662);
and U1304 (N_1304,N_129,N_660);
xnor U1305 (N_1305,N_11,N_824);
or U1306 (N_1306,N_33,N_64);
and U1307 (N_1307,N_513,N_228);
nor U1308 (N_1308,N_60,N_158);
or U1309 (N_1309,N_858,N_832);
and U1310 (N_1310,N_642,N_385);
or U1311 (N_1311,N_124,N_898);
and U1312 (N_1312,N_84,N_143);
xnor U1313 (N_1313,N_949,N_572);
nor U1314 (N_1314,N_980,N_154);
nor U1315 (N_1315,N_177,N_581);
xor U1316 (N_1316,N_931,N_866);
xor U1317 (N_1317,N_672,N_299);
nor U1318 (N_1318,N_284,N_384);
or U1319 (N_1319,N_207,N_932);
nor U1320 (N_1320,N_975,N_733);
and U1321 (N_1321,N_800,N_667);
and U1322 (N_1322,N_430,N_330);
nor U1323 (N_1323,N_827,N_710);
or U1324 (N_1324,N_487,N_88);
and U1325 (N_1325,N_640,N_181);
nand U1326 (N_1326,N_342,N_225);
nand U1327 (N_1327,N_101,N_8);
or U1328 (N_1328,N_249,N_628);
or U1329 (N_1329,N_999,N_744);
and U1330 (N_1330,N_262,N_511);
nor U1331 (N_1331,N_190,N_781);
and U1332 (N_1332,N_410,N_700);
or U1333 (N_1333,N_499,N_90);
or U1334 (N_1334,N_151,N_120);
and U1335 (N_1335,N_597,N_528);
nor U1336 (N_1336,N_142,N_927);
and U1337 (N_1337,N_861,N_304);
nor U1338 (N_1338,N_532,N_618);
xnor U1339 (N_1339,N_770,N_270);
nor U1340 (N_1340,N_766,N_659);
nand U1341 (N_1341,N_420,N_182);
and U1342 (N_1342,N_54,N_105);
and U1343 (N_1343,N_755,N_344);
and U1344 (N_1344,N_5,N_479);
or U1345 (N_1345,N_272,N_964);
nand U1346 (N_1346,N_77,N_897);
xnor U1347 (N_1347,N_431,N_256);
or U1348 (N_1348,N_10,N_658);
or U1349 (N_1349,N_303,N_826);
and U1350 (N_1350,N_460,N_957);
and U1351 (N_1351,N_12,N_169);
nand U1352 (N_1352,N_598,N_928);
nor U1353 (N_1353,N_74,N_992);
nand U1354 (N_1354,N_53,N_868);
and U1355 (N_1355,N_750,N_952);
nand U1356 (N_1356,N_728,N_7);
nor U1357 (N_1357,N_92,N_291);
or U1358 (N_1358,N_644,N_763);
xor U1359 (N_1359,N_594,N_981);
and U1360 (N_1360,N_909,N_745);
or U1361 (N_1361,N_587,N_172);
xor U1362 (N_1362,N_624,N_567);
nand U1363 (N_1363,N_724,N_300);
nor U1364 (N_1364,N_707,N_421);
nor U1365 (N_1365,N_45,N_984);
nor U1366 (N_1366,N_918,N_333);
or U1367 (N_1367,N_201,N_375);
xor U1368 (N_1368,N_276,N_103);
or U1369 (N_1369,N_841,N_864);
nor U1370 (N_1370,N_590,N_212);
and U1371 (N_1371,N_489,N_641);
nand U1372 (N_1372,N_128,N_802);
nand U1373 (N_1373,N_986,N_387);
and U1374 (N_1374,N_546,N_4);
nor U1375 (N_1375,N_318,N_91);
or U1376 (N_1376,N_59,N_373);
nand U1377 (N_1377,N_38,N_159);
or U1378 (N_1378,N_320,N_191);
or U1379 (N_1379,N_695,N_185);
nor U1380 (N_1380,N_251,N_264);
and U1381 (N_1381,N_509,N_206);
nand U1382 (N_1382,N_398,N_885);
or U1383 (N_1383,N_911,N_737);
and U1384 (N_1384,N_563,N_241);
and U1385 (N_1385,N_863,N_149);
and U1386 (N_1386,N_729,N_693);
and U1387 (N_1387,N_403,N_873);
nor U1388 (N_1388,N_317,N_903);
nand U1389 (N_1389,N_87,N_396);
nor U1390 (N_1390,N_139,N_132);
nand U1391 (N_1391,N_469,N_126);
xor U1392 (N_1392,N_323,N_541);
nor U1393 (N_1393,N_764,N_369);
nand U1394 (N_1394,N_848,N_759);
nand U1395 (N_1395,N_316,N_171);
nor U1396 (N_1396,N_118,N_408);
nand U1397 (N_1397,N_888,N_65);
and U1398 (N_1398,N_684,N_637);
and U1399 (N_1399,N_614,N_666);
and U1400 (N_1400,N_263,N_9);
and U1401 (N_1401,N_816,N_484);
or U1402 (N_1402,N_829,N_706);
nor U1403 (N_1403,N_55,N_273);
nor U1404 (N_1404,N_452,N_345);
or U1405 (N_1405,N_363,N_425);
or U1406 (N_1406,N_82,N_347);
xnor U1407 (N_1407,N_434,N_204);
nor U1408 (N_1408,N_591,N_193);
or U1409 (N_1409,N_243,N_855);
xnor U1410 (N_1410,N_758,N_645);
or U1411 (N_1411,N_174,N_945);
nor U1412 (N_1412,N_298,N_308);
nor U1413 (N_1413,N_279,N_652);
xor U1414 (N_1414,N_227,N_948);
or U1415 (N_1415,N_213,N_526);
or U1416 (N_1416,N_370,N_818);
nand U1417 (N_1417,N_657,N_801);
nand U1418 (N_1418,N_83,N_187);
or U1419 (N_1419,N_872,N_988);
or U1420 (N_1420,N_473,N_921);
and U1421 (N_1421,N_493,N_465);
or U1422 (N_1422,N_294,N_732);
xnor U1423 (N_1423,N_529,N_512);
or U1424 (N_1424,N_495,N_730);
nor U1425 (N_1425,N_822,N_571);
and U1426 (N_1426,N_394,N_257);
nor U1427 (N_1427,N_552,N_653);
and U1428 (N_1428,N_825,N_89);
and U1429 (N_1429,N_222,N_929);
nand U1430 (N_1430,N_266,N_754);
or U1431 (N_1431,N_547,N_562);
or U1432 (N_1432,N_471,N_691);
or U1433 (N_1433,N_907,N_525);
nor U1434 (N_1434,N_589,N_67);
nor U1435 (N_1435,N_574,N_831);
or U1436 (N_1436,N_242,N_424);
nor U1437 (N_1437,N_497,N_548);
and U1438 (N_1438,N_963,N_439);
or U1439 (N_1439,N_351,N_309);
or U1440 (N_1440,N_15,N_515);
and U1441 (N_1441,N_307,N_959);
and U1442 (N_1442,N_723,N_0);
or U1443 (N_1443,N_507,N_458);
and U1444 (N_1444,N_306,N_220);
nor U1445 (N_1445,N_269,N_203);
and U1446 (N_1446,N_895,N_144);
nand U1447 (N_1447,N_783,N_117);
nand U1448 (N_1448,N_234,N_31);
or U1449 (N_1449,N_767,N_670);
nand U1450 (N_1450,N_179,N_834);
nand U1451 (N_1451,N_26,N_620);
or U1452 (N_1452,N_216,N_438);
nor U1453 (N_1453,N_180,N_765);
and U1454 (N_1454,N_165,N_536);
or U1455 (N_1455,N_676,N_476);
and U1456 (N_1456,N_692,N_134);
and U1457 (N_1457,N_913,N_381);
nor U1458 (N_1458,N_219,N_821);
nor U1459 (N_1459,N_16,N_514);
or U1460 (N_1460,N_797,N_711);
and U1461 (N_1461,N_25,N_290);
and U1462 (N_1462,N_757,N_697);
and U1463 (N_1463,N_612,N_148);
or U1464 (N_1464,N_274,N_943);
and U1465 (N_1465,N_752,N_502);
nor U1466 (N_1466,N_412,N_336);
or U1467 (N_1467,N_463,N_388);
and U1468 (N_1468,N_761,N_335);
and U1469 (N_1469,N_651,N_423);
or U1470 (N_1470,N_186,N_27);
xor U1471 (N_1471,N_778,N_331);
or U1472 (N_1472,N_260,N_867);
or U1473 (N_1473,N_443,N_627);
and U1474 (N_1474,N_121,N_69);
and U1475 (N_1475,N_76,N_939);
nand U1476 (N_1476,N_96,N_311);
nand U1477 (N_1477,N_876,N_689);
nand U1478 (N_1478,N_435,N_517);
and U1479 (N_1479,N_753,N_145);
xor U1480 (N_1480,N_488,N_669);
and U1481 (N_1481,N_470,N_542);
and U1482 (N_1482,N_453,N_240);
nand U1483 (N_1483,N_355,N_411);
nand U1484 (N_1484,N_852,N_664);
and U1485 (N_1485,N_474,N_426);
nor U1486 (N_1486,N_751,N_714);
and U1487 (N_1487,N_685,N_713);
or U1488 (N_1488,N_634,N_138);
nand U1489 (N_1489,N_860,N_199);
nand U1490 (N_1490,N_36,N_367);
or U1491 (N_1491,N_218,N_519);
nor U1492 (N_1492,N_93,N_521);
nand U1493 (N_1493,N_835,N_14);
or U1494 (N_1494,N_593,N_736);
nand U1495 (N_1495,N_368,N_906);
xnor U1496 (N_1496,N_705,N_910);
nand U1497 (N_1497,N_147,N_830);
or U1498 (N_1498,N_22,N_953);
and U1499 (N_1499,N_609,N_933);
nor U1500 (N_1500,N_298,N_519);
xor U1501 (N_1501,N_599,N_481);
or U1502 (N_1502,N_353,N_158);
nand U1503 (N_1503,N_245,N_446);
xor U1504 (N_1504,N_688,N_141);
or U1505 (N_1505,N_915,N_184);
or U1506 (N_1506,N_906,N_690);
nand U1507 (N_1507,N_71,N_431);
and U1508 (N_1508,N_295,N_800);
and U1509 (N_1509,N_33,N_882);
nor U1510 (N_1510,N_469,N_127);
nor U1511 (N_1511,N_144,N_377);
and U1512 (N_1512,N_692,N_418);
nor U1513 (N_1513,N_673,N_663);
nor U1514 (N_1514,N_393,N_466);
and U1515 (N_1515,N_248,N_54);
nor U1516 (N_1516,N_868,N_572);
and U1517 (N_1517,N_417,N_142);
nand U1518 (N_1518,N_286,N_669);
nor U1519 (N_1519,N_666,N_416);
and U1520 (N_1520,N_617,N_764);
nor U1521 (N_1521,N_360,N_920);
and U1522 (N_1522,N_409,N_185);
or U1523 (N_1523,N_880,N_442);
nor U1524 (N_1524,N_436,N_337);
nor U1525 (N_1525,N_661,N_317);
xor U1526 (N_1526,N_188,N_746);
nor U1527 (N_1527,N_949,N_803);
or U1528 (N_1528,N_334,N_749);
nand U1529 (N_1529,N_125,N_1);
or U1530 (N_1530,N_57,N_405);
nor U1531 (N_1531,N_816,N_725);
nor U1532 (N_1532,N_630,N_228);
or U1533 (N_1533,N_959,N_948);
nor U1534 (N_1534,N_400,N_680);
xnor U1535 (N_1535,N_872,N_423);
nand U1536 (N_1536,N_348,N_934);
and U1537 (N_1537,N_119,N_380);
or U1538 (N_1538,N_765,N_281);
nor U1539 (N_1539,N_979,N_521);
nand U1540 (N_1540,N_631,N_730);
or U1541 (N_1541,N_768,N_61);
or U1542 (N_1542,N_132,N_824);
nand U1543 (N_1543,N_352,N_489);
xor U1544 (N_1544,N_397,N_29);
nor U1545 (N_1545,N_535,N_491);
nor U1546 (N_1546,N_246,N_108);
nand U1547 (N_1547,N_815,N_931);
and U1548 (N_1548,N_796,N_492);
or U1549 (N_1549,N_344,N_539);
or U1550 (N_1550,N_21,N_436);
and U1551 (N_1551,N_962,N_772);
or U1552 (N_1552,N_668,N_108);
or U1553 (N_1553,N_289,N_163);
nand U1554 (N_1554,N_51,N_928);
or U1555 (N_1555,N_542,N_284);
xor U1556 (N_1556,N_739,N_932);
xor U1557 (N_1557,N_222,N_547);
nor U1558 (N_1558,N_672,N_683);
xnor U1559 (N_1559,N_273,N_667);
nand U1560 (N_1560,N_506,N_197);
nor U1561 (N_1561,N_753,N_211);
nor U1562 (N_1562,N_749,N_847);
and U1563 (N_1563,N_477,N_79);
and U1564 (N_1564,N_480,N_312);
and U1565 (N_1565,N_991,N_324);
nor U1566 (N_1566,N_117,N_306);
and U1567 (N_1567,N_924,N_881);
and U1568 (N_1568,N_122,N_314);
nand U1569 (N_1569,N_93,N_152);
or U1570 (N_1570,N_983,N_744);
and U1571 (N_1571,N_856,N_267);
or U1572 (N_1572,N_467,N_429);
xnor U1573 (N_1573,N_105,N_768);
nor U1574 (N_1574,N_651,N_606);
xnor U1575 (N_1575,N_693,N_110);
nand U1576 (N_1576,N_902,N_91);
nor U1577 (N_1577,N_912,N_980);
nor U1578 (N_1578,N_822,N_703);
or U1579 (N_1579,N_903,N_137);
nand U1580 (N_1580,N_206,N_825);
or U1581 (N_1581,N_447,N_441);
and U1582 (N_1582,N_940,N_508);
nand U1583 (N_1583,N_315,N_947);
and U1584 (N_1584,N_921,N_942);
and U1585 (N_1585,N_598,N_651);
xnor U1586 (N_1586,N_961,N_698);
or U1587 (N_1587,N_353,N_172);
nand U1588 (N_1588,N_520,N_712);
or U1589 (N_1589,N_738,N_859);
xnor U1590 (N_1590,N_324,N_640);
and U1591 (N_1591,N_763,N_27);
or U1592 (N_1592,N_513,N_38);
xnor U1593 (N_1593,N_926,N_394);
nand U1594 (N_1594,N_19,N_695);
or U1595 (N_1595,N_125,N_645);
and U1596 (N_1596,N_54,N_477);
and U1597 (N_1597,N_575,N_848);
nor U1598 (N_1598,N_780,N_309);
and U1599 (N_1599,N_855,N_615);
nor U1600 (N_1600,N_26,N_420);
xor U1601 (N_1601,N_880,N_337);
nor U1602 (N_1602,N_310,N_919);
or U1603 (N_1603,N_23,N_835);
xor U1604 (N_1604,N_513,N_823);
nor U1605 (N_1605,N_973,N_560);
or U1606 (N_1606,N_284,N_711);
nor U1607 (N_1607,N_725,N_823);
nand U1608 (N_1608,N_18,N_206);
nor U1609 (N_1609,N_142,N_561);
nor U1610 (N_1610,N_184,N_832);
nor U1611 (N_1611,N_429,N_649);
or U1612 (N_1612,N_354,N_403);
nor U1613 (N_1613,N_783,N_360);
and U1614 (N_1614,N_92,N_3);
and U1615 (N_1615,N_304,N_481);
and U1616 (N_1616,N_193,N_885);
nand U1617 (N_1617,N_640,N_813);
or U1618 (N_1618,N_909,N_693);
or U1619 (N_1619,N_495,N_881);
and U1620 (N_1620,N_220,N_204);
and U1621 (N_1621,N_671,N_797);
or U1622 (N_1622,N_381,N_751);
xor U1623 (N_1623,N_585,N_669);
or U1624 (N_1624,N_778,N_898);
nor U1625 (N_1625,N_299,N_261);
nand U1626 (N_1626,N_199,N_992);
and U1627 (N_1627,N_201,N_900);
nor U1628 (N_1628,N_396,N_290);
xnor U1629 (N_1629,N_288,N_880);
and U1630 (N_1630,N_332,N_807);
nor U1631 (N_1631,N_368,N_106);
nor U1632 (N_1632,N_739,N_148);
and U1633 (N_1633,N_171,N_599);
or U1634 (N_1634,N_852,N_803);
or U1635 (N_1635,N_260,N_651);
nor U1636 (N_1636,N_291,N_979);
xor U1637 (N_1637,N_488,N_327);
nand U1638 (N_1638,N_243,N_854);
or U1639 (N_1639,N_262,N_210);
nand U1640 (N_1640,N_56,N_227);
and U1641 (N_1641,N_850,N_869);
nand U1642 (N_1642,N_78,N_793);
nor U1643 (N_1643,N_404,N_103);
and U1644 (N_1644,N_225,N_129);
nor U1645 (N_1645,N_702,N_98);
or U1646 (N_1646,N_233,N_904);
xnor U1647 (N_1647,N_940,N_465);
or U1648 (N_1648,N_17,N_719);
nor U1649 (N_1649,N_516,N_29);
nor U1650 (N_1650,N_68,N_422);
xnor U1651 (N_1651,N_491,N_740);
or U1652 (N_1652,N_617,N_34);
and U1653 (N_1653,N_105,N_322);
nand U1654 (N_1654,N_697,N_270);
nor U1655 (N_1655,N_892,N_807);
nor U1656 (N_1656,N_79,N_381);
xor U1657 (N_1657,N_934,N_652);
or U1658 (N_1658,N_663,N_151);
nand U1659 (N_1659,N_426,N_151);
or U1660 (N_1660,N_726,N_512);
xor U1661 (N_1661,N_809,N_235);
nor U1662 (N_1662,N_229,N_291);
and U1663 (N_1663,N_352,N_853);
xor U1664 (N_1664,N_176,N_14);
nand U1665 (N_1665,N_919,N_438);
nor U1666 (N_1666,N_144,N_806);
nand U1667 (N_1667,N_18,N_166);
xnor U1668 (N_1668,N_218,N_509);
nand U1669 (N_1669,N_387,N_816);
nand U1670 (N_1670,N_330,N_837);
xor U1671 (N_1671,N_658,N_374);
and U1672 (N_1672,N_97,N_66);
nand U1673 (N_1673,N_525,N_894);
nor U1674 (N_1674,N_801,N_316);
xnor U1675 (N_1675,N_301,N_997);
or U1676 (N_1676,N_196,N_430);
and U1677 (N_1677,N_229,N_670);
or U1678 (N_1678,N_391,N_853);
or U1679 (N_1679,N_406,N_927);
nand U1680 (N_1680,N_795,N_972);
nor U1681 (N_1681,N_925,N_926);
and U1682 (N_1682,N_215,N_494);
nand U1683 (N_1683,N_777,N_534);
nor U1684 (N_1684,N_700,N_891);
nand U1685 (N_1685,N_944,N_674);
or U1686 (N_1686,N_716,N_694);
xnor U1687 (N_1687,N_161,N_108);
or U1688 (N_1688,N_557,N_707);
and U1689 (N_1689,N_5,N_532);
and U1690 (N_1690,N_218,N_406);
and U1691 (N_1691,N_164,N_992);
or U1692 (N_1692,N_808,N_157);
nor U1693 (N_1693,N_819,N_738);
nand U1694 (N_1694,N_795,N_519);
or U1695 (N_1695,N_765,N_599);
xor U1696 (N_1696,N_154,N_955);
nand U1697 (N_1697,N_718,N_829);
and U1698 (N_1698,N_176,N_609);
nor U1699 (N_1699,N_885,N_911);
nand U1700 (N_1700,N_977,N_441);
or U1701 (N_1701,N_177,N_574);
nand U1702 (N_1702,N_674,N_244);
or U1703 (N_1703,N_955,N_693);
or U1704 (N_1704,N_441,N_705);
and U1705 (N_1705,N_128,N_546);
or U1706 (N_1706,N_945,N_553);
and U1707 (N_1707,N_422,N_51);
or U1708 (N_1708,N_611,N_206);
nor U1709 (N_1709,N_385,N_58);
or U1710 (N_1710,N_544,N_653);
nor U1711 (N_1711,N_293,N_643);
nor U1712 (N_1712,N_790,N_119);
xnor U1713 (N_1713,N_155,N_152);
or U1714 (N_1714,N_968,N_748);
xnor U1715 (N_1715,N_219,N_561);
or U1716 (N_1716,N_103,N_856);
nand U1717 (N_1717,N_469,N_815);
xnor U1718 (N_1718,N_635,N_660);
nand U1719 (N_1719,N_491,N_502);
or U1720 (N_1720,N_141,N_543);
nor U1721 (N_1721,N_557,N_944);
or U1722 (N_1722,N_179,N_785);
or U1723 (N_1723,N_64,N_771);
or U1724 (N_1724,N_575,N_570);
and U1725 (N_1725,N_665,N_262);
nand U1726 (N_1726,N_876,N_773);
and U1727 (N_1727,N_494,N_576);
nand U1728 (N_1728,N_323,N_264);
xnor U1729 (N_1729,N_720,N_523);
or U1730 (N_1730,N_113,N_396);
nand U1731 (N_1731,N_79,N_434);
nor U1732 (N_1732,N_476,N_230);
nand U1733 (N_1733,N_982,N_876);
nand U1734 (N_1734,N_314,N_373);
nand U1735 (N_1735,N_898,N_685);
nand U1736 (N_1736,N_871,N_640);
nor U1737 (N_1737,N_374,N_107);
nor U1738 (N_1738,N_438,N_483);
and U1739 (N_1739,N_65,N_245);
nor U1740 (N_1740,N_747,N_543);
nand U1741 (N_1741,N_598,N_953);
nand U1742 (N_1742,N_361,N_547);
nor U1743 (N_1743,N_50,N_2);
or U1744 (N_1744,N_36,N_609);
xnor U1745 (N_1745,N_642,N_21);
nor U1746 (N_1746,N_67,N_73);
or U1747 (N_1747,N_350,N_401);
nand U1748 (N_1748,N_873,N_454);
xor U1749 (N_1749,N_0,N_699);
nor U1750 (N_1750,N_639,N_104);
and U1751 (N_1751,N_638,N_839);
xor U1752 (N_1752,N_867,N_112);
and U1753 (N_1753,N_562,N_963);
xor U1754 (N_1754,N_749,N_643);
and U1755 (N_1755,N_208,N_595);
and U1756 (N_1756,N_524,N_316);
or U1757 (N_1757,N_175,N_481);
or U1758 (N_1758,N_740,N_314);
nor U1759 (N_1759,N_875,N_319);
xor U1760 (N_1760,N_58,N_301);
or U1761 (N_1761,N_839,N_484);
nor U1762 (N_1762,N_542,N_53);
nor U1763 (N_1763,N_952,N_242);
nand U1764 (N_1764,N_146,N_649);
or U1765 (N_1765,N_336,N_195);
and U1766 (N_1766,N_749,N_139);
or U1767 (N_1767,N_482,N_819);
xor U1768 (N_1768,N_165,N_967);
nand U1769 (N_1769,N_298,N_495);
nand U1770 (N_1770,N_162,N_910);
nand U1771 (N_1771,N_697,N_999);
or U1772 (N_1772,N_25,N_334);
nor U1773 (N_1773,N_85,N_411);
nor U1774 (N_1774,N_628,N_374);
or U1775 (N_1775,N_567,N_922);
xor U1776 (N_1776,N_955,N_864);
or U1777 (N_1777,N_114,N_147);
nand U1778 (N_1778,N_39,N_250);
and U1779 (N_1779,N_497,N_522);
and U1780 (N_1780,N_333,N_450);
nand U1781 (N_1781,N_965,N_478);
xor U1782 (N_1782,N_621,N_411);
and U1783 (N_1783,N_544,N_490);
and U1784 (N_1784,N_830,N_715);
or U1785 (N_1785,N_47,N_272);
nand U1786 (N_1786,N_27,N_787);
xor U1787 (N_1787,N_281,N_426);
nor U1788 (N_1788,N_101,N_347);
or U1789 (N_1789,N_561,N_686);
or U1790 (N_1790,N_429,N_143);
nand U1791 (N_1791,N_607,N_910);
nand U1792 (N_1792,N_725,N_772);
or U1793 (N_1793,N_741,N_218);
or U1794 (N_1794,N_250,N_905);
xor U1795 (N_1795,N_515,N_596);
and U1796 (N_1796,N_155,N_979);
or U1797 (N_1797,N_964,N_125);
and U1798 (N_1798,N_481,N_594);
and U1799 (N_1799,N_746,N_466);
xor U1800 (N_1800,N_653,N_197);
nor U1801 (N_1801,N_403,N_470);
or U1802 (N_1802,N_883,N_618);
or U1803 (N_1803,N_111,N_103);
and U1804 (N_1804,N_360,N_850);
or U1805 (N_1805,N_285,N_922);
nor U1806 (N_1806,N_23,N_657);
nor U1807 (N_1807,N_423,N_102);
or U1808 (N_1808,N_621,N_716);
or U1809 (N_1809,N_806,N_59);
nor U1810 (N_1810,N_412,N_275);
nor U1811 (N_1811,N_438,N_732);
or U1812 (N_1812,N_842,N_425);
nor U1813 (N_1813,N_962,N_582);
and U1814 (N_1814,N_620,N_739);
xor U1815 (N_1815,N_808,N_565);
or U1816 (N_1816,N_488,N_376);
xnor U1817 (N_1817,N_81,N_231);
or U1818 (N_1818,N_46,N_729);
or U1819 (N_1819,N_169,N_65);
nor U1820 (N_1820,N_434,N_572);
or U1821 (N_1821,N_780,N_865);
nor U1822 (N_1822,N_878,N_854);
xor U1823 (N_1823,N_573,N_833);
or U1824 (N_1824,N_799,N_625);
and U1825 (N_1825,N_394,N_169);
or U1826 (N_1826,N_729,N_224);
nor U1827 (N_1827,N_27,N_779);
or U1828 (N_1828,N_73,N_84);
and U1829 (N_1829,N_528,N_599);
nor U1830 (N_1830,N_180,N_387);
nor U1831 (N_1831,N_281,N_437);
nor U1832 (N_1832,N_10,N_103);
nand U1833 (N_1833,N_815,N_2);
or U1834 (N_1834,N_429,N_603);
or U1835 (N_1835,N_764,N_552);
or U1836 (N_1836,N_132,N_811);
and U1837 (N_1837,N_298,N_90);
xnor U1838 (N_1838,N_685,N_687);
xnor U1839 (N_1839,N_146,N_99);
nand U1840 (N_1840,N_349,N_851);
or U1841 (N_1841,N_132,N_551);
nor U1842 (N_1842,N_236,N_779);
and U1843 (N_1843,N_375,N_139);
and U1844 (N_1844,N_35,N_671);
and U1845 (N_1845,N_533,N_442);
xor U1846 (N_1846,N_438,N_401);
or U1847 (N_1847,N_284,N_203);
or U1848 (N_1848,N_957,N_341);
nor U1849 (N_1849,N_949,N_765);
and U1850 (N_1850,N_558,N_576);
nand U1851 (N_1851,N_968,N_16);
or U1852 (N_1852,N_327,N_580);
or U1853 (N_1853,N_171,N_467);
and U1854 (N_1854,N_24,N_732);
nand U1855 (N_1855,N_194,N_704);
nor U1856 (N_1856,N_360,N_754);
nor U1857 (N_1857,N_893,N_100);
nand U1858 (N_1858,N_683,N_592);
or U1859 (N_1859,N_396,N_859);
or U1860 (N_1860,N_982,N_954);
or U1861 (N_1861,N_933,N_316);
nor U1862 (N_1862,N_397,N_649);
nand U1863 (N_1863,N_421,N_621);
nand U1864 (N_1864,N_270,N_510);
or U1865 (N_1865,N_909,N_711);
and U1866 (N_1866,N_647,N_868);
or U1867 (N_1867,N_851,N_130);
or U1868 (N_1868,N_831,N_298);
or U1869 (N_1869,N_275,N_240);
nor U1870 (N_1870,N_254,N_44);
nor U1871 (N_1871,N_231,N_27);
xnor U1872 (N_1872,N_424,N_880);
nand U1873 (N_1873,N_205,N_601);
nand U1874 (N_1874,N_237,N_649);
nand U1875 (N_1875,N_973,N_137);
nor U1876 (N_1876,N_985,N_877);
or U1877 (N_1877,N_805,N_359);
nor U1878 (N_1878,N_138,N_309);
nor U1879 (N_1879,N_528,N_374);
xnor U1880 (N_1880,N_578,N_534);
or U1881 (N_1881,N_184,N_256);
or U1882 (N_1882,N_748,N_980);
or U1883 (N_1883,N_204,N_143);
or U1884 (N_1884,N_204,N_960);
nor U1885 (N_1885,N_73,N_891);
xnor U1886 (N_1886,N_620,N_101);
nor U1887 (N_1887,N_842,N_202);
nor U1888 (N_1888,N_424,N_243);
and U1889 (N_1889,N_322,N_364);
xor U1890 (N_1890,N_872,N_932);
nand U1891 (N_1891,N_534,N_224);
xnor U1892 (N_1892,N_134,N_415);
nand U1893 (N_1893,N_213,N_749);
or U1894 (N_1894,N_541,N_150);
nor U1895 (N_1895,N_40,N_548);
nand U1896 (N_1896,N_322,N_55);
and U1897 (N_1897,N_108,N_462);
and U1898 (N_1898,N_432,N_763);
and U1899 (N_1899,N_141,N_965);
nor U1900 (N_1900,N_482,N_905);
or U1901 (N_1901,N_146,N_335);
or U1902 (N_1902,N_37,N_825);
and U1903 (N_1903,N_310,N_800);
nor U1904 (N_1904,N_496,N_340);
or U1905 (N_1905,N_573,N_167);
nor U1906 (N_1906,N_435,N_494);
and U1907 (N_1907,N_428,N_543);
and U1908 (N_1908,N_61,N_358);
nand U1909 (N_1909,N_693,N_344);
nor U1910 (N_1910,N_526,N_793);
and U1911 (N_1911,N_681,N_112);
or U1912 (N_1912,N_87,N_627);
or U1913 (N_1913,N_556,N_651);
and U1914 (N_1914,N_960,N_864);
xor U1915 (N_1915,N_539,N_280);
and U1916 (N_1916,N_133,N_698);
xor U1917 (N_1917,N_863,N_926);
and U1918 (N_1918,N_176,N_425);
or U1919 (N_1919,N_151,N_960);
nor U1920 (N_1920,N_666,N_928);
or U1921 (N_1921,N_747,N_875);
nor U1922 (N_1922,N_137,N_188);
nor U1923 (N_1923,N_739,N_201);
and U1924 (N_1924,N_788,N_370);
and U1925 (N_1925,N_241,N_191);
nor U1926 (N_1926,N_165,N_48);
nand U1927 (N_1927,N_880,N_192);
nor U1928 (N_1928,N_874,N_343);
nor U1929 (N_1929,N_101,N_865);
or U1930 (N_1930,N_540,N_576);
and U1931 (N_1931,N_830,N_361);
nor U1932 (N_1932,N_488,N_7);
nand U1933 (N_1933,N_627,N_599);
nand U1934 (N_1934,N_365,N_768);
nor U1935 (N_1935,N_614,N_830);
nand U1936 (N_1936,N_999,N_873);
nand U1937 (N_1937,N_910,N_37);
or U1938 (N_1938,N_814,N_559);
nand U1939 (N_1939,N_774,N_364);
xor U1940 (N_1940,N_780,N_550);
or U1941 (N_1941,N_317,N_106);
and U1942 (N_1942,N_476,N_402);
or U1943 (N_1943,N_705,N_455);
nand U1944 (N_1944,N_64,N_287);
or U1945 (N_1945,N_470,N_810);
and U1946 (N_1946,N_50,N_788);
nor U1947 (N_1947,N_940,N_990);
nor U1948 (N_1948,N_700,N_746);
nor U1949 (N_1949,N_267,N_386);
nand U1950 (N_1950,N_873,N_35);
nor U1951 (N_1951,N_191,N_822);
and U1952 (N_1952,N_363,N_573);
or U1953 (N_1953,N_716,N_932);
nand U1954 (N_1954,N_153,N_482);
xor U1955 (N_1955,N_241,N_333);
nor U1956 (N_1956,N_658,N_42);
nor U1957 (N_1957,N_800,N_228);
and U1958 (N_1958,N_381,N_783);
xor U1959 (N_1959,N_20,N_262);
nand U1960 (N_1960,N_309,N_55);
and U1961 (N_1961,N_254,N_111);
or U1962 (N_1962,N_962,N_970);
nor U1963 (N_1963,N_333,N_826);
or U1964 (N_1964,N_246,N_569);
and U1965 (N_1965,N_311,N_230);
and U1966 (N_1966,N_393,N_310);
nand U1967 (N_1967,N_493,N_424);
nor U1968 (N_1968,N_868,N_436);
nand U1969 (N_1969,N_239,N_469);
or U1970 (N_1970,N_443,N_975);
or U1971 (N_1971,N_79,N_570);
nor U1972 (N_1972,N_506,N_333);
nor U1973 (N_1973,N_653,N_650);
xor U1974 (N_1974,N_377,N_148);
or U1975 (N_1975,N_974,N_50);
nor U1976 (N_1976,N_470,N_459);
nand U1977 (N_1977,N_949,N_444);
nor U1978 (N_1978,N_470,N_469);
and U1979 (N_1979,N_703,N_830);
xnor U1980 (N_1980,N_292,N_151);
nor U1981 (N_1981,N_755,N_684);
nor U1982 (N_1982,N_593,N_662);
and U1983 (N_1983,N_203,N_493);
nand U1984 (N_1984,N_880,N_768);
and U1985 (N_1985,N_572,N_919);
or U1986 (N_1986,N_120,N_350);
nor U1987 (N_1987,N_330,N_517);
nand U1988 (N_1988,N_550,N_455);
or U1989 (N_1989,N_493,N_267);
nor U1990 (N_1990,N_490,N_416);
nand U1991 (N_1991,N_475,N_329);
or U1992 (N_1992,N_830,N_26);
or U1993 (N_1993,N_606,N_785);
or U1994 (N_1994,N_659,N_439);
nand U1995 (N_1995,N_752,N_994);
nand U1996 (N_1996,N_761,N_322);
nor U1997 (N_1997,N_700,N_279);
or U1998 (N_1998,N_569,N_996);
and U1999 (N_1999,N_278,N_167);
xor U2000 (N_2000,N_1274,N_1134);
and U2001 (N_2001,N_1273,N_1385);
or U2002 (N_2002,N_1693,N_1847);
or U2003 (N_2003,N_1738,N_1216);
nor U2004 (N_2004,N_1992,N_1700);
or U2005 (N_2005,N_1282,N_1776);
and U2006 (N_2006,N_1380,N_1978);
nand U2007 (N_2007,N_1042,N_1874);
and U2008 (N_2008,N_1606,N_1523);
nor U2009 (N_2009,N_1304,N_1104);
and U2010 (N_2010,N_1245,N_1563);
and U2011 (N_2011,N_1475,N_1399);
and U2012 (N_2012,N_1244,N_1118);
and U2013 (N_2013,N_1966,N_1132);
or U2014 (N_2014,N_1911,N_1593);
nor U2015 (N_2015,N_1542,N_1567);
nand U2016 (N_2016,N_1988,N_1967);
nor U2017 (N_2017,N_1278,N_1692);
nor U2018 (N_2018,N_1075,N_1708);
or U2019 (N_2019,N_1236,N_1972);
nand U2020 (N_2020,N_1286,N_1528);
nand U2021 (N_2021,N_1111,N_1049);
nand U2022 (N_2022,N_1004,N_1177);
or U2023 (N_2023,N_1262,N_1797);
or U2024 (N_2024,N_1509,N_1342);
nor U2025 (N_2025,N_1726,N_1062);
nand U2026 (N_2026,N_1897,N_1570);
nor U2027 (N_2027,N_1665,N_1362);
xor U2028 (N_2028,N_1853,N_1840);
or U2029 (N_2029,N_1101,N_1289);
nand U2030 (N_2030,N_1651,N_1139);
nor U2031 (N_2031,N_1766,N_1729);
nand U2032 (N_2032,N_1389,N_1355);
nor U2033 (N_2033,N_1646,N_1209);
nand U2034 (N_2034,N_1346,N_1571);
and U2035 (N_2035,N_1223,N_1553);
nand U2036 (N_2036,N_1750,N_1788);
nand U2037 (N_2037,N_1085,N_1800);
nor U2038 (N_2038,N_1161,N_1395);
or U2039 (N_2039,N_1224,N_1029);
or U2040 (N_2040,N_1562,N_1271);
xor U2041 (N_2041,N_1295,N_1817);
nor U2042 (N_2042,N_1576,N_1564);
nor U2043 (N_2043,N_1277,N_1283);
nor U2044 (N_2044,N_1065,N_1926);
nand U2045 (N_2045,N_1000,N_1543);
xnor U2046 (N_2046,N_1883,N_1525);
or U2047 (N_2047,N_1672,N_1153);
nand U2048 (N_2048,N_1255,N_1353);
nand U2049 (N_2049,N_1504,N_1269);
or U2050 (N_2050,N_1934,N_1674);
or U2051 (N_2051,N_1705,N_1151);
or U2052 (N_2052,N_1707,N_1035);
and U2053 (N_2053,N_1260,N_1136);
nor U2054 (N_2054,N_1411,N_1036);
or U2055 (N_2055,N_1345,N_1302);
or U2056 (N_2056,N_1586,N_1622);
nand U2057 (N_2057,N_1179,N_1751);
nor U2058 (N_2058,N_1691,N_1069);
and U2059 (N_2059,N_1818,N_1435);
xor U2060 (N_2060,N_1256,N_1092);
or U2061 (N_2061,N_1011,N_1820);
nor U2062 (N_2062,N_1902,N_1514);
nor U2063 (N_2063,N_1696,N_1763);
or U2064 (N_2064,N_1604,N_1685);
nor U2065 (N_2065,N_1814,N_1057);
nand U2066 (N_2066,N_1303,N_1520);
nand U2067 (N_2067,N_1076,N_1601);
and U2068 (N_2068,N_1965,N_1762);
nor U2069 (N_2069,N_1100,N_1739);
and U2070 (N_2070,N_1610,N_1094);
and U2071 (N_2071,N_1550,N_1581);
nor U2072 (N_2072,N_1272,N_1025);
nand U2073 (N_2073,N_1807,N_1854);
nor U2074 (N_2074,N_1861,N_1426);
or U2075 (N_2075,N_1229,N_1595);
or U2076 (N_2076,N_1888,N_1958);
nand U2077 (N_2077,N_1145,N_1645);
nor U2078 (N_2078,N_1243,N_1322);
xor U2079 (N_2079,N_1228,N_1241);
and U2080 (N_2080,N_1333,N_1009);
nand U2081 (N_2081,N_1579,N_1433);
xor U2082 (N_2082,N_1515,N_1876);
nor U2083 (N_2083,N_1044,N_1440);
nand U2084 (N_2084,N_1073,N_1001);
nor U2085 (N_2085,N_1276,N_1975);
nand U2086 (N_2086,N_1313,N_1508);
nor U2087 (N_2087,N_1232,N_1784);
or U2088 (N_2088,N_1741,N_1352);
nand U2089 (N_2089,N_1275,N_1795);
nand U2090 (N_2090,N_1072,N_1698);
or U2091 (N_2091,N_1777,N_1006);
nand U2092 (N_2092,N_1884,N_1656);
nor U2093 (N_2093,N_1721,N_1590);
or U2094 (N_2094,N_1845,N_1825);
nand U2095 (N_2095,N_1003,N_1976);
nor U2096 (N_2096,N_1425,N_1328);
or U2097 (N_2097,N_1218,N_1742);
or U2098 (N_2098,N_1964,N_1048);
nor U2099 (N_2099,N_1625,N_1891);
and U2100 (N_2100,N_1752,N_1439);
and U2101 (N_2101,N_1143,N_1414);
or U2102 (N_2102,N_1026,N_1372);
or U2103 (N_2103,N_1238,N_1248);
nand U2104 (N_2104,N_1673,N_1116);
xor U2105 (N_2105,N_1924,N_1718);
xor U2106 (N_2106,N_1174,N_1533);
nor U2107 (N_2107,N_1046,N_1420);
and U2108 (N_2108,N_1931,N_1841);
nand U2109 (N_2109,N_1501,N_1242);
and U2110 (N_2110,N_1753,N_1996);
xnor U2111 (N_2111,N_1526,N_1666);
nor U2112 (N_2112,N_1253,N_1112);
xor U2113 (N_2113,N_1982,N_1649);
nand U2114 (N_2114,N_1252,N_1157);
nor U2115 (N_2115,N_1909,N_1442);
or U2116 (N_2116,N_1343,N_1944);
nand U2117 (N_2117,N_1540,N_1704);
or U2118 (N_2118,N_1811,N_1192);
and U2119 (N_2119,N_1415,N_1205);
and U2120 (N_2120,N_1714,N_1320);
nand U2121 (N_2121,N_1031,N_1109);
and U2122 (N_2122,N_1667,N_1872);
and U2123 (N_2123,N_1279,N_1749);
xnor U2124 (N_2124,N_1530,N_1558);
and U2125 (N_2125,N_1827,N_1050);
nand U2126 (N_2126,N_1037,N_1487);
nand U2127 (N_2127,N_1324,N_1246);
nor U2128 (N_2128,N_1808,N_1516);
nor U2129 (N_2129,N_1456,N_1974);
nor U2130 (N_2130,N_1512,N_1358);
nor U2131 (N_2131,N_1392,N_1312);
nor U2132 (N_2132,N_1577,N_1844);
and U2133 (N_2133,N_1316,N_1664);
and U2134 (N_2134,N_1306,N_1309);
and U2135 (N_2135,N_1668,N_1162);
and U2136 (N_2136,N_1418,N_1067);
and U2137 (N_2137,N_1915,N_1930);
nand U2138 (N_2138,N_1722,N_1142);
nor U2139 (N_2139,N_1490,N_1794);
and U2140 (N_2140,N_1497,N_1801);
or U2141 (N_2141,N_1918,N_1556);
nor U2142 (N_2142,N_1933,N_1292);
nor U2143 (N_2143,N_1922,N_1819);
nand U2144 (N_2144,N_1837,N_1194);
and U2145 (N_2145,N_1637,N_1616);
nand U2146 (N_2146,N_1431,N_1864);
nor U2147 (N_2147,N_1311,N_1619);
nand U2148 (N_2148,N_1419,N_1164);
and U2149 (N_2149,N_1678,N_1724);
nor U2150 (N_2150,N_1125,N_1899);
xor U2151 (N_2151,N_1652,N_1942);
and U2152 (N_2152,N_1458,N_1921);
or U2153 (N_2153,N_1261,N_1429);
and U2154 (N_2154,N_1310,N_1226);
nor U2155 (N_2155,N_1824,N_1920);
or U2156 (N_2156,N_1812,N_1386);
and U2157 (N_2157,N_1175,N_1621);
xnor U2158 (N_2158,N_1599,N_1822);
or U2159 (N_2159,N_1291,N_1641);
nand U2160 (N_2160,N_1815,N_1603);
nand U2161 (N_2161,N_1082,N_1554);
xor U2162 (N_2162,N_1199,N_1983);
nor U2163 (N_2163,N_1779,N_1488);
or U2164 (N_2164,N_1133,N_1197);
or U2165 (N_2165,N_1400,N_1417);
or U2166 (N_2166,N_1019,N_1064);
nor U2167 (N_2167,N_1171,N_1321);
or U2168 (N_2168,N_1755,N_1013);
or U2169 (N_2169,N_1541,N_1941);
xnor U2170 (N_2170,N_1235,N_1890);
or U2171 (N_2171,N_1258,N_1217);
and U2172 (N_2172,N_1878,N_1331);
and U2173 (N_2173,N_1908,N_1998);
or U2174 (N_2174,N_1764,N_1823);
or U2175 (N_2175,N_1589,N_1860);
or U2176 (N_2176,N_1745,N_1719);
or U2177 (N_2177,N_1551,N_1068);
nor U2178 (N_2178,N_1786,N_1225);
xnor U2179 (N_2179,N_1137,N_1913);
nor U2180 (N_2180,N_1427,N_1140);
nor U2181 (N_2181,N_1731,N_1979);
and U2182 (N_2182,N_1020,N_1478);
nand U2183 (N_2183,N_1880,N_1809);
nand U2184 (N_2184,N_1981,N_1098);
and U2185 (N_2185,N_1444,N_1097);
nand U2186 (N_2186,N_1240,N_1344);
nor U2187 (N_2187,N_1428,N_1829);
xor U2188 (N_2188,N_1851,N_1572);
or U2189 (N_2189,N_1655,N_1802);
and U2190 (N_2190,N_1620,N_1074);
xnor U2191 (N_2191,N_1059,N_1263);
and U2192 (N_2192,N_1122,N_1916);
nor U2193 (N_2193,N_1632,N_1239);
nand U2194 (N_2194,N_1297,N_1498);
nand U2195 (N_2195,N_1191,N_1496);
xor U2196 (N_2196,N_1334,N_1204);
and U2197 (N_2197,N_1128,N_1299);
or U2198 (N_2198,N_1212,N_1464);
xnor U2199 (N_2199,N_1394,N_1524);
nor U2200 (N_2200,N_1120,N_1511);
nor U2201 (N_2201,N_1901,N_1538);
xnor U2202 (N_2202,N_1871,N_1626);
and U2203 (N_2203,N_1643,N_1267);
nor U2204 (N_2204,N_1083,N_1017);
or U2205 (N_2205,N_1155,N_1758);
nand U2206 (N_2206,N_1452,N_1351);
and U2207 (N_2207,N_1557,N_1642);
or U2208 (N_2208,N_1135,N_1898);
and U2209 (N_2209,N_1066,N_1335);
and U2210 (N_2210,N_1560,N_1396);
nand U2211 (N_2211,N_1935,N_1744);
nor U2212 (N_2212,N_1437,N_1183);
nor U2213 (N_2213,N_1713,N_1349);
xnor U2214 (N_2214,N_1091,N_1519);
nand U2215 (N_2215,N_1894,N_1058);
nor U2216 (N_2216,N_1014,N_1465);
and U2217 (N_2217,N_1990,N_1917);
nor U2218 (N_2218,N_1222,N_1866);
or U2219 (N_2219,N_1919,N_1369);
or U2220 (N_2220,N_1482,N_1506);
and U2221 (N_2221,N_1585,N_1522);
nor U2222 (N_2222,N_1141,N_1843);
xnor U2223 (N_2223,N_1736,N_1398);
nor U2224 (N_2224,N_1627,N_1434);
or U2225 (N_2225,N_1018,N_1461);
nand U2226 (N_2226,N_1720,N_1865);
nor U2227 (N_2227,N_1022,N_1886);
and U2228 (N_2228,N_1393,N_1293);
or U2229 (N_2229,N_1485,N_1796);
nor U2230 (N_2230,N_1359,N_1466);
nor U2231 (N_2231,N_1914,N_1079);
nor U2232 (N_2232,N_1756,N_1454);
nand U2233 (N_2233,N_1448,N_1340);
and U2234 (N_2234,N_1500,N_1163);
nand U2235 (N_2235,N_1250,N_1450);
and U2236 (N_2236,N_1638,N_1687);
and U2237 (N_2237,N_1798,N_1378);
nor U2238 (N_2238,N_1290,N_1280);
nand U2239 (N_2239,N_1680,N_1858);
nor U2240 (N_2240,N_1662,N_1928);
or U2241 (N_2241,N_1361,N_1634);
nand U2242 (N_2242,N_1390,N_1657);
nor U2243 (N_2243,N_1727,N_1221);
or U2244 (N_2244,N_1489,N_1539);
nand U2245 (N_2245,N_1503,N_1517);
or U2246 (N_2246,N_1008,N_1181);
nand U2247 (N_2247,N_1451,N_1970);
or U2248 (N_2248,N_1857,N_1937);
nor U2249 (N_2249,N_1071,N_1336);
nand U2250 (N_2250,N_1455,N_1952);
xor U2251 (N_2251,N_1005,N_1987);
nand U2252 (N_2252,N_1357,N_1318);
and U2253 (N_2253,N_1605,N_1534);
nand U2254 (N_2254,N_1715,N_1617);
and U2255 (N_2255,N_1633,N_1281);
nor U2256 (N_2256,N_1374,N_1587);
and U2257 (N_2257,N_1129,N_1828);
nor U2258 (N_2258,N_1614,N_1214);
and U2259 (N_2259,N_1149,N_1184);
nor U2260 (N_2260,N_1778,N_1999);
and U2261 (N_2261,N_1231,N_1470);
or U2262 (N_2262,N_1669,N_1946);
nand U2263 (N_2263,N_1733,N_1821);
and U2264 (N_2264,N_1201,N_1315);
nor U2265 (N_2265,N_1077,N_1015);
or U2266 (N_2266,N_1771,N_1927);
or U2267 (N_2267,N_1939,N_1237);
xnor U2268 (N_2268,N_1033,N_1198);
and U2269 (N_2269,N_1326,N_1573);
nand U2270 (N_2270,N_1936,N_1555);
and U2271 (N_2271,N_1636,N_1086);
or U2272 (N_2272,N_1407,N_1032);
and U2273 (N_2273,N_1505,N_1409);
nor U2274 (N_2274,N_1810,N_1227);
xor U2275 (N_2275,N_1147,N_1117);
nand U2276 (N_2276,N_1115,N_1760);
and U2277 (N_2277,N_1055,N_1391);
nand U2278 (N_2278,N_1618,N_1518);
or U2279 (N_2279,N_1484,N_1087);
and U2280 (N_2280,N_1559,N_1070);
or U2281 (N_2281,N_1723,N_1896);
nand U2282 (N_2282,N_1659,N_1826);
and U2283 (N_2283,N_1681,N_1699);
nor U2284 (N_2284,N_1986,N_1124);
nor U2285 (N_2285,N_1023,N_1773);
nand U2286 (N_2286,N_1196,N_1043);
and U2287 (N_2287,N_1943,N_1364);
xnor U2288 (N_2288,N_1188,N_1210);
nand U2289 (N_2289,N_1735,N_1167);
and U2290 (N_2290,N_1850,N_1010);
nand U2291 (N_2291,N_1690,N_1354);
nor U2292 (N_2292,N_1973,N_1499);
and U2293 (N_2293,N_1200,N_1994);
nor U2294 (N_2294,N_1257,N_1329);
and U2295 (N_2295,N_1156,N_1449);
nand U2296 (N_2296,N_1775,N_1106);
and U2297 (N_2297,N_1102,N_1379);
nand U2298 (N_2298,N_1984,N_1813);
and U2299 (N_2299,N_1038,N_1701);
xor U2300 (N_2300,N_1548,N_1189);
nand U2301 (N_2301,N_1863,N_1028);
nor U2302 (N_2302,N_1296,N_1314);
or U2303 (N_2303,N_1305,N_1549);
nor U2304 (N_2304,N_1711,N_1144);
nand U2305 (N_2305,N_1365,N_1830);
and U2306 (N_2306,N_1373,N_1307);
nor U2307 (N_2307,N_1495,N_1095);
and U2308 (N_2308,N_1300,N_1350);
nor U2309 (N_2309,N_1404,N_1639);
nand U2310 (N_2310,N_1932,N_1940);
nand U2311 (N_2311,N_1848,N_1836);
nand U2312 (N_2312,N_1447,N_1578);
xnor U2313 (N_2313,N_1640,N_1105);
nand U2314 (N_2314,N_1774,N_1607);
nor U2315 (N_2315,N_1012,N_1780);
nand U2316 (N_2316,N_1045,N_1462);
and U2317 (N_2317,N_1873,N_1410);
and U2318 (N_2318,N_1476,N_1234);
and U2319 (N_2319,N_1725,N_1165);
nand U2320 (N_2320,N_1051,N_1989);
and U2321 (N_2321,N_1002,N_1383);
nand U2322 (N_2322,N_1259,N_1471);
nor U2323 (N_2323,N_1623,N_1804);
nor U2324 (N_2324,N_1961,N_1953);
nor U2325 (N_2325,N_1039,N_1180);
nand U2326 (N_2326,N_1403,N_1185);
and U2327 (N_2327,N_1945,N_1955);
or U2328 (N_2328,N_1592,N_1481);
xnor U2329 (N_2329,N_1903,N_1099);
and U2330 (N_2330,N_1925,N_1376);
or U2331 (N_2331,N_1388,N_1759);
and U2332 (N_2332,N_1472,N_1416);
nand U2333 (N_2333,N_1695,N_1624);
nand U2334 (N_2334,N_1980,N_1532);
nand U2335 (N_2335,N_1513,N_1436);
and U2336 (N_2336,N_1170,N_1993);
nor U2337 (N_2337,N_1893,N_1337);
nor U2338 (N_2338,N_1682,N_1007);
nand U2339 (N_2339,N_1991,N_1747);
nor U2340 (N_2340,N_1561,N_1628);
and U2341 (N_2341,N_1088,N_1768);
or U2342 (N_2342,N_1904,N_1284);
or U2343 (N_2343,N_1096,N_1670);
nor U2344 (N_2344,N_1108,N_1658);
nor U2345 (N_2345,N_1566,N_1889);
and U2346 (N_2346,N_1702,N_1787);
nor U2347 (N_2347,N_1270,N_1839);
and U2348 (N_2348,N_1703,N_1612);
and U2349 (N_2349,N_1849,N_1650);
or U2350 (N_2350,N_1089,N_1629);
or U2351 (N_2351,N_1594,N_1406);
nor U2352 (N_2352,N_1178,N_1093);
nor U2353 (N_2353,N_1547,N_1441);
or U2354 (N_2354,N_1568,N_1148);
and U2355 (N_2355,N_1377,N_1971);
or U2356 (N_2356,N_1772,N_1677);
and U2357 (N_2357,N_1368,N_1956);
nand U2358 (N_2358,N_1047,N_1600);
nand U2359 (N_2359,N_1203,N_1885);
nand U2360 (N_2360,N_1569,N_1319);
nor U2361 (N_2361,N_1957,N_1247);
xor U2362 (N_2362,N_1912,N_1190);
nor U2363 (N_2363,N_1789,N_1877);
nor U2364 (N_2364,N_1977,N_1382);
nor U2365 (N_2365,N_1486,N_1867);
nand U2366 (N_2366,N_1215,N_1459);
and U2367 (N_2367,N_1081,N_1938);
nand U2368 (N_2368,N_1831,N_1905);
nand U2369 (N_2369,N_1159,N_1325);
nor U2370 (N_2370,N_1408,N_1882);
and U2371 (N_2371,N_1536,N_1732);
xnor U2372 (N_2372,N_1679,N_1502);
nand U2373 (N_2373,N_1997,N_1683);
nand U2374 (N_2374,N_1929,N_1816);
nand U2375 (N_2375,N_1220,N_1338);
and U2376 (N_2376,N_1483,N_1492);
xnor U2377 (N_2377,N_1962,N_1717);
nor U2378 (N_2378,N_1761,N_1054);
nor U2379 (N_2379,N_1308,N_1949);
nand U2380 (N_2380,N_1947,N_1544);
and U2381 (N_2381,N_1401,N_1584);
nor U2382 (N_2382,N_1480,N_1963);
and U2383 (N_2383,N_1611,N_1413);
nand U2384 (N_2384,N_1366,N_1056);
or U2385 (N_2385,N_1127,N_1661);
nand U2386 (N_2386,N_1716,N_1445);
and U2387 (N_2387,N_1743,N_1521);
or U2388 (N_2388,N_1152,N_1613);
or U2389 (N_2389,N_1090,N_1684);
nor U2390 (N_2390,N_1531,N_1881);
nor U2391 (N_2391,N_1948,N_1330);
or U2392 (N_2392,N_1608,N_1663);
and U2393 (N_2393,N_1412,N_1160);
nor U2394 (N_2394,N_1648,N_1833);
or U2395 (N_2395,N_1347,N_1348);
nand U2396 (N_2396,N_1268,N_1832);
nor U2397 (N_2397,N_1609,N_1474);
or U2398 (N_2398,N_1166,N_1468);
and U2399 (N_2399,N_1688,N_1653);
and U2400 (N_2400,N_1080,N_1384);
xnor U2401 (N_2401,N_1781,N_1107);
nand U2402 (N_2402,N_1529,N_1545);
nor U2403 (N_2403,N_1219,N_1078);
or U2404 (N_2404,N_1438,N_1341);
nor U2405 (N_2405,N_1130,N_1317);
xnor U2406 (N_2406,N_1630,N_1799);
or U2407 (N_2407,N_1387,N_1491);
nand U2408 (N_2408,N_1375,N_1697);
nand U2409 (N_2409,N_1838,N_1770);
nor U2410 (N_2410,N_1785,N_1862);
and U2411 (N_2411,N_1363,N_1654);
or U2412 (N_2412,N_1249,N_1537);
or U2413 (N_2413,N_1792,N_1782);
and U2414 (N_2414,N_1602,N_1169);
nor U2415 (N_2415,N_1575,N_1327);
or U2416 (N_2416,N_1887,N_1367);
xor U2417 (N_2417,N_1154,N_1405);
nor U2418 (N_2418,N_1016,N_1467);
and U2419 (N_2419,N_1846,N_1676);
nand U2420 (N_2420,N_1493,N_1615);
and U2421 (N_2421,N_1879,N_1479);
nand U2422 (N_2422,N_1113,N_1182);
or U2423 (N_2423,N_1790,N_1264);
nor U2424 (N_2424,N_1146,N_1686);
nand U2425 (N_2425,N_1710,N_1868);
nand U2426 (N_2426,N_1875,N_1951);
nor U2427 (N_2427,N_1423,N_1172);
nand U2428 (N_2428,N_1114,N_1859);
nor U2429 (N_2429,N_1754,N_1126);
nor U2430 (N_2430,N_1168,N_1061);
nand U2431 (N_2431,N_1959,N_1208);
and U2432 (N_2432,N_1734,N_1737);
and U2433 (N_2433,N_1598,N_1583);
nand U2434 (N_2434,N_1202,N_1791);
or U2435 (N_2435,N_1211,N_1855);
xnor U2436 (N_2436,N_1034,N_1892);
and U2437 (N_2437,N_1193,N_1206);
nor U2438 (N_2438,N_1803,N_1907);
or U2439 (N_2439,N_1580,N_1360);
nand U2440 (N_2440,N_1460,N_1052);
and U2441 (N_2441,N_1402,N_1371);
nor U2442 (N_2442,N_1103,N_1421);
nand U2443 (N_2443,N_1432,N_1463);
and U2444 (N_2444,N_1631,N_1027);
and U2445 (N_2445,N_1430,N_1596);
and U2446 (N_2446,N_1370,N_1647);
nor U2447 (N_2447,N_1469,N_1024);
nor U2448 (N_2448,N_1453,N_1207);
and U2449 (N_2449,N_1588,N_1969);
and U2450 (N_2450,N_1535,N_1287);
nand U2451 (N_2451,N_1793,N_1150);
and U2452 (N_2452,N_1186,N_1123);
and U2453 (N_2453,N_1381,N_1121);
nand U2454 (N_2454,N_1869,N_1254);
nor U2455 (N_2455,N_1757,N_1689);
or U2456 (N_2456,N_1954,N_1834);
nand U2457 (N_2457,N_1187,N_1709);
xnor U2458 (N_2458,N_1805,N_1852);
and U2459 (N_2459,N_1230,N_1176);
and U2460 (N_2460,N_1856,N_1694);
nor U2461 (N_2461,N_1728,N_1063);
xor U2462 (N_2462,N_1084,N_1356);
and U2463 (N_2463,N_1910,N_1546);
nor U2464 (N_2464,N_1294,N_1397);
xor U2465 (N_2465,N_1060,N_1675);
nand U2466 (N_2466,N_1158,N_1213);
or U2467 (N_2467,N_1494,N_1053);
nand U2468 (N_2468,N_1298,N_1740);
nor U2469 (N_2469,N_1030,N_1968);
and U2470 (N_2470,N_1510,N_1233);
nor U2471 (N_2471,N_1195,N_1285);
nor U2472 (N_2472,N_1923,N_1473);
and U2473 (N_2473,N_1706,N_1138);
or U2474 (N_2474,N_1960,N_1597);
or U2475 (N_2475,N_1842,N_1041);
or U2476 (N_2476,N_1835,N_1131);
nand U2477 (N_2477,N_1288,N_1339);
nand U2478 (N_2478,N_1332,N_1021);
and U2479 (N_2479,N_1660,N_1110);
nor U2480 (N_2480,N_1806,N_1635);
and U2481 (N_2481,N_1765,N_1748);
or U2482 (N_2482,N_1565,N_1950);
nor U2483 (N_2483,N_1671,N_1895);
nor U2484 (N_2484,N_1900,N_1985);
and U2485 (N_2485,N_1783,N_1527);
or U2486 (N_2486,N_1443,N_1906);
or U2487 (N_2487,N_1251,N_1552);
nand U2488 (N_2488,N_1769,N_1422);
nand U2489 (N_2489,N_1582,N_1173);
or U2490 (N_2490,N_1870,N_1574);
and U2491 (N_2491,N_1730,N_1301);
and U2492 (N_2492,N_1265,N_1477);
and U2493 (N_2493,N_1424,N_1644);
xnor U2494 (N_2494,N_1712,N_1457);
nor U2495 (N_2495,N_1995,N_1323);
nor U2496 (N_2496,N_1746,N_1507);
nand U2497 (N_2497,N_1266,N_1040);
and U2498 (N_2498,N_1446,N_1119);
nand U2499 (N_2499,N_1591,N_1767);
and U2500 (N_2500,N_1122,N_1679);
or U2501 (N_2501,N_1995,N_1430);
nor U2502 (N_2502,N_1336,N_1018);
or U2503 (N_2503,N_1434,N_1902);
and U2504 (N_2504,N_1087,N_1058);
nand U2505 (N_2505,N_1997,N_1858);
and U2506 (N_2506,N_1533,N_1639);
nand U2507 (N_2507,N_1560,N_1338);
and U2508 (N_2508,N_1270,N_1090);
nand U2509 (N_2509,N_1287,N_1267);
nor U2510 (N_2510,N_1742,N_1922);
or U2511 (N_2511,N_1580,N_1753);
nor U2512 (N_2512,N_1628,N_1901);
nor U2513 (N_2513,N_1410,N_1380);
and U2514 (N_2514,N_1529,N_1137);
and U2515 (N_2515,N_1859,N_1573);
nor U2516 (N_2516,N_1523,N_1206);
or U2517 (N_2517,N_1133,N_1790);
nor U2518 (N_2518,N_1253,N_1580);
or U2519 (N_2519,N_1397,N_1764);
or U2520 (N_2520,N_1778,N_1472);
nand U2521 (N_2521,N_1530,N_1447);
xor U2522 (N_2522,N_1529,N_1676);
and U2523 (N_2523,N_1935,N_1351);
nor U2524 (N_2524,N_1768,N_1892);
nand U2525 (N_2525,N_1198,N_1364);
nand U2526 (N_2526,N_1125,N_1415);
xnor U2527 (N_2527,N_1910,N_1981);
and U2528 (N_2528,N_1846,N_1974);
and U2529 (N_2529,N_1600,N_1933);
nand U2530 (N_2530,N_1128,N_1328);
nand U2531 (N_2531,N_1697,N_1534);
nor U2532 (N_2532,N_1794,N_1492);
nor U2533 (N_2533,N_1766,N_1567);
xnor U2534 (N_2534,N_1254,N_1917);
or U2535 (N_2535,N_1944,N_1401);
nand U2536 (N_2536,N_1172,N_1922);
nor U2537 (N_2537,N_1602,N_1279);
nor U2538 (N_2538,N_1100,N_1705);
or U2539 (N_2539,N_1302,N_1887);
and U2540 (N_2540,N_1319,N_1175);
or U2541 (N_2541,N_1186,N_1848);
nor U2542 (N_2542,N_1482,N_1614);
nand U2543 (N_2543,N_1534,N_1808);
nor U2544 (N_2544,N_1395,N_1152);
nor U2545 (N_2545,N_1366,N_1487);
nor U2546 (N_2546,N_1758,N_1362);
xnor U2547 (N_2547,N_1293,N_1086);
and U2548 (N_2548,N_1052,N_1915);
and U2549 (N_2549,N_1434,N_1586);
or U2550 (N_2550,N_1451,N_1717);
nand U2551 (N_2551,N_1905,N_1119);
nor U2552 (N_2552,N_1997,N_1987);
and U2553 (N_2553,N_1694,N_1692);
nor U2554 (N_2554,N_1737,N_1209);
or U2555 (N_2555,N_1585,N_1170);
nor U2556 (N_2556,N_1257,N_1871);
xnor U2557 (N_2557,N_1205,N_1716);
and U2558 (N_2558,N_1476,N_1912);
and U2559 (N_2559,N_1984,N_1841);
xor U2560 (N_2560,N_1923,N_1070);
or U2561 (N_2561,N_1763,N_1679);
and U2562 (N_2562,N_1685,N_1285);
nand U2563 (N_2563,N_1654,N_1322);
and U2564 (N_2564,N_1040,N_1252);
nand U2565 (N_2565,N_1539,N_1528);
and U2566 (N_2566,N_1851,N_1046);
nor U2567 (N_2567,N_1856,N_1339);
or U2568 (N_2568,N_1658,N_1912);
and U2569 (N_2569,N_1461,N_1013);
and U2570 (N_2570,N_1463,N_1482);
xnor U2571 (N_2571,N_1026,N_1877);
and U2572 (N_2572,N_1018,N_1392);
and U2573 (N_2573,N_1781,N_1612);
nand U2574 (N_2574,N_1664,N_1603);
or U2575 (N_2575,N_1431,N_1766);
nand U2576 (N_2576,N_1244,N_1002);
nand U2577 (N_2577,N_1899,N_1101);
or U2578 (N_2578,N_1221,N_1579);
nor U2579 (N_2579,N_1479,N_1182);
xnor U2580 (N_2580,N_1599,N_1941);
and U2581 (N_2581,N_1098,N_1349);
nand U2582 (N_2582,N_1109,N_1648);
and U2583 (N_2583,N_1392,N_1488);
nor U2584 (N_2584,N_1876,N_1790);
or U2585 (N_2585,N_1479,N_1440);
xnor U2586 (N_2586,N_1293,N_1629);
or U2587 (N_2587,N_1673,N_1481);
or U2588 (N_2588,N_1352,N_1938);
and U2589 (N_2589,N_1186,N_1319);
nand U2590 (N_2590,N_1371,N_1164);
or U2591 (N_2591,N_1247,N_1728);
nor U2592 (N_2592,N_1771,N_1237);
nand U2593 (N_2593,N_1936,N_1742);
and U2594 (N_2594,N_1913,N_1724);
nor U2595 (N_2595,N_1135,N_1550);
nor U2596 (N_2596,N_1480,N_1874);
and U2597 (N_2597,N_1375,N_1060);
or U2598 (N_2598,N_1231,N_1310);
and U2599 (N_2599,N_1882,N_1978);
nor U2600 (N_2600,N_1738,N_1880);
nand U2601 (N_2601,N_1515,N_1781);
nor U2602 (N_2602,N_1366,N_1661);
nand U2603 (N_2603,N_1367,N_1835);
or U2604 (N_2604,N_1480,N_1200);
nand U2605 (N_2605,N_1437,N_1655);
nor U2606 (N_2606,N_1949,N_1155);
and U2607 (N_2607,N_1777,N_1135);
nand U2608 (N_2608,N_1826,N_1887);
nor U2609 (N_2609,N_1541,N_1154);
nor U2610 (N_2610,N_1066,N_1447);
or U2611 (N_2611,N_1001,N_1431);
nand U2612 (N_2612,N_1332,N_1012);
or U2613 (N_2613,N_1405,N_1585);
or U2614 (N_2614,N_1346,N_1159);
or U2615 (N_2615,N_1482,N_1069);
and U2616 (N_2616,N_1734,N_1836);
and U2617 (N_2617,N_1979,N_1053);
or U2618 (N_2618,N_1785,N_1783);
nor U2619 (N_2619,N_1631,N_1372);
or U2620 (N_2620,N_1302,N_1789);
and U2621 (N_2621,N_1873,N_1085);
and U2622 (N_2622,N_1907,N_1236);
or U2623 (N_2623,N_1831,N_1151);
nand U2624 (N_2624,N_1112,N_1498);
nand U2625 (N_2625,N_1455,N_1755);
or U2626 (N_2626,N_1563,N_1945);
or U2627 (N_2627,N_1041,N_1115);
nand U2628 (N_2628,N_1202,N_1280);
and U2629 (N_2629,N_1898,N_1791);
nor U2630 (N_2630,N_1961,N_1253);
nand U2631 (N_2631,N_1887,N_1455);
or U2632 (N_2632,N_1699,N_1964);
nand U2633 (N_2633,N_1620,N_1480);
and U2634 (N_2634,N_1839,N_1868);
and U2635 (N_2635,N_1147,N_1435);
nor U2636 (N_2636,N_1641,N_1719);
and U2637 (N_2637,N_1006,N_1318);
and U2638 (N_2638,N_1866,N_1610);
nor U2639 (N_2639,N_1654,N_1552);
or U2640 (N_2640,N_1835,N_1342);
or U2641 (N_2641,N_1310,N_1223);
and U2642 (N_2642,N_1209,N_1016);
or U2643 (N_2643,N_1487,N_1135);
nor U2644 (N_2644,N_1950,N_1300);
nor U2645 (N_2645,N_1133,N_1795);
and U2646 (N_2646,N_1489,N_1774);
and U2647 (N_2647,N_1546,N_1511);
xnor U2648 (N_2648,N_1360,N_1274);
nor U2649 (N_2649,N_1057,N_1593);
nand U2650 (N_2650,N_1762,N_1268);
and U2651 (N_2651,N_1204,N_1826);
xnor U2652 (N_2652,N_1104,N_1919);
xor U2653 (N_2653,N_1751,N_1167);
and U2654 (N_2654,N_1435,N_1626);
or U2655 (N_2655,N_1188,N_1663);
and U2656 (N_2656,N_1256,N_1863);
or U2657 (N_2657,N_1520,N_1146);
and U2658 (N_2658,N_1898,N_1051);
nor U2659 (N_2659,N_1052,N_1459);
or U2660 (N_2660,N_1194,N_1708);
and U2661 (N_2661,N_1550,N_1514);
and U2662 (N_2662,N_1219,N_1614);
and U2663 (N_2663,N_1573,N_1655);
and U2664 (N_2664,N_1573,N_1594);
nand U2665 (N_2665,N_1782,N_1802);
and U2666 (N_2666,N_1831,N_1431);
nor U2667 (N_2667,N_1744,N_1621);
and U2668 (N_2668,N_1991,N_1377);
or U2669 (N_2669,N_1836,N_1812);
nand U2670 (N_2670,N_1216,N_1825);
and U2671 (N_2671,N_1670,N_1428);
nor U2672 (N_2672,N_1808,N_1897);
nor U2673 (N_2673,N_1857,N_1101);
and U2674 (N_2674,N_1673,N_1763);
xor U2675 (N_2675,N_1750,N_1503);
and U2676 (N_2676,N_1063,N_1636);
or U2677 (N_2677,N_1867,N_1891);
and U2678 (N_2678,N_1388,N_1130);
and U2679 (N_2679,N_1695,N_1358);
or U2680 (N_2680,N_1530,N_1247);
and U2681 (N_2681,N_1988,N_1574);
nor U2682 (N_2682,N_1322,N_1587);
nor U2683 (N_2683,N_1831,N_1133);
nand U2684 (N_2684,N_1104,N_1142);
or U2685 (N_2685,N_1699,N_1867);
nor U2686 (N_2686,N_1141,N_1027);
and U2687 (N_2687,N_1688,N_1770);
or U2688 (N_2688,N_1934,N_1751);
or U2689 (N_2689,N_1401,N_1507);
and U2690 (N_2690,N_1451,N_1663);
or U2691 (N_2691,N_1187,N_1568);
nor U2692 (N_2692,N_1666,N_1848);
xor U2693 (N_2693,N_1446,N_1190);
and U2694 (N_2694,N_1051,N_1347);
nor U2695 (N_2695,N_1816,N_1316);
nand U2696 (N_2696,N_1220,N_1173);
and U2697 (N_2697,N_1366,N_1764);
xor U2698 (N_2698,N_1911,N_1974);
nor U2699 (N_2699,N_1761,N_1148);
nand U2700 (N_2700,N_1240,N_1973);
nand U2701 (N_2701,N_1905,N_1166);
nor U2702 (N_2702,N_1697,N_1918);
nand U2703 (N_2703,N_1382,N_1985);
or U2704 (N_2704,N_1753,N_1043);
or U2705 (N_2705,N_1413,N_1873);
nor U2706 (N_2706,N_1762,N_1889);
xnor U2707 (N_2707,N_1481,N_1037);
xnor U2708 (N_2708,N_1156,N_1491);
nand U2709 (N_2709,N_1240,N_1965);
or U2710 (N_2710,N_1117,N_1139);
xnor U2711 (N_2711,N_1693,N_1605);
or U2712 (N_2712,N_1066,N_1123);
and U2713 (N_2713,N_1274,N_1538);
nor U2714 (N_2714,N_1430,N_1099);
xnor U2715 (N_2715,N_1746,N_1788);
nor U2716 (N_2716,N_1762,N_1438);
nand U2717 (N_2717,N_1410,N_1748);
xnor U2718 (N_2718,N_1255,N_1254);
or U2719 (N_2719,N_1509,N_1373);
and U2720 (N_2720,N_1450,N_1073);
and U2721 (N_2721,N_1084,N_1581);
nand U2722 (N_2722,N_1393,N_1613);
and U2723 (N_2723,N_1153,N_1409);
nand U2724 (N_2724,N_1979,N_1672);
and U2725 (N_2725,N_1044,N_1483);
nor U2726 (N_2726,N_1239,N_1083);
or U2727 (N_2727,N_1746,N_1476);
and U2728 (N_2728,N_1335,N_1617);
or U2729 (N_2729,N_1233,N_1685);
nand U2730 (N_2730,N_1845,N_1589);
or U2731 (N_2731,N_1885,N_1313);
or U2732 (N_2732,N_1465,N_1125);
and U2733 (N_2733,N_1131,N_1500);
nand U2734 (N_2734,N_1734,N_1090);
or U2735 (N_2735,N_1125,N_1793);
and U2736 (N_2736,N_1896,N_1230);
nand U2737 (N_2737,N_1173,N_1382);
nor U2738 (N_2738,N_1808,N_1490);
nor U2739 (N_2739,N_1630,N_1382);
nor U2740 (N_2740,N_1424,N_1346);
nor U2741 (N_2741,N_1366,N_1395);
nor U2742 (N_2742,N_1246,N_1442);
and U2743 (N_2743,N_1778,N_1485);
and U2744 (N_2744,N_1392,N_1628);
xnor U2745 (N_2745,N_1113,N_1032);
or U2746 (N_2746,N_1466,N_1048);
or U2747 (N_2747,N_1234,N_1867);
xnor U2748 (N_2748,N_1718,N_1034);
and U2749 (N_2749,N_1541,N_1679);
and U2750 (N_2750,N_1178,N_1335);
nand U2751 (N_2751,N_1348,N_1357);
or U2752 (N_2752,N_1000,N_1016);
xor U2753 (N_2753,N_1144,N_1008);
or U2754 (N_2754,N_1085,N_1173);
or U2755 (N_2755,N_1176,N_1083);
nand U2756 (N_2756,N_1695,N_1731);
and U2757 (N_2757,N_1630,N_1880);
and U2758 (N_2758,N_1185,N_1886);
nor U2759 (N_2759,N_1346,N_1799);
nand U2760 (N_2760,N_1603,N_1012);
or U2761 (N_2761,N_1912,N_1880);
nor U2762 (N_2762,N_1536,N_1528);
nand U2763 (N_2763,N_1885,N_1530);
or U2764 (N_2764,N_1485,N_1530);
or U2765 (N_2765,N_1142,N_1559);
and U2766 (N_2766,N_1847,N_1191);
xnor U2767 (N_2767,N_1522,N_1349);
nand U2768 (N_2768,N_1932,N_1621);
or U2769 (N_2769,N_1454,N_1172);
or U2770 (N_2770,N_1164,N_1449);
and U2771 (N_2771,N_1256,N_1514);
nor U2772 (N_2772,N_1189,N_1967);
nor U2773 (N_2773,N_1282,N_1349);
or U2774 (N_2774,N_1656,N_1472);
or U2775 (N_2775,N_1500,N_1783);
nor U2776 (N_2776,N_1963,N_1451);
nand U2777 (N_2777,N_1191,N_1617);
nor U2778 (N_2778,N_1651,N_1799);
and U2779 (N_2779,N_1833,N_1623);
nor U2780 (N_2780,N_1945,N_1198);
nor U2781 (N_2781,N_1497,N_1982);
and U2782 (N_2782,N_1998,N_1853);
nand U2783 (N_2783,N_1094,N_1826);
nand U2784 (N_2784,N_1155,N_1549);
and U2785 (N_2785,N_1696,N_1860);
or U2786 (N_2786,N_1067,N_1769);
and U2787 (N_2787,N_1483,N_1549);
nor U2788 (N_2788,N_1662,N_1181);
xnor U2789 (N_2789,N_1332,N_1661);
or U2790 (N_2790,N_1854,N_1389);
nor U2791 (N_2791,N_1743,N_1956);
nand U2792 (N_2792,N_1664,N_1099);
nand U2793 (N_2793,N_1928,N_1919);
nor U2794 (N_2794,N_1723,N_1669);
or U2795 (N_2795,N_1123,N_1070);
nor U2796 (N_2796,N_1894,N_1696);
and U2797 (N_2797,N_1758,N_1067);
nor U2798 (N_2798,N_1187,N_1754);
nor U2799 (N_2799,N_1982,N_1438);
and U2800 (N_2800,N_1766,N_1016);
and U2801 (N_2801,N_1217,N_1359);
nor U2802 (N_2802,N_1058,N_1060);
nor U2803 (N_2803,N_1355,N_1317);
nor U2804 (N_2804,N_1143,N_1420);
or U2805 (N_2805,N_1859,N_1491);
nand U2806 (N_2806,N_1782,N_1615);
or U2807 (N_2807,N_1634,N_1565);
and U2808 (N_2808,N_1021,N_1928);
nor U2809 (N_2809,N_1352,N_1507);
xnor U2810 (N_2810,N_1889,N_1983);
and U2811 (N_2811,N_1428,N_1499);
nand U2812 (N_2812,N_1338,N_1422);
and U2813 (N_2813,N_1349,N_1844);
xnor U2814 (N_2814,N_1869,N_1701);
xor U2815 (N_2815,N_1881,N_1563);
nor U2816 (N_2816,N_1979,N_1254);
nor U2817 (N_2817,N_1310,N_1103);
nor U2818 (N_2818,N_1985,N_1059);
or U2819 (N_2819,N_1254,N_1515);
nor U2820 (N_2820,N_1588,N_1406);
xor U2821 (N_2821,N_1677,N_1889);
and U2822 (N_2822,N_1268,N_1069);
nor U2823 (N_2823,N_1139,N_1352);
or U2824 (N_2824,N_1227,N_1716);
and U2825 (N_2825,N_1978,N_1231);
nand U2826 (N_2826,N_1072,N_1342);
and U2827 (N_2827,N_1535,N_1421);
or U2828 (N_2828,N_1269,N_1530);
nor U2829 (N_2829,N_1816,N_1281);
or U2830 (N_2830,N_1251,N_1533);
xor U2831 (N_2831,N_1140,N_1852);
nand U2832 (N_2832,N_1986,N_1979);
and U2833 (N_2833,N_1607,N_1942);
nand U2834 (N_2834,N_1392,N_1733);
nor U2835 (N_2835,N_1153,N_1546);
or U2836 (N_2836,N_1417,N_1091);
nor U2837 (N_2837,N_1882,N_1758);
nand U2838 (N_2838,N_1154,N_1813);
xor U2839 (N_2839,N_1476,N_1011);
nand U2840 (N_2840,N_1846,N_1471);
nand U2841 (N_2841,N_1010,N_1440);
nor U2842 (N_2842,N_1025,N_1770);
or U2843 (N_2843,N_1280,N_1031);
or U2844 (N_2844,N_1073,N_1658);
xor U2845 (N_2845,N_1574,N_1194);
nand U2846 (N_2846,N_1283,N_1997);
or U2847 (N_2847,N_1954,N_1072);
or U2848 (N_2848,N_1501,N_1962);
and U2849 (N_2849,N_1944,N_1907);
nand U2850 (N_2850,N_1975,N_1823);
nand U2851 (N_2851,N_1030,N_1087);
nor U2852 (N_2852,N_1300,N_1925);
and U2853 (N_2853,N_1282,N_1152);
nor U2854 (N_2854,N_1250,N_1315);
nand U2855 (N_2855,N_1260,N_1397);
and U2856 (N_2856,N_1472,N_1365);
nor U2857 (N_2857,N_1138,N_1754);
and U2858 (N_2858,N_1837,N_1163);
nand U2859 (N_2859,N_1940,N_1670);
nand U2860 (N_2860,N_1055,N_1797);
and U2861 (N_2861,N_1461,N_1356);
nand U2862 (N_2862,N_1046,N_1122);
and U2863 (N_2863,N_1100,N_1641);
and U2864 (N_2864,N_1814,N_1270);
or U2865 (N_2865,N_1039,N_1443);
or U2866 (N_2866,N_1105,N_1863);
nand U2867 (N_2867,N_1306,N_1864);
and U2868 (N_2868,N_1650,N_1729);
xnor U2869 (N_2869,N_1956,N_1517);
or U2870 (N_2870,N_1643,N_1414);
xnor U2871 (N_2871,N_1187,N_1739);
xnor U2872 (N_2872,N_1109,N_1412);
or U2873 (N_2873,N_1171,N_1719);
nand U2874 (N_2874,N_1432,N_1091);
and U2875 (N_2875,N_1268,N_1907);
nor U2876 (N_2876,N_1561,N_1510);
or U2877 (N_2877,N_1551,N_1102);
and U2878 (N_2878,N_1405,N_1787);
or U2879 (N_2879,N_1371,N_1929);
and U2880 (N_2880,N_1039,N_1673);
xor U2881 (N_2881,N_1360,N_1491);
and U2882 (N_2882,N_1666,N_1115);
or U2883 (N_2883,N_1942,N_1542);
nand U2884 (N_2884,N_1396,N_1837);
nor U2885 (N_2885,N_1633,N_1991);
or U2886 (N_2886,N_1426,N_1087);
nor U2887 (N_2887,N_1951,N_1762);
xnor U2888 (N_2888,N_1513,N_1440);
nand U2889 (N_2889,N_1599,N_1215);
and U2890 (N_2890,N_1959,N_1866);
and U2891 (N_2891,N_1195,N_1392);
and U2892 (N_2892,N_1158,N_1576);
xnor U2893 (N_2893,N_1112,N_1214);
or U2894 (N_2894,N_1700,N_1217);
or U2895 (N_2895,N_1826,N_1025);
nand U2896 (N_2896,N_1447,N_1636);
or U2897 (N_2897,N_1219,N_1560);
nor U2898 (N_2898,N_1731,N_1856);
nand U2899 (N_2899,N_1139,N_1439);
and U2900 (N_2900,N_1329,N_1610);
or U2901 (N_2901,N_1264,N_1139);
nand U2902 (N_2902,N_1666,N_1313);
or U2903 (N_2903,N_1816,N_1330);
nand U2904 (N_2904,N_1769,N_1893);
nand U2905 (N_2905,N_1723,N_1917);
or U2906 (N_2906,N_1568,N_1516);
and U2907 (N_2907,N_1057,N_1038);
or U2908 (N_2908,N_1951,N_1727);
nand U2909 (N_2909,N_1919,N_1781);
or U2910 (N_2910,N_1866,N_1870);
nand U2911 (N_2911,N_1702,N_1535);
and U2912 (N_2912,N_1557,N_1833);
nor U2913 (N_2913,N_1141,N_1533);
nand U2914 (N_2914,N_1878,N_1116);
nand U2915 (N_2915,N_1084,N_1218);
nor U2916 (N_2916,N_1870,N_1011);
nor U2917 (N_2917,N_1910,N_1011);
and U2918 (N_2918,N_1410,N_1014);
or U2919 (N_2919,N_1397,N_1570);
nor U2920 (N_2920,N_1994,N_1347);
and U2921 (N_2921,N_1529,N_1930);
xor U2922 (N_2922,N_1884,N_1336);
and U2923 (N_2923,N_1655,N_1316);
or U2924 (N_2924,N_1510,N_1311);
nand U2925 (N_2925,N_1839,N_1950);
nand U2926 (N_2926,N_1265,N_1347);
nand U2927 (N_2927,N_1551,N_1497);
or U2928 (N_2928,N_1540,N_1216);
nor U2929 (N_2929,N_1829,N_1594);
nand U2930 (N_2930,N_1620,N_1696);
or U2931 (N_2931,N_1451,N_1083);
or U2932 (N_2932,N_1634,N_1944);
nor U2933 (N_2933,N_1167,N_1020);
and U2934 (N_2934,N_1619,N_1824);
or U2935 (N_2935,N_1486,N_1683);
nor U2936 (N_2936,N_1964,N_1279);
nor U2937 (N_2937,N_1361,N_1093);
nand U2938 (N_2938,N_1490,N_1619);
and U2939 (N_2939,N_1715,N_1104);
nand U2940 (N_2940,N_1880,N_1096);
nor U2941 (N_2941,N_1468,N_1465);
or U2942 (N_2942,N_1705,N_1952);
or U2943 (N_2943,N_1308,N_1846);
nand U2944 (N_2944,N_1191,N_1338);
and U2945 (N_2945,N_1774,N_1359);
nand U2946 (N_2946,N_1855,N_1277);
nand U2947 (N_2947,N_1455,N_1331);
nor U2948 (N_2948,N_1424,N_1097);
nand U2949 (N_2949,N_1230,N_1411);
nor U2950 (N_2950,N_1859,N_1085);
nand U2951 (N_2951,N_1155,N_1384);
and U2952 (N_2952,N_1748,N_1255);
nand U2953 (N_2953,N_1640,N_1907);
or U2954 (N_2954,N_1310,N_1314);
xor U2955 (N_2955,N_1391,N_1997);
or U2956 (N_2956,N_1548,N_1553);
nand U2957 (N_2957,N_1135,N_1768);
xor U2958 (N_2958,N_1984,N_1722);
nand U2959 (N_2959,N_1808,N_1036);
nand U2960 (N_2960,N_1313,N_1185);
and U2961 (N_2961,N_1731,N_1215);
and U2962 (N_2962,N_1522,N_1246);
nand U2963 (N_2963,N_1834,N_1449);
or U2964 (N_2964,N_1501,N_1255);
and U2965 (N_2965,N_1271,N_1353);
and U2966 (N_2966,N_1688,N_1018);
nor U2967 (N_2967,N_1503,N_1092);
nand U2968 (N_2968,N_1524,N_1113);
or U2969 (N_2969,N_1963,N_1888);
or U2970 (N_2970,N_1291,N_1257);
nor U2971 (N_2971,N_1884,N_1780);
nand U2972 (N_2972,N_1188,N_1893);
nand U2973 (N_2973,N_1688,N_1305);
nand U2974 (N_2974,N_1350,N_1472);
xnor U2975 (N_2975,N_1013,N_1803);
and U2976 (N_2976,N_1454,N_1421);
nor U2977 (N_2977,N_1143,N_1344);
or U2978 (N_2978,N_1545,N_1547);
nor U2979 (N_2979,N_1962,N_1540);
nand U2980 (N_2980,N_1425,N_1965);
and U2981 (N_2981,N_1100,N_1323);
or U2982 (N_2982,N_1788,N_1078);
nor U2983 (N_2983,N_1343,N_1080);
or U2984 (N_2984,N_1654,N_1630);
nor U2985 (N_2985,N_1622,N_1641);
nor U2986 (N_2986,N_1593,N_1363);
nand U2987 (N_2987,N_1376,N_1000);
or U2988 (N_2988,N_1754,N_1976);
nor U2989 (N_2989,N_1585,N_1349);
and U2990 (N_2990,N_1146,N_1966);
nor U2991 (N_2991,N_1336,N_1424);
nor U2992 (N_2992,N_1849,N_1910);
nor U2993 (N_2993,N_1657,N_1986);
nand U2994 (N_2994,N_1647,N_1146);
or U2995 (N_2995,N_1843,N_1176);
and U2996 (N_2996,N_1131,N_1784);
nand U2997 (N_2997,N_1814,N_1299);
and U2998 (N_2998,N_1121,N_1150);
or U2999 (N_2999,N_1191,N_1254);
nor UO_0 (O_0,N_2037,N_2058);
nor UO_1 (O_1,N_2363,N_2730);
and UO_2 (O_2,N_2340,N_2785);
nor UO_3 (O_3,N_2698,N_2974);
nand UO_4 (O_4,N_2255,N_2151);
xnor UO_5 (O_5,N_2269,N_2288);
nor UO_6 (O_6,N_2757,N_2315);
nor UO_7 (O_7,N_2498,N_2737);
nand UO_8 (O_8,N_2817,N_2782);
nor UO_9 (O_9,N_2432,N_2892);
or UO_10 (O_10,N_2844,N_2992);
or UO_11 (O_11,N_2822,N_2849);
nand UO_12 (O_12,N_2179,N_2679);
xnor UO_13 (O_13,N_2706,N_2192);
and UO_14 (O_14,N_2278,N_2745);
xor UO_15 (O_15,N_2949,N_2240);
and UO_16 (O_16,N_2208,N_2409);
nand UO_17 (O_17,N_2019,N_2811);
or UO_18 (O_18,N_2056,N_2504);
nand UO_19 (O_19,N_2143,N_2160);
xor UO_20 (O_20,N_2222,N_2701);
or UO_21 (O_21,N_2842,N_2705);
nand UO_22 (O_22,N_2631,N_2169);
and UO_23 (O_23,N_2751,N_2346);
nor UO_24 (O_24,N_2680,N_2687);
nand UO_25 (O_25,N_2127,N_2589);
and UO_26 (O_26,N_2867,N_2993);
xor UO_27 (O_27,N_2644,N_2625);
or UO_28 (O_28,N_2365,N_2690);
nor UO_29 (O_29,N_2298,N_2436);
or UO_30 (O_30,N_2233,N_2408);
nand UO_31 (O_31,N_2247,N_2952);
nor UO_32 (O_32,N_2057,N_2248);
nor UO_33 (O_33,N_2493,N_2556);
or UO_34 (O_34,N_2976,N_2547);
nor UO_35 (O_35,N_2743,N_2405);
nor UO_36 (O_36,N_2633,N_2656);
nor UO_37 (O_37,N_2792,N_2774);
nor UO_38 (O_38,N_2845,N_2018);
nor UO_39 (O_39,N_2878,N_2416);
xnor UO_40 (O_40,N_2132,N_2317);
and UO_41 (O_41,N_2765,N_2081);
or UO_42 (O_42,N_2520,N_2804);
nor UO_43 (O_43,N_2271,N_2923);
nor UO_44 (O_44,N_2783,N_2552);
xor UO_45 (O_45,N_2188,N_2479);
nor UO_46 (O_46,N_2137,N_2154);
nand UO_47 (O_47,N_2323,N_2083);
or UO_48 (O_48,N_2906,N_2590);
nand UO_49 (O_49,N_2448,N_2726);
nand UO_50 (O_50,N_2866,N_2527);
nor UO_51 (O_51,N_2860,N_2301);
or UO_52 (O_52,N_2749,N_2823);
and UO_53 (O_53,N_2884,N_2766);
xnor UO_54 (O_54,N_2714,N_2183);
or UO_55 (O_55,N_2533,N_2512);
nor UO_56 (O_56,N_2893,N_2003);
or UO_57 (O_57,N_2102,N_2970);
or UO_58 (O_58,N_2606,N_2322);
nor UO_59 (O_59,N_2929,N_2652);
nand UO_60 (O_60,N_2434,N_2847);
nor UO_61 (O_61,N_2353,N_2772);
or UO_62 (O_62,N_2047,N_2013);
nor UO_63 (O_63,N_2702,N_2664);
and UO_64 (O_64,N_2378,N_2030);
nor UO_65 (O_65,N_2209,N_2517);
nor UO_66 (O_66,N_2708,N_2193);
nor UO_67 (O_67,N_2686,N_2624);
or UO_68 (O_68,N_2380,N_2268);
nor UO_69 (O_69,N_2253,N_2387);
and UO_70 (O_70,N_2050,N_2166);
or UO_71 (O_71,N_2114,N_2910);
or UO_72 (O_72,N_2778,N_2854);
nand UO_73 (O_73,N_2264,N_2456);
nor UO_74 (O_74,N_2367,N_2944);
nand UO_75 (O_75,N_2550,N_2775);
nand UO_76 (O_76,N_2939,N_2296);
nor UO_77 (O_77,N_2808,N_2657);
xnor UO_78 (O_78,N_2699,N_2399);
nand UO_79 (O_79,N_2468,N_2519);
xor UO_80 (O_80,N_2382,N_2523);
xnor UO_81 (O_81,N_2753,N_2276);
or UO_82 (O_82,N_2578,N_2295);
or UO_83 (O_83,N_2470,N_2165);
xor UO_84 (O_84,N_2237,N_2877);
xor UO_85 (O_85,N_2306,N_2677);
or UO_86 (O_86,N_2560,N_2833);
nand UO_87 (O_87,N_2999,N_2942);
or UO_88 (O_88,N_2333,N_2835);
or UO_89 (O_89,N_2961,N_2356);
xnor UO_90 (O_90,N_2928,N_2107);
and UO_91 (O_91,N_2258,N_2443);
nor UO_92 (O_92,N_2350,N_2174);
nor UO_93 (O_93,N_2486,N_2173);
xnor UO_94 (O_94,N_2067,N_2226);
nor UO_95 (O_95,N_2465,N_2735);
nor UO_96 (O_96,N_2500,N_2640);
nand UO_97 (O_97,N_2145,N_2245);
nor UO_98 (O_98,N_2598,N_2403);
nand UO_99 (O_99,N_2922,N_2359);
nor UO_100 (O_100,N_2558,N_2885);
and UO_101 (O_101,N_2423,N_2320);
nor UO_102 (O_102,N_2394,N_2022);
nand UO_103 (O_103,N_2364,N_2559);
or UO_104 (O_104,N_2979,N_2988);
and UO_105 (O_105,N_2947,N_2384);
nand UO_106 (O_106,N_2412,N_2039);
or UO_107 (O_107,N_2292,N_2096);
nor UO_108 (O_108,N_2463,N_2046);
or UO_109 (O_109,N_2587,N_2773);
xnor UO_110 (O_110,N_2951,N_2458);
nor UO_111 (O_111,N_2032,N_2871);
nand UO_112 (O_112,N_2548,N_2312);
nand UO_113 (O_113,N_2829,N_2670);
nor UO_114 (O_114,N_2723,N_2986);
xor UO_115 (O_115,N_2703,N_2881);
nor UO_116 (O_116,N_2139,N_2859);
nand UO_117 (O_117,N_2238,N_2246);
and UO_118 (O_118,N_2424,N_2100);
nand UO_119 (O_119,N_2491,N_2781);
nand UO_120 (O_120,N_2768,N_2676);
and UO_121 (O_121,N_2777,N_2709);
nor UO_122 (O_122,N_2564,N_2510);
nand UO_123 (O_123,N_2840,N_2874);
nor UO_124 (O_124,N_2915,N_2930);
nor UO_125 (O_125,N_2116,N_2594);
nand UO_126 (O_126,N_2369,N_2544);
or UO_127 (O_127,N_2397,N_2953);
nor UO_128 (O_128,N_2880,N_2968);
nand UO_129 (O_129,N_2650,N_2526);
or UO_130 (O_130,N_2712,N_2636);
or UO_131 (O_131,N_2170,N_2117);
nor UO_132 (O_132,N_2616,N_2212);
nor UO_133 (O_133,N_2282,N_2430);
or UO_134 (O_134,N_2573,N_2843);
nand UO_135 (O_135,N_2905,N_2812);
nand UO_136 (O_136,N_2718,N_2125);
nor UO_137 (O_137,N_2713,N_2285);
nor UO_138 (O_138,N_2528,N_2095);
nand UO_139 (O_139,N_2622,N_2960);
and UO_140 (O_140,N_2577,N_2603);
and UO_141 (O_141,N_2916,N_2685);
or UO_142 (O_142,N_2637,N_2545);
nand UO_143 (O_143,N_2009,N_2075);
or UO_144 (O_144,N_2795,N_2227);
nand UO_145 (O_145,N_2541,N_2392);
nor UO_146 (O_146,N_2305,N_2641);
nand UO_147 (O_147,N_2293,N_2062);
and UO_148 (O_148,N_2200,N_2146);
and UO_149 (O_149,N_2284,N_2199);
xor UO_150 (O_150,N_2566,N_2888);
or UO_151 (O_151,N_2155,N_2551);
nor UO_152 (O_152,N_2334,N_2002);
and UO_153 (O_153,N_2626,N_2754);
or UO_154 (O_154,N_2784,N_2549);
nor UO_155 (O_155,N_2776,N_2858);
or UO_156 (O_156,N_2756,N_2150);
and UO_157 (O_157,N_2433,N_2761);
xnor UO_158 (O_158,N_2661,N_2567);
nor UO_159 (O_159,N_2920,N_2647);
nor UO_160 (O_160,N_2239,N_2469);
nand UO_161 (O_161,N_2879,N_2389);
xnor UO_162 (O_162,N_2442,N_2126);
and UO_163 (O_163,N_2026,N_2104);
and UO_164 (O_164,N_2600,N_2715);
and UO_165 (O_165,N_2141,N_2210);
or UO_166 (O_166,N_2336,N_2581);
nand UO_167 (O_167,N_2118,N_2411);
and UO_168 (O_168,N_2575,N_2281);
nand UO_169 (O_169,N_2515,N_2375);
nand UO_170 (O_170,N_2655,N_2406);
and UO_171 (O_171,N_2496,N_2739);
and UO_172 (O_172,N_2144,N_2447);
xor UO_173 (O_173,N_2786,N_2249);
nor UO_174 (O_174,N_2287,N_2054);
nand UO_175 (O_175,N_2351,N_2078);
nor UO_176 (O_176,N_2440,N_2001);
or UO_177 (O_177,N_2530,N_2828);
and UO_178 (O_178,N_2900,N_2088);
and UO_179 (O_179,N_2802,N_2068);
and UO_180 (O_180,N_2668,N_2755);
xor UO_181 (O_181,N_2513,N_2629);
or UO_182 (O_182,N_2328,N_2221);
nor UO_183 (O_183,N_2863,N_2591);
and UO_184 (O_184,N_2908,N_2927);
or UO_185 (O_185,N_2172,N_2085);
or UO_186 (O_186,N_2038,N_2005);
nand UO_187 (O_187,N_2439,N_2450);
nand UO_188 (O_188,N_2147,N_2418);
nand UO_189 (O_189,N_2421,N_2462);
nor UO_190 (O_190,N_2327,N_2826);
and UO_191 (O_191,N_2080,N_2499);
nor UO_192 (O_192,N_2279,N_2648);
nand UO_193 (O_193,N_2902,N_2711);
and UO_194 (O_194,N_2402,N_2136);
nand UO_195 (O_195,N_2220,N_2621);
nand UO_196 (O_196,N_2790,N_2228);
nor UO_197 (O_197,N_2224,N_2987);
nor UO_198 (O_198,N_2256,N_2696);
or UO_199 (O_199,N_2407,N_2934);
and UO_200 (O_200,N_2475,N_2780);
and UO_201 (O_201,N_2615,N_2243);
nand UO_202 (O_202,N_2393,N_2204);
xnor UO_203 (O_203,N_2344,N_2063);
nand UO_204 (O_204,N_2277,N_2620);
nand UO_205 (O_205,N_2383,N_2025);
nor UO_206 (O_206,N_2012,N_2597);
and UO_207 (O_207,N_2427,N_2309);
nand UO_208 (O_208,N_2959,N_2638);
or UO_209 (O_209,N_2954,N_2252);
and UO_210 (O_210,N_2020,N_2033);
nor UO_211 (O_211,N_2171,N_2329);
nor UO_212 (O_212,N_2895,N_2330);
nor UO_213 (O_213,N_2876,N_2779);
and UO_214 (O_214,N_2542,N_2265);
or UO_215 (O_215,N_2689,N_2608);
and UO_216 (O_216,N_2918,N_2827);
nor UO_217 (O_217,N_2634,N_2196);
nand UO_218 (O_218,N_2501,N_2163);
nor UO_219 (O_219,N_2031,N_2788);
or UO_220 (O_220,N_2370,N_2110);
or UO_221 (O_221,N_2752,N_2446);
or UO_222 (O_222,N_2793,N_2070);
and UO_223 (O_223,N_2770,N_2958);
nor UO_224 (O_224,N_2618,N_2921);
or UO_225 (O_225,N_2262,N_2474);
xnor UO_226 (O_226,N_2932,N_2267);
or UO_227 (O_227,N_2481,N_2731);
nor UO_228 (O_228,N_2487,N_2694);
and UO_229 (O_229,N_2926,N_2695);
and UO_230 (O_230,N_2189,N_2355);
xor UO_231 (O_231,N_2607,N_2197);
nor UO_232 (O_232,N_2569,N_2283);
nand UO_233 (O_233,N_2997,N_2534);
nand UO_234 (O_234,N_2994,N_2688);
and UO_235 (O_235,N_2563,N_2800);
and UO_236 (O_236,N_2034,N_2747);
nor UO_237 (O_237,N_2352,N_2602);
and UO_238 (O_238,N_2570,N_2077);
and UO_239 (O_239,N_2805,N_2710);
or UO_240 (O_240,N_2175,N_2758);
xor UO_241 (O_241,N_2272,N_2535);
nor UO_242 (O_242,N_2482,N_2152);
nor UO_243 (O_243,N_2574,N_2941);
or UO_244 (O_244,N_2649,N_2707);
nor UO_245 (O_245,N_2816,N_2990);
nand UO_246 (O_246,N_2693,N_2933);
nand UO_247 (O_247,N_2803,N_2917);
or UO_248 (O_248,N_2646,N_2660);
or UO_249 (O_249,N_2787,N_2257);
nor UO_250 (O_250,N_2215,N_2579);
xor UO_251 (O_251,N_2797,N_2121);
or UO_252 (O_252,N_2157,N_2302);
nand UO_253 (O_253,N_2762,N_2123);
nor UO_254 (O_254,N_2108,N_2400);
or UO_255 (O_255,N_2791,N_2203);
or UO_256 (O_256,N_2011,N_2509);
or UO_257 (O_257,N_2027,N_2936);
nor UO_258 (O_258,N_2593,N_2041);
or UO_259 (O_259,N_2891,N_2206);
or UO_260 (O_260,N_2572,N_2744);
nor UO_261 (O_261,N_2870,N_2796);
or UO_262 (O_262,N_2010,N_2925);
and UO_263 (O_263,N_2242,N_2415);
xnor UO_264 (O_264,N_2194,N_2008);
nand UO_265 (O_265,N_2263,N_2483);
nand UO_266 (O_266,N_2073,N_2069);
and UO_267 (O_267,N_2886,N_2798);
or UO_268 (O_268,N_2857,N_2836);
and UO_269 (O_269,N_2911,N_2304);
nand UO_270 (O_270,N_2914,N_2218);
or UO_271 (O_271,N_2072,N_2021);
and UO_272 (O_272,N_2354,N_2824);
nor UO_273 (O_273,N_2120,N_2675);
and UO_274 (O_274,N_2734,N_2217);
nor UO_275 (O_275,N_2310,N_2307);
nor UO_276 (O_276,N_2103,N_2223);
nand UO_277 (O_277,N_2966,N_2251);
nand UO_278 (O_278,N_2361,N_2938);
and UO_279 (O_279,N_2583,N_2623);
and UO_280 (O_280,N_2429,N_2763);
or UO_281 (O_281,N_2972,N_2896);
and UO_282 (O_282,N_2771,N_2091);
or UO_283 (O_283,N_2040,N_2767);
or UO_284 (O_284,N_2543,N_2946);
xor UO_285 (O_285,N_2862,N_2274);
and UO_286 (O_286,N_2971,N_2043);
or UO_287 (O_287,N_2540,N_2848);
or UO_288 (O_288,N_2887,N_2588);
nand UO_289 (O_289,N_2945,N_2425);
or UO_290 (O_290,N_2130,N_2273);
nand UO_291 (O_291,N_2162,N_2901);
nand UO_292 (O_292,N_2834,N_2082);
or UO_293 (O_293,N_2511,N_2627);
or UO_294 (O_294,N_2831,N_2931);
and UO_295 (O_295,N_2229,N_2505);
nand UO_296 (O_296,N_2349,N_2724);
nor UO_297 (O_297,N_2684,N_2422);
nor UO_298 (O_298,N_2148,N_2149);
and UO_299 (O_299,N_2266,N_2131);
or UO_300 (O_300,N_2357,N_2366);
nand UO_301 (O_301,N_2538,N_2135);
nor UO_302 (O_302,N_2903,N_2856);
nor UO_303 (O_303,N_2662,N_2219);
and UO_304 (O_304,N_2935,N_2207);
nand UO_305 (O_305,N_2729,N_2736);
nor UO_306 (O_306,N_2890,N_2467);
and UO_307 (O_307,N_2586,N_2459);
and UO_308 (O_308,N_2555,N_2546);
nand UO_309 (O_309,N_2000,N_2524);
nand UO_310 (O_310,N_2964,N_2230);
xnor UO_311 (O_311,N_2948,N_2168);
and UO_312 (O_312,N_2825,N_2478);
nand UO_313 (O_313,N_2654,N_2176);
and UO_314 (O_314,N_2379,N_2813);
nor UO_315 (O_315,N_2818,N_2435);
nor UO_316 (O_316,N_2899,N_2099);
xor UO_317 (O_317,N_2728,N_2051);
xor UO_318 (O_318,N_2029,N_2195);
nand UO_319 (O_319,N_2760,N_2841);
nand UO_320 (O_320,N_2466,N_2553);
and UO_321 (O_321,N_2477,N_2973);
and UO_322 (O_322,N_2216,N_2580);
nand UO_323 (O_323,N_2348,N_2372);
and UO_324 (O_324,N_2605,N_2024);
and UO_325 (O_325,N_2963,N_2213);
nor UO_326 (O_326,N_2984,N_2205);
xor UO_327 (O_327,N_2975,N_2830);
nor UO_328 (O_328,N_2846,N_2358);
nor UO_329 (O_329,N_2497,N_2140);
or UO_330 (O_330,N_2628,N_2316);
or UO_331 (O_331,N_2645,N_2294);
and UO_332 (O_332,N_2225,N_2855);
nor UO_333 (O_333,N_2610,N_2683);
or UO_334 (O_334,N_2318,N_2653);
nand UO_335 (O_335,N_2419,N_2396);
nor UO_336 (O_336,N_2506,N_2557);
nand UO_337 (O_337,N_2414,N_2385);
xnor UO_338 (O_338,N_2275,N_2955);
nand UO_339 (O_339,N_2764,N_2682);
or UO_340 (O_340,N_2592,N_2814);
nand UO_341 (O_341,N_2201,N_2977);
and UO_342 (O_342,N_2035,N_2472);
or UO_343 (O_343,N_2630,N_2967);
or UO_344 (O_344,N_2565,N_2250);
and UO_345 (O_345,N_2464,N_2721);
and UO_346 (O_346,N_2438,N_2617);
and UO_347 (O_347,N_2673,N_2321);
nand UO_348 (O_348,N_2554,N_2122);
nand UO_349 (O_349,N_2052,N_2738);
nor UO_350 (O_350,N_2453,N_2769);
and UO_351 (O_351,N_2522,N_2270);
and UO_352 (O_352,N_2733,N_2852);
or UO_353 (O_353,N_2036,N_2853);
or UO_354 (O_354,N_2332,N_2291);
xnor UO_355 (O_355,N_2619,N_2090);
and UO_356 (O_356,N_2894,N_2084);
and UO_357 (O_357,N_2381,N_2585);
nor UO_358 (O_358,N_2410,N_2989);
or UO_359 (O_359,N_2182,N_2665);
or UO_360 (O_360,N_2998,N_2700);
nand UO_361 (O_361,N_2325,N_2865);
or UO_362 (O_362,N_2324,N_2850);
and UO_363 (O_363,N_2105,N_2134);
nor UO_364 (O_364,N_2339,N_2167);
or UO_365 (O_365,N_2601,N_2595);
or UO_366 (O_366,N_2985,N_2234);
and UO_367 (O_367,N_2319,N_2672);
xnor UO_368 (O_368,N_2821,N_2996);
nor UO_369 (O_369,N_2187,N_2875);
and UO_370 (O_370,N_2004,N_2488);
nor UO_371 (O_371,N_2044,N_2741);
nor UO_372 (O_372,N_2014,N_2232);
nand UO_373 (O_373,N_2064,N_2957);
and UO_374 (O_374,N_2161,N_2667);
nor UO_375 (O_375,N_2658,N_2609);
xnor UO_376 (O_376,N_2789,N_2704);
nor UO_377 (O_377,N_2980,N_2065);
nand UO_378 (O_378,N_2473,N_2299);
nor UO_379 (O_379,N_2343,N_2180);
nand UO_380 (O_380,N_2087,N_2806);
nor UO_381 (O_381,N_2460,N_2981);
or UO_382 (O_382,N_2485,N_2398);
xor UO_383 (O_383,N_2851,N_2300);
or UO_384 (O_384,N_2308,N_2074);
and UO_385 (O_385,N_2211,N_2360);
and UO_386 (O_386,N_2426,N_2461);
or UO_387 (O_387,N_2940,N_2373);
and UO_388 (O_388,N_2576,N_2452);
and UO_389 (O_389,N_2897,N_2518);
nor UO_390 (O_390,N_2801,N_2663);
nand UO_391 (O_391,N_2489,N_2156);
and UO_392 (O_392,N_2347,N_2995);
nand UO_393 (O_393,N_2457,N_2331);
nor UO_394 (O_394,N_2431,N_2015);
nor UO_395 (O_395,N_2883,N_2508);
xor UO_396 (O_396,N_2244,N_2691);
or UO_397 (O_397,N_2338,N_2437);
and UO_398 (O_398,N_2674,N_2260);
and UO_399 (O_399,N_2254,N_2725);
nor UO_400 (O_400,N_2599,N_2314);
nor UO_401 (O_401,N_2061,N_2017);
and UO_402 (O_402,N_2839,N_2097);
or UO_403 (O_403,N_2420,N_2133);
xor UO_404 (O_404,N_2525,N_2186);
nor UO_405 (O_405,N_2094,N_2692);
nor UO_406 (O_406,N_2869,N_2503);
xnor UO_407 (O_407,N_2809,N_2112);
nor UO_408 (O_408,N_2115,N_2060);
or UO_409 (O_409,N_2185,N_2717);
or UO_410 (O_410,N_2106,N_2864);
nand UO_411 (O_411,N_2531,N_2391);
nand UO_412 (O_412,N_2666,N_2076);
nor UO_413 (O_413,N_2376,N_2449);
and UO_414 (O_414,N_2476,N_2861);
nor UO_415 (O_415,N_2490,N_2289);
nand UO_416 (O_416,N_2016,N_2158);
and UO_417 (O_417,N_2297,N_2943);
xnor UO_418 (O_418,N_2311,N_2720);
nand UO_419 (O_419,N_2362,N_2502);
nand UO_420 (O_420,N_2374,N_2950);
and UO_421 (O_421,N_2124,N_2342);
nand UO_422 (O_422,N_2820,N_2898);
nand UO_423 (O_423,N_2214,N_2101);
or UO_424 (O_424,N_2907,N_2872);
or UO_425 (O_425,N_2536,N_2562);
nand UO_426 (O_426,N_2740,N_2532);
nand UO_427 (O_427,N_2919,N_2584);
and UO_428 (O_428,N_2582,N_2390);
nand UO_429 (O_429,N_2441,N_2386);
or UO_430 (O_430,N_2401,N_2092);
and UO_431 (O_431,N_2604,N_2129);
nand UO_432 (O_432,N_2962,N_2678);
and UO_433 (O_433,N_2495,N_2303);
or UO_434 (O_434,N_2742,N_2815);
xnor UO_435 (O_435,N_2727,N_2671);
and UO_436 (O_436,N_2937,N_2259);
and UO_437 (O_437,N_2086,N_2261);
or UO_438 (O_438,N_2492,N_2965);
or UO_439 (O_439,N_2049,N_2111);
nand UO_440 (O_440,N_2810,N_2444);
xor UO_441 (O_441,N_2113,N_2159);
and UO_442 (O_442,N_2882,N_2480);
or UO_443 (O_443,N_2611,N_2837);
and UO_444 (O_444,N_2669,N_2007);
nand UO_445 (O_445,N_2202,N_2507);
nand UO_446 (O_446,N_2571,N_2153);
xor UO_447 (O_447,N_2494,N_2529);
or UO_448 (O_448,N_2138,N_2516);
nor UO_449 (O_449,N_2969,N_2345);
nor UO_450 (O_450,N_2006,N_2241);
nand UO_451 (O_451,N_2983,N_2313);
nor UO_452 (O_452,N_2904,N_2807);
and UO_453 (O_453,N_2639,N_2794);
nand UO_454 (O_454,N_2341,N_2514);
nor UO_455 (O_455,N_2748,N_2190);
nand UO_456 (O_456,N_2978,N_2371);
or UO_457 (O_457,N_2991,N_2388);
or UO_458 (O_458,N_2280,N_2286);
or UO_459 (O_459,N_2613,N_2198);
xnor UO_460 (O_460,N_2614,N_2873);
or UO_461 (O_461,N_2290,N_2750);
or UO_462 (O_462,N_2612,N_2484);
xor UO_463 (O_463,N_2404,N_2181);
nor UO_464 (O_464,N_2819,N_2023);
xor UO_465 (O_465,N_2417,N_2048);
or UO_466 (O_466,N_2028,N_2335);
or UO_467 (O_467,N_2838,N_2089);
or UO_468 (O_468,N_2568,N_2521);
and UO_469 (O_469,N_2643,N_2428);
xor UO_470 (O_470,N_2632,N_2451);
nor UO_471 (O_471,N_2178,N_2746);
nand UO_472 (O_472,N_2681,N_2596);
or UO_473 (O_473,N_2079,N_2889);
nor UO_474 (O_474,N_2722,N_2445);
nor UO_475 (O_475,N_2326,N_2093);
nor UO_476 (O_476,N_2719,N_2912);
or UO_477 (O_477,N_2042,N_2537);
nand UO_478 (O_478,N_2799,N_2868);
nor UO_479 (O_479,N_2832,N_2177);
xor UO_480 (O_480,N_2128,N_2455);
nand UO_481 (O_481,N_2337,N_2732);
and UO_482 (O_482,N_2236,N_2913);
or UO_483 (O_483,N_2066,N_2053);
or UO_484 (O_484,N_2659,N_2697);
nand UO_485 (O_485,N_2164,N_2454);
and UO_486 (O_486,N_2651,N_2231);
and UO_487 (O_487,N_2716,N_2413);
xor UO_488 (O_488,N_2184,N_2119);
and UO_489 (O_489,N_2561,N_2759);
nor UO_490 (O_490,N_2982,N_2642);
nor UO_491 (O_491,N_2368,N_2924);
nor UO_492 (O_492,N_2235,N_2142);
and UO_493 (O_493,N_2909,N_2635);
nand UO_494 (O_494,N_2191,N_2059);
and UO_495 (O_495,N_2956,N_2071);
or UO_496 (O_496,N_2471,N_2098);
or UO_497 (O_497,N_2109,N_2045);
and UO_498 (O_498,N_2395,N_2055);
nand UO_499 (O_499,N_2377,N_2539);
endmodule