module basic_3000_30000_3500_60_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_2695,In_2009);
nand U1 (N_1,In_1356,In_2639);
xnor U2 (N_2,In_1079,In_2296);
or U3 (N_3,In_550,In_1757);
xnor U4 (N_4,In_1670,In_2713);
nand U5 (N_5,In_2268,In_2400);
nor U6 (N_6,In_468,In_2339);
or U7 (N_7,In_2261,In_938);
and U8 (N_8,In_1298,In_24);
xor U9 (N_9,In_1693,In_290);
nand U10 (N_10,In_1797,In_504);
nor U11 (N_11,In_1453,In_2195);
nor U12 (N_12,In_2859,In_1138);
and U13 (N_13,In_2371,In_2314);
nor U14 (N_14,In_987,In_216);
xor U15 (N_15,In_1989,In_723);
and U16 (N_16,In_582,In_1069);
nand U17 (N_17,In_1399,In_789);
and U18 (N_18,In_2176,In_1664);
nor U19 (N_19,In_263,In_480);
xnor U20 (N_20,In_678,In_2146);
or U21 (N_21,In_28,In_2003);
or U22 (N_22,In_1835,In_1321);
nand U23 (N_23,In_2379,In_718);
and U24 (N_24,In_351,In_434);
xnor U25 (N_25,In_1563,In_1443);
nand U26 (N_26,In_2868,In_1653);
xor U27 (N_27,In_386,In_81);
nor U28 (N_28,In_1917,In_1235);
nand U29 (N_29,In_2599,In_2735);
nor U30 (N_30,In_834,In_537);
and U31 (N_31,In_2601,In_1018);
or U32 (N_32,In_2205,In_486);
nand U33 (N_33,In_2538,In_1461);
xor U34 (N_34,In_1267,In_2478);
nor U35 (N_35,In_1983,In_2585);
nor U36 (N_36,In_2680,In_2206);
and U37 (N_37,In_883,In_383);
xnor U38 (N_38,In_2793,In_757);
and U39 (N_39,In_17,In_1587);
or U40 (N_40,In_1287,In_59);
nand U41 (N_41,In_679,In_2962);
xnor U42 (N_42,In_1987,In_2246);
nand U43 (N_43,In_1828,In_1569);
or U44 (N_44,In_1866,In_2736);
or U45 (N_45,In_2306,In_1154);
xor U46 (N_46,In_1995,In_1977);
or U47 (N_47,In_606,In_2771);
and U48 (N_48,In_1632,In_1842);
and U49 (N_49,In_2663,In_868);
and U50 (N_50,In_1804,In_41);
and U51 (N_51,In_147,In_127);
nand U52 (N_52,In_684,In_701);
nor U53 (N_53,In_1278,In_2345);
xnor U54 (N_54,In_1617,In_770);
nor U55 (N_55,In_1323,In_1491);
nand U56 (N_56,In_2225,In_620);
nand U57 (N_57,In_1483,In_82);
nor U58 (N_58,In_592,In_19);
nand U59 (N_59,In_2567,In_2689);
xor U60 (N_60,In_2203,In_322);
and U61 (N_61,In_1722,In_2481);
nor U62 (N_62,In_247,In_695);
nor U63 (N_63,In_2323,In_2968);
xnor U64 (N_64,In_96,In_1347);
or U65 (N_65,In_2471,In_612);
nor U66 (N_66,In_1131,In_523);
xnor U67 (N_67,In_2377,In_258);
or U68 (N_68,In_2604,In_274);
xor U69 (N_69,In_1663,In_162);
nor U70 (N_70,In_87,In_2760);
nand U71 (N_71,In_1428,In_1480);
xor U72 (N_72,In_2961,In_926);
nand U73 (N_73,In_907,In_1176);
or U74 (N_74,In_1197,In_1004);
nand U75 (N_75,In_1326,In_2986);
nor U76 (N_76,In_433,In_1529);
and U77 (N_77,In_208,In_2340);
nand U78 (N_78,In_2113,In_2864);
or U79 (N_79,In_281,In_2441);
nor U80 (N_80,In_1495,In_2816);
xnor U81 (N_81,In_1605,In_930);
xnor U82 (N_82,In_385,In_2943);
nand U83 (N_83,In_1971,In_1800);
nand U84 (N_84,In_409,In_2580);
xor U85 (N_85,In_2947,In_1586);
or U86 (N_86,In_2437,In_2933);
nor U87 (N_87,In_2174,In_1059);
nand U88 (N_88,In_458,In_1208);
nand U89 (N_89,In_739,In_1183);
xor U90 (N_90,In_1423,In_1731);
nand U91 (N_91,In_2243,In_2730);
xor U92 (N_92,In_865,In_863);
nand U93 (N_93,In_1787,In_981);
nand U94 (N_94,In_2895,In_1871);
and U95 (N_95,In_974,In_1340);
xor U96 (N_96,In_2955,In_2182);
and U97 (N_97,In_2396,In_697);
nand U98 (N_98,In_2088,In_390);
and U99 (N_99,In_271,In_2332);
or U100 (N_100,In_1872,In_1430);
and U101 (N_101,In_347,In_558);
or U102 (N_102,In_2742,In_2387);
xor U103 (N_103,In_122,In_1745);
xor U104 (N_104,In_2051,In_2410);
nand U105 (N_105,In_1532,In_2833);
and U106 (N_106,In_310,In_158);
and U107 (N_107,In_647,In_1300);
or U108 (N_108,In_867,In_806);
nor U109 (N_109,In_1614,In_2671);
nor U110 (N_110,In_967,In_1230);
and U111 (N_111,In_652,In_839);
xor U112 (N_112,In_878,In_1503);
or U113 (N_113,In_847,In_163);
nor U114 (N_114,In_2924,In_2327);
nand U115 (N_115,In_2389,In_604);
nor U116 (N_116,In_1322,In_677);
or U117 (N_117,In_1581,In_476);
xnor U118 (N_118,In_1623,In_174);
xor U119 (N_119,In_1882,In_2238);
nand U120 (N_120,In_2079,In_2395);
xnor U121 (N_121,In_1224,In_2825);
nor U122 (N_122,In_2098,In_2964);
xor U123 (N_123,In_1202,In_411);
nand U124 (N_124,In_1695,In_342);
and U125 (N_125,In_2770,In_786);
nand U126 (N_126,In_1736,In_2775);
nor U127 (N_127,In_154,In_1525);
nand U128 (N_128,In_1796,In_2245);
nor U129 (N_129,In_2015,In_521);
and U130 (N_130,In_1771,In_2140);
nand U131 (N_131,In_694,In_226);
nor U132 (N_132,In_464,In_1206);
nand U133 (N_133,In_928,In_105);
xor U134 (N_134,In_1972,In_1849);
xor U135 (N_135,In_2401,In_1201);
nand U136 (N_136,In_1658,In_2131);
xor U137 (N_137,In_1134,In_2880);
xor U138 (N_138,In_1629,In_2175);
and U139 (N_139,In_1130,In_1920);
xor U140 (N_140,In_763,In_833);
nand U141 (N_141,In_2152,In_2761);
xnor U142 (N_142,In_1256,In_1816);
and U143 (N_143,In_2013,In_736);
and U144 (N_144,In_4,In_250);
and U145 (N_145,In_2486,In_2526);
and U146 (N_146,In_83,In_2788);
nand U147 (N_147,In_1243,In_1213);
and U148 (N_148,In_1959,In_782);
nor U149 (N_149,In_1967,In_401);
nand U150 (N_150,In_1051,In_2520);
or U151 (N_151,In_966,In_1098);
or U152 (N_152,In_1783,In_2561);
and U153 (N_153,In_1738,In_1549);
xor U154 (N_154,In_1395,In_2315);
nor U155 (N_155,In_2551,In_905);
or U156 (N_156,In_1724,In_1506);
xor U157 (N_157,In_2091,In_1158);
and U158 (N_158,In_1892,In_490);
nand U159 (N_159,In_309,In_68);
and U160 (N_160,In_2221,In_1493);
and U161 (N_161,In_2840,In_578);
and U162 (N_162,In_1937,In_818);
nor U163 (N_163,In_929,In_373);
xnor U164 (N_164,In_2207,In_1472);
xor U165 (N_165,In_1818,In_1439);
nor U166 (N_166,In_1455,In_2021);
nand U167 (N_167,In_2727,In_1332);
and U168 (N_168,In_1271,In_2944);
or U169 (N_169,In_2575,In_725);
nor U170 (N_170,In_2738,In_1950);
and U171 (N_171,In_1388,In_2800);
nor U172 (N_172,In_222,In_2495);
xnor U173 (N_173,In_1275,In_614);
and U174 (N_174,In_79,In_513);
and U175 (N_175,In_2677,In_826);
or U176 (N_176,In_690,In_2064);
and U177 (N_177,In_2367,In_1434);
and U178 (N_178,In_2080,In_1427);
nor U179 (N_179,In_2594,In_1218);
nor U180 (N_180,In_10,In_1358);
nor U181 (N_181,In_2328,In_2666);
or U182 (N_182,In_666,In_2209);
xnor U183 (N_183,In_2465,In_1705);
xor U184 (N_184,In_1638,In_1446);
and U185 (N_185,In_256,In_2706);
nand U186 (N_186,In_175,In_2417);
and U187 (N_187,In_1307,In_783);
and U188 (N_188,In_970,In_2863);
nor U189 (N_189,In_1492,In_221);
xnor U190 (N_190,In_1346,In_2286);
xor U191 (N_191,In_549,In_1755);
nor U192 (N_192,In_2460,In_1073);
xor U193 (N_193,In_1891,In_1254);
and U194 (N_194,In_2996,In_1553);
nor U195 (N_195,In_1246,In_2353);
nand U196 (N_196,In_224,In_740);
nor U197 (N_197,In_1277,In_156);
and U198 (N_198,In_2081,In_1511);
nor U199 (N_199,In_692,In_772);
or U200 (N_200,In_2258,In_484);
nand U201 (N_201,In_1807,In_165);
nor U202 (N_202,In_2305,In_1058);
or U203 (N_203,In_1055,In_2819);
xnor U204 (N_204,In_400,In_2688);
xnor U205 (N_205,In_884,In_1220);
or U206 (N_206,In_2330,In_2732);
and U207 (N_207,In_2240,In_1716);
nor U208 (N_208,In_1824,In_1168);
xor U209 (N_209,In_1257,In_2914);
or U210 (N_210,In_2177,In_1460);
nand U211 (N_211,In_916,In_2568);
xor U212 (N_212,In_1464,In_2300);
xnor U213 (N_213,In_1020,In_532);
xor U214 (N_214,In_2159,In_1970);
xor U215 (N_215,In_2000,In_1885);
nand U216 (N_216,In_2194,In_315);
or U217 (N_217,In_2952,In_1316);
and U218 (N_218,In_328,In_2782);
nor U219 (N_219,In_1504,In_1597);
and U220 (N_220,In_803,In_2154);
nor U221 (N_221,In_910,In_1861);
or U222 (N_222,In_2014,In_730);
nand U223 (N_223,In_2930,In_1540);
nor U224 (N_224,In_2352,In_533);
or U225 (N_225,In_1462,In_76);
nand U226 (N_226,In_827,In_1710);
and U227 (N_227,In_648,In_2762);
nor U228 (N_228,In_2333,In_2096);
xnor U229 (N_229,In_1732,In_84);
and U230 (N_230,In_1893,In_660);
nand U231 (N_231,In_2848,In_2757);
or U232 (N_232,In_116,In_2813);
and U233 (N_233,In_1589,In_2709);
nand U234 (N_234,In_1301,In_1555);
and U235 (N_235,In_2070,In_1988);
xnor U236 (N_236,In_1012,In_2433);
nor U237 (N_237,In_185,In_2126);
nand U238 (N_238,In_1524,In_325);
nor U239 (N_239,In_1507,In_623);
and U240 (N_240,In_619,In_721);
or U241 (N_241,In_542,In_1645);
xnor U242 (N_242,In_564,In_960);
nor U243 (N_243,In_955,In_1204);
nor U244 (N_244,In_851,In_1258);
nor U245 (N_245,In_2334,In_2347);
or U246 (N_246,In_745,In_610);
nand U247 (N_247,In_1252,In_2259);
nor U248 (N_248,In_498,In_2712);
or U249 (N_249,In_1185,In_1558);
xor U250 (N_250,In_2073,In_2045);
nand U251 (N_251,In_2809,In_2617);
xor U252 (N_252,In_983,In_1536);
nand U253 (N_253,In_934,In_790);
nand U254 (N_254,In_2879,In_2630);
nor U255 (N_255,In_191,In_545);
and U256 (N_256,In_1854,In_2262);
nand U257 (N_257,In_625,In_1496);
nand U258 (N_258,In_913,In_1801);
or U259 (N_259,In_2659,In_1000);
and U260 (N_260,In_190,In_1895);
xor U261 (N_261,In_2815,In_2100);
xor U262 (N_262,In_2001,In_1105);
nor U263 (N_263,In_540,In_2278);
or U264 (N_264,In_1010,In_2111);
nor U265 (N_265,In_875,In_2385);
nor U266 (N_266,In_1593,In_2446);
xnor U267 (N_267,In_1016,In_2997);
nand U268 (N_268,In_1671,In_1123);
xor U269 (N_269,In_2728,In_2116);
nor U270 (N_270,In_2544,In_166);
nor U271 (N_271,In_2110,In_2167);
or U272 (N_272,In_1484,In_2479);
and U273 (N_273,In_2628,In_2239);
xor U274 (N_274,In_1171,In_2560);
nor U275 (N_275,In_1320,In_2720);
or U276 (N_276,In_1062,In_534);
xnor U277 (N_277,In_2973,In_2162);
nand U278 (N_278,In_220,In_1898);
xnor U279 (N_279,In_88,In_682);
or U280 (N_280,In_2076,In_706);
nand U281 (N_281,In_1160,In_1808);
xor U282 (N_282,In_2291,In_817);
nand U283 (N_283,In_2425,In_1683);
nor U284 (N_284,In_1251,In_1559);
xnor U285 (N_285,In_601,In_2002);
and U286 (N_286,In_879,In_2418);
xnor U287 (N_287,In_2703,In_337);
nand U288 (N_288,In_2292,In_104);
nor U289 (N_289,In_2573,In_2574);
nor U290 (N_290,In_16,In_2890);
nand U291 (N_291,In_2234,In_1070);
nor U292 (N_292,In_2108,In_2115);
nand U293 (N_293,In_108,In_2447);
nand U294 (N_294,In_1420,In_103);
or U295 (N_295,In_118,In_1215);
xnor U296 (N_296,In_712,In_140);
xnor U297 (N_297,In_1229,In_2360);
xnor U298 (N_298,In_2208,In_959);
and U299 (N_299,In_2834,In_1588);
nand U300 (N_300,In_1268,In_1477);
xor U301 (N_301,In_2769,In_781);
nand U302 (N_302,In_29,In_1474);
xnor U303 (N_303,In_2250,In_1369);
xor U304 (N_304,In_1102,In_734);
xor U305 (N_305,In_1889,In_1718);
and U306 (N_306,In_810,In_1402);
xor U307 (N_307,In_182,In_278);
or U308 (N_308,In_2531,In_2063);
nand U309 (N_309,In_1636,In_144);
xor U310 (N_310,In_121,In_828);
xnor U311 (N_311,In_435,In_2452);
xnor U312 (N_312,In_526,In_2725);
nor U313 (N_313,In_304,In_2321);
xnor U314 (N_314,In_668,In_2189);
nand U315 (N_315,In_1390,In_2104);
xor U316 (N_316,In_636,In_1720);
nand U317 (N_317,In_871,In_2496);
nand U318 (N_318,In_2295,In_985);
nand U319 (N_319,In_2500,In_1936);
nor U320 (N_320,In_769,In_2589);
nand U321 (N_321,In_2831,In_727);
or U322 (N_322,In_98,In_1437);
nor U323 (N_323,In_2411,In_285);
nor U324 (N_324,In_2435,In_1851);
nor U325 (N_325,In_2931,In_2247);
nand U326 (N_326,In_143,In_516);
and U327 (N_327,In_2925,In_206);
or U328 (N_328,In_371,In_482);
and U329 (N_329,In_2990,In_686);
and U330 (N_330,In_756,In_308);
and U331 (N_331,In_937,In_2469);
or U332 (N_332,In_2336,In_671);
xnor U333 (N_333,In_170,In_2785);
xnor U334 (N_334,In_8,In_1573);
nor U335 (N_335,In_1749,In_2641);
or U336 (N_336,In_1371,In_1782);
nor U337 (N_337,In_123,In_2607);
or U338 (N_338,In_345,In_201);
nand U339 (N_339,In_2753,In_135);
nand U340 (N_340,In_2402,In_2739);
xnor U341 (N_341,In_2514,In_1644);
nand U342 (N_342,In_2138,In_747);
nand U343 (N_343,In_2075,In_1233);
and U344 (N_344,In_2214,In_1036);
or U345 (N_345,In_815,In_1698);
or U346 (N_346,In_1719,In_563);
or U347 (N_347,In_119,In_2503);
or U348 (N_348,In_2335,In_1863);
xor U349 (N_349,In_2875,In_2512);
nor U350 (N_350,In_2287,In_1568);
and U351 (N_351,In_2878,In_1711);
or U352 (N_352,In_2984,In_2598);
nand U353 (N_353,In_2505,In_901);
xor U354 (N_354,In_1177,In_60);
and U355 (N_355,In_2749,In_2854);
nand U356 (N_356,In_407,In_387);
nand U357 (N_357,In_2413,In_244);
and U358 (N_358,In_716,In_761);
nor U359 (N_359,In_1875,In_915);
xnor U360 (N_360,In_531,In_1781);
xnor U361 (N_361,In_12,In_811);
and U362 (N_362,In_1289,In_1485);
and U363 (N_363,In_1654,In_2645);
and U364 (N_364,In_573,In_1337);
and U365 (N_365,In_1031,In_167);
xnor U366 (N_366,In_1403,In_909);
nor U367 (N_367,In_1806,In_1038);
and U368 (N_368,In_750,In_2649);
or U369 (N_369,In_635,In_798);
or U370 (N_370,In_2027,In_2988);
nand U371 (N_371,In_357,In_71);
nand U372 (N_372,In_1092,In_1838);
and U373 (N_373,In_752,In_2983);
nor U374 (N_374,In_1922,In_2398);
or U375 (N_375,In_621,In_350);
xor U376 (N_376,In_1409,In_2765);
or U377 (N_377,In_2581,In_297);
nor U378 (N_378,In_2343,In_1157);
nor U379 (N_379,In_1648,In_593);
xnor U380 (N_380,In_2294,In_1148);
xor U381 (N_381,In_1659,In_217);
xor U382 (N_382,In_683,In_2290);
nand U383 (N_383,In_2661,In_141);
nand U384 (N_384,In_1565,In_1375);
xnor U385 (N_385,In_2766,In_2178);
nor U386 (N_386,In_1743,In_2613);
or U387 (N_387,In_1169,In_1030);
and U388 (N_388,In_804,In_1034);
nor U389 (N_389,In_2654,In_1510);
nand U390 (N_390,In_599,In_1577);
and U391 (N_391,In_456,In_1772);
nor U392 (N_392,In_1774,In_1852);
and U393 (N_393,In_2242,In_355);
and U394 (N_394,In_572,In_445);
or U395 (N_395,In_574,In_1378);
or U396 (N_396,In_829,In_774);
nand U397 (N_397,In_1343,In_749);
nand U398 (N_398,In_1063,In_2307);
and U399 (N_399,In_2887,In_1471);
and U400 (N_400,In_1998,In_979);
xor U401 (N_401,In_819,In_988);
nand U402 (N_402,In_1047,In_2230);
and U403 (N_403,In_1406,In_1272);
xor U404 (N_404,In_515,In_1883);
nor U405 (N_405,In_0,In_748);
nor U406 (N_406,In_1119,In_1840);
nand U407 (N_407,In_1211,In_53);
and U408 (N_408,In_1578,In_655);
xor U409 (N_409,In_2744,In_313);
and U410 (N_410,In_2533,In_1915);
xnor U411 (N_411,In_1142,In_2297);
nor U412 (N_412,In_2142,In_2827);
nor U413 (N_413,In_957,In_672);
nor U414 (N_414,In_1468,In_2556);
or U415 (N_415,In_1100,In_2523);
or U416 (N_416,In_2846,In_2674);
or U417 (N_417,In_2464,In_2180);
or U418 (N_418,In_1523,In_948);
nor U419 (N_419,In_579,In_2615);
xnor U420 (N_420,In_1265,In_2032);
nand U421 (N_421,In_1684,In_496);
nor U422 (N_422,In_2789,In_2605);
or U423 (N_423,In_787,In_2625);
or U424 (N_424,In_2274,In_1489);
nand U425 (N_425,In_510,In_2950);
xor U426 (N_426,In_440,In_1310);
or U427 (N_427,In_366,In_2404);
or U428 (N_428,In_396,In_773);
or U429 (N_429,In_2578,In_2651);
nand U430 (N_430,In_2927,In_437);
and U431 (N_431,In_1207,In_1742);
nand U432 (N_432,In_1527,In_935);
or U433 (N_433,In_1377,In_2976);
nand U434 (N_434,In_319,In_1222);
xor U435 (N_435,In_238,In_963);
nor U436 (N_436,In_715,In_1652);
xnor U437 (N_437,In_661,In_2097);
nor U438 (N_438,In_576,In_494);
xor U439 (N_439,In_2191,In_571);
and U440 (N_440,In_2623,In_2093);
nand U441 (N_441,In_662,In_146);
xor U442 (N_442,In_577,In_1539);
or U443 (N_443,In_1159,In_600);
and U444 (N_444,In_997,In_2281);
nand U445 (N_445,In_908,In_2629);
nor U446 (N_446,In_596,In_2037);
nand U447 (N_447,In_2382,In_972);
xor U448 (N_448,In_1276,In_2302);
and U449 (N_449,In_2949,In_1141);
and U450 (N_450,In_2745,In_1096);
nand U451 (N_451,In_2778,In_1822);
and U452 (N_452,In_699,In_1433);
and U453 (N_453,In_1,In_1245);
nand U454 (N_454,In_2384,In_824);
nand U455 (N_455,In_2546,In_1554);
nor U456 (N_456,In_1848,In_2839);
nand U457 (N_457,In_2129,In_1596);
xor U458 (N_458,In_101,In_1675);
nor U459 (N_459,In_203,In_1649);
nor U460 (N_460,In_1550,In_2527);
nand U461 (N_461,In_764,In_2786);
or U462 (N_462,In_2378,In_2752);
nor U463 (N_463,In_1083,In_1608);
nor U464 (N_464,In_180,In_1234);
xor U465 (N_465,In_2822,In_2254);
and U466 (N_466,In_1054,In_1019);
or U467 (N_467,In_1458,In_673);
and U468 (N_468,In_1494,In_26);
and U469 (N_469,In_1613,In_999);
nand U470 (N_470,In_950,In_1717);
or U471 (N_471,In_547,In_1957);
and U472 (N_472,In_1951,In_1162);
nor U473 (N_473,In_268,In_861);
or U474 (N_474,In_1135,In_1619);
nand U475 (N_475,In_2965,In_733);
and U476 (N_476,In_990,In_2493);
or U477 (N_477,In_2515,In_1469);
or U478 (N_478,In_1580,In_2529);
and U479 (N_479,In_1582,In_561);
and U480 (N_480,In_2151,In_200);
xor U481 (N_481,In_86,In_1997);
and U482 (N_482,In_502,In_1499);
and U483 (N_483,In_20,In_1344);
nor U484 (N_484,In_1958,In_941);
nor U485 (N_485,In_2006,In_1583);
xor U486 (N_486,In_2856,In_231);
xor U487 (N_487,In_99,In_1992);
nand U488 (N_488,In_368,In_2781);
nor U489 (N_489,In_1380,In_1389);
nand U490 (N_490,In_1572,In_2423);
nand U491 (N_491,In_1890,In_2843);
or U492 (N_492,In_1793,In_2213);
xnor U493 (N_493,In_265,In_1186);
and U494 (N_494,In_989,In_500);
and U495 (N_495,In_2066,In_1441);
or U496 (N_496,In_1255,In_299);
nand U497 (N_497,In_1934,In_22);
and U498 (N_498,In_1811,In_1026);
nor U499 (N_499,In_2042,In_1981);
or U500 (N_500,In_428,In_2821);
xor U501 (N_501,In_425,In_1081);
nor U502 (N_502,In_626,In_2889);
and U503 (N_503,In_2101,N_98);
nand U504 (N_504,In_1355,In_2403);
and U505 (N_505,N_484,In_1545);
and U506 (N_506,N_426,In_583);
nand U507 (N_507,In_2361,In_1006);
nor U508 (N_508,N_487,In_2210);
and U509 (N_509,In_2256,In_1170);
nor U510 (N_510,In_2249,In_892);
and U511 (N_511,In_2420,In_1878);
nand U512 (N_512,N_121,In_493);
nor U513 (N_513,In_1655,In_1831);
or U514 (N_514,In_1737,In_2528);
xor U515 (N_515,In_289,In_56);
nand U516 (N_516,N_92,In_1642);
and U517 (N_517,In_1149,In_2710);
xor U518 (N_518,In_305,N_336);
nor U519 (N_519,In_1381,In_1436);
or U520 (N_520,In_2795,In_836);
and U521 (N_521,In_1674,In_980);
xnor U522 (N_522,In_2940,In_1188);
xnor U523 (N_523,In_251,In_793);
and U524 (N_524,In_2707,In_1195);
nor U525 (N_525,N_187,In_634);
nand U526 (N_526,In_1190,In_1314);
xnor U527 (N_527,In_2363,In_1841);
nor U528 (N_528,In_427,In_2521);
xor U529 (N_529,In_566,In_1374);
nor U530 (N_530,In_109,In_2694);
xnor U531 (N_531,In_676,In_2723);
xnor U532 (N_532,In_2995,In_352);
xor U533 (N_533,In_667,N_184);
xnor U534 (N_534,In_2280,In_1616);
xor U535 (N_535,N_181,In_2618);
nor U536 (N_536,In_1241,N_344);
and U537 (N_537,In_1604,In_2548);
or U538 (N_538,N_286,In_812);
nand U539 (N_539,In_1859,In_2806);
and U540 (N_540,N_428,In_2095);
xnor U541 (N_541,In_1628,In_287);
nand U542 (N_542,N_258,In_1363);
or U543 (N_543,In_2635,In_2421);
or U544 (N_544,In_665,In_2134);
or U545 (N_545,In_2392,In_32);
nand U546 (N_546,In_1802,In_2266);
xor U547 (N_547,In_442,In_2755);
and U548 (N_548,N_491,N_294);
nand U549 (N_549,In_349,In_1876);
or U550 (N_550,In_2721,In_252);
or U551 (N_551,N_17,N_305);
nor U552 (N_552,N_454,N_485);
nor U553 (N_553,In_1630,In_949);
or U554 (N_554,In_1094,In_376);
xor U555 (N_555,N_430,In_1093);
and U556 (N_556,In_2484,In_2810);
xor U557 (N_557,In_149,In_2086);
xor U558 (N_558,In_1005,In_2444);
or U559 (N_559,In_2700,In_872);
xnor U560 (N_560,In_2053,In_2380);
or U561 (N_561,In_799,In_1888);
xnor U562 (N_562,In_1696,In_567);
and U563 (N_563,In_218,In_1877);
and U564 (N_564,In_1858,N_363);
nor U565 (N_565,In_2160,In_1179);
or U566 (N_566,N_240,N_453);
xor U567 (N_567,In_469,In_259);
and U568 (N_568,In_2679,In_2899);
nor U569 (N_569,In_709,In_2430);
and U570 (N_570,In_229,In_1918);
or U571 (N_571,In_2942,In_2559);
or U572 (N_572,In_2791,N_367);
or U573 (N_573,In_394,In_742);
xnor U574 (N_574,In_2,In_1335);
nor U575 (N_575,In_248,In_2060);
nand U576 (N_576,In_1530,In_1926);
nor U577 (N_577,In_452,In_822);
or U578 (N_578,N_86,N_333);
or U579 (N_579,N_29,In_947);
nor U580 (N_580,In_746,In_554);
nor U581 (N_581,In_2647,In_2358);
nor U582 (N_582,In_1668,In_2708);
and U583 (N_583,N_405,In_613);
nor U584 (N_584,In_100,In_1039);
and U585 (N_585,In_841,N_340);
xnor U586 (N_586,In_110,In_1410);
xor U587 (N_587,In_2966,In_2716);
nand U588 (N_588,In_2870,In_1708);
xnor U589 (N_589,In_2768,N_417);
xnor U590 (N_590,In_188,In_992);
or U591 (N_591,In_2459,In_223);
nand U592 (N_592,In_1172,In_1365);
xnor U593 (N_593,In_136,N_10);
nand U594 (N_594,In_2288,In_1607);
xnor U595 (N_595,In_1360,N_310);
or U596 (N_596,In_2994,In_1167);
and U597 (N_597,In_2284,In_195);
nand U598 (N_598,In_94,In_2701);
or U599 (N_599,In_277,In_646);
and U600 (N_600,In_97,In_2171);
or U601 (N_601,In_975,In_2338);
and U602 (N_602,In_183,In_245);
xor U603 (N_603,N_391,In_831);
nand U604 (N_604,In_199,In_2056);
xnor U605 (N_605,N_107,N_115);
nand U606 (N_606,In_1518,In_741);
nand U607 (N_607,In_2591,In_809);
nor U608 (N_608,N_119,N_467);
xnor U609 (N_609,In_952,In_2124);
nor U610 (N_610,N_163,In_1725);
xnor U611 (N_611,In_1236,In_1763);
nor U612 (N_612,In_2872,In_1544);
and U613 (N_613,N_99,In_467);
or U614 (N_614,N_134,N_388);
nand U615 (N_615,In_2130,In_1767);
and U616 (N_616,In_404,In_415);
nand U617 (N_617,In_73,In_2602);
nand U618 (N_618,N_355,In_1457);
and U619 (N_619,In_2963,In_2584);
xnor U620 (N_620,In_887,In_2900);
nor U621 (N_621,N_243,In_2128);
nand U622 (N_622,In_1414,In_1594);
nand U623 (N_623,In_1238,In_1124);
or U624 (N_624,In_2272,In_1091);
nor U625 (N_625,In_768,In_1962);
or U626 (N_626,In_2301,In_2432);
or U627 (N_627,In_2155,N_167);
or U628 (N_628,In_2276,In_413);
nand U629 (N_629,N_324,N_80);
xor U630 (N_630,In_408,In_638);
nor U631 (N_631,In_1635,In_2767);
and U632 (N_632,N_103,In_917);
nand U633 (N_633,In_2855,In_1897);
xor U634 (N_634,In_895,In_361);
xnor U635 (N_635,In_450,In_1829);
and U636 (N_636,In_1239,In_2980);
nand U637 (N_637,In_944,N_456);
or U638 (N_638,N_106,N_277);
nand U639 (N_639,In_1770,In_1546);
or U640 (N_640,In_1027,In_2547);
nand U641 (N_641,In_511,In_295);
nand U642 (N_642,In_714,In_2698);
xor U643 (N_643,In_2993,N_283);
and U644 (N_644,In_507,In_1886);
nor U645 (N_645,In_2449,In_2971);
xnor U646 (N_646,In_710,N_227);
nor U647 (N_647,In_2485,In_2282);
or U648 (N_648,In_2057,In_1543);
xor U649 (N_649,In_1761,In_2204);
xor U650 (N_650,In_1785,In_2724);
and U651 (N_651,In_1850,In_2704);
or U652 (N_652,In_2147,In_2570);
nor U653 (N_653,In_2048,In_2929);
nand U654 (N_654,N_199,In_2429);
and U655 (N_655,In_439,In_2022);
nor U656 (N_656,N_46,In_269);
nor U657 (N_657,In_2145,In_2267);
and U658 (N_658,In_557,In_2992);
nor U659 (N_659,In_2030,N_322);
nor U660 (N_660,In_998,In_2669);
and U661 (N_661,In_897,In_1490);
or U662 (N_662,In_642,In_1707);
or U663 (N_663,In_1318,In_1107);
nand U664 (N_664,In_1865,N_248);
or U665 (N_665,N_130,In_430);
or U666 (N_666,N_202,In_1090);
and U667 (N_667,N_6,In_62);
and U668 (N_668,In_1121,In_2025);
nor U669 (N_669,N_136,In_1223);
and U670 (N_670,In_946,In_1086);
xor U671 (N_671,In_45,In_1140);
nand U672 (N_672,In_406,In_2837);
nor U673 (N_673,In_410,In_853);
or U674 (N_674,In_1610,N_285);
xor U675 (N_675,N_465,In_2776);
or U676 (N_676,In_2325,In_454);
nor U677 (N_677,In_2069,In_2722);
nor U678 (N_678,N_237,In_854);
xnor U679 (N_679,In_1066,N_32);
nand U680 (N_680,N_330,In_151);
nand U681 (N_681,In_771,In_1431);
and U682 (N_682,In_1526,In_1129);
and U683 (N_683,In_2836,In_2648);
and U684 (N_684,In_2137,In_2726);
nand U685 (N_685,In_1606,N_341);
and U686 (N_686,In_2036,N_83);
or U687 (N_687,N_471,In_2586);
xnor U688 (N_688,In_562,N_200);
nand U689 (N_689,In_850,In_1416);
nor U690 (N_690,N_198,In_120);
or U691 (N_691,In_914,In_821);
nand U692 (N_692,N_188,In_973);
nand U693 (N_693,In_1603,N_316);
nor U694 (N_694,N_386,N_444);
or U695 (N_695,N_139,N_224);
or U696 (N_696,In_1548,In_479);
nor U697 (N_697,N_265,In_2910);
xnor U698 (N_698,In_906,In_2211);
nor U699 (N_699,In_2016,In_1440);
xor U700 (N_700,N_249,In_1907);
xor U701 (N_701,In_2453,In_1067);
and U702 (N_702,In_995,N_169);
or U703 (N_703,In_1810,In_228);
nor U704 (N_704,In_2808,In_1139);
and U705 (N_705,In_262,In_436);
xnor U706 (N_706,In_1727,In_2657);
and U707 (N_707,In_1014,In_737);
nand U708 (N_708,In_2555,N_79);
xor U709 (N_709,N_241,In_1052);
and U710 (N_710,In_283,In_1685);
and U711 (N_711,In_1964,N_89);
and U712 (N_712,In_2849,N_247);
and U713 (N_713,N_66,N_353);
or U714 (N_714,In_1283,In_2099);
or U715 (N_715,N_164,In_2874);
and U716 (N_716,In_888,In_2731);
nand U717 (N_717,N_255,In_379);
and U718 (N_718,In_2912,In_1466);
or U719 (N_719,In_845,In_2342);
and U720 (N_720,In_2365,In_1405);
and U721 (N_721,In_2893,In_1873);
and U722 (N_722,In_1315,In_2906);
and U723 (N_723,In_124,In_2455);
xnor U724 (N_724,N_172,In_2161);
or U725 (N_725,In_1221,N_175);
xnor U726 (N_726,In_1912,In_2945);
xnor U727 (N_727,In_1291,In_2192);
nor U728 (N_728,In_2886,In_1820);
nand U729 (N_729,In_1113,N_102);
and U730 (N_730,In_2244,In_2841);
nor U731 (N_731,In_148,In_2381);
and U732 (N_732,In_1452,In_117);
xor U733 (N_733,In_2083,In_1015);
or U734 (N_734,N_424,In_2283);
or U735 (N_735,In_38,In_1250);
or U736 (N_736,N_358,N_362);
or U737 (N_737,In_70,In_202);
nand U738 (N_738,N_141,In_1279);
or U739 (N_739,In_2346,In_581);
nand U740 (N_740,In_2638,N_315);
nand U741 (N_741,In_1994,In_2085);
nor U742 (N_742,N_53,In_2541);
and U743 (N_743,In_1844,In_569);
xnor U744 (N_744,In_2375,In_2273);
nor U745 (N_745,In_1327,In_2609);
nor U746 (N_746,In_1217,In_1101);
nand U747 (N_747,In_1042,In_1826);
nor U748 (N_748,In_1999,In_1881);
and U749 (N_749,In_230,In_2024);
and U750 (N_750,In_1151,In_528);
nand U751 (N_751,In_31,In_294);
nor U752 (N_752,In_1445,In_1910);
or U753 (N_753,In_1687,In_2067);
nand U754 (N_754,In_344,N_496);
nand U755 (N_755,N_156,In_128);
xnor U756 (N_756,In_2351,In_2368);
nand U757 (N_757,In_675,In_1857);
xor U758 (N_758,In_2165,In_1752);
or U759 (N_759,In_1242,In_1419);
nor U760 (N_760,In_1114,In_1522);
nand U761 (N_761,In_1626,In_2196);
or U762 (N_762,N_111,In_1592);
nor U763 (N_763,In_2007,In_2803);
or U764 (N_764,N_489,In_2139);
xor U765 (N_765,In_2691,In_1599);
nor U766 (N_766,In_1681,In_2579);
or U767 (N_767,In_481,In_2466);
xor U768 (N_768,In_2236,In_1661);
xor U769 (N_769,In_2241,In_2506);
xor U770 (N_770,In_575,In_2911);
nor U771 (N_771,In_1678,In_1656);
xor U772 (N_772,In_1762,In_424);
nand U773 (N_773,In_1155,In_1709);
nor U774 (N_774,N_71,In_336);
and U775 (N_775,N_311,In_2811);
and U776 (N_776,In_943,N_72);
xor U777 (N_777,In_1050,In_1579);
or U778 (N_778,N_90,In_2489);
or U779 (N_779,In_1435,In_1570);
or U780 (N_780,In_412,In_1324);
nor U781 (N_781,In_1385,In_2975);
nand U782 (N_782,In_2896,In_314);
xor U783 (N_783,In_2522,N_392);
or U784 (N_784,In_114,In_2374);
xnor U785 (N_785,In_1341,In_1013);
nor U786 (N_786,N_185,In_1750);
or U787 (N_787,In_2033,In_13);
or U788 (N_788,In_14,In_2119);
nor U789 (N_789,In_1429,In_785);
nor U790 (N_790,In_1163,N_273);
or U791 (N_791,N_75,N_421);
or U792 (N_792,In_874,In_1147);
or U793 (N_793,In_1990,In_2600);
nor U794 (N_794,In_176,In_1813);
xnor U795 (N_795,In_2135,In_2876);
nor U796 (N_796,In_2170,In_2289);
xnor U797 (N_797,In_1986,In_1913);
xnor U798 (N_798,In_775,In_470);
or U799 (N_799,In_1679,In_282);
xnor U800 (N_800,In_242,In_2564);
or U801 (N_801,In_1422,In_2109);
xor U802 (N_802,In_2457,In_1266);
xnor U803 (N_803,In_1712,In_1397);
or U804 (N_804,In_1516,In_438);
and U805 (N_805,N_55,In_986);
nor U806 (N_806,In_2587,In_27);
nor U807 (N_807,In_139,In_1312);
xor U808 (N_808,In_288,In_266);
nor U809 (N_809,In_2640,In_585);
nor U810 (N_810,In_2123,In_2319);
or U811 (N_811,In_2422,In_632);
nor U812 (N_812,N_261,In_58);
and U813 (N_813,In_2937,In_463);
and U814 (N_814,In_514,In_1566);
xor U815 (N_815,In_844,In_996);
xor U816 (N_816,In_138,In_508);
and U817 (N_817,N_372,In_2917);
xnor U818 (N_818,N_234,In_2492);
or U819 (N_819,N_342,N_398);
and U820 (N_820,In_1662,In_2608);
nor U821 (N_821,In_2553,In_2916);
nand U822 (N_822,In_1513,N_382);
nor U823 (N_823,In_2316,N_82);
or U824 (N_824,N_266,In_2077);
and U825 (N_825,In_341,In_1293);
or U826 (N_826,In_1786,In_2857);
nor U827 (N_827,N_412,N_37);
or U828 (N_828,N_2,In_34);
nand U829 (N_829,In_2658,In_1021);
xor U830 (N_830,In_1789,In_15);
and U831 (N_831,In_911,In_2005);
nor U832 (N_832,In_1906,N_127);
and U833 (N_833,In_2491,In_280);
and U834 (N_834,N_289,In_982);
xor U835 (N_835,In_2697,N_153);
xor U836 (N_836,In_378,In_1126);
nand U837 (N_837,In_243,N_443);
and U838 (N_838,In_876,In_432);
nor U839 (N_839,In_2168,N_78);
or U840 (N_840,In_1601,In_2035);
nor U841 (N_841,In_2303,In_145);
or U842 (N_842,In_1896,In_2606);
or U843 (N_843,In_1210,In_1189);
nand U844 (N_844,In_1145,In_2366);
and U845 (N_845,In_153,In_306);
and U846 (N_846,In_133,In_825);
xor U847 (N_847,In_1751,In_1305);
xnor U848 (N_848,In_1991,In_2227);
xnor U849 (N_849,In_453,In_2427);
or U850 (N_850,In_1942,In_2516);
nand U851 (N_851,In_2029,In_246);
nor U852 (N_852,In_2894,In_74);
and U853 (N_853,In_609,In_977);
xnor U854 (N_854,In_2792,In_2480);
or U855 (N_855,N_168,In_1706);
nand U856 (N_856,In_2909,In_1136);
nor U857 (N_857,In_1284,In_422);
or U858 (N_858,N_262,In_1677);
or U859 (N_859,In_115,In_544);
and U860 (N_860,In_1993,In_529);
xor U861 (N_861,N_235,In_2122);
or U862 (N_862,In_272,N_117);
xnor U863 (N_863,In_2612,N_36);
nand U864 (N_864,In_2627,In_1699);
xnor U865 (N_865,In_2780,N_290);
and U866 (N_866,In_2882,In_44);
xor U867 (N_867,In_5,In_1641);
or U868 (N_868,N_442,In_2102);
nor U869 (N_869,In_2673,N_365);
or U870 (N_870,In_1775,In_1676);
nor U871 (N_871,In_491,In_968);
xor U872 (N_872,In_1394,N_406);
and U873 (N_873,In_181,In_520);
nand U874 (N_874,In_112,N_14);
nor U875 (N_875,In_296,In_1978);
xor U876 (N_876,In_2977,N_334);
or U877 (N_877,In_377,In_1379);
nor U878 (N_878,In_172,In_1133);
or U879 (N_879,In_688,In_2163);
or U880 (N_880,In_37,N_380);
and U881 (N_881,In_276,In_1639);
xor U882 (N_882,In_2852,In_1760);
xor U883 (N_883,In_1564,N_396);
nand U884 (N_884,In_1225,In_1146);
and U885 (N_885,In_779,In_2383);
and U886 (N_886,N_345,In_899);
xnor U887 (N_887,In_1740,In_2416);
or U888 (N_888,In_213,In_2678);
xor U889 (N_889,In_197,In_505);
and U890 (N_890,In_1103,In_2536);
xor U891 (N_891,In_525,In_707);
or U892 (N_892,In_2068,In_2817);
nand U893 (N_893,In_46,In_1280);
xnor U894 (N_894,In_1805,In_2185);
and U895 (N_895,In_1449,N_77);
nand U896 (N_896,In_2164,N_41);
nand U897 (N_897,In_2084,In_2610);
nor U898 (N_898,In_1308,N_288);
nor U899 (N_899,In_1631,In_849);
or U900 (N_900,In_729,In_1174);
and U901 (N_901,In_784,In_1112);
nand U902 (N_902,In_568,In_2237);
or U903 (N_903,N_201,N_219);
or U904 (N_904,In_2953,N_390);
nor U905 (N_905,N_320,In_2373);
and U906 (N_906,In_2668,In_1575);
nor U907 (N_907,In_2845,N_230);
or U908 (N_908,In_971,In_615);
and U909 (N_909,In_2740,In_298);
nand U910 (N_910,In_732,N_360);
and U911 (N_911,N_174,In_1396);
xor U912 (N_912,N_154,N_226);
xnor U913 (N_913,In_1354,In_2967);
or U914 (N_914,In_1860,In_1285);
and U915 (N_915,In_184,In_1966);
nand U916 (N_916,In_1068,In_2071);
xnor U917 (N_917,In_2595,In_2224);
and U918 (N_918,In_2577,In_1943);
or U919 (N_919,In_1969,In_241);
xnor U920 (N_920,In_808,In_1325);
xor U921 (N_921,In_207,In_1667);
xor U922 (N_922,In_1302,In_2143);
or U923 (N_923,In_2474,In_1033);
or U924 (N_924,In_2660,N_495);
xor U925 (N_925,In_1196,In_517);
or U926 (N_926,In_1088,In_1156);
nand U927 (N_927,In_1794,N_1);
nand U928 (N_928,In_1087,In_2399);
nor U929 (N_929,In_23,In_364);
or U930 (N_930,In_2542,In_2285);
nor U931 (N_931,In_1862,In_735);
and U932 (N_932,In_249,In_89);
nor U933 (N_933,In_1764,In_657);
nor U934 (N_934,N_132,In_760);
nor U935 (N_935,In_951,In_1448);
or U936 (N_936,In_1908,In_2054);
nor U937 (N_937,In_2524,In_1384);
nand U938 (N_938,In_1192,In_212);
and U939 (N_939,In_2044,N_173);
nand U940 (N_940,In_1944,In_2349);
nor U941 (N_941,N_196,N_429);
xnor U942 (N_942,In_1071,In_327);
and U943 (N_943,In_316,In_1048);
or U944 (N_944,In_759,In_645);
xor U945 (N_945,In_859,In_2913);
nor U946 (N_946,In_275,In_1152);
and U947 (N_947,N_420,N_4);
xor U948 (N_948,In_2059,In_171);
xor U949 (N_949,In_2456,N_157);
xor U950 (N_950,In_1584,In_1924);
nor U951 (N_951,In_2797,In_485);
or U952 (N_952,In_1065,In_1319);
and U953 (N_953,In_317,In_1205);
and U954 (N_954,N_313,In_597);
xnor U955 (N_955,In_2978,N_158);
and U956 (N_956,In_2652,In_680);
and U957 (N_957,N_371,In_1349);
or U958 (N_958,In_2644,In_301);
nor U959 (N_959,In_559,In_1296);
xor U960 (N_960,In_2891,In_2226);
nand U961 (N_961,In_405,In_1836);
nand U962 (N_962,In_2557,In_11);
nand U963 (N_963,In_2662,In_2264);
and U964 (N_964,In_198,In_717);
nand U965 (N_965,In_375,In_885);
and U966 (N_966,N_109,In_1292);
or U967 (N_967,In_795,In_2188);
nor U968 (N_968,In_1921,In_2756);
nand U969 (N_969,N_483,In_556);
and U970 (N_970,N_463,In_976);
and U971 (N_971,In_2884,In_2072);
xor U972 (N_972,N_461,In_1615);
and U973 (N_973,In_39,N_312);
nor U974 (N_974,In_2888,In_2153);
nor U975 (N_975,N_20,In_852);
xor U976 (N_976,In_300,N_165);
nand U977 (N_977,In_2031,In_838);
or U978 (N_978,In_2087,N_33);
nor U979 (N_979,In_896,In_869);
or U980 (N_980,N_26,In_2257);
nand U981 (N_981,N_138,In_920);
nand U982 (N_982,In_338,In_962);
nand U983 (N_983,In_2233,In_726);
or U984 (N_984,N_400,In_455);
nand U985 (N_985,In_2948,In_2684);
xor U986 (N_986,In_2393,N_474);
or U987 (N_987,In_1576,In_2621);
or U988 (N_988,In_1456,In_2269);
and U989 (N_989,In_2038,In_474);
nor U990 (N_990,In_106,N_143);
or U991 (N_991,In_555,In_840);
and U992 (N_992,In_1714,In_2907);
or U993 (N_993,N_124,In_1214);
nand U994 (N_994,N_293,In_1352);
nand U995 (N_995,In_2414,In_429);
nand U996 (N_996,N_15,In_2120);
and U997 (N_997,In_2318,In_1184);
or U998 (N_998,In_2409,N_329);
nand U999 (N_999,N_120,N_97);
nand U1000 (N_1000,N_794,N_512);
and U1001 (N_1001,In_2218,N_960);
and U1002 (N_1002,N_784,In_49);
and U1003 (N_1003,In_270,In_2198);
xnor U1004 (N_1004,N_620,In_332);
xor U1005 (N_1005,In_1187,In_1520);
xnor U1006 (N_1006,In_402,N_662);
nor U1007 (N_1007,N_499,In_2956);
nor U1008 (N_1008,In_2921,N_628);
and U1009 (N_1009,In_1741,N_85);
or U1010 (N_1010,In_696,N_900);
or U1011 (N_1011,N_950,In_1487);
xnor U1012 (N_1012,N_395,N_800);
xor U1013 (N_1013,N_547,N_318);
nand U1014 (N_1014,In_711,N_559);
xor U1015 (N_1015,In_2026,In_1476);
or U1016 (N_1016,In_1528,In_93);
nor U1017 (N_1017,In_2959,In_1618);
or U1018 (N_1018,In_2838,In_374);
nor U1019 (N_1019,In_292,In_169);
nor U1020 (N_1020,In_2620,In_1497);
nor U1021 (N_1021,N_690,N_770);
or U1022 (N_1022,In_2592,In_1383);
xor U1023 (N_1023,N_928,In_2969);
and U1024 (N_1024,N_688,In_1040);
xnor U1025 (N_1025,N_566,In_1328);
xnor U1026 (N_1026,N_629,In_589);
and U1027 (N_1027,In_776,In_2344);
xor U1028 (N_1028,In_179,In_767);
and U1029 (N_1029,N_212,N_445);
nor U1030 (N_1030,N_588,N_296);
xnor U1031 (N_1031,In_335,In_2299);
nor U1032 (N_1032,In_1624,In_329);
and U1033 (N_1033,In_1952,N_271);
or U1034 (N_1034,N_549,In_1551);
xnor U1035 (N_1035,In_2473,In_2828);
or U1036 (N_1036,In_367,In_1274);
xnor U1037 (N_1037,In_553,N_408);
nor U1038 (N_1038,N_870,In_2202);
nor U1039 (N_1039,In_1120,N_644);
nor U1040 (N_1040,In_2255,N_686);
or U1041 (N_1041,N_128,N_700);
nor U1042 (N_1042,In_2751,In_2918);
nor U1043 (N_1043,In_477,N_221);
and U1044 (N_1044,N_706,N_675);
or U1045 (N_1045,N_519,In_2619);
xor U1046 (N_1046,N_793,In_2125);
xor U1047 (N_1047,In_1273,In_227);
nand U1048 (N_1048,In_923,In_1342);
nand U1049 (N_1049,N_571,In_2293);
xor U1050 (N_1050,N_192,In_2488);
and U1051 (N_1051,In_1538,In_2475);
or U1052 (N_1052,In_2830,In_1046);
nand U1053 (N_1053,In_2702,N_632);
nand U1054 (N_1054,In_2923,In_2451);
and U1055 (N_1055,In_2772,N_835);
and U1056 (N_1056,In_2046,In_1643);
and U1057 (N_1057,In_36,In_1415);
nand U1058 (N_1058,N_44,N_81);
nor U1059 (N_1059,In_2260,N_730);
or U1060 (N_1060,N_609,N_350);
and U1061 (N_1061,In_1226,In_1759);
or U1062 (N_1062,In_1798,In_2220);
xor U1063 (N_1063,N_28,N_811);
nand U1064 (N_1064,In_2186,In_2507);
and U1065 (N_1065,In_1776,N_3);
or U1066 (N_1066,N_741,N_778);
xor U1067 (N_1067,In_2777,In_2304);
or U1068 (N_1068,In_2743,N_681);
xor U1069 (N_1069,N_116,In_685);
and U1070 (N_1070,N_307,N_397);
and U1071 (N_1071,In_1928,In_518);
and U1072 (N_1072,In_2885,N_570);
nand U1073 (N_1073,In_2232,N_69);
nor U1074 (N_1074,In_1057,N_481);
or U1075 (N_1075,N_972,In_2847);
and U1076 (N_1076,In_1173,In_681);
xor U1077 (N_1077,N_711,In_2711);
or U1078 (N_1078,N_8,In_2989);
nor U1079 (N_1079,N_954,In_603);
nor U1080 (N_1080,In_1704,N_100);
or U1081 (N_1081,In_92,N_713);
or U1082 (N_1082,N_957,In_214);
or U1083 (N_1083,In_323,In_539);
xnor U1084 (N_1084,N_785,In_257);
and U1085 (N_1085,In_66,In_580);
or U1086 (N_1086,N_653,N_771);
nand U1087 (N_1087,In_205,In_1486);
nor U1088 (N_1088,N_510,In_2593);
nor U1089 (N_1089,In_2552,In_2172);
nor U1090 (N_1090,In_720,N_869);
and U1091 (N_1091,In_2832,In_1450);
or U1092 (N_1092,N_921,In_326);
nor U1093 (N_1093,In_2364,In_363);
or U1094 (N_1094,In_1248,In_2331);
nor U1095 (N_1095,N_149,In_2415);
or U1096 (N_1096,In_1945,N_611);
and U1097 (N_1097,In_1930,In_2881);
and U1098 (N_1098,N_193,N_938);
nand U1099 (N_1099,In_777,In_1311);
or U1100 (N_1100,In_2133,N_142);
or U1101 (N_1101,In_846,N_671);
xnor U1102 (N_1102,N_695,In_1542);
nor U1103 (N_1103,In_2157,N_634);
nand U1104 (N_1104,In_1911,In_1075);
nor U1105 (N_1105,N_742,In_1502);
nor U1106 (N_1106,N_792,In_64);
nand U1107 (N_1107,In_1728,In_1203);
or U1108 (N_1108,In_2877,N_663);
nand U1109 (N_1109,In_1933,In_1118);
nand U1110 (N_1110,N_551,In_1778);
nor U1111 (N_1111,In_1219,In_993);
nor U1112 (N_1112,In_1900,N_338);
nor U1113 (N_1113,In_2571,In_903);
and U1114 (N_1114,In_2588,In_1473);
or U1115 (N_1115,In_1412,In_2582);
nor U1116 (N_1116,In_2041,N_446);
xnor U1117 (N_1117,In_918,In_2866);
or U1118 (N_1118,N_804,N_744);
and U1119 (N_1119,In_1463,In_155);
nor U1120 (N_1120,In_1451,N_843);
nand U1121 (N_1121,In_2169,N_801);
or U1122 (N_1122,In_1932,N_451);
and U1123 (N_1123,In_51,In_311);
nand U1124 (N_1124,N_905,N_473);
and U1125 (N_1125,N_655,N_601);
xnor U1126 (N_1126,In_267,In_924);
nand U1127 (N_1127,N_351,In_1682);
xnor U1128 (N_1128,In_1673,In_2078);
nor U1129 (N_1129,In_1869,In_1927);
xor U1130 (N_1130,N_60,N_970);
nand U1131 (N_1131,In_1843,In_622);
nand U1132 (N_1132,In_2179,In_168);
and U1133 (N_1133,N_593,N_978);
xor U1134 (N_1134,N_104,N_849);
xor U1135 (N_1135,N_245,In_2631);
nor U1136 (N_1136,In_2934,N_739);
and U1137 (N_1137,N_375,N_981);
xnor U1138 (N_1138,N_812,In_1931);
and U1139 (N_1139,N_608,In_2946);
or U1140 (N_1140,N_833,N_934);
nand U1141 (N_1141,In_1240,N_546);
nand U1142 (N_1142,N_971,N_458);
and U1143 (N_1143,N_359,In_2535);
or U1144 (N_1144,In_72,In_1777);
or U1145 (N_1145,N_162,In_881);
or U1146 (N_1146,In_1562,N_225);
xnor U1147 (N_1147,N_238,In_211);
xnor U1148 (N_1148,In_254,In_2583);
nor U1149 (N_1149,In_2390,In_2317);
nand U1150 (N_1150,N_328,N_592);
and U1151 (N_1151,In_1024,N_874);
xor U1152 (N_1152,N_821,In_2867);
nand U1153 (N_1153,In_2540,In_1037);
nand U1154 (N_1154,N_679,N_466);
xor U1155 (N_1155,N_579,In_475);
xor U1156 (N_1156,N_246,N_21);
nand U1157 (N_1157,N_683,N_685);
and U1158 (N_1158,In_403,N_684);
and U1159 (N_1159,N_384,N_822);
nor U1160 (N_1160,N_795,N_478);
xnor U1161 (N_1161,N_303,N_949);
and U1162 (N_1162,N_698,In_125);
and U1163 (N_1163,N_511,N_543);
nand U1164 (N_1164,N_976,In_936);
nand U1165 (N_1165,In_194,N_737);
nor U1166 (N_1166,N_58,In_1085);
or U1167 (N_1167,In_598,In_2919);
or U1168 (N_1168,In_2510,N_278);
and U1169 (N_1169,In_2690,In_2010);
nand U1170 (N_1170,In_462,In_2905);
xor U1171 (N_1171,In_2263,In_2733);
xor U1172 (N_1172,In_2183,N_694);
nand U1173 (N_1173,In_2957,In_2871);
nand U1174 (N_1174,N_990,In_546);
nand U1175 (N_1175,In_2074,N_563);
nor U1176 (N_1176,N_880,N_231);
nor U1177 (N_1177,In_663,In_1200);
and U1178 (N_1178,In_570,In_2039);
or U1179 (N_1179,N_455,In_877);
xor U1180 (N_1180,N_834,In_1290);
xnor U1181 (N_1181,N_595,N_147);
or U1182 (N_1182,N_114,N_468);
nor U1183 (N_1183,N_749,In_2424);
or U1184 (N_1184,N_775,In_2748);
and U1185 (N_1185,In_1077,In_137);
nand U1186 (N_1186,N_719,N_61);
xnor U1187 (N_1187,In_1309,In_643);
nor U1188 (N_1188,In_2298,In_2103);
or U1189 (N_1189,In_2497,In_1938);
nand U1190 (N_1190,In_797,N_179);
nor U1191 (N_1191,In_2936,In_2814);
or U1192 (N_1192,In_423,In_1833);
nand U1193 (N_1193,N_847,N_643);
nor U1194 (N_1194,In_1795,N_497);
or U1195 (N_1195,N_947,In_1125);
and U1196 (N_1196,In_1819,N_924);
nand U1197 (N_1197,N_462,In_1002);
xor U1198 (N_1198,In_2898,N_940);
nor U1199 (N_1199,In_2693,In_1270);
xnor U1200 (N_1200,In_2566,In_560);
nand U1201 (N_1201,In_1295,N_540);
nor U1202 (N_1202,In_43,In_1697);
and U1203 (N_1203,N_746,In_2428);
or U1204 (N_1204,In_2107,N_799);
nand U1205 (N_1205,N_250,N_951);
and U1206 (N_1206,N_531,N_76);
or U1207 (N_1207,N_150,In_1084);
nand U1208 (N_1208,In_416,N_689);
xnor U1209 (N_1209,N_917,In_1953);
xor U1210 (N_1210,In_1590,N_475);
and U1211 (N_1211,In_1199,In_2974);
xnor U1212 (N_1212,N_7,In_535);
nand U1213 (N_1213,In_1056,In_630);
nor U1214 (N_1214,N_524,N_740);
nor U1215 (N_1215,In_501,In_744);
xor U1216 (N_1216,In_1976,In_894);
nor U1217 (N_1217,N_645,In_2590);
xnor U1218 (N_1218,N_418,In_1814);
nand U1219 (N_1219,In_2626,In_536);
nor U1220 (N_1220,In_1756,In_842);
xor U1221 (N_1221,In_2650,N_734);
or U1222 (N_1222,N_640,In_1447);
or U1223 (N_1223,N_817,In_2028);
xor U1224 (N_1224,N_625,In_2055);
and U1225 (N_1225,In_1637,In_1161);
nand U1226 (N_1226,In_1166,N_166);
or U1227 (N_1227,In_2322,N_534);
xor U1228 (N_1228,In_860,In_2181);
nor U1229 (N_1229,In_588,In_616);
nand U1230 (N_1230,N_180,In_1313);
and U1231 (N_1231,In_925,In_902);
xor U1232 (N_1232,In_389,In_50);
or U1233 (N_1233,N_284,In_1903);
nand U1234 (N_1234,N_766,N_892);
xor U1235 (N_1235,In_2049,In_755);
nor U1236 (N_1236,In_1744,In_611);
nor U1237 (N_1237,N_140,N_999);
nor U1238 (N_1238,N_674,In_2802);
xor U1239 (N_1239,N_422,N_427);
and U1240 (N_1240,N_267,N_754);
and U1241 (N_1241,In_978,In_512);
xnor U1242 (N_1242,N_878,N_850);
and U1243 (N_1243,N_370,In_1571);
nand U1244 (N_1244,In_1498,In_708);
nand U1245 (N_1245,In_2908,N_717);
nor U1246 (N_1246,In_2320,In_360);
nand U1247 (N_1247,N_993,In_942);
xnor U1248 (N_1248,N_545,In_2090);
and U1249 (N_1249,In_1692,In_2737);
nand U1250 (N_1250,N_197,In_932);
xor U1251 (N_1251,In_1209,N_926);
nor U1252 (N_1252,N_24,In_1723);
xor U1253 (N_1253,N_263,N_317);
nor U1254 (N_1254,In_1739,In_543);
nor U1255 (N_1255,In_2805,N_431);
or U1256 (N_1256,In_497,In_2311);
nand U1257 (N_1257,In_2426,N_558);
nor U1258 (N_1258,In_1979,In_159);
nor U1259 (N_1259,N_191,In_880);
xor U1260 (N_1260,N_0,In_538);
nand U1261 (N_1261,In_2862,In_2603);
or U1262 (N_1262,N_659,In_1017);
nand U1263 (N_1263,In_369,N_493);
or U1264 (N_1264,In_1413,N_832);
nor U1265 (N_1265,N_859,N_987);
nor U1266 (N_1266,In_348,In_1557);
and U1267 (N_1267,In_1702,N_35);
xnor U1268 (N_1268,In_2774,In_2633);
xnor U1269 (N_1269,In_2011,N_726);
xnor U1270 (N_1270,In_584,In_813);
or U1271 (N_1271,In_1622,In_1237);
xor U1272 (N_1272,In_2928,N_666);
nand U1273 (N_1273,N_789,In_1095);
nor U1274 (N_1274,In_691,In_1856);
or U1275 (N_1275,In_1475,N_881);
and U1276 (N_1276,N_752,In_1418);
or U1277 (N_1277,In_1282,N_251);
nor U1278 (N_1278,N_875,In_397);
xor U1279 (N_1279,N_707,N_300);
xor U1280 (N_1280,N_642,N_963);
nand U1281 (N_1281,N_983,In_2434);
xnor U1282 (N_1282,In_639,N_639);
nand U1283 (N_1283,N_780,N_863);
and U1284 (N_1284,N_379,N_480);
nand U1285 (N_1285,In_1791,In_1909);
or U1286 (N_1286,N_407,N_399);
nand U1287 (N_1287,In_1672,N_904);
xor U1288 (N_1288,In_1904,In_1366);
xor U1289 (N_1289,N_802,N_871);
xnor U1290 (N_1290,In_856,N_916);
nor U1291 (N_1291,In_35,N_577);
and U1292 (N_1292,In_2454,In_1625);
or U1293 (N_1293,In_713,N_743);
or U1294 (N_1294,In_1984,In_1110);
nor U1295 (N_1295,In_2764,In_2407);
xor U1296 (N_1296,In_67,In_689);
or U1297 (N_1297,In_1968,In_1111);
nor U1298 (N_1298,N_439,N_572);
nand U1299 (N_1299,In_1620,In_2275);
or U1300 (N_1300,N_708,N_228);
or U1301 (N_1301,In_1061,In_857);
nand U1302 (N_1302,N_206,N_701);
or U1303 (N_1303,In_2445,In_1531);
xor U1304 (N_1304,In_933,In_719);
and U1305 (N_1305,N_118,In_2699);
and U1306 (N_1306,N_948,N_292);
xor U1307 (N_1307,N_530,In_2820);
nor U1308 (N_1308,In_731,N_244);
nor U1309 (N_1309,N_898,In_356);
xnor U1310 (N_1310,In_1025,In_1758);
and U1311 (N_1311,In_234,In_1032);
and U1312 (N_1312,N_88,In_1426);
and U1313 (N_1313,N_930,In_487);
and U1314 (N_1314,In_2686,In_134);
and U1315 (N_1315,In_215,N_973);
nand U1316 (N_1316,In_1688,In_382);
nor U1317 (N_1317,In_1348,In_807);
nor U1318 (N_1318,In_362,In_1263);
nand U1319 (N_1319,In_2883,In_2860);
nor U1320 (N_1320,In_2558,In_835);
and U1321 (N_1321,In_1260,N_383);
nor U1322 (N_1322,N_9,In_1815);
nand U1323 (N_1323,In_2223,In_1386);
nor U1324 (N_1324,In_273,In_858);
and U1325 (N_1325,N_845,In_2614);
or U1326 (N_1326,In_331,N_486);
or U1327 (N_1327,N_989,In_794);
nor U1328 (N_1328,In_1022,N_30);
and U1329 (N_1329,N_457,N_542);
nand U1330 (N_1330,In_2667,In_1404);
or U1331 (N_1331,N_887,In_1509);
xnor U1332 (N_1332,In_2504,In_1180);
nand U1333 (N_1333,In_2675,N_393);
or U1334 (N_1334,In_637,In_2461);
nor U1335 (N_1335,N_846,N_682);
nor U1336 (N_1336,N_56,In_2222);
or U1337 (N_1337,In_2939,In_855);
and U1338 (N_1338,N_415,In_1846);
nand U1339 (N_1339,In_1574,N_50);
nor U1340 (N_1340,N_419,N_937);
and U1341 (N_1341,N_762,N_669);
nor U1342 (N_1342,In_1080,In_449);
nand U1343 (N_1343,In_703,N_48);
nor U1344 (N_1344,In_1803,In_431);
nand U1345 (N_1345,N_515,N_189);
or U1346 (N_1346,N_918,N_774);
or U1347 (N_1347,N_757,In_1249);
nor U1348 (N_1348,N_631,N_64);
or U1349 (N_1349,In_2388,N_190);
xnor U1350 (N_1350,N_16,N_349);
or U1351 (N_1351,In_522,In_2216);
xor U1352 (N_1352,In_48,In_2796);
nand U1353 (N_1353,In_1060,In_751);
or U1354 (N_1354,In_2784,N_433);
nor U1355 (N_1355,N_220,N_272);
nor U1356 (N_1356,N_460,N_553);
nand U1357 (N_1357,In_1350,N_54);
nor U1358 (N_1358,In_457,In_2490);
nand U1359 (N_1359,In_1003,In_2121);
and U1360 (N_1360,In_958,N_818);
or U1361 (N_1361,N_280,In_2094);
and U1362 (N_1362,In_1164,In_2554);
and U1363 (N_1363,In_2922,In_1264);
nor U1364 (N_1364,N_995,N_105);
xor U1365 (N_1365,In_991,In_2718);
or U1366 (N_1366,N_638,In_2458);
xnor U1367 (N_1367,N_969,In_2047);
and U1368 (N_1368,In_354,In_2518);
nand U1369 (N_1369,N_233,In_2023);
xor U1370 (N_1370,N_872,In_650);
nand U1371 (N_1371,In_969,N_13);
or U1372 (N_1372,N_678,N_729);
nor U1373 (N_1373,N_621,In_333);
nand U1374 (N_1374,In_1690,N_980);
nor U1375 (N_1375,In_57,N_617);
nor U1376 (N_1376,In_2356,In_2794);
or U1377 (N_1377,N_884,In_624);
nor U1378 (N_1378,N_74,In_443);
nand U1379 (N_1379,N_823,N_888);
nand U1380 (N_1380,N_194,N_858);
nand U1381 (N_1381,In_418,N_808);
or U1382 (N_1382,In_2773,In_2981);
or U1383 (N_1383,In_2337,In_471);
xor U1384 (N_1384,N_541,In_2664);
and U1385 (N_1385,In_447,In_321);
or U1386 (N_1386,N_62,N_536);
xor U1387 (N_1387,In_2519,N_504);
and U1388 (N_1388,N_615,In_1259);
or U1389 (N_1389,In_1830,In_1150);
and U1390 (N_1390,N_866,In_129);
and U1391 (N_1391,In_2670,N_654);
or U1392 (N_1392,In_2487,N_438);
nand U1393 (N_1393,N_660,N_155);
nand U1394 (N_1394,In_2851,In_1627);
and U1395 (N_1395,In_2201,In_893);
nand U1396 (N_1396,In_2397,In_2991);
nor U1397 (N_1397,N_909,In_629);
or U1398 (N_1398,N_517,In_631);
xnor U1399 (N_1399,In_2065,In_1053);
or U1400 (N_1400,N_482,In_279);
or U1401 (N_1401,N_661,In_1864);
nand U1402 (N_1402,N_177,N_829);
xnor U1403 (N_1403,N_523,In_814);
nand U1404 (N_1404,N_657,In_2040);
nor U1405 (N_1405,In_602,In_586);
xnor U1406 (N_1406,N_984,In_85);
nor U1407 (N_1407,N_939,N_665);
nor U1408 (N_1408,N_452,N_992);
and U1409 (N_1409,In_1231,N_605);
or U1410 (N_1410,N_529,N_810);
or U1411 (N_1411,In_1533,In_1288);
nor U1412 (N_1412,In_608,N_668);
and U1413 (N_1413,In_2443,In_1834);
nor U1414 (N_1414,N_944,N_366);
nand U1415 (N_1415,In_47,N_647);
xor U1416 (N_1416,N_502,N_712);
and U1417 (N_1417,N_985,In_1634);
or U1418 (N_1418,In_260,In_30);
nand U1419 (N_1419,N_298,In_489);
or U1420 (N_1420,In_1261,In_738);
or U1421 (N_1421,In_788,N_703);
nand U1422 (N_1422,N_368,In_2004);
xor U1423 (N_1423,In_2502,In_2798);
nand U1424 (N_1424,In_91,N_902);
nand U1425 (N_1425,N_844,In_649);
or U1426 (N_1426,N_646,N_738);
or U1427 (N_1427,In_832,N_213);
xnor U1428 (N_1428,In_307,N_434);
nor U1429 (N_1429,In_1306,In_1078);
nand U1430 (N_1430,In_2807,In_2779);
or U1431 (N_1431,In_1400,In_2279);
nor U1432 (N_1432,In_2173,In_126);
nor U1433 (N_1433,N_796,In_862);
xnor U1434 (N_1434,In_891,In_2632);
nand U1435 (N_1435,In_2715,N_448);
or U1436 (N_1436,In_2901,In_1899);
and U1437 (N_1437,N_721,N_895);
xnor U1438 (N_1438,In_1747,In_2062);
xor U1439 (N_1439,In_503,N_574);
and U1440 (N_1440,In_1143,N_513);
and U1441 (N_1441,In_2132,N_988);
or U1442 (N_1442,N_538,N_264);
or U1443 (N_1443,In_2501,In_2350);
and U1444 (N_1444,In_2190,In_1505);
xor U1445 (N_1445,N_323,N_319);
or U1446 (N_1446,In_1076,In_758);
nand U1447 (N_1447,In_882,N_925);
xnor U1448 (N_1448,N_525,In_837);
xnor U1449 (N_1449,In_1855,N_920);
nor U1450 (N_1450,In_669,In_1768);
or U1451 (N_1451,In_187,In_1408);
nor U1452 (N_1452,N_600,N_152);
xor U1453 (N_1453,N_299,N_210);
nand U1454 (N_1454,N_854,In_2271);
nor U1455 (N_1455,In_380,In_1729);
nor U1456 (N_1456,N_648,In_2643);
nand U1457 (N_1457,N_160,In_1973);
nand U1458 (N_1458,N_101,In_541);
and U1459 (N_1459,In_1665,N_133);
nand U1460 (N_1460,In_2842,In_889);
nand U1461 (N_1461,N_348,In_664);
xor U1462 (N_1462,In_2853,In_318);
xnor U1463 (N_1463,N_95,In_233);
nand U1464 (N_1464,N_718,In_1432);
nor U1465 (N_1465,In_1089,N_827);
nor U1466 (N_1466,In_1082,In_830);
or U1467 (N_1467,In_2537,In_820);
nor U1468 (N_1468,In_2248,In_2998);
or U1469 (N_1469,In_1784,In_483);
or U1470 (N_1470,In_800,N_38);
or U1471 (N_1471,N_893,In_2467);
nor U1472 (N_1472,N_636,In_495);
or U1473 (N_1473,N_19,In_1916);
xnor U1474 (N_1474,In_1521,In_177);
nand U1475 (N_1475,N_997,N_325);
nand U1476 (N_1476,N_508,In_1072);
nor U1477 (N_1477,N_47,In_1122);
nand U1478 (N_1478,N_11,In_393);
nor U1479 (N_1479,In_1064,In_1382);
xnor U1480 (N_1480,In_1175,In_524);
or U1481 (N_1481,In_2228,In_189);
nand U1482 (N_1482,In_886,In_2436);
nor U1483 (N_1483,In_2470,In_1339);
xor U1484 (N_1484,In_2759,In_1600);
and U1485 (N_1485,In_1832,N_302);
nand U1486 (N_1486,N_568,N_346);
and U1487 (N_1487,In_1097,In_2513);
nor U1488 (N_1488,N_637,N_603);
and U1489 (N_1489,In_286,In_728);
nand U1490 (N_1490,N_494,In_2509);
nor U1491 (N_1491,N_612,In_2850);
and U1492 (N_1492,In_2118,In_2563);
xor U1493 (N_1493,In_330,In_1996);
or U1494 (N_1494,In_235,N_129);
nand U1495 (N_1495,N_959,N_215);
xor U1496 (N_1496,In_324,In_1376);
or U1497 (N_1497,In_1049,In_2166);
nand U1498 (N_1498,In_2970,N_450);
nor U1499 (N_1499,In_2999,In_2818);
xnor U1500 (N_1500,N_1196,N_1171);
nand U1501 (N_1501,In_75,N_1302);
xnor U1502 (N_1502,N_1425,In_426);
nor U1503 (N_1503,N_624,N_899);
or U1504 (N_1504,N_1111,N_936);
or U1505 (N_1505,N_618,N_1107);
or U1506 (N_1506,N_414,In_113);
nor U1507 (N_1507,N_381,In_1792);
nand U1508 (N_1508,N_906,N_1031);
nor U1509 (N_1509,In_961,N_1319);
nor U1510 (N_1510,In_157,N_1463);
and U1511 (N_1511,N_357,N_1443);
or U1512 (N_1512,In_359,N_146);
xnor U1513 (N_1513,N_394,In_2369);
nor U1514 (N_1514,N_282,In_1417);
nand U1515 (N_1515,In_2008,N_1051);
or U1516 (N_1516,N_1184,In_1894);
nand U1517 (N_1517,N_1094,In_77);
or U1518 (N_1518,In_2746,In_381);
xnor U1519 (N_1519,In_1216,In_674);
nor U1520 (N_1520,In_111,N_1197);
xor U1521 (N_1521,N_522,N_123);
nand U1522 (N_1522,N_556,N_369);
nand U1523 (N_1523,In_1884,In_1286);
nand U1524 (N_1524,N_986,N_1104);
xnor U1525 (N_1525,N_1121,N_377);
nor U1526 (N_1526,N_890,N_720);
nand U1527 (N_1527,In_132,In_1753);
or U1528 (N_1528,N_1233,In_1879);
xor U1529 (N_1529,N_763,N_1312);
nor U1530 (N_1530,N_1317,In_2511);
nor U1531 (N_1531,N_974,N_339);
or U1532 (N_1532,N_1376,N_945);
or U1533 (N_1533,N_1056,In_2448);
nand U1534 (N_1534,In_687,In_2359);
nand U1535 (N_1535,In_792,N_1239);
nand U1536 (N_1536,N_469,N_779);
nor U1537 (N_1537,In_261,In_1914);
nor U1538 (N_1538,In_2903,N_696);
or U1539 (N_1539,N_1260,N_1025);
or U1540 (N_1540,N_387,In_2987);
and U1541 (N_1541,N_1473,N_1354);
and U1542 (N_1542,N_435,In_102);
nand U1543 (N_1543,N_1498,N_1267);
or U1544 (N_1544,N_1261,N_137);
xor U1545 (N_1545,N_376,N_787);
nor U1546 (N_1546,N_923,N_1398);
nor U1547 (N_1547,N_314,N_1296);
and U1548 (N_1548,N_769,N_1371);
or U1549 (N_1549,In_765,N_943);
nor U1550 (N_1550,In_931,N_423);
or U1551 (N_1551,N_891,N_1393);
nand U1552 (N_1552,N_1098,N_1339);
nand U1553 (N_1553,N_1136,In_2127);
and U1554 (N_1554,In_2034,N_548);
xnor U1555 (N_1555,N_1399,N_616);
and U1556 (N_1556,In_1880,In_2212);
or U1557 (N_1557,N_304,N_1346);
nor U1558 (N_1558,In_2020,In_2058);
or U1559 (N_1559,N_52,N_1245);
and U1560 (N_1560,N_1269,N_1206);
xnor U1561 (N_1561,In_743,N_561);
xnor U1562 (N_1562,N_756,N_1347);
xor U1563 (N_1563,In_2483,In_2926);
or U1564 (N_1564,N_1235,N_1004);
nand U1565 (N_1565,N_1357,N_211);
and U1566 (N_1566,In_2017,N_509);
and U1567 (N_1567,N_1385,In_2012);
nand U1568 (N_1568,N_1112,In_178);
or U1569 (N_1569,N_23,N_1274);
xnor U1570 (N_1570,N_1226,N_912);
xor U1571 (N_1571,In_2634,In_446);
xor U1572 (N_1572,In_1333,In_225);
and U1573 (N_1573,In_2141,N_327);
xnor U1574 (N_1574,N_1360,In_1949);
nor U1575 (N_1575,N_1442,In_1561);
or U1576 (N_1576,N_604,N_623);
or U1577 (N_1577,N_797,In_465);
or U1578 (N_1578,In_2326,N_1424);
nand U1579 (N_1579,In_1650,N_1365);
and U1580 (N_1580,In_488,In_2187);
xnor U1581 (N_1581,N_786,In_340);
and U1582 (N_1582,In_1043,N_1223);
and U1583 (N_1583,N_1165,N_1210);
and U1584 (N_1584,N_732,N_1194);
nand U1585 (N_1585,In_618,N_1328);
xnor U1586 (N_1586,N_1258,N_148);
nor U1587 (N_1587,N_1152,In_2431);
xnor U1588 (N_1588,In_2861,N_205);
or U1589 (N_1589,N_1237,N_1096);
nand U1590 (N_1590,N_1423,N_1079);
nor U1591 (N_1591,N_1038,In_1181);
or U1592 (N_1592,In_1009,In_1144);
xor U1593 (N_1593,N_229,N_1071);
nand U1594 (N_1594,N_1147,N_753);
or U1595 (N_1595,In_1975,In_2611);
and U1596 (N_1596,In_2758,N_557);
and U1597 (N_1597,N_544,In_2826);
nor U1598 (N_1598,N_40,In_1501);
nor U1599 (N_1599,In_2199,In_1640);
xor U1600 (N_1600,In_1874,N_65);
nand U1601 (N_1601,N_1007,N_1311);
or U1602 (N_1602,N_1192,In_78);
and U1603 (N_1603,In_1612,In_919);
and U1604 (N_1604,N_1097,N_1040);
nor U1605 (N_1605,In_2270,N_1340);
nand U1606 (N_1606,N_526,In_2219);
xor U1607 (N_1607,In_870,N_865);
xor U1608 (N_1608,In_2089,N_853);
and U1609 (N_1609,In_1330,N_619);
and U1610 (N_1610,N_1234,In_1294);
nand U1611 (N_1611,N_964,N_911);
xor U1612 (N_1612,N_798,N_958);
and U1613 (N_1613,N_1125,In_2646);
nor U1614 (N_1614,In_1228,N_1084);
xor U1615 (N_1615,N_555,In_1281);
xnor U1616 (N_1616,N_977,N_1316);
xor U1617 (N_1617,N_910,In_2960);
or U1618 (N_1618,In_1459,N_1428);
nor U1619 (N_1619,N_1409,N_1497);
nor U1620 (N_1620,N_222,N_1276);
nor U1621 (N_1621,N_326,N_1461);
or U1622 (N_1622,N_354,In_1299);
or U1623 (N_1623,N_1236,N_1222);
and U1624 (N_1624,In_2217,N_1167);
and U1625 (N_1625,N_820,In_816);
or U1626 (N_1626,N_436,N_1127);
and U1627 (N_1627,N_877,N_216);
xnor U1628 (N_1628,N_1366,N_807);
and U1629 (N_1629,N_1065,In_2696);
nor U1630 (N_1630,N_472,N_1413);
nand U1631 (N_1631,N_760,N_1188);
nor U1632 (N_1632,N_1157,N_946);
nand U1633 (N_1633,In_2549,N_1080);
nand U1634 (N_1634,N_236,In_530);
xor U1635 (N_1635,In_291,N_1088);
nand U1636 (N_1636,In_1595,In_55);
and U1637 (N_1637,In_2150,In_2106);
nor U1638 (N_1638,In_2655,In_698);
nand U1639 (N_1639,In_54,In_1980);
xnor U1640 (N_1640,In_343,In_595);
and U1641 (N_1641,N_861,In_1481);
nand U1642 (N_1642,N_814,In_2941);
nor U1643 (N_1643,In_1870,In_2897);
and U1644 (N_1644,N_1395,N_67);
xnor U1645 (N_1645,N_836,N_1087);
and U1646 (N_1646,In_1853,N_49);
xnor U1647 (N_1647,N_1294,In_3);
xor U1648 (N_1648,In_1329,N_710);
and U1649 (N_1649,In_1401,In_302);
xor U1650 (N_1650,N_602,In_658);
or U1651 (N_1651,N_1337,N_907);
nor U1652 (N_1652,In_253,In_1001);
nor U1653 (N_1653,In_591,In_2844);
and U1654 (N_1654,N_1481,In_1028);
or U1655 (N_1655,N_1462,N_1213);
or U1656 (N_1656,N_967,N_1073);
and U1657 (N_1657,N_1465,N_1003);
or U1658 (N_1658,N_1085,N_1266);
and U1659 (N_1659,N_1288,N_1297);
nand U1660 (N_1660,N_782,N_1429);
or U1661 (N_1661,N_1492,N_501);
nor U1662 (N_1662,In_1598,N_673);
xnor U1663 (N_1663,N_965,N_1299);
nor U1664 (N_1664,In_548,In_984);
nor U1665 (N_1665,N_1420,N_941);
nand U1666 (N_1666,N_514,N_565);
nand U1667 (N_1667,N_151,In_1198);
xnor U1668 (N_1668,In_900,N_1050);
nand U1669 (N_1669,N_1190,In_1227);
nand U1670 (N_1670,N_828,In_791);
or U1671 (N_1671,In_1317,In_2043);
nand U1672 (N_1672,N_25,N_1055);
xnor U1673 (N_1673,N_1449,In_204);
nor U1674 (N_1674,N_747,In_2954);
xnor U1675 (N_1675,N_1042,In_2391);
nor U1676 (N_1676,N_492,N_308);
or U1677 (N_1677,In_1901,N_1467);
or U1678 (N_1678,In_1552,In_421);
or U1679 (N_1679,N_715,N_1259);
nor U1680 (N_1680,N_1200,N_256);
nor U1681 (N_1681,In_2687,N_335);
and U1682 (N_1682,In_954,In_2442);
or U1683 (N_1683,N_1006,In_2835);
or U1684 (N_1684,N_1058,In_2370);
xor U1685 (N_1685,N_281,In_864);
or U1686 (N_1686,N_432,In_1470);
nor U1687 (N_1687,N_1209,N_1384);
nor U1688 (N_1688,In_1269,In_1514);
nand U1689 (N_1689,N_1392,N_43);
nor U1690 (N_1690,N_1349,N_1304);
nor U1691 (N_1691,N_864,N_1370);
nor U1692 (N_1692,N_1394,In_1398);
or U1693 (N_1693,N_1397,N_1091);
or U1694 (N_1694,In_1837,In_519);
xnor U1695 (N_1695,In_21,In_1519);
xor U1696 (N_1696,N_705,In_1372);
xnor U1697 (N_1697,N_614,N_781);
xor U1698 (N_1698,In_150,N_1252);
nor U1699 (N_1699,N_1381,In_617);
xnor U1700 (N_1700,N_1135,N_1027);
nand U1701 (N_1701,N_862,N_1156);
nor U1702 (N_1702,In_1351,N_479);
and U1703 (N_1703,N_5,In_131);
or U1704 (N_1704,In_1547,In_659);
or U1705 (N_1705,In_1232,In_2061);
or U1706 (N_1706,In_1488,N_51);
and U1707 (N_1707,N_1407,N_692);
xnor U1708 (N_1708,N_1478,N_1015);
nor U1709 (N_1709,N_96,In_898);
nand U1710 (N_1710,N_1019,N_1453);
nand U1711 (N_1711,In_2920,N_613);
and U1712 (N_1712,N_1179,N_759);
and U1713 (N_1713,N_567,In_2184);
or U1714 (N_1714,N_411,In_2308);
and U1715 (N_1715,In_1941,N_842);
nor U1716 (N_1716,N_598,N_1437);
and U1717 (N_1717,N_1375,In_2019);
or U1718 (N_1718,N_1292,N_1202);
xnor U1719 (N_1719,N_1023,N_1103);
and U1720 (N_1720,In_2253,N_1102);
or U1721 (N_1721,In_945,In_644);
xnor U1722 (N_1722,N_584,N_378);
or U1723 (N_1723,In_1923,N_361);
nor U1724 (N_1724,N_590,N_1321);
and U1725 (N_1725,N_837,In_2355);
or U1726 (N_1726,N_622,N_1132);
xor U1727 (N_1727,N_1369,N_1355);
xnor U1728 (N_1728,In_1303,In_1646);
nor U1729 (N_1729,N_159,N_125);
or U1730 (N_1730,In_1393,In_1099);
and U1731 (N_1731,In_1868,N_1128);
nand U1732 (N_1732,N_532,N_1289);
or U1733 (N_1733,N_309,In_499);
or U1734 (N_1734,N_1279,N_1352);
nor U1735 (N_1735,In_1691,N_223);
nor U1736 (N_1736,In_1669,In_1754);
and U1737 (N_1737,N_750,In_2683);
nor U1738 (N_1738,N_1275,In_2405);
and U1739 (N_1739,N_1363,N_1487);
or U1740 (N_1740,In_1535,N_727);
nor U1741 (N_1741,N_1468,In_7);
xor U1742 (N_1742,N_882,N_1396);
nand U1743 (N_1743,In_2951,In_236);
or U1744 (N_1744,N_57,N_933);
or U1745 (N_1745,N_1219,N_1066);
and U1746 (N_1746,In_1769,In_1336);
nor U1747 (N_1747,In_320,N_239);
or U1748 (N_1748,N_1383,N_724);
nand U1749 (N_1749,In_448,N_488);
or U1750 (N_1750,N_824,In_2865);
nor U1751 (N_1751,N_59,N_1265);
nor U1752 (N_1752,N_606,In_33);
nor U1753 (N_1753,In_2156,In_1780);
and U1754 (N_1754,N_287,N_569);
or U1755 (N_1755,N_1009,In_2763);
xor U1756 (N_1756,In_2468,N_1183);
and U1757 (N_1757,N_1262,N_1263);
and U1758 (N_1758,In_2717,N_1491);
and U1759 (N_1759,N_500,In_312);
nor U1760 (N_1760,In_1633,N_1201);
nor U1761 (N_1761,N_1310,In_1585);
and U1762 (N_1762,N_1187,N_573);
or U1763 (N_1763,In_2265,N_1387);
xor U1764 (N_1764,In_1827,N_404);
xor U1765 (N_1765,In_2935,In_656);
or U1766 (N_1766,N_1224,In_1647);
nand U1767 (N_1767,N_1246,N_1047);
xnor U1768 (N_1768,N_922,In_419);
xor U1769 (N_1769,N_1158,N_1464);
or U1770 (N_1770,N_1014,N_364);
or U1771 (N_1771,In_778,N_1182);
nor U1772 (N_1772,N_1335,In_90);
xnor U1773 (N_1773,In_1029,In_1919);
nand U1774 (N_1774,In_2018,N_840);
nor U1775 (N_1775,N_1030,N_670);
and U1776 (N_1776,N_1060,N_586);
or U1777 (N_1777,In_1482,N_1020);
and U1778 (N_1778,N_1203,In_2636);
or U1779 (N_1779,In_2750,N_758);
nor U1780 (N_1780,In_2050,N_1290);
xnor U1781 (N_1781,N_332,N_352);
xnor U1782 (N_1782,In_2215,N_1212);
and U1783 (N_1783,N_1248,In_1823);
and U1784 (N_1784,In_52,N_254);
nand U1785 (N_1785,N_1460,N_932);
and U1786 (N_1786,N_765,In_2790);
nor U1787 (N_1787,In_2498,N_1277);
or U1788 (N_1788,N_702,N_897);
and U1789 (N_1789,N_704,In_1425);
nor U1790 (N_1790,N_385,In_186);
and U1791 (N_1791,In_1809,N_1140);
nor U1792 (N_1792,In_2754,In_1935);
nor U1793 (N_1793,In_651,In_1508);
or U1794 (N_1794,In_1262,In_2869);
and U1795 (N_1795,N_1083,In_2982);
nand U1796 (N_1796,In_1689,In_1424);
and U1797 (N_1797,N_1000,N_1480);
or U1798 (N_1798,In_1534,In_1902);
or U1799 (N_1799,In_1392,N_952);
and U1800 (N_1800,In_551,N_1013);
xnor U1801 (N_1801,In_395,N_1496);
nand U1802 (N_1802,N_1100,In_1839);
nand U1803 (N_1803,N_1490,N_1314);
nor U1804 (N_1804,In_420,In_1602);
nand U1805 (N_1805,N_1124,In_705);
and U1806 (N_1806,N_723,In_1867);
or U1807 (N_1807,In_1657,In_18);
nor U1808 (N_1808,N_806,N_1048);
or U1809 (N_1809,N_1457,N_830);
or U1810 (N_1810,N_755,N_1122);
and U1811 (N_1811,In_2419,N_1332);
or U1812 (N_1812,In_2348,N_672);
nand U1813 (N_1813,N_1482,N_1113);
or U1814 (N_1814,N_733,N_809);
nor U1815 (N_1815,N_498,In_2114);
and U1816 (N_1816,In_303,In_372);
and U1817 (N_1817,N_135,In_590);
or U1818 (N_1818,In_1790,N_1086);
or U1819 (N_1819,In_2672,N_1011);
or U1820 (N_1820,N_94,N_1388);
nor U1821 (N_1821,N_1181,N_1475);
or U1822 (N_1822,N_1391,N_1456);
nand U1823 (N_1823,N_868,N_1422);
xnor U1824 (N_1824,N_680,N_1307);
nand U1825 (N_1825,N_825,In_193);
nor U1826 (N_1826,N_883,In_2406);
nor U1827 (N_1827,In_2979,N_1318);
or U1828 (N_1828,N_1489,N_1336);
xor U1829 (N_1829,In_1799,N_968);
or U1830 (N_1830,N_1139,In_1345);
nor U1831 (N_1831,In_2408,N_982);
or U1832 (N_1832,In_1500,In_940);
and U1833 (N_1833,N_1110,N_1217);
nand U1834 (N_1834,In_2193,In_704);
and U1835 (N_1835,In_1947,N_1470);
and U1836 (N_1836,N_1198,N_1195);
nand U1837 (N_1837,In_2200,N_1046);
nand U1838 (N_1838,In_2729,In_2747);
nor U1839 (N_1839,In_670,N_1238);
nand U1840 (N_1840,N_994,In_964);
and U1841 (N_1841,In_2902,In_1773);
xnor U1842 (N_1842,N_1255,In_1701);
and U1843 (N_1843,N_204,In_160);
nand U1844 (N_1844,In_912,In_1297);
or U1845 (N_1845,N_126,In_1974);
or U1846 (N_1846,N_667,N_1166);
nand U1847 (N_1847,N_1488,N_585);
and U1848 (N_1848,In_1334,N_1227);
and U1849 (N_1849,N_1151,N_403);
or U1850 (N_1850,In_1364,N_1438);
or U1851 (N_1851,N_505,N_112);
xnor U1852 (N_1852,In_2545,N_1295);
nor U1853 (N_1853,In_780,In_2642);
xor U1854 (N_1854,N_855,In_388);
nand U1855 (N_1855,N_1039,In_1212);
nor U1856 (N_1856,N_1012,In_2362);
and U1857 (N_1857,In_441,In_2823);
and U1858 (N_1858,N_996,N_1469);
xor U1859 (N_1859,N_321,N_1451);
xor U1860 (N_1860,N_913,N_1441);
or U1861 (N_1861,In_527,N_641);
xor U1862 (N_1862,N_1315,N_1035);
nand U1863 (N_1863,N_1325,N_552);
xor U1864 (N_1864,In_2144,In_796);
nand U1865 (N_1865,N_1215,N_1483);
xnor U1866 (N_1866,N_1402,In_473);
nand U1867 (N_1867,N_1145,In_398);
nor U1868 (N_1868,In_2824,In_1127);
or U1869 (N_1869,N_767,In_1517);
and U1870 (N_1870,N_852,In_2354);
nor U1871 (N_1871,In_1117,In_1845);
nand U1872 (N_1872,N_1257,In_1735);
nand U1873 (N_1873,N_176,N_374);
and U1874 (N_1874,In_2812,N_1185);
nor U1875 (N_1875,In_1454,In_152);
or U1876 (N_1876,In_722,N_1010);
nand U1877 (N_1877,N_857,In_1734);
nor U1878 (N_1878,N_1075,In_1961);
or U1879 (N_1879,In_1788,In_1700);
nor U1880 (N_1880,N_1372,N_687);
and U1881 (N_1881,In_1373,In_654);
nand U1882 (N_1882,N_1175,In_1370);
xnor U1883 (N_1883,In_2251,In_1651);
xnor U1884 (N_1884,N_1057,In_2499);
nand U1885 (N_1885,In_2117,N_1495);
or U1886 (N_1886,N_274,N_889);
or U1887 (N_1887,In_9,In_6);
or U1888 (N_1888,N_39,N_1204);
nand U1889 (N_1889,In_417,N_503);
nor U1890 (N_1890,N_1231,N_1106);
xnor U1891 (N_1891,N_1105,N_788);
xnor U1892 (N_1892,In_1109,N_297);
nand U1893 (N_1893,N_1356,In_365);
nor U1894 (N_1894,In_1244,In_1556);
nor U1895 (N_1895,In_2532,In_953);
nand U1896 (N_1896,In_823,N_1123);
xor U1897 (N_1897,N_70,N_1115);
xor U1898 (N_1898,N_1330,N_1300);
or U1899 (N_1899,N_677,N_1404);
nand U1900 (N_1900,N_1242,In_2543);
nand U1901 (N_1901,N_1323,In_693);
xor U1902 (N_1902,N_1414,In_1948);
nand U1903 (N_1903,N_1143,N_728);
or U1904 (N_1904,N_1280,N_961);
nand U1905 (N_1905,In_2829,In_921);
or U1906 (N_1906,N_1286,N_791);
and U1907 (N_1907,N_955,N_751);
nand U1908 (N_1908,In_2438,N_1329);
nor U1909 (N_1909,In_890,N_373);
or U1910 (N_1910,In_1887,In_1331);
and U1911 (N_1911,N_1411,N_1455);
and U1912 (N_1912,N_819,N_1164);
and U1913 (N_1913,N_1240,N_1142);
or U1914 (N_1914,N_1281,In_1011);
and U1915 (N_1915,In_605,In_2637);
and U1916 (N_1916,N_144,N_1241);
and U1917 (N_1917,N_1089,In_2783);
nand U1918 (N_1918,In_2341,N_1434);
and U1919 (N_1919,In_1609,N_630);
nand U1920 (N_1920,N_908,In_414);
and U1921 (N_1921,N_1309,In_2565);
xnor U1922 (N_1922,N_1153,N_91);
and U1923 (N_1923,N_1002,In_209);
and U1924 (N_1924,N_1022,N_18);
nand U1925 (N_1925,In_1193,In_1925);
and U1926 (N_1926,N_1308,In_466);
and U1927 (N_1927,In_2277,N_1028);
or U1928 (N_1928,N_736,In_2482);
nand U1929 (N_1929,N_1220,N_1001);
nand U1930 (N_1930,N_848,N_12);
nand U1931 (N_1931,In_1680,In_1128);
nor U1932 (N_1932,N_1069,In_2904);
and U1933 (N_1933,N_409,In_633);
xor U1934 (N_1934,In_2310,In_2149);
and U1935 (N_1935,N_275,N_440);
or U1936 (N_1936,N_599,In_873);
nand U1937 (N_1937,N_1092,N_1389);
nand U1938 (N_1938,In_1165,In_1421);
nand U1939 (N_1939,N_1477,In_2105);
and U1940 (N_1940,In_552,In_391);
xnor U1941 (N_1941,In_2534,N_93);
and U1942 (N_1942,N_1033,In_700);
nand U1943 (N_1943,In_702,N_1444);
xor U1944 (N_1944,In_1730,In_2972);
nand U1945 (N_1945,N_31,In_2494);
nand U1946 (N_1946,N_161,N_1432);
nor U1947 (N_1947,In_1746,N_1408);
xnor U1948 (N_1948,In_939,N_578);
or U1949 (N_1949,In_2476,In_2092);
nand U1950 (N_1950,In_1960,N_1161);
or U1951 (N_1951,In_594,N_269);
nand U1952 (N_1952,N_268,N_186);
nand U1953 (N_1953,N_217,N_1137);
xnor U1954 (N_1954,In_1153,N_195);
nor U1955 (N_1955,N_1141,In_1304);
nand U1956 (N_1956,N_550,In_2719);
xnor U1957 (N_1957,N_1493,N_633);
xnor U1958 (N_1958,N_1247,N_276);
or U1959 (N_1959,N_773,N_1458);
nor U1960 (N_1960,In_284,N_477);
or U1961 (N_1961,In_346,N_1074);
and U1962 (N_1962,N_533,N_1272);
nor U1963 (N_1963,N_1078,In_2985);
nand U1964 (N_1964,N_714,N_1322);
nor U1965 (N_1965,N_1400,N_1036);
nor U1966 (N_1966,N_1454,N_527);
and U1967 (N_1967,N_635,In_565);
nor U1968 (N_1968,N_182,N_539);
and U1969 (N_1969,N_1082,In_1391);
nand U1970 (N_1970,N_554,In_2741);
nand U1971 (N_1971,N_560,N_761);
or U1972 (N_1972,In_2477,In_1963);
xnor U1973 (N_1973,In_2550,N_113);
xor U1974 (N_1974,N_699,N_232);
xnor U1975 (N_1975,N_596,In_1567);
or U1976 (N_1976,In_1965,In_1955);
nand U1977 (N_1977,N_260,N_343);
and U1978 (N_1978,N_1344,In_904);
nand U1979 (N_1979,In_173,In_264);
and U1980 (N_1980,N_45,In_1387);
or U1981 (N_1981,In_1035,N_1418);
nor U1982 (N_1982,N_1364,N_1447);
and U1983 (N_1983,N_1101,In_753);
or U1984 (N_1984,N_1016,In_1686);
xnor U1985 (N_1985,N_122,In_63);
or U1986 (N_1986,N_1313,N_1271);
xnor U1987 (N_1987,N_975,N_935);
nor U1988 (N_1988,N_1117,In_2858);
or U1989 (N_1989,In_994,N_748);
and U1990 (N_1990,N_1421,N_815);
nor U1991 (N_1991,In_1694,N_1431);
and U1992 (N_1992,In_192,N_1479);
xor U1993 (N_1993,N_518,N_1334);
or U1994 (N_1994,N_953,In_358);
or U1995 (N_1995,N_929,In_866);
nand U1996 (N_1996,In_509,In_42);
and U1997 (N_1997,In_1178,In_2576);
nor U1998 (N_1998,N_63,In_1817);
or U1999 (N_1999,In_506,N_1150);
nand U2000 (N_2000,In_2569,N_1960);
nand U2001 (N_2001,N_1351,In_1905);
or U2002 (N_2002,N_1282,N_1941);
and U2003 (N_2003,N_1927,N_1591);
nand U2004 (N_2004,N_1726,N_1944);
nor U2005 (N_2005,N_1640,N_1534);
and U2006 (N_2006,N_1787,N_1459);
nand U2007 (N_2007,In_1726,N_658);
nor U2008 (N_2008,N_1953,N_1708);
or U2009 (N_2009,N_347,In_2597);
or U2010 (N_2010,N_1807,N_1811);
nor U2011 (N_2011,N_1757,N_1915);
and U2012 (N_2012,N_656,N_1264);
nor U2013 (N_2013,N_1580,N_1064);
xnor U2014 (N_2014,N_1788,N_664);
nor U2015 (N_2015,N_1568,In_2082);
xor U2016 (N_2016,In_2804,In_1515);
nor U2017 (N_2017,N_1138,N_676);
and U2018 (N_2018,N_1923,N_1694);
nand U2019 (N_2019,N_1606,In_1541);
and U2020 (N_2020,N_1575,N_1528);
xor U2021 (N_2021,N_1913,N_1228);
xnor U2022 (N_2022,N_1954,N_1577);
xnor U2023 (N_2023,N_1026,N_459);
or U2024 (N_2024,N_1790,N_1624);
nor U2025 (N_2025,N_1613,N_1542);
xnor U2026 (N_2026,N_1625,N_1540);
nand U2027 (N_2027,In_1703,N_1052);
and U2028 (N_2028,N_1169,N_1635);
xnor U2029 (N_2029,N_1662,In_2530);
and U2030 (N_2030,N_731,N_208);
or U2031 (N_2031,N_1712,In_164);
xor U2032 (N_2032,In_461,In_640);
xnor U2033 (N_2033,N_1829,N_1942);
nor U2034 (N_2034,N_1551,In_2472);
and U2035 (N_2035,N_1162,N_1653);
nor U2036 (N_2036,N_1992,N_1484);
and U2037 (N_2037,N_1967,N_1326);
nor U2038 (N_2038,N_1964,N_1005);
nor U2039 (N_2039,N_1576,In_2682);
nand U2040 (N_2040,N_1738,N_1985);
xnor U2041 (N_2041,N_1367,N_1604);
and U2042 (N_2042,N_1343,N_214);
xor U2043 (N_2043,N_1341,N_1844);
nor U2044 (N_2044,N_576,In_2158);
or U2045 (N_2045,N_1972,N_1849);
nand U2046 (N_2046,N_1524,In_2681);
or U2047 (N_2047,N_1472,N_1845);
xor U2048 (N_2048,N_1663,In_1779);
and U2049 (N_2049,N_1759,In_2412);
and U2050 (N_2050,N_1616,N_1514);
nand U2051 (N_2051,N_1390,N_506);
nor U2052 (N_2052,N_1999,N_1560);
or U2053 (N_2053,In_2235,N_1386);
and U2054 (N_2054,In_802,N_1987);
xor U2055 (N_2055,N_1148,In_255);
or U2056 (N_2056,N_1714,N_1543);
or U2057 (N_2057,N_1872,N_1513);
or U2058 (N_2058,N_1908,N_1692);
or U2059 (N_2059,N_1903,N_1049);
and U2060 (N_2060,In_848,N_1705);
nor U2061 (N_2061,N_1362,N_1564);
xor U2062 (N_2062,In_1044,N_1403);
nor U2063 (N_2063,In_1041,In_2562);
nand U2064 (N_2064,N_1621,N_1695);
and U2065 (N_2065,N_1417,N_562);
nor U2066 (N_2066,N_1126,N_270);
nor U2067 (N_2067,N_1523,N_1794);
nor U2068 (N_2068,N_1850,In_1954);
xnor U2069 (N_2069,N_1120,N_1701);
or U2070 (N_2070,In_965,In_2440);
and U2071 (N_2071,In_161,N_1634);
nand U2072 (N_2072,N_1186,N_1305);
or U2073 (N_2073,N_1921,N_1937);
xor U2074 (N_2074,N_1072,N_1781);
nand U2075 (N_2075,N_1586,N_1607);
or U2076 (N_2076,N_1032,N_1584);
and U2077 (N_2077,In_237,In_1115);
nand U2078 (N_2078,In_1956,N_1129);
nand U2079 (N_2079,N_1301,N_1966);
xnor U2080 (N_2080,N_1814,In_1733);
and U2081 (N_2081,In_1765,N_1746);
xor U2082 (N_2082,N_1029,N_587);
or U2083 (N_2083,N_1700,N_1857);
nor U2084 (N_2084,N_291,N_583);
and U2085 (N_2085,N_537,N_1884);
nand U2086 (N_2086,N_1727,N_1656);
nand U2087 (N_2087,N_535,N_1650);
nor U2088 (N_2088,N_582,N_1798);
xnor U2089 (N_2089,N_1660,N_1155);
and U2090 (N_2090,N_691,N_1889);
xnor U2091 (N_2091,N_437,N_1862);
xor U2092 (N_2092,N_1793,N_1864);
nor U2093 (N_2093,N_1199,N_1525);
nor U2094 (N_2094,N_1933,N_1991);
or U2095 (N_2095,In_239,N_1792);
and U2096 (N_2096,N_1044,In_339);
and U2097 (N_2097,In_2357,N_1956);
or U2098 (N_2098,N_1208,In_627);
or U2099 (N_2099,N_1785,N_1626);
and U2100 (N_2100,N_1838,N_1632);
nor U2101 (N_2101,In_607,N_1880);
nand U2102 (N_2102,N_1214,N_927);
nand U2103 (N_2103,In_1106,N_1707);
and U2104 (N_2104,N_1552,In_2439);
or U2105 (N_2105,N_1852,In_1359);
or U2106 (N_2106,N_1062,N_1801);
nand U2107 (N_2107,N_1017,N_1627);
nor U2108 (N_2108,N_1846,N_564);
or U2109 (N_2109,N_108,N_1130);
nor U2110 (N_2110,N_1614,In_1721);
or U2111 (N_2111,N_1957,N_1518);
and U2112 (N_2112,N_1891,In_1438);
nor U2113 (N_2113,N_1909,N_1936);
or U2114 (N_2114,N_1597,N_1912);
nor U2115 (N_2115,N_1679,In_801);
and U2116 (N_2116,N_1611,N_649);
nand U2117 (N_2117,N_1766,N_306);
xor U2118 (N_2118,In_1368,N_1521);
nand U2119 (N_2119,In_1465,N_1892);
or U2120 (N_2120,N_1170,N_1860);
xor U2121 (N_2121,N_1863,N_1377);
nand U2122 (N_2122,N_1791,N_1191);
nor U2123 (N_2123,In_1825,N_1439);
nand U2124 (N_2124,N_1303,In_334);
or U2125 (N_2125,N_1928,N_1715);
nand U2126 (N_2126,N_1853,N_1740);
nand U2127 (N_2127,N_1914,N_1610);
or U2128 (N_2128,N_1043,N_1587);
nand U2129 (N_2129,N_1116,N_838);
and U2130 (N_2130,N_1361,N_1934);
xor U2131 (N_2131,N_1767,N_425);
nor U2132 (N_2132,N_110,In_1713);
xor U2133 (N_2133,In_142,N_1578);
xnor U2134 (N_2134,In_2932,N_1416);
xnor U2135 (N_2135,N_1688,N_1869);
nand U2136 (N_2136,N_1734,N_131);
and U2137 (N_2137,N_816,N_1571);
nor U2138 (N_2138,N_1873,N_1511);
nor U2139 (N_2139,N_1063,In_444);
or U2140 (N_2140,N_1486,N_1879);
or U2141 (N_2141,N_879,N_1762);
xnor U2142 (N_2142,N_1948,N_745);
and U2143 (N_2143,N_1951,N_1796);
nor U2144 (N_2144,N_1592,In_1357);
nand U2145 (N_2145,N_716,In_2309);
xor U2146 (N_2146,N_1981,N_1189);
xor U2147 (N_2147,N_1585,N_1681);
xnor U2148 (N_2148,N_1229,N_1628);
nand U2149 (N_2149,N_1902,N_1955);
nand U2150 (N_2150,N_764,N_1093);
and U2151 (N_2151,N_178,In_2801);
or U2152 (N_2152,N_1333,N_1882);
nor U2153 (N_2153,N_1986,N_1218);
xnor U2154 (N_2154,N_1779,In_1766);
nand U2155 (N_2155,N_1615,N_841);
nand U2156 (N_2156,N_1230,In_2463);
nor U2157 (N_2157,N_1601,N_1994);
xnor U2158 (N_2158,N_1566,In_2665);
nand U2159 (N_2159,N_1930,N_581);
nand U2160 (N_2160,N_1878,N_1871);
or U2161 (N_2161,N_1225,N_1988);
nor U2162 (N_2162,N_1803,N_1841);
nand U2163 (N_2163,N_1515,N_1516);
and U2164 (N_2164,N_1327,N_1920);
or U2165 (N_2165,In_2229,In_1008);
nor U2166 (N_2166,N_1168,In_1560);
or U2167 (N_2167,N_1984,N_1919);
or U2168 (N_2168,N_1962,N_1824);
nor U2169 (N_2169,N_1883,N_1298);
nor U2170 (N_2170,N_1353,N_1893);
xnor U2171 (N_2171,In_2653,N_1553);
or U2172 (N_2172,N_337,N_1526);
xor U2173 (N_2173,N_279,N_1639);
or U2174 (N_2174,In_2892,N_1505);
nor U2175 (N_2175,N_1885,N_1683);
nor U2176 (N_2176,N_68,In_1108);
or U2177 (N_2177,N_1581,N_528);
xor U2178 (N_2178,In_1621,N_1406);
xnor U2179 (N_2179,In_2539,N_1753);
xor U2180 (N_2180,In_1591,In_1512);
nand U2181 (N_2181,N_979,N_1881);
nand U2182 (N_2182,N_1527,N_1594);
nand U2183 (N_2183,N_1821,N_1745);
and U2184 (N_2184,In_25,N_1783);
and U2185 (N_2185,N_209,N_1978);
and U2186 (N_2186,N_1777,N_1494);
or U2187 (N_2187,In_459,N_1929);
or U2188 (N_2188,N_1596,N_1865);
and U2189 (N_2189,N_1723,N_507);
or U2190 (N_2190,N_1761,N_722);
nand U2191 (N_2191,N_1812,N_447);
nor U2192 (N_2192,N_1737,N_693);
and U2193 (N_2193,N_1427,N_34);
xnor U2194 (N_2194,In_762,N_1672);
and U2195 (N_2195,N_1870,N_1251);
or U2196 (N_2196,N_851,N_253);
xnor U2197 (N_2197,N_1648,N_1743);
nor U2198 (N_2198,In_478,N_1702);
nand U2199 (N_2199,N_1691,N_1532);
xor U2200 (N_2200,In_2656,N_1720);
or U2201 (N_2201,In_293,N_1795);
nand U2202 (N_2202,N_331,N_1963);
or U2203 (N_2203,N_1926,N_1866);
xor U2204 (N_2204,N_1799,N_1858);
nand U2205 (N_2205,N_516,N_1818);
nand U2206 (N_2206,In_843,N_1947);
nand U2207 (N_2207,In_1946,In_1478);
or U2208 (N_2208,N_1699,N_1041);
and U2209 (N_2209,N_1670,N_87);
and U2210 (N_2210,In_1367,N_1935);
and U2211 (N_2211,N_1851,N_1901);
xnor U2212 (N_2212,In_2148,N_1177);
or U2213 (N_2213,N_1582,N_1907);
nor U2214 (N_2214,In_1611,N_1544);
nor U2215 (N_2215,N_1897,In_1939);
nor U2216 (N_2216,In_2938,In_2313);
nand U2217 (N_2217,N_1925,N_1760);
and U2218 (N_2218,In_1985,In_240);
nor U2219 (N_2219,In_927,N_1731);
nand U2220 (N_2220,N_413,N_1682);
and U2221 (N_2221,N_1244,N_1243);
nand U2222 (N_2222,N_1959,N_966);
xnor U2223 (N_2223,N_295,In_1444);
or U2224 (N_2224,In_1411,N_1977);
and U2225 (N_2225,N_1270,N_1667);
nand U2226 (N_2226,N_1374,N_1674);
nand U2227 (N_2227,N_1471,N_1159);
nor U2228 (N_2228,N_1780,N_1061);
and U2229 (N_2229,N_1729,N_1368);
or U2230 (N_2230,In_2714,N_1822);
xnor U2231 (N_2231,N_1751,N_1278);
nand U2232 (N_2232,N_1952,In_2136);
nand U2233 (N_2233,N_1180,In_754);
nand U2234 (N_2234,N_915,N_1602);
nor U2235 (N_2235,N_1644,N_998);
xnor U2236 (N_2236,N_1539,N_1287);
nand U2237 (N_2237,N_1837,N_1412);
nand U2238 (N_2238,N_1034,N_1160);
nand U2239 (N_2239,N_1742,N_1661);
nand U2240 (N_2240,N_1764,N_1830);
or U2241 (N_2241,N_1756,N_1569);
xnor U2242 (N_2242,N_1512,N_1348);
nor U2243 (N_2243,N_1598,In_1023);
nor U2244 (N_2244,In_2692,N_1433);
and U2245 (N_2245,N_1430,In_922);
nor U2246 (N_2246,N_1982,N_1636);
nor U2247 (N_2247,In_492,N_1689);
nor U2248 (N_2248,In_61,N_1713);
xnor U2249 (N_2249,N_1998,In_80);
xor U2250 (N_2250,N_1530,N_476);
nor U2251 (N_2251,N_1536,N_1283);
and U2252 (N_2252,N_1782,N_203);
nor U2253 (N_2253,N_1426,In_2685);
nand U2254 (N_2254,N_651,N_813);
nand U2255 (N_2255,N_183,N_956);
or U2256 (N_2256,N_1600,N_896);
nand U2257 (N_2257,N_790,N_1547);
xnor U2258 (N_2258,N_1109,N_1546);
nor U2259 (N_2259,N_1996,N_1599);
and U2260 (N_2260,N_1843,N_1918);
nand U2261 (N_2261,N_1995,N_1721);
nor U2262 (N_2262,N_1382,N_1874);
nor U2263 (N_2263,N_171,N_1608);
or U2264 (N_2264,N_1549,N_1205);
and U2265 (N_2265,N_1509,N_1149);
xnor U2266 (N_2266,N_1784,N_520);
nand U2267 (N_2267,N_1410,N_1968);
and U2268 (N_2268,In_384,N_1077);
nor U2269 (N_2269,N_1517,N_1989);
and U2270 (N_2270,In_1660,N_1059);
nor U2271 (N_2271,In_232,N_1917);
and U2272 (N_2272,N_1932,N_1859);
and U2273 (N_2273,N_42,N_1890);
nand U2274 (N_2274,N_1193,N_1797);
xnor U2275 (N_2275,N_831,N_1938);
and U2276 (N_2276,In_2450,N_1207);
xnor U2277 (N_2277,N_1831,In_641);
nor U2278 (N_2278,N_1570,N_1637);
nand U2279 (N_2279,N_1946,N_777);
xnor U2280 (N_2280,In_2231,N_410);
nand U2281 (N_2281,N_1520,N_1216);
and U2282 (N_2282,N_1706,N_1506);
nor U2283 (N_2283,N_826,N_1696);
nor U2284 (N_2284,N_1645,N_1969);
xor U2285 (N_2285,N_1178,N_356);
nand U2286 (N_2286,N_1067,N_1008);
or U2287 (N_2287,In_1132,N_1595);
and U2288 (N_2288,N_1076,In_370);
or U2289 (N_2289,N_1211,N_1114);
or U2290 (N_2290,N_1541,In_399);
or U2291 (N_2291,In_2734,N_1898);
xnor U2292 (N_2292,N_1519,N_1847);
nor U2293 (N_2293,N_735,N_1620);
nand U2294 (N_2294,N_650,N_1693);
nor U2295 (N_2295,In_1361,N_1823);
or U2296 (N_2296,In_653,N_1752);
nor U2297 (N_2297,N_1572,In_2958);
nor U2298 (N_2298,In_1253,N_1819);
nand U2299 (N_2299,In_2624,N_1646);
nor U2300 (N_2300,N_449,N_1345);
xor U2301 (N_2301,N_1711,N_903);
nand U2302 (N_2302,N_1896,N_1253);
nor U2303 (N_2303,N_1744,N_1816);
or U2304 (N_2304,N_1895,N_1045);
nor U2305 (N_2305,N_1778,In_956);
or U2306 (N_2306,N_1500,N_401);
nand U2307 (N_2307,N_697,N_1979);
nor U2308 (N_2308,N_1993,N_1476);
xor U2309 (N_2309,N_1842,N_1504);
or U2310 (N_2310,N_1817,N_1538);
xor U2311 (N_2311,N_1537,N_1976);
nand U2312 (N_2312,In_2112,N_1671);
xor U2313 (N_2313,In_1982,In_2705);
nor U2314 (N_2314,N_464,In_766);
nor U2315 (N_2315,N_1665,In_1194);
or U2316 (N_2316,N_1154,N_1666);
nand U2317 (N_2317,N_441,N_1502);
xor U2318 (N_2318,In_451,N_1379);
and U2319 (N_2319,N_867,N_1380);
or U2320 (N_2320,N_1474,N_1970);
and U2321 (N_2321,N_1118,N_1561);
nand U2322 (N_2322,N_1359,N_1675);
and U2323 (N_2323,N_1834,N_1749);
or U2324 (N_2324,N_1401,In_2376);
xnor U2325 (N_2325,N_885,N_1350);
xnor U2326 (N_2326,N_610,N_1659);
nor U2327 (N_2327,In_219,In_472);
nand U2328 (N_2328,N_931,N_1593);
nand U2329 (N_2329,N_1623,N_1612);
or U2330 (N_2330,N_402,N_1754);
or U2331 (N_2331,N_914,N_1436);
nand U2332 (N_2332,In_392,N_1588);
or U2333 (N_2333,In_2915,In_69);
or U2334 (N_2334,N_1867,N_1293);
and U2335 (N_2335,N_1173,In_1007);
nand U2336 (N_2336,N_1685,N_1415);
or U2337 (N_2337,N_1789,N_1619);
and U2338 (N_2338,N_1658,N_1657);
nor U2339 (N_2339,N_1622,N_416);
and U2340 (N_2340,N_1273,N_1939);
xor U2341 (N_2341,N_1747,N_856);
nor U2342 (N_2342,In_2508,N_1144);
nand U2343 (N_2343,N_1755,N_772);
and U2344 (N_2344,N_1647,N_1054);
and U2345 (N_2345,N_1974,N_301);
and U2346 (N_2346,N_1848,In_1467);
nand U2347 (N_2347,N_1943,N_1809);
nand U2348 (N_2348,In_2616,N_1466);
or U2349 (N_2349,N_1554,N_1342);
or U2350 (N_2350,N_1961,N_860);
nand U2351 (N_2351,N_1836,N_839);
or U2352 (N_2352,N_589,N_1765);
nand U2353 (N_2353,N_1609,N_1802);
and U2354 (N_2354,N_1854,N_1768);
nand U2355 (N_2355,N_1324,In_1929);
or U2356 (N_2356,N_1669,N_1750);
and U2357 (N_2357,N_1736,N_1652);
xnor U2358 (N_2358,N_22,N_1133);
nand U2359 (N_2359,N_1771,In_2517);
nor U2360 (N_2360,In_2394,N_1786);
nand U2361 (N_2361,N_1642,N_1769);
or U2362 (N_2362,In_65,N_1664);
xor U2363 (N_2363,In_2386,N_1284);
and U2364 (N_2364,N_145,N_626);
or U2365 (N_2365,N_1905,N_803);
nand U2366 (N_2366,N_1748,N_1770);
nor U2367 (N_2367,N_1081,N_1567);
nand U2368 (N_2368,In_1812,N_1940);
nand U2369 (N_2369,N_1555,N_1741);
and U2370 (N_2370,In_2197,N_1583);
xnor U2371 (N_2371,N_1291,N_1563);
nand U2372 (N_2372,In_587,N_1557);
xnor U2373 (N_2373,N_1531,N_1617);
nor U2374 (N_2374,N_1900,In_2252);
and U2375 (N_2375,N_1805,In_2462);
and U2376 (N_2376,N_1373,N_1268);
xor U2377 (N_2377,N_1800,In_2596);
nor U2378 (N_2378,In_1442,N_1131);
or U2379 (N_2379,N_1828,N_1709);
or U2380 (N_2380,N_1924,N_1668);
nor U2381 (N_2381,N_991,N_1655);
and U2382 (N_2382,In_1074,N_1888);
and U2383 (N_2383,N_627,N_1868);
or U2384 (N_2384,N_1550,In_1479);
nor U2385 (N_2385,N_1808,In_2799);
xnor U2386 (N_2386,In_1116,N_1510);
or U2387 (N_2387,N_259,In_353);
or U2388 (N_2388,N_470,In_1748);
nor U2389 (N_2389,N_886,N_1916);
or U2390 (N_2390,N_207,N_1710);
nor U2391 (N_2391,N_1176,N_1501);
nor U2392 (N_2392,N_1910,N_1965);
nand U2393 (N_2393,N_1684,N_1589);
nor U2394 (N_2394,N_1507,N_1630);
nand U2395 (N_2395,N_1826,In_1362);
xor U2396 (N_2396,N_1773,N_1906);
or U2397 (N_2397,In_2572,In_1104);
nand U2398 (N_2398,N_521,N_1839);
or U2399 (N_2399,N_1090,In_1247);
xnor U2400 (N_2400,N_1503,N_1163);
xnor U2401 (N_2401,N_1232,In_1847);
xor U2402 (N_2402,N_1931,N_1250);
or U2403 (N_2403,N_1285,N_1558);
or U2404 (N_2404,N_1249,N_768);
and U2405 (N_2405,N_1146,N_1722);
nand U2406 (N_2406,N_1678,N_1070);
xnor U2407 (N_2407,In_107,In_2787);
xor U2408 (N_2408,N_1698,N_73);
nand U2409 (N_2409,N_894,N_1703);
nand U2410 (N_2410,N_1574,In_2324);
nand U2411 (N_2411,N_591,N_1728);
nor U2412 (N_2412,N_1559,N_1562);
or U2413 (N_2413,N_1638,N_1037);
and U2414 (N_2414,N_1680,N_1911);
xnor U2415 (N_2415,N_1774,N_876);
and U2416 (N_2416,N_919,In_1666);
nand U2417 (N_2417,N_1565,N_1522);
and U2418 (N_2418,N_1832,N_1716);
nor U2419 (N_2419,N_1810,N_1649);
or U2420 (N_2420,N_1922,N_1629);
and U2421 (N_2421,N_1338,N_1775);
nand U2422 (N_2422,N_1320,N_1579);
or U2423 (N_2423,N_1446,N_170);
nand U2424 (N_2424,N_1899,N_1633);
or U2425 (N_2425,N_1735,N_1983);
or U2426 (N_2426,N_1804,N_1687);
and U2427 (N_2427,N_1448,N_1813);
and U2428 (N_2428,In_130,N_580);
xor U2429 (N_2429,N_652,In_1338);
and U2430 (N_2430,N_1997,N_1548);
nor U2431 (N_2431,N_709,N_1018);
nor U2432 (N_2432,N_1405,In_1940);
nand U2433 (N_2433,N_1221,In_95);
or U2434 (N_2434,N_1654,N_1256);
and U2435 (N_2435,N_1306,N_1875);
nor U2436 (N_2436,N_1827,In_2052);
nor U2437 (N_2437,N_1973,In_40);
nand U2438 (N_2438,In_1353,N_1053);
nand U2439 (N_2439,N_218,N_1835);
xnor U2440 (N_2440,N_942,N_1605);
nand U2441 (N_2441,In_2676,N_1445);
and U2442 (N_2442,N_1573,N_1958);
nand U2443 (N_2443,N_1980,N_257);
xnor U2444 (N_2444,N_1021,N_607);
xor U2445 (N_2445,N_1174,N_1254);
nand U2446 (N_2446,N_1833,N_1631);
xnor U2447 (N_2447,In_1182,N_1825);
and U2448 (N_2448,N_1590,N_783);
nand U2449 (N_2449,N_1945,In_2329);
or U2450 (N_2450,N_1739,In_724);
nor U2451 (N_2451,N_1529,N_1099);
xnor U2452 (N_2452,N_1725,N_1450);
nor U2453 (N_2453,N_490,In_805);
and U2454 (N_2454,In_2372,N_1718);
and U2455 (N_2455,N_1772,N_1618);
nor U2456 (N_2456,In_2525,N_1673);
or U2457 (N_2457,N_1806,In_1821);
nand U2458 (N_2458,N_776,In_1537);
nand U2459 (N_2459,N_242,N_1452);
nor U2460 (N_2460,In_2622,In_1715);
and U2461 (N_2461,N_1440,N_1134);
xor U2462 (N_2462,N_1887,N_1776);
or U2463 (N_2463,N_1095,N_1533);
nand U2464 (N_2464,In_2873,N_1971);
nor U2465 (N_2465,N_1815,N_1904);
or U2466 (N_2466,N_1358,N_805);
or U2467 (N_2467,N_1719,N_84);
nor U2468 (N_2468,N_1690,N_1677);
or U2469 (N_2469,N_962,N_594);
nand U2470 (N_2470,N_1876,N_1732);
and U2471 (N_2471,N_1641,In_628);
nor U2472 (N_2472,N_1485,N_1643);
nand U2473 (N_2473,In_1407,N_1758);
nand U2474 (N_2474,N_1603,N_1119);
nor U2475 (N_2475,N_1886,In_2312);
nor U2476 (N_2476,N_252,N_1331);
and U2477 (N_2477,N_27,In_460);
and U2478 (N_2478,N_1435,N_1378);
or U2479 (N_2479,N_1108,N_1855);
or U2480 (N_2480,N_575,N_1508);
xor U2481 (N_2481,In_1191,N_1686);
nand U2482 (N_2482,N_1651,In_1045);
xnor U2483 (N_2483,In_210,In_1137);
xnor U2484 (N_2484,N_1556,N_1975);
nor U2485 (N_2485,N_1068,N_901);
or U2486 (N_2486,N_1697,N_1733);
or U2487 (N_2487,N_1877,N_1704);
nor U2488 (N_2488,N_1024,N_1990);
nor U2489 (N_2489,N_1717,N_1545);
and U2490 (N_2490,N_1861,N_1499);
or U2491 (N_2491,N_1950,N_1763);
xor U2492 (N_2492,N_1840,N_1730);
nor U2493 (N_2493,N_1856,N_1820);
or U2494 (N_2494,N_1949,N_1419);
xor U2495 (N_2495,N_1894,N_725);
xnor U2496 (N_2496,In_196,N_1676);
xor U2497 (N_2497,N_1535,N_1172);
or U2498 (N_2498,N_873,N_389);
and U2499 (N_2499,N_597,N_1724);
xnor U2500 (N_2500,N_2147,N_2090);
nand U2501 (N_2501,N_2344,N_2263);
and U2502 (N_2502,N_2370,N_2029);
nor U2503 (N_2503,N_2021,N_2430);
and U2504 (N_2504,N_2374,N_2129);
nand U2505 (N_2505,N_2326,N_2395);
nor U2506 (N_2506,N_2142,N_2163);
xor U2507 (N_2507,N_2382,N_2281);
nand U2508 (N_2508,N_2205,N_2448);
nand U2509 (N_2509,N_2412,N_2099);
and U2510 (N_2510,N_2324,N_2237);
nor U2511 (N_2511,N_2118,N_2075);
nor U2512 (N_2512,N_2091,N_2053);
xnor U2513 (N_2513,N_2188,N_2016);
nand U2514 (N_2514,N_2162,N_2478);
nor U2515 (N_2515,N_2069,N_2458);
nand U2516 (N_2516,N_2042,N_2233);
and U2517 (N_2517,N_2332,N_2336);
and U2518 (N_2518,N_2104,N_2445);
or U2519 (N_2519,N_2339,N_2404);
and U2520 (N_2520,N_2360,N_2413);
xor U2521 (N_2521,N_2290,N_2072);
and U2522 (N_2522,N_2411,N_2298);
or U2523 (N_2523,N_2182,N_2416);
xnor U2524 (N_2524,N_2187,N_2422);
or U2525 (N_2525,N_2451,N_2319);
or U2526 (N_2526,N_2056,N_2432);
and U2527 (N_2527,N_2301,N_2128);
or U2528 (N_2528,N_2452,N_2394);
and U2529 (N_2529,N_2041,N_2171);
and U2530 (N_2530,N_2175,N_2481);
xnor U2531 (N_2531,N_2212,N_2408);
or U2532 (N_2532,N_2185,N_2225);
or U2533 (N_2533,N_2011,N_2073);
nor U2534 (N_2534,N_2294,N_2122);
and U2535 (N_2535,N_2035,N_2059);
and U2536 (N_2536,N_2363,N_2084);
xnor U2537 (N_2537,N_2476,N_2489);
nor U2538 (N_2538,N_2207,N_2247);
nor U2539 (N_2539,N_2031,N_2383);
or U2540 (N_2540,N_2189,N_2334);
and U2541 (N_2541,N_2004,N_2252);
and U2542 (N_2542,N_2295,N_2357);
and U2543 (N_2543,N_2231,N_2077);
or U2544 (N_2544,N_2454,N_2347);
or U2545 (N_2545,N_2353,N_2093);
nand U2546 (N_2546,N_2457,N_2181);
or U2547 (N_2547,N_2495,N_2241);
xnor U2548 (N_2548,N_2268,N_2364);
xor U2549 (N_2549,N_2169,N_2485);
xnor U2550 (N_2550,N_2446,N_2480);
and U2551 (N_2551,N_2190,N_2107);
xor U2552 (N_2552,N_2352,N_2277);
or U2553 (N_2553,N_2322,N_2019);
and U2554 (N_2554,N_2372,N_2100);
xnor U2555 (N_2555,N_2229,N_2381);
or U2556 (N_2556,N_2482,N_2032);
and U2557 (N_2557,N_2111,N_2327);
nor U2558 (N_2558,N_2284,N_2096);
or U2559 (N_2559,N_2170,N_2425);
and U2560 (N_2560,N_2401,N_2282);
xnor U2561 (N_2561,N_2393,N_2191);
and U2562 (N_2562,N_2257,N_2137);
and U2563 (N_2563,N_2442,N_2392);
xnor U2564 (N_2564,N_2160,N_2330);
xor U2565 (N_2565,N_2375,N_2272);
nand U2566 (N_2566,N_2167,N_2245);
xnor U2567 (N_2567,N_2151,N_2119);
xnor U2568 (N_2568,N_2376,N_2496);
xnor U2569 (N_2569,N_2255,N_2467);
nor U2570 (N_2570,N_2251,N_2343);
and U2571 (N_2571,N_2062,N_2434);
nor U2572 (N_2572,N_2331,N_2045);
or U2573 (N_2573,N_2070,N_2354);
nor U2574 (N_2574,N_2057,N_2218);
nand U2575 (N_2575,N_2260,N_2438);
nand U2576 (N_2576,N_2384,N_2391);
nor U2577 (N_2577,N_2450,N_2017);
and U2578 (N_2578,N_2009,N_2397);
nand U2579 (N_2579,N_2387,N_2208);
nor U2580 (N_2580,N_2079,N_2399);
and U2581 (N_2581,N_2407,N_2222);
nor U2582 (N_2582,N_2039,N_2195);
nor U2583 (N_2583,N_2051,N_2465);
nor U2584 (N_2584,N_2010,N_2064);
or U2585 (N_2585,N_2289,N_2377);
xnor U2586 (N_2586,N_2025,N_2293);
and U2587 (N_2587,N_2048,N_2020);
nor U2588 (N_2588,N_2150,N_2477);
nand U2589 (N_2589,N_2429,N_2197);
nand U2590 (N_2590,N_2213,N_2497);
or U2591 (N_2591,N_2177,N_2491);
nand U2592 (N_2592,N_2155,N_2192);
nor U2593 (N_2593,N_2215,N_2082);
nor U2594 (N_2594,N_2203,N_2306);
nor U2595 (N_2595,N_2316,N_2424);
xor U2596 (N_2596,N_2437,N_2464);
or U2597 (N_2597,N_2441,N_2466);
and U2598 (N_2598,N_2012,N_2089);
nor U2599 (N_2599,N_2380,N_2351);
nand U2600 (N_2600,N_2002,N_2078);
or U2601 (N_2601,N_2223,N_2378);
nand U2602 (N_2602,N_2369,N_2499);
nor U2603 (N_2603,N_2270,N_2309);
nand U2604 (N_2604,N_2204,N_2300);
or U2605 (N_2605,N_2148,N_2052);
or U2606 (N_2606,N_2174,N_2217);
and U2607 (N_2607,N_2049,N_2341);
nor U2608 (N_2608,N_2061,N_2068);
xor U2609 (N_2609,N_2456,N_2108);
and U2610 (N_2610,N_2279,N_2101);
nand U2611 (N_2611,N_2013,N_2325);
nor U2612 (N_2612,N_2367,N_2472);
nand U2613 (N_2613,N_2179,N_2135);
nor U2614 (N_2614,N_2033,N_2487);
xor U2615 (N_2615,N_2239,N_2202);
xor U2616 (N_2616,N_2435,N_2304);
nor U2617 (N_2617,N_2386,N_2333);
and U2618 (N_2618,N_2299,N_2498);
or U2619 (N_2619,N_2116,N_2200);
nand U2620 (N_2620,N_2427,N_2243);
nand U2621 (N_2621,N_2242,N_2307);
xnor U2622 (N_2622,N_2198,N_2368);
or U2623 (N_2623,N_2409,N_2153);
xor U2624 (N_2624,N_2066,N_2259);
and U2625 (N_2625,N_2166,N_2356);
or U2626 (N_2626,N_2055,N_2023);
or U2627 (N_2627,N_2085,N_2366);
nor U2628 (N_2628,N_2313,N_2355);
nand U2629 (N_2629,N_2287,N_2373);
or U2630 (N_2630,N_2105,N_2494);
or U2631 (N_2631,N_2314,N_2134);
and U2632 (N_2632,N_2302,N_2214);
and U2633 (N_2633,N_2027,N_2092);
nor U2634 (N_2634,N_2342,N_2337);
and U2635 (N_2635,N_2349,N_2471);
and U2636 (N_2636,N_2156,N_2415);
nand U2637 (N_2637,N_2140,N_2288);
or U2638 (N_2638,N_2071,N_2276);
xor U2639 (N_2639,N_2246,N_2419);
and U2640 (N_2640,N_2262,N_2402);
nor U2641 (N_2641,N_2158,N_2060);
or U2642 (N_2642,N_2463,N_2254);
and U2643 (N_2643,N_2220,N_2462);
nor U2644 (N_2644,N_2256,N_2178);
nand U2645 (N_2645,N_2297,N_2001);
xor U2646 (N_2646,N_2486,N_2273);
and U2647 (N_2647,N_2034,N_2280);
nor U2648 (N_2648,N_2083,N_2038);
or U2649 (N_2649,N_2067,N_2328);
or U2650 (N_2650,N_2120,N_2470);
nand U2651 (N_2651,N_2455,N_2219);
xor U2652 (N_2652,N_2428,N_2453);
xor U2653 (N_2653,N_2121,N_2007);
nand U2654 (N_2654,N_2022,N_2444);
and U2655 (N_2655,N_2232,N_2040);
nor U2656 (N_2656,N_2248,N_2461);
and U2657 (N_2657,N_2000,N_2046);
or U2658 (N_2658,N_2113,N_2026);
nand U2659 (N_2659,N_2224,N_2123);
and U2660 (N_2660,N_2184,N_2440);
xnor U2661 (N_2661,N_2303,N_2348);
xor U2662 (N_2662,N_2350,N_2139);
nor U2663 (N_2663,N_2274,N_2469);
and U2664 (N_2664,N_2358,N_2228);
xnor U2665 (N_2665,N_2087,N_2157);
or U2666 (N_2666,N_2249,N_2389);
xnor U2667 (N_2667,N_2421,N_2005);
xor U2668 (N_2668,N_2238,N_2346);
nor U2669 (N_2669,N_2312,N_2145);
or U2670 (N_2670,N_2400,N_2131);
nor U2671 (N_2671,N_2474,N_2015);
nor U2672 (N_2672,N_2318,N_2194);
nor U2673 (N_2673,N_2164,N_2371);
xor U2674 (N_2674,N_2406,N_2426);
and U2675 (N_2675,N_2475,N_2149);
xnor U2676 (N_2676,N_2112,N_2138);
xnor U2677 (N_2677,N_2144,N_2165);
nand U2678 (N_2678,N_2186,N_2266);
xor U2679 (N_2679,N_2436,N_2168);
nor U2680 (N_2680,N_2240,N_2417);
nor U2681 (N_2681,N_2345,N_2117);
and U2682 (N_2682,N_2127,N_2275);
or U2683 (N_2683,N_2047,N_2114);
nor U2684 (N_2684,N_2076,N_2172);
or U2685 (N_2685,N_2315,N_2103);
xor U2686 (N_2686,N_2283,N_2335);
nand U2687 (N_2687,N_2044,N_2054);
and U2688 (N_2688,N_2431,N_2365);
or U2689 (N_2689,N_2216,N_2320);
and U2690 (N_2690,N_2193,N_2278);
nor U2691 (N_2691,N_2058,N_2080);
nor U2692 (N_2692,N_2115,N_2180);
nand U2693 (N_2693,N_2414,N_2292);
and U2694 (N_2694,N_2008,N_2271);
or U2695 (N_2695,N_2396,N_2449);
or U2696 (N_2696,N_2490,N_2418);
nor U2697 (N_2697,N_2018,N_2003);
xor U2698 (N_2698,N_2261,N_2183);
nor U2699 (N_2699,N_2014,N_2065);
xnor U2700 (N_2700,N_2483,N_2269);
nor U2701 (N_2701,N_2028,N_2385);
and U2702 (N_2702,N_2265,N_2201);
xor U2703 (N_2703,N_2329,N_2405);
nand U2704 (N_2704,N_2338,N_2209);
or U2705 (N_2705,N_2063,N_2102);
and U2706 (N_2706,N_2176,N_2433);
xnor U2707 (N_2707,N_2492,N_2086);
and U2708 (N_2708,N_2484,N_2291);
xor U2709 (N_2709,N_2199,N_2264);
or U2710 (N_2710,N_2479,N_2146);
nor U2711 (N_2711,N_2226,N_2109);
and U2712 (N_2712,N_2141,N_2210);
xnor U2713 (N_2713,N_2493,N_2323);
nor U2714 (N_2714,N_2286,N_2459);
xnor U2715 (N_2715,N_2468,N_2036);
xor U2716 (N_2716,N_2152,N_2081);
nor U2717 (N_2717,N_2143,N_2074);
nor U2718 (N_2718,N_2136,N_2443);
and U2719 (N_2719,N_2124,N_2043);
xor U2720 (N_2720,N_2361,N_2230);
and U2721 (N_2721,N_2030,N_2095);
nor U2722 (N_2722,N_2097,N_2388);
or U2723 (N_2723,N_2420,N_2379);
nand U2724 (N_2724,N_2050,N_2236);
nor U2725 (N_2725,N_2488,N_2285);
nor U2726 (N_2726,N_2296,N_2098);
or U2727 (N_2727,N_2398,N_2258);
and U2728 (N_2728,N_2460,N_2154);
nand U2729 (N_2729,N_2037,N_2310);
nor U2730 (N_2730,N_2110,N_2024);
xor U2731 (N_2731,N_2094,N_2447);
nor U2732 (N_2732,N_2159,N_2410);
and U2733 (N_2733,N_2227,N_2340);
nand U2734 (N_2734,N_2305,N_2423);
nand U2735 (N_2735,N_2267,N_2088);
or U2736 (N_2736,N_2161,N_2403);
nor U2737 (N_2737,N_2253,N_2106);
or U2738 (N_2738,N_2390,N_2126);
or U2739 (N_2739,N_2359,N_2234);
and U2740 (N_2740,N_2321,N_2250);
nand U2741 (N_2741,N_2133,N_2211);
and U2742 (N_2742,N_2132,N_2006);
nand U2743 (N_2743,N_2221,N_2473);
and U2744 (N_2744,N_2439,N_2206);
or U2745 (N_2745,N_2244,N_2235);
or U2746 (N_2746,N_2317,N_2125);
or U2747 (N_2747,N_2196,N_2311);
xor U2748 (N_2748,N_2130,N_2173);
nand U2749 (N_2749,N_2362,N_2308);
nor U2750 (N_2750,N_2479,N_2363);
or U2751 (N_2751,N_2077,N_2320);
xnor U2752 (N_2752,N_2115,N_2234);
or U2753 (N_2753,N_2118,N_2046);
nand U2754 (N_2754,N_2135,N_2114);
nor U2755 (N_2755,N_2466,N_2428);
nand U2756 (N_2756,N_2054,N_2091);
xnor U2757 (N_2757,N_2492,N_2283);
or U2758 (N_2758,N_2036,N_2347);
nor U2759 (N_2759,N_2471,N_2355);
nand U2760 (N_2760,N_2049,N_2013);
or U2761 (N_2761,N_2365,N_2281);
nor U2762 (N_2762,N_2024,N_2474);
xor U2763 (N_2763,N_2071,N_2284);
nand U2764 (N_2764,N_2415,N_2260);
nor U2765 (N_2765,N_2295,N_2482);
xor U2766 (N_2766,N_2093,N_2139);
xnor U2767 (N_2767,N_2225,N_2421);
and U2768 (N_2768,N_2348,N_2438);
and U2769 (N_2769,N_2092,N_2013);
and U2770 (N_2770,N_2006,N_2048);
nor U2771 (N_2771,N_2384,N_2257);
nand U2772 (N_2772,N_2150,N_2103);
or U2773 (N_2773,N_2319,N_2197);
nand U2774 (N_2774,N_2185,N_2378);
xor U2775 (N_2775,N_2175,N_2011);
xnor U2776 (N_2776,N_2320,N_2410);
nand U2777 (N_2777,N_2307,N_2058);
or U2778 (N_2778,N_2110,N_2135);
or U2779 (N_2779,N_2430,N_2072);
and U2780 (N_2780,N_2300,N_2068);
xor U2781 (N_2781,N_2417,N_2112);
nor U2782 (N_2782,N_2166,N_2268);
nor U2783 (N_2783,N_2055,N_2392);
nor U2784 (N_2784,N_2003,N_2352);
and U2785 (N_2785,N_2014,N_2044);
nor U2786 (N_2786,N_2430,N_2038);
nand U2787 (N_2787,N_2279,N_2124);
or U2788 (N_2788,N_2115,N_2239);
or U2789 (N_2789,N_2250,N_2491);
nand U2790 (N_2790,N_2494,N_2355);
xor U2791 (N_2791,N_2094,N_2119);
and U2792 (N_2792,N_2100,N_2313);
nor U2793 (N_2793,N_2168,N_2480);
nor U2794 (N_2794,N_2109,N_2342);
or U2795 (N_2795,N_2466,N_2150);
or U2796 (N_2796,N_2242,N_2222);
and U2797 (N_2797,N_2221,N_2066);
and U2798 (N_2798,N_2338,N_2445);
nor U2799 (N_2799,N_2349,N_2445);
xnor U2800 (N_2800,N_2427,N_2475);
or U2801 (N_2801,N_2385,N_2346);
or U2802 (N_2802,N_2344,N_2371);
and U2803 (N_2803,N_2150,N_2050);
nand U2804 (N_2804,N_2089,N_2126);
or U2805 (N_2805,N_2074,N_2336);
and U2806 (N_2806,N_2396,N_2054);
nor U2807 (N_2807,N_2336,N_2495);
and U2808 (N_2808,N_2404,N_2255);
nor U2809 (N_2809,N_2333,N_2275);
xor U2810 (N_2810,N_2295,N_2050);
nand U2811 (N_2811,N_2080,N_2093);
nor U2812 (N_2812,N_2334,N_2075);
nor U2813 (N_2813,N_2418,N_2491);
and U2814 (N_2814,N_2027,N_2433);
xor U2815 (N_2815,N_2283,N_2300);
or U2816 (N_2816,N_2180,N_2450);
and U2817 (N_2817,N_2485,N_2287);
xnor U2818 (N_2818,N_2084,N_2101);
and U2819 (N_2819,N_2399,N_2021);
or U2820 (N_2820,N_2076,N_2367);
xnor U2821 (N_2821,N_2121,N_2389);
nand U2822 (N_2822,N_2200,N_2462);
and U2823 (N_2823,N_2247,N_2159);
xnor U2824 (N_2824,N_2061,N_2138);
nor U2825 (N_2825,N_2349,N_2347);
and U2826 (N_2826,N_2447,N_2404);
and U2827 (N_2827,N_2349,N_2417);
nand U2828 (N_2828,N_2408,N_2395);
and U2829 (N_2829,N_2353,N_2013);
nor U2830 (N_2830,N_2278,N_2133);
and U2831 (N_2831,N_2041,N_2156);
xor U2832 (N_2832,N_2188,N_2354);
and U2833 (N_2833,N_2197,N_2258);
xor U2834 (N_2834,N_2121,N_2004);
xnor U2835 (N_2835,N_2091,N_2257);
nor U2836 (N_2836,N_2478,N_2380);
nand U2837 (N_2837,N_2076,N_2486);
and U2838 (N_2838,N_2212,N_2304);
and U2839 (N_2839,N_2311,N_2187);
nor U2840 (N_2840,N_2269,N_2359);
xor U2841 (N_2841,N_2343,N_2045);
xnor U2842 (N_2842,N_2010,N_2325);
and U2843 (N_2843,N_2184,N_2006);
and U2844 (N_2844,N_2471,N_2321);
nand U2845 (N_2845,N_2330,N_2331);
and U2846 (N_2846,N_2341,N_2356);
nor U2847 (N_2847,N_2107,N_2413);
xnor U2848 (N_2848,N_2496,N_2018);
nor U2849 (N_2849,N_2465,N_2298);
xor U2850 (N_2850,N_2053,N_2435);
or U2851 (N_2851,N_2163,N_2010);
or U2852 (N_2852,N_2299,N_2296);
xnor U2853 (N_2853,N_2266,N_2406);
and U2854 (N_2854,N_2374,N_2081);
or U2855 (N_2855,N_2316,N_2444);
or U2856 (N_2856,N_2015,N_2184);
nor U2857 (N_2857,N_2059,N_2098);
and U2858 (N_2858,N_2108,N_2420);
nor U2859 (N_2859,N_2424,N_2095);
nor U2860 (N_2860,N_2482,N_2033);
nand U2861 (N_2861,N_2037,N_2164);
nor U2862 (N_2862,N_2319,N_2365);
nand U2863 (N_2863,N_2157,N_2344);
nand U2864 (N_2864,N_2032,N_2019);
or U2865 (N_2865,N_2321,N_2330);
nor U2866 (N_2866,N_2016,N_2228);
nor U2867 (N_2867,N_2028,N_2322);
nand U2868 (N_2868,N_2088,N_2117);
and U2869 (N_2869,N_2360,N_2020);
xor U2870 (N_2870,N_2095,N_2448);
xor U2871 (N_2871,N_2065,N_2206);
nand U2872 (N_2872,N_2308,N_2298);
xnor U2873 (N_2873,N_2082,N_2057);
or U2874 (N_2874,N_2141,N_2268);
nor U2875 (N_2875,N_2263,N_2177);
and U2876 (N_2876,N_2360,N_2493);
nor U2877 (N_2877,N_2450,N_2171);
nor U2878 (N_2878,N_2268,N_2280);
nand U2879 (N_2879,N_2476,N_2149);
or U2880 (N_2880,N_2340,N_2389);
or U2881 (N_2881,N_2368,N_2058);
or U2882 (N_2882,N_2022,N_2236);
or U2883 (N_2883,N_2267,N_2414);
nor U2884 (N_2884,N_2266,N_2047);
nand U2885 (N_2885,N_2256,N_2292);
and U2886 (N_2886,N_2009,N_2019);
or U2887 (N_2887,N_2154,N_2011);
and U2888 (N_2888,N_2139,N_2052);
and U2889 (N_2889,N_2460,N_2199);
nor U2890 (N_2890,N_2288,N_2031);
and U2891 (N_2891,N_2470,N_2158);
nor U2892 (N_2892,N_2310,N_2406);
or U2893 (N_2893,N_2448,N_2329);
and U2894 (N_2894,N_2070,N_2284);
nand U2895 (N_2895,N_2385,N_2343);
and U2896 (N_2896,N_2362,N_2237);
and U2897 (N_2897,N_2149,N_2486);
or U2898 (N_2898,N_2361,N_2161);
nor U2899 (N_2899,N_2249,N_2009);
xor U2900 (N_2900,N_2069,N_2240);
xnor U2901 (N_2901,N_2127,N_2483);
and U2902 (N_2902,N_2177,N_2122);
and U2903 (N_2903,N_2143,N_2140);
nand U2904 (N_2904,N_2166,N_2019);
nand U2905 (N_2905,N_2091,N_2355);
and U2906 (N_2906,N_2380,N_2043);
nor U2907 (N_2907,N_2260,N_2230);
and U2908 (N_2908,N_2217,N_2307);
and U2909 (N_2909,N_2374,N_2261);
xor U2910 (N_2910,N_2002,N_2099);
or U2911 (N_2911,N_2463,N_2444);
and U2912 (N_2912,N_2429,N_2497);
nor U2913 (N_2913,N_2004,N_2402);
nand U2914 (N_2914,N_2067,N_2482);
or U2915 (N_2915,N_2364,N_2360);
nor U2916 (N_2916,N_2104,N_2401);
and U2917 (N_2917,N_2305,N_2397);
or U2918 (N_2918,N_2307,N_2405);
xor U2919 (N_2919,N_2099,N_2125);
or U2920 (N_2920,N_2073,N_2352);
and U2921 (N_2921,N_2250,N_2189);
nand U2922 (N_2922,N_2004,N_2263);
or U2923 (N_2923,N_2045,N_2251);
nor U2924 (N_2924,N_2434,N_2313);
nand U2925 (N_2925,N_2424,N_2161);
and U2926 (N_2926,N_2452,N_2025);
xor U2927 (N_2927,N_2115,N_2285);
or U2928 (N_2928,N_2447,N_2439);
or U2929 (N_2929,N_2168,N_2171);
nand U2930 (N_2930,N_2123,N_2070);
nor U2931 (N_2931,N_2132,N_2230);
and U2932 (N_2932,N_2164,N_2481);
nand U2933 (N_2933,N_2268,N_2498);
and U2934 (N_2934,N_2312,N_2492);
nor U2935 (N_2935,N_2000,N_2319);
nand U2936 (N_2936,N_2279,N_2130);
or U2937 (N_2937,N_2485,N_2403);
and U2938 (N_2938,N_2142,N_2455);
nor U2939 (N_2939,N_2484,N_2354);
nand U2940 (N_2940,N_2459,N_2225);
nand U2941 (N_2941,N_2346,N_2224);
nor U2942 (N_2942,N_2073,N_2228);
xnor U2943 (N_2943,N_2076,N_2111);
or U2944 (N_2944,N_2298,N_2293);
and U2945 (N_2945,N_2489,N_2260);
nor U2946 (N_2946,N_2279,N_2269);
or U2947 (N_2947,N_2239,N_2482);
nor U2948 (N_2948,N_2182,N_2169);
or U2949 (N_2949,N_2355,N_2014);
xnor U2950 (N_2950,N_2050,N_2320);
and U2951 (N_2951,N_2153,N_2090);
or U2952 (N_2952,N_2498,N_2080);
xnor U2953 (N_2953,N_2280,N_2054);
or U2954 (N_2954,N_2248,N_2180);
and U2955 (N_2955,N_2021,N_2414);
or U2956 (N_2956,N_2408,N_2274);
or U2957 (N_2957,N_2494,N_2361);
xnor U2958 (N_2958,N_2242,N_2205);
nand U2959 (N_2959,N_2142,N_2483);
and U2960 (N_2960,N_2241,N_2194);
xnor U2961 (N_2961,N_2495,N_2008);
or U2962 (N_2962,N_2456,N_2297);
xor U2963 (N_2963,N_2057,N_2440);
nor U2964 (N_2964,N_2251,N_2050);
and U2965 (N_2965,N_2231,N_2398);
nor U2966 (N_2966,N_2051,N_2415);
and U2967 (N_2967,N_2341,N_2275);
nor U2968 (N_2968,N_2064,N_2459);
xnor U2969 (N_2969,N_2334,N_2018);
and U2970 (N_2970,N_2304,N_2434);
and U2971 (N_2971,N_2045,N_2032);
and U2972 (N_2972,N_2341,N_2428);
and U2973 (N_2973,N_2306,N_2199);
or U2974 (N_2974,N_2480,N_2221);
nand U2975 (N_2975,N_2438,N_2225);
xnor U2976 (N_2976,N_2417,N_2050);
nor U2977 (N_2977,N_2283,N_2416);
nor U2978 (N_2978,N_2173,N_2387);
or U2979 (N_2979,N_2108,N_2289);
xor U2980 (N_2980,N_2046,N_2175);
xor U2981 (N_2981,N_2292,N_2138);
xor U2982 (N_2982,N_2393,N_2434);
xnor U2983 (N_2983,N_2182,N_2042);
or U2984 (N_2984,N_2365,N_2404);
nor U2985 (N_2985,N_2062,N_2161);
nand U2986 (N_2986,N_2011,N_2220);
xor U2987 (N_2987,N_2306,N_2105);
and U2988 (N_2988,N_2035,N_2024);
and U2989 (N_2989,N_2290,N_2478);
xor U2990 (N_2990,N_2189,N_2024);
or U2991 (N_2991,N_2186,N_2479);
xor U2992 (N_2992,N_2425,N_2437);
nor U2993 (N_2993,N_2433,N_2203);
nor U2994 (N_2994,N_2467,N_2147);
and U2995 (N_2995,N_2305,N_2189);
or U2996 (N_2996,N_2072,N_2460);
nor U2997 (N_2997,N_2292,N_2031);
nor U2998 (N_2998,N_2175,N_2201);
nor U2999 (N_2999,N_2488,N_2333);
nand U3000 (N_3000,N_2598,N_2961);
nand U3001 (N_3001,N_2653,N_2935);
nor U3002 (N_3002,N_2742,N_2983);
and U3003 (N_3003,N_2712,N_2543);
or U3004 (N_3004,N_2876,N_2869);
xor U3005 (N_3005,N_2557,N_2515);
and U3006 (N_3006,N_2868,N_2574);
nor U3007 (N_3007,N_2536,N_2615);
nor U3008 (N_3008,N_2786,N_2747);
or U3009 (N_3009,N_2859,N_2528);
nor U3010 (N_3010,N_2630,N_2668);
or U3011 (N_3011,N_2544,N_2632);
or U3012 (N_3012,N_2828,N_2877);
and U3013 (N_3013,N_2817,N_2784);
xor U3014 (N_3014,N_2753,N_2959);
nor U3015 (N_3015,N_2622,N_2607);
or U3016 (N_3016,N_2778,N_2699);
or U3017 (N_3017,N_2643,N_2863);
nor U3018 (N_3018,N_2678,N_2902);
or U3019 (N_3019,N_2531,N_2822);
nand U3020 (N_3020,N_2954,N_2864);
nor U3021 (N_3021,N_2546,N_2882);
or U3022 (N_3022,N_2586,N_2942);
nand U3023 (N_3023,N_2922,N_2808);
or U3024 (N_3024,N_2693,N_2625);
and U3025 (N_3025,N_2656,N_2760);
nand U3026 (N_3026,N_2949,N_2579);
nand U3027 (N_3027,N_2620,N_2895);
nand U3028 (N_3028,N_2960,N_2969);
nand U3029 (N_3029,N_2683,N_2564);
or U3030 (N_3030,N_2852,N_2988);
nand U3031 (N_3031,N_2737,N_2707);
or U3032 (N_3032,N_2991,N_2793);
xnor U3033 (N_3033,N_2659,N_2724);
xor U3034 (N_3034,N_2601,N_2913);
nand U3035 (N_3035,N_2754,N_2700);
or U3036 (N_3036,N_2533,N_2865);
or U3037 (N_3037,N_2795,N_2931);
xnor U3038 (N_3038,N_2611,N_2788);
nand U3039 (N_3039,N_2676,N_2987);
nor U3040 (N_3040,N_2705,N_2534);
and U3041 (N_3041,N_2673,N_2513);
or U3042 (N_3042,N_2777,N_2981);
nand U3043 (N_3043,N_2592,N_2989);
nand U3044 (N_3044,N_2571,N_2684);
and U3045 (N_3045,N_2792,N_2558);
nand U3046 (N_3046,N_2925,N_2519);
and U3047 (N_3047,N_2875,N_2905);
and U3048 (N_3048,N_2727,N_2530);
and U3049 (N_3049,N_2901,N_2870);
nor U3050 (N_3050,N_2797,N_2888);
and U3051 (N_3051,N_2702,N_2701);
nor U3052 (N_3052,N_2810,N_2597);
and U3053 (N_3053,N_2749,N_2994);
nand U3054 (N_3054,N_2892,N_2851);
xnor U3055 (N_3055,N_2578,N_2997);
or U3056 (N_3056,N_2722,N_2860);
and U3057 (N_3057,N_2841,N_2614);
nor U3058 (N_3058,N_2899,N_2772);
nor U3059 (N_3059,N_2524,N_2569);
and U3060 (N_3060,N_2921,N_2617);
nand U3061 (N_3061,N_2561,N_2646);
nand U3062 (N_3062,N_2638,N_2733);
nand U3063 (N_3063,N_2674,N_2773);
xor U3064 (N_3064,N_2685,N_2896);
or U3065 (N_3065,N_2590,N_2890);
or U3066 (N_3066,N_2956,N_2919);
or U3067 (N_3067,N_2984,N_2781);
nor U3068 (N_3068,N_2583,N_2679);
nor U3069 (N_3069,N_2556,N_2605);
nor U3070 (N_3070,N_2770,N_2929);
xnor U3071 (N_3071,N_2974,N_2540);
or U3072 (N_3072,N_2985,N_2884);
xor U3073 (N_3073,N_2553,N_2924);
nor U3074 (N_3074,N_2835,N_2972);
xnor U3075 (N_3075,N_2849,N_2789);
xnor U3076 (N_3076,N_2559,N_2500);
nor U3077 (N_3077,N_2631,N_2833);
xor U3078 (N_3078,N_2726,N_2745);
and U3079 (N_3079,N_2514,N_2594);
nor U3080 (N_3080,N_2599,N_2937);
or U3081 (N_3081,N_2776,N_2591);
nor U3082 (N_3082,N_2541,N_2746);
or U3083 (N_3083,N_2838,N_2672);
xor U3084 (N_3084,N_2669,N_2651);
nor U3085 (N_3085,N_2775,N_2680);
and U3086 (N_3086,N_2977,N_2823);
and U3087 (N_3087,N_2648,N_2866);
and U3088 (N_3088,N_2986,N_2610);
nand U3089 (N_3089,N_2714,N_2719);
xnor U3090 (N_3090,N_2799,N_2640);
and U3091 (N_3091,N_2549,N_2535);
nand U3092 (N_3092,N_2511,N_2764);
nand U3093 (N_3093,N_2883,N_2744);
and U3094 (N_3094,N_2768,N_2711);
xor U3095 (N_3095,N_2522,N_2873);
and U3096 (N_3096,N_2872,N_2509);
nand U3097 (N_3097,N_2967,N_2940);
or U3098 (N_3098,N_2527,N_2554);
and U3099 (N_3099,N_2609,N_2505);
or U3100 (N_3100,N_2769,N_2743);
nor U3101 (N_3101,N_2600,N_2552);
xor U3102 (N_3102,N_2918,N_2785);
nor U3103 (N_3103,N_2565,N_2794);
or U3104 (N_3104,N_2846,N_2758);
nand U3105 (N_3105,N_2624,N_2867);
nand U3106 (N_3106,N_2703,N_2734);
nand U3107 (N_3107,N_2504,N_2616);
nor U3108 (N_3108,N_2850,N_2572);
nand U3109 (N_3109,N_2621,N_2965);
or U3110 (N_3110,N_2887,N_2862);
and U3111 (N_3111,N_2802,N_2812);
xor U3112 (N_3112,N_2608,N_2821);
xor U3113 (N_3113,N_2635,N_2805);
nand U3114 (N_3114,N_2825,N_2577);
nor U3115 (N_3115,N_2933,N_2520);
nor U3116 (N_3116,N_2654,N_2813);
nor U3117 (N_3117,N_2928,N_2881);
xor U3118 (N_3118,N_2762,N_2824);
nand U3119 (N_3119,N_2976,N_2633);
and U3120 (N_3120,N_2717,N_2998);
nand U3121 (N_3121,N_2735,N_2508);
and U3122 (N_3122,N_2946,N_2613);
and U3123 (N_3123,N_2593,N_2783);
nor U3124 (N_3124,N_2964,N_2510);
nand U3125 (N_3125,N_2966,N_2950);
nand U3126 (N_3126,N_2765,N_2767);
or U3127 (N_3127,N_2807,N_2641);
or U3128 (N_3128,N_2944,N_2791);
nor U3129 (N_3129,N_2800,N_2912);
xor U3130 (N_3130,N_2993,N_2885);
and U3131 (N_3131,N_2708,N_2897);
xor U3132 (N_3132,N_2771,N_2819);
or U3133 (N_3133,N_2827,N_2661);
nand U3134 (N_3134,N_2687,N_2682);
xor U3135 (N_3135,N_2501,N_2843);
nand U3136 (N_3136,N_2506,N_2982);
and U3137 (N_3137,N_2575,N_2739);
or U3138 (N_3138,N_2740,N_2858);
nand U3139 (N_3139,N_2750,N_2731);
nand U3140 (N_3140,N_2650,N_2644);
xnor U3141 (N_3141,N_2526,N_2704);
and U3142 (N_3142,N_2798,N_2955);
or U3143 (N_3143,N_2716,N_2803);
nor U3144 (N_3144,N_2652,N_2539);
or U3145 (N_3145,N_2932,N_2698);
nor U3146 (N_3146,N_2715,N_2952);
xor U3147 (N_3147,N_2507,N_2962);
xor U3148 (N_3148,N_2879,N_2634);
xnor U3149 (N_3149,N_2830,N_2662);
nor U3150 (N_3150,N_2926,N_2755);
or U3151 (N_3151,N_2796,N_2681);
xor U3152 (N_3152,N_2857,N_2971);
nor U3153 (N_3153,N_2930,N_2990);
xnor U3154 (N_3154,N_2752,N_2667);
nor U3155 (N_3155,N_2915,N_2645);
and U3156 (N_3156,N_2815,N_2898);
and U3157 (N_3157,N_2904,N_2502);
xor U3158 (N_3158,N_2589,N_2709);
nor U3159 (N_3159,N_2580,N_2670);
xnor U3160 (N_3160,N_2936,N_2671);
or U3161 (N_3161,N_2560,N_2854);
nand U3162 (N_3162,N_2837,N_2663);
nor U3163 (N_3163,N_2562,N_2893);
or U3164 (N_3164,N_2545,N_2910);
and U3165 (N_3165,N_2538,N_2780);
xnor U3166 (N_3166,N_2706,N_2878);
or U3167 (N_3167,N_2525,N_2532);
xor U3168 (N_3168,N_2958,N_2801);
xor U3169 (N_3169,N_2871,N_2839);
xor U3170 (N_3170,N_2551,N_2957);
or U3171 (N_3171,N_2806,N_2820);
or U3172 (N_3172,N_2665,N_2563);
xnor U3173 (N_3173,N_2874,N_2555);
nand U3174 (N_3174,N_2941,N_2523);
nand U3175 (N_3175,N_2736,N_2710);
or U3176 (N_3176,N_2690,N_2729);
xnor U3177 (N_3177,N_2720,N_2548);
and U3178 (N_3178,N_2880,N_2618);
xnor U3179 (N_3179,N_2891,N_2804);
nor U3180 (N_3180,N_2923,N_2861);
xnor U3181 (N_3181,N_2547,N_2660);
and U3182 (N_3182,N_2761,N_2999);
or U3183 (N_3183,N_2938,N_2516);
nand U3184 (N_3184,N_2748,N_2853);
xnor U3185 (N_3185,N_2756,N_2686);
and U3186 (N_3186,N_2939,N_2816);
or U3187 (N_3187,N_2629,N_2732);
and U3188 (N_3188,N_2550,N_2963);
nor U3189 (N_3189,N_2596,N_2692);
or U3190 (N_3190,N_2948,N_2741);
nand U3191 (N_3191,N_2995,N_2666);
and U3192 (N_3192,N_2811,N_2582);
xor U3193 (N_3193,N_2738,N_2832);
xnor U3194 (N_3194,N_2657,N_2602);
nand U3195 (N_3195,N_2836,N_2623);
or U3196 (N_3196,N_2980,N_2908);
nor U3197 (N_3197,N_2818,N_2920);
or U3198 (N_3198,N_2675,N_2581);
xnor U3199 (N_3199,N_2697,N_2518);
nor U3200 (N_3200,N_2992,N_2691);
nand U3201 (N_3201,N_2721,N_2834);
and U3202 (N_3202,N_2537,N_2689);
or U3203 (N_3203,N_2521,N_2636);
nor U3204 (N_3204,N_2576,N_2566);
xnor U3205 (N_3205,N_2759,N_2573);
nor U3206 (N_3206,N_2570,N_2723);
nor U3207 (N_3207,N_2647,N_2695);
or U3208 (N_3208,N_2911,N_2628);
or U3209 (N_3209,N_2848,N_2917);
and U3210 (N_3210,N_2655,N_2943);
and U3211 (N_3211,N_2763,N_2728);
xor U3212 (N_3212,N_2642,N_2725);
nand U3213 (N_3213,N_2847,N_2782);
xor U3214 (N_3214,N_2585,N_2677);
or U3215 (N_3215,N_2975,N_2664);
xnor U3216 (N_3216,N_2909,N_2814);
or U3217 (N_3217,N_2637,N_2934);
nand U3218 (N_3218,N_2840,N_2588);
nor U3219 (N_3219,N_2603,N_2757);
xor U3220 (N_3220,N_2903,N_2996);
or U3221 (N_3221,N_2945,N_2713);
or U3222 (N_3222,N_2889,N_2856);
nor U3223 (N_3223,N_2831,N_2826);
or U3224 (N_3224,N_2906,N_2694);
nor U3225 (N_3225,N_2787,N_2529);
xnor U3226 (N_3226,N_2696,N_2970);
or U3227 (N_3227,N_2914,N_2730);
nor U3228 (N_3228,N_2842,N_2844);
and U3229 (N_3229,N_2790,N_2751);
nand U3230 (N_3230,N_2953,N_2626);
or U3231 (N_3231,N_2774,N_2894);
nor U3232 (N_3232,N_2649,N_2916);
nand U3233 (N_3233,N_2907,N_2612);
xor U3234 (N_3234,N_2779,N_2627);
nor U3235 (N_3235,N_2829,N_2639);
nand U3236 (N_3236,N_2584,N_2568);
and U3237 (N_3237,N_2718,N_2809);
xnor U3238 (N_3238,N_2979,N_2512);
nand U3239 (N_3239,N_2503,N_2595);
or U3240 (N_3240,N_2688,N_2845);
xor U3241 (N_3241,N_2766,N_2947);
and U3242 (N_3242,N_2973,N_2587);
xnor U3243 (N_3243,N_2567,N_2978);
nand U3244 (N_3244,N_2606,N_2658);
and U3245 (N_3245,N_2886,N_2951);
and U3246 (N_3246,N_2855,N_2900);
xnor U3247 (N_3247,N_2927,N_2619);
and U3248 (N_3248,N_2604,N_2968);
and U3249 (N_3249,N_2517,N_2542);
nor U3250 (N_3250,N_2838,N_2669);
and U3251 (N_3251,N_2975,N_2876);
nor U3252 (N_3252,N_2635,N_2588);
or U3253 (N_3253,N_2802,N_2725);
xnor U3254 (N_3254,N_2730,N_2540);
and U3255 (N_3255,N_2679,N_2936);
nand U3256 (N_3256,N_2701,N_2974);
nor U3257 (N_3257,N_2652,N_2972);
and U3258 (N_3258,N_2904,N_2671);
nor U3259 (N_3259,N_2814,N_2978);
or U3260 (N_3260,N_2803,N_2737);
and U3261 (N_3261,N_2874,N_2780);
or U3262 (N_3262,N_2889,N_2747);
nand U3263 (N_3263,N_2692,N_2706);
nor U3264 (N_3264,N_2904,N_2544);
or U3265 (N_3265,N_2759,N_2815);
nor U3266 (N_3266,N_2744,N_2569);
or U3267 (N_3267,N_2963,N_2889);
or U3268 (N_3268,N_2814,N_2740);
nand U3269 (N_3269,N_2686,N_2613);
or U3270 (N_3270,N_2783,N_2966);
or U3271 (N_3271,N_2797,N_2523);
and U3272 (N_3272,N_2872,N_2778);
xor U3273 (N_3273,N_2598,N_2773);
xor U3274 (N_3274,N_2880,N_2651);
nand U3275 (N_3275,N_2810,N_2819);
xnor U3276 (N_3276,N_2517,N_2900);
nand U3277 (N_3277,N_2983,N_2781);
or U3278 (N_3278,N_2879,N_2843);
or U3279 (N_3279,N_2921,N_2586);
and U3280 (N_3280,N_2771,N_2582);
xor U3281 (N_3281,N_2774,N_2576);
or U3282 (N_3282,N_2707,N_2958);
xor U3283 (N_3283,N_2917,N_2911);
nor U3284 (N_3284,N_2533,N_2695);
or U3285 (N_3285,N_2634,N_2796);
nand U3286 (N_3286,N_2831,N_2793);
xor U3287 (N_3287,N_2665,N_2741);
nand U3288 (N_3288,N_2757,N_2805);
xor U3289 (N_3289,N_2784,N_2581);
nand U3290 (N_3290,N_2807,N_2722);
nand U3291 (N_3291,N_2897,N_2628);
or U3292 (N_3292,N_2753,N_2783);
and U3293 (N_3293,N_2602,N_2579);
or U3294 (N_3294,N_2950,N_2662);
nand U3295 (N_3295,N_2999,N_2785);
nand U3296 (N_3296,N_2595,N_2801);
xnor U3297 (N_3297,N_2613,N_2675);
nand U3298 (N_3298,N_2959,N_2535);
or U3299 (N_3299,N_2999,N_2967);
or U3300 (N_3300,N_2582,N_2777);
xor U3301 (N_3301,N_2602,N_2791);
nand U3302 (N_3302,N_2573,N_2558);
nor U3303 (N_3303,N_2970,N_2962);
nor U3304 (N_3304,N_2671,N_2952);
or U3305 (N_3305,N_2511,N_2593);
and U3306 (N_3306,N_2851,N_2753);
nor U3307 (N_3307,N_2659,N_2746);
and U3308 (N_3308,N_2652,N_2631);
nand U3309 (N_3309,N_2561,N_2514);
nand U3310 (N_3310,N_2558,N_2863);
nor U3311 (N_3311,N_2540,N_2780);
or U3312 (N_3312,N_2549,N_2899);
nand U3313 (N_3313,N_2845,N_2903);
nor U3314 (N_3314,N_2744,N_2779);
xor U3315 (N_3315,N_2589,N_2597);
nor U3316 (N_3316,N_2514,N_2965);
xor U3317 (N_3317,N_2944,N_2972);
xnor U3318 (N_3318,N_2716,N_2871);
or U3319 (N_3319,N_2893,N_2537);
nand U3320 (N_3320,N_2731,N_2940);
nor U3321 (N_3321,N_2781,N_2613);
or U3322 (N_3322,N_2803,N_2605);
nand U3323 (N_3323,N_2935,N_2995);
nor U3324 (N_3324,N_2508,N_2776);
or U3325 (N_3325,N_2989,N_2871);
and U3326 (N_3326,N_2515,N_2671);
or U3327 (N_3327,N_2766,N_2592);
xor U3328 (N_3328,N_2964,N_2987);
and U3329 (N_3329,N_2795,N_2970);
xor U3330 (N_3330,N_2764,N_2913);
or U3331 (N_3331,N_2925,N_2809);
or U3332 (N_3332,N_2822,N_2824);
nor U3333 (N_3333,N_2871,N_2967);
nand U3334 (N_3334,N_2887,N_2618);
nor U3335 (N_3335,N_2520,N_2723);
nor U3336 (N_3336,N_2629,N_2806);
and U3337 (N_3337,N_2700,N_2871);
nor U3338 (N_3338,N_2693,N_2576);
nand U3339 (N_3339,N_2767,N_2676);
xor U3340 (N_3340,N_2978,N_2779);
nor U3341 (N_3341,N_2509,N_2969);
nor U3342 (N_3342,N_2893,N_2722);
nor U3343 (N_3343,N_2784,N_2993);
xor U3344 (N_3344,N_2603,N_2722);
xnor U3345 (N_3345,N_2827,N_2636);
or U3346 (N_3346,N_2644,N_2676);
and U3347 (N_3347,N_2670,N_2798);
nand U3348 (N_3348,N_2931,N_2696);
nor U3349 (N_3349,N_2841,N_2793);
nand U3350 (N_3350,N_2848,N_2795);
nor U3351 (N_3351,N_2745,N_2525);
nor U3352 (N_3352,N_2908,N_2719);
and U3353 (N_3353,N_2965,N_2750);
nand U3354 (N_3354,N_2822,N_2722);
and U3355 (N_3355,N_2549,N_2511);
nand U3356 (N_3356,N_2699,N_2753);
xor U3357 (N_3357,N_2612,N_2867);
xnor U3358 (N_3358,N_2622,N_2754);
nand U3359 (N_3359,N_2927,N_2854);
nand U3360 (N_3360,N_2820,N_2800);
nor U3361 (N_3361,N_2739,N_2933);
xnor U3362 (N_3362,N_2500,N_2516);
nand U3363 (N_3363,N_2737,N_2939);
and U3364 (N_3364,N_2621,N_2792);
xor U3365 (N_3365,N_2510,N_2858);
nand U3366 (N_3366,N_2525,N_2713);
or U3367 (N_3367,N_2729,N_2816);
xor U3368 (N_3368,N_2507,N_2800);
and U3369 (N_3369,N_2563,N_2548);
nand U3370 (N_3370,N_2715,N_2683);
and U3371 (N_3371,N_2598,N_2915);
and U3372 (N_3372,N_2992,N_2788);
or U3373 (N_3373,N_2795,N_2693);
xnor U3374 (N_3374,N_2953,N_2721);
and U3375 (N_3375,N_2580,N_2989);
nand U3376 (N_3376,N_2629,N_2893);
or U3377 (N_3377,N_2548,N_2800);
or U3378 (N_3378,N_2649,N_2565);
nor U3379 (N_3379,N_2853,N_2730);
nor U3380 (N_3380,N_2818,N_2597);
or U3381 (N_3381,N_2621,N_2735);
nor U3382 (N_3382,N_2599,N_2891);
nor U3383 (N_3383,N_2653,N_2529);
and U3384 (N_3384,N_2635,N_2867);
nor U3385 (N_3385,N_2711,N_2804);
nor U3386 (N_3386,N_2932,N_2586);
xnor U3387 (N_3387,N_2986,N_2602);
nand U3388 (N_3388,N_2560,N_2617);
or U3389 (N_3389,N_2730,N_2944);
nor U3390 (N_3390,N_2545,N_2513);
xnor U3391 (N_3391,N_2678,N_2763);
xor U3392 (N_3392,N_2522,N_2694);
or U3393 (N_3393,N_2835,N_2624);
or U3394 (N_3394,N_2735,N_2967);
and U3395 (N_3395,N_2575,N_2920);
xor U3396 (N_3396,N_2804,N_2524);
xor U3397 (N_3397,N_2923,N_2991);
nor U3398 (N_3398,N_2875,N_2701);
and U3399 (N_3399,N_2816,N_2789);
xnor U3400 (N_3400,N_2537,N_2956);
xor U3401 (N_3401,N_2644,N_2570);
xnor U3402 (N_3402,N_2512,N_2796);
and U3403 (N_3403,N_2769,N_2500);
xnor U3404 (N_3404,N_2878,N_2948);
nor U3405 (N_3405,N_2573,N_2738);
nand U3406 (N_3406,N_2566,N_2649);
nand U3407 (N_3407,N_2508,N_2694);
or U3408 (N_3408,N_2887,N_2821);
or U3409 (N_3409,N_2554,N_2692);
and U3410 (N_3410,N_2500,N_2570);
or U3411 (N_3411,N_2917,N_2541);
nand U3412 (N_3412,N_2775,N_2617);
xor U3413 (N_3413,N_2897,N_2792);
or U3414 (N_3414,N_2836,N_2653);
and U3415 (N_3415,N_2751,N_2868);
nand U3416 (N_3416,N_2696,N_2730);
and U3417 (N_3417,N_2688,N_2707);
xor U3418 (N_3418,N_2934,N_2833);
nand U3419 (N_3419,N_2913,N_2777);
or U3420 (N_3420,N_2963,N_2897);
or U3421 (N_3421,N_2918,N_2804);
and U3422 (N_3422,N_2588,N_2561);
xor U3423 (N_3423,N_2609,N_2674);
nand U3424 (N_3424,N_2649,N_2783);
or U3425 (N_3425,N_2700,N_2899);
xnor U3426 (N_3426,N_2758,N_2871);
and U3427 (N_3427,N_2870,N_2748);
or U3428 (N_3428,N_2992,N_2804);
xor U3429 (N_3429,N_2632,N_2840);
and U3430 (N_3430,N_2556,N_2553);
nand U3431 (N_3431,N_2792,N_2847);
nor U3432 (N_3432,N_2607,N_2515);
nor U3433 (N_3433,N_2686,N_2517);
and U3434 (N_3434,N_2758,N_2836);
nand U3435 (N_3435,N_2794,N_2613);
xnor U3436 (N_3436,N_2530,N_2562);
nand U3437 (N_3437,N_2764,N_2688);
nand U3438 (N_3438,N_2559,N_2615);
and U3439 (N_3439,N_2752,N_2956);
nand U3440 (N_3440,N_2803,N_2646);
and U3441 (N_3441,N_2829,N_2522);
and U3442 (N_3442,N_2996,N_2832);
xnor U3443 (N_3443,N_2554,N_2714);
nor U3444 (N_3444,N_2600,N_2690);
or U3445 (N_3445,N_2621,N_2513);
nor U3446 (N_3446,N_2501,N_2520);
nand U3447 (N_3447,N_2840,N_2920);
nor U3448 (N_3448,N_2621,N_2730);
xnor U3449 (N_3449,N_2719,N_2815);
xnor U3450 (N_3450,N_2708,N_2770);
or U3451 (N_3451,N_2942,N_2615);
and U3452 (N_3452,N_2773,N_2896);
nor U3453 (N_3453,N_2671,N_2557);
nor U3454 (N_3454,N_2533,N_2540);
or U3455 (N_3455,N_2873,N_2506);
nor U3456 (N_3456,N_2767,N_2973);
nor U3457 (N_3457,N_2705,N_2523);
and U3458 (N_3458,N_2572,N_2939);
and U3459 (N_3459,N_2823,N_2784);
nor U3460 (N_3460,N_2781,N_2609);
xnor U3461 (N_3461,N_2620,N_2654);
xnor U3462 (N_3462,N_2839,N_2520);
nand U3463 (N_3463,N_2714,N_2747);
nor U3464 (N_3464,N_2944,N_2507);
nor U3465 (N_3465,N_2500,N_2755);
nand U3466 (N_3466,N_2831,N_2923);
nor U3467 (N_3467,N_2985,N_2628);
xnor U3468 (N_3468,N_2504,N_2817);
and U3469 (N_3469,N_2735,N_2647);
nor U3470 (N_3470,N_2638,N_2979);
and U3471 (N_3471,N_2874,N_2730);
and U3472 (N_3472,N_2614,N_2737);
nand U3473 (N_3473,N_2504,N_2939);
xnor U3474 (N_3474,N_2949,N_2569);
nor U3475 (N_3475,N_2761,N_2922);
nor U3476 (N_3476,N_2610,N_2835);
and U3477 (N_3477,N_2598,N_2819);
nor U3478 (N_3478,N_2785,N_2571);
and U3479 (N_3479,N_2885,N_2577);
nor U3480 (N_3480,N_2741,N_2977);
nand U3481 (N_3481,N_2989,N_2646);
and U3482 (N_3482,N_2906,N_2947);
xnor U3483 (N_3483,N_2813,N_2609);
nand U3484 (N_3484,N_2819,N_2792);
or U3485 (N_3485,N_2778,N_2785);
and U3486 (N_3486,N_2931,N_2845);
nand U3487 (N_3487,N_2942,N_2594);
nand U3488 (N_3488,N_2727,N_2684);
xnor U3489 (N_3489,N_2766,N_2659);
or U3490 (N_3490,N_2942,N_2698);
xor U3491 (N_3491,N_2601,N_2974);
or U3492 (N_3492,N_2815,N_2624);
nor U3493 (N_3493,N_2916,N_2612);
nand U3494 (N_3494,N_2620,N_2761);
xnor U3495 (N_3495,N_2930,N_2881);
nand U3496 (N_3496,N_2707,N_2723);
nand U3497 (N_3497,N_2941,N_2559);
or U3498 (N_3498,N_2693,N_2700);
or U3499 (N_3499,N_2733,N_2870);
or U3500 (N_3500,N_3234,N_3299);
nand U3501 (N_3501,N_3454,N_3209);
xnor U3502 (N_3502,N_3248,N_3144);
nor U3503 (N_3503,N_3380,N_3170);
nor U3504 (N_3504,N_3354,N_3168);
nand U3505 (N_3505,N_3003,N_3439);
xnor U3506 (N_3506,N_3072,N_3115);
nand U3507 (N_3507,N_3479,N_3236);
nand U3508 (N_3508,N_3239,N_3330);
nor U3509 (N_3509,N_3445,N_3455);
and U3510 (N_3510,N_3240,N_3040);
or U3511 (N_3511,N_3220,N_3147);
or U3512 (N_3512,N_3148,N_3250);
nand U3513 (N_3513,N_3276,N_3070);
or U3514 (N_3514,N_3389,N_3368);
or U3515 (N_3515,N_3223,N_3405);
xnor U3516 (N_3516,N_3030,N_3121);
and U3517 (N_3517,N_3136,N_3300);
nor U3518 (N_3518,N_3202,N_3359);
nor U3519 (N_3519,N_3082,N_3016);
nand U3520 (N_3520,N_3397,N_3160);
xnor U3521 (N_3521,N_3139,N_3018);
xnor U3522 (N_3522,N_3000,N_3080);
or U3523 (N_3523,N_3289,N_3425);
and U3524 (N_3524,N_3279,N_3015);
xor U3525 (N_3525,N_3198,N_3317);
nor U3526 (N_3526,N_3367,N_3177);
and U3527 (N_3527,N_3378,N_3322);
nor U3528 (N_3528,N_3131,N_3460);
and U3529 (N_3529,N_3435,N_3247);
nand U3530 (N_3530,N_3415,N_3403);
or U3531 (N_3531,N_3012,N_3058);
and U3532 (N_3532,N_3320,N_3426);
xnor U3533 (N_3533,N_3241,N_3112);
nor U3534 (N_3534,N_3061,N_3088);
and U3535 (N_3535,N_3008,N_3039);
nor U3536 (N_3536,N_3482,N_3258);
xor U3537 (N_3537,N_3163,N_3001);
and U3538 (N_3538,N_3078,N_3379);
xnor U3539 (N_3539,N_3085,N_3382);
and U3540 (N_3540,N_3164,N_3023);
nand U3541 (N_3541,N_3461,N_3295);
nor U3542 (N_3542,N_3208,N_3325);
or U3543 (N_3543,N_3283,N_3494);
and U3544 (N_3544,N_3087,N_3476);
or U3545 (N_3545,N_3235,N_3022);
nor U3546 (N_3546,N_3029,N_3488);
nor U3547 (N_3547,N_3233,N_3173);
xnor U3548 (N_3548,N_3057,N_3268);
and U3549 (N_3549,N_3069,N_3485);
nor U3550 (N_3550,N_3178,N_3211);
nand U3551 (N_3551,N_3338,N_3358);
xor U3552 (N_3552,N_3365,N_3033);
xor U3553 (N_3553,N_3274,N_3370);
nand U3554 (N_3554,N_3327,N_3360);
and U3555 (N_3555,N_3324,N_3210);
or U3556 (N_3556,N_3434,N_3282);
or U3557 (N_3557,N_3315,N_3407);
or U3558 (N_3558,N_3344,N_3459);
nor U3559 (N_3559,N_3103,N_3026);
nor U3560 (N_3560,N_3073,N_3064);
or U3561 (N_3561,N_3138,N_3270);
and U3562 (N_3562,N_3277,N_3404);
nand U3563 (N_3563,N_3393,N_3371);
nand U3564 (N_3564,N_3127,N_3132);
and U3565 (N_3565,N_3025,N_3428);
or U3566 (N_3566,N_3134,N_3284);
nor U3567 (N_3567,N_3414,N_3312);
xnor U3568 (N_3568,N_3395,N_3199);
and U3569 (N_3569,N_3364,N_3205);
or U3570 (N_3570,N_3419,N_3224);
nand U3571 (N_3571,N_3060,N_3158);
xnor U3572 (N_3572,N_3383,N_3099);
nor U3573 (N_3573,N_3049,N_3129);
and U3574 (N_3574,N_3465,N_3418);
xor U3575 (N_3575,N_3185,N_3417);
xor U3576 (N_3576,N_3413,N_3478);
or U3577 (N_3577,N_3167,N_3111);
nand U3578 (N_3578,N_3204,N_3334);
or U3579 (N_3579,N_3498,N_3273);
nor U3580 (N_3580,N_3318,N_3114);
nor U3581 (N_3581,N_3411,N_3155);
and U3582 (N_3582,N_3310,N_3089);
nor U3583 (N_3583,N_3497,N_3021);
nor U3584 (N_3584,N_3095,N_3302);
xor U3585 (N_3585,N_3451,N_3120);
or U3586 (N_3586,N_3468,N_3253);
nor U3587 (N_3587,N_3492,N_3188);
xor U3588 (N_3588,N_3339,N_3162);
or U3589 (N_3589,N_3385,N_3375);
nand U3590 (N_3590,N_3079,N_3218);
or U3591 (N_3591,N_3091,N_3196);
nor U3592 (N_3592,N_3493,N_3424);
or U3593 (N_3593,N_3441,N_3142);
nor U3594 (N_3594,N_3288,N_3225);
and U3595 (N_3595,N_3059,N_3217);
xnor U3596 (N_3596,N_3377,N_3409);
nand U3597 (N_3597,N_3341,N_3146);
nand U3598 (N_3598,N_3067,N_3052);
nand U3599 (N_3599,N_3108,N_3183);
or U3600 (N_3600,N_3350,N_3332);
nor U3601 (N_3601,N_3376,N_3055);
and U3602 (N_3602,N_3293,N_3184);
nand U3603 (N_3603,N_3402,N_3449);
nand U3604 (N_3604,N_3093,N_3106);
nand U3605 (N_3605,N_3214,N_3427);
and U3606 (N_3606,N_3400,N_3422);
nand U3607 (N_3607,N_3249,N_3092);
xor U3608 (N_3608,N_3361,N_3453);
and U3609 (N_3609,N_3362,N_3104);
or U3610 (N_3610,N_3431,N_3294);
or U3611 (N_3611,N_3291,N_3065);
and U3612 (N_3612,N_3372,N_3083);
and U3613 (N_3613,N_3031,N_3396);
nor U3614 (N_3614,N_3232,N_3336);
nor U3615 (N_3615,N_3333,N_3017);
or U3616 (N_3616,N_3452,N_3014);
xor U3617 (N_3617,N_3495,N_3237);
xor U3618 (N_3618,N_3243,N_3047);
and U3619 (N_3619,N_3213,N_3062);
and U3620 (N_3620,N_3216,N_3256);
xor U3621 (N_3621,N_3477,N_3051);
nor U3622 (N_3622,N_3130,N_3296);
nor U3623 (N_3623,N_3471,N_3470);
nand U3624 (N_3624,N_3118,N_3174);
or U3625 (N_3625,N_3257,N_3309);
xnor U3626 (N_3626,N_3458,N_3187);
nor U3627 (N_3627,N_3145,N_3194);
xor U3628 (N_3628,N_3032,N_3009);
nor U3629 (N_3629,N_3019,N_3036);
xor U3630 (N_3630,N_3227,N_3440);
and U3631 (N_3631,N_3063,N_3212);
xor U3632 (N_3632,N_3489,N_3412);
nand U3633 (N_3633,N_3190,N_3394);
or U3634 (N_3634,N_3221,N_3171);
and U3635 (N_3635,N_3392,N_3245);
and U3636 (N_3636,N_3263,N_3319);
nand U3637 (N_3637,N_3024,N_3286);
nand U3638 (N_3638,N_3469,N_3043);
nor U3639 (N_3639,N_3481,N_3443);
nor U3640 (N_3640,N_3222,N_3399);
nand U3641 (N_3641,N_3448,N_3457);
nor U3642 (N_3642,N_3125,N_3335);
and U3643 (N_3643,N_3094,N_3084);
nor U3644 (N_3644,N_3005,N_3007);
nor U3645 (N_3645,N_3181,N_3436);
nand U3646 (N_3646,N_3119,N_3182);
nand U3647 (N_3647,N_3328,N_3391);
or U3648 (N_3648,N_3352,N_3126);
or U3649 (N_3649,N_3433,N_3159);
nand U3650 (N_3650,N_3207,N_3262);
nand U3651 (N_3651,N_3045,N_3373);
and U3652 (N_3652,N_3437,N_3430);
nand U3653 (N_3653,N_3323,N_3381);
or U3654 (N_3654,N_3447,N_3165);
nor U3655 (N_3655,N_3046,N_3363);
nor U3656 (N_3656,N_3002,N_3107);
xor U3657 (N_3657,N_3117,N_3272);
and U3658 (N_3658,N_3462,N_3035);
xnor U3659 (N_3659,N_3483,N_3133);
or U3660 (N_3660,N_3346,N_3201);
and U3661 (N_3661,N_3305,N_3275);
nor U3662 (N_3662,N_3011,N_3444);
nand U3663 (N_3663,N_3311,N_3280);
nor U3664 (N_3664,N_3416,N_3244);
or U3665 (N_3665,N_3480,N_3186);
nand U3666 (N_3666,N_3281,N_3356);
nor U3667 (N_3667,N_3077,N_3486);
or U3668 (N_3668,N_3020,N_3450);
nand U3669 (N_3669,N_3304,N_3464);
nor U3670 (N_3670,N_3137,N_3096);
nor U3671 (N_3671,N_3326,N_3068);
xnor U3672 (N_3672,N_3071,N_3410);
nor U3673 (N_3673,N_3342,N_3347);
and U3674 (N_3674,N_3348,N_3251);
nand U3675 (N_3675,N_3287,N_3390);
and U3676 (N_3676,N_3042,N_3466);
xor U3677 (N_3677,N_3484,N_3278);
nand U3678 (N_3678,N_3406,N_3343);
or U3679 (N_3679,N_3074,N_3496);
or U3680 (N_3680,N_3123,N_3313);
and U3681 (N_3681,N_3056,N_3307);
nor U3682 (N_3682,N_3135,N_3456);
or U3683 (N_3683,N_3285,N_3374);
or U3684 (N_3684,N_3321,N_3166);
nand U3685 (N_3685,N_3122,N_3140);
xor U3686 (N_3686,N_3200,N_3006);
or U3687 (N_3687,N_3028,N_3329);
and U3688 (N_3688,N_3487,N_3401);
and U3689 (N_3689,N_3044,N_3421);
nor U3690 (N_3690,N_3366,N_3066);
or U3691 (N_3691,N_3053,N_3349);
nand U3692 (N_3692,N_3113,N_3226);
nor U3693 (N_3693,N_3105,N_3191);
nor U3694 (N_3694,N_3161,N_3151);
or U3695 (N_3695,N_3442,N_3152);
and U3696 (N_3696,N_3475,N_3189);
nand U3697 (N_3697,N_3473,N_3292);
xnor U3698 (N_3698,N_3195,N_3252);
xnor U3699 (N_3699,N_3308,N_3491);
nor U3700 (N_3700,N_3149,N_3150);
xor U3701 (N_3701,N_3467,N_3128);
xnor U3702 (N_3702,N_3314,N_3169);
nand U3703 (N_3703,N_3420,N_3306);
and U3704 (N_3704,N_3499,N_3331);
nor U3705 (N_3705,N_3098,N_3446);
nand U3706 (N_3706,N_3355,N_3141);
and U3707 (N_3707,N_3298,N_3238);
or U3708 (N_3708,N_3260,N_3353);
xnor U3709 (N_3709,N_3387,N_3153);
nand U3710 (N_3710,N_3197,N_3301);
nand U3711 (N_3711,N_3027,N_3340);
nand U3712 (N_3712,N_3271,N_3041);
nand U3713 (N_3713,N_3219,N_3013);
or U3714 (N_3714,N_3143,N_3100);
nand U3715 (N_3715,N_3242,N_3228);
or U3716 (N_3716,N_3176,N_3180);
nand U3717 (N_3717,N_3097,N_3081);
xnor U3718 (N_3718,N_3490,N_3038);
and U3719 (N_3719,N_3050,N_3246);
nand U3720 (N_3720,N_3034,N_3432);
nor U3721 (N_3721,N_3388,N_3154);
or U3722 (N_3722,N_3345,N_3254);
or U3723 (N_3723,N_3102,N_3297);
xor U3724 (N_3724,N_3203,N_3386);
or U3725 (N_3725,N_3316,N_3179);
nor U3726 (N_3726,N_3230,N_3357);
nand U3727 (N_3727,N_3408,N_3090);
and U3728 (N_3728,N_3398,N_3175);
nor U3729 (N_3729,N_3192,N_3172);
and U3730 (N_3730,N_3110,N_3231);
or U3731 (N_3731,N_3076,N_3206);
xnor U3732 (N_3732,N_3267,N_3264);
nand U3733 (N_3733,N_3429,N_3337);
or U3734 (N_3734,N_3255,N_3259);
and U3735 (N_3735,N_3124,N_3369);
nand U3736 (N_3736,N_3438,N_3290);
nor U3737 (N_3737,N_3086,N_3269);
nor U3738 (N_3738,N_3010,N_3229);
nor U3739 (N_3739,N_3215,N_3048);
or U3740 (N_3740,N_3266,N_3193);
nor U3741 (N_3741,N_3384,N_3004);
xor U3742 (N_3742,N_3109,N_3054);
nand U3743 (N_3743,N_3156,N_3075);
or U3744 (N_3744,N_3303,N_3116);
and U3745 (N_3745,N_3101,N_3157);
nand U3746 (N_3746,N_3463,N_3423);
xor U3747 (N_3747,N_3261,N_3351);
and U3748 (N_3748,N_3265,N_3474);
nor U3749 (N_3749,N_3037,N_3472);
and U3750 (N_3750,N_3452,N_3065);
nand U3751 (N_3751,N_3134,N_3118);
xor U3752 (N_3752,N_3332,N_3098);
and U3753 (N_3753,N_3063,N_3355);
or U3754 (N_3754,N_3456,N_3405);
or U3755 (N_3755,N_3376,N_3159);
or U3756 (N_3756,N_3241,N_3023);
nor U3757 (N_3757,N_3173,N_3214);
nand U3758 (N_3758,N_3166,N_3490);
nor U3759 (N_3759,N_3471,N_3228);
nand U3760 (N_3760,N_3461,N_3066);
nor U3761 (N_3761,N_3266,N_3362);
nand U3762 (N_3762,N_3173,N_3168);
and U3763 (N_3763,N_3060,N_3441);
and U3764 (N_3764,N_3192,N_3087);
and U3765 (N_3765,N_3151,N_3325);
nand U3766 (N_3766,N_3215,N_3031);
nor U3767 (N_3767,N_3132,N_3099);
nand U3768 (N_3768,N_3482,N_3493);
and U3769 (N_3769,N_3227,N_3272);
xor U3770 (N_3770,N_3455,N_3019);
nor U3771 (N_3771,N_3136,N_3493);
nand U3772 (N_3772,N_3482,N_3313);
xnor U3773 (N_3773,N_3301,N_3162);
and U3774 (N_3774,N_3168,N_3326);
nor U3775 (N_3775,N_3282,N_3206);
and U3776 (N_3776,N_3387,N_3104);
or U3777 (N_3777,N_3449,N_3461);
or U3778 (N_3778,N_3331,N_3208);
xnor U3779 (N_3779,N_3253,N_3250);
nor U3780 (N_3780,N_3333,N_3201);
or U3781 (N_3781,N_3063,N_3183);
xnor U3782 (N_3782,N_3351,N_3484);
and U3783 (N_3783,N_3312,N_3435);
nand U3784 (N_3784,N_3410,N_3147);
xnor U3785 (N_3785,N_3385,N_3086);
nand U3786 (N_3786,N_3398,N_3492);
xor U3787 (N_3787,N_3024,N_3199);
xnor U3788 (N_3788,N_3342,N_3004);
and U3789 (N_3789,N_3220,N_3469);
nand U3790 (N_3790,N_3059,N_3176);
nor U3791 (N_3791,N_3155,N_3121);
or U3792 (N_3792,N_3224,N_3066);
or U3793 (N_3793,N_3032,N_3149);
nor U3794 (N_3794,N_3100,N_3092);
or U3795 (N_3795,N_3004,N_3428);
and U3796 (N_3796,N_3089,N_3473);
nor U3797 (N_3797,N_3418,N_3412);
nand U3798 (N_3798,N_3338,N_3008);
nor U3799 (N_3799,N_3079,N_3272);
or U3800 (N_3800,N_3162,N_3282);
nor U3801 (N_3801,N_3426,N_3495);
nor U3802 (N_3802,N_3352,N_3096);
nor U3803 (N_3803,N_3412,N_3313);
nand U3804 (N_3804,N_3085,N_3196);
and U3805 (N_3805,N_3056,N_3373);
xor U3806 (N_3806,N_3351,N_3265);
and U3807 (N_3807,N_3039,N_3179);
nor U3808 (N_3808,N_3480,N_3496);
or U3809 (N_3809,N_3295,N_3154);
or U3810 (N_3810,N_3029,N_3383);
nor U3811 (N_3811,N_3291,N_3420);
xor U3812 (N_3812,N_3030,N_3366);
or U3813 (N_3813,N_3021,N_3141);
nand U3814 (N_3814,N_3090,N_3006);
xnor U3815 (N_3815,N_3217,N_3210);
or U3816 (N_3816,N_3104,N_3454);
and U3817 (N_3817,N_3094,N_3089);
or U3818 (N_3818,N_3128,N_3122);
xor U3819 (N_3819,N_3234,N_3073);
or U3820 (N_3820,N_3424,N_3143);
nor U3821 (N_3821,N_3484,N_3068);
and U3822 (N_3822,N_3335,N_3017);
nand U3823 (N_3823,N_3284,N_3278);
nor U3824 (N_3824,N_3050,N_3484);
and U3825 (N_3825,N_3269,N_3487);
nand U3826 (N_3826,N_3358,N_3461);
and U3827 (N_3827,N_3266,N_3119);
or U3828 (N_3828,N_3133,N_3321);
nand U3829 (N_3829,N_3168,N_3274);
and U3830 (N_3830,N_3320,N_3193);
or U3831 (N_3831,N_3350,N_3397);
or U3832 (N_3832,N_3110,N_3187);
nand U3833 (N_3833,N_3058,N_3287);
or U3834 (N_3834,N_3303,N_3198);
or U3835 (N_3835,N_3182,N_3150);
or U3836 (N_3836,N_3125,N_3443);
or U3837 (N_3837,N_3240,N_3166);
and U3838 (N_3838,N_3399,N_3185);
and U3839 (N_3839,N_3291,N_3386);
and U3840 (N_3840,N_3465,N_3417);
or U3841 (N_3841,N_3230,N_3111);
nor U3842 (N_3842,N_3359,N_3228);
nor U3843 (N_3843,N_3380,N_3223);
nor U3844 (N_3844,N_3406,N_3030);
nor U3845 (N_3845,N_3333,N_3024);
xnor U3846 (N_3846,N_3415,N_3170);
xnor U3847 (N_3847,N_3375,N_3350);
xnor U3848 (N_3848,N_3180,N_3270);
nor U3849 (N_3849,N_3061,N_3149);
nor U3850 (N_3850,N_3250,N_3180);
xor U3851 (N_3851,N_3234,N_3216);
nand U3852 (N_3852,N_3294,N_3281);
nor U3853 (N_3853,N_3042,N_3171);
and U3854 (N_3854,N_3395,N_3460);
nor U3855 (N_3855,N_3373,N_3209);
xor U3856 (N_3856,N_3167,N_3170);
nor U3857 (N_3857,N_3422,N_3444);
nand U3858 (N_3858,N_3348,N_3431);
nor U3859 (N_3859,N_3081,N_3409);
or U3860 (N_3860,N_3336,N_3357);
xor U3861 (N_3861,N_3484,N_3301);
xor U3862 (N_3862,N_3155,N_3474);
and U3863 (N_3863,N_3271,N_3012);
or U3864 (N_3864,N_3261,N_3443);
xor U3865 (N_3865,N_3152,N_3411);
nor U3866 (N_3866,N_3458,N_3160);
or U3867 (N_3867,N_3020,N_3357);
nand U3868 (N_3868,N_3309,N_3397);
xor U3869 (N_3869,N_3395,N_3177);
xor U3870 (N_3870,N_3150,N_3198);
nor U3871 (N_3871,N_3173,N_3352);
or U3872 (N_3872,N_3099,N_3103);
and U3873 (N_3873,N_3470,N_3112);
and U3874 (N_3874,N_3230,N_3051);
xnor U3875 (N_3875,N_3483,N_3057);
and U3876 (N_3876,N_3132,N_3399);
nor U3877 (N_3877,N_3402,N_3201);
and U3878 (N_3878,N_3292,N_3469);
xnor U3879 (N_3879,N_3035,N_3097);
and U3880 (N_3880,N_3222,N_3029);
nor U3881 (N_3881,N_3333,N_3300);
or U3882 (N_3882,N_3326,N_3398);
or U3883 (N_3883,N_3246,N_3243);
xor U3884 (N_3884,N_3167,N_3176);
nand U3885 (N_3885,N_3236,N_3449);
nor U3886 (N_3886,N_3167,N_3190);
nor U3887 (N_3887,N_3201,N_3409);
and U3888 (N_3888,N_3364,N_3051);
and U3889 (N_3889,N_3132,N_3227);
and U3890 (N_3890,N_3031,N_3459);
nor U3891 (N_3891,N_3273,N_3158);
xor U3892 (N_3892,N_3035,N_3051);
nor U3893 (N_3893,N_3307,N_3068);
xor U3894 (N_3894,N_3172,N_3042);
xnor U3895 (N_3895,N_3300,N_3187);
xor U3896 (N_3896,N_3120,N_3308);
nand U3897 (N_3897,N_3101,N_3377);
or U3898 (N_3898,N_3329,N_3421);
xor U3899 (N_3899,N_3407,N_3437);
nor U3900 (N_3900,N_3489,N_3046);
nor U3901 (N_3901,N_3038,N_3145);
nand U3902 (N_3902,N_3121,N_3406);
and U3903 (N_3903,N_3285,N_3279);
xor U3904 (N_3904,N_3230,N_3001);
xnor U3905 (N_3905,N_3350,N_3056);
xnor U3906 (N_3906,N_3029,N_3201);
xor U3907 (N_3907,N_3306,N_3250);
xor U3908 (N_3908,N_3237,N_3029);
nor U3909 (N_3909,N_3441,N_3055);
xor U3910 (N_3910,N_3350,N_3262);
or U3911 (N_3911,N_3175,N_3456);
nand U3912 (N_3912,N_3308,N_3180);
or U3913 (N_3913,N_3345,N_3128);
and U3914 (N_3914,N_3449,N_3108);
or U3915 (N_3915,N_3337,N_3173);
or U3916 (N_3916,N_3386,N_3435);
and U3917 (N_3917,N_3306,N_3129);
nor U3918 (N_3918,N_3124,N_3427);
and U3919 (N_3919,N_3261,N_3452);
nand U3920 (N_3920,N_3127,N_3282);
xnor U3921 (N_3921,N_3119,N_3167);
nor U3922 (N_3922,N_3290,N_3333);
or U3923 (N_3923,N_3147,N_3120);
nor U3924 (N_3924,N_3308,N_3469);
xor U3925 (N_3925,N_3495,N_3139);
nor U3926 (N_3926,N_3029,N_3357);
xor U3927 (N_3927,N_3451,N_3155);
and U3928 (N_3928,N_3289,N_3272);
nand U3929 (N_3929,N_3276,N_3074);
xor U3930 (N_3930,N_3305,N_3376);
nand U3931 (N_3931,N_3210,N_3077);
nor U3932 (N_3932,N_3021,N_3205);
nor U3933 (N_3933,N_3273,N_3262);
xor U3934 (N_3934,N_3045,N_3076);
or U3935 (N_3935,N_3036,N_3071);
and U3936 (N_3936,N_3303,N_3168);
xor U3937 (N_3937,N_3052,N_3436);
and U3938 (N_3938,N_3432,N_3284);
and U3939 (N_3939,N_3255,N_3451);
xnor U3940 (N_3940,N_3078,N_3412);
nand U3941 (N_3941,N_3086,N_3120);
xnor U3942 (N_3942,N_3038,N_3051);
xnor U3943 (N_3943,N_3394,N_3092);
xnor U3944 (N_3944,N_3156,N_3273);
and U3945 (N_3945,N_3283,N_3105);
or U3946 (N_3946,N_3209,N_3383);
and U3947 (N_3947,N_3339,N_3072);
nand U3948 (N_3948,N_3341,N_3074);
and U3949 (N_3949,N_3152,N_3441);
or U3950 (N_3950,N_3142,N_3099);
nand U3951 (N_3951,N_3494,N_3379);
or U3952 (N_3952,N_3205,N_3143);
or U3953 (N_3953,N_3076,N_3466);
nor U3954 (N_3954,N_3475,N_3460);
nand U3955 (N_3955,N_3449,N_3104);
or U3956 (N_3956,N_3454,N_3117);
nor U3957 (N_3957,N_3372,N_3456);
xnor U3958 (N_3958,N_3342,N_3282);
and U3959 (N_3959,N_3107,N_3171);
or U3960 (N_3960,N_3406,N_3244);
nand U3961 (N_3961,N_3142,N_3340);
or U3962 (N_3962,N_3014,N_3174);
xnor U3963 (N_3963,N_3359,N_3273);
xor U3964 (N_3964,N_3382,N_3308);
nor U3965 (N_3965,N_3310,N_3127);
nor U3966 (N_3966,N_3480,N_3464);
or U3967 (N_3967,N_3350,N_3187);
nor U3968 (N_3968,N_3209,N_3239);
or U3969 (N_3969,N_3466,N_3447);
nor U3970 (N_3970,N_3487,N_3434);
or U3971 (N_3971,N_3304,N_3422);
or U3972 (N_3972,N_3170,N_3358);
or U3973 (N_3973,N_3249,N_3000);
and U3974 (N_3974,N_3216,N_3164);
and U3975 (N_3975,N_3163,N_3262);
nand U3976 (N_3976,N_3136,N_3356);
nor U3977 (N_3977,N_3379,N_3199);
or U3978 (N_3978,N_3023,N_3372);
and U3979 (N_3979,N_3018,N_3020);
nand U3980 (N_3980,N_3135,N_3367);
xor U3981 (N_3981,N_3095,N_3488);
or U3982 (N_3982,N_3382,N_3364);
nand U3983 (N_3983,N_3317,N_3402);
nand U3984 (N_3984,N_3406,N_3226);
xnor U3985 (N_3985,N_3466,N_3295);
xnor U3986 (N_3986,N_3095,N_3129);
xnor U3987 (N_3987,N_3188,N_3032);
xnor U3988 (N_3988,N_3259,N_3381);
and U3989 (N_3989,N_3163,N_3464);
and U3990 (N_3990,N_3379,N_3027);
or U3991 (N_3991,N_3127,N_3124);
or U3992 (N_3992,N_3179,N_3056);
nand U3993 (N_3993,N_3385,N_3111);
or U3994 (N_3994,N_3058,N_3262);
or U3995 (N_3995,N_3132,N_3490);
and U3996 (N_3996,N_3048,N_3376);
nand U3997 (N_3997,N_3481,N_3210);
nand U3998 (N_3998,N_3498,N_3284);
nor U3999 (N_3999,N_3305,N_3037);
nand U4000 (N_4000,N_3845,N_3967);
xnor U4001 (N_4001,N_3997,N_3918);
nor U4002 (N_4002,N_3765,N_3783);
nor U4003 (N_4003,N_3907,N_3771);
and U4004 (N_4004,N_3640,N_3915);
and U4005 (N_4005,N_3697,N_3549);
and U4006 (N_4006,N_3841,N_3763);
and U4007 (N_4007,N_3725,N_3564);
and U4008 (N_4008,N_3834,N_3682);
nand U4009 (N_4009,N_3579,N_3539);
nand U4010 (N_4010,N_3795,N_3869);
xnor U4011 (N_4011,N_3751,N_3840);
or U4012 (N_4012,N_3599,N_3591);
xor U4013 (N_4013,N_3936,N_3571);
nor U4014 (N_4014,N_3729,N_3502);
nand U4015 (N_4015,N_3961,N_3891);
and U4016 (N_4016,N_3919,N_3605);
nand U4017 (N_4017,N_3780,N_3755);
or U4018 (N_4018,N_3817,N_3576);
and U4019 (N_4019,N_3596,N_3636);
and U4020 (N_4020,N_3506,N_3542);
nand U4021 (N_4021,N_3732,N_3882);
or U4022 (N_4022,N_3673,N_3857);
nor U4023 (N_4023,N_3581,N_3876);
and U4024 (N_4024,N_3554,N_3730);
nand U4025 (N_4025,N_3672,N_3828);
and U4026 (N_4026,N_3886,N_3735);
or U4027 (N_4027,N_3505,N_3566);
nand U4028 (N_4028,N_3597,N_3894);
or U4029 (N_4029,N_3509,N_3519);
xnor U4030 (N_4030,N_3706,N_3692);
or U4031 (N_4031,N_3601,N_3777);
or U4032 (N_4032,N_3609,N_3525);
nand U4033 (N_4033,N_3635,N_3943);
or U4034 (N_4034,N_3626,N_3529);
nand U4035 (N_4035,N_3719,N_3563);
xnor U4036 (N_4036,N_3871,N_3955);
nand U4037 (N_4037,N_3810,N_3741);
nor U4038 (N_4038,N_3880,N_3799);
nor U4039 (N_4039,N_3931,N_3518);
nand U4040 (N_4040,N_3990,N_3790);
nand U4041 (N_4041,N_3911,N_3717);
nor U4042 (N_4042,N_3973,N_3612);
nand U4043 (N_4043,N_3941,N_3949);
nor U4044 (N_4044,N_3514,N_3813);
nor U4045 (N_4045,N_3649,N_3785);
and U4046 (N_4046,N_3831,N_3541);
nor U4047 (N_4047,N_3701,N_3690);
nand U4048 (N_4048,N_3570,N_3711);
and U4049 (N_4049,N_3504,N_3957);
or U4050 (N_4050,N_3675,N_3913);
and U4051 (N_4051,N_3996,N_3586);
nor U4052 (N_4052,N_3698,N_3677);
and U4053 (N_4053,N_3522,N_3778);
nor U4054 (N_4054,N_3801,N_3602);
xnor U4055 (N_4055,N_3528,N_3663);
nor U4056 (N_4056,N_3708,N_3513);
xnor U4057 (N_4057,N_3829,N_3971);
or U4058 (N_4058,N_3510,N_3854);
or U4059 (N_4059,N_3569,N_3620);
or U4060 (N_4060,N_3629,N_3800);
xor U4061 (N_4061,N_3768,N_3760);
nand U4062 (N_4062,N_3945,N_3809);
or U4063 (N_4063,N_3912,N_3753);
nand U4064 (N_4064,N_3835,N_3986);
and U4065 (N_4065,N_3762,N_3713);
and U4066 (N_4066,N_3885,N_3979);
nand U4067 (N_4067,N_3865,N_3926);
xnor U4068 (N_4068,N_3664,N_3921);
or U4069 (N_4069,N_3822,N_3733);
or U4070 (N_4070,N_3544,N_3534);
nand U4071 (N_4071,N_3639,N_3842);
xor U4072 (N_4072,N_3693,N_3736);
or U4073 (N_4073,N_3665,N_3545);
nand U4074 (N_4074,N_3982,N_3547);
xor U4075 (N_4075,N_3781,N_3740);
or U4076 (N_4076,N_3896,N_3798);
xor U4077 (N_4077,N_3653,N_3685);
nor U4078 (N_4078,N_3618,N_3718);
nor U4079 (N_4079,N_3844,N_3981);
and U4080 (N_4080,N_3860,N_3747);
or U4081 (N_4081,N_3978,N_3558);
and U4082 (N_4082,N_3657,N_3999);
xnor U4083 (N_4083,N_3577,N_3917);
and U4084 (N_4084,N_3826,N_3786);
xor U4085 (N_4085,N_3695,N_3723);
nand U4086 (N_4086,N_3952,N_3895);
xnor U4087 (N_4087,N_3775,N_3802);
nand U4088 (N_4088,N_3816,N_3501);
or U4089 (N_4089,N_3633,N_3807);
or U4090 (N_4090,N_3617,N_3744);
nand U4091 (N_4091,N_3565,N_3739);
nand U4092 (N_4092,N_3646,N_3837);
nand U4093 (N_4093,N_3779,N_3870);
xor U4094 (N_4094,N_3856,N_3500);
xnor U4095 (N_4095,N_3988,N_3772);
and U4096 (N_4096,N_3667,N_3658);
nand U4097 (N_4097,N_3937,N_3940);
xnor U4098 (N_4098,N_3587,N_3552);
xnor U4099 (N_4099,N_3622,N_3855);
and U4100 (N_4100,N_3866,N_3625);
nand U4101 (N_4101,N_3980,N_3811);
nand U4102 (N_4102,N_3890,N_3964);
or U4103 (N_4103,N_3742,N_3787);
and U4104 (N_4104,N_3696,N_3903);
nor U4105 (N_4105,N_3796,N_3849);
nand U4106 (N_4106,N_3608,N_3909);
or U4107 (N_4107,N_3852,N_3572);
nor U4108 (N_4108,N_3950,N_3976);
nand U4109 (N_4109,N_3606,N_3580);
xnor U4110 (N_4110,N_3887,N_3864);
nor U4111 (N_4111,N_3604,N_3645);
xnor U4112 (N_4112,N_3647,N_3968);
nor U4113 (N_4113,N_3610,N_3823);
nand U4114 (N_4114,N_3648,N_3704);
nand U4115 (N_4115,N_3881,N_3557);
and U4116 (N_4116,N_3536,N_3707);
or U4117 (N_4117,N_3910,N_3676);
or U4118 (N_4118,N_3644,N_3944);
or U4119 (N_4119,N_3818,N_3517);
xnor U4120 (N_4120,N_3769,N_3963);
or U4121 (N_4121,N_3562,N_3630);
xnor U4122 (N_4122,N_3899,N_3641);
and U4123 (N_4123,N_3992,N_3767);
or U4124 (N_4124,N_3995,N_3590);
nor U4125 (N_4125,N_3638,N_3752);
and U4126 (N_4126,N_3589,N_3947);
and U4127 (N_4127,N_3819,N_3958);
nor U4128 (N_4128,N_3642,N_3731);
nand U4129 (N_4129,N_3862,N_3898);
and U4130 (N_4130,N_3593,N_3803);
and U4131 (N_4131,N_3948,N_3508);
or U4132 (N_4132,N_3567,N_3627);
or U4133 (N_4133,N_3993,N_3634);
nand U4134 (N_4134,N_3678,N_3594);
nor U4135 (N_4135,N_3836,N_3754);
xor U4136 (N_4136,N_3619,N_3843);
nor U4137 (N_4137,N_3600,N_3651);
and U4138 (N_4138,N_3660,N_3575);
nand U4139 (N_4139,N_3928,N_3812);
xnor U4140 (N_4140,N_3994,N_3724);
or U4141 (N_4141,N_3537,N_3598);
nor U4142 (N_4142,N_3561,N_3684);
or U4143 (N_4143,N_3868,N_3694);
nand U4144 (N_4144,N_3942,N_3671);
and U4145 (N_4145,N_3776,N_3901);
nand U4146 (N_4146,N_3616,N_3543);
nand U4147 (N_4147,N_3867,N_3592);
xor U4148 (N_4148,N_3631,N_3923);
nand U4149 (N_4149,N_3987,N_3861);
nand U4150 (N_4150,N_3998,N_3535);
nor U4151 (N_4151,N_3878,N_3568);
xnor U4152 (N_4152,N_3965,N_3797);
nand U4153 (N_4153,N_3839,N_3656);
nand U4154 (N_4154,N_3766,N_3689);
nor U4155 (N_4155,N_3975,N_3532);
nand U4156 (N_4156,N_3661,N_3560);
or U4157 (N_4157,N_3832,N_3956);
nand U4158 (N_4158,N_3905,N_3615);
nand U4159 (N_4159,N_3520,N_3873);
xnor U4160 (N_4160,N_3756,N_3749);
and U4161 (N_4161,N_3850,N_3573);
or U4162 (N_4162,N_3827,N_3582);
xnor U4163 (N_4163,N_3916,N_3794);
xnor U4164 (N_4164,N_3788,N_3507);
xnor U4165 (N_4165,N_3897,N_3720);
and U4166 (N_4166,N_3659,N_3924);
and U4167 (N_4167,N_3691,N_3515);
and U4168 (N_4168,N_3674,N_3847);
nand U4169 (N_4169,N_3530,N_3974);
xnor U4170 (N_4170,N_3516,N_3546);
nor U4171 (N_4171,N_3578,N_3758);
nor U4172 (N_4172,N_3521,N_3551);
xor U4173 (N_4173,N_3621,N_3884);
nand U4174 (N_4174,N_3970,N_3791);
and U4175 (N_4175,N_3666,N_3585);
or U4176 (N_4176,N_3683,N_3709);
nand U4177 (N_4177,N_3538,N_3574);
or U4178 (N_4178,N_3726,N_3938);
nor U4179 (N_4179,N_3746,N_3681);
nor U4180 (N_4180,N_3652,N_3548);
nor U4181 (N_4181,N_3748,N_3833);
and U4182 (N_4182,N_3523,N_3670);
nor U4183 (N_4183,N_3906,N_3699);
or U4184 (N_4184,N_3728,N_3983);
nor U4185 (N_4185,N_3904,N_3680);
xnor U4186 (N_4186,N_3888,N_3930);
nand U4187 (N_4187,N_3556,N_3782);
xor U4188 (N_4188,N_3784,N_3902);
and U4189 (N_4189,N_3959,N_3705);
nand U4190 (N_4190,N_3972,N_3738);
xnor U4191 (N_4191,N_3929,N_3792);
and U4192 (N_4192,N_3679,N_3757);
xor U4193 (N_4193,N_3553,N_3511);
nor U4194 (N_4194,N_3951,N_3820);
and U4195 (N_4195,N_3774,N_3700);
xor U4196 (N_4196,N_3540,N_3946);
or U4197 (N_4197,N_3848,N_3814);
nand U4198 (N_4198,N_3623,N_3650);
nand U4199 (N_4199,N_3991,N_3922);
nand U4200 (N_4200,N_3953,N_3628);
and U4201 (N_4201,N_3584,N_3858);
and U4202 (N_4202,N_3927,N_3688);
or U4203 (N_4203,N_3825,N_3703);
nor U4204 (N_4204,N_3875,N_3874);
xor U4205 (N_4205,N_3607,N_3550);
nand U4206 (N_4206,N_3984,N_3893);
nand U4207 (N_4207,N_3512,N_3863);
or U4208 (N_4208,N_3687,N_3734);
nor U4209 (N_4209,N_3555,N_3883);
xnor U4210 (N_4210,N_3824,N_3595);
nor U4211 (N_4211,N_3533,N_3889);
xor U4212 (N_4212,N_3808,N_3613);
nor U4213 (N_4213,N_3770,N_3830);
xnor U4214 (N_4214,N_3804,N_3920);
xor U4215 (N_4215,N_3846,N_3892);
xor U4216 (N_4216,N_3686,N_3524);
xor U4217 (N_4217,N_3908,N_3727);
and U4218 (N_4218,N_3851,N_3935);
or U4219 (N_4219,N_3603,N_3900);
nor U4220 (N_4220,N_3531,N_3722);
nor U4221 (N_4221,N_3714,N_3614);
nor U4222 (N_4222,N_3793,N_3933);
nor U4223 (N_4223,N_3872,N_3526);
nand U4224 (N_4224,N_3669,N_3962);
or U4225 (N_4225,N_3702,N_3914);
nand U4226 (N_4226,N_3815,N_3668);
and U4227 (N_4227,N_3838,N_3662);
or U4228 (N_4228,N_3806,N_3503);
nand U4229 (N_4229,N_3934,N_3637);
nor U4230 (N_4230,N_3712,N_3737);
nor U4231 (N_4231,N_3977,N_3716);
or U4232 (N_4232,N_3939,N_3527);
and U4233 (N_4233,N_3932,N_3710);
or U4234 (N_4234,N_3721,N_3960);
nand U4235 (N_4235,N_3821,N_3877);
or U4236 (N_4236,N_3750,N_3925);
or U4237 (N_4237,N_3853,N_3583);
nand U4238 (N_4238,N_3879,N_3632);
nand U4239 (N_4239,N_3655,N_3759);
xnor U4240 (N_4240,N_3985,N_3643);
nor U4241 (N_4241,N_3745,N_3859);
nor U4242 (N_4242,N_3764,N_3624);
or U4243 (N_4243,N_3954,N_3773);
and U4244 (N_4244,N_3654,N_3966);
xor U4245 (N_4245,N_3805,N_3789);
xor U4246 (N_4246,N_3559,N_3588);
or U4247 (N_4247,N_3611,N_3969);
or U4248 (N_4248,N_3761,N_3743);
xnor U4249 (N_4249,N_3715,N_3989);
xor U4250 (N_4250,N_3882,N_3870);
and U4251 (N_4251,N_3670,N_3739);
nor U4252 (N_4252,N_3922,N_3740);
or U4253 (N_4253,N_3978,N_3777);
nor U4254 (N_4254,N_3505,N_3709);
and U4255 (N_4255,N_3834,N_3769);
xnor U4256 (N_4256,N_3633,N_3902);
nor U4257 (N_4257,N_3522,N_3916);
or U4258 (N_4258,N_3792,N_3721);
xnor U4259 (N_4259,N_3928,N_3666);
and U4260 (N_4260,N_3947,N_3844);
nor U4261 (N_4261,N_3934,N_3825);
xnor U4262 (N_4262,N_3764,N_3549);
or U4263 (N_4263,N_3578,N_3763);
or U4264 (N_4264,N_3569,N_3688);
or U4265 (N_4265,N_3652,N_3881);
xnor U4266 (N_4266,N_3783,N_3928);
or U4267 (N_4267,N_3995,N_3589);
or U4268 (N_4268,N_3721,N_3568);
nor U4269 (N_4269,N_3682,N_3977);
or U4270 (N_4270,N_3731,N_3783);
xor U4271 (N_4271,N_3721,N_3765);
or U4272 (N_4272,N_3798,N_3826);
or U4273 (N_4273,N_3735,N_3750);
nor U4274 (N_4274,N_3824,N_3851);
and U4275 (N_4275,N_3960,N_3843);
nand U4276 (N_4276,N_3762,N_3543);
nand U4277 (N_4277,N_3905,N_3611);
xnor U4278 (N_4278,N_3696,N_3967);
xnor U4279 (N_4279,N_3850,N_3720);
nor U4280 (N_4280,N_3707,N_3887);
nand U4281 (N_4281,N_3848,N_3569);
nor U4282 (N_4282,N_3782,N_3851);
and U4283 (N_4283,N_3903,N_3647);
xnor U4284 (N_4284,N_3877,N_3768);
nand U4285 (N_4285,N_3806,N_3708);
xor U4286 (N_4286,N_3686,N_3671);
nand U4287 (N_4287,N_3731,N_3741);
nor U4288 (N_4288,N_3909,N_3763);
or U4289 (N_4289,N_3841,N_3993);
nand U4290 (N_4290,N_3906,N_3662);
and U4291 (N_4291,N_3578,N_3702);
or U4292 (N_4292,N_3573,N_3840);
nand U4293 (N_4293,N_3948,N_3986);
nor U4294 (N_4294,N_3906,N_3668);
or U4295 (N_4295,N_3576,N_3849);
nor U4296 (N_4296,N_3677,N_3754);
and U4297 (N_4297,N_3917,N_3593);
and U4298 (N_4298,N_3791,N_3634);
or U4299 (N_4299,N_3524,N_3819);
and U4300 (N_4300,N_3896,N_3925);
xnor U4301 (N_4301,N_3911,N_3528);
or U4302 (N_4302,N_3726,N_3878);
and U4303 (N_4303,N_3945,N_3916);
xor U4304 (N_4304,N_3864,N_3741);
nand U4305 (N_4305,N_3725,N_3917);
nor U4306 (N_4306,N_3887,N_3617);
nor U4307 (N_4307,N_3722,N_3500);
xor U4308 (N_4308,N_3772,N_3817);
and U4309 (N_4309,N_3542,N_3838);
and U4310 (N_4310,N_3560,N_3686);
or U4311 (N_4311,N_3566,N_3670);
nand U4312 (N_4312,N_3738,N_3508);
xnor U4313 (N_4313,N_3650,N_3877);
nand U4314 (N_4314,N_3814,N_3524);
or U4315 (N_4315,N_3942,N_3532);
nand U4316 (N_4316,N_3958,N_3667);
and U4317 (N_4317,N_3559,N_3743);
xor U4318 (N_4318,N_3863,N_3534);
and U4319 (N_4319,N_3691,N_3999);
nor U4320 (N_4320,N_3954,N_3604);
nor U4321 (N_4321,N_3962,N_3686);
nand U4322 (N_4322,N_3533,N_3880);
nor U4323 (N_4323,N_3986,N_3527);
and U4324 (N_4324,N_3914,N_3627);
nor U4325 (N_4325,N_3522,N_3856);
nor U4326 (N_4326,N_3917,N_3633);
nor U4327 (N_4327,N_3909,N_3619);
nor U4328 (N_4328,N_3992,N_3646);
xor U4329 (N_4329,N_3926,N_3582);
nand U4330 (N_4330,N_3954,N_3538);
xor U4331 (N_4331,N_3856,N_3640);
nor U4332 (N_4332,N_3833,N_3669);
or U4333 (N_4333,N_3717,N_3622);
or U4334 (N_4334,N_3675,N_3829);
xnor U4335 (N_4335,N_3752,N_3820);
or U4336 (N_4336,N_3960,N_3738);
and U4337 (N_4337,N_3702,N_3509);
xnor U4338 (N_4338,N_3872,N_3592);
or U4339 (N_4339,N_3635,N_3968);
and U4340 (N_4340,N_3669,N_3748);
xnor U4341 (N_4341,N_3750,N_3815);
and U4342 (N_4342,N_3739,N_3815);
xor U4343 (N_4343,N_3756,N_3697);
nand U4344 (N_4344,N_3569,N_3868);
or U4345 (N_4345,N_3814,N_3892);
nand U4346 (N_4346,N_3636,N_3971);
xnor U4347 (N_4347,N_3531,N_3832);
nor U4348 (N_4348,N_3840,N_3741);
xnor U4349 (N_4349,N_3777,N_3977);
nand U4350 (N_4350,N_3739,N_3737);
and U4351 (N_4351,N_3644,N_3551);
or U4352 (N_4352,N_3694,N_3562);
xnor U4353 (N_4353,N_3999,N_3514);
xnor U4354 (N_4354,N_3948,N_3800);
or U4355 (N_4355,N_3896,N_3953);
or U4356 (N_4356,N_3648,N_3952);
nand U4357 (N_4357,N_3999,N_3554);
or U4358 (N_4358,N_3539,N_3914);
nor U4359 (N_4359,N_3602,N_3792);
nor U4360 (N_4360,N_3500,N_3909);
nand U4361 (N_4361,N_3626,N_3784);
nand U4362 (N_4362,N_3963,N_3597);
nand U4363 (N_4363,N_3949,N_3530);
xor U4364 (N_4364,N_3778,N_3887);
and U4365 (N_4365,N_3613,N_3771);
nand U4366 (N_4366,N_3688,N_3892);
or U4367 (N_4367,N_3719,N_3883);
nor U4368 (N_4368,N_3544,N_3538);
xor U4369 (N_4369,N_3641,N_3605);
or U4370 (N_4370,N_3761,N_3946);
nand U4371 (N_4371,N_3569,N_3797);
and U4372 (N_4372,N_3580,N_3690);
or U4373 (N_4373,N_3561,N_3883);
nor U4374 (N_4374,N_3996,N_3810);
xnor U4375 (N_4375,N_3873,N_3797);
or U4376 (N_4376,N_3964,N_3938);
nor U4377 (N_4377,N_3766,N_3909);
nand U4378 (N_4378,N_3757,N_3799);
xnor U4379 (N_4379,N_3882,N_3939);
nor U4380 (N_4380,N_3567,N_3884);
nand U4381 (N_4381,N_3609,N_3666);
or U4382 (N_4382,N_3841,N_3657);
or U4383 (N_4383,N_3929,N_3651);
nand U4384 (N_4384,N_3885,N_3592);
and U4385 (N_4385,N_3523,N_3626);
xor U4386 (N_4386,N_3713,N_3978);
or U4387 (N_4387,N_3998,N_3789);
nor U4388 (N_4388,N_3709,N_3993);
nor U4389 (N_4389,N_3905,N_3888);
or U4390 (N_4390,N_3791,N_3995);
nor U4391 (N_4391,N_3988,N_3538);
nor U4392 (N_4392,N_3506,N_3807);
or U4393 (N_4393,N_3790,N_3808);
nor U4394 (N_4394,N_3806,N_3900);
nand U4395 (N_4395,N_3704,N_3501);
and U4396 (N_4396,N_3968,N_3960);
or U4397 (N_4397,N_3848,N_3923);
nand U4398 (N_4398,N_3782,N_3947);
nand U4399 (N_4399,N_3513,N_3831);
xor U4400 (N_4400,N_3804,N_3528);
xnor U4401 (N_4401,N_3588,N_3856);
nand U4402 (N_4402,N_3698,N_3648);
and U4403 (N_4403,N_3829,N_3863);
xor U4404 (N_4404,N_3556,N_3913);
and U4405 (N_4405,N_3823,N_3791);
xnor U4406 (N_4406,N_3927,N_3898);
nand U4407 (N_4407,N_3834,N_3651);
or U4408 (N_4408,N_3779,N_3557);
xnor U4409 (N_4409,N_3589,N_3801);
and U4410 (N_4410,N_3807,N_3761);
xnor U4411 (N_4411,N_3862,N_3731);
nand U4412 (N_4412,N_3699,N_3898);
nand U4413 (N_4413,N_3600,N_3883);
nor U4414 (N_4414,N_3697,N_3874);
nor U4415 (N_4415,N_3670,N_3775);
or U4416 (N_4416,N_3917,N_3874);
xnor U4417 (N_4417,N_3643,N_3905);
and U4418 (N_4418,N_3962,N_3600);
nand U4419 (N_4419,N_3700,N_3944);
nor U4420 (N_4420,N_3940,N_3934);
xor U4421 (N_4421,N_3906,N_3707);
nand U4422 (N_4422,N_3862,N_3965);
nand U4423 (N_4423,N_3789,N_3601);
xnor U4424 (N_4424,N_3732,N_3915);
or U4425 (N_4425,N_3999,N_3804);
nor U4426 (N_4426,N_3671,N_3735);
or U4427 (N_4427,N_3798,N_3863);
nand U4428 (N_4428,N_3596,N_3888);
nor U4429 (N_4429,N_3500,N_3761);
xnor U4430 (N_4430,N_3612,N_3546);
nor U4431 (N_4431,N_3984,N_3599);
or U4432 (N_4432,N_3803,N_3926);
nor U4433 (N_4433,N_3941,N_3729);
and U4434 (N_4434,N_3961,N_3535);
nor U4435 (N_4435,N_3786,N_3749);
nand U4436 (N_4436,N_3610,N_3914);
and U4437 (N_4437,N_3970,N_3782);
nand U4438 (N_4438,N_3795,N_3815);
xnor U4439 (N_4439,N_3702,N_3737);
or U4440 (N_4440,N_3821,N_3800);
nor U4441 (N_4441,N_3619,N_3788);
and U4442 (N_4442,N_3575,N_3652);
nand U4443 (N_4443,N_3803,N_3798);
nand U4444 (N_4444,N_3929,N_3902);
or U4445 (N_4445,N_3825,N_3603);
nand U4446 (N_4446,N_3835,N_3886);
nor U4447 (N_4447,N_3962,N_3984);
and U4448 (N_4448,N_3724,N_3891);
xor U4449 (N_4449,N_3677,N_3792);
or U4450 (N_4450,N_3594,N_3860);
and U4451 (N_4451,N_3952,N_3533);
nor U4452 (N_4452,N_3696,N_3643);
and U4453 (N_4453,N_3849,N_3851);
or U4454 (N_4454,N_3673,N_3601);
and U4455 (N_4455,N_3583,N_3773);
or U4456 (N_4456,N_3989,N_3916);
or U4457 (N_4457,N_3819,N_3861);
xor U4458 (N_4458,N_3691,N_3681);
or U4459 (N_4459,N_3720,N_3860);
nand U4460 (N_4460,N_3961,N_3645);
xnor U4461 (N_4461,N_3858,N_3552);
nor U4462 (N_4462,N_3970,N_3717);
and U4463 (N_4463,N_3682,N_3646);
xor U4464 (N_4464,N_3981,N_3901);
nor U4465 (N_4465,N_3561,N_3731);
or U4466 (N_4466,N_3632,N_3903);
xnor U4467 (N_4467,N_3987,N_3858);
xnor U4468 (N_4468,N_3987,N_3542);
and U4469 (N_4469,N_3582,N_3777);
xnor U4470 (N_4470,N_3976,N_3669);
nand U4471 (N_4471,N_3953,N_3624);
xor U4472 (N_4472,N_3932,N_3928);
or U4473 (N_4473,N_3537,N_3863);
nand U4474 (N_4474,N_3840,N_3774);
xor U4475 (N_4475,N_3934,N_3998);
and U4476 (N_4476,N_3978,N_3969);
xnor U4477 (N_4477,N_3526,N_3607);
or U4478 (N_4478,N_3956,N_3997);
nor U4479 (N_4479,N_3730,N_3697);
xnor U4480 (N_4480,N_3790,N_3700);
nand U4481 (N_4481,N_3741,N_3671);
and U4482 (N_4482,N_3859,N_3856);
nor U4483 (N_4483,N_3917,N_3642);
nand U4484 (N_4484,N_3580,N_3955);
xnor U4485 (N_4485,N_3705,N_3710);
nand U4486 (N_4486,N_3942,N_3983);
or U4487 (N_4487,N_3630,N_3981);
nand U4488 (N_4488,N_3656,N_3772);
and U4489 (N_4489,N_3563,N_3527);
and U4490 (N_4490,N_3677,N_3782);
or U4491 (N_4491,N_3912,N_3738);
nand U4492 (N_4492,N_3963,N_3979);
or U4493 (N_4493,N_3535,N_3756);
nand U4494 (N_4494,N_3714,N_3968);
nor U4495 (N_4495,N_3786,N_3723);
xor U4496 (N_4496,N_3590,N_3610);
and U4497 (N_4497,N_3768,N_3620);
nor U4498 (N_4498,N_3881,N_3813);
xnor U4499 (N_4499,N_3582,N_3603);
xnor U4500 (N_4500,N_4200,N_4275);
and U4501 (N_4501,N_4298,N_4420);
and U4502 (N_4502,N_4234,N_4262);
nor U4503 (N_4503,N_4170,N_4155);
xor U4504 (N_4504,N_4021,N_4294);
nand U4505 (N_4505,N_4401,N_4154);
nor U4506 (N_4506,N_4403,N_4457);
nand U4507 (N_4507,N_4141,N_4211);
xnor U4508 (N_4508,N_4304,N_4243);
or U4509 (N_4509,N_4491,N_4138);
xnor U4510 (N_4510,N_4425,N_4173);
xnor U4511 (N_4511,N_4269,N_4383);
nand U4512 (N_4512,N_4185,N_4108);
nand U4513 (N_4513,N_4373,N_4033);
or U4514 (N_4514,N_4288,N_4448);
xnor U4515 (N_4515,N_4086,N_4410);
nand U4516 (N_4516,N_4011,N_4067);
or U4517 (N_4517,N_4120,N_4007);
xor U4518 (N_4518,N_4219,N_4048);
and U4519 (N_4519,N_4010,N_4441);
or U4520 (N_4520,N_4017,N_4259);
nand U4521 (N_4521,N_4334,N_4140);
or U4522 (N_4522,N_4359,N_4081);
and U4523 (N_4523,N_4100,N_4488);
and U4524 (N_4524,N_4476,N_4110);
or U4525 (N_4525,N_4146,N_4054);
or U4526 (N_4526,N_4272,N_4064);
nor U4527 (N_4527,N_4443,N_4295);
nand U4528 (N_4528,N_4088,N_4467);
or U4529 (N_4529,N_4169,N_4144);
nor U4530 (N_4530,N_4254,N_4193);
or U4531 (N_4531,N_4437,N_4228);
nor U4532 (N_4532,N_4096,N_4050);
and U4533 (N_4533,N_4418,N_4014);
nand U4534 (N_4534,N_4280,N_4332);
nor U4535 (N_4535,N_4343,N_4182);
nand U4536 (N_4536,N_4092,N_4498);
or U4537 (N_4537,N_4492,N_4245);
and U4538 (N_4538,N_4205,N_4263);
and U4539 (N_4539,N_4112,N_4020);
xnor U4540 (N_4540,N_4106,N_4432);
or U4541 (N_4541,N_4416,N_4206);
nor U4542 (N_4542,N_4306,N_4315);
nor U4543 (N_4543,N_4151,N_4352);
nor U4544 (N_4544,N_4013,N_4123);
and U4545 (N_4545,N_4345,N_4271);
or U4546 (N_4546,N_4446,N_4019);
nor U4547 (N_4547,N_4232,N_4479);
nor U4548 (N_4548,N_4411,N_4134);
nor U4549 (N_4549,N_4415,N_4355);
nor U4550 (N_4550,N_4028,N_4165);
xnor U4551 (N_4551,N_4047,N_4284);
and U4552 (N_4552,N_4133,N_4237);
nand U4553 (N_4553,N_4122,N_4408);
nand U4554 (N_4554,N_4235,N_4117);
or U4555 (N_4555,N_4392,N_4236);
and U4556 (N_4556,N_4043,N_4220);
nor U4557 (N_4557,N_4402,N_4209);
or U4558 (N_4558,N_4319,N_4227);
nor U4559 (N_4559,N_4389,N_4059);
xnor U4560 (N_4560,N_4396,N_4353);
and U4561 (N_4561,N_4147,N_4356);
or U4562 (N_4562,N_4070,N_4285);
and U4563 (N_4563,N_4176,N_4366);
or U4564 (N_4564,N_4296,N_4222);
xor U4565 (N_4565,N_4022,N_4004);
xnor U4566 (N_4566,N_4468,N_4341);
and U4567 (N_4567,N_4082,N_4247);
nand U4568 (N_4568,N_4426,N_4102);
and U4569 (N_4569,N_4367,N_4063);
nor U4570 (N_4570,N_4481,N_4368);
xnor U4571 (N_4571,N_4148,N_4281);
nor U4572 (N_4572,N_4060,N_4335);
nor U4573 (N_4573,N_4489,N_4210);
and U4574 (N_4574,N_4150,N_4436);
nand U4575 (N_4575,N_4453,N_4429);
nor U4576 (N_4576,N_4089,N_4208);
or U4577 (N_4577,N_4461,N_4384);
nor U4578 (N_4578,N_4286,N_4174);
or U4579 (N_4579,N_4080,N_4217);
and U4580 (N_4580,N_4034,N_4257);
and U4581 (N_4581,N_4338,N_4199);
nand U4582 (N_4582,N_4459,N_4202);
or U4583 (N_4583,N_4053,N_4390);
and U4584 (N_4584,N_4129,N_4455);
nand U4585 (N_4585,N_4238,N_4339);
nor U4586 (N_4586,N_4029,N_4330);
nand U4587 (N_4587,N_4291,N_4204);
xnor U4588 (N_4588,N_4466,N_4472);
nand U4589 (N_4589,N_4031,N_4454);
nor U4590 (N_4590,N_4253,N_4103);
and U4591 (N_4591,N_4023,N_4172);
nand U4592 (N_4592,N_4090,N_4186);
and U4593 (N_4593,N_4119,N_4276);
xor U4594 (N_4594,N_4270,N_4215);
xor U4595 (N_4595,N_4486,N_4136);
nand U4596 (N_4596,N_4268,N_4423);
nor U4597 (N_4597,N_4362,N_4166);
xor U4598 (N_4598,N_4221,N_4087);
xnor U4599 (N_4599,N_4252,N_4201);
and U4600 (N_4600,N_4282,N_4084);
nand U4601 (N_4601,N_4142,N_4349);
nor U4602 (N_4602,N_4231,N_4414);
and U4603 (N_4603,N_4171,N_4462);
nand U4604 (N_4604,N_4274,N_4449);
and U4605 (N_4605,N_4451,N_4195);
or U4606 (N_4606,N_4440,N_4159);
xor U4607 (N_4607,N_4124,N_4073);
nor U4608 (N_4608,N_4036,N_4260);
or U4609 (N_4609,N_4399,N_4125);
nand U4610 (N_4610,N_4027,N_4385);
nand U4611 (N_4611,N_4323,N_4207);
xnor U4612 (N_4612,N_4214,N_4483);
nand U4613 (N_4613,N_4340,N_4152);
nand U4614 (N_4614,N_4393,N_4091);
or U4615 (N_4615,N_4044,N_4248);
and U4616 (N_4616,N_4075,N_4445);
nand U4617 (N_4617,N_4283,N_4485);
nor U4618 (N_4618,N_4380,N_4265);
and U4619 (N_4619,N_4458,N_4061);
nand U4620 (N_4620,N_4413,N_4024);
nor U4621 (N_4621,N_4351,N_4377);
and U4622 (N_4622,N_4246,N_4342);
or U4623 (N_4623,N_4055,N_4379);
and U4624 (N_4624,N_4181,N_4465);
nand U4625 (N_4625,N_4395,N_4072);
nor U4626 (N_4626,N_4032,N_4289);
nand U4627 (N_4627,N_4212,N_4016);
or U4628 (N_4628,N_4085,N_4167);
nor U4629 (N_4629,N_4109,N_4192);
or U4630 (N_4630,N_4287,N_4127);
or U4631 (N_4631,N_4115,N_4198);
nand U4632 (N_4632,N_4037,N_4224);
nand U4633 (N_4633,N_4290,N_4318);
nor U4634 (N_4634,N_4003,N_4376);
or U4635 (N_4635,N_4083,N_4143);
xor U4636 (N_4636,N_4098,N_4095);
nor U4637 (N_4637,N_4374,N_4194);
nor U4638 (N_4638,N_4052,N_4417);
and U4639 (N_4639,N_4187,N_4251);
or U4640 (N_4640,N_4494,N_4378);
nor U4641 (N_4641,N_4386,N_4039);
and U4642 (N_4642,N_4229,N_4406);
nor U4643 (N_4643,N_4371,N_4331);
nor U4644 (N_4644,N_4424,N_4471);
nand U4645 (N_4645,N_4469,N_4012);
and U4646 (N_4646,N_4321,N_4068);
xor U4647 (N_4647,N_4430,N_4153);
xor U4648 (N_4648,N_4308,N_4038);
nor U4649 (N_4649,N_4365,N_4196);
and U4650 (N_4650,N_4470,N_4114);
nor U4651 (N_4651,N_4266,N_4300);
nor U4652 (N_4652,N_4104,N_4175);
or U4653 (N_4653,N_4057,N_4030);
and U4654 (N_4654,N_4347,N_4372);
xor U4655 (N_4655,N_4316,N_4293);
and U4656 (N_4656,N_4421,N_4069);
or U4657 (N_4657,N_4157,N_4482);
nor U4658 (N_4658,N_4358,N_4277);
nand U4659 (N_4659,N_4005,N_4314);
nand U4660 (N_4660,N_4357,N_4387);
and U4661 (N_4661,N_4398,N_4137);
xnor U4662 (N_4662,N_4191,N_4118);
xnor U4663 (N_4663,N_4346,N_4161);
nand U4664 (N_4664,N_4213,N_4225);
nor U4665 (N_4665,N_4404,N_4101);
xnor U4666 (N_4666,N_4139,N_4099);
and U4667 (N_4667,N_4438,N_4250);
xor U4668 (N_4668,N_4241,N_4363);
nor U4669 (N_4669,N_4310,N_4233);
xor U4670 (N_4670,N_4452,N_4107);
nand U4671 (N_4671,N_4001,N_4434);
xnor U4672 (N_4672,N_4388,N_4326);
or U4673 (N_4673,N_4336,N_4348);
or U4674 (N_4674,N_4297,N_4015);
nand U4675 (N_4675,N_4071,N_4435);
and U4676 (N_4676,N_4442,N_4132);
or U4677 (N_4677,N_4261,N_4267);
xor U4678 (N_4678,N_4369,N_4477);
nand U4679 (N_4679,N_4474,N_4375);
nand U4680 (N_4680,N_4325,N_4065);
nor U4681 (N_4681,N_4394,N_4444);
or U4682 (N_4682,N_4475,N_4299);
nand U4683 (N_4683,N_4484,N_4499);
nand U4684 (N_4684,N_4242,N_4066);
nand U4685 (N_4685,N_4273,N_4062);
nor U4686 (N_4686,N_4344,N_4058);
or U4687 (N_4687,N_4006,N_4049);
xnor U4688 (N_4688,N_4145,N_4322);
or U4689 (N_4689,N_4163,N_4177);
nand U4690 (N_4690,N_4076,N_4422);
nand U4691 (N_4691,N_4490,N_4478);
or U4692 (N_4692,N_4302,N_4258);
nor U4693 (N_4693,N_4350,N_4240);
nand U4694 (N_4694,N_4400,N_4324);
nor U4695 (N_4695,N_4264,N_4183);
and U4696 (N_4696,N_4464,N_4409);
nand U4697 (N_4697,N_4189,N_4309);
xor U4698 (N_4698,N_4190,N_4495);
xnor U4699 (N_4699,N_4188,N_4244);
nor U4700 (N_4700,N_4111,N_4078);
and U4701 (N_4701,N_4391,N_4292);
nor U4702 (N_4702,N_4431,N_4135);
nor U4703 (N_4703,N_4407,N_4223);
nor U4704 (N_4704,N_4184,N_4128);
nand U4705 (N_4705,N_4361,N_4439);
or U4706 (N_4706,N_4164,N_4249);
or U4707 (N_4707,N_4301,N_4113);
nand U4708 (N_4708,N_4008,N_4354);
nand U4709 (N_4709,N_4463,N_4493);
and U4710 (N_4710,N_4035,N_4412);
or U4711 (N_4711,N_4307,N_4168);
xnor U4712 (N_4712,N_4130,N_4473);
nor U4713 (N_4713,N_4480,N_4041);
and U4714 (N_4714,N_4364,N_4131);
or U4715 (N_4715,N_4256,N_4226);
and U4716 (N_4716,N_4025,N_4230);
and U4717 (N_4717,N_4456,N_4381);
nand U4718 (N_4718,N_4160,N_4018);
nor U4719 (N_4719,N_4497,N_4428);
or U4720 (N_4720,N_4311,N_4427);
xnor U4721 (N_4721,N_4312,N_4329);
nor U4722 (N_4722,N_4487,N_4239);
and U4723 (N_4723,N_4026,N_4051);
xor U4724 (N_4724,N_4000,N_4333);
nor U4725 (N_4725,N_4216,N_4203);
xor U4726 (N_4726,N_4278,N_4419);
and U4727 (N_4727,N_4156,N_4317);
and U4728 (N_4728,N_4433,N_4279);
nor U4729 (N_4729,N_4040,N_4178);
xnor U4730 (N_4730,N_4097,N_4218);
and U4731 (N_4731,N_4447,N_4042);
or U4732 (N_4732,N_4360,N_4158);
or U4733 (N_4733,N_4397,N_4079);
and U4734 (N_4734,N_4382,N_4320);
and U4735 (N_4735,N_4303,N_4094);
nor U4736 (N_4736,N_4074,N_4255);
nor U4737 (N_4737,N_4009,N_4046);
or U4738 (N_4738,N_4370,N_4077);
nand U4739 (N_4739,N_4328,N_4313);
xnor U4740 (N_4740,N_4337,N_4305);
nand U4741 (N_4741,N_4197,N_4105);
nor U4742 (N_4742,N_4496,N_4149);
and U4743 (N_4743,N_4327,N_4093);
nand U4744 (N_4744,N_4162,N_4002);
nor U4745 (N_4745,N_4126,N_4179);
nand U4746 (N_4746,N_4045,N_4180);
nand U4747 (N_4747,N_4405,N_4450);
nand U4748 (N_4748,N_4121,N_4116);
and U4749 (N_4749,N_4460,N_4056);
xnor U4750 (N_4750,N_4414,N_4271);
xnor U4751 (N_4751,N_4320,N_4491);
and U4752 (N_4752,N_4189,N_4123);
nor U4753 (N_4753,N_4301,N_4166);
or U4754 (N_4754,N_4067,N_4224);
or U4755 (N_4755,N_4204,N_4132);
nand U4756 (N_4756,N_4325,N_4257);
and U4757 (N_4757,N_4259,N_4071);
nand U4758 (N_4758,N_4470,N_4318);
nand U4759 (N_4759,N_4235,N_4173);
nor U4760 (N_4760,N_4138,N_4063);
or U4761 (N_4761,N_4017,N_4012);
nor U4762 (N_4762,N_4378,N_4295);
and U4763 (N_4763,N_4214,N_4393);
nor U4764 (N_4764,N_4128,N_4401);
nor U4765 (N_4765,N_4347,N_4161);
xor U4766 (N_4766,N_4176,N_4495);
nor U4767 (N_4767,N_4179,N_4286);
nand U4768 (N_4768,N_4162,N_4096);
xor U4769 (N_4769,N_4263,N_4466);
and U4770 (N_4770,N_4441,N_4357);
or U4771 (N_4771,N_4417,N_4447);
or U4772 (N_4772,N_4039,N_4478);
xor U4773 (N_4773,N_4004,N_4064);
xor U4774 (N_4774,N_4197,N_4249);
nand U4775 (N_4775,N_4234,N_4378);
or U4776 (N_4776,N_4237,N_4393);
and U4777 (N_4777,N_4261,N_4079);
nor U4778 (N_4778,N_4128,N_4437);
or U4779 (N_4779,N_4464,N_4330);
xor U4780 (N_4780,N_4327,N_4010);
xor U4781 (N_4781,N_4281,N_4347);
nand U4782 (N_4782,N_4411,N_4063);
or U4783 (N_4783,N_4169,N_4242);
xnor U4784 (N_4784,N_4182,N_4420);
nand U4785 (N_4785,N_4383,N_4452);
nand U4786 (N_4786,N_4181,N_4421);
xor U4787 (N_4787,N_4322,N_4085);
nand U4788 (N_4788,N_4053,N_4024);
and U4789 (N_4789,N_4169,N_4112);
or U4790 (N_4790,N_4375,N_4397);
nand U4791 (N_4791,N_4036,N_4422);
nor U4792 (N_4792,N_4055,N_4077);
or U4793 (N_4793,N_4028,N_4210);
nor U4794 (N_4794,N_4415,N_4278);
and U4795 (N_4795,N_4327,N_4461);
nor U4796 (N_4796,N_4283,N_4143);
nor U4797 (N_4797,N_4151,N_4060);
or U4798 (N_4798,N_4091,N_4029);
xnor U4799 (N_4799,N_4077,N_4326);
xnor U4800 (N_4800,N_4300,N_4133);
nand U4801 (N_4801,N_4475,N_4291);
nor U4802 (N_4802,N_4261,N_4453);
xor U4803 (N_4803,N_4422,N_4436);
nand U4804 (N_4804,N_4034,N_4316);
xor U4805 (N_4805,N_4456,N_4386);
or U4806 (N_4806,N_4091,N_4049);
and U4807 (N_4807,N_4204,N_4243);
nand U4808 (N_4808,N_4368,N_4115);
or U4809 (N_4809,N_4110,N_4082);
nor U4810 (N_4810,N_4100,N_4034);
or U4811 (N_4811,N_4176,N_4284);
nor U4812 (N_4812,N_4240,N_4182);
nand U4813 (N_4813,N_4264,N_4445);
and U4814 (N_4814,N_4244,N_4314);
or U4815 (N_4815,N_4096,N_4354);
nand U4816 (N_4816,N_4024,N_4044);
nor U4817 (N_4817,N_4420,N_4220);
or U4818 (N_4818,N_4439,N_4101);
and U4819 (N_4819,N_4073,N_4011);
or U4820 (N_4820,N_4088,N_4014);
and U4821 (N_4821,N_4281,N_4025);
and U4822 (N_4822,N_4055,N_4113);
nor U4823 (N_4823,N_4437,N_4326);
nand U4824 (N_4824,N_4260,N_4142);
nand U4825 (N_4825,N_4174,N_4096);
nand U4826 (N_4826,N_4180,N_4399);
and U4827 (N_4827,N_4042,N_4091);
xnor U4828 (N_4828,N_4193,N_4259);
xnor U4829 (N_4829,N_4184,N_4118);
xnor U4830 (N_4830,N_4047,N_4421);
and U4831 (N_4831,N_4461,N_4342);
nor U4832 (N_4832,N_4366,N_4165);
nor U4833 (N_4833,N_4442,N_4257);
nor U4834 (N_4834,N_4047,N_4059);
nor U4835 (N_4835,N_4052,N_4438);
xnor U4836 (N_4836,N_4373,N_4462);
xnor U4837 (N_4837,N_4395,N_4201);
nor U4838 (N_4838,N_4475,N_4002);
nor U4839 (N_4839,N_4322,N_4471);
nand U4840 (N_4840,N_4075,N_4310);
nand U4841 (N_4841,N_4241,N_4235);
xnor U4842 (N_4842,N_4452,N_4149);
nor U4843 (N_4843,N_4048,N_4208);
and U4844 (N_4844,N_4245,N_4086);
nor U4845 (N_4845,N_4058,N_4207);
and U4846 (N_4846,N_4447,N_4037);
xor U4847 (N_4847,N_4065,N_4029);
nand U4848 (N_4848,N_4191,N_4122);
nand U4849 (N_4849,N_4472,N_4250);
or U4850 (N_4850,N_4258,N_4287);
and U4851 (N_4851,N_4341,N_4316);
and U4852 (N_4852,N_4217,N_4289);
or U4853 (N_4853,N_4020,N_4325);
or U4854 (N_4854,N_4400,N_4053);
and U4855 (N_4855,N_4405,N_4134);
nand U4856 (N_4856,N_4198,N_4206);
xnor U4857 (N_4857,N_4263,N_4300);
or U4858 (N_4858,N_4121,N_4417);
or U4859 (N_4859,N_4396,N_4043);
xnor U4860 (N_4860,N_4243,N_4036);
xor U4861 (N_4861,N_4456,N_4295);
or U4862 (N_4862,N_4213,N_4208);
or U4863 (N_4863,N_4339,N_4333);
nor U4864 (N_4864,N_4126,N_4263);
xnor U4865 (N_4865,N_4063,N_4498);
and U4866 (N_4866,N_4425,N_4472);
or U4867 (N_4867,N_4438,N_4475);
and U4868 (N_4868,N_4280,N_4451);
and U4869 (N_4869,N_4187,N_4017);
nand U4870 (N_4870,N_4315,N_4479);
nor U4871 (N_4871,N_4212,N_4325);
and U4872 (N_4872,N_4401,N_4435);
nor U4873 (N_4873,N_4387,N_4035);
and U4874 (N_4874,N_4498,N_4354);
or U4875 (N_4875,N_4228,N_4314);
and U4876 (N_4876,N_4457,N_4001);
or U4877 (N_4877,N_4384,N_4264);
nand U4878 (N_4878,N_4314,N_4100);
nand U4879 (N_4879,N_4018,N_4098);
nor U4880 (N_4880,N_4479,N_4155);
nand U4881 (N_4881,N_4219,N_4032);
nand U4882 (N_4882,N_4476,N_4015);
or U4883 (N_4883,N_4342,N_4361);
xor U4884 (N_4884,N_4309,N_4094);
and U4885 (N_4885,N_4415,N_4204);
xnor U4886 (N_4886,N_4032,N_4342);
xnor U4887 (N_4887,N_4315,N_4476);
nor U4888 (N_4888,N_4350,N_4209);
nand U4889 (N_4889,N_4181,N_4106);
nand U4890 (N_4890,N_4242,N_4389);
nand U4891 (N_4891,N_4461,N_4435);
xor U4892 (N_4892,N_4436,N_4082);
nor U4893 (N_4893,N_4393,N_4398);
xor U4894 (N_4894,N_4263,N_4018);
nor U4895 (N_4895,N_4430,N_4187);
nor U4896 (N_4896,N_4223,N_4409);
nand U4897 (N_4897,N_4140,N_4398);
or U4898 (N_4898,N_4360,N_4124);
nor U4899 (N_4899,N_4450,N_4375);
nand U4900 (N_4900,N_4326,N_4346);
and U4901 (N_4901,N_4047,N_4191);
nor U4902 (N_4902,N_4219,N_4272);
nand U4903 (N_4903,N_4339,N_4466);
xnor U4904 (N_4904,N_4032,N_4142);
or U4905 (N_4905,N_4369,N_4211);
nor U4906 (N_4906,N_4241,N_4269);
or U4907 (N_4907,N_4019,N_4121);
or U4908 (N_4908,N_4056,N_4410);
nor U4909 (N_4909,N_4266,N_4481);
nor U4910 (N_4910,N_4182,N_4424);
nor U4911 (N_4911,N_4415,N_4123);
nand U4912 (N_4912,N_4275,N_4418);
and U4913 (N_4913,N_4046,N_4349);
xnor U4914 (N_4914,N_4293,N_4330);
or U4915 (N_4915,N_4065,N_4313);
nand U4916 (N_4916,N_4118,N_4433);
xor U4917 (N_4917,N_4384,N_4101);
nor U4918 (N_4918,N_4319,N_4170);
nand U4919 (N_4919,N_4276,N_4044);
xnor U4920 (N_4920,N_4357,N_4434);
and U4921 (N_4921,N_4017,N_4402);
and U4922 (N_4922,N_4209,N_4086);
or U4923 (N_4923,N_4204,N_4091);
or U4924 (N_4924,N_4494,N_4128);
or U4925 (N_4925,N_4132,N_4393);
xor U4926 (N_4926,N_4026,N_4419);
nand U4927 (N_4927,N_4207,N_4447);
or U4928 (N_4928,N_4071,N_4310);
or U4929 (N_4929,N_4401,N_4397);
nand U4930 (N_4930,N_4374,N_4281);
nand U4931 (N_4931,N_4472,N_4164);
xor U4932 (N_4932,N_4122,N_4368);
nor U4933 (N_4933,N_4016,N_4132);
xor U4934 (N_4934,N_4442,N_4271);
nand U4935 (N_4935,N_4026,N_4435);
and U4936 (N_4936,N_4464,N_4110);
xnor U4937 (N_4937,N_4239,N_4126);
nor U4938 (N_4938,N_4462,N_4114);
or U4939 (N_4939,N_4298,N_4122);
and U4940 (N_4940,N_4358,N_4022);
xor U4941 (N_4941,N_4329,N_4094);
xor U4942 (N_4942,N_4406,N_4172);
nor U4943 (N_4943,N_4466,N_4015);
nand U4944 (N_4944,N_4413,N_4331);
and U4945 (N_4945,N_4386,N_4387);
and U4946 (N_4946,N_4467,N_4404);
or U4947 (N_4947,N_4082,N_4460);
or U4948 (N_4948,N_4115,N_4140);
nand U4949 (N_4949,N_4185,N_4327);
nand U4950 (N_4950,N_4048,N_4191);
xnor U4951 (N_4951,N_4340,N_4156);
nor U4952 (N_4952,N_4441,N_4431);
nand U4953 (N_4953,N_4234,N_4321);
nand U4954 (N_4954,N_4496,N_4024);
nand U4955 (N_4955,N_4408,N_4192);
xnor U4956 (N_4956,N_4369,N_4484);
nor U4957 (N_4957,N_4172,N_4146);
xor U4958 (N_4958,N_4432,N_4128);
nand U4959 (N_4959,N_4232,N_4109);
or U4960 (N_4960,N_4287,N_4037);
xor U4961 (N_4961,N_4041,N_4156);
and U4962 (N_4962,N_4236,N_4225);
nor U4963 (N_4963,N_4154,N_4389);
and U4964 (N_4964,N_4140,N_4263);
xnor U4965 (N_4965,N_4217,N_4074);
or U4966 (N_4966,N_4261,N_4135);
nor U4967 (N_4967,N_4188,N_4053);
nand U4968 (N_4968,N_4288,N_4286);
or U4969 (N_4969,N_4196,N_4464);
nor U4970 (N_4970,N_4498,N_4177);
nor U4971 (N_4971,N_4463,N_4153);
and U4972 (N_4972,N_4202,N_4236);
xor U4973 (N_4973,N_4002,N_4318);
nand U4974 (N_4974,N_4317,N_4382);
or U4975 (N_4975,N_4437,N_4444);
nor U4976 (N_4976,N_4022,N_4275);
and U4977 (N_4977,N_4333,N_4480);
or U4978 (N_4978,N_4344,N_4462);
xor U4979 (N_4979,N_4354,N_4279);
nand U4980 (N_4980,N_4251,N_4391);
and U4981 (N_4981,N_4132,N_4008);
nor U4982 (N_4982,N_4153,N_4022);
nor U4983 (N_4983,N_4012,N_4243);
or U4984 (N_4984,N_4076,N_4135);
xor U4985 (N_4985,N_4451,N_4033);
or U4986 (N_4986,N_4087,N_4147);
or U4987 (N_4987,N_4026,N_4288);
nand U4988 (N_4988,N_4184,N_4229);
nand U4989 (N_4989,N_4086,N_4014);
and U4990 (N_4990,N_4041,N_4007);
and U4991 (N_4991,N_4437,N_4166);
nor U4992 (N_4992,N_4415,N_4343);
nand U4993 (N_4993,N_4495,N_4356);
xnor U4994 (N_4994,N_4055,N_4464);
nor U4995 (N_4995,N_4161,N_4488);
or U4996 (N_4996,N_4057,N_4032);
nand U4997 (N_4997,N_4094,N_4175);
or U4998 (N_4998,N_4128,N_4322);
xor U4999 (N_4999,N_4430,N_4272);
nand U5000 (N_5000,N_4903,N_4933);
xor U5001 (N_5001,N_4857,N_4677);
xor U5002 (N_5002,N_4734,N_4944);
nand U5003 (N_5003,N_4748,N_4629);
xor U5004 (N_5004,N_4625,N_4759);
and U5005 (N_5005,N_4988,N_4541);
nor U5006 (N_5006,N_4926,N_4714);
and U5007 (N_5007,N_4647,N_4543);
or U5008 (N_5008,N_4695,N_4994);
nand U5009 (N_5009,N_4614,N_4902);
and U5010 (N_5010,N_4630,N_4579);
nand U5011 (N_5011,N_4825,N_4712);
or U5012 (N_5012,N_4648,N_4869);
nor U5013 (N_5013,N_4989,N_4990);
or U5014 (N_5014,N_4900,N_4584);
nor U5015 (N_5015,N_4941,N_4892);
nand U5016 (N_5016,N_4899,N_4793);
or U5017 (N_5017,N_4942,N_4826);
and U5018 (N_5018,N_4688,N_4963);
nand U5019 (N_5019,N_4744,N_4707);
and U5020 (N_5020,N_4583,N_4645);
xor U5021 (N_5021,N_4795,N_4739);
nand U5022 (N_5022,N_4884,N_4682);
or U5023 (N_5023,N_4701,N_4929);
or U5024 (N_5024,N_4567,N_4711);
or U5025 (N_5025,N_4724,N_4580);
xor U5026 (N_5026,N_4937,N_4849);
nor U5027 (N_5027,N_4755,N_4607);
nand U5028 (N_5028,N_4888,N_4626);
nor U5029 (N_5029,N_4841,N_4732);
nor U5030 (N_5030,N_4861,N_4608);
nor U5031 (N_5031,N_4754,N_4635);
xor U5032 (N_5032,N_4954,N_4997);
nor U5033 (N_5033,N_4823,N_4995);
nor U5034 (N_5034,N_4896,N_4502);
or U5035 (N_5035,N_4500,N_4773);
and U5036 (N_5036,N_4750,N_4805);
or U5037 (N_5037,N_4588,N_4611);
xnor U5038 (N_5038,N_4906,N_4642);
xor U5039 (N_5039,N_4723,N_4603);
or U5040 (N_5040,N_4980,N_4915);
xor U5041 (N_5041,N_4779,N_4991);
xor U5042 (N_5042,N_4575,N_4831);
and U5043 (N_5043,N_4889,N_4545);
nand U5044 (N_5044,N_4563,N_4881);
nand U5045 (N_5045,N_4919,N_4939);
nand U5046 (N_5046,N_4658,N_4961);
nor U5047 (N_5047,N_4532,N_4753);
nor U5048 (N_5048,N_4751,N_4801);
nand U5049 (N_5049,N_4736,N_4574);
nand U5050 (N_5050,N_4761,N_4566);
nand U5051 (N_5051,N_4927,N_4993);
nand U5052 (N_5052,N_4662,N_4572);
and U5053 (N_5053,N_4968,N_4974);
nor U5054 (N_5054,N_4894,N_4747);
xor U5055 (N_5055,N_4887,N_4778);
and U5056 (N_5056,N_4581,N_4769);
xor U5057 (N_5057,N_4912,N_4535);
nor U5058 (N_5058,N_4719,N_4897);
and U5059 (N_5059,N_4838,N_4726);
nor U5060 (N_5060,N_4780,N_4704);
nor U5061 (N_5061,N_4556,N_4890);
and U5062 (N_5062,N_4800,N_4512);
nor U5063 (N_5063,N_4516,N_4537);
nand U5064 (N_5064,N_4871,N_4848);
nand U5065 (N_5065,N_4882,N_4758);
or U5066 (N_5066,N_4945,N_4519);
nor U5067 (N_5067,N_4710,N_4760);
nor U5068 (N_5068,N_4864,N_4696);
xnor U5069 (N_5069,N_4713,N_4598);
and U5070 (N_5070,N_4716,N_4576);
and U5071 (N_5071,N_4507,N_4699);
and U5072 (N_5072,N_4967,N_4534);
nor U5073 (N_5073,N_4810,N_4615);
and U5074 (N_5074,N_4797,N_4819);
xor U5075 (N_5075,N_4785,N_4975);
xor U5076 (N_5076,N_4922,N_4782);
or U5077 (N_5077,N_4947,N_4846);
and U5078 (N_5078,N_4757,N_4943);
and U5079 (N_5079,N_4542,N_4589);
or U5080 (N_5080,N_4982,N_4987);
nand U5081 (N_5081,N_4544,N_4513);
or U5082 (N_5082,N_4876,N_4664);
xnor U5083 (N_5083,N_4686,N_4908);
and U5084 (N_5084,N_4594,N_4597);
nand U5085 (N_5085,N_4646,N_4845);
nor U5086 (N_5086,N_4621,N_4665);
xnor U5087 (N_5087,N_4957,N_4955);
xor U5088 (N_5088,N_4986,N_4693);
nor U5089 (N_5089,N_4705,N_4798);
nor U5090 (N_5090,N_4738,N_4730);
and U5091 (N_5091,N_4632,N_4840);
and U5092 (N_5092,N_4764,N_4875);
nand U5093 (N_5093,N_4533,N_4930);
or U5094 (N_5094,N_4909,N_4850);
or U5095 (N_5095,N_4873,N_4827);
or U5096 (N_5096,N_4820,N_4552);
nand U5097 (N_5097,N_4959,N_4851);
nor U5098 (N_5098,N_4934,N_4700);
xnor U5099 (N_5099,N_4839,N_4938);
nor U5100 (N_5100,N_4853,N_4940);
nand U5101 (N_5101,N_4517,N_4879);
xnor U5102 (N_5102,N_4668,N_4860);
or U5103 (N_5103,N_4911,N_4565);
or U5104 (N_5104,N_4692,N_4680);
nor U5105 (N_5105,N_4546,N_4774);
nand U5106 (N_5106,N_4679,N_4643);
xnor U5107 (N_5107,N_4816,N_4654);
xor U5108 (N_5108,N_4573,N_4766);
xor U5109 (N_5109,N_4592,N_4554);
nor U5110 (N_5110,N_4717,N_4807);
nand U5111 (N_5111,N_4706,N_4638);
xnor U5112 (N_5112,N_4746,N_4983);
nand U5113 (N_5113,N_4880,N_4960);
xnor U5114 (N_5114,N_4687,N_4708);
and U5115 (N_5115,N_4756,N_4950);
xor U5116 (N_5116,N_4557,N_4669);
nor U5117 (N_5117,N_4878,N_4972);
nand U5118 (N_5118,N_4952,N_4728);
nand U5119 (N_5119,N_4866,N_4539);
xnor U5120 (N_5120,N_4858,N_4657);
or U5121 (N_5121,N_4854,N_4837);
and U5122 (N_5122,N_4582,N_4538);
and U5123 (N_5123,N_4661,N_4777);
xor U5124 (N_5124,N_4787,N_4653);
xor U5125 (N_5125,N_4735,N_4762);
nor U5126 (N_5126,N_4676,N_4709);
nand U5127 (N_5127,N_4577,N_4720);
xnor U5128 (N_5128,N_4783,N_4770);
nand U5129 (N_5129,N_4685,N_4616);
nand U5130 (N_5130,N_4949,N_4935);
xor U5131 (N_5131,N_4794,N_4652);
nand U5132 (N_5132,N_4733,N_4920);
nor U5133 (N_5133,N_4969,N_4796);
or U5134 (N_5134,N_4691,N_4548);
xor U5135 (N_5135,N_4844,N_4872);
nor U5136 (N_5136,N_4536,N_4637);
and U5137 (N_5137,N_4984,N_4596);
nor U5138 (N_5138,N_4870,N_4867);
or U5139 (N_5139,N_4765,N_4893);
or U5140 (N_5140,N_4530,N_4511);
nand U5141 (N_5141,N_4962,N_4979);
xor U5142 (N_5142,N_4956,N_4784);
or U5143 (N_5143,N_4886,N_4815);
nor U5144 (N_5144,N_4569,N_4528);
nand U5145 (N_5145,N_4606,N_4558);
xnor U5146 (N_5146,N_4649,N_4817);
and U5147 (N_5147,N_4768,N_4865);
nor U5148 (N_5148,N_4775,N_4981);
and U5149 (N_5149,N_4731,N_4718);
xor U5150 (N_5150,N_4602,N_4924);
and U5151 (N_5151,N_4821,N_4996);
and U5152 (N_5152,N_4802,N_4901);
xor U5153 (N_5153,N_4593,N_4612);
nand U5154 (N_5154,N_4812,N_4727);
nor U5155 (N_5155,N_4948,N_4740);
and U5156 (N_5156,N_4958,N_4828);
nand U5157 (N_5157,N_4623,N_4634);
nand U5158 (N_5158,N_4540,N_4971);
and U5159 (N_5159,N_4789,N_4504);
nand U5160 (N_5160,N_4697,N_4913);
nand U5161 (N_5161,N_4619,N_4862);
nor U5162 (N_5162,N_4604,N_4650);
nand U5163 (N_5163,N_4560,N_4752);
xor U5164 (N_5164,N_4521,N_4928);
nor U5165 (N_5165,N_4824,N_4618);
nor U5166 (N_5166,N_4885,N_4660);
nor U5167 (N_5167,N_4586,N_4681);
nor U5168 (N_5168,N_4672,N_4745);
and U5169 (N_5169,N_4587,N_4836);
and U5170 (N_5170,N_4620,N_4855);
nor U5171 (N_5171,N_4628,N_4624);
or U5172 (N_5172,N_4559,N_4741);
xor U5173 (N_5173,N_4946,N_4561);
nor U5174 (N_5174,N_4992,N_4999);
or U5175 (N_5175,N_4523,N_4767);
or U5176 (N_5176,N_4891,N_4508);
and U5177 (N_5177,N_4703,N_4804);
xor U5178 (N_5178,N_4639,N_4527);
and U5179 (N_5179,N_4631,N_4898);
nor U5180 (N_5180,N_4863,N_4842);
xor U5181 (N_5181,N_4830,N_4847);
and U5182 (N_5182,N_4690,N_4595);
nand U5183 (N_5183,N_4932,N_4931);
xor U5184 (N_5184,N_4781,N_4918);
and U5185 (N_5185,N_4613,N_4910);
xor U5186 (N_5186,N_4667,N_4564);
nand U5187 (N_5187,N_4689,N_4834);
or U5188 (N_5188,N_4683,N_4678);
nand U5189 (N_5189,N_4791,N_4788);
xnor U5190 (N_5190,N_4663,N_4524);
nand U5191 (N_5191,N_4749,N_4822);
xor U5192 (N_5192,N_4671,N_4674);
and U5193 (N_5193,N_4998,N_4585);
or U5194 (N_5194,N_4923,N_4833);
or U5195 (N_5195,N_4953,N_4636);
xnor U5196 (N_5196,N_4895,N_4790);
nand U5197 (N_5197,N_4973,N_4609);
and U5198 (N_5198,N_4786,N_4925);
and U5199 (N_5199,N_4905,N_4951);
and U5200 (N_5200,N_4976,N_4529);
xnor U5201 (N_5201,N_4916,N_4852);
and U5202 (N_5202,N_4966,N_4673);
nor U5203 (N_5203,N_4694,N_4809);
nor U5204 (N_5204,N_4698,N_4506);
xnor U5205 (N_5205,N_4715,N_4549);
nand U5206 (N_5206,N_4666,N_4814);
or U5207 (N_5207,N_4531,N_4684);
nand U5208 (N_5208,N_4551,N_4868);
xor U5209 (N_5209,N_4562,N_4725);
xor U5210 (N_5210,N_4675,N_4729);
xnor U5211 (N_5211,N_4722,N_4644);
nand U5212 (N_5212,N_4525,N_4550);
or U5213 (N_5213,N_4590,N_4829);
nand U5214 (N_5214,N_4832,N_4806);
xnor U5215 (N_5215,N_4743,N_4856);
and U5216 (N_5216,N_4568,N_4601);
xor U5217 (N_5217,N_4985,N_4803);
nor U5218 (N_5218,N_4883,N_4904);
nor U5219 (N_5219,N_4514,N_4763);
and U5220 (N_5220,N_4617,N_4917);
nand U5221 (N_5221,N_4651,N_4570);
and U5222 (N_5222,N_4509,N_4771);
nor U5223 (N_5223,N_4578,N_4600);
nand U5224 (N_5224,N_4505,N_4811);
and U5225 (N_5225,N_4605,N_4877);
or U5226 (N_5226,N_4978,N_4522);
or U5227 (N_5227,N_4622,N_4591);
xor U5228 (N_5228,N_4977,N_4518);
nor U5229 (N_5229,N_4808,N_4555);
nor U5230 (N_5230,N_4641,N_4859);
or U5231 (N_5231,N_4702,N_4659);
or U5232 (N_5232,N_4510,N_4610);
or U5233 (N_5233,N_4627,N_4599);
and U5234 (N_5234,N_4640,N_4843);
nand U5235 (N_5235,N_4520,N_4526);
and U5236 (N_5236,N_4964,N_4655);
or U5237 (N_5237,N_4936,N_4874);
xor U5238 (N_5238,N_4813,N_4553);
nor U5239 (N_5239,N_4970,N_4776);
and U5240 (N_5240,N_4515,N_4965);
nor U5241 (N_5241,N_4921,N_4721);
and U5242 (N_5242,N_4670,N_4914);
nand U5243 (N_5243,N_4835,N_4799);
nand U5244 (N_5244,N_4742,N_4656);
nor U5245 (N_5245,N_4501,N_4792);
and U5246 (N_5246,N_4633,N_4503);
and U5247 (N_5247,N_4571,N_4547);
nor U5248 (N_5248,N_4818,N_4737);
nor U5249 (N_5249,N_4772,N_4907);
and U5250 (N_5250,N_4748,N_4822);
nor U5251 (N_5251,N_4686,N_4860);
xor U5252 (N_5252,N_4555,N_4856);
xnor U5253 (N_5253,N_4875,N_4620);
or U5254 (N_5254,N_4532,N_4591);
and U5255 (N_5255,N_4875,N_4997);
and U5256 (N_5256,N_4576,N_4810);
xor U5257 (N_5257,N_4829,N_4917);
nand U5258 (N_5258,N_4527,N_4582);
or U5259 (N_5259,N_4935,N_4613);
nand U5260 (N_5260,N_4705,N_4963);
nor U5261 (N_5261,N_4514,N_4974);
and U5262 (N_5262,N_4882,N_4871);
nand U5263 (N_5263,N_4891,N_4754);
nand U5264 (N_5264,N_4786,N_4651);
and U5265 (N_5265,N_4552,N_4533);
nand U5266 (N_5266,N_4585,N_4915);
xnor U5267 (N_5267,N_4944,N_4546);
or U5268 (N_5268,N_4516,N_4870);
nand U5269 (N_5269,N_4741,N_4981);
nor U5270 (N_5270,N_4967,N_4540);
xnor U5271 (N_5271,N_4888,N_4848);
nand U5272 (N_5272,N_4500,N_4502);
nor U5273 (N_5273,N_4846,N_4697);
nor U5274 (N_5274,N_4740,N_4636);
nor U5275 (N_5275,N_4678,N_4736);
and U5276 (N_5276,N_4646,N_4502);
nor U5277 (N_5277,N_4976,N_4906);
and U5278 (N_5278,N_4846,N_4558);
or U5279 (N_5279,N_4935,N_4993);
or U5280 (N_5280,N_4990,N_4806);
nand U5281 (N_5281,N_4566,N_4522);
xor U5282 (N_5282,N_4616,N_4982);
xnor U5283 (N_5283,N_4567,N_4577);
xor U5284 (N_5284,N_4821,N_4899);
xnor U5285 (N_5285,N_4677,N_4515);
or U5286 (N_5286,N_4679,N_4555);
nor U5287 (N_5287,N_4980,N_4630);
nor U5288 (N_5288,N_4678,N_4925);
or U5289 (N_5289,N_4750,N_4851);
nand U5290 (N_5290,N_4774,N_4591);
and U5291 (N_5291,N_4643,N_4641);
nor U5292 (N_5292,N_4844,N_4782);
nor U5293 (N_5293,N_4918,N_4862);
xnor U5294 (N_5294,N_4649,N_4887);
nand U5295 (N_5295,N_4622,N_4889);
xor U5296 (N_5296,N_4961,N_4941);
nor U5297 (N_5297,N_4844,N_4963);
and U5298 (N_5298,N_4918,N_4875);
or U5299 (N_5299,N_4934,N_4883);
xnor U5300 (N_5300,N_4890,N_4876);
nor U5301 (N_5301,N_4824,N_4693);
and U5302 (N_5302,N_4914,N_4731);
xnor U5303 (N_5303,N_4878,N_4725);
nand U5304 (N_5304,N_4998,N_4921);
and U5305 (N_5305,N_4640,N_4914);
xnor U5306 (N_5306,N_4770,N_4680);
nand U5307 (N_5307,N_4510,N_4783);
or U5308 (N_5308,N_4913,N_4901);
nor U5309 (N_5309,N_4759,N_4950);
and U5310 (N_5310,N_4853,N_4863);
or U5311 (N_5311,N_4678,N_4756);
nor U5312 (N_5312,N_4732,N_4577);
xnor U5313 (N_5313,N_4527,N_4549);
and U5314 (N_5314,N_4528,N_4692);
nor U5315 (N_5315,N_4869,N_4761);
xnor U5316 (N_5316,N_4500,N_4562);
nor U5317 (N_5317,N_4878,N_4686);
and U5318 (N_5318,N_4647,N_4834);
nand U5319 (N_5319,N_4503,N_4768);
xnor U5320 (N_5320,N_4595,N_4809);
nand U5321 (N_5321,N_4561,N_4816);
nand U5322 (N_5322,N_4538,N_4687);
xnor U5323 (N_5323,N_4640,N_4905);
or U5324 (N_5324,N_4834,N_4902);
nand U5325 (N_5325,N_4772,N_4884);
or U5326 (N_5326,N_4525,N_4676);
and U5327 (N_5327,N_4775,N_4529);
nor U5328 (N_5328,N_4995,N_4857);
and U5329 (N_5329,N_4833,N_4552);
nor U5330 (N_5330,N_4962,N_4693);
nor U5331 (N_5331,N_4602,N_4665);
xnor U5332 (N_5332,N_4973,N_4731);
xor U5333 (N_5333,N_4977,N_4507);
and U5334 (N_5334,N_4899,N_4748);
nor U5335 (N_5335,N_4716,N_4991);
or U5336 (N_5336,N_4907,N_4564);
and U5337 (N_5337,N_4843,N_4819);
nor U5338 (N_5338,N_4996,N_4720);
nand U5339 (N_5339,N_4567,N_4531);
or U5340 (N_5340,N_4836,N_4862);
nand U5341 (N_5341,N_4818,N_4580);
nor U5342 (N_5342,N_4624,N_4858);
and U5343 (N_5343,N_4728,N_4615);
and U5344 (N_5344,N_4711,N_4663);
nand U5345 (N_5345,N_4680,N_4777);
nand U5346 (N_5346,N_4940,N_4718);
or U5347 (N_5347,N_4674,N_4693);
nor U5348 (N_5348,N_4699,N_4565);
and U5349 (N_5349,N_4815,N_4758);
nand U5350 (N_5350,N_4501,N_4558);
and U5351 (N_5351,N_4566,N_4717);
xor U5352 (N_5352,N_4848,N_4720);
nor U5353 (N_5353,N_4541,N_4837);
nand U5354 (N_5354,N_4595,N_4796);
or U5355 (N_5355,N_4626,N_4830);
xnor U5356 (N_5356,N_4883,N_4568);
xnor U5357 (N_5357,N_4892,N_4603);
and U5358 (N_5358,N_4564,N_4607);
nand U5359 (N_5359,N_4843,N_4670);
nand U5360 (N_5360,N_4659,N_4557);
nor U5361 (N_5361,N_4680,N_4646);
xor U5362 (N_5362,N_4936,N_4993);
and U5363 (N_5363,N_4869,N_4970);
or U5364 (N_5364,N_4782,N_4699);
xor U5365 (N_5365,N_4552,N_4723);
or U5366 (N_5366,N_4794,N_4589);
xnor U5367 (N_5367,N_4782,N_4959);
and U5368 (N_5368,N_4678,N_4884);
nand U5369 (N_5369,N_4883,N_4774);
nor U5370 (N_5370,N_4741,N_4826);
or U5371 (N_5371,N_4914,N_4589);
nor U5372 (N_5372,N_4583,N_4981);
nand U5373 (N_5373,N_4932,N_4519);
xor U5374 (N_5374,N_4876,N_4815);
and U5375 (N_5375,N_4591,N_4956);
or U5376 (N_5376,N_4916,N_4740);
nand U5377 (N_5377,N_4562,N_4926);
xnor U5378 (N_5378,N_4626,N_4999);
or U5379 (N_5379,N_4729,N_4642);
nor U5380 (N_5380,N_4913,N_4702);
or U5381 (N_5381,N_4610,N_4765);
nor U5382 (N_5382,N_4710,N_4886);
xor U5383 (N_5383,N_4970,N_4794);
xor U5384 (N_5384,N_4679,N_4811);
nand U5385 (N_5385,N_4686,N_4810);
and U5386 (N_5386,N_4724,N_4886);
or U5387 (N_5387,N_4701,N_4555);
or U5388 (N_5388,N_4633,N_4951);
or U5389 (N_5389,N_4690,N_4771);
or U5390 (N_5390,N_4832,N_4941);
nor U5391 (N_5391,N_4656,N_4999);
nor U5392 (N_5392,N_4866,N_4594);
and U5393 (N_5393,N_4765,N_4894);
or U5394 (N_5394,N_4987,N_4709);
xor U5395 (N_5395,N_4950,N_4587);
xor U5396 (N_5396,N_4871,N_4919);
and U5397 (N_5397,N_4865,N_4752);
xnor U5398 (N_5398,N_4618,N_4567);
nor U5399 (N_5399,N_4575,N_4701);
nand U5400 (N_5400,N_4945,N_4725);
xor U5401 (N_5401,N_4860,N_4972);
nand U5402 (N_5402,N_4626,N_4818);
and U5403 (N_5403,N_4767,N_4733);
nor U5404 (N_5404,N_4545,N_4715);
xnor U5405 (N_5405,N_4648,N_4749);
nor U5406 (N_5406,N_4925,N_4647);
xnor U5407 (N_5407,N_4545,N_4989);
xnor U5408 (N_5408,N_4811,N_4872);
or U5409 (N_5409,N_4970,N_4846);
nor U5410 (N_5410,N_4946,N_4804);
or U5411 (N_5411,N_4668,N_4972);
nor U5412 (N_5412,N_4827,N_4874);
and U5413 (N_5413,N_4999,N_4979);
nor U5414 (N_5414,N_4970,N_4972);
and U5415 (N_5415,N_4921,N_4588);
nand U5416 (N_5416,N_4809,N_4929);
xor U5417 (N_5417,N_4616,N_4557);
or U5418 (N_5418,N_4799,N_4911);
and U5419 (N_5419,N_4977,N_4876);
nor U5420 (N_5420,N_4736,N_4740);
nand U5421 (N_5421,N_4519,N_4514);
xor U5422 (N_5422,N_4837,N_4518);
xnor U5423 (N_5423,N_4827,N_4658);
or U5424 (N_5424,N_4722,N_4663);
nor U5425 (N_5425,N_4584,N_4641);
nor U5426 (N_5426,N_4835,N_4760);
xnor U5427 (N_5427,N_4937,N_4622);
nor U5428 (N_5428,N_4811,N_4788);
and U5429 (N_5429,N_4769,N_4602);
and U5430 (N_5430,N_4590,N_4797);
nand U5431 (N_5431,N_4749,N_4656);
nor U5432 (N_5432,N_4992,N_4630);
nor U5433 (N_5433,N_4916,N_4506);
and U5434 (N_5434,N_4588,N_4732);
and U5435 (N_5435,N_4905,N_4661);
xnor U5436 (N_5436,N_4665,N_4623);
xor U5437 (N_5437,N_4928,N_4855);
nand U5438 (N_5438,N_4892,N_4534);
nor U5439 (N_5439,N_4536,N_4595);
nor U5440 (N_5440,N_4861,N_4970);
xor U5441 (N_5441,N_4940,N_4658);
or U5442 (N_5442,N_4605,N_4997);
xor U5443 (N_5443,N_4887,N_4791);
xor U5444 (N_5444,N_4719,N_4765);
or U5445 (N_5445,N_4555,N_4774);
nor U5446 (N_5446,N_4783,N_4678);
or U5447 (N_5447,N_4892,N_4925);
and U5448 (N_5448,N_4940,N_4941);
xnor U5449 (N_5449,N_4863,N_4544);
xnor U5450 (N_5450,N_4762,N_4639);
nor U5451 (N_5451,N_4897,N_4840);
and U5452 (N_5452,N_4571,N_4802);
nand U5453 (N_5453,N_4955,N_4534);
nand U5454 (N_5454,N_4729,N_4979);
or U5455 (N_5455,N_4962,N_4815);
or U5456 (N_5456,N_4858,N_4885);
nor U5457 (N_5457,N_4572,N_4916);
xor U5458 (N_5458,N_4927,N_4790);
and U5459 (N_5459,N_4677,N_4788);
xnor U5460 (N_5460,N_4829,N_4896);
nor U5461 (N_5461,N_4978,N_4546);
or U5462 (N_5462,N_4562,N_4820);
nand U5463 (N_5463,N_4880,N_4708);
xor U5464 (N_5464,N_4797,N_4884);
xor U5465 (N_5465,N_4663,N_4758);
and U5466 (N_5466,N_4564,N_4566);
nand U5467 (N_5467,N_4717,N_4623);
and U5468 (N_5468,N_4795,N_4684);
nand U5469 (N_5469,N_4550,N_4874);
or U5470 (N_5470,N_4612,N_4535);
and U5471 (N_5471,N_4760,N_4728);
or U5472 (N_5472,N_4946,N_4815);
or U5473 (N_5473,N_4704,N_4921);
nor U5474 (N_5474,N_4552,N_4775);
nand U5475 (N_5475,N_4900,N_4872);
or U5476 (N_5476,N_4581,N_4629);
nand U5477 (N_5477,N_4787,N_4686);
nor U5478 (N_5478,N_4608,N_4694);
and U5479 (N_5479,N_4591,N_4562);
or U5480 (N_5480,N_4727,N_4987);
or U5481 (N_5481,N_4596,N_4634);
xnor U5482 (N_5482,N_4610,N_4749);
or U5483 (N_5483,N_4913,N_4621);
nand U5484 (N_5484,N_4936,N_4588);
and U5485 (N_5485,N_4919,N_4606);
nor U5486 (N_5486,N_4960,N_4782);
xnor U5487 (N_5487,N_4868,N_4675);
and U5488 (N_5488,N_4958,N_4975);
or U5489 (N_5489,N_4658,N_4569);
xnor U5490 (N_5490,N_4702,N_4662);
nand U5491 (N_5491,N_4747,N_4835);
and U5492 (N_5492,N_4833,N_4873);
nand U5493 (N_5493,N_4605,N_4769);
nand U5494 (N_5494,N_4549,N_4783);
nand U5495 (N_5495,N_4761,N_4963);
nor U5496 (N_5496,N_4571,N_4681);
xor U5497 (N_5497,N_4508,N_4838);
nor U5498 (N_5498,N_4507,N_4643);
and U5499 (N_5499,N_4563,N_4809);
xnor U5500 (N_5500,N_5315,N_5262);
or U5501 (N_5501,N_5385,N_5448);
xnor U5502 (N_5502,N_5074,N_5342);
xnor U5503 (N_5503,N_5126,N_5192);
nor U5504 (N_5504,N_5169,N_5333);
xnor U5505 (N_5505,N_5305,N_5316);
and U5506 (N_5506,N_5129,N_5021);
and U5507 (N_5507,N_5038,N_5302);
nor U5508 (N_5508,N_5450,N_5304);
nor U5509 (N_5509,N_5405,N_5391);
or U5510 (N_5510,N_5407,N_5243);
xor U5511 (N_5511,N_5242,N_5040);
and U5512 (N_5512,N_5202,N_5390);
xnor U5513 (N_5513,N_5494,N_5370);
nand U5514 (N_5514,N_5053,N_5201);
xor U5515 (N_5515,N_5125,N_5272);
nor U5516 (N_5516,N_5257,N_5331);
xnor U5517 (N_5517,N_5488,N_5255);
or U5518 (N_5518,N_5499,N_5468);
and U5519 (N_5519,N_5303,N_5051);
nor U5520 (N_5520,N_5057,N_5470);
xor U5521 (N_5521,N_5235,N_5211);
nand U5522 (N_5522,N_5052,N_5377);
xnor U5523 (N_5523,N_5019,N_5193);
and U5524 (N_5524,N_5206,N_5352);
nand U5525 (N_5525,N_5250,N_5491);
nor U5526 (N_5526,N_5068,N_5217);
xnor U5527 (N_5527,N_5080,N_5170);
xnor U5528 (N_5528,N_5419,N_5449);
and U5529 (N_5529,N_5395,N_5138);
xnor U5530 (N_5530,N_5137,N_5279);
or U5531 (N_5531,N_5416,N_5381);
xor U5532 (N_5532,N_5064,N_5456);
xor U5533 (N_5533,N_5236,N_5451);
nor U5534 (N_5534,N_5152,N_5199);
nand U5535 (N_5535,N_5018,N_5042);
nand U5536 (N_5536,N_5301,N_5384);
nand U5537 (N_5537,N_5127,N_5288);
nor U5538 (N_5538,N_5299,N_5066);
xnor U5539 (N_5539,N_5411,N_5072);
and U5540 (N_5540,N_5266,N_5160);
or U5541 (N_5541,N_5404,N_5022);
xnor U5542 (N_5542,N_5088,N_5106);
or U5543 (N_5543,N_5130,N_5097);
nor U5544 (N_5544,N_5372,N_5163);
nand U5545 (N_5545,N_5007,N_5189);
or U5546 (N_5546,N_5026,N_5062);
nor U5547 (N_5547,N_5147,N_5002);
or U5548 (N_5548,N_5270,N_5135);
or U5549 (N_5549,N_5228,N_5350);
and U5550 (N_5550,N_5086,N_5082);
nor U5551 (N_5551,N_5161,N_5267);
and U5552 (N_5552,N_5368,N_5308);
nor U5553 (N_5553,N_5162,N_5183);
and U5554 (N_5554,N_5108,N_5076);
xnor U5555 (N_5555,N_5406,N_5083);
or U5556 (N_5556,N_5179,N_5004);
or U5557 (N_5557,N_5265,N_5196);
xor U5558 (N_5558,N_5188,N_5409);
xor U5559 (N_5559,N_5421,N_5037);
nor U5560 (N_5560,N_5222,N_5226);
nand U5561 (N_5561,N_5166,N_5480);
and U5562 (N_5562,N_5209,N_5017);
or U5563 (N_5563,N_5340,N_5223);
xnor U5564 (N_5564,N_5043,N_5477);
nand U5565 (N_5565,N_5447,N_5387);
nand U5566 (N_5566,N_5173,N_5020);
xor U5567 (N_5567,N_5109,N_5273);
nor U5568 (N_5568,N_5133,N_5280);
nor U5569 (N_5569,N_5092,N_5212);
xnor U5570 (N_5570,N_5149,N_5458);
xor U5571 (N_5571,N_5048,N_5438);
xnor U5572 (N_5572,N_5141,N_5357);
nand U5573 (N_5573,N_5124,N_5087);
and U5574 (N_5574,N_5346,N_5113);
and U5575 (N_5575,N_5142,N_5112);
xor U5576 (N_5576,N_5306,N_5165);
nor U5577 (N_5577,N_5444,N_5177);
nor U5578 (N_5578,N_5362,N_5376);
nand U5579 (N_5579,N_5420,N_5056);
and U5580 (N_5580,N_5261,N_5495);
and U5581 (N_5581,N_5032,N_5093);
xor U5582 (N_5582,N_5297,N_5281);
and U5583 (N_5583,N_5207,N_5187);
or U5584 (N_5584,N_5184,N_5401);
xnor U5585 (N_5585,N_5122,N_5107);
nor U5586 (N_5586,N_5388,N_5023);
or U5587 (N_5587,N_5389,N_5361);
and U5588 (N_5588,N_5329,N_5492);
and U5589 (N_5589,N_5213,N_5114);
nand U5590 (N_5590,N_5498,N_5383);
nor U5591 (N_5591,N_5335,N_5039);
or U5592 (N_5592,N_5237,N_5356);
or U5593 (N_5593,N_5230,N_5324);
and U5594 (N_5594,N_5460,N_5013);
and U5595 (N_5595,N_5185,N_5099);
nand U5596 (N_5596,N_5290,N_5485);
and U5597 (N_5597,N_5318,N_5061);
nor U5598 (N_5598,N_5474,N_5285);
nor U5599 (N_5599,N_5168,N_5360);
nand U5600 (N_5600,N_5031,N_5435);
nand U5601 (N_5601,N_5232,N_5428);
nand U5602 (N_5602,N_5364,N_5067);
and U5603 (N_5603,N_5172,N_5059);
nor U5604 (N_5604,N_5075,N_5328);
and U5605 (N_5605,N_5143,N_5454);
or U5606 (N_5606,N_5200,N_5497);
nor U5607 (N_5607,N_5144,N_5311);
and U5608 (N_5608,N_5476,N_5153);
or U5609 (N_5609,N_5229,N_5493);
or U5610 (N_5610,N_5176,N_5220);
nand U5611 (N_5611,N_5227,N_5483);
and U5612 (N_5612,N_5487,N_5289);
nand U5613 (N_5613,N_5060,N_5215);
xnor U5614 (N_5614,N_5365,N_5041);
nand U5615 (N_5615,N_5481,N_5089);
xnor U5616 (N_5616,N_5320,N_5269);
or U5617 (N_5617,N_5446,N_5218);
xnor U5618 (N_5618,N_5219,N_5374);
and U5619 (N_5619,N_5128,N_5055);
xnor U5620 (N_5620,N_5245,N_5392);
and U5621 (N_5621,N_5412,N_5256);
or U5622 (N_5622,N_5400,N_5422);
nor U5623 (N_5623,N_5371,N_5459);
xor U5624 (N_5624,N_5490,N_5065);
xnor U5625 (N_5625,N_5140,N_5102);
nor U5626 (N_5626,N_5465,N_5084);
nand U5627 (N_5627,N_5224,N_5115);
nand U5628 (N_5628,N_5131,N_5096);
nand U5629 (N_5629,N_5208,N_5095);
and U5630 (N_5630,N_5047,N_5001);
xnor U5631 (N_5631,N_5418,N_5035);
nor U5632 (N_5632,N_5314,N_5312);
nand U5633 (N_5633,N_5175,N_5054);
xnor U5634 (N_5634,N_5063,N_5073);
or U5635 (N_5635,N_5393,N_5445);
or U5636 (N_5636,N_5378,N_5249);
or U5637 (N_5637,N_5210,N_5496);
nand U5638 (N_5638,N_5367,N_5146);
nand U5639 (N_5639,N_5380,N_5337);
nor U5640 (N_5640,N_5134,N_5339);
nor U5641 (N_5641,N_5295,N_5292);
nand U5642 (N_5642,N_5413,N_5327);
nor U5643 (N_5643,N_5247,N_5101);
nor U5644 (N_5644,N_5085,N_5033);
nand U5645 (N_5645,N_5284,N_5355);
or U5646 (N_5646,N_5070,N_5348);
xnor U5647 (N_5647,N_5472,N_5330);
or U5648 (N_5648,N_5427,N_5046);
nor U5649 (N_5649,N_5464,N_5466);
xor U5650 (N_5650,N_5439,N_5091);
xor U5651 (N_5651,N_5251,N_5174);
nand U5652 (N_5652,N_5011,N_5349);
or U5653 (N_5653,N_5186,N_5473);
nor U5654 (N_5654,N_5443,N_5319);
or U5655 (N_5655,N_5424,N_5015);
and U5656 (N_5656,N_5440,N_5467);
and U5657 (N_5657,N_5027,N_5198);
or U5658 (N_5658,N_5426,N_5069);
nand U5659 (N_5659,N_5171,N_5478);
xor U5660 (N_5660,N_5382,N_5225);
and U5661 (N_5661,N_5034,N_5325);
nand U5662 (N_5662,N_5276,N_5167);
or U5663 (N_5663,N_5414,N_5151);
and U5664 (N_5664,N_5341,N_5111);
or U5665 (N_5665,N_5205,N_5351);
nor U5666 (N_5666,N_5323,N_5240);
or U5667 (N_5667,N_5486,N_5036);
nor U5668 (N_5668,N_5334,N_5058);
nand U5669 (N_5669,N_5252,N_5386);
or U5670 (N_5670,N_5136,N_5110);
or U5671 (N_5671,N_5397,N_5214);
xnor U5672 (N_5672,N_5132,N_5009);
or U5673 (N_5673,N_5090,N_5050);
or U5674 (N_5674,N_5359,N_5309);
and U5675 (N_5675,N_5078,N_5434);
and U5676 (N_5676,N_5442,N_5436);
nor U5677 (N_5677,N_5332,N_5430);
nand U5678 (N_5678,N_5118,N_5121);
or U5679 (N_5679,N_5307,N_5455);
or U5680 (N_5680,N_5344,N_5441);
xnor U5681 (N_5681,N_5238,N_5461);
xor U5682 (N_5682,N_5028,N_5234);
and U5683 (N_5683,N_5000,N_5159);
nand U5684 (N_5684,N_5016,N_5181);
xnor U5685 (N_5685,N_5024,N_5408);
nor U5686 (N_5686,N_5484,N_5313);
and U5687 (N_5687,N_5194,N_5429);
nand U5688 (N_5688,N_5336,N_5012);
xnor U5689 (N_5689,N_5182,N_5204);
nand U5690 (N_5690,N_5403,N_5150);
nand U5691 (N_5691,N_5119,N_5283);
nor U5692 (N_5692,N_5298,N_5231);
nand U5693 (N_5693,N_5010,N_5098);
xnor U5694 (N_5694,N_5216,N_5402);
nand U5695 (N_5695,N_5398,N_5433);
xor U5696 (N_5696,N_5094,N_5326);
xnor U5697 (N_5697,N_5275,N_5338);
nor U5698 (N_5698,N_5154,N_5100);
nor U5699 (N_5699,N_5258,N_5233);
nand U5700 (N_5700,N_5437,N_5025);
xnor U5701 (N_5701,N_5452,N_5294);
nand U5702 (N_5702,N_5241,N_5103);
nand U5703 (N_5703,N_5157,N_5071);
or U5704 (N_5704,N_5286,N_5139);
or U5705 (N_5705,N_5203,N_5432);
nand U5706 (N_5706,N_5369,N_5347);
and U5707 (N_5707,N_5417,N_5014);
and U5708 (N_5708,N_5379,N_5423);
nor U5709 (N_5709,N_5277,N_5471);
and U5710 (N_5710,N_5008,N_5264);
and U5711 (N_5711,N_5415,N_5463);
nand U5712 (N_5712,N_5006,N_5268);
nor U5713 (N_5713,N_5296,N_5253);
or U5714 (N_5714,N_5221,N_5489);
or U5715 (N_5715,N_5399,N_5271);
or U5716 (N_5716,N_5353,N_5195);
or U5717 (N_5717,N_5254,N_5322);
xor U5718 (N_5718,N_5366,N_5343);
nor U5719 (N_5719,N_5148,N_5164);
nand U5720 (N_5720,N_5310,N_5293);
and U5721 (N_5721,N_5354,N_5248);
nand U5722 (N_5722,N_5239,N_5300);
and U5723 (N_5723,N_5081,N_5317);
xnor U5724 (N_5724,N_5105,N_5278);
nand U5725 (N_5725,N_5117,N_5425);
nor U5726 (N_5726,N_5246,N_5263);
xor U5727 (N_5727,N_5191,N_5363);
and U5728 (N_5728,N_5190,N_5291);
and U5729 (N_5729,N_5197,N_5005);
nor U5730 (N_5730,N_5244,N_5457);
or U5731 (N_5731,N_5180,N_5431);
xor U5732 (N_5732,N_5321,N_5373);
and U5733 (N_5733,N_5158,N_5475);
nand U5734 (N_5734,N_5482,N_5120);
nand U5735 (N_5735,N_5282,N_5259);
or U5736 (N_5736,N_5123,N_5178);
xnor U5737 (N_5737,N_5155,N_5116);
or U5738 (N_5738,N_5396,N_5029);
or U5739 (N_5739,N_5462,N_5049);
nand U5740 (N_5740,N_5453,N_5003);
xnor U5741 (N_5741,N_5287,N_5044);
and U5742 (N_5742,N_5079,N_5274);
and U5743 (N_5743,N_5077,N_5469);
and U5744 (N_5744,N_5358,N_5045);
and U5745 (N_5745,N_5479,N_5345);
and U5746 (N_5746,N_5145,N_5394);
nor U5747 (N_5747,N_5410,N_5030);
or U5748 (N_5748,N_5104,N_5375);
nand U5749 (N_5749,N_5260,N_5156);
nand U5750 (N_5750,N_5166,N_5022);
xor U5751 (N_5751,N_5417,N_5095);
nand U5752 (N_5752,N_5489,N_5085);
and U5753 (N_5753,N_5094,N_5000);
or U5754 (N_5754,N_5294,N_5497);
xnor U5755 (N_5755,N_5153,N_5450);
nor U5756 (N_5756,N_5298,N_5143);
and U5757 (N_5757,N_5281,N_5395);
xnor U5758 (N_5758,N_5375,N_5075);
and U5759 (N_5759,N_5077,N_5002);
and U5760 (N_5760,N_5225,N_5338);
nor U5761 (N_5761,N_5196,N_5335);
nand U5762 (N_5762,N_5176,N_5181);
xnor U5763 (N_5763,N_5059,N_5425);
and U5764 (N_5764,N_5305,N_5319);
or U5765 (N_5765,N_5455,N_5333);
xor U5766 (N_5766,N_5361,N_5111);
nand U5767 (N_5767,N_5059,N_5019);
and U5768 (N_5768,N_5376,N_5025);
and U5769 (N_5769,N_5066,N_5354);
nand U5770 (N_5770,N_5344,N_5249);
and U5771 (N_5771,N_5207,N_5325);
xor U5772 (N_5772,N_5174,N_5290);
nand U5773 (N_5773,N_5016,N_5072);
nand U5774 (N_5774,N_5429,N_5369);
and U5775 (N_5775,N_5169,N_5484);
nor U5776 (N_5776,N_5307,N_5008);
nor U5777 (N_5777,N_5029,N_5463);
and U5778 (N_5778,N_5385,N_5205);
nor U5779 (N_5779,N_5459,N_5168);
and U5780 (N_5780,N_5476,N_5031);
or U5781 (N_5781,N_5325,N_5200);
and U5782 (N_5782,N_5059,N_5091);
xor U5783 (N_5783,N_5154,N_5044);
nor U5784 (N_5784,N_5417,N_5462);
or U5785 (N_5785,N_5379,N_5099);
nor U5786 (N_5786,N_5074,N_5246);
xor U5787 (N_5787,N_5177,N_5000);
xnor U5788 (N_5788,N_5046,N_5401);
nand U5789 (N_5789,N_5000,N_5266);
xor U5790 (N_5790,N_5380,N_5270);
and U5791 (N_5791,N_5406,N_5317);
xnor U5792 (N_5792,N_5266,N_5142);
xor U5793 (N_5793,N_5411,N_5403);
and U5794 (N_5794,N_5467,N_5366);
or U5795 (N_5795,N_5213,N_5322);
or U5796 (N_5796,N_5462,N_5489);
or U5797 (N_5797,N_5198,N_5434);
nand U5798 (N_5798,N_5252,N_5101);
nand U5799 (N_5799,N_5241,N_5250);
or U5800 (N_5800,N_5006,N_5137);
nor U5801 (N_5801,N_5361,N_5396);
and U5802 (N_5802,N_5291,N_5301);
or U5803 (N_5803,N_5245,N_5402);
nand U5804 (N_5804,N_5117,N_5157);
nand U5805 (N_5805,N_5099,N_5221);
xnor U5806 (N_5806,N_5082,N_5112);
and U5807 (N_5807,N_5433,N_5198);
nor U5808 (N_5808,N_5436,N_5086);
and U5809 (N_5809,N_5273,N_5411);
nand U5810 (N_5810,N_5321,N_5428);
and U5811 (N_5811,N_5354,N_5276);
nor U5812 (N_5812,N_5033,N_5428);
nand U5813 (N_5813,N_5058,N_5426);
or U5814 (N_5814,N_5293,N_5215);
nor U5815 (N_5815,N_5090,N_5126);
nor U5816 (N_5816,N_5098,N_5130);
or U5817 (N_5817,N_5316,N_5177);
nand U5818 (N_5818,N_5034,N_5320);
nor U5819 (N_5819,N_5452,N_5407);
and U5820 (N_5820,N_5055,N_5292);
xor U5821 (N_5821,N_5153,N_5130);
xor U5822 (N_5822,N_5327,N_5178);
xnor U5823 (N_5823,N_5284,N_5307);
or U5824 (N_5824,N_5038,N_5409);
nor U5825 (N_5825,N_5253,N_5341);
xor U5826 (N_5826,N_5193,N_5164);
and U5827 (N_5827,N_5229,N_5188);
nor U5828 (N_5828,N_5175,N_5082);
and U5829 (N_5829,N_5035,N_5166);
nand U5830 (N_5830,N_5448,N_5331);
nor U5831 (N_5831,N_5430,N_5288);
or U5832 (N_5832,N_5333,N_5042);
and U5833 (N_5833,N_5468,N_5196);
nor U5834 (N_5834,N_5103,N_5099);
xor U5835 (N_5835,N_5172,N_5434);
xnor U5836 (N_5836,N_5226,N_5028);
and U5837 (N_5837,N_5014,N_5486);
or U5838 (N_5838,N_5408,N_5493);
nor U5839 (N_5839,N_5136,N_5471);
and U5840 (N_5840,N_5069,N_5206);
nor U5841 (N_5841,N_5126,N_5488);
or U5842 (N_5842,N_5394,N_5442);
nand U5843 (N_5843,N_5416,N_5147);
and U5844 (N_5844,N_5270,N_5245);
and U5845 (N_5845,N_5213,N_5411);
or U5846 (N_5846,N_5006,N_5122);
or U5847 (N_5847,N_5402,N_5438);
xor U5848 (N_5848,N_5237,N_5233);
xor U5849 (N_5849,N_5245,N_5397);
nand U5850 (N_5850,N_5004,N_5390);
and U5851 (N_5851,N_5366,N_5145);
and U5852 (N_5852,N_5455,N_5141);
or U5853 (N_5853,N_5196,N_5493);
nand U5854 (N_5854,N_5318,N_5275);
and U5855 (N_5855,N_5329,N_5430);
nand U5856 (N_5856,N_5403,N_5342);
nand U5857 (N_5857,N_5082,N_5018);
nor U5858 (N_5858,N_5064,N_5489);
or U5859 (N_5859,N_5247,N_5237);
and U5860 (N_5860,N_5102,N_5391);
and U5861 (N_5861,N_5277,N_5246);
nor U5862 (N_5862,N_5193,N_5131);
and U5863 (N_5863,N_5232,N_5016);
or U5864 (N_5864,N_5408,N_5046);
and U5865 (N_5865,N_5313,N_5104);
or U5866 (N_5866,N_5484,N_5181);
or U5867 (N_5867,N_5032,N_5484);
and U5868 (N_5868,N_5262,N_5384);
nand U5869 (N_5869,N_5255,N_5161);
and U5870 (N_5870,N_5259,N_5281);
or U5871 (N_5871,N_5021,N_5316);
and U5872 (N_5872,N_5149,N_5466);
xnor U5873 (N_5873,N_5250,N_5041);
or U5874 (N_5874,N_5252,N_5034);
or U5875 (N_5875,N_5364,N_5041);
nand U5876 (N_5876,N_5143,N_5030);
or U5877 (N_5877,N_5410,N_5345);
nor U5878 (N_5878,N_5197,N_5404);
and U5879 (N_5879,N_5309,N_5026);
or U5880 (N_5880,N_5470,N_5417);
xor U5881 (N_5881,N_5007,N_5177);
and U5882 (N_5882,N_5481,N_5174);
nand U5883 (N_5883,N_5342,N_5123);
nor U5884 (N_5884,N_5144,N_5356);
and U5885 (N_5885,N_5357,N_5450);
nand U5886 (N_5886,N_5465,N_5332);
nor U5887 (N_5887,N_5370,N_5435);
xnor U5888 (N_5888,N_5444,N_5338);
and U5889 (N_5889,N_5219,N_5067);
nand U5890 (N_5890,N_5425,N_5338);
and U5891 (N_5891,N_5023,N_5480);
or U5892 (N_5892,N_5103,N_5289);
and U5893 (N_5893,N_5474,N_5085);
and U5894 (N_5894,N_5135,N_5238);
and U5895 (N_5895,N_5295,N_5003);
or U5896 (N_5896,N_5015,N_5476);
or U5897 (N_5897,N_5173,N_5145);
nor U5898 (N_5898,N_5006,N_5319);
nor U5899 (N_5899,N_5471,N_5164);
nor U5900 (N_5900,N_5075,N_5103);
and U5901 (N_5901,N_5371,N_5014);
or U5902 (N_5902,N_5209,N_5267);
xor U5903 (N_5903,N_5203,N_5354);
and U5904 (N_5904,N_5170,N_5086);
nand U5905 (N_5905,N_5083,N_5040);
nor U5906 (N_5906,N_5092,N_5154);
nand U5907 (N_5907,N_5043,N_5401);
xnor U5908 (N_5908,N_5321,N_5265);
nand U5909 (N_5909,N_5296,N_5184);
xor U5910 (N_5910,N_5066,N_5128);
nor U5911 (N_5911,N_5483,N_5028);
or U5912 (N_5912,N_5120,N_5362);
nand U5913 (N_5913,N_5375,N_5226);
and U5914 (N_5914,N_5096,N_5016);
nor U5915 (N_5915,N_5332,N_5195);
nand U5916 (N_5916,N_5465,N_5486);
nand U5917 (N_5917,N_5343,N_5348);
and U5918 (N_5918,N_5259,N_5457);
xnor U5919 (N_5919,N_5342,N_5092);
and U5920 (N_5920,N_5037,N_5324);
nand U5921 (N_5921,N_5381,N_5495);
xnor U5922 (N_5922,N_5205,N_5159);
or U5923 (N_5923,N_5423,N_5351);
xnor U5924 (N_5924,N_5439,N_5293);
or U5925 (N_5925,N_5368,N_5457);
and U5926 (N_5926,N_5038,N_5029);
nand U5927 (N_5927,N_5351,N_5378);
or U5928 (N_5928,N_5051,N_5306);
nand U5929 (N_5929,N_5028,N_5274);
and U5930 (N_5930,N_5008,N_5257);
nor U5931 (N_5931,N_5270,N_5228);
and U5932 (N_5932,N_5228,N_5486);
or U5933 (N_5933,N_5087,N_5389);
and U5934 (N_5934,N_5177,N_5222);
and U5935 (N_5935,N_5427,N_5455);
nor U5936 (N_5936,N_5368,N_5085);
and U5937 (N_5937,N_5379,N_5285);
or U5938 (N_5938,N_5007,N_5253);
nand U5939 (N_5939,N_5402,N_5415);
xor U5940 (N_5940,N_5177,N_5073);
nand U5941 (N_5941,N_5369,N_5492);
nor U5942 (N_5942,N_5441,N_5127);
nand U5943 (N_5943,N_5160,N_5261);
nor U5944 (N_5944,N_5438,N_5086);
xor U5945 (N_5945,N_5426,N_5360);
nand U5946 (N_5946,N_5040,N_5179);
nor U5947 (N_5947,N_5460,N_5110);
or U5948 (N_5948,N_5224,N_5090);
nand U5949 (N_5949,N_5040,N_5255);
and U5950 (N_5950,N_5480,N_5171);
nand U5951 (N_5951,N_5158,N_5191);
xnor U5952 (N_5952,N_5458,N_5202);
nand U5953 (N_5953,N_5237,N_5248);
nor U5954 (N_5954,N_5471,N_5309);
and U5955 (N_5955,N_5085,N_5011);
xnor U5956 (N_5956,N_5309,N_5241);
and U5957 (N_5957,N_5391,N_5303);
xnor U5958 (N_5958,N_5363,N_5189);
and U5959 (N_5959,N_5030,N_5317);
or U5960 (N_5960,N_5354,N_5040);
nand U5961 (N_5961,N_5343,N_5248);
nand U5962 (N_5962,N_5452,N_5320);
nor U5963 (N_5963,N_5234,N_5342);
xnor U5964 (N_5964,N_5355,N_5220);
and U5965 (N_5965,N_5158,N_5314);
nor U5966 (N_5966,N_5137,N_5286);
and U5967 (N_5967,N_5466,N_5230);
or U5968 (N_5968,N_5124,N_5455);
nor U5969 (N_5969,N_5243,N_5021);
xnor U5970 (N_5970,N_5141,N_5010);
nand U5971 (N_5971,N_5227,N_5219);
or U5972 (N_5972,N_5079,N_5263);
nand U5973 (N_5973,N_5031,N_5043);
xnor U5974 (N_5974,N_5048,N_5331);
or U5975 (N_5975,N_5010,N_5382);
nand U5976 (N_5976,N_5218,N_5117);
or U5977 (N_5977,N_5000,N_5270);
and U5978 (N_5978,N_5081,N_5106);
xor U5979 (N_5979,N_5250,N_5474);
nand U5980 (N_5980,N_5003,N_5301);
xor U5981 (N_5981,N_5012,N_5302);
nand U5982 (N_5982,N_5179,N_5130);
or U5983 (N_5983,N_5107,N_5197);
and U5984 (N_5984,N_5326,N_5354);
xnor U5985 (N_5985,N_5184,N_5199);
nor U5986 (N_5986,N_5010,N_5437);
or U5987 (N_5987,N_5282,N_5300);
nand U5988 (N_5988,N_5461,N_5165);
or U5989 (N_5989,N_5031,N_5236);
nor U5990 (N_5990,N_5372,N_5384);
xnor U5991 (N_5991,N_5181,N_5023);
xor U5992 (N_5992,N_5165,N_5422);
nand U5993 (N_5993,N_5341,N_5029);
or U5994 (N_5994,N_5348,N_5025);
and U5995 (N_5995,N_5054,N_5180);
nand U5996 (N_5996,N_5218,N_5158);
and U5997 (N_5997,N_5491,N_5011);
and U5998 (N_5998,N_5053,N_5228);
nand U5999 (N_5999,N_5172,N_5394);
nor U6000 (N_6000,N_5790,N_5858);
and U6001 (N_6001,N_5728,N_5609);
nand U6002 (N_6002,N_5710,N_5791);
and U6003 (N_6003,N_5962,N_5949);
or U6004 (N_6004,N_5652,N_5562);
nor U6005 (N_6005,N_5509,N_5620);
nand U6006 (N_6006,N_5785,N_5892);
xor U6007 (N_6007,N_5912,N_5686);
nand U6008 (N_6008,N_5715,N_5586);
or U6009 (N_6009,N_5544,N_5991);
and U6010 (N_6010,N_5999,N_5532);
xnor U6011 (N_6011,N_5902,N_5923);
nor U6012 (N_6012,N_5665,N_5657);
nand U6013 (N_6013,N_5663,N_5582);
nor U6014 (N_6014,N_5674,N_5914);
xnor U6015 (N_6015,N_5700,N_5784);
nand U6016 (N_6016,N_5805,N_5617);
and U6017 (N_6017,N_5897,N_5824);
and U6018 (N_6018,N_5636,N_5577);
and U6019 (N_6019,N_5653,N_5862);
and U6020 (N_6020,N_5878,N_5597);
and U6021 (N_6021,N_5554,N_5740);
nor U6022 (N_6022,N_5865,N_5987);
xor U6023 (N_6023,N_5573,N_5781);
nand U6024 (N_6024,N_5520,N_5706);
xnor U6025 (N_6025,N_5720,N_5990);
xnor U6026 (N_6026,N_5519,N_5551);
nand U6027 (N_6027,N_5697,N_5887);
nand U6028 (N_6028,N_5623,N_5545);
or U6029 (N_6029,N_5813,N_5789);
and U6030 (N_6030,N_5753,N_5548);
nor U6031 (N_6031,N_5901,N_5927);
or U6032 (N_6032,N_5560,N_5794);
xnor U6033 (N_6033,N_5922,N_5803);
and U6034 (N_6034,N_5846,N_5632);
and U6035 (N_6035,N_5527,N_5518);
nand U6036 (N_6036,N_5667,N_5910);
and U6037 (N_6037,N_5589,N_5960);
and U6038 (N_6038,N_5648,N_5777);
xnor U6039 (N_6039,N_5644,N_5564);
or U6040 (N_6040,N_5875,N_5553);
or U6041 (N_6041,N_5646,N_5619);
xor U6042 (N_6042,N_5977,N_5868);
xor U6043 (N_6043,N_5935,N_5951);
and U6044 (N_6044,N_5861,N_5825);
and U6045 (N_6045,N_5963,N_5613);
nand U6046 (N_6046,N_5832,N_5621);
nand U6047 (N_6047,N_5570,N_5507);
and U6048 (N_6048,N_5880,N_5886);
and U6049 (N_6049,N_5952,N_5978);
and U6050 (N_6050,N_5762,N_5581);
xnor U6051 (N_6051,N_5655,N_5747);
nor U6052 (N_6052,N_5983,N_5967);
nand U6053 (N_6053,N_5847,N_5894);
xnor U6054 (N_6054,N_5684,N_5917);
xor U6055 (N_6055,N_5647,N_5682);
and U6056 (N_6056,N_5763,N_5840);
or U6057 (N_6057,N_5871,N_5662);
nand U6058 (N_6058,N_5543,N_5919);
xor U6059 (N_6059,N_5766,N_5516);
or U6060 (N_6060,N_5680,N_5826);
or U6061 (N_6061,N_5556,N_5976);
nor U6062 (N_6062,N_5523,N_5735);
nand U6063 (N_6063,N_5515,N_5678);
nor U6064 (N_6064,N_5957,N_5968);
nor U6065 (N_6065,N_5721,N_5725);
and U6066 (N_6066,N_5585,N_5669);
xor U6067 (N_6067,N_5637,N_5691);
nor U6068 (N_6068,N_5618,N_5932);
nand U6069 (N_6069,N_5925,N_5607);
or U6070 (N_6070,N_5852,N_5659);
nor U6071 (N_6071,N_5526,N_5679);
or U6072 (N_6072,N_5881,N_5676);
nor U6073 (N_6073,N_5822,N_5997);
nor U6074 (N_6074,N_5729,N_5671);
nor U6075 (N_6075,N_5816,N_5883);
xnor U6076 (N_6076,N_5734,N_5829);
or U6077 (N_6077,N_5797,N_5546);
and U6078 (N_6078,N_5780,N_5599);
nand U6079 (N_6079,N_5630,N_5774);
nand U6080 (N_6080,N_5749,N_5578);
xnor U6081 (N_6081,N_5773,N_5614);
nor U6082 (N_6082,N_5939,N_5755);
xor U6083 (N_6083,N_5696,N_5907);
nor U6084 (N_6084,N_5699,N_5895);
xnor U6085 (N_6085,N_5786,N_5973);
and U6086 (N_6086,N_5770,N_5835);
nand U6087 (N_6087,N_5661,N_5966);
and U6088 (N_6088,N_5579,N_5827);
and U6089 (N_6089,N_5672,N_5645);
xor U6090 (N_6090,N_5675,N_5702);
xor U6091 (N_6091,N_5819,N_5559);
nand U6092 (N_6092,N_5857,N_5802);
and U6093 (N_6093,N_5779,N_5870);
or U6094 (N_6094,N_5792,N_5535);
xor U6095 (N_6095,N_5558,N_5701);
or U6096 (N_6096,N_5771,N_5956);
nand U6097 (N_6097,N_5521,N_5529);
nor U6098 (N_6098,N_5838,N_5542);
and U6099 (N_6099,N_5508,N_5530);
and U6100 (N_6100,N_5948,N_5909);
or U6101 (N_6101,N_5555,N_5600);
nor U6102 (N_6102,N_5622,N_5800);
nand U6103 (N_6103,N_5574,N_5944);
and U6104 (N_6104,N_5920,N_5764);
nor U6105 (N_6105,N_5685,N_5591);
nor U6106 (N_6106,N_5566,N_5795);
and U6107 (N_6107,N_5673,N_5627);
and U6108 (N_6108,N_5760,N_5732);
xor U6109 (N_6109,N_5538,N_5929);
or U6110 (N_6110,N_5534,N_5612);
and U6111 (N_6111,N_5565,N_5756);
xnor U6112 (N_6112,N_5851,N_5751);
or U6113 (N_6113,N_5714,N_5666);
xnor U6114 (N_6114,N_5945,N_5890);
nand U6115 (N_6115,N_5950,N_5658);
xnor U6116 (N_6116,N_5668,N_5514);
nand U6117 (N_6117,N_5568,N_5693);
xor U6118 (N_6118,N_5758,N_5955);
or U6119 (N_6119,N_5730,N_5596);
xor U6120 (N_6120,N_5921,N_5717);
nor U6121 (N_6121,N_5625,N_5831);
or U6122 (N_6122,N_5629,N_5841);
xnor U6123 (N_6123,N_5814,N_5801);
and U6124 (N_6124,N_5818,N_5635);
xor U6125 (N_6125,N_5873,N_5593);
nor U6126 (N_6126,N_5884,N_5694);
or U6127 (N_6127,N_5782,N_5634);
or U6128 (N_6128,N_5876,N_5745);
and U6129 (N_6129,N_5640,N_5913);
xor U6130 (N_6130,N_5736,N_5830);
xnor U6131 (N_6131,N_5754,N_5930);
nor U6132 (N_6132,N_5744,N_5848);
and U6133 (N_6133,N_5820,N_5569);
nand U6134 (N_6134,N_5850,N_5934);
xor U6135 (N_6135,N_5712,N_5650);
nor U6136 (N_6136,N_5810,N_5624);
xnor U6137 (N_6137,N_5525,N_5995);
xnor U6138 (N_6138,N_5726,N_5752);
nor U6139 (N_6139,N_5550,N_5692);
xnor U6140 (N_6140,N_5988,N_5704);
nand U6141 (N_6141,N_5812,N_5855);
and U6142 (N_6142,N_5787,N_5727);
or U6143 (N_6143,N_5849,N_5877);
or U6144 (N_6144,N_5903,N_5961);
nand U6145 (N_6145,N_5687,N_5683);
or U6146 (N_6146,N_5711,N_5946);
xnor U6147 (N_6147,N_5759,N_5761);
xor U6148 (N_6148,N_5750,N_5874);
xor U6149 (N_6149,N_5842,N_5911);
xor U6150 (N_6150,N_5567,N_5972);
xor U6151 (N_6151,N_5866,N_5608);
xor U6152 (N_6152,N_5943,N_5867);
nand U6153 (N_6153,N_5998,N_5722);
or U6154 (N_6154,N_5746,N_5821);
nand U6155 (N_6155,N_5718,N_5601);
and U6156 (N_6156,N_5808,N_5924);
nand U6157 (N_6157,N_5985,N_5788);
or U6158 (N_6158,N_5709,N_5954);
or U6159 (N_6159,N_5575,N_5641);
or U6160 (N_6160,N_5626,N_5860);
and U6161 (N_6161,N_5522,N_5888);
and U6162 (N_6162,N_5859,N_5615);
nor U6163 (N_6163,N_5768,N_5992);
xor U6164 (N_6164,N_5941,N_5980);
nand U6165 (N_6165,N_5708,N_5643);
and U6166 (N_6166,N_5879,N_5572);
nor U6167 (N_6167,N_5833,N_5681);
nand U6168 (N_6168,N_5500,N_5900);
and U6169 (N_6169,N_5703,N_5864);
or U6170 (N_6170,N_5937,N_5970);
nand U6171 (N_6171,N_5723,N_5834);
nand U6172 (N_6172,N_5656,N_5811);
or U6173 (N_6173,N_5670,N_5605);
and U6174 (N_6174,N_5796,N_5505);
nor U6175 (N_6175,N_5926,N_5885);
xnor U6176 (N_6176,N_5539,N_5537);
or U6177 (N_6177,N_5610,N_5513);
nor U6178 (N_6178,N_5843,N_5936);
nand U6179 (N_6179,N_5767,N_5837);
nand U6180 (N_6180,N_5975,N_5738);
or U6181 (N_6181,N_5677,N_5631);
and U6182 (N_6182,N_5982,N_5517);
and U6183 (N_6183,N_5893,N_5651);
nand U6184 (N_6184,N_5844,N_5733);
xnor U6185 (N_6185,N_5896,N_5965);
nor U6186 (N_6186,N_5953,N_5815);
and U6187 (N_6187,N_5898,N_5611);
nor U6188 (N_6188,N_5695,N_5828);
and U6189 (N_6189,N_5511,N_5969);
nand U6190 (N_6190,N_5775,N_5856);
nand U6191 (N_6191,N_5510,N_5845);
and U6192 (N_6192,N_5642,N_5882);
nand U6193 (N_6193,N_5915,N_5595);
or U6194 (N_6194,N_5716,N_5616);
nand U6195 (N_6195,N_5904,N_5504);
xnor U6196 (N_6196,N_5928,N_5664);
nand U6197 (N_6197,N_5869,N_5590);
xor U6198 (N_6198,N_5793,N_5571);
xnor U6199 (N_6199,N_5724,N_5501);
nand U6200 (N_6200,N_5552,N_5958);
and U6201 (N_6201,N_5576,N_5549);
nand U6202 (N_6202,N_5713,N_5563);
and U6203 (N_6203,N_5541,N_5776);
nor U6204 (N_6204,N_5528,N_5839);
or U6205 (N_6205,N_5743,N_5817);
xor U6206 (N_6206,N_5964,N_5986);
or U6207 (N_6207,N_5778,N_5707);
and U6208 (N_6208,N_5587,N_5654);
and U6209 (N_6209,N_5592,N_5540);
nor U6210 (N_6210,N_5804,N_5561);
xnor U6211 (N_6211,N_5916,N_5971);
or U6212 (N_6212,N_5698,N_5604);
or U6213 (N_6213,N_5905,N_5979);
and U6214 (N_6214,N_5606,N_5628);
or U6215 (N_6215,N_5602,N_5889);
and U6216 (N_6216,N_5854,N_5947);
nor U6217 (N_6217,N_5993,N_5731);
nand U6218 (N_6218,N_5741,N_5739);
nand U6219 (N_6219,N_5639,N_5547);
and U6220 (N_6220,N_5772,N_5942);
nor U6221 (N_6221,N_5584,N_5769);
nand U6222 (N_6222,N_5959,N_5503);
and U6223 (N_6223,N_5918,N_5853);
nor U6224 (N_6224,N_5836,N_5583);
nor U6225 (N_6225,N_5580,N_5533);
nand U6226 (N_6226,N_5633,N_5807);
nor U6227 (N_6227,N_5649,N_5688);
nor U6228 (N_6228,N_5594,N_5719);
nor U6229 (N_6229,N_5524,N_5502);
nand U6230 (N_6230,N_5863,N_5536);
and U6231 (N_6231,N_5891,N_5981);
nor U6232 (N_6232,N_5742,N_5799);
nand U6233 (N_6233,N_5872,N_5933);
nor U6234 (N_6234,N_5931,N_5603);
nand U6235 (N_6235,N_5798,N_5908);
xnor U6236 (N_6236,N_5809,N_5989);
xor U6237 (N_6237,N_5938,N_5757);
nand U6238 (N_6238,N_5748,N_5690);
nor U6239 (N_6239,N_5906,N_5598);
nand U6240 (N_6240,N_5899,N_5660);
xnor U6241 (N_6241,N_5940,N_5984);
or U6242 (N_6242,N_5765,N_5737);
or U6243 (N_6243,N_5996,N_5638);
nor U6244 (N_6244,N_5689,N_5506);
or U6245 (N_6245,N_5806,N_5557);
nor U6246 (N_6246,N_5588,N_5705);
nor U6247 (N_6247,N_5512,N_5531);
nor U6248 (N_6248,N_5783,N_5823);
nor U6249 (N_6249,N_5994,N_5974);
and U6250 (N_6250,N_5862,N_5919);
xor U6251 (N_6251,N_5574,N_5663);
nor U6252 (N_6252,N_5655,N_5596);
xnor U6253 (N_6253,N_5892,N_5953);
or U6254 (N_6254,N_5641,N_5770);
nand U6255 (N_6255,N_5574,N_5963);
nor U6256 (N_6256,N_5659,N_5616);
nand U6257 (N_6257,N_5543,N_5508);
nor U6258 (N_6258,N_5915,N_5828);
and U6259 (N_6259,N_5682,N_5953);
xnor U6260 (N_6260,N_5837,N_5819);
xor U6261 (N_6261,N_5844,N_5913);
or U6262 (N_6262,N_5900,N_5846);
and U6263 (N_6263,N_5957,N_5863);
nand U6264 (N_6264,N_5858,N_5511);
nor U6265 (N_6265,N_5616,N_5895);
and U6266 (N_6266,N_5752,N_5912);
nand U6267 (N_6267,N_5513,N_5727);
nand U6268 (N_6268,N_5996,N_5970);
xnor U6269 (N_6269,N_5799,N_5950);
nand U6270 (N_6270,N_5897,N_5605);
nand U6271 (N_6271,N_5638,N_5510);
and U6272 (N_6272,N_5516,N_5509);
nand U6273 (N_6273,N_5752,N_5668);
and U6274 (N_6274,N_5643,N_5611);
nand U6275 (N_6275,N_5922,N_5852);
or U6276 (N_6276,N_5671,N_5870);
nand U6277 (N_6277,N_5647,N_5921);
nor U6278 (N_6278,N_5581,N_5913);
or U6279 (N_6279,N_5774,N_5745);
and U6280 (N_6280,N_5824,N_5919);
and U6281 (N_6281,N_5598,N_5553);
xnor U6282 (N_6282,N_5794,N_5606);
and U6283 (N_6283,N_5921,N_5898);
and U6284 (N_6284,N_5996,N_5550);
nand U6285 (N_6285,N_5972,N_5795);
nand U6286 (N_6286,N_5655,N_5616);
xnor U6287 (N_6287,N_5968,N_5643);
and U6288 (N_6288,N_5795,N_5892);
xor U6289 (N_6289,N_5573,N_5902);
nand U6290 (N_6290,N_5820,N_5695);
and U6291 (N_6291,N_5656,N_5878);
nand U6292 (N_6292,N_5656,N_5951);
or U6293 (N_6293,N_5842,N_5985);
or U6294 (N_6294,N_5999,N_5627);
or U6295 (N_6295,N_5765,N_5598);
and U6296 (N_6296,N_5633,N_5615);
nand U6297 (N_6297,N_5569,N_5502);
and U6298 (N_6298,N_5587,N_5708);
nor U6299 (N_6299,N_5741,N_5908);
and U6300 (N_6300,N_5778,N_5585);
nor U6301 (N_6301,N_5568,N_5949);
nor U6302 (N_6302,N_5770,N_5546);
or U6303 (N_6303,N_5655,N_5959);
and U6304 (N_6304,N_5997,N_5872);
and U6305 (N_6305,N_5553,N_5821);
xor U6306 (N_6306,N_5745,N_5637);
or U6307 (N_6307,N_5755,N_5572);
or U6308 (N_6308,N_5918,N_5531);
xnor U6309 (N_6309,N_5699,N_5525);
and U6310 (N_6310,N_5588,N_5736);
nor U6311 (N_6311,N_5997,N_5620);
nor U6312 (N_6312,N_5961,N_5877);
nand U6313 (N_6313,N_5558,N_5879);
nor U6314 (N_6314,N_5508,N_5741);
nand U6315 (N_6315,N_5838,N_5903);
and U6316 (N_6316,N_5858,N_5577);
or U6317 (N_6317,N_5617,N_5955);
and U6318 (N_6318,N_5969,N_5534);
nor U6319 (N_6319,N_5503,N_5819);
xor U6320 (N_6320,N_5820,N_5884);
and U6321 (N_6321,N_5760,N_5892);
nor U6322 (N_6322,N_5937,N_5950);
nor U6323 (N_6323,N_5759,N_5585);
nand U6324 (N_6324,N_5712,N_5731);
nor U6325 (N_6325,N_5935,N_5855);
or U6326 (N_6326,N_5529,N_5798);
and U6327 (N_6327,N_5653,N_5774);
and U6328 (N_6328,N_5629,N_5829);
and U6329 (N_6329,N_5785,N_5974);
nor U6330 (N_6330,N_5802,N_5640);
nor U6331 (N_6331,N_5820,N_5650);
or U6332 (N_6332,N_5759,N_5738);
and U6333 (N_6333,N_5930,N_5518);
nor U6334 (N_6334,N_5811,N_5884);
or U6335 (N_6335,N_5904,N_5901);
nand U6336 (N_6336,N_5987,N_5884);
nor U6337 (N_6337,N_5536,N_5735);
nor U6338 (N_6338,N_5628,N_5517);
and U6339 (N_6339,N_5699,N_5723);
or U6340 (N_6340,N_5718,N_5819);
and U6341 (N_6341,N_5597,N_5634);
nor U6342 (N_6342,N_5672,N_5886);
xor U6343 (N_6343,N_5806,N_5918);
xnor U6344 (N_6344,N_5696,N_5743);
xor U6345 (N_6345,N_5667,N_5974);
or U6346 (N_6346,N_5954,N_5618);
or U6347 (N_6347,N_5837,N_5860);
xor U6348 (N_6348,N_5685,N_5565);
nand U6349 (N_6349,N_5803,N_5733);
or U6350 (N_6350,N_5570,N_5534);
or U6351 (N_6351,N_5571,N_5875);
xor U6352 (N_6352,N_5735,N_5785);
xnor U6353 (N_6353,N_5957,N_5562);
xnor U6354 (N_6354,N_5763,N_5729);
nand U6355 (N_6355,N_5842,N_5510);
nor U6356 (N_6356,N_5798,N_5829);
and U6357 (N_6357,N_5873,N_5905);
or U6358 (N_6358,N_5877,N_5567);
or U6359 (N_6359,N_5744,N_5865);
nor U6360 (N_6360,N_5507,N_5805);
xor U6361 (N_6361,N_5799,N_5559);
nor U6362 (N_6362,N_5840,N_5618);
nand U6363 (N_6363,N_5567,N_5738);
xnor U6364 (N_6364,N_5530,N_5562);
or U6365 (N_6365,N_5672,N_5859);
xor U6366 (N_6366,N_5813,N_5726);
and U6367 (N_6367,N_5946,N_5955);
nand U6368 (N_6368,N_5618,N_5893);
or U6369 (N_6369,N_5952,N_5597);
xnor U6370 (N_6370,N_5975,N_5551);
nand U6371 (N_6371,N_5992,N_5721);
xor U6372 (N_6372,N_5899,N_5722);
xor U6373 (N_6373,N_5777,N_5978);
or U6374 (N_6374,N_5564,N_5654);
nor U6375 (N_6375,N_5614,N_5823);
nand U6376 (N_6376,N_5572,N_5916);
nor U6377 (N_6377,N_5834,N_5552);
and U6378 (N_6378,N_5505,N_5532);
and U6379 (N_6379,N_5821,N_5563);
and U6380 (N_6380,N_5844,N_5591);
nor U6381 (N_6381,N_5594,N_5530);
or U6382 (N_6382,N_5975,N_5511);
xnor U6383 (N_6383,N_5626,N_5683);
nor U6384 (N_6384,N_5639,N_5710);
nor U6385 (N_6385,N_5848,N_5767);
nor U6386 (N_6386,N_5577,N_5826);
or U6387 (N_6387,N_5568,N_5953);
nand U6388 (N_6388,N_5595,N_5827);
xor U6389 (N_6389,N_5728,N_5964);
nand U6390 (N_6390,N_5519,N_5581);
or U6391 (N_6391,N_5752,N_5939);
xnor U6392 (N_6392,N_5981,N_5628);
nor U6393 (N_6393,N_5721,N_5746);
nand U6394 (N_6394,N_5884,N_5617);
xnor U6395 (N_6395,N_5593,N_5825);
and U6396 (N_6396,N_5917,N_5925);
nand U6397 (N_6397,N_5934,N_5758);
nand U6398 (N_6398,N_5877,N_5664);
nor U6399 (N_6399,N_5959,N_5785);
xnor U6400 (N_6400,N_5620,N_5754);
nand U6401 (N_6401,N_5544,N_5831);
nor U6402 (N_6402,N_5614,N_5704);
xnor U6403 (N_6403,N_5620,N_5892);
nor U6404 (N_6404,N_5672,N_5899);
xnor U6405 (N_6405,N_5809,N_5570);
or U6406 (N_6406,N_5783,N_5549);
and U6407 (N_6407,N_5869,N_5611);
nand U6408 (N_6408,N_5517,N_5590);
xor U6409 (N_6409,N_5559,N_5960);
nor U6410 (N_6410,N_5615,N_5667);
or U6411 (N_6411,N_5943,N_5892);
nand U6412 (N_6412,N_5669,N_5977);
nor U6413 (N_6413,N_5900,N_5966);
and U6414 (N_6414,N_5690,N_5991);
nor U6415 (N_6415,N_5962,N_5573);
or U6416 (N_6416,N_5768,N_5633);
or U6417 (N_6417,N_5795,N_5737);
nand U6418 (N_6418,N_5808,N_5668);
xor U6419 (N_6419,N_5928,N_5921);
nand U6420 (N_6420,N_5982,N_5657);
xnor U6421 (N_6421,N_5632,N_5774);
xor U6422 (N_6422,N_5995,N_5630);
and U6423 (N_6423,N_5534,N_5580);
or U6424 (N_6424,N_5936,N_5548);
or U6425 (N_6425,N_5752,N_5801);
or U6426 (N_6426,N_5894,N_5713);
nand U6427 (N_6427,N_5860,N_5595);
nand U6428 (N_6428,N_5805,N_5762);
nand U6429 (N_6429,N_5712,N_5509);
and U6430 (N_6430,N_5852,N_5582);
nor U6431 (N_6431,N_5775,N_5886);
or U6432 (N_6432,N_5619,N_5808);
nand U6433 (N_6433,N_5821,N_5869);
nor U6434 (N_6434,N_5911,N_5869);
xor U6435 (N_6435,N_5649,N_5639);
xnor U6436 (N_6436,N_5932,N_5919);
nand U6437 (N_6437,N_5652,N_5923);
nand U6438 (N_6438,N_5893,N_5746);
or U6439 (N_6439,N_5874,N_5762);
and U6440 (N_6440,N_5678,N_5619);
xnor U6441 (N_6441,N_5733,N_5601);
and U6442 (N_6442,N_5713,N_5595);
nor U6443 (N_6443,N_5549,N_5691);
or U6444 (N_6444,N_5598,N_5834);
xnor U6445 (N_6445,N_5908,N_5855);
xor U6446 (N_6446,N_5731,N_5537);
nor U6447 (N_6447,N_5541,N_5706);
or U6448 (N_6448,N_5562,N_5817);
nor U6449 (N_6449,N_5602,N_5947);
or U6450 (N_6450,N_5857,N_5970);
nand U6451 (N_6451,N_5564,N_5903);
and U6452 (N_6452,N_5653,N_5880);
and U6453 (N_6453,N_5520,N_5795);
nor U6454 (N_6454,N_5939,N_5854);
and U6455 (N_6455,N_5815,N_5731);
nand U6456 (N_6456,N_5939,N_5628);
xor U6457 (N_6457,N_5692,N_5602);
nor U6458 (N_6458,N_5949,N_5912);
or U6459 (N_6459,N_5581,N_5888);
nand U6460 (N_6460,N_5952,N_5918);
nand U6461 (N_6461,N_5692,N_5641);
nand U6462 (N_6462,N_5751,N_5582);
and U6463 (N_6463,N_5959,N_5696);
xnor U6464 (N_6464,N_5715,N_5817);
xnor U6465 (N_6465,N_5795,N_5740);
xnor U6466 (N_6466,N_5945,N_5744);
and U6467 (N_6467,N_5798,N_5685);
nand U6468 (N_6468,N_5932,N_5607);
nand U6469 (N_6469,N_5729,N_5580);
xor U6470 (N_6470,N_5752,N_5867);
or U6471 (N_6471,N_5706,N_5786);
nor U6472 (N_6472,N_5888,N_5992);
or U6473 (N_6473,N_5924,N_5996);
and U6474 (N_6474,N_5616,N_5553);
and U6475 (N_6475,N_5717,N_5962);
and U6476 (N_6476,N_5898,N_5753);
or U6477 (N_6477,N_5792,N_5744);
nor U6478 (N_6478,N_5974,N_5591);
nor U6479 (N_6479,N_5589,N_5977);
or U6480 (N_6480,N_5593,N_5988);
and U6481 (N_6481,N_5772,N_5570);
nand U6482 (N_6482,N_5780,N_5605);
and U6483 (N_6483,N_5636,N_5818);
nand U6484 (N_6484,N_5660,N_5978);
xor U6485 (N_6485,N_5569,N_5819);
nor U6486 (N_6486,N_5962,N_5519);
xnor U6487 (N_6487,N_5942,N_5875);
nand U6488 (N_6488,N_5628,N_5955);
or U6489 (N_6489,N_5676,N_5847);
or U6490 (N_6490,N_5886,N_5617);
nor U6491 (N_6491,N_5551,N_5882);
xnor U6492 (N_6492,N_5534,N_5840);
nor U6493 (N_6493,N_5978,N_5629);
xor U6494 (N_6494,N_5657,N_5607);
xor U6495 (N_6495,N_5542,N_5978);
nand U6496 (N_6496,N_5623,N_5921);
and U6497 (N_6497,N_5955,N_5760);
or U6498 (N_6498,N_5549,N_5748);
xor U6499 (N_6499,N_5804,N_5788);
and U6500 (N_6500,N_6067,N_6439);
nand U6501 (N_6501,N_6109,N_6223);
nor U6502 (N_6502,N_6485,N_6353);
nand U6503 (N_6503,N_6203,N_6409);
or U6504 (N_6504,N_6257,N_6123);
or U6505 (N_6505,N_6086,N_6133);
and U6506 (N_6506,N_6476,N_6204);
or U6507 (N_6507,N_6225,N_6479);
or U6508 (N_6508,N_6141,N_6105);
xnor U6509 (N_6509,N_6000,N_6333);
nor U6510 (N_6510,N_6192,N_6402);
nand U6511 (N_6511,N_6443,N_6101);
or U6512 (N_6512,N_6156,N_6302);
xor U6513 (N_6513,N_6447,N_6279);
and U6514 (N_6514,N_6200,N_6288);
nor U6515 (N_6515,N_6088,N_6209);
nor U6516 (N_6516,N_6287,N_6326);
or U6517 (N_6517,N_6382,N_6037);
nor U6518 (N_6518,N_6117,N_6325);
nor U6519 (N_6519,N_6280,N_6072);
xnor U6520 (N_6520,N_6081,N_6051);
nand U6521 (N_6521,N_6172,N_6110);
and U6522 (N_6522,N_6481,N_6456);
and U6523 (N_6523,N_6189,N_6301);
nor U6524 (N_6524,N_6313,N_6399);
and U6525 (N_6525,N_6422,N_6036);
xnor U6526 (N_6526,N_6102,N_6059);
or U6527 (N_6527,N_6263,N_6367);
nand U6528 (N_6528,N_6342,N_6498);
nor U6529 (N_6529,N_6258,N_6355);
and U6530 (N_6530,N_6347,N_6079);
nor U6531 (N_6531,N_6467,N_6094);
and U6532 (N_6532,N_6416,N_6398);
nor U6533 (N_6533,N_6457,N_6495);
nor U6534 (N_6534,N_6145,N_6368);
and U6535 (N_6535,N_6262,N_6320);
nand U6536 (N_6536,N_6104,N_6232);
or U6537 (N_6537,N_6208,N_6369);
nand U6538 (N_6538,N_6264,N_6354);
nand U6539 (N_6539,N_6162,N_6274);
nand U6540 (N_6540,N_6103,N_6154);
xor U6541 (N_6541,N_6095,N_6484);
xnor U6542 (N_6542,N_6337,N_6230);
xnor U6543 (N_6543,N_6020,N_6489);
nor U6544 (N_6544,N_6229,N_6240);
xor U6545 (N_6545,N_6047,N_6314);
xor U6546 (N_6546,N_6419,N_6214);
xor U6547 (N_6547,N_6448,N_6480);
and U6548 (N_6548,N_6423,N_6030);
and U6549 (N_6549,N_6207,N_6217);
or U6550 (N_6550,N_6271,N_6384);
xnor U6551 (N_6551,N_6268,N_6055);
nand U6552 (N_6552,N_6159,N_6026);
or U6553 (N_6553,N_6491,N_6074);
nor U6554 (N_6554,N_6089,N_6222);
or U6555 (N_6555,N_6451,N_6391);
nand U6556 (N_6556,N_6310,N_6362);
nor U6557 (N_6557,N_6256,N_6176);
and U6558 (N_6558,N_6064,N_6373);
or U6559 (N_6559,N_6085,N_6116);
or U6560 (N_6560,N_6188,N_6428);
nor U6561 (N_6561,N_6323,N_6125);
nor U6562 (N_6562,N_6475,N_6245);
or U6563 (N_6563,N_6374,N_6294);
and U6564 (N_6564,N_6282,N_6427);
or U6565 (N_6565,N_6458,N_6297);
nor U6566 (N_6566,N_6014,N_6041);
or U6567 (N_6567,N_6388,N_6468);
and U6568 (N_6568,N_6164,N_6330);
xnor U6569 (N_6569,N_6408,N_6472);
or U6570 (N_6570,N_6140,N_6052);
xnor U6571 (N_6571,N_6437,N_6238);
and U6572 (N_6572,N_6487,N_6289);
xor U6573 (N_6573,N_6254,N_6380);
nor U6574 (N_6574,N_6370,N_6108);
nand U6575 (N_6575,N_6197,N_6425);
nand U6576 (N_6576,N_6132,N_6025);
xor U6577 (N_6577,N_6194,N_6247);
and U6578 (N_6578,N_6273,N_6016);
xnor U6579 (N_6579,N_6115,N_6019);
or U6580 (N_6580,N_6007,N_6334);
xnor U6581 (N_6581,N_6364,N_6168);
nand U6582 (N_6582,N_6376,N_6069);
xor U6583 (N_6583,N_6415,N_6488);
nor U6584 (N_6584,N_6292,N_6252);
nand U6585 (N_6585,N_6177,N_6058);
xor U6586 (N_6586,N_6351,N_6122);
nand U6587 (N_6587,N_6454,N_6028);
nand U6588 (N_6588,N_6411,N_6446);
nor U6589 (N_6589,N_6253,N_6449);
or U6590 (N_6590,N_6331,N_6191);
xnor U6591 (N_6591,N_6358,N_6434);
or U6592 (N_6592,N_6265,N_6002);
xor U6593 (N_6593,N_6250,N_6015);
nand U6594 (N_6594,N_6436,N_6234);
or U6595 (N_6595,N_6006,N_6082);
and U6596 (N_6596,N_6352,N_6295);
nor U6597 (N_6597,N_6012,N_6486);
xor U6598 (N_6598,N_6004,N_6236);
and U6599 (N_6599,N_6142,N_6226);
nand U6600 (N_6600,N_6414,N_6417);
xnor U6601 (N_6601,N_6442,N_6385);
or U6602 (N_6602,N_6185,N_6182);
nor U6603 (N_6603,N_6111,N_6260);
or U6604 (N_6604,N_6336,N_6403);
xor U6605 (N_6605,N_6453,N_6034);
xor U6606 (N_6606,N_6418,N_6243);
xor U6607 (N_6607,N_6119,N_6056);
nor U6608 (N_6608,N_6220,N_6219);
nor U6609 (N_6609,N_6163,N_6013);
nand U6610 (N_6610,N_6100,N_6131);
and U6611 (N_6611,N_6474,N_6401);
xor U6612 (N_6612,N_6068,N_6075);
xnor U6613 (N_6613,N_6478,N_6477);
nand U6614 (N_6614,N_6461,N_6039);
or U6615 (N_6615,N_6450,N_6193);
and U6616 (N_6616,N_6357,N_6057);
and U6617 (N_6617,N_6270,N_6393);
xnor U6618 (N_6618,N_6251,N_6304);
nor U6619 (N_6619,N_6285,N_6024);
nand U6620 (N_6620,N_6078,N_6473);
nand U6621 (N_6621,N_6017,N_6183);
nor U6622 (N_6622,N_6235,N_6202);
xor U6623 (N_6623,N_6483,N_6216);
or U6624 (N_6624,N_6308,N_6315);
or U6625 (N_6625,N_6490,N_6063);
and U6626 (N_6626,N_6341,N_6113);
nand U6627 (N_6627,N_6377,N_6212);
xor U6628 (N_6628,N_6213,N_6150);
nor U6629 (N_6629,N_6307,N_6322);
or U6630 (N_6630,N_6345,N_6317);
nand U6631 (N_6631,N_6494,N_6171);
xnor U6632 (N_6632,N_6174,N_6405);
nor U6633 (N_6633,N_6379,N_6206);
nand U6634 (N_6634,N_6137,N_6309);
or U6635 (N_6635,N_6211,N_6138);
or U6636 (N_6636,N_6077,N_6165);
nand U6637 (N_6637,N_6239,N_6143);
nor U6638 (N_6638,N_6318,N_6149);
xor U6639 (N_6639,N_6018,N_6210);
or U6640 (N_6640,N_6107,N_6244);
and U6641 (N_6641,N_6413,N_6324);
xnor U6642 (N_6642,N_6184,N_6255);
and U6643 (N_6643,N_6361,N_6412);
xor U6644 (N_6644,N_6146,N_6196);
nor U6645 (N_6645,N_6462,N_6332);
xor U6646 (N_6646,N_6091,N_6126);
nand U6647 (N_6647,N_6061,N_6346);
nand U6648 (N_6648,N_6375,N_6042);
and U6649 (N_6649,N_6135,N_6452);
and U6650 (N_6650,N_6060,N_6070);
nand U6651 (N_6651,N_6033,N_6387);
nand U6652 (N_6652,N_6073,N_6106);
nand U6653 (N_6653,N_6249,N_6180);
and U6654 (N_6654,N_6350,N_6464);
or U6655 (N_6655,N_6435,N_6493);
nor U6656 (N_6656,N_6029,N_6492);
or U6657 (N_6657,N_6242,N_6035);
xor U6658 (N_6658,N_6366,N_6083);
and U6659 (N_6659,N_6394,N_6008);
xnor U6660 (N_6660,N_6306,N_6460);
nor U6661 (N_6661,N_6321,N_6097);
or U6662 (N_6662,N_6429,N_6118);
nor U6663 (N_6663,N_6300,N_6343);
nand U6664 (N_6664,N_6062,N_6023);
xnor U6665 (N_6665,N_6372,N_6269);
nand U6666 (N_6666,N_6084,N_6397);
nand U6667 (N_6667,N_6166,N_6124);
nor U6668 (N_6668,N_6360,N_6195);
nor U6669 (N_6669,N_6134,N_6231);
or U6670 (N_6670,N_6395,N_6046);
xor U6671 (N_6671,N_6120,N_6406);
xnor U6672 (N_6672,N_6031,N_6112);
nand U6673 (N_6673,N_6291,N_6303);
nand U6674 (N_6674,N_6128,N_6246);
xor U6675 (N_6675,N_6227,N_6499);
nand U6676 (N_6676,N_6040,N_6179);
and U6677 (N_6677,N_6283,N_6396);
or U6678 (N_6678,N_6293,N_6050);
nor U6679 (N_6679,N_6277,N_6432);
nand U6680 (N_6680,N_6275,N_6121);
or U6681 (N_6681,N_6298,N_6400);
nand U6682 (N_6682,N_6001,N_6378);
nand U6683 (N_6683,N_6440,N_6459);
and U6684 (N_6684,N_6129,N_6224);
nor U6685 (N_6685,N_6363,N_6153);
nor U6686 (N_6686,N_6139,N_6045);
nor U6687 (N_6687,N_6173,N_6284);
and U6688 (N_6688,N_6096,N_6114);
or U6689 (N_6689,N_6038,N_6455);
nor U6690 (N_6690,N_6421,N_6438);
and U6691 (N_6691,N_6444,N_6259);
or U6692 (N_6692,N_6158,N_6261);
nand U6693 (N_6693,N_6130,N_6092);
or U6694 (N_6694,N_6445,N_6186);
or U6695 (N_6695,N_6410,N_6248);
nor U6696 (N_6696,N_6344,N_6148);
nor U6697 (N_6697,N_6152,N_6349);
and U6698 (N_6698,N_6497,N_6328);
or U6699 (N_6699,N_6144,N_6340);
and U6700 (N_6700,N_6312,N_6147);
xor U6701 (N_6701,N_6470,N_6087);
xnor U6702 (N_6702,N_6076,N_6272);
or U6703 (N_6703,N_6431,N_6299);
xor U6704 (N_6704,N_6199,N_6228);
and U6705 (N_6705,N_6441,N_6065);
nor U6706 (N_6706,N_6286,N_6335);
nor U6707 (N_6707,N_6010,N_6338);
xnor U6708 (N_6708,N_6215,N_6003);
nand U6709 (N_6709,N_6266,N_6161);
or U6710 (N_6710,N_6407,N_6430);
or U6711 (N_6711,N_6027,N_6359);
and U6712 (N_6712,N_6469,N_6044);
or U6713 (N_6713,N_6383,N_6316);
or U6714 (N_6714,N_6276,N_6049);
xnor U6715 (N_6715,N_6021,N_6433);
nand U6716 (N_6716,N_6099,N_6201);
and U6717 (N_6717,N_6424,N_6011);
nand U6718 (N_6718,N_6319,N_6281);
or U6719 (N_6719,N_6386,N_6233);
or U6720 (N_6720,N_6426,N_6181);
nor U6721 (N_6721,N_6496,N_6290);
nor U6722 (N_6722,N_6218,N_6169);
xor U6723 (N_6723,N_6389,N_6160);
and U6724 (N_6724,N_6190,N_6296);
xor U6725 (N_6725,N_6365,N_6167);
xnor U6726 (N_6726,N_6043,N_6466);
and U6727 (N_6727,N_6066,N_6032);
nand U6728 (N_6728,N_6221,N_6267);
nand U6729 (N_6729,N_6371,N_6127);
and U6730 (N_6730,N_6465,N_6053);
or U6731 (N_6731,N_6009,N_6327);
xnor U6732 (N_6732,N_6348,N_6155);
and U6733 (N_6733,N_6157,N_6420);
nand U6734 (N_6734,N_6237,N_6381);
xor U6735 (N_6735,N_6356,N_6339);
xor U6736 (N_6736,N_6205,N_6241);
or U6737 (N_6737,N_6175,N_6005);
or U6738 (N_6738,N_6392,N_6404);
nor U6739 (N_6739,N_6311,N_6178);
nand U6740 (N_6740,N_6305,N_6170);
or U6741 (N_6741,N_6390,N_6151);
or U6742 (N_6742,N_6482,N_6054);
or U6743 (N_6743,N_6463,N_6098);
nand U6744 (N_6744,N_6048,N_6022);
nor U6745 (N_6745,N_6187,N_6071);
nand U6746 (N_6746,N_6471,N_6198);
nand U6747 (N_6747,N_6329,N_6090);
xnor U6748 (N_6748,N_6278,N_6080);
nor U6749 (N_6749,N_6093,N_6136);
nor U6750 (N_6750,N_6037,N_6270);
nand U6751 (N_6751,N_6451,N_6085);
or U6752 (N_6752,N_6365,N_6131);
and U6753 (N_6753,N_6364,N_6459);
nand U6754 (N_6754,N_6384,N_6317);
and U6755 (N_6755,N_6354,N_6307);
nor U6756 (N_6756,N_6209,N_6429);
nor U6757 (N_6757,N_6210,N_6286);
xor U6758 (N_6758,N_6312,N_6355);
and U6759 (N_6759,N_6465,N_6354);
and U6760 (N_6760,N_6353,N_6116);
nand U6761 (N_6761,N_6355,N_6088);
and U6762 (N_6762,N_6455,N_6493);
or U6763 (N_6763,N_6247,N_6181);
xnor U6764 (N_6764,N_6330,N_6096);
xor U6765 (N_6765,N_6324,N_6357);
xor U6766 (N_6766,N_6372,N_6452);
nor U6767 (N_6767,N_6168,N_6432);
or U6768 (N_6768,N_6175,N_6133);
xnor U6769 (N_6769,N_6388,N_6319);
nor U6770 (N_6770,N_6478,N_6000);
nand U6771 (N_6771,N_6085,N_6437);
nor U6772 (N_6772,N_6202,N_6238);
nor U6773 (N_6773,N_6451,N_6307);
or U6774 (N_6774,N_6183,N_6269);
and U6775 (N_6775,N_6450,N_6092);
xor U6776 (N_6776,N_6088,N_6253);
or U6777 (N_6777,N_6100,N_6110);
and U6778 (N_6778,N_6033,N_6269);
xnor U6779 (N_6779,N_6121,N_6473);
and U6780 (N_6780,N_6377,N_6173);
or U6781 (N_6781,N_6452,N_6423);
or U6782 (N_6782,N_6398,N_6393);
xnor U6783 (N_6783,N_6373,N_6172);
nor U6784 (N_6784,N_6064,N_6377);
nor U6785 (N_6785,N_6271,N_6138);
or U6786 (N_6786,N_6303,N_6400);
or U6787 (N_6787,N_6255,N_6336);
xor U6788 (N_6788,N_6454,N_6378);
or U6789 (N_6789,N_6098,N_6466);
nand U6790 (N_6790,N_6351,N_6387);
nor U6791 (N_6791,N_6405,N_6353);
or U6792 (N_6792,N_6375,N_6022);
and U6793 (N_6793,N_6120,N_6240);
xor U6794 (N_6794,N_6155,N_6258);
xnor U6795 (N_6795,N_6384,N_6098);
nand U6796 (N_6796,N_6240,N_6038);
and U6797 (N_6797,N_6285,N_6349);
nand U6798 (N_6798,N_6424,N_6279);
nand U6799 (N_6799,N_6496,N_6403);
nand U6800 (N_6800,N_6034,N_6452);
xnor U6801 (N_6801,N_6097,N_6370);
nand U6802 (N_6802,N_6267,N_6118);
and U6803 (N_6803,N_6412,N_6431);
or U6804 (N_6804,N_6157,N_6338);
nand U6805 (N_6805,N_6418,N_6170);
and U6806 (N_6806,N_6009,N_6339);
or U6807 (N_6807,N_6231,N_6090);
and U6808 (N_6808,N_6257,N_6039);
and U6809 (N_6809,N_6376,N_6438);
and U6810 (N_6810,N_6128,N_6038);
xor U6811 (N_6811,N_6110,N_6030);
xor U6812 (N_6812,N_6256,N_6044);
or U6813 (N_6813,N_6429,N_6449);
and U6814 (N_6814,N_6010,N_6068);
and U6815 (N_6815,N_6478,N_6331);
and U6816 (N_6816,N_6375,N_6426);
and U6817 (N_6817,N_6160,N_6345);
and U6818 (N_6818,N_6175,N_6117);
or U6819 (N_6819,N_6461,N_6465);
nand U6820 (N_6820,N_6310,N_6392);
or U6821 (N_6821,N_6421,N_6446);
xnor U6822 (N_6822,N_6248,N_6307);
and U6823 (N_6823,N_6275,N_6374);
xor U6824 (N_6824,N_6089,N_6014);
or U6825 (N_6825,N_6344,N_6191);
xnor U6826 (N_6826,N_6100,N_6252);
nand U6827 (N_6827,N_6005,N_6202);
and U6828 (N_6828,N_6447,N_6452);
and U6829 (N_6829,N_6127,N_6475);
xor U6830 (N_6830,N_6365,N_6478);
and U6831 (N_6831,N_6159,N_6070);
xnor U6832 (N_6832,N_6116,N_6251);
or U6833 (N_6833,N_6209,N_6326);
or U6834 (N_6834,N_6421,N_6327);
or U6835 (N_6835,N_6144,N_6200);
and U6836 (N_6836,N_6093,N_6261);
nand U6837 (N_6837,N_6193,N_6063);
nor U6838 (N_6838,N_6397,N_6380);
xor U6839 (N_6839,N_6435,N_6380);
nor U6840 (N_6840,N_6451,N_6328);
and U6841 (N_6841,N_6237,N_6459);
nand U6842 (N_6842,N_6450,N_6232);
nor U6843 (N_6843,N_6210,N_6268);
nand U6844 (N_6844,N_6488,N_6310);
and U6845 (N_6845,N_6247,N_6227);
and U6846 (N_6846,N_6456,N_6161);
nand U6847 (N_6847,N_6171,N_6106);
nor U6848 (N_6848,N_6446,N_6427);
or U6849 (N_6849,N_6415,N_6335);
and U6850 (N_6850,N_6077,N_6281);
xor U6851 (N_6851,N_6162,N_6060);
nand U6852 (N_6852,N_6465,N_6457);
nand U6853 (N_6853,N_6418,N_6304);
or U6854 (N_6854,N_6206,N_6064);
nand U6855 (N_6855,N_6240,N_6262);
nor U6856 (N_6856,N_6353,N_6133);
xnor U6857 (N_6857,N_6067,N_6225);
xnor U6858 (N_6858,N_6301,N_6175);
and U6859 (N_6859,N_6271,N_6473);
or U6860 (N_6860,N_6486,N_6221);
and U6861 (N_6861,N_6065,N_6193);
nor U6862 (N_6862,N_6254,N_6136);
nand U6863 (N_6863,N_6241,N_6095);
xor U6864 (N_6864,N_6448,N_6214);
and U6865 (N_6865,N_6364,N_6273);
xnor U6866 (N_6866,N_6165,N_6139);
nand U6867 (N_6867,N_6263,N_6129);
and U6868 (N_6868,N_6075,N_6166);
or U6869 (N_6869,N_6352,N_6209);
nand U6870 (N_6870,N_6261,N_6281);
nand U6871 (N_6871,N_6205,N_6178);
nand U6872 (N_6872,N_6436,N_6220);
and U6873 (N_6873,N_6312,N_6089);
nand U6874 (N_6874,N_6303,N_6073);
or U6875 (N_6875,N_6227,N_6035);
and U6876 (N_6876,N_6253,N_6320);
nand U6877 (N_6877,N_6477,N_6448);
or U6878 (N_6878,N_6192,N_6134);
and U6879 (N_6879,N_6445,N_6420);
and U6880 (N_6880,N_6149,N_6330);
nor U6881 (N_6881,N_6371,N_6421);
xnor U6882 (N_6882,N_6472,N_6393);
and U6883 (N_6883,N_6344,N_6491);
xnor U6884 (N_6884,N_6034,N_6467);
nor U6885 (N_6885,N_6329,N_6426);
or U6886 (N_6886,N_6153,N_6132);
or U6887 (N_6887,N_6476,N_6104);
xor U6888 (N_6888,N_6211,N_6002);
nand U6889 (N_6889,N_6468,N_6499);
nand U6890 (N_6890,N_6488,N_6324);
and U6891 (N_6891,N_6390,N_6065);
nand U6892 (N_6892,N_6468,N_6039);
and U6893 (N_6893,N_6086,N_6262);
nand U6894 (N_6894,N_6026,N_6123);
or U6895 (N_6895,N_6419,N_6205);
xnor U6896 (N_6896,N_6476,N_6148);
nor U6897 (N_6897,N_6208,N_6189);
and U6898 (N_6898,N_6374,N_6256);
xnor U6899 (N_6899,N_6139,N_6030);
xnor U6900 (N_6900,N_6153,N_6347);
and U6901 (N_6901,N_6278,N_6150);
nand U6902 (N_6902,N_6339,N_6225);
nand U6903 (N_6903,N_6277,N_6354);
or U6904 (N_6904,N_6333,N_6121);
nor U6905 (N_6905,N_6406,N_6389);
nand U6906 (N_6906,N_6118,N_6108);
nand U6907 (N_6907,N_6139,N_6192);
nand U6908 (N_6908,N_6150,N_6420);
nor U6909 (N_6909,N_6409,N_6134);
nand U6910 (N_6910,N_6412,N_6382);
xor U6911 (N_6911,N_6440,N_6236);
nor U6912 (N_6912,N_6388,N_6288);
and U6913 (N_6913,N_6139,N_6305);
nor U6914 (N_6914,N_6186,N_6167);
or U6915 (N_6915,N_6012,N_6132);
nor U6916 (N_6916,N_6469,N_6252);
or U6917 (N_6917,N_6452,N_6104);
xnor U6918 (N_6918,N_6188,N_6482);
nand U6919 (N_6919,N_6412,N_6167);
xnor U6920 (N_6920,N_6098,N_6100);
and U6921 (N_6921,N_6358,N_6306);
and U6922 (N_6922,N_6120,N_6476);
and U6923 (N_6923,N_6417,N_6203);
xnor U6924 (N_6924,N_6080,N_6214);
and U6925 (N_6925,N_6026,N_6196);
nand U6926 (N_6926,N_6468,N_6347);
and U6927 (N_6927,N_6036,N_6170);
nor U6928 (N_6928,N_6114,N_6270);
xor U6929 (N_6929,N_6107,N_6147);
or U6930 (N_6930,N_6404,N_6015);
or U6931 (N_6931,N_6069,N_6306);
and U6932 (N_6932,N_6114,N_6397);
nor U6933 (N_6933,N_6488,N_6198);
and U6934 (N_6934,N_6180,N_6392);
or U6935 (N_6935,N_6383,N_6161);
and U6936 (N_6936,N_6067,N_6278);
or U6937 (N_6937,N_6087,N_6272);
xnor U6938 (N_6938,N_6279,N_6021);
nor U6939 (N_6939,N_6098,N_6004);
xnor U6940 (N_6940,N_6314,N_6118);
nand U6941 (N_6941,N_6136,N_6459);
xor U6942 (N_6942,N_6156,N_6332);
nand U6943 (N_6943,N_6158,N_6462);
nor U6944 (N_6944,N_6302,N_6487);
nand U6945 (N_6945,N_6418,N_6038);
and U6946 (N_6946,N_6175,N_6178);
or U6947 (N_6947,N_6348,N_6118);
or U6948 (N_6948,N_6144,N_6149);
xnor U6949 (N_6949,N_6437,N_6098);
or U6950 (N_6950,N_6053,N_6381);
nor U6951 (N_6951,N_6357,N_6141);
nand U6952 (N_6952,N_6292,N_6115);
nor U6953 (N_6953,N_6324,N_6093);
nor U6954 (N_6954,N_6201,N_6409);
nand U6955 (N_6955,N_6365,N_6472);
and U6956 (N_6956,N_6471,N_6151);
or U6957 (N_6957,N_6121,N_6097);
or U6958 (N_6958,N_6444,N_6391);
or U6959 (N_6959,N_6130,N_6010);
nor U6960 (N_6960,N_6408,N_6412);
xnor U6961 (N_6961,N_6380,N_6457);
or U6962 (N_6962,N_6452,N_6049);
nand U6963 (N_6963,N_6358,N_6281);
and U6964 (N_6964,N_6033,N_6054);
or U6965 (N_6965,N_6164,N_6055);
nor U6966 (N_6966,N_6306,N_6101);
nor U6967 (N_6967,N_6405,N_6396);
nor U6968 (N_6968,N_6073,N_6471);
and U6969 (N_6969,N_6029,N_6458);
nand U6970 (N_6970,N_6321,N_6090);
nand U6971 (N_6971,N_6263,N_6039);
and U6972 (N_6972,N_6166,N_6174);
xor U6973 (N_6973,N_6090,N_6019);
or U6974 (N_6974,N_6186,N_6391);
nor U6975 (N_6975,N_6171,N_6317);
or U6976 (N_6976,N_6484,N_6145);
xor U6977 (N_6977,N_6430,N_6230);
nand U6978 (N_6978,N_6289,N_6129);
nor U6979 (N_6979,N_6420,N_6308);
and U6980 (N_6980,N_6342,N_6248);
and U6981 (N_6981,N_6418,N_6466);
or U6982 (N_6982,N_6466,N_6277);
xnor U6983 (N_6983,N_6140,N_6065);
and U6984 (N_6984,N_6166,N_6315);
xor U6985 (N_6985,N_6256,N_6397);
nor U6986 (N_6986,N_6159,N_6231);
nor U6987 (N_6987,N_6216,N_6080);
nor U6988 (N_6988,N_6033,N_6022);
nor U6989 (N_6989,N_6101,N_6217);
or U6990 (N_6990,N_6109,N_6142);
and U6991 (N_6991,N_6037,N_6348);
xor U6992 (N_6992,N_6364,N_6179);
nand U6993 (N_6993,N_6149,N_6218);
nor U6994 (N_6994,N_6259,N_6179);
nand U6995 (N_6995,N_6188,N_6268);
xor U6996 (N_6996,N_6179,N_6431);
or U6997 (N_6997,N_6181,N_6052);
or U6998 (N_6998,N_6204,N_6424);
or U6999 (N_6999,N_6199,N_6447);
and U7000 (N_7000,N_6609,N_6687);
nand U7001 (N_7001,N_6994,N_6971);
nor U7002 (N_7002,N_6969,N_6879);
or U7003 (N_7003,N_6912,N_6800);
xnor U7004 (N_7004,N_6831,N_6787);
and U7005 (N_7005,N_6623,N_6773);
and U7006 (N_7006,N_6607,N_6728);
and U7007 (N_7007,N_6677,N_6752);
xnor U7008 (N_7008,N_6931,N_6901);
and U7009 (N_7009,N_6727,N_6759);
nor U7010 (N_7010,N_6576,N_6970);
or U7011 (N_7011,N_6988,N_6921);
nor U7012 (N_7012,N_6881,N_6649);
or U7013 (N_7013,N_6980,N_6619);
or U7014 (N_7014,N_6720,N_6534);
nand U7015 (N_7015,N_6566,N_6679);
nand U7016 (N_7016,N_6716,N_6575);
and U7017 (N_7017,N_6648,N_6775);
and U7018 (N_7018,N_6768,N_6870);
or U7019 (N_7019,N_6662,N_6674);
nand U7020 (N_7020,N_6528,N_6794);
and U7021 (N_7021,N_6793,N_6580);
xnor U7022 (N_7022,N_6976,N_6890);
xnor U7023 (N_7023,N_6837,N_6610);
and U7024 (N_7024,N_6908,N_6981);
xor U7025 (N_7025,N_6854,N_6845);
or U7026 (N_7026,N_6832,N_6664);
or U7027 (N_7027,N_6585,N_6671);
or U7028 (N_7028,N_6710,N_6742);
and U7029 (N_7029,N_6657,N_6616);
xnor U7030 (N_7030,N_6629,N_6659);
nand U7031 (N_7031,N_6626,N_6920);
nor U7032 (N_7032,N_6911,N_6945);
and U7033 (N_7033,N_6681,N_6682);
xor U7034 (N_7034,N_6544,N_6586);
xnor U7035 (N_7035,N_6798,N_6507);
nand U7036 (N_7036,N_6871,N_6909);
and U7037 (N_7037,N_6696,N_6725);
nand U7038 (N_7038,N_6836,N_6884);
or U7039 (N_7039,N_6972,N_6606);
nand U7040 (N_7040,N_6982,N_6844);
nor U7041 (N_7041,N_6525,N_6906);
nand U7042 (N_7042,N_6635,N_6695);
nor U7043 (N_7043,N_6964,N_6955);
xnor U7044 (N_7044,N_6591,N_6676);
or U7045 (N_7045,N_6579,N_6833);
or U7046 (N_7046,N_6552,N_6807);
xor U7047 (N_7047,N_6786,N_6622);
and U7048 (N_7048,N_6847,N_6509);
nor U7049 (N_7049,N_6843,N_6684);
xnor U7050 (N_7050,N_6957,N_6590);
or U7051 (N_7051,N_6803,N_6743);
or U7052 (N_7052,N_6875,N_6708);
and U7053 (N_7053,N_6531,N_6526);
and U7054 (N_7054,N_6925,N_6675);
nor U7055 (N_7055,N_6949,N_6650);
or U7056 (N_7056,N_6736,N_6732);
nand U7057 (N_7057,N_6688,N_6809);
xnor U7058 (N_7058,N_6919,N_6788);
nand U7059 (N_7059,N_6571,N_6930);
nand U7060 (N_7060,N_6717,N_6715);
xnor U7061 (N_7061,N_6838,N_6733);
xor U7062 (N_7062,N_6928,N_6532);
and U7063 (N_7063,N_6781,N_6588);
and U7064 (N_7064,N_6817,N_6501);
nor U7065 (N_7065,N_6864,N_6791);
or U7066 (N_7066,N_6738,N_6802);
and U7067 (N_7067,N_6608,N_6652);
or U7068 (N_7068,N_6685,N_6850);
or U7069 (N_7069,N_6672,N_6617);
nand U7070 (N_7070,N_6853,N_6667);
xnor U7071 (N_7071,N_6641,N_6943);
xnor U7072 (N_7072,N_6751,N_6618);
nand U7073 (N_7073,N_6706,N_6973);
and U7074 (N_7074,N_6562,N_6805);
xnor U7075 (N_7075,N_6842,N_6886);
and U7076 (N_7076,N_6907,N_6746);
nand U7077 (N_7077,N_6916,N_6653);
and U7078 (N_7078,N_6523,N_6551);
nand U7079 (N_7079,N_6554,N_6730);
nand U7080 (N_7080,N_6574,N_6997);
nor U7081 (N_7081,N_6801,N_6922);
and U7082 (N_7082,N_6582,N_6663);
and U7083 (N_7083,N_6874,N_6992);
xnor U7084 (N_7084,N_6785,N_6859);
nor U7085 (N_7085,N_6754,N_6639);
or U7086 (N_7086,N_6863,N_6968);
nand U7087 (N_7087,N_6985,N_6600);
nand U7088 (N_7088,N_6578,N_6683);
and U7089 (N_7089,N_6790,N_6612);
and U7090 (N_7090,N_6570,N_6825);
and U7091 (N_7091,N_6535,N_6573);
xor U7092 (N_7092,N_6839,N_6537);
nor U7093 (N_7093,N_6504,N_6821);
xor U7094 (N_7094,N_6974,N_6789);
and U7095 (N_7095,N_6757,N_6515);
or U7096 (N_7096,N_6915,N_6548);
xor U7097 (N_7097,N_6950,N_6624);
xor U7098 (N_7098,N_6638,N_6704);
nand U7099 (N_7099,N_6699,N_6512);
xnor U7100 (N_7100,N_6707,N_6745);
nor U7101 (N_7101,N_6977,N_6934);
nand U7102 (N_7102,N_6940,N_6904);
xnor U7103 (N_7103,N_6991,N_6959);
and U7104 (N_7104,N_6818,N_6656);
and U7105 (N_7105,N_6625,N_6633);
nor U7106 (N_7106,N_6953,N_6691);
nand U7107 (N_7107,N_6929,N_6690);
nor U7108 (N_7108,N_6866,N_6729);
xnor U7109 (N_7109,N_6520,N_6924);
nor U7110 (N_7110,N_6851,N_6846);
xnor U7111 (N_7111,N_6748,N_6651);
and U7112 (N_7112,N_6714,N_6894);
xnor U7113 (N_7113,N_6694,N_6712);
nand U7114 (N_7114,N_6880,N_6883);
and U7115 (N_7115,N_6784,N_6634);
nor U7116 (N_7116,N_6860,N_6819);
xnor U7117 (N_7117,N_6693,N_6952);
nor U7118 (N_7118,N_6776,N_6724);
and U7119 (N_7119,N_6975,N_6830);
xnor U7120 (N_7120,N_6778,N_6636);
nand U7121 (N_7121,N_6810,N_6902);
nor U7122 (N_7122,N_6637,N_6530);
xnor U7123 (N_7123,N_6923,N_6852);
or U7124 (N_7124,N_6877,N_6581);
or U7125 (N_7125,N_6686,N_6918);
nor U7126 (N_7126,N_6967,N_6739);
and U7127 (N_7127,N_6654,N_6620);
or U7128 (N_7128,N_6927,N_6896);
and U7129 (N_7129,N_6521,N_6673);
nand U7130 (N_7130,N_6697,N_6948);
or U7131 (N_7131,N_6557,N_6529);
or U7132 (N_7132,N_6848,N_6995);
xor U7133 (N_7133,N_6737,N_6646);
xor U7134 (N_7134,N_6627,N_6893);
or U7135 (N_7135,N_6841,N_6577);
nand U7136 (N_7136,N_6546,N_6829);
nand U7137 (N_7137,N_6796,N_6840);
nor U7138 (N_7138,N_6771,N_6865);
and U7139 (N_7139,N_6867,N_6539);
xnor U7140 (N_7140,N_6753,N_6603);
nor U7141 (N_7141,N_6584,N_6792);
or U7142 (N_7142,N_6806,N_6599);
nand U7143 (N_7143,N_6721,N_6958);
nor U7144 (N_7144,N_6986,N_6761);
nor U7145 (N_7145,N_6965,N_6910);
and U7146 (N_7146,N_6705,N_6522);
xnor U7147 (N_7147,N_6799,N_6917);
or U7148 (N_7148,N_6569,N_6631);
or U7149 (N_7149,N_6777,N_6868);
or U7150 (N_7150,N_6614,N_6872);
and U7151 (N_7151,N_6524,N_6700);
or U7152 (N_7152,N_6655,N_6932);
xnor U7153 (N_7153,N_6804,N_6795);
nand U7154 (N_7154,N_6999,N_6698);
xor U7155 (N_7155,N_6758,N_6508);
nor U7156 (N_7156,N_6961,N_6835);
nand U7157 (N_7157,N_6767,N_6774);
nand U7158 (N_7158,N_6540,N_6645);
or U7159 (N_7159,N_6926,N_6740);
or U7160 (N_7160,N_6563,N_6678);
nand U7161 (N_7161,N_6518,N_6749);
nor U7162 (N_7162,N_6665,N_6760);
nor U7163 (N_7163,N_6514,N_6783);
xnor U7164 (N_7164,N_6723,N_6892);
or U7165 (N_7165,N_6545,N_6680);
and U7166 (N_7166,N_6937,N_6628);
and U7167 (N_7167,N_6538,N_6891);
nand U7168 (N_7168,N_6561,N_6718);
and U7169 (N_7169,N_6913,N_6701);
nand U7170 (N_7170,N_6939,N_6861);
nor U7171 (N_7171,N_6947,N_6595);
nor U7172 (N_7172,N_6989,N_6811);
nor U7173 (N_7173,N_6604,N_6756);
and U7174 (N_7174,N_6542,N_6503);
and U7175 (N_7175,N_6984,N_6527);
or U7176 (N_7176,N_6898,N_6764);
nand U7177 (N_7177,N_6857,N_6747);
and U7178 (N_7178,N_6513,N_6593);
and U7179 (N_7179,N_6519,N_6589);
nand U7180 (N_7180,N_6936,N_6862);
and U7181 (N_7181,N_6808,N_6899);
nand U7182 (N_7182,N_6613,N_6782);
xnor U7183 (N_7183,N_6640,N_6549);
and U7184 (N_7184,N_6647,N_6914);
xnor U7185 (N_7185,N_6885,N_6556);
xnor U7186 (N_7186,N_6643,N_6954);
nand U7187 (N_7187,N_6726,N_6849);
nand U7188 (N_7188,N_6564,N_6812);
and U7189 (N_7189,N_6734,N_6543);
xnor U7190 (N_7190,N_6709,N_6516);
or U7191 (N_7191,N_6719,N_6703);
or U7192 (N_7192,N_6731,N_6689);
xnor U7193 (N_7193,N_6935,N_6661);
nand U7194 (N_7194,N_6630,N_6744);
nor U7195 (N_7195,N_6547,N_6770);
xnor U7196 (N_7196,N_6553,N_6873);
or U7197 (N_7197,N_6722,N_6966);
nor U7198 (N_7198,N_6597,N_6766);
nand U7199 (N_7199,N_6658,N_6882);
or U7200 (N_7200,N_6938,N_6824);
or U7201 (N_7201,N_6941,N_6692);
or U7202 (N_7202,N_6615,N_6814);
or U7203 (N_7203,N_6669,N_6632);
nand U7204 (N_7204,N_6755,N_6741);
or U7205 (N_7205,N_6666,N_6670);
xnor U7206 (N_7206,N_6888,N_6702);
xnor U7207 (N_7207,N_6572,N_6979);
and U7208 (N_7208,N_6711,N_6900);
or U7209 (N_7209,N_6876,N_6956);
or U7210 (N_7210,N_6541,N_6878);
or U7211 (N_7211,N_6558,N_6780);
xnor U7212 (N_7212,N_6944,N_6951);
or U7213 (N_7213,N_6834,N_6897);
or U7214 (N_7214,N_6605,N_6536);
xor U7215 (N_7215,N_6996,N_6828);
nor U7216 (N_7216,N_6815,N_6978);
and U7217 (N_7217,N_6502,N_6660);
xor U7218 (N_7218,N_6601,N_6642);
nor U7219 (N_7219,N_6933,N_6500);
or U7220 (N_7220,N_6713,N_6510);
and U7221 (N_7221,N_6762,N_6960);
or U7222 (N_7222,N_6602,N_6826);
nand U7223 (N_7223,N_6820,N_6735);
nand U7224 (N_7224,N_6550,N_6779);
nor U7225 (N_7225,N_6644,N_6905);
xor U7226 (N_7226,N_6987,N_6506);
nor U7227 (N_7227,N_6895,N_6769);
xnor U7228 (N_7228,N_6621,N_6813);
nor U7229 (N_7229,N_6889,N_6856);
and U7230 (N_7230,N_6797,N_6983);
nor U7231 (N_7231,N_6855,N_6869);
or U7232 (N_7232,N_6823,N_6962);
and U7233 (N_7233,N_6942,N_6993);
and U7234 (N_7234,N_6946,N_6598);
or U7235 (N_7235,N_6887,N_6567);
xor U7236 (N_7236,N_6772,N_6587);
or U7237 (N_7237,N_6822,N_6827);
or U7238 (N_7238,N_6903,N_6517);
xnor U7239 (N_7239,N_6533,N_6555);
nand U7240 (N_7240,N_6505,N_6560);
nor U7241 (N_7241,N_6596,N_6750);
or U7242 (N_7242,N_6583,N_6668);
nand U7243 (N_7243,N_6998,N_6559);
and U7244 (N_7244,N_6568,N_6990);
nor U7245 (N_7245,N_6816,N_6592);
xor U7246 (N_7246,N_6763,N_6858);
nor U7247 (N_7247,N_6511,N_6594);
or U7248 (N_7248,N_6565,N_6765);
or U7249 (N_7249,N_6611,N_6963);
nor U7250 (N_7250,N_6704,N_6600);
nor U7251 (N_7251,N_6762,N_6995);
or U7252 (N_7252,N_6784,N_6582);
nor U7253 (N_7253,N_6787,N_6569);
nor U7254 (N_7254,N_6650,N_6542);
or U7255 (N_7255,N_6712,N_6904);
and U7256 (N_7256,N_6552,N_6899);
nor U7257 (N_7257,N_6671,N_6881);
xor U7258 (N_7258,N_6678,N_6885);
and U7259 (N_7259,N_6632,N_6807);
and U7260 (N_7260,N_6835,N_6505);
nor U7261 (N_7261,N_6966,N_6820);
or U7262 (N_7262,N_6622,N_6884);
or U7263 (N_7263,N_6823,N_6825);
and U7264 (N_7264,N_6784,N_6600);
nand U7265 (N_7265,N_6665,N_6974);
xnor U7266 (N_7266,N_6664,N_6654);
and U7267 (N_7267,N_6788,N_6822);
xnor U7268 (N_7268,N_6991,N_6509);
nor U7269 (N_7269,N_6731,N_6817);
xor U7270 (N_7270,N_6549,N_6823);
or U7271 (N_7271,N_6827,N_6560);
xor U7272 (N_7272,N_6799,N_6628);
and U7273 (N_7273,N_6584,N_6898);
nand U7274 (N_7274,N_6788,N_6978);
and U7275 (N_7275,N_6596,N_6608);
and U7276 (N_7276,N_6891,N_6999);
or U7277 (N_7277,N_6753,N_6918);
and U7278 (N_7278,N_6771,N_6555);
nor U7279 (N_7279,N_6760,N_6778);
or U7280 (N_7280,N_6550,N_6652);
or U7281 (N_7281,N_6689,N_6665);
nand U7282 (N_7282,N_6742,N_6874);
nor U7283 (N_7283,N_6503,N_6735);
nor U7284 (N_7284,N_6512,N_6575);
nor U7285 (N_7285,N_6918,N_6905);
or U7286 (N_7286,N_6914,N_6569);
or U7287 (N_7287,N_6579,N_6607);
and U7288 (N_7288,N_6878,N_6937);
and U7289 (N_7289,N_6678,N_6719);
nor U7290 (N_7290,N_6696,N_6913);
nor U7291 (N_7291,N_6570,N_6767);
nand U7292 (N_7292,N_6838,N_6622);
or U7293 (N_7293,N_6916,N_6748);
and U7294 (N_7294,N_6530,N_6798);
nand U7295 (N_7295,N_6729,N_6583);
xnor U7296 (N_7296,N_6870,N_6917);
nand U7297 (N_7297,N_6665,N_6751);
and U7298 (N_7298,N_6906,N_6784);
nand U7299 (N_7299,N_6850,N_6882);
nor U7300 (N_7300,N_6642,N_6538);
and U7301 (N_7301,N_6960,N_6763);
or U7302 (N_7302,N_6992,N_6967);
xnor U7303 (N_7303,N_6631,N_6521);
nand U7304 (N_7304,N_6559,N_6754);
xor U7305 (N_7305,N_6631,N_6551);
or U7306 (N_7306,N_6649,N_6983);
nor U7307 (N_7307,N_6791,N_6558);
and U7308 (N_7308,N_6628,N_6741);
nor U7309 (N_7309,N_6950,N_6949);
nor U7310 (N_7310,N_6826,N_6948);
xnor U7311 (N_7311,N_6729,N_6802);
or U7312 (N_7312,N_6700,N_6547);
or U7313 (N_7313,N_6852,N_6556);
or U7314 (N_7314,N_6840,N_6625);
nand U7315 (N_7315,N_6770,N_6751);
xor U7316 (N_7316,N_6679,N_6746);
nand U7317 (N_7317,N_6579,N_6700);
nand U7318 (N_7318,N_6861,N_6579);
or U7319 (N_7319,N_6543,N_6736);
xor U7320 (N_7320,N_6569,N_6882);
nor U7321 (N_7321,N_6908,N_6663);
nand U7322 (N_7322,N_6791,N_6706);
or U7323 (N_7323,N_6882,N_6875);
nor U7324 (N_7324,N_6538,N_6519);
nand U7325 (N_7325,N_6560,N_6644);
or U7326 (N_7326,N_6558,N_6671);
or U7327 (N_7327,N_6838,N_6511);
xor U7328 (N_7328,N_6800,N_6960);
and U7329 (N_7329,N_6958,N_6642);
nand U7330 (N_7330,N_6557,N_6592);
and U7331 (N_7331,N_6973,N_6634);
and U7332 (N_7332,N_6918,N_6954);
or U7333 (N_7333,N_6604,N_6613);
nor U7334 (N_7334,N_6771,N_6793);
nor U7335 (N_7335,N_6559,N_6680);
and U7336 (N_7336,N_6803,N_6748);
nor U7337 (N_7337,N_6515,N_6830);
nor U7338 (N_7338,N_6821,N_6860);
nor U7339 (N_7339,N_6941,N_6785);
nor U7340 (N_7340,N_6597,N_6807);
xnor U7341 (N_7341,N_6808,N_6530);
or U7342 (N_7342,N_6952,N_6817);
nand U7343 (N_7343,N_6590,N_6979);
or U7344 (N_7344,N_6979,N_6635);
and U7345 (N_7345,N_6807,N_6573);
xor U7346 (N_7346,N_6503,N_6971);
and U7347 (N_7347,N_6928,N_6886);
nand U7348 (N_7348,N_6574,N_6626);
nor U7349 (N_7349,N_6625,N_6913);
xor U7350 (N_7350,N_6842,N_6916);
nand U7351 (N_7351,N_6679,N_6503);
xnor U7352 (N_7352,N_6621,N_6914);
xor U7353 (N_7353,N_6821,N_6989);
nor U7354 (N_7354,N_6605,N_6852);
xnor U7355 (N_7355,N_6510,N_6857);
nand U7356 (N_7356,N_6764,N_6696);
nor U7357 (N_7357,N_6943,N_6718);
or U7358 (N_7358,N_6695,N_6767);
or U7359 (N_7359,N_6675,N_6715);
nor U7360 (N_7360,N_6786,N_6581);
nor U7361 (N_7361,N_6607,N_6664);
nor U7362 (N_7362,N_6857,N_6748);
nor U7363 (N_7363,N_6806,N_6690);
or U7364 (N_7364,N_6537,N_6662);
and U7365 (N_7365,N_6623,N_6564);
or U7366 (N_7366,N_6803,N_6569);
xnor U7367 (N_7367,N_6542,N_6915);
nand U7368 (N_7368,N_6708,N_6642);
nor U7369 (N_7369,N_6858,N_6674);
and U7370 (N_7370,N_6568,N_6862);
nor U7371 (N_7371,N_6591,N_6553);
nor U7372 (N_7372,N_6654,N_6793);
or U7373 (N_7373,N_6988,N_6779);
or U7374 (N_7374,N_6850,N_6663);
nor U7375 (N_7375,N_6632,N_6662);
nand U7376 (N_7376,N_6552,N_6979);
nor U7377 (N_7377,N_6551,N_6937);
xor U7378 (N_7378,N_6924,N_6932);
and U7379 (N_7379,N_6660,N_6710);
or U7380 (N_7380,N_6657,N_6559);
xor U7381 (N_7381,N_6694,N_6884);
or U7382 (N_7382,N_6620,N_6684);
and U7383 (N_7383,N_6551,N_6956);
nor U7384 (N_7384,N_6575,N_6729);
or U7385 (N_7385,N_6523,N_6962);
nor U7386 (N_7386,N_6822,N_6730);
or U7387 (N_7387,N_6613,N_6957);
nand U7388 (N_7388,N_6980,N_6507);
and U7389 (N_7389,N_6586,N_6774);
nand U7390 (N_7390,N_6586,N_6840);
or U7391 (N_7391,N_6857,N_6784);
nor U7392 (N_7392,N_6865,N_6947);
or U7393 (N_7393,N_6839,N_6787);
or U7394 (N_7394,N_6998,N_6991);
and U7395 (N_7395,N_6696,N_6924);
nand U7396 (N_7396,N_6574,N_6766);
nand U7397 (N_7397,N_6811,N_6573);
nor U7398 (N_7398,N_6635,N_6950);
and U7399 (N_7399,N_6513,N_6557);
or U7400 (N_7400,N_6974,N_6755);
nor U7401 (N_7401,N_6781,N_6798);
or U7402 (N_7402,N_6715,N_6547);
and U7403 (N_7403,N_6873,N_6716);
or U7404 (N_7404,N_6901,N_6608);
nand U7405 (N_7405,N_6934,N_6787);
xor U7406 (N_7406,N_6551,N_6844);
xnor U7407 (N_7407,N_6589,N_6852);
and U7408 (N_7408,N_6629,N_6869);
or U7409 (N_7409,N_6573,N_6698);
nor U7410 (N_7410,N_6843,N_6625);
or U7411 (N_7411,N_6677,N_6602);
xor U7412 (N_7412,N_6980,N_6918);
and U7413 (N_7413,N_6711,N_6861);
nand U7414 (N_7414,N_6533,N_6833);
nand U7415 (N_7415,N_6589,N_6933);
and U7416 (N_7416,N_6838,N_6797);
and U7417 (N_7417,N_6711,N_6769);
xnor U7418 (N_7418,N_6563,N_6829);
nor U7419 (N_7419,N_6994,N_6795);
or U7420 (N_7420,N_6504,N_6569);
or U7421 (N_7421,N_6533,N_6909);
nor U7422 (N_7422,N_6540,N_6849);
nor U7423 (N_7423,N_6621,N_6939);
xnor U7424 (N_7424,N_6973,N_6652);
or U7425 (N_7425,N_6973,N_6969);
or U7426 (N_7426,N_6710,N_6672);
and U7427 (N_7427,N_6826,N_6892);
nand U7428 (N_7428,N_6618,N_6635);
or U7429 (N_7429,N_6977,N_6596);
or U7430 (N_7430,N_6993,N_6719);
and U7431 (N_7431,N_6613,N_6870);
or U7432 (N_7432,N_6547,N_6690);
or U7433 (N_7433,N_6790,N_6658);
nand U7434 (N_7434,N_6912,N_6911);
xor U7435 (N_7435,N_6969,N_6568);
and U7436 (N_7436,N_6823,N_6837);
nor U7437 (N_7437,N_6986,N_6804);
and U7438 (N_7438,N_6595,N_6720);
xnor U7439 (N_7439,N_6655,N_6884);
nand U7440 (N_7440,N_6968,N_6843);
or U7441 (N_7441,N_6590,N_6778);
xor U7442 (N_7442,N_6781,N_6589);
xnor U7443 (N_7443,N_6708,N_6995);
nor U7444 (N_7444,N_6849,N_6657);
and U7445 (N_7445,N_6755,N_6763);
and U7446 (N_7446,N_6547,N_6718);
and U7447 (N_7447,N_6770,N_6982);
and U7448 (N_7448,N_6871,N_6795);
nor U7449 (N_7449,N_6956,N_6957);
and U7450 (N_7450,N_6831,N_6653);
and U7451 (N_7451,N_6795,N_6649);
nor U7452 (N_7452,N_6608,N_6597);
nor U7453 (N_7453,N_6625,N_6669);
nor U7454 (N_7454,N_6940,N_6660);
or U7455 (N_7455,N_6821,N_6927);
xor U7456 (N_7456,N_6646,N_6679);
nor U7457 (N_7457,N_6649,N_6602);
nor U7458 (N_7458,N_6932,N_6918);
xnor U7459 (N_7459,N_6868,N_6584);
nor U7460 (N_7460,N_6823,N_6784);
and U7461 (N_7461,N_6698,N_6614);
xor U7462 (N_7462,N_6973,N_6713);
nor U7463 (N_7463,N_6692,N_6604);
nand U7464 (N_7464,N_6841,N_6709);
nand U7465 (N_7465,N_6554,N_6770);
and U7466 (N_7466,N_6597,N_6859);
nand U7467 (N_7467,N_6501,N_6608);
and U7468 (N_7468,N_6714,N_6549);
nand U7469 (N_7469,N_6909,N_6891);
nand U7470 (N_7470,N_6509,N_6748);
or U7471 (N_7471,N_6821,N_6611);
nor U7472 (N_7472,N_6620,N_6647);
nand U7473 (N_7473,N_6940,N_6919);
nand U7474 (N_7474,N_6902,N_6670);
nor U7475 (N_7475,N_6863,N_6574);
nor U7476 (N_7476,N_6867,N_6860);
or U7477 (N_7477,N_6523,N_6888);
nor U7478 (N_7478,N_6708,N_6795);
nand U7479 (N_7479,N_6787,N_6700);
xor U7480 (N_7480,N_6647,N_6987);
or U7481 (N_7481,N_6777,N_6575);
nand U7482 (N_7482,N_6509,N_6635);
and U7483 (N_7483,N_6772,N_6932);
nor U7484 (N_7484,N_6790,N_6564);
nand U7485 (N_7485,N_6643,N_6681);
nor U7486 (N_7486,N_6855,N_6725);
xor U7487 (N_7487,N_6969,N_6550);
nand U7488 (N_7488,N_6948,N_6795);
xnor U7489 (N_7489,N_6871,N_6985);
nor U7490 (N_7490,N_6959,N_6552);
and U7491 (N_7491,N_6813,N_6898);
nor U7492 (N_7492,N_6643,N_6720);
nor U7493 (N_7493,N_6769,N_6564);
or U7494 (N_7494,N_6870,N_6988);
and U7495 (N_7495,N_6738,N_6830);
xor U7496 (N_7496,N_6722,N_6822);
or U7497 (N_7497,N_6794,N_6662);
or U7498 (N_7498,N_6837,N_6769);
nor U7499 (N_7499,N_6559,N_6714);
nand U7500 (N_7500,N_7156,N_7114);
and U7501 (N_7501,N_7006,N_7427);
or U7502 (N_7502,N_7194,N_7395);
nor U7503 (N_7503,N_7401,N_7371);
nor U7504 (N_7504,N_7181,N_7319);
nor U7505 (N_7505,N_7465,N_7226);
nor U7506 (N_7506,N_7212,N_7163);
xor U7507 (N_7507,N_7313,N_7169);
xnor U7508 (N_7508,N_7013,N_7357);
xor U7509 (N_7509,N_7483,N_7306);
or U7510 (N_7510,N_7283,N_7148);
xor U7511 (N_7511,N_7215,N_7019);
xor U7512 (N_7512,N_7213,N_7354);
or U7513 (N_7513,N_7278,N_7466);
nor U7514 (N_7514,N_7254,N_7164);
nor U7515 (N_7515,N_7462,N_7280);
xnor U7516 (N_7516,N_7391,N_7286);
nor U7517 (N_7517,N_7311,N_7291);
or U7518 (N_7518,N_7025,N_7364);
xor U7519 (N_7519,N_7358,N_7491);
nand U7520 (N_7520,N_7201,N_7482);
or U7521 (N_7521,N_7033,N_7071);
nor U7522 (N_7522,N_7330,N_7032);
xnor U7523 (N_7523,N_7109,N_7110);
or U7524 (N_7524,N_7302,N_7374);
nor U7525 (N_7525,N_7487,N_7485);
xor U7526 (N_7526,N_7446,N_7091);
nor U7527 (N_7527,N_7328,N_7209);
nand U7528 (N_7528,N_7267,N_7017);
and U7529 (N_7529,N_7259,N_7062);
or U7530 (N_7530,N_7376,N_7162);
or U7531 (N_7531,N_7469,N_7285);
and U7532 (N_7532,N_7179,N_7356);
or U7533 (N_7533,N_7276,N_7447);
xnor U7534 (N_7534,N_7092,N_7347);
nor U7535 (N_7535,N_7230,N_7412);
xor U7536 (N_7536,N_7293,N_7024);
nor U7537 (N_7537,N_7386,N_7012);
nor U7538 (N_7538,N_7288,N_7477);
or U7539 (N_7539,N_7143,N_7296);
nor U7540 (N_7540,N_7431,N_7284);
nand U7541 (N_7541,N_7223,N_7041);
or U7542 (N_7542,N_7224,N_7097);
or U7543 (N_7543,N_7255,N_7074);
and U7544 (N_7544,N_7424,N_7204);
nor U7545 (N_7545,N_7198,N_7021);
nand U7546 (N_7546,N_7337,N_7272);
or U7547 (N_7547,N_7115,N_7359);
xnor U7548 (N_7548,N_7154,N_7035);
nor U7549 (N_7549,N_7027,N_7435);
nor U7550 (N_7550,N_7449,N_7234);
xor U7551 (N_7551,N_7433,N_7461);
nand U7552 (N_7552,N_7152,N_7063);
nand U7553 (N_7553,N_7233,N_7494);
nand U7554 (N_7554,N_7105,N_7060);
or U7555 (N_7555,N_7031,N_7387);
xnor U7556 (N_7556,N_7136,N_7093);
and U7557 (N_7557,N_7274,N_7192);
xnor U7558 (N_7558,N_7208,N_7177);
nand U7559 (N_7559,N_7452,N_7474);
and U7560 (N_7560,N_7235,N_7326);
xnor U7561 (N_7561,N_7398,N_7489);
or U7562 (N_7562,N_7420,N_7004);
xnor U7563 (N_7563,N_7422,N_7150);
nor U7564 (N_7564,N_7367,N_7498);
nand U7565 (N_7565,N_7287,N_7108);
nor U7566 (N_7566,N_7053,N_7340);
nand U7567 (N_7567,N_7432,N_7368);
xnor U7568 (N_7568,N_7122,N_7200);
nand U7569 (N_7569,N_7083,N_7244);
nor U7570 (N_7570,N_7327,N_7382);
xnor U7571 (N_7571,N_7210,N_7300);
or U7572 (N_7572,N_7101,N_7082);
nor U7573 (N_7573,N_7098,N_7409);
or U7574 (N_7574,N_7059,N_7172);
nand U7575 (N_7575,N_7301,N_7043);
or U7576 (N_7576,N_7282,N_7068);
xnor U7577 (N_7577,N_7185,N_7430);
or U7578 (N_7578,N_7318,N_7001);
xor U7579 (N_7579,N_7086,N_7463);
or U7580 (N_7580,N_7457,N_7436);
nor U7581 (N_7581,N_7023,N_7178);
and U7582 (N_7582,N_7094,N_7471);
xnor U7583 (N_7583,N_7137,N_7403);
xnor U7584 (N_7584,N_7155,N_7250);
xor U7585 (N_7585,N_7247,N_7348);
or U7586 (N_7586,N_7478,N_7252);
xnor U7587 (N_7587,N_7362,N_7381);
and U7588 (N_7588,N_7481,N_7183);
or U7589 (N_7589,N_7049,N_7052);
nor U7590 (N_7590,N_7444,N_7046);
or U7591 (N_7591,N_7044,N_7125);
xnor U7592 (N_7592,N_7089,N_7281);
xor U7593 (N_7593,N_7321,N_7197);
nand U7594 (N_7594,N_7051,N_7170);
and U7595 (N_7595,N_7232,N_7499);
nand U7596 (N_7596,N_7355,N_7275);
or U7597 (N_7597,N_7324,N_7456);
and U7598 (N_7598,N_7190,N_7270);
xnor U7599 (N_7599,N_7417,N_7138);
nand U7600 (N_7600,N_7440,N_7495);
xor U7601 (N_7601,N_7222,N_7058);
or U7602 (N_7602,N_7455,N_7249);
and U7603 (N_7603,N_7383,N_7385);
nor U7604 (N_7604,N_7407,N_7390);
xnor U7605 (N_7605,N_7087,N_7026);
or U7606 (N_7606,N_7076,N_7206);
nand U7607 (N_7607,N_7425,N_7126);
xnor U7608 (N_7608,N_7048,N_7149);
nand U7609 (N_7609,N_7221,N_7472);
or U7610 (N_7610,N_7139,N_7072);
or U7611 (N_7611,N_7069,N_7040);
nor U7612 (N_7612,N_7199,N_7442);
nand U7613 (N_7613,N_7344,N_7323);
nand U7614 (N_7614,N_7251,N_7184);
and U7615 (N_7615,N_7257,N_7265);
or U7616 (N_7616,N_7158,N_7405);
nand U7617 (N_7617,N_7140,N_7145);
nand U7618 (N_7618,N_7207,N_7258);
nor U7619 (N_7619,N_7341,N_7002);
nand U7620 (N_7620,N_7345,N_7490);
xor U7621 (N_7621,N_7171,N_7146);
xnor U7622 (N_7622,N_7339,N_7279);
or U7623 (N_7623,N_7396,N_7066);
or U7624 (N_7624,N_7182,N_7470);
and U7625 (N_7625,N_7392,N_7174);
or U7626 (N_7626,N_7262,N_7413);
xnor U7627 (N_7627,N_7034,N_7402);
nor U7628 (N_7628,N_7127,N_7246);
nor U7629 (N_7629,N_7315,N_7373);
nand U7630 (N_7630,N_7193,N_7473);
or U7631 (N_7631,N_7384,N_7073);
xnor U7632 (N_7632,N_7191,N_7428);
xor U7633 (N_7633,N_7151,N_7099);
or U7634 (N_7634,N_7240,N_7410);
xor U7635 (N_7635,N_7061,N_7353);
nor U7636 (N_7636,N_7176,N_7277);
xnor U7637 (N_7637,N_7379,N_7266);
xnor U7638 (N_7638,N_7070,N_7103);
and U7639 (N_7639,N_7480,N_7123);
nand U7640 (N_7640,N_7468,N_7458);
and U7641 (N_7641,N_7443,N_7366);
nand U7642 (N_7642,N_7010,N_7329);
and U7643 (N_7643,N_7426,N_7116);
nand U7644 (N_7644,N_7029,N_7370);
nor U7645 (N_7645,N_7256,N_7352);
nor U7646 (N_7646,N_7335,N_7312);
nand U7647 (N_7647,N_7134,N_7187);
nor U7648 (N_7648,N_7018,N_7451);
nor U7649 (N_7649,N_7338,N_7022);
nor U7650 (N_7650,N_7441,N_7346);
and U7651 (N_7651,N_7118,N_7408);
nor U7652 (N_7652,N_7037,N_7106);
and U7653 (N_7653,N_7448,N_7445);
nand U7654 (N_7654,N_7237,N_7055);
or U7655 (N_7655,N_7078,N_7394);
and U7656 (N_7656,N_7450,N_7294);
and U7657 (N_7657,N_7225,N_7493);
nand U7658 (N_7658,N_7389,N_7400);
and U7659 (N_7659,N_7363,N_7241);
nor U7660 (N_7660,N_7057,N_7459);
or U7661 (N_7661,N_7476,N_7121);
nand U7662 (N_7662,N_7167,N_7434);
nor U7663 (N_7663,N_7332,N_7333);
nor U7664 (N_7664,N_7304,N_7414);
or U7665 (N_7665,N_7119,N_7297);
xnor U7666 (N_7666,N_7292,N_7261);
nor U7667 (N_7667,N_7111,N_7438);
nand U7668 (N_7668,N_7336,N_7080);
nand U7669 (N_7669,N_7299,N_7310);
nor U7670 (N_7670,N_7406,N_7128);
nor U7671 (N_7671,N_7075,N_7227);
xor U7672 (N_7672,N_7175,N_7000);
xnor U7673 (N_7673,N_7039,N_7065);
or U7674 (N_7674,N_7289,N_7100);
xor U7675 (N_7675,N_7016,N_7273);
nand U7676 (N_7676,N_7011,N_7211);
nand U7677 (N_7677,N_7248,N_7325);
nor U7678 (N_7678,N_7160,N_7264);
nor U7679 (N_7679,N_7236,N_7369);
or U7680 (N_7680,N_7014,N_7064);
nor U7681 (N_7681,N_7050,N_7195);
or U7682 (N_7682,N_7090,N_7467);
nor U7683 (N_7683,N_7005,N_7129);
or U7684 (N_7684,N_7186,N_7404);
nand U7685 (N_7685,N_7030,N_7334);
or U7686 (N_7686,N_7102,N_7077);
xnor U7687 (N_7687,N_7497,N_7484);
nor U7688 (N_7688,N_7377,N_7421);
nand U7689 (N_7689,N_7454,N_7263);
nor U7690 (N_7690,N_7268,N_7439);
and U7691 (N_7691,N_7088,N_7219);
and U7692 (N_7692,N_7416,N_7375);
and U7693 (N_7693,N_7141,N_7214);
xnor U7694 (N_7694,N_7113,N_7218);
xor U7695 (N_7695,N_7216,N_7492);
nor U7696 (N_7696,N_7488,N_7168);
and U7697 (N_7697,N_7243,N_7202);
xor U7698 (N_7698,N_7153,N_7423);
xor U7699 (N_7699,N_7008,N_7120);
nor U7700 (N_7700,N_7229,N_7189);
or U7701 (N_7701,N_7343,N_7161);
xor U7702 (N_7702,N_7144,N_7173);
nand U7703 (N_7703,N_7453,N_7196);
and U7704 (N_7704,N_7429,N_7308);
or U7705 (N_7705,N_7361,N_7349);
nand U7706 (N_7706,N_7331,N_7054);
nand U7707 (N_7707,N_7003,N_7295);
nand U7708 (N_7708,N_7085,N_7096);
nand U7709 (N_7709,N_7350,N_7378);
nand U7710 (N_7710,N_7038,N_7132);
nand U7711 (N_7711,N_7042,N_7271);
nand U7712 (N_7712,N_7496,N_7290);
and U7713 (N_7713,N_7317,N_7117);
and U7714 (N_7714,N_7351,N_7245);
nor U7715 (N_7715,N_7260,N_7081);
nand U7716 (N_7716,N_7231,N_7124);
or U7717 (N_7717,N_7079,N_7415);
or U7718 (N_7718,N_7166,N_7388);
nand U7719 (N_7719,N_7112,N_7217);
nand U7720 (N_7720,N_7220,N_7411);
and U7721 (N_7721,N_7056,N_7320);
or U7722 (N_7722,N_7399,N_7307);
xnor U7723 (N_7723,N_7130,N_7159);
nor U7724 (N_7724,N_7418,N_7437);
nor U7725 (N_7725,N_7203,N_7007);
nand U7726 (N_7726,N_7460,N_7479);
xnor U7727 (N_7727,N_7135,N_7045);
nor U7728 (N_7728,N_7147,N_7393);
xnor U7729 (N_7729,N_7380,N_7165);
and U7730 (N_7730,N_7372,N_7239);
or U7731 (N_7731,N_7342,N_7309);
nand U7732 (N_7732,N_7228,N_7020);
or U7733 (N_7733,N_7095,N_7142);
nand U7734 (N_7734,N_7419,N_7133);
nor U7735 (N_7735,N_7131,N_7067);
and U7736 (N_7736,N_7475,N_7242);
nor U7737 (N_7737,N_7015,N_7009);
or U7738 (N_7738,N_7036,N_7269);
and U7739 (N_7739,N_7084,N_7298);
nand U7740 (N_7740,N_7322,N_7305);
nand U7741 (N_7741,N_7028,N_7303);
or U7742 (N_7742,N_7464,N_7180);
nor U7743 (N_7743,N_7486,N_7360);
or U7744 (N_7744,N_7365,N_7397);
and U7745 (N_7745,N_7107,N_7188);
and U7746 (N_7746,N_7253,N_7205);
xnor U7747 (N_7747,N_7314,N_7104);
xnor U7748 (N_7748,N_7238,N_7047);
nand U7749 (N_7749,N_7157,N_7316);
nor U7750 (N_7750,N_7411,N_7030);
xnor U7751 (N_7751,N_7371,N_7404);
and U7752 (N_7752,N_7209,N_7310);
and U7753 (N_7753,N_7492,N_7453);
xor U7754 (N_7754,N_7264,N_7204);
nor U7755 (N_7755,N_7432,N_7145);
or U7756 (N_7756,N_7426,N_7468);
and U7757 (N_7757,N_7139,N_7090);
xor U7758 (N_7758,N_7447,N_7073);
nand U7759 (N_7759,N_7325,N_7453);
and U7760 (N_7760,N_7107,N_7000);
xor U7761 (N_7761,N_7009,N_7064);
nor U7762 (N_7762,N_7302,N_7245);
xor U7763 (N_7763,N_7321,N_7487);
and U7764 (N_7764,N_7137,N_7383);
and U7765 (N_7765,N_7058,N_7072);
xnor U7766 (N_7766,N_7381,N_7250);
nand U7767 (N_7767,N_7478,N_7475);
xnor U7768 (N_7768,N_7329,N_7394);
or U7769 (N_7769,N_7130,N_7156);
or U7770 (N_7770,N_7413,N_7457);
xor U7771 (N_7771,N_7178,N_7036);
nor U7772 (N_7772,N_7010,N_7438);
nor U7773 (N_7773,N_7208,N_7414);
nand U7774 (N_7774,N_7440,N_7403);
nand U7775 (N_7775,N_7454,N_7393);
nor U7776 (N_7776,N_7256,N_7086);
xor U7777 (N_7777,N_7486,N_7226);
xor U7778 (N_7778,N_7402,N_7371);
or U7779 (N_7779,N_7190,N_7492);
nand U7780 (N_7780,N_7206,N_7378);
and U7781 (N_7781,N_7486,N_7016);
xor U7782 (N_7782,N_7034,N_7003);
or U7783 (N_7783,N_7122,N_7013);
xnor U7784 (N_7784,N_7455,N_7108);
nor U7785 (N_7785,N_7485,N_7343);
xnor U7786 (N_7786,N_7265,N_7132);
or U7787 (N_7787,N_7412,N_7339);
nand U7788 (N_7788,N_7209,N_7093);
xnor U7789 (N_7789,N_7035,N_7463);
xnor U7790 (N_7790,N_7169,N_7314);
nand U7791 (N_7791,N_7348,N_7011);
or U7792 (N_7792,N_7181,N_7009);
and U7793 (N_7793,N_7458,N_7325);
nor U7794 (N_7794,N_7195,N_7456);
or U7795 (N_7795,N_7256,N_7390);
or U7796 (N_7796,N_7396,N_7380);
or U7797 (N_7797,N_7303,N_7329);
xnor U7798 (N_7798,N_7017,N_7019);
xor U7799 (N_7799,N_7332,N_7329);
nor U7800 (N_7800,N_7340,N_7139);
nand U7801 (N_7801,N_7440,N_7448);
nor U7802 (N_7802,N_7403,N_7165);
or U7803 (N_7803,N_7169,N_7321);
nand U7804 (N_7804,N_7192,N_7293);
xnor U7805 (N_7805,N_7268,N_7326);
nor U7806 (N_7806,N_7018,N_7221);
xnor U7807 (N_7807,N_7459,N_7205);
xnor U7808 (N_7808,N_7453,N_7386);
xnor U7809 (N_7809,N_7084,N_7401);
nand U7810 (N_7810,N_7197,N_7057);
nand U7811 (N_7811,N_7119,N_7337);
xnor U7812 (N_7812,N_7082,N_7340);
and U7813 (N_7813,N_7276,N_7399);
xnor U7814 (N_7814,N_7321,N_7216);
nand U7815 (N_7815,N_7323,N_7413);
or U7816 (N_7816,N_7205,N_7241);
or U7817 (N_7817,N_7430,N_7326);
nand U7818 (N_7818,N_7141,N_7139);
and U7819 (N_7819,N_7250,N_7098);
and U7820 (N_7820,N_7435,N_7148);
nand U7821 (N_7821,N_7306,N_7274);
or U7822 (N_7822,N_7018,N_7010);
or U7823 (N_7823,N_7011,N_7131);
nand U7824 (N_7824,N_7160,N_7448);
or U7825 (N_7825,N_7256,N_7446);
or U7826 (N_7826,N_7406,N_7284);
xnor U7827 (N_7827,N_7074,N_7098);
xnor U7828 (N_7828,N_7351,N_7335);
nand U7829 (N_7829,N_7337,N_7088);
xnor U7830 (N_7830,N_7347,N_7181);
and U7831 (N_7831,N_7435,N_7220);
xnor U7832 (N_7832,N_7450,N_7424);
or U7833 (N_7833,N_7109,N_7064);
nand U7834 (N_7834,N_7385,N_7132);
xor U7835 (N_7835,N_7118,N_7199);
xor U7836 (N_7836,N_7384,N_7350);
xnor U7837 (N_7837,N_7270,N_7344);
or U7838 (N_7838,N_7128,N_7287);
nor U7839 (N_7839,N_7056,N_7289);
xnor U7840 (N_7840,N_7189,N_7221);
nand U7841 (N_7841,N_7337,N_7370);
xor U7842 (N_7842,N_7270,N_7377);
or U7843 (N_7843,N_7199,N_7222);
nand U7844 (N_7844,N_7315,N_7148);
xnor U7845 (N_7845,N_7432,N_7398);
and U7846 (N_7846,N_7170,N_7284);
or U7847 (N_7847,N_7340,N_7032);
nand U7848 (N_7848,N_7298,N_7375);
or U7849 (N_7849,N_7359,N_7286);
or U7850 (N_7850,N_7394,N_7447);
or U7851 (N_7851,N_7160,N_7099);
nor U7852 (N_7852,N_7079,N_7110);
or U7853 (N_7853,N_7483,N_7213);
and U7854 (N_7854,N_7243,N_7463);
xor U7855 (N_7855,N_7086,N_7483);
xnor U7856 (N_7856,N_7115,N_7456);
nor U7857 (N_7857,N_7467,N_7204);
nor U7858 (N_7858,N_7470,N_7105);
or U7859 (N_7859,N_7244,N_7342);
or U7860 (N_7860,N_7203,N_7128);
nand U7861 (N_7861,N_7145,N_7350);
nand U7862 (N_7862,N_7058,N_7206);
xor U7863 (N_7863,N_7076,N_7148);
and U7864 (N_7864,N_7113,N_7258);
or U7865 (N_7865,N_7184,N_7289);
xor U7866 (N_7866,N_7198,N_7207);
nand U7867 (N_7867,N_7265,N_7380);
xnor U7868 (N_7868,N_7357,N_7258);
nor U7869 (N_7869,N_7037,N_7088);
xnor U7870 (N_7870,N_7303,N_7389);
nor U7871 (N_7871,N_7032,N_7274);
nand U7872 (N_7872,N_7488,N_7359);
nor U7873 (N_7873,N_7009,N_7437);
or U7874 (N_7874,N_7297,N_7378);
nor U7875 (N_7875,N_7277,N_7448);
xor U7876 (N_7876,N_7142,N_7257);
nor U7877 (N_7877,N_7447,N_7370);
nor U7878 (N_7878,N_7220,N_7061);
or U7879 (N_7879,N_7309,N_7453);
xnor U7880 (N_7880,N_7171,N_7075);
nand U7881 (N_7881,N_7149,N_7329);
and U7882 (N_7882,N_7282,N_7121);
and U7883 (N_7883,N_7214,N_7398);
and U7884 (N_7884,N_7436,N_7021);
xor U7885 (N_7885,N_7103,N_7492);
or U7886 (N_7886,N_7372,N_7131);
nand U7887 (N_7887,N_7220,N_7097);
or U7888 (N_7888,N_7257,N_7333);
xor U7889 (N_7889,N_7273,N_7321);
nor U7890 (N_7890,N_7477,N_7321);
xnor U7891 (N_7891,N_7079,N_7314);
xnor U7892 (N_7892,N_7076,N_7249);
or U7893 (N_7893,N_7381,N_7490);
nand U7894 (N_7894,N_7302,N_7434);
nor U7895 (N_7895,N_7121,N_7410);
or U7896 (N_7896,N_7061,N_7293);
or U7897 (N_7897,N_7038,N_7170);
xor U7898 (N_7898,N_7061,N_7253);
and U7899 (N_7899,N_7074,N_7436);
nand U7900 (N_7900,N_7209,N_7327);
nor U7901 (N_7901,N_7034,N_7302);
nor U7902 (N_7902,N_7426,N_7361);
nor U7903 (N_7903,N_7296,N_7428);
and U7904 (N_7904,N_7015,N_7178);
xor U7905 (N_7905,N_7130,N_7315);
nor U7906 (N_7906,N_7209,N_7346);
xor U7907 (N_7907,N_7267,N_7245);
nand U7908 (N_7908,N_7105,N_7025);
nor U7909 (N_7909,N_7152,N_7470);
nand U7910 (N_7910,N_7417,N_7079);
nor U7911 (N_7911,N_7210,N_7303);
xor U7912 (N_7912,N_7179,N_7013);
nor U7913 (N_7913,N_7089,N_7040);
or U7914 (N_7914,N_7057,N_7442);
xnor U7915 (N_7915,N_7093,N_7222);
nor U7916 (N_7916,N_7461,N_7114);
xnor U7917 (N_7917,N_7176,N_7114);
nor U7918 (N_7918,N_7179,N_7150);
xnor U7919 (N_7919,N_7193,N_7143);
xnor U7920 (N_7920,N_7252,N_7146);
and U7921 (N_7921,N_7310,N_7219);
xnor U7922 (N_7922,N_7280,N_7382);
and U7923 (N_7923,N_7297,N_7105);
nor U7924 (N_7924,N_7195,N_7447);
nand U7925 (N_7925,N_7141,N_7443);
xor U7926 (N_7926,N_7095,N_7060);
nor U7927 (N_7927,N_7419,N_7486);
nand U7928 (N_7928,N_7207,N_7162);
and U7929 (N_7929,N_7194,N_7336);
xor U7930 (N_7930,N_7119,N_7394);
nor U7931 (N_7931,N_7482,N_7002);
xor U7932 (N_7932,N_7041,N_7263);
and U7933 (N_7933,N_7024,N_7048);
and U7934 (N_7934,N_7055,N_7340);
xnor U7935 (N_7935,N_7301,N_7482);
nand U7936 (N_7936,N_7001,N_7380);
nor U7937 (N_7937,N_7134,N_7286);
xor U7938 (N_7938,N_7029,N_7030);
xnor U7939 (N_7939,N_7048,N_7147);
nor U7940 (N_7940,N_7140,N_7217);
nor U7941 (N_7941,N_7259,N_7261);
nor U7942 (N_7942,N_7074,N_7073);
nor U7943 (N_7943,N_7442,N_7100);
nor U7944 (N_7944,N_7229,N_7253);
and U7945 (N_7945,N_7448,N_7326);
or U7946 (N_7946,N_7489,N_7292);
or U7947 (N_7947,N_7264,N_7024);
nand U7948 (N_7948,N_7420,N_7125);
nor U7949 (N_7949,N_7234,N_7043);
nand U7950 (N_7950,N_7484,N_7213);
nand U7951 (N_7951,N_7105,N_7370);
or U7952 (N_7952,N_7342,N_7364);
xnor U7953 (N_7953,N_7482,N_7449);
nand U7954 (N_7954,N_7286,N_7305);
and U7955 (N_7955,N_7497,N_7018);
xnor U7956 (N_7956,N_7311,N_7160);
or U7957 (N_7957,N_7087,N_7357);
nor U7958 (N_7958,N_7390,N_7284);
and U7959 (N_7959,N_7380,N_7291);
and U7960 (N_7960,N_7350,N_7371);
xor U7961 (N_7961,N_7332,N_7108);
nand U7962 (N_7962,N_7240,N_7271);
and U7963 (N_7963,N_7495,N_7368);
nor U7964 (N_7964,N_7285,N_7085);
nand U7965 (N_7965,N_7429,N_7059);
and U7966 (N_7966,N_7049,N_7082);
nand U7967 (N_7967,N_7231,N_7230);
nand U7968 (N_7968,N_7478,N_7201);
and U7969 (N_7969,N_7203,N_7255);
or U7970 (N_7970,N_7213,N_7318);
nand U7971 (N_7971,N_7011,N_7017);
and U7972 (N_7972,N_7457,N_7452);
nor U7973 (N_7973,N_7063,N_7498);
nand U7974 (N_7974,N_7285,N_7490);
or U7975 (N_7975,N_7223,N_7428);
nor U7976 (N_7976,N_7198,N_7417);
xnor U7977 (N_7977,N_7078,N_7361);
nor U7978 (N_7978,N_7119,N_7253);
nand U7979 (N_7979,N_7233,N_7084);
or U7980 (N_7980,N_7352,N_7210);
nand U7981 (N_7981,N_7118,N_7112);
or U7982 (N_7982,N_7267,N_7094);
and U7983 (N_7983,N_7371,N_7170);
nor U7984 (N_7984,N_7224,N_7460);
or U7985 (N_7985,N_7289,N_7387);
nand U7986 (N_7986,N_7452,N_7169);
nor U7987 (N_7987,N_7410,N_7236);
nor U7988 (N_7988,N_7042,N_7101);
xor U7989 (N_7989,N_7389,N_7101);
or U7990 (N_7990,N_7057,N_7133);
nand U7991 (N_7991,N_7359,N_7164);
nand U7992 (N_7992,N_7404,N_7051);
nor U7993 (N_7993,N_7489,N_7272);
or U7994 (N_7994,N_7271,N_7006);
or U7995 (N_7995,N_7117,N_7218);
xnor U7996 (N_7996,N_7351,N_7276);
xnor U7997 (N_7997,N_7235,N_7159);
xnor U7998 (N_7998,N_7423,N_7264);
or U7999 (N_7999,N_7400,N_7242);
and U8000 (N_8000,N_7884,N_7674);
nor U8001 (N_8001,N_7999,N_7617);
nand U8002 (N_8002,N_7577,N_7893);
and U8003 (N_8003,N_7722,N_7525);
and U8004 (N_8004,N_7826,N_7548);
xnor U8005 (N_8005,N_7558,N_7915);
xnor U8006 (N_8006,N_7518,N_7941);
nand U8007 (N_8007,N_7638,N_7951);
or U8008 (N_8008,N_7543,N_7760);
and U8009 (N_8009,N_7631,N_7624);
nor U8010 (N_8010,N_7758,N_7730);
and U8011 (N_8011,N_7653,N_7850);
and U8012 (N_8012,N_7594,N_7662);
or U8013 (N_8013,N_7928,N_7569);
xor U8014 (N_8014,N_7926,N_7879);
nor U8015 (N_8015,N_7847,N_7554);
xor U8016 (N_8016,N_7901,N_7959);
xor U8017 (N_8017,N_7509,N_7922);
or U8018 (N_8018,N_7817,N_7632);
nor U8019 (N_8019,N_7687,N_7640);
and U8020 (N_8020,N_7995,N_7774);
or U8021 (N_8021,N_7610,N_7769);
xnor U8022 (N_8022,N_7627,N_7968);
nor U8023 (N_8023,N_7710,N_7652);
nand U8024 (N_8024,N_7547,N_7564);
xnor U8025 (N_8025,N_7675,N_7742);
and U8026 (N_8026,N_7511,N_7764);
or U8027 (N_8027,N_7700,N_7500);
nand U8028 (N_8028,N_7855,N_7816);
nor U8029 (N_8029,N_7669,N_7861);
and U8030 (N_8030,N_7852,N_7780);
or U8031 (N_8031,N_7940,N_7596);
or U8032 (N_8032,N_7524,N_7683);
xor U8033 (N_8033,N_7967,N_7641);
nor U8034 (N_8034,N_7949,N_7909);
nand U8035 (N_8035,N_7567,N_7581);
or U8036 (N_8036,N_7705,N_7923);
or U8037 (N_8037,N_7727,N_7728);
nand U8038 (N_8038,N_7680,N_7813);
nand U8039 (N_8039,N_7930,N_7910);
and U8040 (N_8040,N_7835,N_7782);
and U8041 (N_8041,N_7794,N_7693);
and U8042 (N_8042,N_7553,N_7920);
and U8043 (N_8043,N_7744,N_7749);
and U8044 (N_8044,N_7888,N_7745);
or U8045 (N_8045,N_7906,N_7833);
nand U8046 (N_8046,N_7766,N_7536);
nand U8047 (N_8047,N_7899,N_7838);
nor U8048 (N_8048,N_7917,N_7682);
nand U8049 (N_8049,N_7840,N_7649);
and U8050 (N_8050,N_7592,N_7831);
or U8051 (N_8051,N_7880,N_7666);
and U8052 (N_8052,N_7613,N_7796);
and U8053 (N_8053,N_7903,N_7507);
or U8054 (N_8054,N_7797,N_7656);
xor U8055 (N_8055,N_7714,N_7534);
nor U8056 (N_8056,N_7799,N_7828);
nand U8057 (N_8057,N_7668,N_7887);
nor U8058 (N_8058,N_7998,N_7751);
nand U8059 (N_8059,N_7528,N_7827);
and U8060 (N_8060,N_7695,N_7869);
or U8061 (N_8061,N_7535,N_7609);
nand U8062 (N_8062,N_7542,N_7932);
or U8063 (N_8063,N_7529,N_7538);
nor U8064 (N_8064,N_7900,N_7818);
or U8065 (N_8065,N_7800,N_7913);
nand U8066 (N_8066,N_7723,N_7713);
nor U8067 (N_8067,N_7561,N_7974);
nor U8068 (N_8068,N_7508,N_7986);
and U8069 (N_8069,N_7946,N_7767);
or U8070 (N_8070,N_7905,N_7757);
and U8071 (N_8071,N_7512,N_7788);
xor U8072 (N_8072,N_7801,N_7778);
and U8073 (N_8073,N_7977,N_7619);
and U8074 (N_8074,N_7697,N_7886);
xnor U8075 (N_8075,N_7731,N_7587);
xor U8076 (N_8076,N_7600,N_7639);
or U8077 (N_8077,N_7980,N_7732);
nor U8078 (N_8078,N_7936,N_7964);
and U8079 (N_8079,N_7925,N_7625);
nand U8080 (N_8080,N_7615,N_7911);
xor U8081 (N_8081,N_7702,N_7939);
xnor U8082 (N_8082,N_7614,N_7891);
and U8083 (N_8083,N_7636,N_7725);
and U8084 (N_8084,N_7907,N_7779);
nor U8085 (N_8085,N_7866,N_7657);
xor U8086 (N_8086,N_7621,N_7804);
and U8087 (N_8087,N_7792,N_7551);
nor U8088 (N_8088,N_7950,N_7918);
nor U8089 (N_8089,N_7517,N_7622);
and U8090 (N_8090,N_7692,N_7606);
and U8091 (N_8091,N_7985,N_7570);
and U8092 (N_8092,N_7785,N_7962);
nor U8093 (N_8093,N_7608,N_7793);
and U8094 (N_8094,N_7618,N_7571);
or U8095 (N_8095,N_7862,N_7844);
nor U8096 (N_8096,N_7821,N_7783);
nand U8097 (N_8097,N_7952,N_7841);
and U8098 (N_8098,N_7895,N_7765);
xnor U8099 (N_8099,N_7521,N_7832);
nand U8100 (N_8100,N_7597,N_7948);
and U8101 (N_8101,N_7768,N_7672);
nand U8102 (N_8102,N_7503,N_7527);
and U8103 (N_8103,N_7890,N_7882);
and U8104 (N_8104,N_7556,N_7753);
xor U8105 (N_8105,N_7676,N_7784);
or U8106 (N_8106,N_7781,N_7699);
nand U8107 (N_8107,N_7659,N_7563);
or U8108 (N_8108,N_7791,N_7960);
and U8109 (N_8109,N_7634,N_7715);
and U8110 (N_8110,N_7726,N_7670);
xor U8111 (N_8111,N_7679,N_7754);
xor U8112 (N_8112,N_7963,N_7604);
nor U8113 (N_8113,N_7759,N_7510);
xnor U8114 (N_8114,N_7858,N_7593);
nor U8115 (N_8115,N_7501,N_7867);
nor U8116 (N_8116,N_7642,N_7979);
xnor U8117 (N_8117,N_7790,N_7537);
and U8118 (N_8118,N_7989,N_7802);
and U8119 (N_8119,N_7736,N_7557);
nor U8120 (N_8120,N_7568,N_7660);
and U8121 (N_8121,N_7513,N_7506);
or U8122 (N_8122,N_7856,N_7973);
and U8123 (N_8123,N_7544,N_7969);
and U8124 (N_8124,N_7738,N_7647);
xnor U8125 (N_8125,N_7805,N_7750);
nand U8126 (N_8126,N_7756,N_7830);
xnor U8127 (N_8127,N_7583,N_7868);
or U8128 (N_8128,N_7916,N_7643);
xor U8129 (N_8129,N_7740,N_7580);
nand U8130 (N_8130,N_7601,N_7530);
nand U8131 (N_8131,N_7650,N_7752);
nor U8132 (N_8132,N_7771,N_7540);
nor U8133 (N_8133,N_7881,N_7770);
or U8134 (N_8134,N_7681,N_7651);
xnor U8135 (N_8135,N_7665,N_7896);
nor U8136 (N_8136,N_7739,N_7822);
xnor U8137 (N_8137,N_7935,N_7874);
xnor U8138 (N_8138,N_7629,N_7573);
and U8139 (N_8139,N_7644,N_7843);
and U8140 (N_8140,N_7684,N_7845);
and U8141 (N_8141,N_7971,N_7914);
or U8142 (N_8142,N_7599,N_7836);
and U8143 (N_8143,N_7904,N_7648);
xor U8144 (N_8144,N_7626,N_7533);
nor U8145 (N_8145,N_7719,N_7942);
and U8146 (N_8146,N_7630,N_7953);
or U8147 (N_8147,N_7958,N_7814);
and U8148 (N_8148,N_7696,N_7834);
xnor U8149 (N_8149,N_7663,N_7761);
and U8150 (N_8150,N_7546,N_7853);
or U8151 (N_8151,N_7851,N_7701);
xor U8152 (N_8152,N_7504,N_7612);
nand U8153 (N_8153,N_7772,N_7937);
nor U8154 (N_8154,N_7691,N_7798);
nand U8155 (N_8155,N_7755,N_7854);
nor U8156 (N_8156,N_7545,N_7823);
and U8157 (N_8157,N_7611,N_7902);
and U8158 (N_8158,N_7934,N_7775);
and U8159 (N_8159,N_7820,N_7897);
nor U8160 (N_8160,N_7743,N_7961);
xnor U8161 (N_8161,N_7966,N_7720);
nand U8162 (N_8162,N_7812,N_7735);
or U8163 (N_8163,N_7531,N_7724);
and U8164 (N_8164,N_7921,N_7709);
and U8165 (N_8165,N_7839,N_7562);
xor U8166 (N_8166,N_7992,N_7819);
and U8167 (N_8167,N_7747,N_7846);
or U8168 (N_8168,N_7655,N_7717);
nand U8169 (N_8169,N_7671,N_7689);
xor U8170 (N_8170,N_7585,N_7582);
xor U8171 (N_8171,N_7678,N_7707);
and U8172 (N_8172,N_7924,N_7633);
nand U8173 (N_8173,N_7628,N_7541);
nand U8174 (N_8174,N_7677,N_7807);
and U8175 (N_8175,N_7616,N_7523);
and U8176 (N_8176,N_7876,N_7894);
or U8177 (N_8177,N_7877,N_7944);
and U8178 (N_8178,N_7620,N_7815);
xor U8179 (N_8179,N_7803,N_7708);
xor U8180 (N_8180,N_7912,N_7889);
and U8181 (N_8181,N_7806,N_7982);
or U8182 (N_8182,N_7983,N_7996);
nand U8183 (N_8183,N_7860,N_7810);
and U8184 (N_8184,N_7970,N_7703);
xor U8185 (N_8185,N_7829,N_7865);
nor U8186 (N_8186,N_7842,N_7824);
nand U8187 (N_8187,N_7808,N_7965);
nor U8188 (N_8188,N_7635,N_7947);
or U8189 (N_8189,N_7704,N_7908);
or U8190 (N_8190,N_7623,N_7502);
nor U8191 (N_8191,N_7892,N_7872);
xnor U8192 (N_8192,N_7938,N_7565);
nor U8193 (N_8193,N_7737,N_7591);
and U8194 (N_8194,N_7933,N_7955);
nand U8195 (N_8195,N_7721,N_7733);
and U8196 (N_8196,N_7848,N_7688);
nand U8197 (N_8197,N_7787,N_7987);
or U8198 (N_8198,N_7519,N_7574);
and U8199 (N_8199,N_7646,N_7870);
nor U8200 (N_8200,N_7716,N_7931);
and U8201 (N_8201,N_7898,N_7712);
nor U8202 (N_8202,N_7686,N_7514);
nor U8203 (N_8203,N_7589,N_7539);
or U8204 (N_8204,N_7584,N_7595);
and U8205 (N_8205,N_7729,N_7990);
or U8206 (N_8206,N_7929,N_7871);
xor U8207 (N_8207,N_7776,N_7972);
nor U8208 (N_8208,N_7988,N_7505);
or U8209 (N_8209,N_7811,N_7711);
or U8210 (N_8210,N_7825,N_7706);
and U8211 (N_8211,N_7746,N_7549);
nor U8212 (N_8212,N_7976,N_7605);
and U8213 (N_8213,N_7637,N_7809);
and U8214 (N_8214,N_7863,N_7919);
or U8215 (N_8215,N_7698,N_7873);
xnor U8216 (N_8216,N_7748,N_7575);
xnor U8217 (N_8217,N_7997,N_7578);
or U8218 (N_8218,N_7673,N_7588);
or U8219 (N_8219,N_7885,N_7883);
or U8220 (N_8220,N_7993,N_7576);
xnor U8221 (N_8221,N_7520,N_7991);
and U8222 (N_8222,N_7849,N_7566);
xnor U8223 (N_8223,N_7586,N_7994);
nand U8224 (N_8224,N_7837,N_7685);
nor U8225 (N_8225,N_7786,N_7795);
nor U8226 (N_8226,N_7734,N_7602);
nor U8227 (N_8227,N_7661,N_7658);
nor U8228 (N_8228,N_7607,N_7559);
or U8229 (N_8229,N_7572,N_7943);
nand U8230 (N_8230,N_7603,N_7532);
or U8231 (N_8231,N_7598,N_7526);
nor U8232 (N_8232,N_7957,N_7694);
or U8233 (N_8233,N_7859,N_7857);
or U8234 (N_8234,N_7954,N_7555);
or U8235 (N_8235,N_7875,N_7864);
or U8236 (N_8236,N_7789,N_7956);
and U8237 (N_8237,N_7762,N_7927);
nand U8238 (N_8238,N_7718,N_7515);
nand U8239 (N_8239,N_7664,N_7590);
nand U8240 (N_8240,N_7579,N_7552);
xor U8241 (N_8241,N_7975,N_7978);
and U8242 (N_8242,N_7773,N_7981);
nor U8243 (N_8243,N_7516,N_7645);
xor U8244 (N_8244,N_7878,N_7667);
xnor U8245 (N_8245,N_7763,N_7690);
or U8246 (N_8246,N_7560,N_7550);
nor U8247 (N_8247,N_7945,N_7654);
xnor U8248 (N_8248,N_7741,N_7777);
or U8249 (N_8249,N_7984,N_7522);
and U8250 (N_8250,N_7940,N_7981);
or U8251 (N_8251,N_7879,N_7774);
nor U8252 (N_8252,N_7882,N_7943);
xor U8253 (N_8253,N_7717,N_7661);
and U8254 (N_8254,N_7678,N_7663);
nor U8255 (N_8255,N_7806,N_7901);
xnor U8256 (N_8256,N_7666,N_7635);
nor U8257 (N_8257,N_7713,N_7550);
nor U8258 (N_8258,N_7539,N_7962);
and U8259 (N_8259,N_7965,N_7957);
nor U8260 (N_8260,N_7931,N_7938);
xor U8261 (N_8261,N_7996,N_7559);
nand U8262 (N_8262,N_7556,N_7572);
nand U8263 (N_8263,N_7636,N_7913);
nor U8264 (N_8264,N_7836,N_7716);
and U8265 (N_8265,N_7692,N_7586);
xnor U8266 (N_8266,N_7524,N_7801);
and U8267 (N_8267,N_7583,N_7703);
nor U8268 (N_8268,N_7603,N_7706);
xor U8269 (N_8269,N_7725,N_7908);
nand U8270 (N_8270,N_7940,N_7890);
and U8271 (N_8271,N_7520,N_7648);
or U8272 (N_8272,N_7835,N_7793);
xor U8273 (N_8273,N_7511,N_7818);
and U8274 (N_8274,N_7822,N_7516);
xor U8275 (N_8275,N_7855,N_7827);
or U8276 (N_8276,N_7675,N_7588);
or U8277 (N_8277,N_7776,N_7927);
nor U8278 (N_8278,N_7652,N_7729);
nand U8279 (N_8279,N_7850,N_7607);
nand U8280 (N_8280,N_7963,N_7704);
and U8281 (N_8281,N_7523,N_7742);
xnor U8282 (N_8282,N_7946,N_7963);
or U8283 (N_8283,N_7940,N_7987);
nor U8284 (N_8284,N_7884,N_7960);
and U8285 (N_8285,N_7733,N_7643);
and U8286 (N_8286,N_7900,N_7677);
and U8287 (N_8287,N_7674,N_7813);
nand U8288 (N_8288,N_7527,N_7732);
xnor U8289 (N_8289,N_7729,N_7789);
and U8290 (N_8290,N_7759,N_7808);
nor U8291 (N_8291,N_7875,N_7811);
xor U8292 (N_8292,N_7606,N_7590);
xnor U8293 (N_8293,N_7697,N_7511);
or U8294 (N_8294,N_7890,N_7887);
and U8295 (N_8295,N_7732,N_7998);
nand U8296 (N_8296,N_7587,N_7868);
and U8297 (N_8297,N_7693,N_7524);
nand U8298 (N_8298,N_7638,N_7773);
nand U8299 (N_8299,N_7841,N_7507);
and U8300 (N_8300,N_7803,N_7551);
nor U8301 (N_8301,N_7861,N_7734);
or U8302 (N_8302,N_7718,N_7774);
or U8303 (N_8303,N_7811,N_7527);
nor U8304 (N_8304,N_7682,N_7615);
or U8305 (N_8305,N_7523,N_7503);
xnor U8306 (N_8306,N_7734,N_7622);
or U8307 (N_8307,N_7907,N_7601);
nor U8308 (N_8308,N_7592,N_7969);
or U8309 (N_8309,N_7611,N_7793);
nor U8310 (N_8310,N_7987,N_7846);
or U8311 (N_8311,N_7987,N_7924);
or U8312 (N_8312,N_7850,N_7939);
nor U8313 (N_8313,N_7680,N_7806);
nor U8314 (N_8314,N_7913,N_7814);
and U8315 (N_8315,N_7776,N_7639);
and U8316 (N_8316,N_7546,N_7793);
xor U8317 (N_8317,N_7962,N_7906);
xor U8318 (N_8318,N_7995,N_7821);
and U8319 (N_8319,N_7868,N_7598);
xnor U8320 (N_8320,N_7855,N_7641);
and U8321 (N_8321,N_7978,N_7730);
xnor U8322 (N_8322,N_7869,N_7512);
and U8323 (N_8323,N_7538,N_7880);
or U8324 (N_8324,N_7700,N_7994);
nor U8325 (N_8325,N_7904,N_7540);
or U8326 (N_8326,N_7642,N_7789);
xnor U8327 (N_8327,N_7506,N_7914);
or U8328 (N_8328,N_7938,N_7598);
and U8329 (N_8329,N_7870,N_7871);
and U8330 (N_8330,N_7929,N_7727);
nand U8331 (N_8331,N_7775,N_7948);
nand U8332 (N_8332,N_7972,N_7988);
nor U8333 (N_8333,N_7773,N_7827);
nand U8334 (N_8334,N_7815,N_7752);
and U8335 (N_8335,N_7662,N_7899);
nor U8336 (N_8336,N_7933,N_7608);
nor U8337 (N_8337,N_7668,N_7510);
xor U8338 (N_8338,N_7836,N_7852);
or U8339 (N_8339,N_7950,N_7656);
or U8340 (N_8340,N_7887,N_7882);
and U8341 (N_8341,N_7947,N_7549);
xor U8342 (N_8342,N_7785,N_7701);
or U8343 (N_8343,N_7895,N_7866);
nor U8344 (N_8344,N_7593,N_7897);
nor U8345 (N_8345,N_7684,N_7671);
nand U8346 (N_8346,N_7602,N_7591);
xnor U8347 (N_8347,N_7528,N_7642);
or U8348 (N_8348,N_7719,N_7897);
xnor U8349 (N_8349,N_7542,N_7923);
nor U8350 (N_8350,N_7799,N_7588);
or U8351 (N_8351,N_7744,N_7903);
and U8352 (N_8352,N_7860,N_7506);
xnor U8353 (N_8353,N_7953,N_7797);
and U8354 (N_8354,N_7623,N_7859);
and U8355 (N_8355,N_7557,N_7888);
nor U8356 (N_8356,N_7889,N_7742);
nand U8357 (N_8357,N_7976,N_7810);
xnor U8358 (N_8358,N_7982,N_7988);
or U8359 (N_8359,N_7614,N_7818);
nor U8360 (N_8360,N_7815,N_7903);
and U8361 (N_8361,N_7735,N_7647);
nor U8362 (N_8362,N_7915,N_7792);
or U8363 (N_8363,N_7919,N_7642);
nor U8364 (N_8364,N_7850,N_7997);
or U8365 (N_8365,N_7963,N_7876);
and U8366 (N_8366,N_7767,N_7672);
or U8367 (N_8367,N_7756,N_7770);
nor U8368 (N_8368,N_7814,N_7533);
or U8369 (N_8369,N_7665,N_7624);
nor U8370 (N_8370,N_7819,N_7961);
xnor U8371 (N_8371,N_7766,N_7583);
xor U8372 (N_8372,N_7866,N_7857);
nor U8373 (N_8373,N_7926,N_7610);
nand U8374 (N_8374,N_7602,N_7616);
nor U8375 (N_8375,N_7593,N_7973);
or U8376 (N_8376,N_7848,N_7520);
nor U8377 (N_8377,N_7902,N_7963);
or U8378 (N_8378,N_7871,N_7906);
xor U8379 (N_8379,N_7650,N_7654);
xnor U8380 (N_8380,N_7641,N_7531);
nor U8381 (N_8381,N_7710,N_7827);
xnor U8382 (N_8382,N_7901,N_7965);
or U8383 (N_8383,N_7639,N_7737);
nor U8384 (N_8384,N_7882,N_7852);
nand U8385 (N_8385,N_7716,N_7632);
nor U8386 (N_8386,N_7822,N_7580);
or U8387 (N_8387,N_7900,N_7684);
xnor U8388 (N_8388,N_7681,N_7775);
nand U8389 (N_8389,N_7541,N_7977);
nor U8390 (N_8390,N_7559,N_7991);
nor U8391 (N_8391,N_7649,N_7987);
nor U8392 (N_8392,N_7563,N_7841);
and U8393 (N_8393,N_7991,N_7725);
or U8394 (N_8394,N_7504,N_7949);
or U8395 (N_8395,N_7503,N_7707);
nand U8396 (N_8396,N_7986,N_7684);
nor U8397 (N_8397,N_7721,N_7952);
xnor U8398 (N_8398,N_7657,N_7759);
nor U8399 (N_8399,N_7853,N_7745);
nor U8400 (N_8400,N_7949,N_7515);
xnor U8401 (N_8401,N_7994,N_7537);
xor U8402 (N_8402,N_7793,N_7836);
nor U8403 (N_8403,N_7549,N_7606);
nand U8404 (N_8404,N_7890,N_7733);
nand U8405 (N_8405,N_7680,N_7649);
xor U8406 (N_8406,N_7820,N_7720);
and U8407 (N_8407,N_7880,N_7575);
or U8408 (N_8408,N_7748,N_7774);
and U8409 (N_8409,N_7881,N_7769);
xnor U8410 (N_8410,N_7502,N_7990);
or U8411 (N_8411,N_7926,N_7817);
or U8412 (N_8412,N_7503,N_7802);
xnor U8413 (N_8413,N_7972,N_7531);
or U8414 (N_8414,N_7552,N_7591);
and U8415 (N_8415,N_7962,N_7926);
xnor U8416 (N_8416,N_7875,N_7809);
xnor U8417 (N_8417,N_7934,N_7621);
xor U8418 (N_8418,N_7840,N_7632);
nor U8419 (N_8419,N_7943,N_7525);
nor U8420 (N_8420,N_7738,N_7839);
and U8421 (N_8421,N_7728,N_7706);
or U8422 (N_8422,N_7635,N_7859);
and U8423 (N_8423,N_7541,N_7797);
nor U8424 (N_8424,N_7810,N_7605);
and U8425 (N_8425,N_7866,N_7722);
xor U8426 (N_8426,N_7564,N_7888);
nor U8427 (N_8427,N_7776,N_7503);
xnor U8428 (N_8428,N_7818,N_7879);
and U8429 (N_8429,N_7677,N_7979);
or U8430 (N_8430,N_7562,N_7889);
xor U8431 (N_8431,N_7508,N_7754);
and U8432 (N_8432,N_7551,N_7787);
or U8433 (N_8433,N_7743,N_7988);
nand U8434 (N_8434,N_7686,N_7915);
xnor U8435 (N_8435,N_7756,N_7505);
nor U8436 (N_8436,N_7833,N_7710);
or U8437 (N_8437,N_7989,N_7764);
nand U8438 (N_8438,N_7652,N_7849);
and U8439 (N_8439,N_7550,N_7549);
and U8440 (N_8440,N_7598,N_7786);
nand U8441 (N_8441,N_7953,N_7724);
nor U8442 (N_8442,N_7507,N_7536);
nor U8443 (N_8443,N_7642,N_7688);
or U8444 (N_8444,N_7660,N_7811);
and U8445 (N_8445,N_7858,N_7796);
or U8446 (N_8446,N_7991,N_7920);
nand U8447 (N_8447,N_7924,N_7737);
or U8448 (N_8448,N_7977,N_7738);
or U8449 (N_8449,N_7964,N_7688);
and U8450 (N_8450,N_7917,N_7873);
nor U8451 (N_8451,N_7981,N_7529);
and U8452 (N_8452,N_7633,N_7855);
xor U8453 (N_8453,N_7743,N_7519);
nor U8454 (N_8454,N_7772,N_7990);
nor U8455 (N_8455,N_7957,N_7859);
or U8456 (N_8456,N_7627,N_7893);
xor U8457 (N_8457,N_7509,N_7859);
nand U8458 (N_8458,N_7992,N_7514);
and U8459 (N_8459,N_7798,N_7999);
nor U8460 (N_8460,N_7760,N_7691);
nor U8461 (N_8461,N_7592,N_7637);
and U8462 (N_8462,N_7789,N_7648);
xnor U8463 (N_8463,N_7999,N_7522);
or U8464 (N_8464,N_7938,N_7694);
xor U8465 (N_8465,N_7532,N_7735);
nor U8466 (N_8466,N_7528,N_7768);
and U8467 (N_8467,N_7840,N_7844);
and U8468 (N_8468,N_7517,N_7711);
xor U8469 (N_8469,N_7809,N_7595);
xnor U8470 (N_8470,N_7821,N_7564);
nor U8471 (N_8471,N_7681,N_7828);
or U8472 (N_8472,N_7532,N_7979);
xor U8473 (N_8473,N_7587,N_7824);
nor U8474 (N_8474,N_7967,N_7522);
or U8475 (N_8475,N_7606,N_7733);
xnor U8476 (N_8476,N_7525,N_7882);
or U8477 (N_8477,N_7537,N_7723);
xor U8478 (N_8478,N_7914,N_7836);
nand U8479 (N_8479,N_7509,N_7588);
and U8480 (N_8480,N_7743,N_7730);
or U8481 (N_8481,N_7616,N_7721);
xnor U8482 (N_8482,N_7796,N_7957);
nor U8483 (N_8483,N_7571,N_7872);
nor U8484 (N_8484,N_7574,N_7798);
nand U8485 (N_8485,N_7976,N_7803);
nor U8486 (N_8486,N_7710,N_7787);
or U8487 (N_8487,N_7972,N_7755);
or U8488 (N_8488,N_7684,N_7613);
or U8489 (N_8489,N_7558,N_7934);
and U8490 (N_8490,N_7911,N_7562);
nor U8491 (N_8491,N_7822,N_7986);
or U8492 (N_8492,N_7675,N_7536);
and U8493 (N_8493,N_7864,N_7985);
or U8494 (N_8494,N_7620,N_7882);
or U8495 (N_8495,N_7949,N_7857);
nor U8496 (N_8496,N_7709,N_7995);
nor U8497 (N_8497,N_7517,N_7910);
and U8498 (N_8498,N_7673,N_7740);
nand U8499 (N_8499,N_7601,N_7511);
or U8500 (N_8500,N_8215,N_8444);
or U8501 (N_8501,N_8009,N_8211);
nand U8502 (N_8502,N_8259,N_8164);
nor U8503 (N_8503,N_8248,N_8396);
nand U8504 (N_8504,N_8468,N_8306);
or U8505 (N_8505,N_8350,N_8068);
nor U8506 (N_8506,N_8162,N_8261);
or U8507 (N_8507,N_8447,N_8325);
nand U8508 (N_8508,N_8385,N_8286);
nand U8509 (N_8509,N_8253,N_8270);
and U8510 (N_8510,N_8207,N_8356);
nand U8511 (N_8511,N_8199,N_8373);
and U8512 (N_8512,N_8171,N_8170);
or U8513 (N_8513,N_8242,N_8332);
xnor U8514 (N_8514,N_8172,N_8069);
nand U8515 (N_8515,N_8309,N_8065);
and U8516 (N_8516,N_8456,N_8222);
xnor U8517 (N_8517,N_8056,N_8363);
xor U8518 (N_8518,N_8369,N_8123);
nor U8519 (N_8519,N_8320,N_8094);
and U8520 (N_8520,N_8487,N_8036);
and U8521 (N_8521,N_8146,N_8438);
nor U8522 (N_8522,N_8221,N_8074);
nor U8523 (N_8523,N_8187,N_8347);
nand U8524 (N_8524,N_8186,N_8359);
or U8525 (N_8525,N_8411,N_8459);
nor U8526 (N_8526,N_8218,N_8430);
and U8527 (N_8527,N_8158,N_8257);
and U8528 (N_8528,N_8434,N_8011);
and U8529 (N_8529,N_8498,N_8395);
and U8530 (N_8530,N_8001,N_8446);
nand U8531 (N_8531,N_8081,N_8274);
and U8532 (N_8532,N_8156,N_8103);
nor U8533 (N_8533,N_8338,N_8079);
nand U8534 (N_8534,N_8279,N_8098);
or U8535 (N_8535,N_8161,N_8254);
nor U8536 (N_8536,N_8108,N_8436);
nand U8537 (N_8537,N_8165,N_8097);
and U8538 (N_8538,N_8497,N_8002);
and U8539 (N_8539,N_8071,N_8299);
xor U8540 (N_8540,N_8173,N_8365);
xnor U8541 (N_8541,N_8155,N_8387);
xnor U8542 (N_8542,N_8390,N_8475);
nand U8543 (N_8543,N_8301,N_8063);
or U8544 (N_8544,N_8424,N_8083);
nand U8545 (N_8545,N_8303,N_8185);
nor U8546 (N_8546,N_8288,N_8157);
and U8547 (N_8547,N_8217,N_8489);
nor U8548 (N_8548,N_8085,N_8353);
and U8549 (N_8549,N_8361,N_8314);
nor U8550 (N_8550,N_8372,N_8328);
xor U8551 (N_8551,N_8159,N_8141);
xnor U8552 (N_8552,N_8180,N_8029);
or U8553 (N_8553,N_8110,N_8214);
nor U8554 (N_8554,N_8250,N_8375);
xor U8555 (N_8555,N_8414,N_8048);
nand U8556 (N_8556,N_8023,N_8357);
nand U8557 (N_8557,N_8236,N_8243);
xnor U8558 (N_8558,N_8428,N_8174);
nor U8559 (N_8559,N_8417,N_8310);
nand U8560 (N_8560,N_8256,N_8196);
nand U8561 (N_8561,N_8143,N_8037);
or U8562 (N_8562,N_8179,N_8017);
nor U8563 (N_8563,N_8234,N_8084);
or U8564 (N_8564,N_8008,N_8419);
and U8565 (N_8565,N_8095,N_8488);
nand U8566 (N_8566,N_8479,N_8154);
nand U8567 (N_8567,N_8160,N_8412);
or U8568 (N_8568,N_8176,N_8483);
nor U8569 (N_8569,N_8491,N_8241);
xor U8570 (N_8570,N_8038,N_8282);
nand U8571 (N_8571,N_8237,N_8111);
xor U8572 (N_8572,N_8461,N_8151);
nand U8573 (N_8573,N_8230,N_8007);
nor U8574 (N_8574,N_8404,N_8202);
xnor U8575 (N_8575,N_8478,N_8235);
nor U8576 (N_8576,N_8484,N_8142);
xnor U8577 (N_8577,N_8093,N_8399);
xnor U8578 (N_8578,N_8408,N_8219);
nand U8579 (N_8579,N_8284,N_8169);
nand U8580 (N_8580,N_8494,N_8140);
nor U8581 (N_8581,N_8255,N_8191);
nor U8582 (N_8582,N_8311,N_8358);
xor U8583 (N_8583,N_8272,N_8212);
nor U8584 (N_8584,N_8178,N_8465);
and U8585 (N_8585,N_8400,N_8200);
nand U8586 (N_8586,N_8067,N_8326);
xnor U8587 (N_8587,N_8490,N_8495);
nor U8588 (N_8588,N_8120,N_8443);
or U8589 (N_8589,N_8440,N_8295);
or U8590 (N_8590,N_8062,N_8226);
and U8591 (N_8591,N_8168,N_8109);
nand U8592 (N_8592,N_8124,N_8289);
nor U8593 (N_8593,N_8045,N_8485);
xor U8594 (N_8594,N_8136,N_8360);
and U8595 (N_8595,N_8264,N_8405);
or U8596 (N_8596,N_8030,N_8294);
nand U8597 (N_8597,N_8184,N_8113);
and U8598 (N_8598,N_8188,N_8476);
or U8599 (N_8599,N_8026,N_8285);
xnor U8600 (N_8600,N_8381,N_8075);
or U8601 (N_8601,N_8371,N_8380);
and U8602 (N_8602,N_8216,N_8132);
xnor U8603 (N_8603,N_8334,N_8394);
nand U8604 (N_8604,N_8182,N_8383);
and U8605 (N_8605,N_8229,N_8398);
or U8606 (N_8606,N_8177,N_8096);
nor U8607 (N_8607,N_8304,N_8046);
or U8608 (N_8608,N_8072,N_8031);
nand U8609 (N_8609,N_8016,N_8416);
xor U8610 (N_8610,N_8148,N_8102);
or U8611 (N_8611,N_8402,N_8233);
or U8612 (N_8612,N_8342,N_8413);
nand U8613 (N_8613,N_8238,N_8344);
and U8614 (N_8614,N_8025,N_8379);
nand U8615 (N_8615,N_8251,N_8189);
or U8616 (N_8616,N_8422,N_8429);
nor U8617 (N_8617,N_8013,N_8175);
nand U8618 (N_8618,N_8012,N_8442);
or U8619 (N_8619,N_8327,N_8492);
xnor U8620 (N_8620,N_8323,N_8228);
and U8621 (N_8621,N_8335,N_8122);
xnor U8622 (N_8622,N_8374,N_8100);
xor U8623 (N_8623,N_8450,N_8015);
nor U8624 (N_8624,N_8376,N_8496);
nor U8625 (N_8625,N_8198,N_8423);
nor U8626 (N_8626,N_8252,N_8104);
nor U8627 (N_8627,N_8280,N_8401);
nor U8628 (N_8628,N_8076,N_8433);
or U8629 (N_8629,N_8336,N_8138);
or U8630 (N_8630,N_8339,N_8277);
and U8631 (N_8631,N_8115,N_8203);
xnor U8632 (N_8632,N_8147,N_8055);
and U8633 (N_8633,N_8354,N_8066);
or U8634 (N_8634,N_8051,N_8239);
or U8635 (N_8635,N_8089,N_8437);
and U8636 (N_8636,N_8266,N_8206);
and U8637 (N_8637,N_8119,N_8366);
or U8638 (N_8638,N_8149,N_8471);
or U8639 (N_8639,N_8118,N_8027);
nor U8640 (N_8640,N_8054,N_8247);
nor U8641 (N_8641,N_8273,N_8091);
or U8642 (N_8642,N_8061,N_8127);
nand U8643 (N_8643,N_8477,N_8397);
and U8644 (N_8644,N_8302,N_8137);
nor U8645 (N_8645,N_8033,N_8278);
and U8646 (N_8646,N_8153,N_8192);
nor U8647 (N_8647,N_8425,N_8034);
or U8648 (N_8648,N_8106,N_8349);
nor U8649 (N_8649,N_8486,N_8355);
and U8650 (N_8650,N_8362,N_8070);
nor U8651 (N_8651,N_8393,N_8469);
xnor U8652 (N_8652,N_8409,N_8205);
xor U8653 (N_8653,N_8297,N_8194);
and U8654 (N_8654,N_8117,N_8445);
xor U8655 (N_8655,N_8004,N_8131);
or U8656 (N_8656,N_8467,N_8080);
nor U8657 (N_8657,N_8455,N_8466);
or U8658 (N_8658,N_8453,N_8431);
nor U8659 (N_8659,N_8145,N_8300);
xor U8660 (N_8660,N_8032,N_8305);
and U8661 (N_8661,N_8435,N_8204);
or U8662 (N_8662,N_8249,N_8193);
nand U8663 (N_8663,N_8276,N_8293);
and U8664 (N_8664,N_8324,N_8421);
xnor U8665 (N_8665,N_8190,N_8322);
or U8666 (N_8666,N_8042,N_8386);
nor U8667 (N_8667,N_8480,N_8473);
nor U8668 (N_8668,N_8377,N_8415);
or U8669 (N_8669,N_8078,N_8000);
or U8670 (N_8670,N_8384,N_8316);
and U8671 (N_8671,N_8364,N_8059);
or U8672 (N_8672,N_8368,N_8317);
and U8673 (N_8673,N_8114,N_8290);
and U8674 (N_8674,N_8382,N_8116);
or U8675 (N_8675,N_8197,N_8039);
nand U8676 (N_8676,N_8313,N_8462);
xor U8677 (N_8677,N_8246,N_8135);
xnor U8678 (N_8678,N_8296,N_8225);
nor U8679 (N_8679,N_8125,N_8133);
or U8680 (N_8680,N_8082,N_8406);
xnor U8681 (N_8681,N_8343,N_8245);
and U8682 (N_8682,N_8231,N_8150);
nand U8683 (N_8683,N_8112,N_8121);
nor U8684 (N_8684,N_8315,N_8057);
and U8685 (N_8685,N_8128,N_8265);
nand U8686 (N_8686,N_8099,N_8060);
or U8687 (N_8687,N_8018,N_8024);
and U8688 (N_8688,N_8388,N_8318);
and U8689 (N_8689,N_8307,N_8333);
nand U8690 (N_8690,N_8134,N_8474);
and U8691 (N_8691,N_8268,N_8014);
and U8692 (N_8692,N_8454,N_8427);
xor U8693 (N_8693,N_8053,N_8420);
xor U8694 (N_8694,N_8352,N_8041);
and U8695 (N_8695,N_8292,N_8210);
nor U8696 (N_8696,N_8232,N_8020);
and U8697 (N_8697,N_8040,N_8224);
nand U8698 (N_8698,N_8340,N_8298);
and U8699 (N_8699,N_8482,N_8330);
and U8700 (N_8700,N_8052,N_8345);
nor U8701 (N_8701,N_8463,N_8451);
or U8702 (N_8702,N_8064,N_8403);
or U8703 (N_8703,N_8088,N_8077);
or U8704 (N_8704,N_8003,N_8049);
nand U8705 (N_8705,N_8346,N_8432);
and U8706 (N_8706,N_8472,N_8439);
or U8707 (N_8707,N_8107,N_8418);
nand U8708 (N_8708,N_8329,N_8050);
nand U8709 (N_8709,N_8129,N_8367);
xnor U8710 (N_8710,N_8308,N_8321);
or U8711 (N_8711,N_8281,N_8258);
nor U8712 (N_8712,N_8220,N_8341);
xnor U8713 (N_8713,N_8043,N_8044);
xnor U8714 (N_8714,N_8319,N_8458);
or U8715 (N_8715,N_8410,N_8240);
nor U8716 (N_8716,N_8152,N_8092);
and U8717 (N_8717,N_8005,N_8021);
xnor U8718 (N_8718,N_8378,N_8105);
nor U8719 (N_8719,N_8337,N_8291);
xnor U8720 (N_8720,N_8260,N_8213);
nand U8721 (N_8721,N_8389,N_8262);
xnor U8722 (N_8722,N_8201,N_8181);
nand U8723 (N_8723,N_8195,N_8167);
xnor U8724 (N_8724,N_8087,N_8275);
nor U8725 (N_8725,N_8287,N_8441);
or U8726 (N_8726,N_8392,N_8090);
and U8727 (N_8727,N_8139,N_8058);
or U8728 (N_8728,N_8035,N_8022);
nand U8729 (N_8729,N_8348,N_8460);
nand U8730 (N_8730,N_8144,N_8163);
and U8731 (N_8731,N_8209,N_8227);
nor U8732 (N_8732,N_8166,N_8493);
or U8733 (N_8733,N_8331,N_8183);
xor U8734 (N_8734,N_8267,N_8499);
and U8735 (N_8735,N_8208,N_8426);
and U8736 (N_8736,N_8073,N_8047);
and U8737 (N_8737,N_8312,N_8101);
xnor U8738 (N_8738,N_8028,N_8126);
and U8739 (N_8739,N_8223,N_8086);
xor U8740 (N_8740,N_8351,N_8464);
xnor U8741 (N_8741,N_8470,N_8010);
or U8742 (N_8742,N_8452,N_8019);
nand U8743 (N_8743,N_8271,N_8391);
nand U8744 (N_8744,N_8006,N_8370);
and U8745 (N_8745,N_8269,N_8244);
and U8746 (N_8746,N_8448,N_8130);
and U8747 (N_8747,N_8449,N_8457);
or U8748 (N_8748,N_8407,N_8263);
or U8749 (N_8749,N_8283,N_8481);
or U8750 (N_8750,N_8339,N_8045);
or U8751 (N_8751,N_8499,N_8189);
xor U8752 (N_8752,N_8367,N_8481);
or U8753 (N_8753,N_8077,N_8294);
and U8754 (N_8754,N_8237,N_8204);
and U8755 (N_8755,N_8142,N_8279);
nor U8756 (N_8756,N_8119,N_8341);
nor U8757 (N_8757,N_8225,N_8473);
nor U8758 (N_8758,N_8363,N_8060);
nand U8759 (N_8759,N_8167,N_8162);
nor U8760 (N_8760,N_8303,N_8238);
xnor U8761 (N_8761,N_8057,N_8178);
and U8762 (N_8762,N_8009,N_8049);
and U8763 (N_8763,N_8143,N_8291);
or U8764 (N_8764,N_8207,N_8126);
and U8765 (N_8765,N_8363,N_8112);
nand U8766 (N_8766,N_8272,N_8048);
nand U8767 (N_8767,N_8085,N_8205);
or U8768 (N_8768,N_8298,N_8495);
nand U8769 (N_8769,N_8071,N_8261);
or U8770 (N_8770,N_8248,N_8268);
nand U8771 (N_8771,N_8006,N_8186);
or U8772 (N_8772,N_8379,N_8448);
xor U8773 (N_8773,N_8475,N_8221);
xor U8774 (N_8774,N_8283,N_8331);
or U8775 (N_8775,N_8194,N_8461);
and U8776 (N_8776,N_8006,N_8079);
and U8777 (N_8777,N_8275,N_8145);
nor U8778 (N_8778,N_8348,N_8344);
and U8779 (N_8779,N_8231,N_8115);
nor U8780 (N_8780,N_8483,N_8152);
and U8781 (N_8781,N_8072,N_8207);
nand U8782 (N_8782,N_8427,N_8452);
xor U8783 (N_8783,N_8300,N_8204);
nor U8784 (N_8784,N_8323,N_8269);
or U8785 (N_8785,N_8041,N_8248);
nor U8786 (N_8786,N_8207,N_8073);
xnor U8787 (N_8787,N_8201,N_8358);
xnor U8788 (N_8788,N_8189,N_8459);
nand U8789 (N_8789,N_8309,N_8195);
and U8790 (N_8790,N_8371,N_8259);
or U8791 (N_8791,N_8290,N_8192);
nand U8792 (N_8792,N_8085,N_8069);
and U8793 (N_8793,N_8284,N_8303);
nor U8794 (N_8794,N_8442,N_8207);
or U8795 (N_8795,N_8201,N_8250);
nand U8796 (N_8796,N_8432,N_8349);
xnor U8797 (N_8797,N_8210,N_8192);
nor U8798 (N_8798,N_8494,N_8417);
nor U8799 (N_8799,N_8327,N_8477);
nor U8800 (N_8800,N_8037,N_8106);
nor U8801 (N_8801,N_8455,N_8083);
and U8802 (N_8802,N_8115,N_8140);
xor U8803 (N_8803,N_8068,N_8241);
or U8804 (N_8804,N_8424,N_8007);
nand U8805 (N_8805,N_8233,N_8388);
nand U8806 (N_8806,N_8473,N_8070);
xor U8807 (N_8807,N_8459,N_8436);
or U8808 (N_8808,N_8118,N_8285);
xnor U8809 (N_8809,N_8329,N_8100);
and U8810 (N_8810,N_8113,N_8329);
nor U8811 (N_8811,N_8310,N_8416);
xor U8812 (N_8812,N_8480,N_8377);
xnor U8813 (N_8813,N_8280,N_8028);
or U8814 (N_8814,N_8210,N_8140);
or U8815 (N_8815,N_8332,N_8247);
nor U8816 (N_8816,N_8362,N_8272);
nor U8817 (N_8817,N_8180,N_8362);
or U8818 (N_8818,N_8410,N_8428);
and U8819 (N_8819,N_8330,N_8231);
xnor U8820 (N_8820,N_8186,N_8083);
xor U8821 (N_8821,N_8014,N_8222);
xor U8822 (N_8822,N_8397,N_8430);
or U8823 (N_8823,N_8159,N_8329);
or U8824 (N_8824,N_8025,N_8322);
nor U8825 (N_8825,N_8323,N_8170);
nand U8826 (N_8826,N_8232,N_8119);
nor U8827 (N_8827,N_8347,N_8406);
nand U8828 (N_8828,N_8323,N_8482);
xor U8829 (N_8829,N_8251,N_8382);
or U8830 (N_8830,N_8075,N_8303);
and U8831 (N_8831,N_8033,N_8457);
nor U8832 (N_8832,N_8061,N_8450);
and U8833 (N_8833,N_8479,N_8028);
nand U8834 (N_8834,N_8156,N_8242);
nor U8835 (N_8835,N_8299,N_8376);
xnor U8836 (N_8836,N_8219,N_8180);
and U8837 (N_8837,N_8065,N_8130);
xnor U8838 (N_8838,N_8412,N_8435);
and U8839 (N_8839,N_8324,N_8088);
and U8840 (N_8840,N_8092,N_8389);
nor U8841 (N_8841,N_8262,N_8248);
nor U8842 (N_8842,N_8135,N_8264);
nor U8843 (N_8843,N_8279,N_8478);
nor U8844 (N_8844,N_8103,N_8405);
nor U8845 (N_8845,N_8006,N_8409);
xnor U8846 (N_8846,N_8300,N_8047);
nor U8847 (N_8847,N_8029,N_8451);
nand U8848 (N_8848,N_8015,N_8000);
nor U8849 (N_8849,N_8467,N_8073);
or U8850 (N_8850,N_8082,N_8277);
nand U8851 (N_8851,N_8241,N_8073);
and U8852 (N_8852,N_8243,N_8396);
or U8853 (N_8853,N_8300,N_8376);
and U8854 (N_8854,N_8064,N_8071);
nor U8855 (N_8855,N_8340,N_8110);
nor U8856 (N_8856,N_8183,N_8353);
nor U8857 (N_8857,N_8353,N_8454);
nand U8858 (N_8858,N_8355,N_8284);
and U8859 (N_8859,N_8227,N_8037);
xnor U8860 (N_8860,N_8143,N_8452);
and U8861 (N_8861,N_8037,N_8468);
xnor U8862 (N_8862,N_8484,N_8274);
or U8863 (N_8863,N_8148,N_8283);
nor U8864 (N_8864,N_8067,N_8380);
and U8865 (N_8865,N_8118,N_8274);
or U8866 (N_8866,N_8299,N_8027);
or U8867 (N_8867,N_8048,N_8421);
nor U8868 (N_8868,N_8118,N_8070);
xnor U8869 (N_8869,N_8166,N_8221);
and U8870 (N_8870,N_8473,N_8395);
or U8871 (N_8871,N_8479,N_8049);
and U8872 (N_8872,N_8082,N_8231);
and U8873 (N_8873,N_8344,N_8116);
xor U8874 (N_8874,N_8487,N_8454);
and U8875 (N_8875,N_8094,N_8372);
xor U8876 (N_8876,N_8334,N_8161);
or U8877 (N_8877,N_8209,N_8233);
or U8878 (N_8878,N_8270,N_8420);
xnor U8879 (N_8879,N_8124,N_8472);
and U8880 (N_8880,N_8342,N_8035);
nand U8881 (N_8881,N_8211,N_8010);
xor U8882 (N_8882,N_8151,N_8021);
or U8883 (N_8883,N_8436,N_8359);
and U8884 (N_8884,N_8182,N_8099);
or U8885 (N_8885,N_8139,N_8364);
nor U8886 (N_8886,N_8343,N_8023);
and U8887 (N_8887,N_8334,N_8066);
and U8888 (N_8888,N_8425,N_8279);
nor U8889 (N_8889,N_8470,N_8103);
and U8890 (N_8890,N_8068,N_8204);
nor U8891 (N_8891,N_8134,N_8185);
and U8892 (N_8892,N_8443,N_8143);
nor U8893 (N_8893,N_8029,N_8034);
nand U8894 (N_8894,N_8423,N_8251);
or U8895 (N_8895,N_8262,N_8111);
nand U8896 (N_8896,N_8014,N_8478);
xor U8897 (N_8897,N_8353,N_8191);
xor U8898 (N_8898,N_8081,N_8341);
nor U8899 (N_8899,N_8011,N_8378);
nor U8900 (N_8900,N_8058,N_8166);
nor U8901 (N_8901,N_8154,N_8449);
nor U8902 (N_8902,N_8348,N_8162);
nand U8903 (N_8903,N_8226,N_8121);
or U8904 (N_8904,N_8189,N_8299);
nand U8905 (N_8905,N_8164,N_8100);
and U8906 (N_8906,N_8195,N_8291);
nand U8907 (N_8907,N_8484,N_8343);
xor U8908 (N_8908,N_8442,N_8412);
or U8909 (N_8909,N_8428,N_8203);
nand U8910 (N_8910,N_8399,N_8011);
or U8911 (N_8911,N_8357,N_8281);
nand U8912 (N_8912,N_8071,N_8003);
or U8913 (N_8913,N_8087,N_8430);
xor U8914 (N_8914,N_8482,N_8175);
or U8915 (N_8915,N_8129,N_8103);
or U8916 (N_8916,N_8053,N_8193);
nand U8917 (N_8917,N_8257,N_8318);
xnor U8918 (N_8918,N_8320,N_8427);
nand U8919 (N_8919,N_8078,N_8247);
and U8920 (N_8920,N_8103,N_8111);
and U8921 (N_8921,N_8425,N_8255);
xor U8922 (N_8922,N_8239,N_8019);
nor U8923 (N_8923,N_8104,N_8321);
and U8924 (N_8924,N_8239,N_8283);
or U8925 (N_8925,N_8313,N_8420);
or U8926 (N_8926,N_8354,N_8333);
or U8927 (N_8927,N_8152,N_8201);
or U8928 (N_8928,N_8157,N_8252);
xnor U8929 (N_8929,N_8067,N_8288);
or U8930 (N_8930,N_8244,N_8072);
nand U8931 (N_8931,N_8336,N_8273);
or U8932 (N_8932,N_8420,N_8080);
nor U8933 (N_8933,N_8176,N_8351);
nand U8934 (N_8934,N_8460,N_8117);
xor U8935 (N_8935,N_8407,N_8302);
or U8936 (N_8936,N_8305,N_8397);
or U8937 (N_8937,N_8187,N_8273);
or U8938 (N_8938,N_8468,N_8491);
or U8939 (N_8939,N_8481,N_8336);
nand U8940 (N_8940,N_8493,N_8127);
and U8941 (N_8941,N_8201,N_8456);
nand U8942 (N_8942,N_8108,N_8203);
nor U8943 (N_8943,N_8354,N_8053);
xnor U8944 (N_8944,N_8256,N_8105);
nand U8945 (N_8945,N_8369,N_8405);
nand U8946 (N_8946,N_8080,N_8349);
xnor U8947 (N_8947,N_8070,N_8471);
nor U8948 (N_8948,N_8253,N_8308);
or U8949 (N_8949,N_8072,N_8018);
or U8950 (N_8950,N_8323,N_8313);
xnor U8951 (N_8951,N_8360,N_8004);
xnor U8952 (N_8952,N_8302,N_8085);
or U8953 (N_8953,N_8468,N_8458);
or U8954 (N_8954,N_8152,N_8145);
nor U8955 (N_8955,N_8373,N_8472);
or U8956 (N_8956,N_8004,N_8471);
nor U8957 (N_8957,N_8085,N_8468);
and U8958 (N_8958,N_8084,N_8207);
or U8959 (N_8959,N_8443,N_8073);
nand U8960 (N_8960,N_8053,N_8360);
and U8961 (N_8961,N_8128,N_8017);
xnor U8962 (N_8962,N_8338,N_8038);
nor U8963 (N_8963,N_8127,N_8217);
nor U8964 (N_8964,N_8176,N_8481);
nor U8965 (N_8965,N_8022,N_8191);
xnor U8966 (N_8966,N_8172,N_8098);
nor U8967 (N_8967,N_8173,N_8180);
and U8968 (N_8968,N_8037,N_8490);
and U8969 (N_8969,N_8473,N_8324);
xor U8970 (N_8970,N_8162,N_8108);
and U8971 (N_8971,N_8414,N_8188);
nor U8972 (N_8972,N_8476,N_8370);
or U8973 (N_8973,N_8064,N_8424);
nand U8974 (N_8974,N_8172,N_8327);
or U8975 (N_8975,N_8216,N_8487);
nand U8976 (N_8976,N_8190,N_8256);
xnor U8977 (N_8977,N_8205,N_8477);
xor U8978 (N_8978,N_8335,N_8130);
nand U8979 (N_8979,N_8373,N_8142);
nor U8980 (N_8980,N_8277,N_8286);
xor U8981 (N_8981,N_8211,N_8225);
and U8982 (N_8982,N_8054,N_8087);
and U8983 (N_8983,N_8319,N_8394);
or U8984 (N_8984,N_8079,N_8346);
nand U8985 (N_8985,N_8487,N_8423);
xnor U8986 (N_8986,N_8435,N_8230);
or U8987 (N_8987,N_8494,N_8054);
nor U8988 (N_8988,N_8315,N_8389);
or U8989 (N_8989,N_8230,N_8042);
and U8990 (N_8990,N_8265,N_8152);
nand U8991 (N_8991,N_8054,N_8223);
nand U8992 (N_8992,N_8409,N_8034);
and U8993 (N_8993,N_8490,N_8390);
nor U8994 (N_8994,N_8126,N_8414);
nand U8995 (N_8995,N_8292,N_8437);
and U8996 (N_8996,N_8147,N_8218);
and U8997 (N_8997,N_8392,N_8394);
nor U8998 (N_8998,N_8121,N_8275);
xnor U8999 (N_8999,N_8050,N_8438);
nor U9000 (N_9000,N_8524,N_8895);
nand U9001 (N_9001,N_8617,N_8729);
nor U9002 (N_9002,N_8937,N_8784);
or U9003 (N_9003,N_8667,N_8938);
nor U9004 (N_9004,N_8654,N_8745);
nand U9005 (N_9005,N_8616,N_8810);
and U9006 (N_9006,N_8849,N_8580);
nor U9007 (N_9007,N_8546,N_8522);
and U9008 (N_9008,N_8866,N_8998);
and U9009 (N_9009,N_8827,N_8981);
nor U9010 (N_9010,N_8591,N_8531);
and U9011 (N_9011,N_8668,N_8909);
or U9012 (N_9012,N_8852,N_8741);
xor U9013 (N_9013,N_8821,N_8641);
or U9014 (N_9014,N_8525,N_8693);
nand U9015 (N_9015,N_8569,N_8578);
or U9016 (N_9016,N_8588,N_8999);
or U9017 (N_9017,N_8519,N_8664);
nor U9018 (N_9018,N_8747,N_8996);
nand U9019 (N_9019,N_8595,N_8606);
nand U9020 (N_9020,N_8631,N_8990);
nor U9021 (N_9021,N_8708,N_8924);
nand U9022 (N_9022,N_8872,N_8671);
and U9023 (N_9023,N_8750,N_8598);
nand U9024 (N_9024,N_8891,N_8587);
or U9025 (N_9025,N_8828,N_8626);
or U9026 (N_9026,N_8857,N_8893);
nor U9027 (N_9027,N_8984,N_8926);
nand U9028 (N_9028,N_8913,N_8644);
nor U9029 (N_9029,N_8740,N_8607);
nand U9030 (N_9030,N_8545,N_8679);
and U9031 (N_9031,N_8819,N_8972);
and U9032 (N_9032,N_8533,N_8608);
and U9033 (N_9033,N_8503,N_8841);
and U9034 (N_9034,N_8725,N_8783);
nor U9035 (N_9035,N_8513,N_8839);
xor U9036 (N_9036,N_8860,N_8848);
nor U9037 (N_9037,N_8912,N_8951);
nor U9038 (N_9038,N_8798,N_8842);
nor U9039 (N_9039,N_8613,N_8771);
nor U9040 (N_9040,N_8597,N_8734);
nand U9041 (N_9041,N_8730,N_8583);
nor U9042 (N_9042,N_8619,N_8553);
xnor U9043 (N_9043,N_8562,N_8892);
or U9044 (N_9044,N_8831,N_8551);
or U9045 (N_9045,N_8888,N_8901);
or U9046 (N_9046,N_8712,N_8635);
nand U9047 (N_9047,N_8801,N_8838);
and U9048 (N_9048,N_8956,N_8584);
nand U9049 (N_9049,N_8820,N_8911);
nor U9050 (N_9050,N_8690,N_8976);
or U9051 (N_9051,N_8508,N_8518);
nand U9052 (N_9052,N_8510,N_8705);
nand U9053 (N_9053,N_8925,N_8601);
or U9054 (N_9054,N_8694,N_8931);
nor U9055 (N_9055,N_8878,N_8772);
xor U9056 (N_9056,N_8794,N_8769);
nand U9057 (N_9057,N_8719,N_8565);
xnor U9058 (N_9058,N_8630,N_8582);
or U9059 (N_9059,N_8793,N_8709);
and U9060 (N_9060,N_8920,N_8670);
nor U9061 (N_9061,N_8677,N_8995);
nand U9062 (N_9062,N_8855,N_8986);
or U9063 (N_9063,N_8536,N_8941);
nor U9064 (N_9064,N_8555,N_8977);
xor U9065 (N_9065,N_8899,N_8908);
and U9066 (N_9066,N_8685,N_8672);
or U9067 (N_9067,N_8916,N_8678);
nor U9068 (N_9068,N_8614,N_8814);
nor U9069 (N_9069,N_8970,N_8540);
nand U9070 (N_9070,N_8564,N_8826);
and U9071 (N_9071,N_8952,N_8516);
nand U9072 (N_9072,N_8538,N_8835);
xor U9073 (N_9073,N_8549,N_8944);
nor U9074 (N_9074,N_8770,N_8577);
and U9075 (N_9075,N_8773,N_8706);
and U9076 (N_9076,N_8684,N_8890);
and U9077 (N_9077,N_8966,N_8816);
xnor U9078 (N_9078,N_8699,N_8700);
or U9079 (N_9079,N_8505,N_8586);
or U9080 (N_9080,N_8932,N_8638);
and U9081 (N_9081,N_8746,N_8596);
nand U9082 (N_9082,N_8779,N_8877);
xnor U9083 (N_9083,N_8713,N_8789);
xnor U9084 (N_9084,N_8876,N_8550);
nand U9085 (N_9085,N_8942,N_8830);
nor U9086 (N_9086,N_8864,N_8581);
nand U9087 (N_9087,N_8882,N_8721);
xnor U9088 (N_9088,N_8558,N_8948);
nand U9089 (N_9089,N_8620,N_8874);
xor U9090 (N_9090,N_8547,N_8760);
or U9091 (N_9091,N_8632,N_8526);
and U9092 (N_9092,N_8680,N_8755);
nand U9093 (N_9093,N_8511,N_8724);
nor U9094 (N_9094,N_8930,N_8529);
nand U9095 (N_9095,N_8949,N_8718);
nand U9096 (N_9096,N_8844,N_8959);
nor U9097 (N_9097,N_8947,N_8845);
and U9098 (N_9098,N_8714,N_8850);
nor U9099 (N_9099,N_8994,N_8824);
and U9100 (N_9100,N_8840,N_8940);
nor U9101 (N_9101,N_8862,N_8572);
nor U9102 (N_9102,N_8665,N_8687);
and U9103 (N_9103,N_8707,N_8504);
nand U9104 (N_9104,N_8957,N_8918);
or U9105 (N_9105,N_8961,N_8590);
nand U9106 (N_9106,N_8650,N_8711);
nor U9107 (N_9107,N_8813,N_8846);
or U9108 (N_9108,N_8847,N_8958);
nand U9109 (N_9109,N_8933,N_8871);
nor U9110 (N_9110,N_8702,N_8946);
nor U9111 (N_9111,N_8682,N_8921);
and U9112 (N_9112,N_8800,N_8557);
and U9113 (N_9113,N_8865,N_8753);
and U9114 (N_9114,N_8535,N_8778);
nor U9115 (N_9115,N_8615,N_8731);
nor U9116 (N_9116,N_8870,N_8715);
nor U9117 (N_9117,N_8738,N_8589);
and U9118 (N_9118,N_8736,N_8894);
nor U9119 (N_9119,N_8649,N_8853);
xor U9120 (N_9120,N_8543,N_8502);
or U9121 (N_9121,N_8744,N_8752);
or U9122 (N_9122,N_8636,N_8517);
nor U9123 (N_9123,N_8610,N_8811);
nor U9124 (N_9124,N_8861,N_8863);
xor U9125 (N_9125,N_8809,N_8657);
and U9126 (N_9126,N_8867,N_8599);
xor U9127 (N_9127,N_8560,N_8544);
nand U9128 (N_9128,N_8960,N_8919);
xnor U9129 (N_9129,N_8927,N_8663);
xor U9130 (N_9130,N_8646,N_8879);
nor U9131 (N_9131,N_8559,N_8506);
nand U9132 (N_9132,N_8751,N_8868);
and U9133 (N_9133,N_8762,N_8640);
nand U9134 (N_9134,N_8507,N_8812);
and U9135 (N_9135,N_8950,N_8757);
nor U9136 (N_9136,N_8997,N_8903);
xor U9137 (N_9137,N_8885,N_8501);
and U9138 (N_9138,N_8897,N_8808);
and U9139 (N_9139,N_8833,N_8520);
nor U9140 (N_9140,N_8603,N_8929);
nand U9141 (N_9141,N_8576,N_8600);
and U9142 (N_9142,N_8799,N_8775);
nor U9143 (N_9143,N_8655,N_8733);
and U9144 (N_9144,N_8509,N_8548);
nand U9145 (N_9145,N_8829,N_8629);
nor U9146 (N_9146,N_8987,N_8945);
or U9147 (N_9147,N_8628,N_8807);
nor U9148 (N_9148,N_8964,N_8859);
and U9149 (N_9149,N_8943,N_8910);
xnor U9150 (N_9150,N_8686,N_8723);
and U9151 (N_9151,N_8634,N_8735);
and U9152 (N_9152,N_8612,N_8716);
and U9153 (N_9153,N_8962,N_8659);
nor U9154 (N_9154,N_8902,N_8579);
and U9155 (N_9155,N_8817,N_8669);
nand U9156 (N_9156,N_8886,N_8537);
xor U9157 (N_9157,N_8512,N_8914);
nor U9158 (N_9158,N_8873,N_8554);
xnor U9159 (N_9159,N_8818,N_8532);
or U9160 (N_9160,N_8652,N_8561);
nor U9161 (N_9161,N_8983,N_8673);
or U9162 (N_9162,N_8623,N_8790);
xor U9163 (N_9163,N_8688,N_8627);
or U9164 (N_9164,N_8720,N_8796);
xor U9165 (N_9165,N_8749,N_8954);
xor U9166 (N_9166,N_8566,N_8993);
xnor U9167 (N_9167,N_8701,N_8975);
xnor U9168 (N_9168,N_8523,N_8500);
nor U9169 (N_9169,N_8661,N_8765);
xnor U9170 (N_9170,N_8756,N_8776);
xor U9171 (N_9171,N_8530,N_8515);
or U9172 (N_9172,N_8574,N_8832);
xor U9173 (N_9173,N_8806,N_8568);
nand U9174 (N_9174,N_8917,N_8887);
and U9175 (N_9175,N_8697,N_8823);
and U9176 (N_9176,N_8639,N_8955);
nor U9177 (N_9177,N_8889,N_8898);
and U9178 (N_9178,N_8834,N_8633);
nand U9179 (N_9179,N_8737,N_8689);
or U9180 (N_9180,N_8928,N_8739);
xor U9181 (N_9181,N_8856,N_8843);
nor U9182 (N_9182,N_8777,N_8567);
nor U9183 (N_9183,N_8974,N_8980);
xnor U9184 (N_9184,N_8978,N_8774);
nand U9185 (N_9185,N_8556,N_8764);
and U9186 (N_9186,N_8754,N_8674);
or U9187 (N_9187,N_8896,N_8732);
nand U9188 (N_9188,N_8988,N_8781);
xor U9189 (N_9189,N_8869,N_8728);
nand U9190 (N_9190,N_8906,N_8683);
nand U9191 (N_9191,N_8883,N_8971);
nor U9192 (N_9192,N_8825,N_8973);
xnor U9193 (N_9193,N_8645,N_8609);
or U9194 (N_9194,N_8982,N_8618);
xor U9195 (N_9195,N_8875,N_8802);
nor U9196 (N_9196,N_8815,N_8726);
nor U9197 (N_9197,N_8768,N_8624);
xnor U9198 (N_9198,N_8851,N_8521);
and U9199 (N_9199,N_8953,N_8662);
xor U9200 (N_9200,N_8743,N_8965);
or U9201 (N_9201,N_8884,N_8904);
nand U9202 (N_9202,N_8611,N_8643);
or U9203 (N_9203,N_8681,N_8822);
xnor U9204 (N_9204,N_8785,N_8722);
and U9205 (N_9205,N_8880,N_8923);
or U9206 (N_9206,N_8967,N_8787);
nor U9207 (N_9207,N_8935,N_8985);
and U9208 (N_9208,N_8979,N_8622);
nor U9209 (N_9209,N_8534,N_8991);
or U9210 (N_9210,N_8936,N_8660);
or U9211 (N_9211,N_8621,N_8858);
nand U9212 (N_9212,N_8593,N_8788);
nor U9213 (N_9213,N_8552,N_8570);
or U9214 (N_9214,N_8767,N_8881);
or U9215 (N_9215,N_8594,N_8642);
xor U9216 (N_9216,N_8695,N_8541);
xor U9217 (N_9217,N_8696,N_8915);
xnor U9218 (N_9218,N_8792,N_8571);
xor U9219 (N_9219,N_8963,N_8648);
and U9220 (N_9220,N_8786,N_8656);
nor U9221 (N_9221,N_8795,N_8761);
or U9222 (N_9222,N_8675,N_8585);
nand U9223 (N_9223,N_8804,N_8758);
or U9224 (N_9224,N_8922,N_8766);
or U9225 (N_9225,N_8698,N_8563);
and U9226 (N_9226,N_8900,N_8637);
xnor U9227 (N_9227,N_8780,N_8836);
nand U9228 (N_9228,N_8748,N_8514);
nand U9229 (N_9229,N_8527,N_8797);
nor U9230 (N_9230,N_8907,N_8969);
and U9231 (N_9231,N_8803,N_8666);
and U9232 (N_9232,N_8717,N_8592);
and U9233 (N_9233,N_8542,N_8605);
nand U9234 (N_9234,N_8968,N_8854);
nand U9235 (N_9235,N_8837,N_8528);
xor U9236 (N_9236,N_8905,N_8604);
xnor U9237 (N_9237,N_8704,N_8692);
and U9238 (N_9238,N_8791,N_8727);
nand U9239 (N_9239,N_8658,N_8602);
nand U9240 (N_9240,N_8989,N_8573);
xor U9241 (N_9241,N_8651,N_8782);
nor U9242 (N_9242,N_8742,N_8759);
or U9243 (N_9243,N_8763,N_8992);
or U9244 (N_9244,N_8653,N_8625);
or U9245 (N_9245,N_8710,N_8676);
xor U9246 (N_9246,N_8939,N_8691);
and U9247 (N_9247,N_8539,N_8934);
or U9248 (N_9248,N_8703,N_8805);
nor U9249 (N_9249,N_8647,N_8575);
nand U9250 (N_9250,N_8883,N_8536);
nor U9251 (N_9251,N_8543,N_8531);
nand U9252 (N_9252,N_8869,N_8603);
nor U9253 (N_9253,N_8971,N_8897);
and U9254 (N_9254,N_8819,N_8886);
nand U9255 (N_9255,N_8855,N_8590);
xor U9256 (N_9256,N_8845,N_8916);
or U9257 (N_9257,N_8706,N_8820);
xor U9258 (N_9258,N_8754,N_8614);
nor U9259 (N_9259,N_8627,N_8577);
nand U9260 (N_9260,N_8890,N_8823);
or U9261 (N_9261,N_8797,N_8518);
nand U9262 (N_9262,N_8646,N_8774);
nand U9263 (N_9263,N_8852,N_8893);
xnor U9264 (N_9264,N_8901,N_8514);
xnor U9265 (N_9265,N_8765,N_8997);
nand U9266 (N_9266,N_8528,N_8968);
and U9267 (N_9267,N_8650,N_8985);
nor U9268 (N_9268,N_8657,N_8804);
xor U9269 (N_9269,N_8511,N_8585);
and U9270 (N_9270,N_8737,N_8816);
nand U9271 (N_9271,N_8667,N_8665);
xnor U9272 (N_9272,N_8660,N_8980);
or U9273 (N_9273,N_8972,N_8627);
xnor U9274 (N_9274,N_8938,N_8996);
nand U9275 (N_9275,N_8652,N_8735);
nor U9276 (N_9276,N_8729,N_8733);
and U9277 (N_9277,N_8537,N_8746);
and U9278 (N_9278,N_8803,N_8688);
xnor U9279 (N_9279,N_8634,N_8851);
xnor U9280 (N_9280,N_8645,N_8621);
nor U9281 (N_9281,N_8674,N_8701);
nor U9282 (N_9282,N_8593,N_8507);
xor U9283 (N_9283,N_8986,N_8690);
or U9284 (N_9284,N_8524,N_8854);
xnor U9285 (N_9285,N_8825,N_8932);
and U9286 (N_9286,N_8916,N_8609);
xor U9287 (N_9287,N_8540,N_8893);
xnor U9288 (N_9288,N_8723,N_8524);
xnor U9289 (N_9289,N_8712,N_8693);
xnor U9290 (N_9290,N_8638,N_8620);
nor U9291 (N_9291,N_8590,N_8864);
xnor U9292 (N_9292,N_8989,N_8652);
xor U9293 (N_9293,N_8693,N_8858);
and U9294 (N_9294,N_8640,N_8544);
nand U9295 (N_9295,N_8612,N_8503);
and U9296 (N_9296,N_8809,N_8830);
xnor U9297 (N_9297,N_8701,N_8828);
nor U9298 (N_9298,N_8881,N_8786);
and U9299 (N_9299,N_8795,N_8991);
nor U9300 (N_9300,N_8820,N_8891);
xor U9301 (N_9301,N_8517,N_8747);
xnor U9302 (N_9302,N_8597,N_8571);
nand U9303 (N_9303,N_8778,N_8569);
nor U9304 (N_9304,N_8654,N_8752);
or U9305 (N_9305,N_8755,N_8511);
and U9306 (N_9306,N_8532,N_8624);
or U9307 (N_9307,N_8739,N_8520);
and U9308 (N_9308,N_8514,N_8688);
xor U9309 (N_9309,N_8747,N_8575);
or U9310 (N_9310,N_8986,N_8528);
and U9311 (N_9311,N_8617,N_8669);
nor U9312 (N_9312,N_8640,N_8803);
nand U9313 (N_9313,N_8505,N_8689);
or U9314 (N_9314,N_8517,N_8908);
nor U9315 (N_9315,N_8981,N_8557);
xor U9316 (N_9316,N_8848,N_8742);
nand U9317 (N_9317,N_8544,N_8524);
xnor U9318 (N_9318,N_8854,N_8697);
and U9319 (N_9319,N_8726,N_8580);
nor U9320 (N_9320,N_8934,N_8665);
or U9321 (N_9321,N_8700,N_8813);
xnor U9322 (N_9322,N_8767,N_8850);
and U9323 (N_9323,N_8742,N_8863);
nor U9324 (N_9324,N_8764,N_8951);
and U9325 (N_9325,N_8568,N_8772);
nor U9326 (N_9326,N_8570,N_8594);
or U9327 (N_9327,N_8951,N_8954);
nand U9328 (N_9328,N_8569,N_8764);
or U9329 (N_9329,N_8865,N_8851);
nand U9330 (N_9330,N_8532,N_8738);
nor U9331 (N_9331,N_8576,N_8975);
nor U9332 (N_9332,N_8586,N_8821);
and U9333 (N_9333,N_8821,N_8908);
nor U9334 (N_9334,N_8757,N_8944);
xor U9335 (N_9335,N_8800,N_8823);
nor U9336 (N_9336,N_8990,N_8678);
nand U9337 (N_9337,N_8592,N_8926);
and U9338 (N_9338,N_8608,N_8844);
xor U9339 (N_9339,N_8513,N_8626);
or U9340 (N_9340,N_8579,N_8749);
and U9341 (N_9341,N_8799,N_8778);
xor U9342 (N_9342,N_8657,N_8704);
and U9343 (N_9343,N_8577,N_8990);
nor U9344 (N_9344,N_8937,N_8741);
xnor U9345 (N_9345,N_8835,N_8530);
and U9346 (N_9346,N_8903,N_8662);
nand U9347 (N_9347,N_8621,N_8771);
and U9348 (N_9348,N_8800,N_8751);
nor U9349 (N_9349,N_8931,N_8607);
nor U9350 (N_9350,N_8855,N_8966);
xor U9351 (N_9351,N_8691,N_8784);
xor U9352 (N_9352,N_8606,N_8779);
xor U9353 (N_9353,N_8961,N_8640);
or U9354 (N_9354,N_8920,N_8751);
nor U9355 (N_9355,N_8960,N_8633);
nor U9356 (N_9356,N_8874,N_8576);
and U9357 (N_9357,N_8829,N_8547);
nand U9358 (N_9358,N_8781,N_8515);
nor U9359 (N_9359,N_8664,N_8718);
and U9360 (N_9360,N_8592,N_8685);
nor U9361 (N_9361,N_8854,N_8988);
nand U9362 (N_9362,N_8825,N_8502);
and U9363 (N_9363,N_8693,N_8807);
and U9364 (N_9364,N_8938,N_8829);
or U9365 (N_9365,N_8790,N_8938);
and U9366 (N_9366,N_8938,N_8934);
and U9367 (N_9367,N_8692,N_8785);
nand U9368 (N_9368,N_8535,N_8514);
or U9369 (N_9369,N_8837,N_8657);
nor U9370 (N_9370,N_8921,N_8945);
xnor U9371 (N_9371,N_8897,N_8532);
xor U9372 (N_9372,N_8824,N_8769);
or U9373 (N_9373,N_8666,N_8574);
nor U9374 (N_9374,N_8814,N_8952);
nor U9375 (N_9375,N_8585,N_8602);
or U9376 (N_9376,N_8603,N_8755);
and U9377 (N_9377,N_8635,N_8682);
or U9378 (N_9378,N_8734,N_8703);
nor U9379 (N_9379,N_8880,N_8670);
nor U9380 (N_9380,N_8781,N_8792);
xnor U9381 (N_9381,N_8870,N_8622);
nor U9382 (N_9382,N_8940,N_8988);
xnor U9383 (N_9383,N_8782,N_8981);
nand U9384 (N_9384,N_8519,N_8962);
nor U9385 (N_9385,N_8632,N_8517);
nand U9386 (N_9386,N_8875,N_8973);
and U9387 (N_9387,N_8562,N_8563);
or U9388 (N_9388,N_8921,N_8897);
or U9389 (N_9389,N_8889,N_8776);
or U9390 (N_9390,N_8519,N_8710);
nand U9391 (N_9391,N_8863,N_8882);
xor U9392 (N_9392,N_8841,N_8507);
or U9393 (N_9393,N_8721,N_8891);
xor U9394 (N_9394,N_8783,N_8785);
nand U9395 (N_9395,N_8571,N_8666);
and U9396 (N_9396,N_8682,N_8782);
and U9397 (N_9397,N_8802,N_8974);
nor U9398 (N_9398,N_8965,N_8810);
nor U9399 (N_9399,N_8661,N_8810);
and U9400 (N_9400,N_8913,N_8571);
nor U9401 (N_9401,N_8800,N_8704);
or U9402 (N_9402,N_8827,N_8944);
xor U9403 (N_9403,N_8685,N_8855);
xor U9404 (N_9404,N_8652,N_8617);
nor U9405 (N_9405,N_8876,N_8953);
and U9406 (N_9406,N_8897,N_8870);
and U9407 (N_9407,N_8970,N_8662);
and U9408 (N_9408,N_8960,N_8669);
xnor U9409 (N_9409,N_8842,N_8557);
or U9410 (N_9410,N_8876,N_8580);
nor U9411 (N_9411,N_8843,N_8562);
and U9412 (N_9412,N_8829,N_8743);
nor U9413 (N_9413,N_8651,N_8580);
or U9414 (N_9414,N_8670,N_8824);
xor U9415 (N_9415,N_8829,N_8559);
nor U9416 (N_9416,N_8619,N_8833);
xnor U9417 (N_9417,N_8766,N_8837);
and U9418 (N_9418,N_8768,N_8593);
and U9419 (N_9419,N_8942,N_8571);
or U9420 (N_9420,N_8822,N_8921);
nand U9421 (N_9421,N_8808,N_8927);
or U9422 (N_9422,N_8823,N_8543);
xor U9423 (N_9423,N_8883,N_8932);
nand U9424 (N_9424,N_8557,N_8625);
and U9425 (N_9425,N_8836,N_8994);
nor U9426 (N_9426,N_8569,N_8562);
xor U9427 (N_9427,N_8813,N_8859);
nand U9428 (N_9428,N_8516,N_8838);
and U9429 (N_9429,N_8826,N_8570);
xor U9430 (N_9430,N_8974,N_8836);
or U9431 (N_9431,N_8688,N_8586);
or U9432 (N_9432,N_8708,N_8719);
and U9433 (N_9433,N_8921,N_8704);
or U9434 (N_9434,N_8977,N_8725);
or U9435 (N_9435,N_8664,N_8560);
nor U9436 (N_9436,N_8656,N_8744);
xnor U9437 (N_9437,N_8948,N_8512);
xnor U9438 (N_9438,N_8507,N_8526);
and U9439 (N_9439,N_8684,N_8904);
nand U9440 (N_9440,N_8573,N_8533);
nor U9441 (N_9441,N_8723,N_8583);
or U9442 (N_9442,N_8747,N_8756);
nor U9443 (N_9443,N_8710,N_8916);
xor U9444 (N_9444,N_8596,N_8897);
and U9445 (N_9445,N_8911,N_8763);
xnor U9446 (N_9446,N_8792,N_8511);
and U9447 (N_9447,N_8922,N_8999);
and U9448 (N_9448,N_8551,N_8724);
or U9449 (N_9449,N_8765,N_8719);
and U9450 (N_9450,N_8998,N_8809);
and U9451 (N_9451,N_8720,N_8575);
nor U9452 (N_9452,N_8509,N_8664);
or U9453 (N_9453,N_8511,N_8519);
and U9454 (N_9454,N_8851,N_8999);
xor U9455 (N_9455,N_8874,N_8579);
and U9456 (N_9456,N_8553,N_8594);
nand U9457 (N_9457,N_8827,N_8529);
xor U9458 (N_9458,N_8958,N_8671);
xor U9459 (N_9459,N_8558,N_8938);
xnor U9460 (N_9460,N_8808,N_8964);
nand U9461 (N_9461,N_8745,N_8800);
or U9462 (N_9462,N_8807,N_8605);
xor U9463 (N_9463,N_8585,N_8628);
and U9464 (N_9464,N_8791,N_8526);
and U9465 (N_9465,N_8942,N_8909);
and U9466 (N_9466,N_8903,N_8515);
nor U9467 (N_9467,N_8574,N_8875);
nand U9468 (N_9468,N_8843,N_8530);
xor U9469 (N_9469,N_8698,N_8734);
xor U9470 (N_9470,N_8795,N_8941);
xor U9471 (N_9471,N_8628,N_8528);
or U9472 (N_9472,N_8939,N_8739);
or U9473 (N_9473,N_8624,N_8891);
and U9474 (N_9474,N_8777,N_8760);
or U9475 (N_9475,N_8612,N_8771);
or U9476 (N_9476,N_8610,N_8783);
xnor U9477 (N_9477,N_8782,N_8539);
nand U9478 (N_9478,N_8978,N_8879);
nor U9479 (N_9479,N_8810,N_8559);
or U9480 (N_9480,N_8890,N_8512);
and U9481 (N_9481,N_8974,N_8666);
xnor U9482 (N_9482,N_8629,N_8568);
xor U9483 (N_9483,N_8866,N_8884);
or U9484 (N_9484,N_8677,N_8585);
or U9485 (N_9485,N_8949,N_8626);
and U9486 (N_9486,N_8844,N_8634);
nor U9487 (N_9487,N_8676,N_8711);
or U9488 (N_9488,N_8576,N_8635);
nor U9489 (N_9489,N_8878,N_8631);
nand U9490 (N_9490,N_8881,N_8567);
or U9491 (N_9491,N_8905,N_8797);
or U9492 (N_9492,N_8691,N_8847);
nor U9493 (N_9493,N_8908,N_8863);
nor U9494 (N_9494,N_8802,N_8961);
and U9495 (N_9495,N_8595,N_8752);
or U9496 (N_9496,N_8633,N_8726);
nand U9497 (N_9497,N_8611,N_8862);
nand U9498 (N_9498,N_8999,N_8839);
nor U9499 (N_9499,N_8951,N_8658);
xnor U9500 (N_9500,N_9281,N_9270);
xor U9501 (N_9501,N_9071,N_9291);
nor U9502 (N_9502,N_9351,N_9364);
and U9503 (N_9503,N_9297,N_9221);
and U9504 (N_9504,N_9305,N_9278);
or U9505 (N_9505,N_9358,N_9078);
nor U9506 (N_9506,N_9186,N_9198);
and U9507 (N_9507,N_9331,N_9347);
and U9508 (N_9508,N_9150,N_9032);
nand U9509 (N_9509,N_9010,N_9246);
and U9510 (N_9510,N_9176,N_9427);
or U9511 (N_9511,N_9315,N_9195);
nor U9512 (N_9512,N_9169,N_9011);
xnor U9513 (N_9513,N_9040,N_9422);
xor U9514 (N_9514,N_9335,N_9452);
nand U9515 (N_9515,N_9109,N_9435);
or U9516 (N_9516,N_9251,N_9482);
and U9517 (N_9517,N_9408,N_9185);
xor U9518 (N_9518,N_9495,N_9135);
or U9519 (N_9519,N_9374,N_9065);
or U9520 (N_9520,N_9208,N_9342);
nand U9521 (N_9521,N_9451,N_9122);
and U9522 (N_9522,N_9031,N_9229);
and U9523 (N_9523,N_9120,N_9289);
nor U9524 (N_9524,N_9379,N_9036);
or U9525 (N_9525,N_9133,N_9403);
nand U9526 (N_9526,N_9405,N_9022);
nor U9527 (N_9527,N_9253,N_9354);
nand U9528 (N_9528,N_9287,N_9077);
and U9529 (N_9529,N_9153,N_9345);
nor U9530 (N_9530,N_9476,N_9144);
and U9531 (N_9531,N_9441,N_9477);
nor U9532 (N_9532,N_9458,N_9045);
nor U9533 (N_9533,N_9430,N_9432);
and U9534 (N_9534,N_9163,N_9230);
nor U9535 (N_9535,N_9444,N_9324);
nand U9536 (N_9536,N_9202,N_9142);
nor U9537 (N_9537,N_9114,N_9419);
and U9538 (N_9538,N_9247,N_9394);
or U9539 (N_9539,N_9279,N_9353);
and U9540 (N_9540,N_9241,N_9099);
or U9541 (N_9541,N_9485,N_9009);
nor U9542 (N_9542,N_9325,N_9119);
or U9543 (N_9543,N_9035,N_9480);
or U9544 (N_9544,N_9004,N_9124);
or U9545 (N_9545,N_9296,N_9172);
xnor U9546 (N_9546,N_9410,N_9129);
or U9547 (N_9547,N_9412,N_9243);
xor U9548 (N_9548,N_9283,N_9396);
and U9549 (N_9549,N_9140,N_9267);
xor U9550 (N_9550,N_9361,N_9222);
nor U9551 (N_9551,N_9062,N_9041);
or U9552 (N_9552,N_9234,N_9029);
and U9553 (N_9553,N_9393,N_9258);
xnor U9554 (N_9554,N_9350,N_9426);
nor U9555 (N_9555,N_9357,N_9164);
nand U9556 (N_9556,N_9486,N_9141);
or U9557 (N_9557,N_9468,N_9170);
and U9558 (N_9558,N_9066,N_9034);
or U9559 (N_9559,N_9276,N_9192);
xor U9560 (N_9560,N_9095,N_9404);
nand U9561 (N_9561,N_9248,N_9074);
nand U9562 (N_9562,N_9388,N_9242);
and U9563 (N_9563,N_9470,N_9178);
and U9564 (N_9564,N_9446,N_9382);
and U9565 (N_9565,N_9064,N_9338);
or U9566 (N_9566,N_9376,N_9337);
or U9567 (N_9567,N_9117,N_9171);
and U9568 (N_9568,N_9021,N_9254);
or U9569 (N_9569,N_9175,N_9341);
xor U9570 (N_9570,N_9151,N_9260);
or U9571 (N_9571,N_9105,N_9323);
or U9572 (N_9572,N_9355,N_9227);
xnor U9573 (N_9573,N_9380,N_9496);
or U9574 (N_9574,N_9216,N_9106);
nor U9575 (N_9575,N_9012,N_9081);
and U9576 (N_9576,N_9282,N_9488);
and U9577 (N_9577,N_9481,N_9235);
nor U9578 (N_9578,N_9413,N_9218);
or U9579 (N_9579,N_9069,N_9056);
nor U9580 (N_9580,N_9052,N_9043);
and U9581 (N_9581,N_9401,N_9453);
and U9582 (N_9582,N_9210,N_9274);
and U9583 (N_9583,N_9344,N_9138);
nand U9584 (N_9584,N_9326,N_9499);
and U9585 (N_9585,N_9256,N_9431);
or U9586 (N_9586,N_9359,N_9205);
nor U9587 (N_9587,N_9424,N_9306);
nand U9588 (N_9588,N_9197,N_9360);
nor U9589 (N_9589,N_9181,N_9352);
nand U9590 (N_9590,N_9107,N_9390);
nand U9591 (N_9591,N_9318,N_9409);
or U9592 (N_9592,N_9113,N_9220);
nor U9593 (N_9593,N_9188,N_9149);
xor U9594 (N_9594,N_9319,N_9059);
nand U9595 (N_9595,N_9094,N_9193);
and U9596 (N_9596,N_9042,N_9311);
nor U9597 (N_9597,N_9051,N_9086);
or U9598 (N_9598,N_9333,N_9136);
or U9599 (N_9599,N_9203,N_9407);
and U9600 (N_9600,N_9255,N_9327);
xnor U9601 (N_9601,N_9005,N_9295);
nor U9602 (N_9602,N_9162,N_9067);
nor U9603 (N_9603,N_9494,N_9356);
or U9604 (N_9604,N_9037,N_9087);
or U9605 (N_9605,N_9317,N_9159);
nor U9606 (N_9606,N_9116,N_9475);
nand U9607 (N_9607,N_9252,N_9284);
nand U9608 (N_9608,N_9083,N_9228);
xor U9609 (N_9609,N_9111,N_9329);
xnor U9610 (N_9610,N_9085,N_9439);
or U9611 (N_9611,N_9101,N_9214);
and U9612 (N_9612,N_9154,N_9006);
nand U9613 (N_9613,N_9349,N_9157);
nand U9614 (N_9614,N_9442,N_9212);
nand U9615 (N_9615,N_9414,N_9240);
nor U9616 (N_9616,N_9402,N_9123);
and U9617 (N_9617,N_9266,N_9058);
and U9618 (N_9618,N_9013,N_9304);
xnor U9619 (N_9619,N_9183,N_9008);
xor U9620 (N_9620,N_9023,N_9148);
nand U9621 (N_9621,N_9425,N_9348);
nor U9622 (N_9622,N_9072,N_9398);
or U9623 (N_9623,N_9118,N_9076);
and U9624 (N_9624,N_9108,N_9082);
nor U9625 (N_9625,N_9238,N_9363);
and U9626 (N_9626,N_9190,N_9201);
and U9627 (N_9627,N_9262,N_9084);
xor U9628 (N_9628,N_9244,N_9060);
and U9629 (N_9629,N_9492,N_9054);
or U9630 (N_9630,N_9307,N_9381);
or U9631 (N_9631,N_9286,N_9204);
xor U9632 (N_9632,N_9265,N_9039);
or U9633 (N_9633,N_9207,N_9303);
nand U9634 (N_9634,N_9182,N_9490);
nand U9635 (N_9635,N_9098,N_9025);
nand U9636 (N_9636,N_9389,N_9301);
and U9637 (N_9637,N_9314,N_9020);
nand U9638 (N_9638,N_9002,N_9237);
or U9639 (N_9639,N_9090,N_9454);
xor U9640 (N_9640,N_9130,N_9395);
nor U9641 (N_9641,N_9434,N_9132);
xnor U9642 (N_9642,N_9433,N_9075);
and U9643 (N_9643,N_9299,N_9316);
nand U9644 (N_9644,N_9156,N_9309);
and U9645 (N_9645,N_9177,N_9330);
or U9646 (N_9646,N_9158,N_9466);
nor U9647 (N_9647,N_9019,N_9196);
nand U9648 (N_9648,N_9383,N_9257);
nor U9649 (N_9649,N_9384,N_9200);
xnor U9650 (N_9650,N_9160,N_9417);
xor U9651 (N_9651,N_9017,N_9450);
nor U9652 (N_9652,N_9143,N_9225);
or U9653 (N_9653,N_9343,N_9100);
nor U9654 (N_9654,N_9102,N_9092);
and U9655 (N_9655,N_9112,N_9493);
nor U9656 (N_9656,N_9302,N_9464);
or U9657 (N_9657,N_9079,N_9027);
and U9658 (N_9658,N_9397,N_9224);
xor U9659 (N_9659,N_9263,N_9165);
nand U9660 (N_9660,N_9217,N_9459);
xor U9661 (N_9661,N_9498,N_9428);
nand U9662 (N_9662,N_9044,N_9211);
xor U9663 (N_9663,N_9440,N_9313);
and U9664 (N_9664,N_9024,N_9231);
or U9665 (N_9665,N_9377,N_9061);
xnor U9666 (N_9666,N_9473,N_9420);
or U9667 (N_9667,N_9047,N_9445);
xnor U9668 (N_9668,N_9128,N_9049);
nor U9669 (N_9669,N_9269,N_9055);
nand U9670 (N_9670,N_9298,N_9187);
nor U9671 (N_9671,N_9063,N_9239);
xnor U9672 (N_9672,N_9001,N_9334);
nor U9673 (N_9673,N_9179,N_9479);
nor U9674 (N_9674,N_9294,N_9411);
and U9675 (N_9675,N_9015,N_9199);
nand U9676 (N_9676,N_9366,N_9336);
and U9677 (N_9677,N_9018,N_9030);
xor U9678 (N_9678,N_9406,N_9073);
xnor U9679 (N_9679,N_9484,N_9497);
nor U9680 (N_9680,N_9455,N_9139);
and U9681 (N_9681,N_9290,N_9438);
or U9682 (N_9682,N_9308,N_9386);
or U9683 (N_9683,N_9489,N_9321);
nor U9684 (N_9684,N_9213,N_9339);
xor U9685 (N_9685,N_9145,N_9028);
or U9686 (N_9686,N_9368,N_9093);
and U9687 (N_9687,N_9166,N_9026);
or U9688 (N_9688,N_9104,N_9264);
or U9689 (N_9689,N_9416,N_9483);
nor U9690 (N_9690,N_9168,N_9249);
xor U9691 (N_9691,N_9194,N_9371);
nand U9692 (N_9692,N_9134,N_9180);
xor U9693 (N_9693,N_9173,N_9460);
nand U9694 (N_9694,N_9385,N_9285);
nor U9695 (N_9695,N_9320,N_9373);
nor U9696 (N_9696,N_9209,N_9191);
nand U9697 (N_9697,N_9288,N_9223);
nor U9698 (N_9698,N_9378,N_9400);
or U9699 (N_9699,N_9206,N_9057);
nand U9700 (N_9700,N_9007,N_9415);
nor U9701 (N_9701,N_9322,N_9399);
nand U9702 (N_9702,N_9226,N_9250);
nor U9703 (N_9703,N_9070,N_9003);
or U9704 (N_9704,N_9469,N_9233);
and U9705 (N_9705,N_9174,N_9272);
xor U9706 (N_9706,N_9467,N_9152);
or U9707 (N_9707,N_9370,N_9300);
or U9708 (N_9708,N_9436,N_9088);
nor U9709 (N_9709,N_9219,N_9392);
nor U9710 (N_9710,N_9465,N_9277);
and U9711 (N_9711,N_9103,N_9462);
xor U9712 (N_9712,N_9391,N_9184);
or U9713 (N_9713,N_9089,N_9280);
nor U9714 (N_9714,N_9312,N_9293);
nor U9715 (N_9715,N_9491,N_9421);
or U9716 (N_9716,N_9155,N_9000);
nor U9717 (N_9717,N_9046,N_9097);
nor U9718 (N_9718,N_9096,N_9091);
and U9719 (N_9719,N_9448,N_9340);
nand U9720 (N_9720,N_9271,N_9332);
and U9721 (N_9721,N_9131,N_9292);
nor U9722 (N_9722,N_9456,N_9259);
or U9723 (N_9723,N_9369,N_9447);
xnor U9724 (N_9724,N_9115,N_9429);
and U9725 (N_9725,N_9437,N_9273);
or U9726 (N_9726,N_9048,N_9275);
and U9727 (N_9727,N_9068,N_9236);
and U9728 (N_9728,N_9033,N_9418);
or U9729 (N_9729,N_9110,N_9457);
or U9730 (N_9730,N_9125,N_9137);
and U9731 (N_9731,N_9050,N_9038);
xnor U9732 (N_9732,N_9423,N_9346);
or U9733 (N_9733,N_9167,N_9443);
nor U9734 (N_9734,N_9189,N_9375);
and U9735 (N_9735,N_9478,N_9474);
or U9736 (N_9736,N_9449,N_9261);
and U9737 (N_9737,N_9127,N_9161);
xor U9738 (N_9738,N_9014,N_9268);
nand U9739 (N_9739,N_9463,N_9080);
nand U9740 (N_9740,N_9487,N_9472);
nand U9741 (N_9741,N_9365,N_9461);
or U9742 (N_9742,N_9387,N_9310);
nor U9743 (N_9743,N_9471,N_9362);
and U9744 (N_9744,N_9053,N_9016);
or U9745 (N_9745,N_9367,N_9147);
or U9746 (N_9746,N_9121,N_9372);
or U9747 (N_9747,N_9146,N_9126);
nand U9748 (N_9748,N_9328,N_9232);
or U9749 (N_9749,N_9215,N_9245);
nor U9750 (N_9750,N_9211,N_9202);
nor U9751 (N_9751,N_9105,N_9030);
nand U9752 (N_9752,N_9422,N_9461);
or U9753 (N_9753,N_9495,N_9318);
xor U9754 (N_9754,N_9478,N_9388);
or U9755 (N_9755,N_9475,N_9435);
xnor U9756 (N_9756,N_9063,N_9287);
nor U9757 (N_9757,N_9065,N_9187);
nand U9758 (N_9758,N_9146,N_9414);
xnor U9759 (N_9759,N_9152,N_9243);
and U9760 (N_9760,N_9350,N_9126);
nand U9761 (N_9761,N_9129,N_9158);
nand U9762 (N_9762,N_9308,N_9019);
xnor U9763 (N_9763,N_9337,N_9355);
xor U9764 (N_9764,N_9149,N_9486);
nor U9765 (N_9765,N_9122,N_9193);
nor U9766 (N_9766,N_9396,N_9128);
xnor U9767 (N_9767,N_9476,N_9455);
nand U9768 (N_9768,N_9479,N_9414);
nand U9769 (N_9769,N_9292,N_9357);
nor U9770 (N_9770,N_9233,N_9372);
and U9771 (N_9771,N_9407,N_9457);
nand U9772 (N_9772,N_9153,N_9166);
nand U9773 (N_9773,N_9352,N_9149);
or U9774 (N_9774,N_9000,N_9410);
xnor U9775 (N_9775,N_9085,N_9268);
or U9776 (N_9776,N_9485,N_9081);
xnor U9777 (N_9777,N_9159,N_9390);
nand U9778 (N_9778,N_9344,N_9021);
nand U9779 (N_9779,N_9224,N_9458);
and U9780 (N_9780,N_9016,N_9136);
xor U9781 (N_9781,N_9197,N_9394);
or U9782 (N_9782,N_9009,N_9045);
nor U9783 (N_9783,N_9042,N_9419);
nand U9784 (N_9784,N_9214,N_9027);
or U9785 (N_9785,N_9134,N_9346);
or U9786 (N_9786,N_9354,N_9429);
xnor U9787 (N_9787,N_9222,N_9275);
xnor U9788 (N_9788,N_9158,N_9463);
or U9789 (N_9789,N_9214,N_9090);
and U9790 (N_9790,N_9037,N_9184);
and U9791 (N_9791,N_9256,N_9320);
and U9792 (N_9792,N_9416,N_9061);
nor U9793 (N_9793,N_9269,N_9284);
xor U9794 (N_9794,N_9205,N_9408);
or U9795 (N_9795,N_9392,N_9193);
nand U9796 (N_9796,N_9014,N_9131);
xnor U9797 (N_9797,N_9459,N_9449);
and U9798 (N_9798,N_9198,N_9472);
nand U9799 (N_9799,N_9494,N_9292);
and U9800 (N_9800,N_9123,N_9292);
nor U9801 (N_9801,N_9063,N_9094);
xnor U9802 (N_9802,N_9219,N_9163);
or U9803 (N_9803,N_9256,N_9439);
nand U9804 (N_9804,N_9008,N_9099);
xor U9805 (N_9805,N_9074,N_9370);
and U9806 (N_9806,N_9178,N_9315);
nand U9807 (N_9807,N_9393,N_9184);
nand U9808 (N_9808,N_9273,N_9132);
or U9809 (N_9809,N_9411,N_9255);
nor U9810 (N_9810,N_9092,N_9440);
or U9811 (N_9811,N_9222,N_9046);
or U9812 (N_9812,N_9298,N_9097);
or U9813 (N_9813,N_9486,N_9303);
and U9814 (N_9814,N_9141,N_9281);
nand U9815 (N_9815,N_9079,N_9348);
nor U9816 (N_9816,N_9154,N_9199);
or U9817 (N_9817,N_9072,N_9130);
nor U9818 (N_9818,N_9130,N_9007);
nand U9819 (N_9819,N_9085,N_9098);
nor U9820 (N_9820,N_9432,N_9376);
nand U9821 (N_9821,N_9113,N_9100);
nand U9822 (N_9822,N_9255,N_9037);
nor U9823 (N_9823,N_9185,N_9454);
xor U9824 (N_9824,N_9294,N_9260);
and U9825 (N_9825,N_9314,N_9397);
nand U9826 (N_9826,N_9283,N_9192);
nor U9827 (N_9827,N_9073,N_9235);
nor U9828 (N_9828,N_9020,N_9426);
or U9829 (N_9829,N_9216,N_9191);
or U9830 (N_9830,N_9436,N_9349);
xnor U9831 (N_9831,N_9240,N_9422);
nor U9832 (N_9832,N_9283,N_9035);
xnor U9833 (N_9833,N_9488,N_9483);
or U9834 (N_9834,N_9374,N_9493);
nor U9835 (N_9835,N_9358,N_9072);
nand U9836 (N_9836,N_9316,N_9189);
nand U9837 (N_9837,N_9077,N_9217);
nand U9838 (N_9838,N_9126,N_9480);
or U9839 (N_9839,N_9371,N_9264);
and U9840 (N_9840,N_9078,N_9048);
and U9841 (N_9841,N_9026,N_9456);
xnor U9842 (N_9842,N_9167,N_9262);
or U9843 (N_9843,N_9461,N_9294);
nand U9844 (N_9844,N_9399,N_9446);
nor U9845 (N_9845,N_9180,N_9241);
nand U9846 (N_9846,N_9360,N_9114);
and U9847 (N_9847,N_9429,N_9118);
and U9848 (N_9848,N_9250,N_9187);
nand U9849 (N_9849,N_9449,N_9228);
nor U9850 (N_9850,N_9401,N_9334);
nor U9851 (N_9851,N_9497,N_9459);
or U9852 (N_9852,N_9131,N_9435);
or U9853 (N_9853,N_9300,N_9101);
and U9854 (N_9854,N_9437,N_9153);
nor U9855 (N_9855,N_9042,N_9487);
nand U9856 (N_9856,N_9025,N_9254);
xor U9857 (N_9857,N_9193,N_9030);
xor U9858 (N_9858,N_9058,N_9349);
nand U9859 (N_9859,N_9115,N_9341);
or U9860 (N_9860,N_9499,N_9291);
nand U9861 (N_9861,N_9462,N_9239);
xor U9862 (N_9862,N_9342,N_9489);
nor U9863 (N_9863,N_9116,N_9002);
and U9864 (N_9864,N_9474,N_9430);
and U9865 (N_9865,N_9092,N_9286);
xor U9866 (N_9866,N_9222,N_9362);
and U9867 (N_9867,N_9294,N_9097);
and U9868 (N_9868,N_9411,N_9345);
xor U9869 (N_9869,N_9329,N_9408);
xor U9870 (N_9870,N_9297,N_9467);
or U9871 (N_9871,N_9326,N_9218);
nor U9872 (N_9872,N_9464,N_9200);
nor U9873 (N_9873,N_9446,N_9395);
xnor U9874 (N_9874,N_9358,N_9401);
nor U9875 (N_9875,N_9392,N_9433);
or U9876 (N_9876,N_9366,N_9455);
nor U9877 (N_9877,N_9204,N_9422);
or U9878 (N_9878,N_9395,N_9034);
nor U9879 (N_9879,N_9358,N_9280);
and U9880 (N_9880,N_9171,N_9183);
xnor U9881 (N_9881,N_9232,N_9314);
xnor U9882 (N_9882,N_9224,N_9306);
xor U9883 (N_9883,N_9147,N_9392);
xor U9884 (N_9884,N_9256,N_9194);
nand U9885 (N_9885,N_9423,N_9195);
or U9886 (N_9886,N_9128,N_9245);
and U9887 (N_9887,N_9272,N_9322);
nor U9888 (N_9888,N_9382,N_9117);
nand U9889 (N_9889,N_9195,N_9324);
and U9890 (N_9890,N_9324,N_9078);
nand U9891 (N_9891,N_9097,N_9176);
nand U9892 (N_9892,N_9241,N_9344);
nor U9893 (N_9893,N_9234,N_9418);
nor U9894 (N_9894,N_9285,N_9411);
or U9895 (N_9895,N_9089,N_9306);
or U9896 (N_9896,N_9117,N_9116);
xor U9897 (N_9897,N_9048,N_9326);
or U9898 (N_9898,N_9179,N_9482);
or U9899 (N_9899,N_9378,N_9414);
xor U9900 (N_9900,N_9211,N_9245);
nor U9901 (N_9901,N_9450,N_9038);
and U9902 (N_9902,N_9266,N_9169);
nor U9903 (N_9903,N_9226,N_9447);
nor U9904 (N_9904,N_9038,N_9352);
xnor U9905 (N_9905,N_9324,N_9399);
and U9906 (N_9906,N_9149,N_9333);
nand U9907 (N_9907,N_9375,N_9058);
nand U9908 (N_9908,N_9185,N_9165);
nand U9909 (N_9909,N_9226,N_9438);
nand U9910 (N_9910,N_9091,N_9266);
xor U9911 (N_9911,N_9104,N_9496);
nand U9912 (N_9912,N_9392,N_9313);
nor U9913 (N_9913,N_9294,N_9427);
nor U9914 (N_9914,N_9281,N_9412);
nor U9915 (N_9915,N_9011,N_9484);
xnor U9916 (N_9916,N_9486,N_9389);
nand U9917 (N_9917,N_9348,N_9270);
or U9918 (N_9918,N_9215,N_9172);
and U9919 (N_9919,N_9274,N_9363);
and U9920 (N_9920,N_9220,N_9201);
nor U9921 (N_9921,N_9051,N_9236);
xor U9922 (N_9922,N_9308,N_9142);
nand U9923 (N_9923,N_9330,N_9286);
xor U9924 (N_9924,N_9475,N_9004);
nand U9925 (N_9925,N_9095,N_9431);
and U9926 (N_9926,N_9052,N_9375);
nand U9927 (N_9927,N_9019,N_9235);
or U9928 (N_9928,N_9262,N_9307);
nand U9929 (N_9929,N_9261,N_9350);
or U9930 (N_9930,N_9322,N_9302);
xnor U9931 (N_9931,N_9104,N_9468);
or U9932 (N_9932,N_9218,N_9228);
nor U9933 (N_9933,N_9217,N_9428);
nor U9934 (N_9934,N_9381,N_9377);
nand U9935 (N_9935,N_9217,N_9034);
nor U9936 (N_9936,N_9062,N_9051);
nand U9937 (N_9937,N_9240,N_9355);
nor U9938 (N_9938,N_9320,N_9015);
xor U9939 (N_9939,N_9370,N_9068);
xor U9940 (N_9940,N_9391,N_9071);
xnor U9941 (N_9941,N_9218,N_9498);
xnor U9942 (N_9942,N_9470,N_9493);
and U9943 (N_9943,N_9205,N_9177);
and U9944 (N_9944,N_9100,N_9042);
nor U9945 (N_9945,N_9173,N_9402);
and U9946 (N_9946,N_9200,N_9434);
nand U9947 (N_9947,N_9326,N_9316);
nor U9948 (N_9948,N_9359,N_9388);
xor U9949 (N_9949,N_9489,N_9431);
and U9950 (N_9950,N_9234,N_9415);
and U9951 (N_9951,N_9148,N_9398);
nand U9952 (N_9952,N_9292,N_9270);
and U9953 (N_9953,N_9357,N_9171);
nand U9954 (N_9954,N_9414,N_9170);
xnor U9955 (N_9955,N_9313,N_9419);
nor U9956 (N_9956,N_9109,N_9374);
nor U9957 (N_9957,N_9480,N_9340);
nor U9958 (N_9958,N_9413,N_9147);
or U9959 (N_9959,N_9324,N_9164);
and U9960 (N_9960,N_9354,N_9478);
xor U9961 (N_9961,N_9086,N_9337);
xor U9962 (N_9962,N_9285,N_9406);
nor U9963 (N_9963,N_9465,N_9306);
nor U9964 (N_9964,N_9435,N_9291);
xnor U9965 (N_9965,N_9235,N_9211);
and U9966 (N_9966,N_9352,N_9353);
and U9967 (N_9967,N_9096,N_9051);
or U9968 (N_9968,N_9390,N_9204);
nand U9969 (N_9969,N_9194,N_9157);
nand U9970 (N_9970,N_9499,N_9129);
xor U9971 (N_9971,N_9406,N_9417);
xnor U9972 (N_9972,N_9108,N_9408);
nand U9973 (N_9973,N_9066,N_9076);
or U9974 (N_9974,N_9137,N_9335);
nor U9975 (N_9975,N_9037,N_9066);
and U9976 (N_9976,N_9220,N_9489);
xor U9977 (N_9977,N_9006,N_9491);
or U9978 (N_9978,N_9227,N_9246);
nand U9979 (N_9979,N_9300,N_9085);
nor U9980 (N_9980,N_9039,N_9031);
or U9981 (N_9981,N_9115,N_9317);
nor U9982 (N_9982,N_9135,N_9234);
nor U9983 (N_9983,N_9105,N_9330);
xor U9984 (N_9984,N_9409,N_9405);
xnor U9985 (N_9985,N_9405,N_9393);
or U9986 (N_9986,N_9293,N_9443);
nor U9987 (N_9987,N_9032,N_9091);
nand U9988 (N_9988,N_9334,N_9333);
nor U9989 (N_9989,N_9189,N_9013);
nand U9990 (N_9990,N_9440,N_9208);
nand U9991 (N_9991,N_9280,N_9243);
or U9992 (N_9992,N_9053,N_9055);
or U9993 (N_9993,N_9213,N_9353);
or U9994 (N_9994,N_9053,N_9336);
or U9995 (N_9995,N_9326,N_9292);
nor U9996 (N_9996,N_9066,N_9114);
nand U9997 (N_9997,N_9169,N_9405);
and U9998 (N_9998,N_9177,N_9371);
or U9999 (N_9999,N_9326,N_9100);
and U10000 (N_10000,N_9687,N_9720);
or U10001 (N_10001,N_9990,N_9949);
nand U10002 (N_10002,N_9946,N_9807);
nor U10003 (N_10003,N_9832,N_9940);
and U10004 (N_10004,N_9831,N_9876);
and U10005 (N_10005,N_9508,N_9746);
or U10006 (N_10006,N_9922,N_9863);
nand U10007 (N_10007,N_9663,N_9523);
nand U10008 (N_10008,N_9972,N_9700);
or U10009 (N_10009,N_9613,N_9809);
nor U10010 (N_10010,N_9742,N_9906);
xnor U10011 (N_10011,N_9651,N_9822);
nor U10012 (N_10012,N_9821,N_9964);
nand U10013 (N_10013,N_9642,N_9704);
or U10014 (N_10014,N_9723,N_9935);
nor U10015 (N_10015,N_9686,N_9997);
xor U10016 (N_10016,N_9971,N_9799);
nor U10017 (N_10017,N_9612,N_9713);
xnor U10018 (N_10018,N_9977,N_9769);
xnor U10019 (N_10019,N_9790,N_9852);
xnor U10020 (N_10020,N_9767,N_9796);
nor U10021 (N_10021,N_9614,N_9744);
and U10022 (N_10022,N_9661,N_9657);
xnor U10023 (N_10023,N_9930,N_9593);
nor U10024 (N_10024,N_9509,N_9762);
nor U10025 (N_10025,N_9816,N_9524);
and U10026 (N_10026,N_9859,N_9953);
or U10027 (N_10027,N_9645,N_9794);
and U10028 (N_10028,N_9679,N_9552);
or U10029 (N_10029,N_9758,N_9888);
xor U10030 (N_10030,N_9916,N_9502);
nor U10031 (N_10031,N_9621,N_9518);
nand U10032 (N_10032,N_9868,N_9564);
and U10033 (N_10033,N_9510,N_9900);
nor U10034 (N_10034,N_9543,N_9941);
and U10035 (N_10035,N_9725,N_9588);
xnor U10036 (N_10036,N_9670,N_9842);
xor U10037 (N_10037,N_9843,N_9748);
nand U10038 (N_10038,N_9681,N_9881);
and U10039 (N_10039,N_9948,N_9653);
xnor U10040 (N_10040,N_9546,N_9622);
and U10041 (N_10041,N_9853,N_9785);
and U10042 (N_10042,N_9995,N_9501);
or U10043 (N_10043,N_9706,N_9715);
and U10044 (N_10044,N_9838,N_9649);
nand U10045 (N_10045,N_9628,N_9553);
nor U10046 (N_10046,N_9895,N_9851);
and U10047 (N_10047,N_9837,N_9734);
and U10048 (N_10048,N_9727,N_9584);
or U10049 (N_10049,N_9560,N_9820);
and U10050 (N_10050,N_9994,N_9992);
and U10051 (N_10051,N_9556,N_9936);
nor U10052 (N_10052,N_9521,N_9908);
and U10053 (N_10053,N_9596,N_9675);
and U10054 (N_10054,N_9591,N_9970);
nor U10055 (N_10055,N_9676,N_9652);
or U10056 (N_10056,N_9824,N_9673);
nor U10057 (N_10057,N_9750,N_9566);
or U10058 (N_10058,N_9708,N_9671);
and U10059 (N_10059,N_9680,N_9893);
and U10060 (N_10060,N_9536,N_9618);
nor U10061 (N_10061,N_9685,N_9656);
and U10062 (N_10062,N_9878,N_9913);
nand U10063 (N_10063,N_9978,N_9860);
xnor U10064 (N_10064,N_9786,N_9836);
nand U10065 (N_10065,N_9697,N_9754);
or U10066 (N_10066,N_9749,N_9619);
xnor U10067 (N_10067,N_9586,N_9782);
nand U10068 (N_10068,N_9915,N_9590);
xor U10069 (N_10069,N_9635,N_9714);
nor U10070 (N_10070,N_9540,N_9846);
nor U10071 (N_10071,N_9887,N_9945);
and U10072 (N_10072,N_9541,N_9818);
and U10073 (N_10073,N_9811,N_9665);
and U10074 (N_10074,N_9629,N_9694);
or U10075 (N_10075,N_9787,N_9610);
and U10076 (N_10076,N_9677,N_9520);
or U10077 (N_10077,N_9531,N_9736);
xor U10078 (N_10078,N_9574,N_9500);
nor U10079 (N_10079,N_9691,N_9827);
xnor U10080 (N_10080,N_9667,N_9793);
nand U10081 (N_10081,N_9624,N_9517);
and U10082 (N_10082,N_9896,N_9587);
nor U10083 (N_10083,N_9885,N_9600);
and U10084 (N_10084,N_9963,N_9766);
or U10085 (N_10085,N_9719,N_9514);
or U10086 (N_10086,N_9578,N_9774);
xor U10087 (N_10087,N_9866,N_9698);
xor U10088 (N_10088,N_9513,N_9639);
nand U10089 (N_10089,N_9542,N_9506);
or U10090 (N_10090,N_9861,N_9530);
and U10091 (N_10091,N_9996,N_9892);
xnor U10092 (N_10092,N_9924,N_9696);
or U10093 (N_10093,N_9711,N_9638);
nand U10094 (N_10094,N_9815,N_9788);
or U10095 (N_10095,N_9538,N_9733);
xnor U10096 (N_10096,N_9801,N_9987);
and U10097 (N_10097,N_9683,N_9575);
xor U10098 (N_10098,N_9780,N_9601);
nor U10099 (N_10099,N_9862,N_9732);
nand U10100 (N_10100,N_9933,N_9874);
nand U10101 (N_10101,N_9839,N_9741);
and U10102 (N_10102,N_9731,N_9561);
xnor U10103 (N_10103,N_9646,N_9898);
nand U10104 (N_10104,N_9738,N_9756);
or U10105 (N_10105,N_9974,N_9841);
nor U10106 (N_10106,N_9737,N_9849);
nor U10107 (N_10107,N_9594,N_9765);
nor U10108 (N_10108,N_9519,N_9966);
nand U10109 (N_10109,N_9961,N_9505);
or U10110 (N_10110,N_9928,N_9802);
nor U10111 (N_10111,N_9558,N_9877);
or U10112 (N_10112,N_9592,N_9772);
and U10113 (N_10113,N_9976,N_9828);
nor U10114 (N_10114,N_9595,N_9724);
nor U10115 (N_10115,N_9636,N_9515);
and U10116 (N_10116,N_9812,N_9773);
xnor U10117 (N_10117,N_9598,N_9739);
or U10118 (N_10118,N_9599,N_9902);
nand U10119 (N_10119,N_9701,N_9938);
or U10120 (N_10120,N_9919,N_9999);
and U10121 (N_10121,N_9779,N_9848);
xor U10122 (N_10122,N_9692,N_9985);
nor U10123 (N_10123,N_9761,N_9835);
and U10124 (N_10124,N_9993,N_9886);
nor U10125 (N_10125,N_9699,N_9817);
xor U10126 (N_10126,N_9979,N_9712);
or U10127 (N_10127,N_9950,N_9764);
nand U10128 (N_10128,N_9504,N_9813);
or U10129 (N_10129,N_9954,N_9927);
nand U10130 (N_10130,N_9729,N_9666);
nor U10131 (N_10131,N_9753,N_9989);
nand U10132 (N_10132,N_9934,N_9525);
or U10133 (N_10133,N_9791,N_9894);
or U10134 (N_10134,N_9641,N_9512);
or U10135 (N_10135,N_9735,N_9583);
xor U10136 (N_10136,N_9923,N_9939);
xnor U10137 (N_10137,N_9830,N_9899);
nand U10138 (N_10138,N_9907,N_9689);
xnor U10139 (N_10139,N_9721,N_9969);
nor U10140 (N_10140,N_9528,N_9882);
nor U10141 (N_10141,N_9983,N_9804);
nor U10142 (N_10142,N_9883,N_9951);
and U10143 (N_10143,N_9722,N_9571);
nand U10144 (N_10144,N_9891,N_9548);
or U10145 (N_10145,N_9570,N_9728);
nand U10146 (N_10146,N_9984,N_9909);
nor U10147 (N_10147,N_9937,N_9965);
or U10148 (N_10148,N_9559,N_9823);
xnor U10149 (N_10149,N_9833,N_9630);
or U10150 (N_10150,N_9959,N_9549);
nor U10151 (N_10151,N_9760,N_9917);
nor U10152 (N_10152,N_9576,N_9751);
or U10153 (N_10153,N_9770,N_9745);
nand U10154 (N_10154,N_9975,N_9633);
and U10155 (N_10155,N_9579,N_9879);
and U10156 (N_10156,N_9942,N_9664);
or U10157 (N_10157,N_9529,N_9957);
xnor U10158 (N_10158,N_9844,N_9625);
and U10159 (N_10159,N_9855,N_9511);
or U10160 (N_10160,N_9623,N_9943);
xor U10161 (N_10161,N_9805,N_9800);
or U10162 (N_10162,N_9932,N_9752);
or U10163 (N_10163,N_9981,N_9929);
nand U10164 (N_10164,N_9674,N_9562);
and U10165 (N_10165,N_9768,N_9555);
nand U10166 (N_10166,N_9608,N_9650);
xor U10167 (N_10167,N_9710,N_9632);
nand U10168 (N_10168,N_9952,N_9707);
and U10169 (N_10169,N_9889,N_9709);
xor U10170 (N_10170,N_9740,N_9897);
xnor U10171 (N_10171,N_9781,N_9778);
nor U10172 (N_10172,N_9703,N_9798);
and U10173 (N_10173,N_9585,N_9516);
xnor U10174 (N_10174,N_9567,N_9806);
xor U10175 (N_10175,N_9551,N_9615);
or U10176 (N_10176,N_9856,N_9718);
nor U10177 (N_10177,N_9668,N_9944);
nand U10178 (N_10178,N_9537,N_9626);
or U10179 (N_10179,N_9991,N_9544);
nor U10180 (N_10180,N_9682,N_9678);
or U10181 (N_10181,N_9534,N_9693);
or U10182 (N_10182,N_9643,N_9602);
and U10183 (N_10183,N_9533,N_9783);
or U10184 (N_10184,N_9955,N_9757);
nor U10185 (N_10185,N_9730,N_9637);
nand U10186 (N_10186,N_9609,N_9865);
nand U10187 (N_10187,N_9926,N_9925);
nand U10188 (N_10188,N_9627,N_9705);
or U10189 (N_10189,N_9931,N_9763);
nand U10190 (N_10190,N_9920,N_9911);
or U10191 (N_10191,N_9998,N_9690);
and U10192 (N_10192,N_9545,N_9755);
xor U10193 (N_10193,N_9577,N_9535);
nor U10194 (N_10194,N_9507,N_9903);
nor U10195 (N_10195,N_9988,N_9960);
nor U10196 (N_10196,N_9947,N_9702);
xnor U10197 (N_10197,N_9648,N_9797);
xor U10198 (N_10198,N_9962,N_9647);
or U10199 (N_10199,N_9611,N_9864);
and U10200 (N_10200,N_9634,N_9914);
nor U10201 (N_10201,N_9726,N_9973);
nor U10202 (N_10202,N_9854,N_9871);
or U10203 (N_10203,N_9829,N_9771);
and U10204 (N_10204,N_9968,N_9554);
or U10205 (N_10205,N_9967,N_9550);
or U10206 (N_10206,N_9688,N_9503);
or U10207 (N_10207,N_9532,N_9921);
xor U10208 (N_10208,N_9858,N_9910);
and U10209 (N_10209,N_9867,N_9526);
nor U10210 (N_10210,N_9644,N_9901);
and U10211 (N_10211,N_9958,N_9617);
nand U10212 (N_10212,N_9655,N_9563);
nor U10213 (N_10213,N_9986,N_9695);
nand U10214 (N_10214,N_9547,N_9759);
xor U10215 (N_10215,N_9880,N_9716);
and U10216 (N_10216,N_9684,N_9569);
xor U10217 (N_10217,N_9825,N_9869);
nand U10218 (N_10218,N_9845,N_9557);
xnor U10219 (N_10219,N_9565,N_9803);
and U10220 (N_10220,N_9884,N_9573);
or U10221 (N_10221,N_9980,N_9572);
nand U10222 (N_10222,N_9912,N_9607);
nor U10223 (N_10223,N_9875,N_9808);
or U10224 (N_10224,N_9776,N_9834);
and U10225 (N_10225,N_9589,N_9597);
xnor U10226 (N_10226,N_9840,N_9603);
and U10227 (N_10227,N_9795,N_9660);
xnor U10228 (N_10228,N_9847,N_9857);
nand U10229 (N_10229,N_9850,N_9640);
nor U10230 (N_10230,N_9982,N_9826);
or U10231 (N_10231,N_9890,N_9905);
xor U10232 (N_10232,N_9747,N_9870);
xor U10233 (N_10233,N_9616,N_9792);
nor U10234 (N_10234,N_9672,N_9581);
or U10235 (N_10235,N_9904,N_9659);
nor U10236 (N_10236,N_9604,N_9789);
and U10237 (N_10237,N_9717,N_9810);
and U10238 (N_10238,N_9539,N_9580);
and U10239 (N_10239,N_9522,N_9606);
nor U10240 (N_10240,N_9775,N_9669);
and U10241 (N_10241,N_9658,N_9568);
nand U10242 (N_10242,N_9956,N_9527);
xor U10243 (N_10243,N_9662,N_9631);
nor U10244 (N_10244,N_9918,N_9777);
xor U10245 (N_10245,N_9872,N_9819);
or U10246 (N_10246,N_9654,N_9873);
nor U10247 (N_10247,N_9582,N_9743);
or U10248 (N_10248,N_9620,N_9814);
xor U10249 (N_10249,N_9605,N_9784);
and U10250 (N_10250,N_9939,N_9786);
or U10251 (N_10251,N_9770,N_9851);
or U10252 (N_10252,N_9554,N_9654);
or U10253 (N_10253,N_9886,N_9506);
or U10254 (N_10254,N_9516,N_9592);
or U10255 (N_10255,N_9963,N_9893);
or U10256 (N_10256,N_9520,N_9936);
and U10257 (N_10257,N_9837,N_9662);
xor U10258 (N_10258,N_9578,N_9795);
nand U10259 (N_10259,N_9738,N_9791);
nor U10260 (N_10260,N_9528,N_9922);
and U10261 (N_10261,N_9930,N_9526);
xor U10262 (N_10262,N_9624,N_9919);
and U10263 (N_10263,N_9878,N_9717);
nand U10264 (N_10264,N_9652,N_9572);
nand U10265 (N_10265,N_9527,N_9703);
nor U10266 (N_10266,N_9888,N_9743);
or U10267 (N_10267,N_9823,N_9841);
nand U10268 (N_10268,N_9629,N_9650);
and U10269 (N_10269,N_9512,N_9936);
nor U10270 (N_10270,N_9788,N_9809);
nand U10271 (N_10271,N_9691,N_9867);
nor U10272 (N_10272,N_9523,N_9558);
or U10273 (N_10273,N_9531,N_9845);
and U10274 (N_10274,N_9898,N_9663);
nand U10275 (N_10275,N_9865,N_9940);
and U10276 (N_10276,N_9957,N_9544);
or U10277 (N_10277,N_9746,N_9674);
and U10278 (N_10278,N_9910,N_9986);
nand U10279 (N_10279,N_9860,N_9715);
xor U10280 (N_10280,N_9580,N_9860);
xor U10281 (N_10281,N_9848,N_9570);
nand U10282 (N_10282,N_9839,N_9524);
nand U10283 (N_10283,N_9901,N_9986);
or U10284 (N_10284,N_9854,N_9993);
xor U10285 (N_10285,N_9867,N_9730);
or U10286 (N_10286,N_9802,N_9640);
and U10287 (N_10287,N_9947,N_9941);
nand U10288 (N_10288,N_9845,N_9591);
and U10289 (N_10289,N_9989,N_9564);
and U10290 (N_10290,N_9818,N_9763);
nor U10291 (N_10291,N_9591,N_9887);
nor U10292 (N_10292,N_9794,N_9751);
and U10293 (N_10293,N_9829,N_9834);
or U10294 (N_10294,N_9737,N_9855);
nor U10295 (N_10295,N_9614,N_9881);
nor U10296 (N_10296,N_9873,N_9529);
nand U10297 (N_10297,N_9811,N_9580);
nor U10298 (N_10298,N_9741,N_9670);
xnor U10299 (N_10299,N_9793,N_9600);
xor U10300 (N_10300,N_9932,N_9553);
nand U10301 (N_10301,N_9948,N_9632);
nor U10302 (N_10302,N_9519,N_9852);
xnor U10303 (N_10303,N_9543,N_9723);
nor U10304 (N_10304,N_9974,N_9746);
nor U10305 (N_10305,N_9742,N_9753);
nor U10306 (N_10306,N_9800,N_9911);
nand U10307 (N_10307,N_9641,N_9568);
xnor U10308 (N_10308,N_9927,N_9911);
or U10309 (N_10309,N_9611,N_9772);
or U10310 (N_10310,N_9998,N_9894);
xnor U10311 (N_10311,N_9870,N_9746);
or U10312 (N_10312,N_9971,N_9672);
nand U10313 (N_10313,N_9791,N_9906);
xnor U10314 (N_10314,N_9862,N_9742);
or U10315 (N_10315,N_9541,N_9809);
nor U10316 (N_10316,N_9606,N_9937);
xnor U10317 (N_10317,N_9763,N_9938);
nor U10318 (N_10318,N_9660,N_9826);
and U10319 (N_10319,N_9827,N_9842);
nor U10320 (N_10320,N_9989,N_9507);
xor U10321 (N_10321,N_9684,N_9992);
and U10322 (N_10322,N_9922,N_9569);
xnor U10323 (N_10323,N_9777,N_9776);
or U10324 (N_10324,N_9716,N_9572);
nor U10325 (N_10325,N_9557,N_9842);
or U10326 (N_10326,N_9807,N_9577);
nand U10327 (N_10327,N_9723,N_9712);
nor U10328 (N_10328,N_9525,N_9854);
nand U10329 (N_10329,N_9613,N_9662);
xnor U10330 (N_10330,N_9974,N_9799);
or U10331 (N_10331,N_9923,N_9680);
nor U10332 (N_10332,N_9550,N_9725);
nand U10333 (N_10333,N_9633,N_9897);
or U10334 (N_10334,N_9794,N_9875);
nand U10335 (N_10335,N_9535,N_9831);
or U10336 (N_10336,N_9657,N_9721);
nor U10337 (N_10337,N_9827,N_9812);
and U10338 (N_10338,N_9788,N_9892);
or U10339 (N_10339,N_9643,N_9856);
xor U10340 (N_10340,N_9727,N_9832);
nor U10341 (N_10341,N_9617,N_9587);
xor U10342 (N_10342,N_9832,N_9576);
nand U10343 (N_10343,N_9554,N_9716);
and U10344 (N_10344,N_9982,N_9956);
nand U10345 (N_10345,N_9799,N_9566);
nor U10346 (N_10346,N_9574,N_9642);
nand U10347 (N_10347,N_9804,N_9570);
nor U10348 (N_10348,N_9820,N_9596);
nor U10349 (N_10349,N_9542,N_9806);
and U10350 (N_10350,N_9562,N_9945);
or U10351 (N_10351,N_9684,N_9658);
or U10352 (N_10352,N_9651,N_9606);
xor U10353 (N_10353,N_9536,N_9754);
xnor U10354 (N_10354,N_9969,N_9608);
and U10355 (N_10355,N_9563,N_9603);
and U10356 (N_10356,N_9818,N_9888);
nor U10357 (N_10357,N_9690,N_9971);
xor U10358 (N_10358,N_9908,N_9655);
nor U10359 (N_10359,N_9811,N_9522);
or U10360 (N_10360,N_9784,N_9749);
and U10361 (N_10361,N_9853,N_9696);
xor U10362 (N_10362,N_9663,N_9812);
nor U10363 (N_10363,N_9855,N_9871);
or U10364 (N_10364,N_9664,N_9560);
xnor U10365 (N_10365,N_9646,N_9675);
or U10366 (N_10366,N_9844,N_9852);
xor U10367 (N_10367,N_9757,N_9805);
and U10368 (N_10368,N_9888,N_9504);
and U10369 (N_10369,N_9667,N_9712);
nand U10370 (N_10370,N_9736,N_9679);
or U10371 (N_10371,N_9831,N_9952);
or U10372 (N_10372,N_9947,N_9765);
nor U10373 (N_10373,N_9816,N_9622);
or U10374 (N_10374,N_9716,N_9732);
nor U10375 (N_10375,N_9701,N_9957);
xor U10376 (N_10376,N_9982,N_9876);
or U10377 (N_10377,N_9945,N_9750);
xnor U10378 (N_10378,N_9639,N_9543);
nor U10379 (N_10379,N_9975,N_9588);
nand U10380 (N_10380,N_9910,N_9907);
or U10381 (N_10381,N_9917,N_9948);
nor U10382 (N_10382,N_9676,N_9959);
nor U10383 (N_10383,N_9949,N_9858);
or U10384 (N_10384,N_9660,N_9510);
and U10385 (N_10385,N_9737,N_9740);
xor U10386 (N_10386,N_9916,N_9685);
or U10387 (N_10387,N_9979,N_9732);
nor U10388 (N_10388,N_9681,N_9641);
and U10389 (N_10389,N_9690,N_9659);
nor U10390 (N_10390,N_9656,N_9529);
and U10391 (N_10391,N_9972,N_9534);
xnor U10392 (N_10392,N_9591,N_9748);
xnor U10393 (N_10393,N_9535,N_9675);
nor U10394 (N_10394,N_9797,N_9682);
nand U10395 (N_10395,N_9750,N_9511);
xor U10396 (N_10396,N_9865,N_9521);
xnor U10397 (N_10397,N_9990,N_9745);
xnor U10398 (N_10398,N_9953,N_9642);
nand U10399 (N_10399,N_9752,N_9637);
nor U10400 (N_10400,N_9505,N_9866);
and U10401 (N_10401,N_9812,N_9542);
and U10402 (N_10402,N_9682,N_9512);
nand U10403 (N_10403,N_9725,N_9523);
nor U10404 (N_10404,N_9918,N_9832);
or U10405 (N_10405,N_9971,N_9591);
and U10406 (N_10406,N_9639,N_9506);
or U10407 (N_10407,N_9861,N_9915);
nor U10408 (N_10408,N_9903,N_9721);
nor U10409 (N_10409,N_9536,N_9985);
and U10410 (N_10410,N_9626,N_9534);
nor U10411 (N_10411,N_9931,N_9746);
nand U10412 (N_10412,N_9998,N_9806);
or U10413 (N_10413,N_9666,N_9511);
and U10414 (N_10414,N_9795,N_9761);
nand U10415 (N_10415,N_9893,N_9750);
nor U10416 (N_10416,N_9842,N_9923);
nand U10417 (N_10417,N_9916,N_9755);
or U10418 (N_10418,N_9696,N_9678);
nand U10419 (N_10419,N_9521,N_9597);
nand U10420 (N_10420,N_9796,N_9798);
and U10421 (N_10421,N_9954,N_9596);
nand U10422 (N_10422,N_9507,N_9637);
or U10423 (N_10423,N_9754,N_9982);
or U10424 (N_10424,N_9778,N_9796);
and U10425 (N_10425,N_9828,N_9891);
or U10426 (N_10426,N_9687,N_9902);
nand U10427 (N_10427,N_9933,N_9640);
nor U10428 (N_10428,N_9606,N_9602);
xnor U10429 (N_10429,N_9846,N_9921);
xnor U10430 (N_10430,N_9730,N_9688);
xor U10431 (N_10431,N_9551,N_9961);
xor U10432 (N_10432,N_9562,N_9593);
or U10433 (N_10433,N_9505,N_9864);
nand U10434 (N_10434,N_9595,N_9592);
nor U10435 (N_10435,N_9732,N_9766);
xor U10436 (N_10436,N_9547,N_9835);
xor U10437 (N_10437,N_9998,N_9648);
xnor U10438 (N_10438,N_9707,N_9881);
and U10439 (N_10439,N_9557,N_9509);
nand U10440 (N_10440,N_9611,N_9622);
xnor U10441 (N_10441,N_9981,N_9668);
or U10442 (N_10442,N_9558,N_9717);
and U10443 (N_10443,N_9956,N_9875);
nand U10444 (N_10444,N_9813,N_9553);
or U10445 (N_10445,N_9815,N_9555);
and U10446 (N_10446,N_9558,N_9673);
and U10447 (N_10447,N_9637,N_9511);
and U10448 (N_10448,N_9710,N_9593);
nand U10449 (N_10449,N_9713,N_9849);
nor U10450 (N_10450,N_9617,N_9554);
or U10451 (N_10451,N_9874,N_9759);
xnor U10452 (N_10452,N_9938,N_9606);
xor U10453 (N_10453,N_9825,N_9968);
and U10454 (N_10454,N_9867,N_9821);
xor U10455 (N_10455,N_9908,N_9587);
or U10456 (N_10456,N_9856,N_9745);
xor U10457 (N_10457,N_9972,N_9992);
nand U10458 (N_10458,N_9562,N_9698);
nor U10459 (N_10459,N_9740,N_9775);
and U10460 (N_10460,N_9555,N_9749);
and U10461 (N_10461,N_9746,N_9723);
or U10462 (N_10462,N_9984,N_9530);
and U10463 (N_10463,N_9805,N_9968);
nor U10464 (N_10464,N_9794,N_9708);
or U10465 (N_10465,N_9606,N_9751);
or U10466 (N_10466,N_9700,N_9630);
nor U10467 (N_10467,N_9879,N_9659);
or U10468 (N_10468,N_9731,N_9820);
nor U10469 (N_10469,N_9650,N_9669);
or U10470 (N_10470,N_9897,N_9646);
nand U10471 (N_10471,N_9909,N_9705);
nor U10472 (N_10472,N_9572,N_9563);
nand U10473 (N_10473,N_9794,N_9838);
nand U10474 (N_10474,N_9747,N_9913);
nor U10475 (N_10475,N_9723,N_9958);
and U10476 (N_10476,N_9916,N_9894);
or U10477 (N_10477,N_9613,N_9846);
xor U10478 (N_10478,N_9629,N_9810);
xnor U10479 (N_10479,N_9713,N_9573);
xnor U10480 (N_10480,N_9885,N_9874);
nand U10481 (N_10481,N_9517,N_9893);
nand U10482 (N_10482,N_9820,N_9546);
xor U10483 (N_10483,N_9500,N_9689);
nand U10484 (N_10484,N_9848,N_9602);
or U10485 (N_10485,N_9620,N_9985);
nor U10486 (N_10486,N_9702,N_9618);
nand U10487 (N_10487,N_9852,N_9826);
nand U10488 (N_10488,N_9724,N_9928);
and U10489 (N_10489,N_9974,N_9566);
xor U10490 (N_10490,N_9794,N_9601);
nor U10491 (N_10491,N_9951,N_9921);
and U10492 (N_10492,N_9992,N_9667);
and U10493 (N_10493,N_9610,N_9526);
xnor U10494 (N_10494,N_9504,N_9526);
nand U10495 (N_10495,N_9708,N_9788);
nand U10496 (N_10496,N_9990,N_9624);
or U10497 (N_10497,N_9964,N_9872);
and U10498 (N_10498,N_9788,N_9958);
xnor U10499 (N_10499,N_9809,N_9891);
nor U10500 (N_10500,N_10009,N_10440);
or U10501 (N_10501,N_10479,N_10451);
xor U10502 (N_10502,N_10228,N_10028);
xnor U10503 (N_10503,N_10220,N_10326);
nor U10504 (N_10504,N_10386,N_10454);
and U10505 (N_10505,N_10329,N_10414);
or U10506 (N_10506,N_10060,N_10472);
nor U10507 (N_10507,N_10116,N_10047);
or U10508 (N_10508,N_10018,N_10283);
and U10509 (N_10509,N_10193,N_10237);
nor U10510 (N_10510,N_10302,N_10195);
and U10511 (N_10511,N_10126,N_10477);
nand U10512 (N_10512,N_10172,N_10474);
and U10513 (N_10513,N_10258,N_10410);
nand U10514 (N_10514,N_10269,N_10233);
or U10515 (N_10515,N_10354,N_10282);
nand U10516 (N_10516,N_10373,N_10345);
and U10517 (N_10517,N_10475,N_10162);
and U10518 (N_10518,N_10291,N_10095);
nor U10519 (N_10519,N_10311,N_10024);
nor U10520 (N_10520,N_10064,N_10249);
and U10521 (N_10521,N_10308,N_10005);
nand U10522 (N_10522,N_10498,N_10313);
and U10523 (N_10523,N_10418,N_10052);
and U10524 (N_10524,N_10265,N_10154);
and U10525 (N_10525,N_10156,N_10389);
or U10526 (N_10526,N_10148,N_10099);
and U10527 (N_10527,N_10203,N_10341);
xnor U10528 (N_10528,N_10388,N_10076);
xor U10529 (N_10529,N_10419,N_10007);
nand U10530 (N_10530,N_10387,N_10381);
nand U10531 (N_10531,N_10279,N_10407);
and U10532 (N_10532,N_10369,N_10000);
nand U10533 (N_10533,N_10039,N_10245);
nand U10534 (N_10534,N_10190,N_10216);
nand U10535 (N_10535,N_10392,N_10281);
xor U10536 (N_10536,N_10048,N_10417);
or U10537 (N_10537,N_10432,N_10171);
or U10538 (N_10538,N_10010,N_10358);
and U10539 (N_10539,N_10086,N_10301);
or U10540 (N_10540,N_10334,N_10306);
xnor U10541 (N_10541,N_10114,N_10055);
xnor U10542 (N_10542,N_10470,N_10316);
nand U10543 (N_10543,N_10385,N_10490);
and U10544 (N_10544,N_10176,N_10123);
xnor U10545 (N_10545,N_10458,N_10088);
or U10546 (N_10546,N_10420,N_10017);
xor U10547 (N_10547,N_10207,N_10166);
and U10548 (N_10548,N_10142,N_10063);
nor U10549 (N_10549,N_10314,N_10330);
or U10550 (N_10550,N_10307,N_10038);
xnor U10551 (N_10551,N_10137,N_10140);
or U10552 (N_10552,N_10217,N_10328);
xor U10553 (N_10553,N_10486,N_10080);
and U10554 (N_10554,N_10270,N_10436);
or U10555 (N_10555,N_10160,N_10003);
nor U10556 (N_10556,N_10247,N_10011);
or U10557 (N_10557,N_10037,N_10045);
or U10558 (N_10558,N_10315,N_10438);
nor U10559 (N_10559,N_10318,N_10101);
and U10560 (N_10560,N_10327,N_10285);
or U10561 (N_10561,N_10084,N_10209);
or U10562 (N_10562,N_10189,N_10421);
xor U10563 (N_10563,N_10180,N_10351);
xnor U10564 (N_10564,N_10393,N_10029);
or U10565 (N_10565,N_10428,N_10023);
and U10566 (N_10566,N_10336,N_10104);
xor U10567 (N_10567,N_10259,N_10437);
or U10568 (N_10568,N_10449,N_10286);
xor U10569 (N_10569,N_10157,N_10444);
nand U10570 (N_10570,N_10187,N_10107);
nor U10571 (N_10571,N_10134,N_10181);
or U10572 (N_10572,N_10168,N_10067);
xor U10573 (N_10573,N_10248,N_10208);
xnor U10574 (N_10574,N_10355,N_10268);
and U10575 (N_10575,N_10066,N_10004);
nor U10576 (N_10576,N_10464,N_10339);
xor U10577 (N_10577,N_10078,N_10319);
xor U10578 (N_10578,N_10484,N_10002);
xor U10579 (N_10579,N_10225,N_10243);
and U10580 (N_10580,N_10359,N_10499);
or U10581 (N_10581,N_10117,N_10348);
nor U10582 (N_10582,N_10174,N_10109);
nor U10583 (N_10583,N_10020,N_10427);
or U10584 (N_10584,N_10442,N_10439);
or U10585 (N_10585,N_10443,N_10495);
or U10586 (N_10586,N_10033,N_10324);
nor U10587 (N_10587,N_10303,N_10273);
or U10588 (N_10588,N_10058,N_10403);
or U10589 (N_10589,N_10229,N_10362);
xor U10590 (N_10590,N_10480,N_10197);
nor U10591 (N_10591,N_10448,N_10103);
nor U10592 (N_10592,N_10274,N_10275);
xor U10593 (N_10593,N_10147,N_10072);
nand U10594 (N_10594,N_10264,N_10185);
and U10595 (N_10595,N_10041,N_10360);
nor U10596 (N_10596,N_10413,N_10133);
and U10597 (N_10597,N_10074,N_10129);
nor U10598 (N_10598,N_10416,N_10347);
nor U10599 (N_10599,N_10459,N_10277);
nor U10600 (N_10600,N_10353,N_10158);
nor U10601 (N_10601,N_10222,N_10138);
and U10602 (N_10602,N_10150,N_10092);
and U10603 (N_10603,N_10040,N_10292);
or U10604 (N_10604,N_10320,N_10256);
nand U10605 (N_10605,N_10165,N_10212);
and U10606 (N_10606,N_10423,N_10065);
or U10607 (N_10607,N_10143,N_10136);
nor U10608 (N_10608,N_10124,N_10473);
xor U10609 (N_10609,N_10276,N_10435);
nand U10610 (N_10610,N_10272,N_10120);
and U10611 (N_10611,N_10068,N_10404);
nand U10612 (N_10612,N_10030,N_10422);
nand U10613 (N_10613,N_10186,N_10219);
and U10614 (N_10614,N_10118,N_10132);
and U10615 (N_10615,N_10238,N_10170);
nand U10616 (N_10616,N_10242,N_10332);
and U10617 (N_10617,N_10194,N_10322);
nand U10618 (N_10618,N_10461,N_10411);
nor U10619 (N_10619,N_10481,N_10201);
xnor U10620 (N_10620,N_10361,N_10253);
nor U10621 (N_10621,N_10412,N_10398);
xor U10622 (N_10622,N_10091,N_10331);
xnor U10623 (N_10623,N_10462,N_10382);
nand U10624 (N_10624,N_10075,N_10415);
xnor U10625 (N_10625,N_10497,N_10034);
and U10626 (N_10626,N_10478,N_10297);
nand U10627 (N_10627,N_10085,N_10325);
xnor U10628 (N_10628,N_10183,N_10251);
or U10629 (N_10629,N_10450,N_10049);
nand U10630 (N_10630,N_10062,N_10053);
nand U10631 (N_10631,N_10016,N_10298);
and U10632 (N_10632,N_10399,N_10081);
xor U10633 (N_10633,N_10246,N_10070);
or U10634 (N_10634,N_10232,N_10340);
or U10635 (N_10635,N_10487,N_10130);
nand U10636 (N_10636,N_10200,N_10210);
nand U10637 (N_10637,N_10184,N_10321);
xnor U10638 (N_10638,N_10447,N_10098);
nand U10639 (N_10639,N_10240,N_10202);
xnor U10640 (N_10640,N_10239,N_10278);
nand U10641 (N_10641,N_10296,N_10192);
and U10642 (N_10642,N_10406,N_10198);
nor U10643 (N_10643,N_10375,N_10234);
nand U10644 (N_10644,N_10342,N_10008);
xnor U10645 (N_10645,N_10384,N_10352);
nand U10646 (N_10646,N_10395,N_10289);
nor U10647 (N_10647,N_10012,N_10214);
xnor U10648 (N_10648,N_10021,N_10350);
and U10649 (N_10649,N_10469,N_10257);
or U10650 (N_10650,N_10346,N_10042);
nand U10651 (N_10651,N_10400,N_10155);
nor U10652 (N_10652,N_10044,N_10367);
xor U10653 (N_10653,N_10108,N_10433);
nor U10654 (N_10654,N_10266,N_10230);
or U10655 (N_10655,N_10396,N_10372);
xnor U10656 (N_10656,N_10218,N_10179);
xnor U10657 (N_10657,N_10383,N_10139);
nor U10658 (N_10658,N_10061,N_10119);
or U10659 (N_10659,N_10463,N_10241);
nor U10660 (N_10660,N_10090,N_10335);
xnor U10661 (N_10661,N_10299,N_10261);
or U10662 (N_10662,N_10429,N_10013);
and U10663 (N_10663,N_10149,N_10294);
and U10664 (N_10664,N_10161,N_10485);
xor U10665 (N_10665,N_10343,N_10226);
nor U10666 (N_10666,N_10022,N_10056);
and U10667 (N_10667,N_10169,N_10204);
xor U10668 (N_10668,N_10111,N_10051);
or U10669 (N_10669,N_10113,N_10173);
or U10670 (N_10670,N_10431,N_10188);
nor U10671 (N_10671,N_10164,N_10496);
nor U10672 (N_10672,N_10163,N_10014);
nor U10673 (N_10673,N_10227,N_10492);
or U10674 (N_10674,N_10380,N_10153);
xnor U10675 (N_10675,N_10363,N_10223);
or U10676 (N_10676,N_10280,N_10083);
nand U10677 (N_10677,N_10096,N_10378);
nand U10678 (N_10678,N_10178,N_10488);
and U10679 (N_10679,N_10263,N_10466);
and U10680 (N_10680,N_10252,N_10110);
nand U10681 (N_10681,N_10106,N_10368);
nand U10682 (N_10682,N_10135,N_10457);
and U10683 (N_10683,N_10043,N_10035);
nand U10684 (N_10684,N_10146,N_10323);
and U10685 (N_10685,N_10452,N_10177);
and U10686 (N_10686,N_10424,N_10267);
nor U10687 (N_10687,N_10491,N_10032);
xor U10688 (N_10688,N_10284,N_10405);
xor U10689 (N_10689,N_10196,N_10102);
and U10690 (N_10690,N_10031,N_10456);
nand U10691 (N_10691,N_10182,N_10205);
nand U10692 (N_10692,N_10131,N_10397);
nor U10693 (N_10693,N_10082,N_10036);
and U10694 (N_10694,N_10025,N_10357);
nand U10695 (N_10695,N_10377,N_10394);
nor U10696 (N_10696,N_10338,N_10206);
xnor U10697 (N_10697,N_10426,N_10374);
and U10698 (N_10698,N_10305,N_10376);
xnor U10699 (N_10699,N_10244,N_10441);
nor U10700 (N_10700,N_10309,N_10356);
nand U10701 (N_10701,N_10015,N_10271);
or U10702 (N_10702,N_10460,N_10401);
nor U10703 (N_10703,N_10494,N_10050);
and U10704 (N_10704,N_10125,N_10402);
and U10705 (N_10705,N_10391,N_10287);
nand U10706 (N_10706,N_10151,N_10434);
nand U10707 (N_10707,N_10260,N_10288);
nand U10708 (N_10708,N_10145,N_10476);
nand U10709 (N_10709,N_10054,N_10310);
and U10710 (N_10710,N_10141,N_10115);
nand U10711 (N_10711,N_10026,N_10027);
or U10712 (N_10712,N_10167,N_10471);
or U10713 (N_10713,N_10019,N_10364);
xnor U10714 (N_10714,N_10489,N_10100);
and U10715 (N_10715,N_10191,N_10337);
xor U10716 (N_10716,N_10453,N_10093);
and U10717 (N_10717,N_10071,N_10371);
xor U10718 (N_10718,N_10366,N_10493);
or U10719 (N_10719,N_10379,N_10231);
or U10720 (N_10720,N_10122,N_10094);
xor U10721 (N_10721,N_10255,N_10112);
or U10722 (N_10722,N_10317,N_10455);
and U10723 (N_10723,N_10224,N_10215);
and U10724 (N_10724,N_10069,N_10059);
and U10725 (N_10725,N_10300,N_10057);
nand U10726 (N_10726,N_10121,N_10089);
nor U10727 (N_10727,N_10312,N_10482);
xnor U10728 (N_10728,N_10127,N_10046);
xor U10729 (N_10729,N_10333,N_10097);
or U10730 (N_10730,N_10001,N_10077);
nor U10731 (N_10731,N_10425,N_10152);
nor U10732 (N_10732,N_10370,N_10235);
and U10733 (N_10733,N_10211,N_10390);
and U10734 (N_10734,N_10465,N_10079);
nor U10735 (N_10735,N_10236,N_10446);
or U10736 (N_10736,N_10213,N_10365);
nand U10737 (N_10737,N_10467,N_10409);
or U10738 (N_10738,N_10006,N_10349);
xor U10739 (N_10739,N_10087,N_10293);
nor U10740 (N_10740,N_10408,N_10221);
and U10741 (N_10741,N_10254,N_10159);
xnor U10742 (N_10742,N_10250,N_10199);
xor U10743 (N_10743,N_10468,N_10290);
and U10744 (N_10744,N_10295,N_10430);
nand U10745 (N_10745,N_10128,N_10344);
nor U10746 (N_10746,N_10262,N_10144);
or U10747 (N_10747,N_10175,N_10105);
or U10748 (N_10748,N_10073,N_10483);
nor U10749 (N_10749,N_10445,N_10304);
nand U10750 (N_10750,N_10479,N_10375);
xor U10751 (N_10751,N_10415,N_10449);
or U10752 (N_10752,N_10204,N_10280);
nor U10753 (N_10753,N_10340,N_10371);
nor U10754 (N_10754,N_10143,N_10269);
nor U10755 (N_10755,N_10317,N_10488);
nand U10756 (N_10756,N_10432,N_10250);
and U10757 (N_10757,N_10180,N_10332);
or U10758 (N_10758,N_10037,N_10118);
nand U10759 (N_10759,N_10397,N_10292);
or U10760 (N_10760,N_10207,N_10116);
xnor U10761 (N_10761,N_10150,N_10065);
nor U10762 (N_10762,N_10436,N_10111);
nor U10763 (N_10763,N_10216,N_10273);
nor U10764 (N_10764,N_10145,N_10211);
or U10765 (N_10765,N_10083,N_10488);
xor U10766 (N_10766,N_10245,N_10355);
and U10767 (N_10767,N_10044,N_10343);
nand U10768 (N_10768,N_10196,N_10395);
nand U10769 (N_10769,N_10461,N_10496);
xnor U10770 (N_10770,N_10382,N_10142);
nor U10771 (N_10771,N_10134,N_10368);
nand U10772 (N_10772,N_10312,N_10461);
nand U10773 (N_10773,N_10432,N_10310);
and U10774 (N_10774,N_10209,N_10011);
or U10775 (N_10775,N_10046,N_10291);
or U10776 (N_10776,N_10228,N_10070);
nor U10777 (N_10777,N_10136,N_10173);
or U10778 (N_10778,N_10379,N_10328);
xor U10779 (N_10779,N_10054,N_10066);
nor U10780 (N_10780,N_10250,N_10075);
or U10781 (N_10781,N_10234,N_10226);
and U10782 (N_10782,N_10442,N_10207);
xor U10783 (N_10783,N_10083,N_10039);
and U10784 (N_10784,N_10421,N_10060);
xnor U10785 (N_10785,N_10158,N_10460);
and U10786 (N_10786,N_10424,N_10203);
or U10787 (N_10787,N_10027,N_10275);
or U10788 (N_10788,N_10201,N_10108);
or U10789 (N_10789,N_10409,N_10359);
or U10790 (N_10790,N_10395,N_10254);
nand U10791 (N_10791,N_10088,N_10187);
or U10792 (N_10792,N_10494,N_10187);
or U10793 (N_10793,N_10453,N_10334);
nor U10794 (N_10794,N_10234,N_10277);
or U10795 (N_10795,N_10233,N_10234);
and U10796 (N_10796,N_10401,N_10366);
or U10797 (N_10797,N_10239,N_10061);
nor U10798 (N_10798,N_10162,N_10006);
or U10799 (N_10799,N_10394,N_10354);
xnor U10800 (N_10800,N_10312,N_10328);
nand U10801 (N_10801,N_10138,N_10350);
and U10802 (N_10802,N_10496,N_10350);
or U10803 (N_10803,N_10107,N_10334);
nand U10804 (N_10804,N_10296,N_10425);
nand U10805 (N_10805,N_10010,N_10287);
nand U10806 (N_10806,N_10237,N_10342);
and U10807 (N_10807,N_10353,N_10333);
xnor U10808 (N_10808,N_10203,N_10174);
nand U10809 (N_10809,N_10372,N_10105);
or U10810 (N_10810,N_10373,N_10447);
and U10811 (N_10811,N_10425,N_10102);
nor U10812 (N_10812,N_10083,N_10391);
nand U10813 (N_10813,N_10315,N_10115);
nor U10814 (N_10814,N_10109,N_10094);
nor U10815 (N_10815,N_10401,N_10321);
and U10816 (N_10816,N_10449,N_10224);
nor U10817 (N_10817,N_10267,N_10085);
and U10818 (N_10818,N_10490,N_10110);
nor U10819 (N_10819,N_10128,N_10175);
and U10820 (N_10820,N_10444,N_10065);
and U10821 (N_10821,N_10197,N_10312);
xor U10822 (N_10822,N_10322,N_10223);
nor U10823 (N_10823,N_10222,N_10353);
or U10824 (N_10824,N_10203,N_10089);
xnor U10825 (N_10825,N_10230,N_10423);
xor U10826 (N_10826,N_10465,N_10341);
and U10827 (N_10827,N_10076,N_10210);
and U10828 (N_10828,N_10246,N_10153);
nor U10829 (N_10829,N_10311,N_10225);
nand U10830 (N_10830,N_10109,N_10414);
or U10831 (N_10831,N_10399,N_10333);
and U10832 (N_10832,N_10440,N_10085);
or U10833 (N_10833,N_10100,N_10391);
or U10834 (N_10834,N_10154,N_10023);
and U10835 (N_10835,N_10435,N_10210);
and U10836 (N_10836,N_10362,N_10275);
and U10837 (N_10837,N_10244,N_10385);
nand U10838 (N_10838,N_10271,N_10481);
nor U10839 (N_10839,N_10068,N_10047);
and U10840 (N_10840,N_10448,N_10178);
nand U10841 (N_10841,N_10090,N_10034);
or U10842 (N_10842,N_10138,N_10148);
nand U10843 (N_10843,N_10030,N_10185);
and U10844 (N_10844,N_10016,N_10182);
and U10845 (N_10845,N_10060,N_10231);
or U10846 (N_10846,N_10093,N_10214);
nor U10847 (N_10847,N_10357,N_10403);
or U10848 (N_10848,N_10256,N_10212);
xnor U10849 (N_10849,N_10233,N_10134);
nand U10850 (N_10850,N_10053,N_10138);
xor U10851 (N_10851,N_10439,N_10152);
or U10852 (N_10852,N_10013,N_10198);
and U10853 (N_10853,N_10329,N_10365);
or U10854 (N_10854,N_10235,N_10070);
and U10855 (N_10855,N_10288,N_10439);
xnor U10856 (N_10856,N_10020,N_10054);
nand U10857 (N_10857,N_10022,N_10137);
and U10858 (N_10858,N_10158,N_10331);
nand U10859 (N_10859,N_10343,N_10200);
or U10860 (N_10860,N_10437,N_10227);
and U10861 (N_10861,N_10332,N_10192);
xor U10862 (N_10862,N_10359,N_10052);
and U10863 (N_10863,N_10263,N_10371);
or U10864 (N_10864,N_10253,N_10098);
nor U10865 (N_10865,N_10446,N_10016);
or U10866 (N_10866,N_10169,N_10081);
nand U10867 (N_10867,N_10350,N_10493);
and U10868 (N_10868,N_10086,N_10410);
or U10869 (N_10869,N_10226,N_10071);
xor U10870 (N_10870,N_10068,N_10044);
or U10871 (N_10871,N_10450,N_10323);
nand U10872 (N_10872,N_10383,N_10259);
xor U10873 (N_10873,N_10476,N_10274);
nand U10874 (N_10874,N_10227,N_10427);
xor U10875 (N_10875,N_10434,N_10106);
xor U10876 (N_10876,N_10189,N_10474);
or U10877 (N_10877,N_10118,N_10179);
or U10878 (N_10878,N_10105,N_10486);
and U10879 (N_10879,N_10294,N_10327);
nor U10880 (N_10880,N_10179,N_10481);
and U10881 (N_10881,N_10497,N_10457);
nand U10882 (N_10882,N_10176,N_10367);
or U10883 (N_10883,N_10367,N_10324);
nand U10884 (N_10884,N_10044,N_10436);
and U10885 (N_10885,N_10453,N_10441);
nand U10886 (N_10886,N_10485,N_10120);
nand U10887 (N_10887,N_10072,N_10293);
xor U10888 (N_10888,N_10237,N_10398);
and U10889 (N_10889,N_10347,N_10266);
nor U10890 (N_10890,N_10027,N_10404);
nand U10891 (N_10891,N_10140,N_10079);
nor U10892 (N_10892,N_10081,N_10109);
or U10893 (N_10893,N_10298,N_10398);
nand U10894 (N_10894,N_10320,N_10277);
or U10895 (N_10895,N_10018,N_10416);
or U10896 (N_10896,N_10487,N_10458);
and U10897 (N_10897,N_10129,N_10369);
or U10898 (N_10898,N_10222,N_10248);
nor U10899 (N_10899,N_10300,N_10475);
or U10900 (N_10900,N_10461,N_10395);
or U10901 (N_10901,N_10104,N_10313);
xnor U10902 (N_10902,N_10009,N_10370);
and U10903 (N_10903,N_10126,N_10301);
or U10904 (N_10904,N_10307,N_10316);
xor U10905 (N_10905,N_10136,N_10315);
and U10906 (N_10906,N_10402,N_10007);
or U10907 (N_10907,N_10293,N_10261);
xnor U10908 (N_10908,N_10229,N_10406);
nand U10909 (N_10909,N_10111,N_10287);
nor U10910 (N_10910,N_10107,N_10194);
nor U10911 (N_10911,N_10488,N_10253);
xnor U10912 (N_10912,N_10293,N_10190);
nand U10913 (N_10913,N_10082,N_10077);
nand U10914 (N_10914,N_10200,N_10081);
nor U10915 (N_10915,N_10346,N_10073);
nor U10916 (N_10916,N_10393,N_10232);
and U10917 (N_10917,N_10302,N_10379);
nand U10918 (N_10918,N_10282,N_10409);
xnor U10919 (N_10919,N_10090,N_10136);
nor U10920 (N_10920,N_10425,N_10219);
and U10921 (N_10921,N_10124,N_10223);
or U10922 (N_10922,N_10129,N_10191);
or U10923 (N_10923,N_10103,N_10207);
or U10924 (N_10924,N_10032,N_10144);
nand U10925 (N_10925,N_10340,N_10217);
nand U10926 (N_10926,N_10098,N_10292);
and U10927 (N_10927,N_10465,N_10116);
nor U10928 (N_10928,N_10291,N_10128);
nor U10929 (N_10929,N_10079,N_10201);
or U10930 (N_10930,N_10329,N_10154);
nand U10931 (N_10931,N_10197,N_10233);
and U10932 (N_10932,N_10108,N_10109);
xnor U10933 (N_10933,N_10275,N_10346);
xnor U10934 (N_10934,N_10009,N_10394);
nand U10935 (N_10935,N_10156,N_10238);
xor U10936 (N_10936,N_10334,N_10168);
and U10937 (N_10937,N_10497,N_10379);
xnor U10938 (N_10938,N_10350,N_10087);
xnor U10939 (N_10939,N_10043,N_10030);
or U10940 (N_10940,N_10412,N_10434);
nand U10941 (N_10941,N_10021,N_10096);
nand U10942 (N_10942,N_10239,N_10421);
and U10943 (N_10943,N_10218,N_10467);
or U10944 (N_10944,N_10345,N_10034);
nand U10945 (N_10945,N_10320,N_10217);
xnor U10946 (N_10946,N_10214,N_10294);
nor U10947 (N_10947,N_10179,N_10419);
nand U10948 (N_10948,N_10061,N_10271);
and U10949 (N_10949,N_10092,N_10444);
nand U10950 (N_10950,N_10323,N_10463);
or U10951 (N_10951,N_10451,N_10338);
xor U10952 (N_10952,N_10256,N_10209);
and U10953 (N_10953,N_10252,N_10463);
xnor U10954 (N_10954,N_10230,N_10246);
nor U10955 (N_10955,N_10211,N_10188);
xnor U10956 (N_10956,N_10492,N_10062);
nand U10957 (N_10957,N_10245,N_10226);
nor U10958 (N_10958,N_10210,N_10066);
xnor U10959 (N_10959,N_10414,N_10083);
and U10960 (N_10960,N_10207,N_10094);
nor U10961 (N_10961,N_10372,N_10374);
xnor U10962 (N_10962,N_10325,N_10205);
or U10963 (N_10963,N_10458,N_10405);
nand U10964 (N_10964,N_10248,N_10327);
or U10965 (N_10965,N_10368,N_10157);
or U10966 (N_10966,N_10123,N_10189);
nand U10967 (N_10967,N_10156,N_10050);
nand U10968 (N_10968,N_10072,N_10093);
nand U10969 (N_10969,N_10460,N_10123);
nor U10970 (N_10970,N_10065,N_10028);
and U10971 (N_10971,N_10163,N_10053);
or U10972 (N_10972,N_10308,N_10079);
or U10973 (N_10973,N_10110,N_10489);
and U10974 (N_10974,N_10163,N_10079);
nor U10975 (N_10975,N_10305,N_10140);
and U10976 (N_10976,N_10225,N_10222);
or U10977 (N_10977,N_10373,N_10476);
and U10978 (N_10978,N_10058,N_10063);
and U10979 (N_10979,N_10186,N_10426);
and U10980 (N_10980,N_10130,N_10461);
nor U10981 (N_10981,N_10022,N_10129);
or U10982 (N_10982,N_10127,N_10495);
and U10983 (N_10983,N_10219,N_10204);
xnor U10984 (N_10984,N_10099,N_10000);
nor U10985 (N_10985,N_10299,N_10157);
or U10986 (N_10986,N_10254,N_10170);
and U10987 (N_10987,N_10113,N_10039);
and U10988 (N_10988,N_10292,N_10214);
or U10989 (N_10989,N_10253,N_10365);
nand U10990 (N_10990,N_10414,N_10333);
xor U10991 (N_10991,N_10460,N_10044);
nand U10992 (N_10992,N_10010,N_10226);
or U10993 (N_10993,N_10324,N_10050);
xor U10994 (N_10994,N_10026,N_10135);
nand U10995 (N_10995,N_10202,N_10348);
nand U10996 (N_10996,N_10366,N_10138);
nand U10997 (N_10997,N_10474,N_10371);
or U10998 (N_10998,N_10040,N_10143);
xor U10999 (N_10999,N_10083,N_10035);
xnor U11000 (N_11000,N_10609,N_10544);
and U11001 (N_11001,N_10515,N_10600);
nor U11002 (N_11002,N_10931,N_10894);
nor U11003 (N_11003,N_10620,N_10511);
or U11004 (N_11004,N_10656,N_10698);
nor U11005 (N_11005,N_10845,N_10781);
nor U11006 (N_11006,N_10624,N_10526);
or U11007 (N_11007,N_10783,N_10696);
nand U11008 (N_11008,N_10785,N_10717);
nor U11009 (N_11009,N_10939,N_10922);
and U11010 (N_11010,N_10854,N_10720);
nand U11011 (N_11011,N_10837,N_10541);
nand U11012 (N_11012,N_10725,N_10738);
and U11013 (N_11013,N_10617,N_10693);
and U11014 (N_11014,N_10942,N_10893);
nand U11015 (N_11015,N_10743,N_10974);
nor U11016 (N_11016,N_10771,N_10571);
xor U11017 (N_11017,N_10561,N_10679);
nand U11018 (N_11018,N_10817,N_10851);
xor U11019 (N_11019,N_10648,N_10749);
nand U11020 (N_11020,N_10674,N_10754);
and U11021 (N_11021,N_10706,N_10638);
or U11022 (N_11022,N_10584,N_10869);
xnor U11023 (N_11023,N_10635,N_10521);
xor U11024 (N_11024,N_10784,N_10677);
nand U11025 (N_11025,N_10752,N_10760);
and U11026 (N_11026,N_10726,N_10659);
or U11027 (N_11027,N_10588,N_10671);
nor U11028 (N_11028,N_10778,N_10923);
or U11029 (N_11029,N_10788,N_10681);
nor U11030 (N_11030,N_10512,N_10753);
nand U11031 (N_11031,N_10791,N_10715);
nand U11032 (N_11032,N_10578,N_10814);
xor U11033 (N_11033,N_10826,N_10874);
or U11034 (N_11034,N_10809,N_10933);
xnor U11035 (N_11035,N_10920,N_10736);
or U11036 (N_11036,N_10870,N_10686);
xor U11037 (N_11037,N_10790,N_10574);
or U11038 (N_11038,N_10524,N_10573);
and U11039 (N_11039,N_10858,N_10957);
and U11040 (N_11040,N_10700,N_10821);
nand U11041 (N_11041,N_10848,N_10678);
nor U11042 (N_11042,N_10560,N_10820);
xor U11043 (N_11043,N_10844,N_10927);
nor U11044 (N_11044,N_10872,N_10775);
xnor U11045 (N_11045,N_10567,N_10772);
and U11046 (N_11046,N_10881,N_10580);
xor U11047 (N_11047,N_10501,N_10506);
xor U11048 (N_11048,N_10568,N_10780);
and U11049 (N_11049,N_10628,N_10908);
and U11050 (N_11050,N_10786,N_10694);
or U11051 (N_11051,N_10513,N_10988);
and U11052 (N_11052,N_10547,N_10570);
and U11053 (N_11053,N_10831,N_10660);
or U11054 (N_11054,N_10556,N_10919);
or U11055 (N_11055,N_10504,N_10950);
or U11056 (N_11056,N_10773,N_10517);
nand U11057 (N_11057,N_10808,N_10711);
nand U11058 (N_11058,N_10618,N_10910);
xnor U11059 (N_11059,N_10739,N_10546);
and U11060 (N_11060,N_10956,N_10868);
and U11061 (N_11061,N_10586,N_10543);
or U11062 (N_11062,N_10719,N_10582);
and U11063 (N_11063,N_10946,N_10597);
xor U11064 (N_11064,N_10748,N_10747);
and U11065 (N_11065,N_10902,N_10776);
nor U11066 (N_11066,N_10834,N_10598);
xnor U11067 (N_11067,N_10904,N_10667);
nor U11068 (N_11068,N_10647,N_10687);
and U11069 (N_11069,N_10959,N_10839);
nand U11070 (N_11070,N_10983,N_10683);
and U11071 (N_11071,N_10998,N_10856);
xor U11072 (N_11072,N_10928,N_10827);
or U11073 (N_11073,N_10622,N_10566);
nand U11074 (N_11074,N_10591,N_10640);
or U11075 (N_11075,N_10800,N_10766);
and U11076 (N_11076,N_10531,N_10673);
or U11077 (N_11077,N_10967,N_10563);
or U11078 (N_11078,N_10599,N_10619);
nor U11079 (N_11079,N_10581,N_10519);
nand U11080 (N_11080,N_10777,N_10680);
and U11081 (N_11081,N_10861,N_10704);
nand U11082 (N_11082,N_10740,N_10873);
and U11083 (N_11083,N_10981,N_10538);
nand U11084 (N_11084,N_10505,N_10976);
nor U11085 (N_11085,N_10921,N_10986);
and U11086 (N_11086,N_10764,N_10966);
nor U11087 (N_11087,N_10852,N_10975);
or U11088 (N_11088,N_10705,N_10987);
and U11089 (N_11089,N_10540,N_10822);
xnor U11090 (N_11090,N_10887,N_10954);
nand U11091 (N_11091,N_10840,N_10746);
nand U11092 (N_11092,N_10914,N_10813);
xor U11093 (N_11093,N_10623,N_10663);
nor U11094 (N_11094,N_10707,N_10735);
nand U11095 (N_11095,N_10758,N_10645);
and U11096 (N_11096,N_10905,N_10880);
or U11097 (N_11097,N_10862,N_10810);
or U11098 (N_11098,N_10968,N_10787);
nor U11099 (N_11099,N_10551,N_10589);
nor U11100 (N_11100,N_10703,N_10621);
or U11101 (N_11101,N_10533,N_10690);
or U11102 (N_11102,N_10793,N_10688);
or U11103 (N_11103,N_10575,N_10522);
nand U11104 (N_11104,N_10565,N_10516);
xor U11105 (N_11105,N_10537,N_10510);
xnor U11106 (N_11106,N_10769,N_10789);
nand U11107 (N_11107,N_10554,N_10549);
xor U11108 (N_11108,N_10828,N_10615);
nand U11109 (N_11109,N_10930,N_10532);
or U11110 (N_11110,N_10611,N_10876);
nand U11111 (N_11111,N_10508,N_10912);
nand U11112 (N_11112,N_10916,N_10523);
nor U11113 (N_11113,N_10951,N_10883);
nand U11114 (N_11114,N_10590,N_10601);
or U11115 (N_11115,N_10884,N_10545);
and U11116 (N_11116,N_10906,N_10909);
and U11117 (N_11117,N_10602,N_10889);
nand U11118 (N_11118,N_10643,N_10666);
nor U11119 (N_11119,N_10982,N_10572);
nand U11120 (N_11120,N_10610,N_10750);
and U11121 (N_11121,N_10964,N_10592);
nand U11122 (N_11122,N_10865,N_10829);
xor U11123 (N_11123,N_10913,N_10702);
and U11124 (N_11124,N_10745,N_10731);
nor U11125 (N_11125,N_10934,N_10938);
or U11126 (N_11126,N_10898,N_10596);
nand U11127 (N_11127,N_10652,N_10733);
nand U11128 (N_11128,N_10836,N_10779);
and U11129 (N_11129,N_10838,N_10960);
and U11130 (N_11130,N_10815,N_10612);
nand U11131 (N_11131,N_10585,N_10606);
and U11132 (N_11132,N_10818,N_10765);
nor U11133 (N_11133,N_10812,N_10972);
nand U11134 (N_11134,N_10634,N_10665);
and U11135 (N_11135,N_10664,N_10802);
or U11136 (N_11136,N_10729,N_10650);
nor U11137 (N_11137,N_10948,N_10973);
nor U11138 (N_11138,N_10768,N_10937);
and U11139 (N_11139,N_10734,N_10692);
and U11140 (N_11140,N_10646,N_10841);
xnor U11141 (N_11141,N_10644,N_10994);
and U11142 (N_11142,N_10708,N_10830);
or U11143 (N_11143,N_10936,N_10535);
or U11144 (N_11144,N_10722,N_10658);
and U11145 (N_11145,N_10728,N_10991);
or U11146 (N_11146,N_10641,N_10629);
xor U11147 (N_11147,N_10662,N_10875);
xnor U11148 (N_11148,N_10853,N_10528);
nand U11149 (N_11149,N_10895,N_10886);
nand U11150 (N_11150,N_10569,N_10925);
nor U11151 (N_11151,N_10855,N_10891);
and U11152 (N_11152,N_10548,N_10917);
or U11153 (N_11153,N_10847,N_10877);
nand U11154 (N_11154,N_10632,N_10672);
nor U11155 (N_11155,N_10943,N_10654);
and U11156 (N_11156,N_10761,N_10542);
and U11157 (N_11157,N_10969,N_10804);
or U11158 (N_11158,N_10605,N_10723);
nor U11159 (N_11159,N_10577,N_10929);
and U11160 (N_11160,N_10849,N_10595);
and U11161 (N_11161,N_10579,N_10944);
nor U11162 (N_11162,N_10799,N_10965);
and U11163 (N_11163,N_10907,N_10732);
nor U11164 (N_11164,N_10801,N_10651);
or U11165 (N_11165,N_10530,N_10742);
xnor U11166 (N_11166,N_10980,N_10500);
nor U11167 (N_11167,N_10721,N_10797);
or U11168 (N_11168,N_10608,N_10899);
nor U11169 (N_11169,N_10774,N_10593);
nor U11170 (N_11170,N_10824,N_10604);
nor U11171 (N_11171,N_10751,N_10724);
nand U11172 (N_11172,N_10805,N_10924);
nand U11173 (N_11173,N_10846,N_10625);
nand U11174 (N_11174,N_10529,N_10866);
nor U11175 (N_11175,N_10555,N_10709);
or U11176 (N_11176,N_10642,N_10863);
xnor U11177 (N_11177,N_10682,N_10657);
and U11178 (N_11178,N_10940,N_10962);
and U11179 (N_11179,N_10819,N_10562);
and U11180 (N_11180,N_10882,N_10900);
nand U11181 (N_11181,N_10878,N_10952);
or U11182 (N_11182,N_10903,N_10896);
xor U11183 (N_11183,N_10557,N_10999);
and U11184 (N_11184,N_10888,N_10767);
or U11185 (N_11185,N_10675,N_10859);
xor U11186 (N_11186,N_10979,N_10661);
nor U11187 (N_11187,N_10639,N_10627);
and U11188 (N_11188,N_10850,N_10718);
and U11189 (N_11189,N_10890,N_10744);
nor U11190 (N_11190,N_10860,N_10762);
nor U11191 (N_11191,N_10993,N_10713);
or U11192 (N_11192,N_10807,N_10811);
and U11193 (N_11193,N_10941,N_10502);
or U11194 (N_11194,N_10684,N_10803);
nor U11195 (N_11195,N_10915,N_10932);
nand U11196 (N_11196,N_10630,N_10564);
nor U11197 (N_11197,N_10971,N_10520);
and U11198 (N_11198,N_10782,N_10885);
xnor U11199 (N_11199,N_10918,N_10961);
and U11200 (N_11200,N_10697,N_10514);
and U11201 (N_11201,N_10871,N_10668);
xor U11202 (N_11202,N_10637,N_10816);
xnor U11203 (N_11203,N_10985,N_10757);
nand U11204 (N_11204,N_10536,N_10741);
xnor U11205 (N_11205,N_10636,N_10984);
xnor U11206 (N_11206,N_10631,N_10992);
or U11207 (N_11207,N_10559,N_10879);
xor U11208 (N_11208,N_10553,N_10716);
xor U11209 (N_11209,N_10970,N_10806);
or U11210 (N_11210,N_10633,N_10503);
nor U11211 (N_11211,N_10958,N_10892);
xnor U11212 (N_11212,N_10756,N_10963);
or U11213 (N_11213,N_10792,N_10949);
nor U11214 (N_11214,N_10653,N_10911);
or U11215 (N_11215,N_10989,N_10867);
and U11216 (N_11216,N_10935,N_10795);
nor U11217 (N_11217,N_10763,N_10507);
xnor U11218 (N_11218,N_10842,N_10897);
nand U11219 (N_11219,N_10737,N_10576);
and U11220 (N_11220,N_10710,N_10835);
xnor U11221 (N_11221,N_10945,N_10685);
xor U11222 (N_11222,N_10539,N_10518);
or U11223 (N_11223,N_10509,N_10953);
or U11224 (N_11224,N_10701,N_10655);
nand U11225 (N_11225,N_10977,N_10857);
xor U11226 (N_11226,N_10712,N_10832);
or U11227 (N_11227,N_10825,N_10759);
or U11228 (N_11228,N_10558,N_10594);
and U11229 (N_11229,N_10997,N_10699);
nand U11230 (N_11230,N_10978,N_10926);
and U11231 (N_11231,N_10607,N_10833);
or U11232 (N_11232,N_10794,N_10996);
xor U11233 (N_11233,N_10730,N_10670);
xor U11234 (N_11234,N_10864,N_10587);
or U11235 (N_11235,N_10603,N_10947);
nand U11236 (N_11236,N_10616,N_10727);
xor U11237 (N_11237,N_10676,N_10552);
and U11238 (N_11238,N_10613,N_10691);
nand U11239 (N_11239,N_10550,N_10525);
or U11240 (N_11240,N_10614,N_10534);
xor U11241 (N_11241,N_10843,N_10714);
or U11242 (N_11242,N_10990,N_10798);
xor U11243 (N_11243,N_10689,N_10755);
nand U11244 (N_11244,N_10823,N_10527);
nor U11245 (N_11245,N_10669,N_10796);
xnor U11246 (N_11246,N_10695,N_10649);
and U11247 (N_11247,N_10583,N_10995);
and U11248 (N_11248,N_10770,N_10901);
nand U11249 (N_11249,N_10955,N_10626);
nor U11250 (N_11250,N_10875,N_10850);
nor U11251 (N_11251,N_10525,N_10745);
or U11252 (N_11252,N_10910,N_10836);
nor U11253 (N_11253,N_10997,N_10612);
xor U11254 (N_11254,N_10607,N_10940);
or U11255 (N_11255,N_10533,N_10597);
nor U11256 (N_11256,N_10726,N_10602);
nand U11257 (N_11257,N_10792,N_10831);
xnor U11258 (N_11258,N_10502,N_10540);
nand U11259 (N_11259,N_10811,N_10575);
or U11260 (N_11260,N_10977,N_10551);
and U11261 (N_11261,N_10610,N_10968);
xnor U11262 (N_11262,N_10570,N_10596);
or U11263 (N_11263,N_10565,N_10776);
nor U11264 (N_11264,N_10700,N_10574);
nor U11265 (N_11265,N_10908,N_10510);
nor U11266 (N_11266,N_10600,N_10899);
nor U11267 (N_11267,N_10813,N_10812);
nand U11268 (N_11268,N_10637,N_10557);
nand U11269 (N_11269,N_10675,N_10746);
nand U11270 (N_11270,N_10838,N_10974);
or U11271 (N_11271,N_10891,N_10905);
and U11272 (N_11272,N_10922,N_10502);
and U11273 (N_11273,N_10536,N_10698);
or U11274 (N_11274,N_10604,N_10944);
or U11275 (N_11275,N_10890,N_10533);
nor U11276 (N_11276,N_10999,N_10753);
or U11277 (N_11277,N_10634,N_10835);
xor U11278 (N_11278,N_10644,N_10589);
xor U11279 (N_11279,N_10978,N_10666);
and U11280 (N_11280,N_10947,N_10901);
or U11281 (N_11281,N_10694,N_10500);
and U11282 (N_11282,N_10865,N_10924);
or U11283 (N_11283,N_10787,N_10688);
or U11284 (N_11284,N_10541,N_10719);
nand U11285 (N_11285,N_10980,N_10832);
xor U11286 (N_11286,N_10907,N_10578);
xor U11287 (N_11287,N_10827,N_10668);
xor U11288 (N_11288,N_10664,N_10740);
xor U11289 (N_11289,N_10596,N_10565);
nand U11290 (N_11290,N_10533,N_10655);
nand U11291 (N_11291,N_10591,N_10955);
and U11292 (N_11292,N_10699,N_10836);
xor U11293 (N_11293,N_10843,N_10544);
or U11294 (N_11294,N_10788,N_10706);
xnor U11295 (N_11295,N_10588,N_10653);
or U11296 (N_11296,N_10698,N_10754);
nor U11297 (N_11297,N_10772,N_10993);
and U11298 (N_11298,N_10668,N_10741);
nor U11299 (N_11299,N_10599,N_10805);
and U11300 (N_11300,N_10741,N_10755);
nor U11301 (N_11301,N_10687,N_10640);
nor U11302 (N_11302,N_10651,N_10827);
nand U11303 (N_11303,N_10872,N_10988);
xnor U11304 (N_11304,N_10769,N_10869);
xnor U11305 (N_11305,N_10688,N_10549);
or U11306 (N_11306,N_10990,N_10813);
and U11307 (N_11307,N_10767,N_10985);
and U11308 (N_11308,N_10901,N_10836);
or U11309 (N_11309,N_10943,N_10617);
and U11310 (N_11310,N_10509,N_10633);
nand U11311 (N_11311,N_10582,N_10773);
and U11312 (N_11312,N_10548,N_10984);
or U11313 (N_11313,N_10976,N_10524);
nand U11314 (N_11314,N_10588,N_10524);
or U11315 (N_11315,N_10720,N_10900);
and U11316 (N_11316,N_10643,N_10740);
nand U11317 (N_11317,N_10856,N_10905);
xor U11318 (N_11318,N_10758,N_10995);
or U11319 (N_11319,N_10900,N_10560);
xnor U11320 (N_11320,N_10987,N_10692);
xor U11321 (N_11321,N_10542,N_10773);
nand U11322 (N_11322,N_10946,N_10885);
and U11323 (N_11323,N_10856,N_10843);
xor U11324 (N_11324,N_10625,N_10859);
nor U11325 (N_11325,N_10658,N_10927);
nor U11326 (N_11326,N_10568,N_10655);
and U11327 (N_11327,N_10661,N_10671);
and U11328 (N_11328,N_10561,N_10857);
nand U11329 (N_11329,N_10982,N_10788);
xor U11330 (N_11330,N_10656,N_10757);
xnor U11331 (N_11331,N_10531,N_10600);
and U11332 (N_11332,N_10990,N_10565);
or U11333 (N_11333,N_10502,N_10648);
nor U11334 (N_11334,N_10960,N_10779);
or U11335 (N_11335,N_10803,N_10667);
or U11336 (N_11336,N_10566,N_10755);
or U11337 (N_11337,N_10725,N_10522);
and U11338 (N_11338,N_10814,N_10885);
nand U11339 (N_11339,N_10571,N_10818);
or U11340 (N_11340,N_10699,N_10735);
and U11341 (N_11341,N_10560,N_10782);
nor U11342 (N_11342,N_10585,N_10912);
and U11343 (N_11343,N_10925,N_10640);
nand U11344 (N_11344,N_10889,N_10871);
xnor U11345 (N_11345,N_10688,N_10872);
or U11346 (N_11346,N_10991,N_10987);
nor U11347 (N_11347,N_10569,N_10720);
or U11348 (N_11348,N_10802,N_10720);
and U11349 (N_11349,N_10721,N_10571);
nand U11350 (N_11350,N_10831,N_10545);
and U11351 (N_11351,N_10815,N_10743);
xor U11352 (N_11352,N_10849,N_10558);
xnor U11353 (N_11353,N_10932,N_10698);
xor U11354 (N_11354,N_10682,N_10837);
or U11355 (N_11355,N_10843,N_10508);
or U11356 (N_11356,N_10909,N_10766);
and U11357 (N_11357,N_10721,N_10836);
nor U11358 (N_11358,N_10819,N_10603);
nand U11359 (N_11359,N_10937,N_10788);
nor U11360 (N_11360,N_10976,N_10757);
and U11361 (N_11361,N_10752,N_10504);
xor U11362 (N_11362,N_10929,N_10821);
nor U11363 (N_11363,N_10860,N_10907);
xnor U11364 (N_11364,N_10753,N_10874);
xor U11365 (N_11365,N_10955,N_10779);
xnor U11366 (N_11366,N_10845,N_10512);
nand U11367 (N_11367,N_10906,N_10935);
and U11368 (N_11368,N_10685,N_10924);
nor U11369 (N_11369,N_10855,N_10567);
nand U11370 (N_11370,N_10906,N_10823);
or U11371 (N_11371,N_10718,N_10689);
xnor U11372 (N_11372,N_10749,N_10897);
xnor U11373 (N_11373,N_10876,N_10751);
nor U11374 (N_11374,N_10772,N_10832);
and U11375 (N_11375,N_10638,N_10761);
and U11376 (N_11376,N_10702,N_10997);
or U11377 (N_11377,N_10991,N_10535);
or U11378 (N_11378,N_10798,N_10841);
nor U11379 (N_11379,N_10628,N_10957);
or U11380 (N_11380,N_10524,N_10953);
nor U11381 (N_11381,N_10578,N_10921);
nor U11382 (N_11382,N_10649,N_10989);
and U11383 (N_11383,N_10645,N_10727);
and U11384 (N_11384,N_10790,N_10645);
or U11385 (N_11385,N_10552,N_10896);
nor U11386 (N_11386,N_10690,N_10620);
or U11387 (N_11387,N_10528,N_10787);
nand U11388 (N_11388,N_10667,N_10548);
nand U11389 (N_11389,N_10730,N_10777);
xnor U11390 (N_11390,N_10669,N_10526);
xnor U11391 (N_11391,N_10972,N_10751);
nor U11392 (N_11392,N_10996,N_10731);
nor U11393 (N_11393,N_10626,N_10686);
or U11394 (N_11394,N_10688,N_10888);
and U11395 (N_11395,N_10503,N_10665);
and U11396 (N_11396,N_10693,N_10788);
nor U11397 (N_11397,N_10878,N_10589);
xor U11398 (N_11398,N_10791,N_10687);
nor U11399 (N_11399,N_10735,N_10763);
or U11400 (N_11400,N_10610,N_10626);
nand U11401 (N_11401,N_10782,N_10959);
nand U11402 (N_11402,N_10868,N_10815);
or U11403 (N_11403,N_10849,N_10807);
nor U11404 (N_11404,N_10592,N_10805);
xor U11405 (N_11405,N_10881,N_10751);
and U11406 (N_11406,N_10520,N_10724);
nor U11407 (N_11407,N_10891,N_10988);
nand U11408 (N_11408,N_10724,N_10640);
or U11409 (N_11409,N_10579,N_10774);
or U11410 (N_11410,N_10919,N_10506);
xnor U11411 (N_11411,N_10567,N_10540);
xnor U11412 (N_11412,N_10652,N_10782);
nor U11413 (N_11413,N_10643,N_10817);
nand U11414 (N_11414,N_10542,N_10768);
and U11415 (N_11415,N_10741,N_10709);
nand U11416 (N_11416,N_10621,N_10624);
nand U11417 (N_11417,N_10749,N_10805);
nor U11418 (N_11418,N_10867,N_10827);
nand U11419 (N_11419,N_10934,N_10743);
and U11420 (N_11420,N_10956,N_10540);
or U11421 (N_11421,N_10978,N_10793);
nand U11422 (N_11422,N_10912,N_10804);
or U11423 (N_11423,N_10813,N_10772);
xnor U11424 (N_11424,N_10736,N_10556);
nand U11425 (N_11425,N_10872,N_10605);
nand U11426 (N_11426,N_10699,N_10639);
nor U11427 (N_11427,N_10576,N_10971);
xor U11428 (N_11428,N_10512,N_10867);
and U11429 (N_11429,N_10889,N_10778);
or U11430 (N_11430,N_10960,N_10985);
or U11431 (N_11431,N_10706,N_10765);
nor U11432 (N_11432,N_10904,N_10694);
and U11433 (N_11433,N_10994,N_10714);
nand U11434 (N_11434,N_10829,N_10979);
nand U11435 (N_11435,N_10891,N_10678);
and U11436 (N_11436,N_10605,N_10680);
and U11437 (N_11437,N_10525,N_10647);
xor U11438 (N_11438,N_10659,N_10639);
or U11439 (N_11439,N_10940,N_10578);
xor U11440 (N_11440,N_10698,N_10554);
nand U11441 (N_11441,N_10892,N_10788);
xor U11442 (N_11442,N_10733,N_10663);
nand U11443 (N_11443,N_10562,N_10966);
nor U11444 (N_11444,N_10810,N_10894);
xnor U11445 (N_11445,N_10581,N_10912);
nor U11446 (N_11446,N_10938,N_10995);
nor U11447 (N_11447,N_10755,N_10879);
or U11448 (N_11448,N_10762,N_10820);
nor U11449 (N_11449,N_10607,N_10783);
or U11450 (N_11450,N_10982,N_10667);
nand U11451 (N_11451,N_10948,N_10520);
or U11452 (N_11452,N_10716,N_10892);
or U11453 (N_11453,N_10811,N_10743);
or U11454 (N_11454,N_10830,N_10674);
and U11455 (N_11455,N_10918,N_10804);
and U11456 (N_11456,N_10859,N_10548);
nor U11457 (N_11457,N_10896,N_10572);
or U11458 (N_11458,N_10957,N_10832);
or U11459 (N_11459,N_10920,N_10799);
and U11460 (N_11460,N_10977,N_10630);
nor U11461 (N_11461,N_10797,N_10542);
xor U11462 (N_11462,N_10859,N_10543);
nand U11463 (N_11463,N_10614,N_10848);
nor U11464 (N_11464,N_10675,N_10750);
and U11465 (N_11465,N_10768,N_10817);
nor U11466 (N_11466,N_10679,N_10925);
xnor U11467 (N_11467,N_10795,N_10538);
and U11468 (N_11468,N_10521,N_10622);
xnor U11469 (N_11469,N_10738,N_10717);
xnor U11470 (N_11470,N_10933,N_10797);
or U11471 (N_11471,N_10765,N_10686);
xor U11472 (N_11472,N_10702,N_10869);
nand U11473 (N_11473,N_10772,N_10537);
nand U11474 (N_11474,N_10916,N_10601);
and U11475 (N_11475,N_10850,N_10687);
nor U11476 (N_11476,N_10609,N_10974);
nand U11477 (N_11477,N_10660,N_10908);
nor U11478 (N_11478,N_10840,N_10708);
nor U11479 (N_11479,N_10690,N_10721);
or U11480 (N_11480,N_10928,N_10546);
nor U11481 (N_11481,N_10683,N_10810);
nand U11482 (N_11482,N_10822,N_10609);
nor U11483 (N_11483,N_10745,N_10526);
nor U11484 (N_11484,N_10882,N_10863);
or U11485 (N_11485,N_10720,N_10978);
xor U11486 (N_11486,N_10710,N_10871);
nor U11487 (N_11487,N_10743,N_10729);
and U11488 (N_11488,N_10905,N_10983);
and U11489 (N_11489,N_10776,N_10731);
nand U11490 (N_11490,N_10741,N_10754);
nand U11491 (N_11491,N_10823,N_10612);
or U11492 (N_11492,N_10653,N_10606);
and U11493 (N_11493,N_10649,N_10506);
and U11494 (N_11494,N_10538,N_10885);
or U11495 (N_11495,N_10520,N_10882);
xnor U11496 (N_11496,N_10598,N_10728);
xnor U11497 (N_11497,N_10879,N_10596);
nor U11498 (N_11498,N_10777,N_10837);
or U11499 (N_11499,N_10951,N_10518);
xnor U11500 (N_11500,N_11133,N_11057);
xor U11501 (N_11501,N_11091,N_11229);
nor U11502 (N_11502,N_11440,N_11230);
nor U11503 (N_11503,N_11312,N_11470);
and U11504 (N_11504,N_11176,N_11203);
nand U11505 (N_11505,N_11194,N_11274);
nor U11506 (N_11506,N_11449,N_11404);
and U11507 (N_11507,N_11188,N_11047);
nor U11508 (N_11508,N_11461,N_11074);
nand U11509 (N_11509,N_11077,N_11307);
xnor U11510 (N_11510,N_11150,N_11345);
and U11511 (N_11511,N_11298,N_11380);
nand U11512 (N_11512,N_11186,N_11370);
xor U11513 (N_11513,N_11116,N_11130);
and U11514 (N_11514,N_11154,N_11008);
nor U11515 (N_11515,N_11488,N_11491);
xor U11516 (N_11516,N_11347,N_11287);
nor U11517 (N_11517,N_11215,N_11143);
and U11518 (N_11518,N_11259,N_11221);
and U11519 (N_11519,N_11368,N_11072);
and U11520 (N_11520,N_11324,N_11463);
nand U11521 (N_11521,N_11196,N_11381);
nor U11522 (N_11522,N_11015,N_11220);
nand U11523 (N_11523,N_11087,N_11019);
xor U11524 (N_11524,N_11457,N_11068);
and U11525 (N_11525,N_11344,N_11302);
xnor U11526 (N_11526,N_11349,N_11026);
xnor U11527 (N_11527,N_11295,N_11290);
nor U11528 (N_11528,N_11299,N_11313);
nor U11529 (N_11529,N_11359,N_11148);
nand U11530 (N_11530,N_11284,N_11331);
nor U11531 (N_11531,N_11139,N_11242);
or U11532 (N_11532,N_11018,N_11371);
nor U11533 (N_11533,N_11180,N_11360);
xnor U11534 (N_11534,N_11403,N_11400);
or U11535 (N_11535,N_11046,N_11235);
xor U11536 (N_11536,N_11320,N_11214);
and U11537 (N_11537,N_11192,N_11064);
nand U11538 (N_11538,N_11459,N_11399);
nand U11539 (N_11539,N_11390,N_11051);
or U11540 (N_11540,N_11498,N_11117);
xor U11541 (N_11541,N_11121,N_11132);
or U11542 (N_11542,N_11474,N_11244);
xor U11543 (N_11543,N_11266,N_11401);
and U11544 (N_11544,N_11469,N_11375);
or U11545 (N_11545,N_11483,N_11078);
nand U11546 (N_11546,N_11282,N_11175);
nor U11547 (N_11547,N_11454,N_11044);
xor U11548 (N_11548,N_11408,N_11279);
xnor U11549 (N_11549,N_11391,N_11138);
xnor U11550 (N_11550,N_11104,N_11387);
or U11551 (N_11551,N_11226,N_11351);
nand U11552 (N_11552,N_11346,N_11092);
nand U11553 (N_11553,N_11246,N_11288);
or U11554 (N_11554,N_11239,N_11329);
and U11555 (N_11555,N_11211,N_11140);
and U11556 (N_11556,N_11445,N_11029);
xnor U11557 (N_11557,N_11361,N_11183);
xor U11558 (N_11558,N_11070,N_11362);
or U11559 (N_11559,N_11115,N_11448);
nand U11560 (N_11560,N_11396,N_11228);
nand U11561 (N_11561,N_11415,N_11450);
and U11562 (N_11562,N_11268,N_11340);
and U11563 (N_11563,N_11350,N_11293);
or U11564 (N_11564,N_11366,N_11159);
or U11565 (N_11565,N_11218,N_11170);
nor U11566 (N_11566,N_11195,N_11248);
or U11567 (N_11567,N_11010,N_11076);
and U11568 (N_11568,N_11128,N_11202);
and U11569 (N_11569,N_11283,N_11304);
or U11570 (N_11570,N_11338,N_11249);
nand U11571 (N_11571,N_11037,N_11405);
and U11572 (N_11572,N_11050,N_11082);
and U11573 (N_11573,N_11069,N_11059);
nand U11574 (N_11574,N_11341,N_11427);
or U11575 (N_11575,N_11199,N_11270);
xor U11576 (N_11576,N_11397,N_11086);
nand U11577 (N_11577,N_11464,N_11099);
or U11578 (N_11578,N_11442,N_11492);
or U11579 (N_11579,N_11061,N_11236);
and U11580 (N_11580,N_11063,N_11152);
xnor U11581 (N_11581,N_11250,N_11447);
xor U11582 (N_11582,N_11004,N_11429);
and U11583 (N_11583,N_11053,N_11308);
and U11584 (N_11584,N_11319,N_11316);
nand U11585 (N_11585,N_11205,N_11093);
or U11586 (N_11586,N_11420,N_11281);
or U11587 (N_11587,N_11422,N_11251);
or U11588 (N_11588,N_11261,N_11042);
and U11589 (N_11589,N_11339,N_11490);
nor U11590 (N_11590,N_11353,N_11499);
or U11591 (N_11591,N_11465,N_11022);
or U11592 (N_11592,N_11437,N_11052);
nand U11593 (N_11593,N_11496,N_11142);
xnor U11594 (N_11594,N_11000,N_11389);
nor U11595 (N_11595,N_11134,N_11267);
nor U11596 (N_11596,N_11164,N_11151);
nand U11597 (N_11597,N_11439,N_11033);
nor U11598 (N_11598,N_11277,N_11455);
nand U11599 (N_11599,N_11446,N_11157);
xnor U11600 (N_11600,N_11210,N_11017);
or U11601 (N_11601,N_11482,N_11342);
or U11602 (N_11602,N_11386,N_11060);
or U11603 (N_11603,N_11145,N_11257);
nor U11604 (N_11604,N_11080,N_11048);
nor U11605 (N_11605,N_11300,N_11125);
nand U11606 (N_11606,N_11275,N_11055);
and U11607 (N_11607,N_11315,N_11385);
or U11608 (N_11608,N_11306,N_11096);
and U11609 (N_11609,N_11326,N_11426);
nand U11610 (N_11610,N_11119,N_11158);
xnor U11611 (N_11611,N_11224,N_11083);
or U11612 (N_11612,N_11468,N_11081);
and U11613 (N_11613,N_11208,N_11146);
or U11614 (N_11614,N_11495,N_11172);
or U11615 (N_11615,N_11460,N_11497);
and U11616 (N_11616,N_11373,N_11179);
and U11617 (N_11617,N_11321,N_11434);
or U11618 (N_11618,N_11206,N_11003);
and U11619 (N_11619,N_11262,N_11184);
nor U11620 (N_11620,N_11101,N_11041);
nor U11621 (N_11621,N_11009,N_11289);
and U11622 (N_11622,N_11038,N_11238);
nand U11623 (N_11623,N_11020,N_11189);
and U11624 (N_11624,N_11173,N_11384);
and U11625 (N_11625,N_11127,N_11040);
or U11626 (N_11626,N_11309,N_11109);
or U11627 (N_11627,N_11278,N_11049);
nand U11628 (N_11628,N_11084,N_11197);
xor U11629 (N_11629,N_11255,N_11365);
xor U11630 (N_11630,N_11475,N_11131);
or U11631 (N_11631,N_11424,N_11054);
and U11632 (N_11632,N_11466,N_11433);
nor U11633 (N_11633,N_11233,N_11322);
xnor U11634 (N_11634,N_11123,N_11379);
xor U11635 (N_11635,N_11398,N_11155);
nor U11636 (N_11636,N_11032,N_11129);
nand U11637 (N_11637,N_11073,N_11471);
nand U11638 (N_11638,N_11178,N_11135);
nor U11639 (N_11639,N_11149,N_11332);
nor U11640 (N_11640,N_11237,N_11147);
and U11641 (N_11641,N_11191,N_11480);
xnor U11642 (N_11642,N_11182,N_11207);
xor U11643 (N_11643,N_11269,N_11122);
nand U11644 (N_11644,N_11436,N_11095);
nand U11645 (N_11645,N_11062,N_11264);
or U11646 (N_11646,N_11328,N_11174);
xnor U11647 (N_11647,N_11413,N_11240);
xor U11648 (N_11648,N_11376,N_11247);
and U11649 (N_11649,N_11271,N_11303);
nor U11650 (N_11650,N_11406,N_11356);
xor U11651 (N_11651,N_11336,N_11355);
nor U11652 (N_11652,N_11486,N_11167);
and U11653 (N_11653,N_11419,N_11161);
and U11654 (N_11654,N_11438,N_11337);
or U11655 (N_11655,N_11007,N_11013);
and U11656 (N_11656,N_11372,N_11011);
or U11657 (N_11657,N_11113,N_11291);
or U11658 (N_11658,N_11169,N_11407);
or U11659 (N_11659,N_11006,N_11036);
and U11660 (N_11660,N_11168,N_11067);
or U11661 (N_11661,N_11014,N_11369);
and U11662 (N_11662,N_11252,N_11079);
and U11663 (N_11663,N_11243,N_11477);
or U11664 (N_11664,N_11108,N_11357);
nor U11665 (N_11665,N_11198,N_11473);
or U11666 (N_11666,N_11330,N_11162);
xnor U11667 (N_11667,N_11035,N_11417);
or U11668 (N_11668,N_11388,N_11034);
xor U11669 (N_11669,N_11023,N_11256);
or U11670 (N_11670,N_11394,N_11212);
and U11671 (N_11671,N_11137,N_11317);
xnor U11672 (N_11672,N_11098,N_11416);
nand U11673 (N_11673,N_11493,N_11421);
or U11674 (N_11674,N_11039,N_11156);
nand U11675 (N_11675,N_11476,N_11343);
nand U11676 (N_11676,N_11335,N_11367);
nand U11677 (N_11677,N_11043,N_11297);
nand U11678 (N_11678,N_11024,N_11441);
and U11679 (N_11679,N_11005,N_11325);
or U11680 (N_11680,N_11352,N_11213);
nor U11681 (N_11681,N_11276,N_11219);
or U11682 (N_11682,N_11412,N_11430);
nor U11683 (N_11683,N_11494,N_11136);
or U11684 (N_11684,N_11310,N_11481);
and U11685 (N_11685,N_11258,N_11395);
or U11686 (N_11686,N_11333,N_11462);
xor U11687 (N_11687,N_11354,N_11432);
nand U11688 (N_11688,N_11012,N_11374);
xor U11689 (N_11689,N_11280,N_11314);
or U11690 (N_11690,N_11444,N_11102);
nand U11691 (N_11691,N_11021,N_11263);
and U11692 (N_11692,N_11204,N_11414);
nor U11693 (N_11693,N_11489,N_11472);
nor U11694 (N_11694,N_11100,N_11253);
and U11695 (N_11695,N_11065,N_11106);
nand U11696 (N_11696,N_11377,N_11364);
nor U11697 (N_11697,N_11285,N_11056);
nor U11698 (N_11698,N_11088,N_11160);
xor U11699 (N_11699,N_11431,N_11286);
nor U11700 (N_11700,N_11058,N_11254);
and U11701 (N_11701,N_11002,N_11232);
nor U11702 (N_11702,N_11292,N_11227);
nor U11703 (N_11703,N_11234,N_11085);
nor U11704 (N_11704,N_11111,N_11045);
or U11705 (N_11705,N_11456,N_11110);
nand U11706 (N_11706,N_11318,N_11141);
nand U11707 (N_11707,N_11435,N_11177);
nand U11708 (N_11708,N_11231,N_11479);
nand U11709 (N_11709,N_11225,N_11423);
nor U11710 (N_11710,N_11209,N_11163);
xor U11711 (N_11711,N_11166,N_11348);
nor U11712 (N_11712,N_11165,N_11071);
and U11713 (N_11713,N_11181,N_11467);
and U11714 (N_11714,N_11443,N_11027);
xnor U11715 (N_11715,N_11066,N_11144);
xor U11716 (N_11716,N_11216,N_11382);
nor U11717 (N_11717,N_11334,N_11112);
xor U11718 (N_11718,N_11031,N_11378);
and U11719 (N_11719,N_11030,N_11296);
nor U11720 (N_11720,N_11458,N_11265);
and U11721 (N_11721,N_11410,N_11323);
and U11722 (N_11722,N_11418,N_11363);
xor U11723 (N_11723,N_11453,N_11305);
nor U11724 (N_11724,N_11025,N_11016);
and U11725 (N_11725,N_11392,N_11311);
nand U11726 (N_11726,N_11223,N_11001);
nor U11727 (N_11727,N_11193,N_11114);
or U11728 (N_11728,N_11245,N_11241);
or U11729 (N_11729,N_11153,N_11478);
xnor U11730 (N_11730,N_11118,N_11393);
and U11731 (N_11731,N_11383,N_11185);
xnor U11732 (N_11732,N_11107,N_11452);
xnor U11733 (N_11733,N_11097,N_11487);
or U11734 (N_11734,N_11217,N_11171);
nor U11735 (N_11735,N_11222,N_11428);
and U11736 (N_11736,N_11451,N_11089);
nand U11737 (N_11737,N_11090,N_11327);
xnor U11738 (N_11738,N_11126,N_11190);
nand U11739 (N_11739,N_11402,N_11260);
or U11740 (N_11740,N_11028,N_11273);
xnor U11741 (N_11741,N_11075,N_11484);
xor U11742 (N_11742,N_11272,N_11200);
nand U11743 (N_11743,N_11124,N_11409);
or U11744 (N_11744,N_11301,N_11485);
nor U11745 (N_11745,N_11187,N_11358);
nor U11746 (N_11746,N_11411,N_11294);
xnor U11747 (N_11747,N_11105,N_11103);
and U11748 (N_11748,N_11120,N_11201);
xnor U11749 (N_11749,N_11425,N_11094);
nor U11750 (N_11750,N_11230,N_11351);
nor U11751 (N_11751,N_11160,N_11318);
xnor U11752 (N_11752,N_11271,N_11350);
nand U11753 (N_11753,N_11112,N_11259);
xnor U11754 (N_11754,N_11446,N_11036);
xor U11755 (N_11755,N_11360,N_11013);
nand U11756 (N_11756,N_11312,N_11095);
nand U11757 (N_11757,N_11461,N_11455);
nor U11758 (N_11758,N_11315,N_11380);
nor U11759 (N_11759,N_11116,N_11153);
nand U11760 (N_11760,N_11013,N_11213);
nand U11761 (N_11761,N_11085,N_11241);
and U11762 (N_11762,N_11146,N_11401);
nand U11763 (N_11763,N_11210,N_11089);
or U11764 (N_11764,N_11292,N_11357);
or U11765 (N_11765,N_11078,N_11213);
xor U11766 (N_11766,N_11475,N_11316);
xor U11767 (N_11767,N_11058,N_11057);
nand U11768 (N_11768,N_11248,N_11170);
or U11769 (N_11769,N_11042,N_11229);
xor U11770 (N_11770,N_11173,N_11273);
nor U11771 (N_11771,N_11168,N_11135);
and U11772 (N_11772,N_11026,N_11223);
or U11773 (N_11773,N_11029,N_11368);
nor U11774 (N_11774,N_11132,N_11276);
nor U11775 (N_11775,N_11112,N_11199);
and U11776 (N_11776,N_11347,N_11257);
xnor U11777 (N_11777,N_11372,N_11284);
nor U11778 (N_11778,N_11150,N_11222);
and U11779 (N_11779,N_11113,N_11379);
xor U11780 (N_11780,N_11488,N_11205);
or U11781 (N_11781,N_11186,N_11223);
xnor U11782 (N_11782,N_11453,N_11340);
nand U11783 (N_11783,N_11353,N_11026);
and U11784 (N_11784,N_11178,N_11020);
nand U11785 (N_11785,N_11288,N_11498);
nor U11786 (N_11786,N_11118,N_11079);
nand U11787 (N_11787,N_11304,N_11118);
and U11788 (N_11788,N_11014,N_11337);
xnor U11789 (N_11789,N_11261,N_11200);
nand U11790 (N_11790,N_11182,N_11251);
xor U11791 (N_11791,N_11168,N_11307);
and U11792 (N_11792,N_11386,N_11126);
and U11793 (N_11793,N_11411,N_11053);
nand U11794 (N_11794,N_11067,N_11192);
and U11795 (N_11795,N_11028,N_11186);
xnor U11796 (N_11796,N_11248,N_11386);
nand U11797 (N_11797,N_11106,N_11374);
xor U11798 (N_11798,N_11282,N_11060);
nor U11799 (N_11799,N_11217,N_11143);
nand U11800 (N_11800,N_11035,N_11076);
nand U11801 (N_11801,N_11437,N_11419);
nand U11802 (N_11802,N_11304,N_11087);
or U11803 (N_11803,N_11385,N_11406);
nor U11804 (N_11804,N_11338,N_11063);
nand U11805 (N_11805,N_11253,N_11237);
nand U11806 (N_11806,N_11397,N_11390);
or U11807 (N_11807,N_11289,N_11126);
and U11808 (N_11808,N_11170,N_11267);
nor U11809 (N_11809,N_11465,N_11015);
nor U11810 (N_11810,N_11309,N_11418);
and U11811 (N_11811,N_11279,N_11088);
nand U11812 (N_11812,N_11431,N_11191);
nor U11813 (N_11813,N_11232,N_11267);
xnor U11814 (N_11814,N_11264,N_11033);
nor U11815 (N_11815,N_11439,N_11023);
and U11816 (N_11816,N_11176,N_11043);
or U11817 (N_11817,N_11456,N_11396);
xor U11818 (N_11818,N_11329,N_11289);
and U11819 (N_11819,N_11357,N_11233);
nand U11820 (N_11820,N_11269,N_11400);
nor U11821 (N_11821,N_11419,N_11429);
xnor U11822 (N_11822,N_11440,N_11226);
nand U11823 (N_11823,N_11470,N_11059);
or U11824 (N_11824,N_11037,N_11128);
nor U11825 (N_11825,N_11430,N_11036);
xnor U11826 (N_11826,N_11307,N_11217);
nor U11827 (N_11827,N_11212,N_11411);
nand U11828 (N_11828,N_11395,N_11110);
nor U11829 (N_11829,N_11218,N_11032);
nand U11830 (N_11830,N_11078,N_11193);
and U11831 (N_11831,N_11115,N_11363);
or U11832 (N_11832,N_11236,N_11146);
and U11833 (N_11833,N_11110,N_11313);
nand U11834 (N_11834,N_11019,N_11295);
xor U11835 (N_11835,N_11438,N_11255);
nor U11836 (N_11836,N_11497,N_11230);
nand U11837 (N_11837,N_11181,N_11278);
nor U11838 (N_11838,N_11008,N_11195);
and U11839 (N_11839,N_11444,N_11084);
nor U11840 (N_11840,N_11360,N_11130);
and U11841 (N_11841,N_11408,N_11367);
nor U11842 (N_11842,N_11141,N_11268);
xnor U11843 (N_11843,N_11146,N_11068);
xnor U11844 (N_11844,N_11158,N_11353);
or U11845 (N_11845,N_11381,N_11408);
nand U11846 (N_11846,N_11211,N_11419);
or U11847 (N_11847,N_11165,N_11428);
nor U11848 (N_11848,N_11050,N_11436);
xnor U11849 (N_11849,N_11078,N_11219);
or U11850 (N_11850,N_11154,N_11313);
xor U11851 (N_11851,N_11235,N_11404);
or U11852 (N_11852,N_11052,N_11002);
or U11853 (N_11853,N_11251,N_11198);
nor U11854 (N_11854,N_11373,N_11340);
or U11855 (N_11855,N_11468,N_11002);
nor U11856 (N_11856,N_11107,N_11051);
nor U11857 (N_11857,N_11244,N_11179);
nor U11858 (N_11858,N_11223,N_11195);
and U11859 (N_11859,N_11130,N_11107);
and U11860 (N_11860,N_11159,N_11125);
and U11861 (N_11861,N_11065,N_11145);
xnor U11862 (N_11862,N_11284,N_11425);
xnor U11863 (N_11863,N_11181,N_11014);
or U11864 (N_11864,N_11236,N_11460);
xor U11865 (N_11865,N_11197,N_11036);
and U11866 (N_11866,N_11294,N_11475);
and U11867 (N_11867,N_11469,N_11295);
nand U11868 (N_11868,N_11167,N_11054);
nand U11869 (N_11869,N_11073,N_11085);
and U11870 (N_11870,N_11387,N_11034);
nand U11871 (N_11871,N_11495,N_11479);
or U11872 (N_11872,N_11418,N_11062);
xnor U11873 (N_11873,N_11218,N_11079);
xnor U11874 (N_11874,N_11481,N_11373);
nor U11875 (N_11875,N_11232,N_11263);
or U11876 (N_11876,N_11068,N_11013);
or U11877 (N_11877,N_11329,N_11197);
nor U11878 (N_11878,N_11381,N_11323);
or U11879 (N_11879,N_11099,N_11405);
and U11880 (N_11880,N_11367,N_11170);
and U11881 (N_11881,N_11359,N_11025);
or U11882 (N_11882,N_11236,N_11189);
nor U11883 (N_11883,N_11419,N_11091);
xor U11884 (N_11884,N_11428,N_11175);
nand U11885 (N_11885,N_11037,N_11365);
xnor U11886 (N_11886,N_11253,N_11198);
nor U11887 (N_11887,N_11308,N_11417);
nor U11888 (N_11888,N_11217,N_11092);
nand U11889 (N_11889,N_11426,N_11307);
and U11890 (N_11890,N_11335,N_11243);
nand U11891 (N_11891,N_11010,N_11061);
and U11892 (N_11892,N_11436,N_11042);
or U11893 (N_11893,N_11055,N_11004);
and U11894 (N_11894,N_11278,N_11227);
and U11895 (N_11895,N_11163,N_11446);
or U11896 (N_11896,N_11069,N_11435);
nor U11897 (N_11897,N_11438,N_11400);
xnor U11898 (N_11898,N_11171,N_11275);
and U11899 (N_11899,N_11361,N_11303);
nand U11900 (N_11900,N_11123,N_11025);
or U11901 (N_11901,N_11391,N_11257);
nand U11902 (N_11902,N_11406,N_11104);
nor U11903 (N_11903,N_11133,N_11490);
nor U11904 (N_11904,N_11020,N_11233);
nor U11905 (N_11905,N_11334,N_11123);
xor U11906 (N_11906,N_11299,N_11155);
xnor U11907 (N_11907,N_11055,N_11017);
xor U11908 (N_11908,N_11179,N_11366);
xnor U11909 (N_11909,N_11435,N_11095);
nor U11910 (N_11910,N_11322,N_11348);
nor U11911 (N_11911,N_11058,N_11166);
and U11912 (N_11912,N_11269,N_11464);
nand U11913 (N_11913,N_11040,N_11296);
nor U11914 (N_11914,N_11137,N_11459);
or U11915 (N_11915,N_11290,N_11486);
xor U11916 (N_11916,N_11458,N_11408);
nand U11917 (N_11917,N_11302,N_11445);
nor U11918 (N_11918,N_11036,N_11473);
nor U11919 (N_11919,N_11027,N_11308);
xor U11920 (N_11920,N_11428,N_11384);
and U11921 (N_11921,N_11251,N_11150);
nand U11922 (N_11922,N_11261,N_11333);
nand U11923 (N_11923,N_11318,N_11360);
nor U11924 (N_11924,N_11017,N_11344);
xor U11925 (N_11925,N_11341,N_11334);
nand U11926 (N_11926,N_11156,N_11117);
nand U11927 (N_11927,N_11072,N_11196);
or U11928 (N_11928,N_11420,N_11043);
nand U11929 (N_11929,N_11447,N_11105);
nand U11930 (N_11930,N_11461,N_11312);
or U11931 (N_11931,N_11004,N_11449);
and U11932 (N_11932,N_11402,N_11106);
nor U11933 (N_11933,N_11354,N_11264);
nor U11934 (N_11934,N_11226,N_11281);
nor U11935 (N_11935,N_11338,N_11425);
and U11936 (N_11936,N_11342,N_11274);
nor U11937 (N_11937,N_11194,N_11067);
nor U11938 (N_11938,N_11019,N_11074);
nand U11939 (N_11939,N_11257,N_11064);
nor U11940 (N_11940,N_11244,N_11040);
nor U11941 (N_11941,N_11479,N_11415);
xnor U11942 (N_11942,N_11158,N_11020);
xor U11943 (N_11943,N_11046,N_11440);
xnor U11944 (N_11944,N_11227,N_11105);
nor U11945 (N_11945,N_11164,N_11006);
nand U11946 (N_11946,N_11178,N_11042);
nand U11947 (N_11947,N_11400,N_11073);
nand U11948 (N_11948,N_11090,N_11005);
nor U11949 (N_11949,N_11284,N_11450);
or U11950 (N_11950,N_11360,N_11190);
nand U11951 (N_11951,N_11247,N_11440);
or U11952 (N_11952,N_11492,N_11305);
nand U11953 (N_11953,N_11369,N_11325);
or U11954 (N_11954,N_11176,N_11096);
and U11955 (N_11955,N_11357,N_11206);
nand U11956 (N_11956,N_11313,N_11381);
nand U11957 (N_11957,N_11207,N_11037);
xnor U11958 (N_11958,N_11077,N_11065);
xor U11959 (N_11959,N_11050,N_11189);
xor U11960 (N_11960,N_11063,N_11331);
nand U11961 (N_11961,N_11380,N_11253);
xnor U11962 (N_11962,N_11409,N_11301);
xnor U11963 (N_11963,N_11389,N_11458);
and U11964 (N_11964,N_11292,N_11344);
nand U11965 (N_11965,N_11204,N_11345);
nand U11966 (N_11966,N_11197,N_11210);
nand U11967 (N_11967,N_11018,N_11239);
and U11968 (N_11968,N_11461,N_11458);
xnor U11969 (N_11969,N_11388,N_11420);
and U11970 (N_11970,N_11292,N_11404);
nand U11971 (N_11971,N_11094,N_11374);
nor U11972 (N_11972,N_11379,N_11185);
and U11973 (N_11973,N_11414,N_11157);
xor U11974 (N_11974,N_11351,N_11364);
xnor U11975 (N_11975,N_11478,N_11158);
nor U11976 (N_11976,N_11253,N_11113);
nand U11977 (N_11977,N_11067,N_11219);
or U11978 (N_11978,N_11206,N_11464);
and U11979 (N_11979,N_11033,N_11114);
and U11980 (N_11980,N_11362,N_11405);
and U11981 (N_11981,N_11138,N_11029);
and U11982 (N_11982,N_11087,N_11163);
nand U11983 (N_11983,N_11366,N_11098);
nor U11984 (N_11984,N_11111,N_11096);
nor U11985 (N_11985,N_11489,N_11425);
nand U11986 (N_11986,N_11166,N_11095);
and U11987 (N_11987,N_11262,N_11379);
nand U11988 (N_11988,N_11190,N_11446);
or U11989 (N_11989,N_11237,N_11338);
or U11990 (N_11990,N_11479,N_11063);
xor U11991 (N_11991,N_11328,N_11386);
nor U11992 (N_11992,N_11438,N_11078);
or U11993 (N_11993,N_11440,N_11190);
and U11994 (N_11994,N_11250,N_11345);
xnor U11995 (N_11995,N_11090,N_11113);
nor U11996 (N_11996,N_11135,N_11046);
xnor U11997 (N_11997,N_11176,N_11174);
nand U11998 (N_11998,N_11141,N_11145);
xor U11999 (N_11999,N_11017,N_11338);
nor U12000 (N_12000,N_11643,N_11614);
xor U12001 (N_12001,N_11872,N_11938);
nand U12002 (N_12002,N_11548,N_11718);
or U12003 (N_12003,N_11734,N_11803);
and U12004 (N_12004,N_11966,N_11521);
xor U12005 (N_12005,N_11895,N_11630);
xnor U12006 (N_12006,N_11645,N_11852);
xor U12007 (N_12007,N_11514,N_11914);
and U12008 (N_12008,N_11880,N_11633);
nand U12009 (N_12009,N_11580,N_11737);
xor U12010 (N_12010,N_11976,N_11573);
xor U12011 (N_12011,N_11807,N_11908);
nor U12012 (N_12012,N_11667,N_11819);
and U12013 (N_12013,N_11970,N_11971);
xnor U12014 (N_12014,N_11528,N_11508);
xor U12015 (N_12015,N_11607,N_11978);
and U12016 (N_12016,N_11663,N_11617);
or U12017 (N_12017,N_11629,N_11652);
and U12018 (N_12018,N_11861,N_11700);
and U12019 (N_12019,N_11958,N_11500);
nand U12020 (N_12020,N_11815,N_11527);
nor U12021 (N_12021,N_11841,N_11790);
and U12022 (N_12022,N_11870,N_11677);
nor U12023 (N_12023,N_11919,N_11632);
and U12024 (N_12024,N_11862,N_11967);
nor U12025 (N_12025,N_11795,N_11986);
nand U12026 (N_12026,N_11741,N_11955);
and U12027 (N_12027,N_11544,N_11798);
and U12028 (N_12028,N_11695,N_11532);
xnor U12029 (N_12029,N_11639,N_11713);
nor U12030 (N_12030,N_11877,N_11930);
xor U12031 (N_12031,N_11811,N_11927);
xnor U12032 (N_12032,N_11937,N_11601);
nor U12033 (N_12033,N_11817,N_11520);
nand U12034 (N_12034,N_11975,N_11826);
or U12035 (N_12035,N_11769,N_11956);
or U12036 (N_12036,N_11511,N_11996);
xor U12037 (N_12037,N_11555,N_11923);
or U12038 (N_12038,N_11689,N_11954);
and U12039 (N_12039,N_11653,N_11805);
and U12040 (N_12040,N_11832,N_11673);
nor U12041 (N_12041,N_11944,N_11507);
nand U12042 (N_12042,N_11712,N_11879);
nor U12043 (N_12043,N_11681,N_11679);
and U12044 (N_12044,N_11744,N_11961);
nand U12045 (N_12045,N_11921,N_11878);
or U12046 (N_12046,N_11813,N_11530);
or U12047 (N_12047,N_11776,N_11503);
nor U12048 (N_12048,N_11788,N_11587);
or U12049 (N_12049,N_11814,N_11567);
xor U12050 (N_12050,N_11786,N_11572);
xor U12051 (N_12051,N_11513,N_11929);
and U12052 (N_12052,N_11721,N_11636);
or U12053 (N_12053,N_11640,N_11605);
xor U12054 (N_12054,N_11594,N_11599);
nor U12055 (N_12055,N_11609,N_11606);
nor U12056 (N_12056,N_11957,N_11538);
nand U12057 (N_12057,N_11922,N_11539);
xnor U12058 (N_12058,N_11896,N_11725);
nand U12059 (N_12059,N_11748,N_11738);
nand U12060 (N_12060,N_11796,N_11899);
nand U12061 (N_12061,N_11684,N_11714);
xnor U12062 (N_12062,N_11926,N_11698);
nor U12063 (N_12063,N_11973,N_11728);
nand U12064 (N_12064,N_11835,N_11886);
nor U12065 (N_12065,N_11924,N_11549);
or U12066 (N_12066,N_11506,N_11952);
nand U12067 (N_12067,N_11512,N_11794);
nor U12068 (N_12068,N_11907,N_11875);
and U12069 (N_12069,N_11551,N_11859);
xor U12070 (N_12070,N_11887,N_11550);
nand U12071 (N_12071,N_11627,N_11889);
or U12072 (N_12072,N_11683,N_11543);
nand U12073 (N_12073,N_11623,N_11591);
nand U12074 (N_12074,N_11766,N_11959);
nor U12075 (N_12075,N_11925,N_11866);
nand U12076 (N_12076,N_11704,N_11767);
xor U12077 (N_12077,N_11916,N_11867);
nor U12078 (N_12078,N_11680,N_11724);
nor U12079 (N_12079,N_11830,N_11563);
and U12080 (N_12080,N_11598,N_11701);
nand U12081 (N_12081,N_11770,N_11736);
xor U12082 (N_12082,N_11509,N_11556);
xnor U12083 (N_12083,N_11780,N_11574);
and U12084 (N_12084,N_11988,N_11746);
and U12085 (N_12085,N_11933,N_11647);
or U12086 (N_12086,N_11934,N_11537);
and U12087 (N_12087,N_11984,N_11545);
nand U12088 (N_12088,N_11827,N_11901);
nor U12089 (N_12089,N_11604,N_11762);
and U12090 (N_12090,N_11840,N_11851);
xor U12091 (N_12091,N_11857,N_11833);
nand U12092 (N_12092,N_11592,N_11611);
xnor U12093 (N_12093,N_11571,N_11804);
nor U12094 (N_12094,N_11999,N_11898);
or U12095 (N_12095,N_11661,N_11995);
nor U12096 (N_12096,N_11517,N_11960);
nand U12097 (N_12097,N_11991,N_11900);
xnor U12098 (N_12098,N_11962,N_11729);
nand U12099 (N_12099,N_11595,N_11529);
or U12100 (N_12100,N_11524,N_11672);
and U12101 (N_12101,N_11932,N_11755);
nor U12102 (N_12102,N_11608,N_11918);
nand U12103 (N_12103,N_11596,N_11874);
and U12104 (N_12104,N_11763,N_11635);
xor U12105 (N_12105,N_11800,N_11818);
xor U12106 (N_12106,N_11660,N_11836);
xor U12107 (N_12107,N_11773,N_11749);
and U12108 (N_12108,N_11553,N_11992);
or U12109 (N_12109,N_11624,N_11651);
xnor U12110 (N_12110,N_11946,N_11733);
nand U12111 (N_12111,N_11579,N_11501);
xor U12112 (N_12112,N_11658,N_11585);
or U12113 (N_12113,N_11847,N_11715);
xnor U12114 (N_12114,N_11759,N_11902);
nor U12115 (N_12115,N_11522,N_11758);
nor U12116 (N_12116,N_11690,N_11732);
or U12117 (N_12117,N_11820,N_11634);
or U12118 (N_12118,N_11742,N_11824);
nand U12119 (N_12119,N_11552,N_11519);
nor U12120 (N_12120,N_11618,N_11903);
nor U12121 (N_12121,N_11829,N_11989);
xor U12122 (N_12122,N_11943,N_11536);
or U12123 (N_12123,N_11883,N_11799);
nand U12124 (N_12124,N_11787,N_11577);
nand U12125 (N_12125,N_11936,N_11590);
nor U12126 (N_12126,N_11757,N_11584);
nand U12127 (N_12127,N_11912,N_11541);
and U12128 (N_12128,N_11842,N_11593);
nor U12129 (N_12129,N_11682,N_11864);
and U12130 (N_12130,N_11793,N_11745);
or U12131 (N_12131,N_11703,N_11910);
and U12132 (N_12132,N_11772,N_11674);
nor U12133 (N_12133,N_11656,N_11863);
and U12134 (N_12134,N_11844,N_11917);
nor U12135 (N_12135,N_11760,N_11822);
xor U12136 (N_12136,N_11823,N_11678);
nor U12137 (N_12137,N_11953,N_11783);
nor U12138 (N_12138,N_11735,N_11638);
and U12139 (N_12139,N_11569,N_11846);
or U12140 (N_12140,N_11982,N_11825);
or U12141 (N_12141,N_11644,N_11687);
nand U12142 (N_12142,N_11810,N_11802);
nor U12143 (N_12143,N_11942,N_11963);
nand U12144 (N_12144,N_11781,N_11565);
or U12145 (N_12145,N_11706,N_11619);
or U12146 (N_12146,N_11650,N_11675);
xor U12147 (N_12147,N_11694,N_11560);
and U12148 (N_12148,N_11777,N_11821);
nand U12149 (N_12149,N_11747,N_11568);
nand U12150 (N_12150,N_11945,N_11588);
and U12151 (N_12151,N_11516,N_11784);
nand U12152 (N_12152,N_11581,N_11646);
nor U12153 (N_12153,N_11950,N_11720);
and U12154 (N_12154,N_11515,N_11968);
nand U12155 (N_12155,N_11535,N_11664);
or U12156 (N_12156,N_11564,N_11985);
or U12157 (N_12157,N_11751,N_11797);
or U12158 (N_12158,N_11994,N_11668);
nand U12159 (N_12159,N_11940,N_11812);
nor U12160 (N_12160,N_11626,N_11727);
or U12161 (N_12161,N_11540,N_11597);
nand U12162 (N_12162,N_11774,N_11981);
and U12163 (N_12163,N_11941,N_11603);
nor U12164 (N_12164,N_11602,N_11890);
xor U12165 (N_12165,N_11709,N_11809);
and U12166 (N_12166,N_11882,N_11719);
and U12167 (N_12167,N_11625,N_11716);
and U12168 (N_12168,N_11974,N_11837);
nand U12169 (N_12169,N_11534,N_11561);
xnor U12170 (N_12170,N_11913,N_11756);
and U12171 (N_12171,N_11613,N_11722);
nor U12172 (N_12172,N_11785,N_11686);
or U12173 (N_12173,N_11616,N_11845);
and U12174 (N_12174,N_11979,N_11685);
and U12175 (N_12175,N_11600,N_11637);
nor U12176 (N_12176,N_11533,N_11723);
nand U12177 (N_12177,N_11881,N_11504);
or U12178 (N_12178,N_11987,N_11909);
or U12179 (N_12179,N_11868,N_11858);
nor U12180 (N_12180,N_11575,N_11764);
and U12181 (N_12181,N_11666,N_11731);
or U12182 (N_12182,N_11849,N_11782);
xor U12183 (N_12183,N_11854,N_11894);
nand U12184 (N_12184,N_11615,N_11775);
nand U12185 (N_12185,N_11642,N_11789);
xor U12186 (N_12186,N_11948,N_11570);
nor U12187 (N_12187,N_11949,N_11993);
or U12188 (N_12188,N_11947,N_11977);
nand U12189 (N_12189,N_11843,N_11920);
nor U12190 (N_12190,N_11885,N_11905);
xnor U12191 (N_12191,N_11693,N_11641);
and U12192 (N_12192,N_11710,N_11939);
and U12193 (N_12193,N_11692,N_11771);
or U12194 (N_12194,N_11865,N_11816);
nor U12195 (N_12195,N_11765,N_11702);
and U12196 (N_12196,N_11891,N_11631);
and U12197 (N_12197,N_11582,N_11649);
nand U12198 (N_12198,N_11998,N_11904);
xor U12199 (N_12199,N_11662,N_11853);
nand U12200 (N_12200,N_11876,N_11965);
nand U12201 (N_12201,N_11557,N_11523);
or U12202 (N_12202,N_11806,N_11951);
or U12203 (N_12203,N_11697,N_11928);
xnor U12204 (N_12204,N_11831,N_11665);
xnor U12205 (N_12205,N_11688,N_11583);
xnor U12206 (N_12206,N_11696,N_11931);
and U12207 (N_12207,N_11502,N_11612);
and U12208 (N_12208,N_11610,N_11911);
xnor U12209 (N_12209,N_11791,N_11670);
or U12210 (N_12210,N_11873,N_11983);
and U12211 (N_12211,N_11622,N_11743);
nor U12212 (N_12212,N_11871,N_11739);
nand U12213 (N_12213,N_11589,N_11547);
or U12214 (N_12214,N_11838,N_11969);
or U12215 (N_12215,N_11620,N_11860);
xor U12216 (N_12216,N_11671,N_11750);
nand U12217 (N_12217,N_11761,N_11518);
xor U12218 (N_12218,N_11669,N_11578);
nand U12219 (N_12219,N_11754,N_11730);
or U12220 (N_12220,N_11768,N_11856);
and U12221 (N_12221,N_11834,N_11542);
xor U12222 (N_12222,N_11997,N_11562);
and U12223 (N_12223,N_11753,N_11808);
or U12224 (N_12224,N_11792,N_11828);
nand U12225 (N_12225,N_11778,N_11699);
nand U12226 (N_12226,N_11855,N_11628);
nand U12227 (N_12227,N_11531,N_11648);
xnor U12228 (N_12228,N_11779,N_11726);
and U12229 (N_12229,N_11505,N_11559);
nor U12230 (N_12230,N_11676,N_11566);
xor U12231 (N_12231,N_11869,N_11526);
xor U12232 (N_12232,N_11708,N_11972);
nand U12233 (N_12233,N_11717,N_11705);
nand U12234 (N_12234,N_11558,N_11752);
xnor U12235 (N_12235,N_11657,N_11850);
or U12236 (N_12236,N_11659,N_11892);
nand U12237 (N_12237,N_11884,N_11848);
and U12238 (N_12238,N_11711,N_11801);
or U12239 (N_12239,N_11691,N_11906);
nor U12240 (N_12240,N_11740,N_11546);
nand U12241 (N_12241,N_11525,N_11888);
and U12242 (N_12242,N_11915,N_11654);
nand U12243 (N_12243,N_11707,N_11964);
nor U12244 (N_12244,N_11586,N_11980);
and U12245 (N_12245,N_11554,N_11935);
xor U12246 (N_12246,N_11576,N_11893);
or U12247 (N_12247,N_11510,N_11897);
or U12248 (N_12248,N_11990,N_11621);
xor U12249 (N_12249,N_11839,N_11655);
nor U12250 (N_12250,N_11619,N_11594);
nor U12251 (N_12251,N_11688,N_11525);
nor U12252 (N_12252,N_11602,N_11761);
nand U12253 (N_12253,N_11925,N_11638);
nor U12254 (N_12254,N_11710,N_11555);
nor U12255 (N_12255,N_11774,N_11667);
and U12256 (N_12256,N_11628,N_11695);
xor U12257 (N_12257,N_11757,N_11913);
nor U12258 (N_12258,N_11591,N_11876);
xnor U12259 (N_12259,N_11557,N_11950);
xnor U12260 (N_12260,N_11674,N_11658);
nand U12261 (N_12261,N_11824,N_11660);
or U12262 (N_12262,N_11760,N_11568);
xor U12263 (N_12263,N_11823,N_11780);
nand U12264 (N_12264,N_11675,N_11797);
nand U12265 (N_12265,N_11949,N_11731);
nor U12266 (N_12266,N_11883,N_11623);
or U12267 (N_12267,N_11563,N_11735);
nand U12268 (N_12268,N_11528,N_11770);
or U12269 (N_12269,N_11557,N_11877);
xnor U12270 (N_12270,N_11920,N_11881);
xor U12271 (N_12271,N_11925,N_11981);
nor U12272 (N_12272,N_11537,N_11996);
nor U12273 (N_12273,N_11861,N_11813);
or U12274 (N_12274,N_11674,N_11926);
nand U12275 (N_12275,N_11907,N_11709);
nand U12276 (N_12276,N_11899,N_11621);
or U12277 (N_12277,N_11858,N_11715);
and U12278 (N_12278,N_11958,N_11560);
nand U12279 (N_12279,N_11841,N_11996);
nand U12280 (N_12280,N_11993,N_11501);
and U12281 (N_12281,N_11662,N_11807);
xnor U12282 (N_12282,N_11692,N_11701);
and U12283 (N_12283,N_11906,N_11742);
or U12284 (N_12284,N_11819,N_11555);
nand U12285 (N_12285,N_11608,N_11862);
nand U12286 (N_12286,N_11942,N_11985);
nand U12287 (N_12287,N_11518,N_11764);
or U12288 (N_12288,N_11902,N_11924);
nor U12289 (N_12289,N_11540,N_11699);
and U12290 (N_12290,N_11695,N_11815);
and U12291 (N_12291,N_11739,N_11697);
nand U12292 (N_12292,N_11915,N_11622);
nor U12293 (N_12293,N_11863,N_11668);
xnor U12294 (N_12294,N_11590,N_11696);
or U12295 (N_12295,N_11655,N_11633);
or U12296 (N_12296,N_11743,N_11747);
nor U12297 (N_12297,N_11544,N_11581);
nand U12298 (N_12298,N_11585,N_11781);
and U12299 (N_12299,N_11510,N_11752);
xor U12300 (N_12300,N_11774,N_11894);
xor U12301 (N_12301,N_11621,N_11585);
nor U12302 (N_12302,N_11963,N_11758);
or U12303 (N_12303,N_11829,N_11642);
nand U12304 (N_12304,N_11578,N_11859);
xnor U12305 (N_12305,N_11772,N_11812);
or U12306 (N_12306,N_11809,N_11559);
or U12307 (N_12307,N_11837,N_11683);
and U12308 (N_12308,N_11816,N_11778);
nand U12309 (N_12309,N_11574,N_11911);
and U12310 (N_12310,N_11936,N_11806);
nand U12311 (N_12311,N_11835,N_11763);
and U12312 (N_12312,N_11949,N_11857);
nand U12313 (N_12313,N_11887,N_11745);
or U12314 (N_12314,N_11844,N_11569);
xor U12315 (N_12315,N_11604,N_11755);
and U12316 (N_12316,N_11685,N_11903);
and U12317 (N_12317,N_11782,N_11736);
nor U12318 (N_12318,N_11869,N_11598);
or U12319 (N_12319,N_11544,N_11977);
or U12320 (N_12320,N_11887,N_11786);
nor U12321 (N_12321,N_11763,N_11582);
nand U12322 (N_12322,N_11957,N_11509);
and U12323 (N_12323,N_11713,N_11597);
nand U12324 (N_12324,N_11922,N_11999);
and U12325 (N_12325,N_11633,N_11726);
nor U12326 (N_12326,N_11914,N_11655);
nand U12327 (N_12327,N_11926,N_11678);
nand U12328 (N_12328,N_11861,N_11666);
and U12329 (N_12329,N_11969,N_11689);
or U12330 (N_12330,N_11918,N_11692);
nor U12331 (N_12331,N_11714,N_11790);
and U12332 (N_12332,N_11926,N_11660);
nand U12333 (N_12333,N_11964,N_11774);
or U12334 (N_12334,N_11981,N_11733);
xor U12335 (N_12335,N_11953,N_11588);
and U12336 (N_12336,N_11696,N_11986);
or U12337 (N_12337,N_11661,N_11531);
nor U12338 (N_12338,N_11698,N_11667);
nor U12339 (N_12339,N_11774,N_11840);
nand U12340 (N_12340,N_11869,N_11769);
xnor U12341 (N_12341,N_11605,N_11802);
nand U12342 (N_12342,N_11938,N_11870);
or U12343 (N_12343,N_11969,N_11587);
or U12344 (N_12344,N_11839,N_11525);
or U12345 (N_12345,N_11589,N_11706);
nor U12346 (N_12346,N_11867,N_11520);
or U12347 (N_12347,N_11580,N_11624);
and U12348 (N_12348,N_11618,N_11780);
nand U12349 (N_12349,N_11869,N_11965);
and U12350 (N_12350,N_11789,N_11879);
or U12351 (N_12351,N_11954,N_11662);
nor U12352 (N_12352,N_11811,N_11744);
and U12353 (N_12353,N_11882,N_11937);
nand U12354 (N_12354,N_11713,N_11664);
and U12355 (N_12355,N_11905,N_11989);
nor U12356 (N_12356,N_11765,N_11793);
or U12357 (N_12357,N_11564,N_11957);
xnor U12358 (N_12358,N_11819,N_11855);
nor U12359 (N_12359,N_11694,N_11955);
xnor U12360 (N_12360,N_11575,N_11658);
and U12361 (N_12361,N_11531,N_11508);
or U12362 (N_12362,N_11955,N_11692);
and U12363 (N_12363,N_11693,N_11618);
nand U12364 (N_12364,N_11720,N_11684);
or U12365 (N_12365,N_11856,N_11661);
xor U12366 (N_12366,N_11744,N_11580);
and U12367 (N_12367,N_11604,N_11915);
nand U12368 (N_12368,N_11742,N_11945);
xnor U12369 (N_12369,N_11948,N_11524);
and U12370 (N_12370,N_11970,N_11728);
or U12371 (N_12371,N_11847,N_11548);
nand U12372 (N_12372,N_11825,N_11518);
and U12373 (N_12373,N_11832,N_11620);
or U12374 (N_12374,N_11802,N_11570);
or U12375 (N_12375,N_11898,N_11713);
nor U12376 (N_12376,N_11681,N_11501);
or U12377 (N_12377,N_11810,N_11595);
or U12378 (N_12378,N_11559,N_11889);
and U12379 (N_12379,N_11700,N_11852);
and U12380 (N_12380,N_11545,N_11678);
nor U12381 (N_12381,N_11780,N_11989);
nand U12382 (N_12382,N_11983,N_11524);
and U12383 (N_12383,N_11860,N_11740);
and U12384 (N_12384,N_11611,N_11618);
and U12385 (N_12385,N_11822,N_11535);
xnor U12386 (N_12386,N_11794,N_11779);
nor U12387 (N_12387,N_11851,N_11645);
nand U12388 (N_12388,N_11523,N_11658);
and U12389 (N_12389,N_11910,N_11648);
or U12390 (N_12390,N_11524,N_11954);
nand U12391 (N_12391,N_11737,N_11683);
xor U12392 (N_12392,N_11984,N_11543);
nor U12393 (N_12393,N_11667,N_11789);
nand U12394 (N_12394,N_11862,N_11649);
nand U12395 (N_12395,N_11917,N_11770);
and U12396 (N_12396,N_11961,N_11553);
nand U12397 (N_12397,N_11909,N_11936);
nand U12398 (N_12398,N_11641,N_11952);
nor U12399 (N_12399,N_11543,N_11570);
nand U12400 (N_12400,N_11840,N_11919);
or U12401 (N_12401,N_11649,N_11993);
nand U12402 (N_12402,N_11964,N_11818);
or U12403 (N_12403,N_11784,N_11985);
nor U12404 (N_12404,N_11863,N_11831);
nand U12405 (N_12405,N_11973,N_11980);
and U12406 (N_12406,N_11944,N_11844);
and U12407 (N_12407,N_11628,N_11858);
xnor U12408 (N_12408,N_11933,N_11850);
xnor U12409 (N_12409,N_11834,N_11519);
or U12410 (N_12410,N_11909,N_11550);
nor U12411 (N_12411,N_11857,N_11884);
and U12412 (N_12412,N_11904,N_11825);
nand U12413 (N_12413,N_11902,N_11741);
and U12414 (N_12414,N_11668,N_11888);
and U12415 (N_12415,N_11936,N_11865);
nor U12416 (N_12416,N_11820,N_11534);
nand U12417 (N_12417,N_11651,N_11927);
or U12418 (N_12418,N_11669,N_11724);
and U12419 (N_12419,N_11897,N_11547);
nand U12420 (N_12420,N_11853,N_11723);
nand U12421 (N_12421,N_11664,N_11827);
xnor U12422 (N_12422,N_11709,N_11666);
nor U12423 (N_12423,N_11693,N_11870);
nand U12424 (N_12424,N_11789,N_11747);
nand U12425 (N_12425,N_11745,N_11743);
nor U12426 (N_12426,N_11881,N_11802);
and U12427 (N_12427,N_11810,N_11633);
xnor U12428 (N_12428,N_11974,N_11663);
nor U12429 (N_12429,N_11972,N_11688);
or U12430 (N_12430,N_11553,N_11725);
and U12431 (N_12431,N_11842,N_11560);
and U12432 (N_12432,N_11943,N_11842);
xor U12433 (N_12433,N_11571,N_11786);
and U12434 (N_12434,N_11663,N_11653);
nor U12435 (N_12435,N_11684,N_11990);
nand U12436 (N_12436,N_11746,N_11703);
or U12437 (N_12437,N_11938,N_11710);
nand U12438 (N_12438,N_11646,N_11721);
nand U12439 (N_12439,N_11567,N_11940);
or U12440 (N_12440,N_11901,N_11932);
or U12441 (N_12441,N_11831,N_11781);
nor U12442 (N_12442,N_11534,N_11593);
xnor U12443 (N_12443,N_11713,N_11875);
nand U12444 (N_12444,N_11906,N_11637);
and U12445 (N_12445,N_11812,N_11749);
nor U12446 (N_12446,N_11777,N_11923);
and U12447 (N_12447,N_11509,N_11765);
nand U12448 (N_12448,N_11943,N_11503);
and U12449 (N_12449,N_11741,N_11543);
and U12450 (N_12450,N_11847,N_11994);
and U12451 (N_12451,N_11930,N_11929);
nand U12452 (N_12452,N_11859,N_11759);
nand U12453 (N_12453,N_11718,N_11532);
nor U12454 (N_12454,N_11847,N_11726);
xnor U12455 (N_12455,N_11933,N_11508);
or U12456 (N_12456,N_11950,N_11722);
xnor U12457 (N_12457,N_11674,N_11673);
and U12458 (N_12458,N_11556,N_11546);
xor U12459 (N_12459,N_11761,N_11624);
or U12460 (N_12460,N_11669,N_11599);
nand U12461 (N_12461,N_11545,N_11705);
or U12462 (N_12462,N_11947,N_11588);
and U12463 (N_12463,N_11734,N_11820);
nor U12464 (N_12464,N_11824,N_11730);
or U12465 (N_12465,N_11563,N_11524);
nand U12466 (N_12466,N_11510,N_11598);
and U12467 (N_12467,N_11811,N_11891);
or U12468 (N_12468,N_11637,N_11792);
nor U12469 (N_12469,N_11801,N_11575);
and U12470 (N_12470,N_11663,N_11681);
and U12471 (N_12471,N_11843,N_11894);
or U12472 (N_12472,N_11684,N_11674);
nand U12473 (N_12473,N_11529,N_11946);
nand U12474 (N_12474,N_11896,N_11579);
xor U12475 (N_12475,N_11503,N_11546);
and U12476 (N_12476,N_11673,N_11612);
xnor U12477 (N_12477,N_11773,N_11933);
nor U12478 (N_12478,N_11836,N_11669);
and U12479 (N_12479,N_11602,N_11959);
or U12480 (N_12480,N_11937,N_11679);
or U12481 (N_12481,N_11655,N_11738);
or U12482 (N_12482,N_11828,N_11924);
or U12483 (N_12483,N_11687,N_11934);
nand U12484 (N_12484,N_11628,N_11847);
and U12485 (N_12485,N_11503,N_11838);
nor U12486 (N_12486,N_11833,N_11728);
nand U12487 (N_12487,N_11981,N_11861);
xor U12488 (N_12488,N_11755,N_11660);
xor U12489 (N_12489,N_11784,N_11801);
nor U12490 (N_12490,N_11664,N_11732);
and U12491 (N_12491,N_11575,N_11977);
xnor U12492 (N_12492,N_11573,N_11798);
and U12493 (N_12493,N_11526,N_11712);
nor U12494 (N_12494,N_11756,N_11827);
or U12495 (N_12495,N_11651,N_11674);
nor U12496 (N_12496,N_11558,N_11747);
and U12497 (N_12497,N_11777,N_11716);
xnor U12498 (N_12498,N_11714,N_11722);
and U12499 (N_12499,N_11815,N_11509);
or U12500 (N_12500,N_12143,N_12258);
or U12501 (N_12501,N_12030,N_12448);
nand U12502 (N_12502,N_12227,N_12126);
nand U12503 (N_12503,N_12025,N_12314);
and U12504 (N_12504,N_12406,N_12272);
and U12505 (N_12505,N_12260,N_12097);
and U12506 (N_12506,N_12400,N_12079);
and U12507 (N_12507,N_12273,N_12212);
xor U12508 (N_12508,N_12282,N_12311);
or U12509 (N_12509,N_12175,N_12007);
xor U12510 (N_12510,N_12027,N_12120);
and U12511 (N_12511,N_12267,N_12067);
and U12512 (N_12512,N_12413,N_12432);
xnor U12513 (N_12513,N_12125,N_12106);
nor U12514 (N_12514,N_12425,N_12041);
xnor U12515 (N_12515,N_12024,N_12317);
nor U12516 (N_12516,N_12006,N_12467);
xor U12517 (N_12517,N_12357,N_12478);
and U12518 (N_12518,N_12042,N_12394);
nand U12519 (N_12519,N_12354,N_12355);
xnor U12520 (N_12520,N_12065,N_12466);
and U12521 (N_12521,N_12319,N_12134);
and U12522 (N_12522,N_12472,N_12276);
or U12523 (N_12523,N_12207,N_12421);
nor U12524 (N_12524,N_12455,N_12071);
nor U12525 (N_12525,N_12312,N_12076);
nor U12526 (N_12526,N_12442,N_12160);
or U12527 (N_12527,N_12046,N_12462);
or U12528 (N_12528,N_12458,N_12476);
and U12529 (N_12529,N_12254,N_12320);
nand U12530 (N_12530,N_12374,N_12147);
nand U12531 (N_12531,N_12220,N_12165);
nand U12532 (N_12532,N_12404,N_12014);
and U12533 (N_12533,N_12446,N_12137);
or U12534 (N_12534,N_12218,N_12345);
and U12535 (N_12535,N_12062,N_12297);
or U12536 (N_12536,N_12149,N_12280);
or U12537 (N_12537,N_12492,N_12367);
nor U12538 (N_12538,N_12241,N_12139);
or U12539 (N_12539,N_12038,N_12373);
nand U12540 (N_12540,N_12410,N_12248);
xnor U12541 (N_12541,N_12082,N_12154);
and U12542 (N_12542,N_12135,N_12368);
or U12543 (N_12543,N_12295,N_12371);
and U12544 (N_12544,N_12127,N_12415);
and U12545 (N_12545,N_12411,N_12454);
or U12546 (N_12546,N_12145,N_12018);
or U12547 (N_12547,N_12200,N_12161);
nor U12548 (N_12548,N_12464,N_12190);
and U12549 (N_12549,N_12337,N_12453);
or U12550 (N_12550,N_12482,N_12329);
nand U12551 (N_12551,N_12445,N_12477);
nand U12552 (N_12552,N_12348,N_12238);
nand U12553 (N_12553,N_12262,N_12128);
or U12554 (N_12554,N_12296,N_12031);
and U12555 (N_12555,N_12063,N_12349);
and U12556 (N_12556,N_12179,N_12269);
nand U12557 (N_12557,N_12109,N_12118);
xnor U12558 (N_12558,N_12047,N_12117);
xor U12559 (N_12559,N_12049,N_12204);
xor U12560 (N_12560,N_12486,N_12235);
or U12561 (N_12561,N_12231,N_12197);
and U12562 (N_12562,N_12393,N_12085);
xor U12563 (N_12563,N_12483,N_12140);
and U12564 (N_12564,N_12073,N_12004);
and U12565 (N_12565,N_12418,N_12171);
nand U12566 (N_12566,N_12327,N_12096);
xnor U12567 (N_12567,N_12121,N_12334);
nand U12568 (N_12568,N_12189,N_12158);
nor U12569 (N_12569,N_12017,N_12495);
nand U12570 (N_12570,N_12366,N_12084);
nand U12571 (N_12571,N_12424,N_12275);
nand U12572 (N_12572,N_12463,N_12291);
xnor U12573 (N_12573,N_12219,N_12229);
nor U12574 (N_12574,N_12182,N_12383);
nand U12575 (N_12575,N_12287,N_12301);
nor U12576 (N_12576,N_12428,N_12470);
nand U12577 (N_12577,N_12068,N_12114);
and U12578 (N_12578,N_12362,N_12372);
nor U12579 (N_12579,N_12378,N_12289);
nor U12580 (N_12580,N_12426,N_12285);
nor U12581 (N_12581,N_12261,N_12361);
nand U12582 (N_12582,N_12060,N_12377);
nor U12583 (N_12583,N_12330,N_12083);
nand U12584 (N_12584,N_12225,N_12045);
nand U12585 (N_12585,N_12256,N_12089);
nand U12586 (N_12586,N_12387,N_12019);
nor U12587 (N_12587,N_12176,N_12304);
and U12588 (N_12588,N_12369,N_12166);
or U12589 (N_12589,N_12222,N_12493);
xnor U12590 (N_12590,N_12288,N_12039);
nand U12591 (N_12591,N_12412,N_12474);
xnor U12592 (N_12592,N_12444,N_12066);
and U12593 (N_12593,N_12257,N_12048);
xor U12594 (N_12594,N_12036,N_12405);
xor U12595 (N_12595,N_12051,N_12469);
xor U12596 (N_12596,N_12102,N_12423);
xor U12597 (N_12597,N_12250,N_12447);
or U12598 (N_12598,N_12278,N_12064);
or U12599 (N_12599,N_12279,N_12183);
xnor U12600 (N_12600,N_12116,N_12211);
xnor U12601 (N_12601,N_12026,N_12359);
nor U12602 (N_12602,N_12223,N_12136);
nor U12603 (N_12603,N_12274,N_12335);
nor U12604 (N_12604,N_12015,N_12035);
or U12605 (N_12605,N_12033,N_12012);
and U12606 (N_12606,N_12325,N_12239);
or U12607 (N_12607,N_12001,N_12437);
or U12608 (N_12608,N_12452,N_12247);
xnor U12609 (N_12609,N_12379,N_12298);
nor U12610 (N_12610,N_12217,N_12305);
nand U12611 (N_12611,N_12230,N_12431);
and U12612 (N_12612,N_12091,N_12214);
and U12613 (N_12613,N_12193,N_12259);
xor U12614 (N_12614,N_12105,N_12384);
nand U12615 (N_12615,N_12005,N_12115);
nor U12616 (N_12616,N_12224,N_12321);
xor U12617 (N_12617,N_12306,N_12093);
nand U12618 (N_12618,N_12110,N_12443);
or U12619 (N_12619,N_12456,N_12098);
nor U12620 (N_12620,N_12465,N_12205);
nor U12621 (N_12621,N_12440,N_12132);
or U12622 (N_12622,N_12020,N_12040);
or U12623 (N_12623,N_12226,N_12055);
xor U12624 (N_12624,N_12313,N_12107);
nor U12625 (N_12625,N_12496,N_12497);
nor U12626 (N_12626,N_12174,N_12403);
xnor U12627 (N_12627,N_12034,N_12308);
xor U12628 (N_12628,N_12188,N_12087);
or U12629 (N_12629,N_12186,N_12245);
nand U12630 (N_12630,N_12092,N_12363);
or U12631 (N_12631,N_12032,N_12488);
nor U12632 (N_12632,N_12309,N_12056);
and U12633 (N_12633,N_12003,N_12080);
and U12634 (N_12634,N_12167,N_12339);
nor U12635 (N_12635,N_12170,N_12449);
or U12636 (N_12636,N_12209,N_12459);
nand U12637 (N_12637,N_12471,N_12481);
nor U12638 (N_12638,N_12061,N_12353);
or U12639 (N_12639,N_12142,N_12475);
or U12640 (N_12640,N_12100,N_12251);
or U12641 (N_12641,N_12324,N_12169);
or U12642 (N_12642,N_12294,N_12385);
nor U12643 (N_12643,N_12008,N_12499);
and U12644 (N_12644,N_12156,N_12441);
xnor U12645 (N_12645,N_12323,N_12131);
and U12646 (N_12646,N_12479,N_12058);
and U12647 (N_12647,N_12162,N_12419);
nor U12648 (N_12648,N_12152,N_12172);
and U12649 (N_12649,N_12489,N_12293);
xnor U12650 (N_12650,N_12234,N_12151);
nor U12651 (N_12651,N_12316,N_12029);
or U12652 (N_12652,N_12157,N_12494);
xnor U12653 (N_12653,N_12081,N_12168);
nor U12654 (N_12654,N_12233,N_12215);
nand U12655 (N_12655,N_12144,N_12360);
or U12656 (N_12656,N_12221,N_12101);
and U12657 (N_12657,N_12281,N_12146);
or U12658 (N_12658,N_12427,N_12201);
nor U12659 (N_12659,N_12375,N_12074);
xnor U12660 (N_12660,N_12263,N_12202);
nor U12661 (N_12661,N_12347,N_12053);
and U12662 (N_12662,N_12075,N_12194);
xnor U12663 (N_12663,N_12302,N_12216);
nand U12664 (N_12664,N_12113,N_12398);
nand U12665 (N_12665,N_12232,N_12228);
xor U12666 (N_12666,N_12346,N_12000);
nor U12667 (N_12667,N_12210,N_12178);
or U12668 (N_12668,N_12416,N_12255);
and U12669 (N_12669,N_12198,N_12365);
and U12670 (N_12670,N_12420,N_12159);
nor U12671 (N_12671,N_12090,N_12252);
nor U12672 (N_12672,N_12155,N_12244);
or U12673 (N_12673,N_12358,N_12356);
or U12674 (N_12674,N_12206,N_12195);
xor U12675 (N_12675,N_12342,N_12108);
nand U12676 (N_12676,N_12173,N_12484);
and U12677 (N_12677,N_12380,N_12208);
nand U12678 (N_12678,N_12119,N_12480);
nor U12679 (N_12679,N_12266,N_12338);
xor U12680 (N_12680,N_12103,N_12290);
xor U12681 (N_12681,N_12264,N_12433);
nor U12682 (N_12682,N_12111,N_12435);
and U12683 (N_12683,N_12485,N_12336);
xor U12684 (N_12684,N_12299,N_12043);
nor U12685 (N_12685,N_12180,N_12016);
xnor U12686 (N_12686,N_12328,N_12088);
xor U12687 (N_12687,N_12271,N_12303);
or U12688 (N_12688,N_12277,N_12364);
and U12689 (N_12689,N_12392,N_12122);
nand U12690 (N_12690,N_12468,N_12191);
xnor U12691 (N_12691,N_12010,N_12307);
nor U12692 (N_12692,N_12099,N_12023);
nand U12693 (N_12693,N_12213,N_12331);
xnor U12694 (N_12694,N_12397,N_12370);
nor U12695 (N_12695,N_12237,N_12414);
nand U12696 (N_12696,N_12242,N_12395);
nand U12697 (N_12697,N_12112,N_12133);
or U12698 (N_12698,N_12070,N_12086);
nor U12699 (N_12699,N_12333,N_12382);
nand U12700 (N_12700,N_12268,N_12192);
nand U12701 (N_12701,N_12434,N_12284);
or U12702 (N_12702,N_12438,N_12332);
or U12703 (N_12703,N_12401,N_12402);
and U12704 (N_12704,N_12141,N_12203);
nor U12705 (N_12705,N_12351,N_12177);
xor U12706 (N_12706,N_12148,N_12386);
or U12707 (N_12707,N_12490,N_12450);
nand U12708 (N_12708,N_12407,N_12391);
xnor U12709 (N_12709,N_12315,N_12199);
nand U12710 (N_12710,N_12072,N_12164);
nor U12711 (N_12711,N_12002,N_12184);
xnor U12712 (N_12712,N_12451,N_12078);
xor U12713 (N_12713,N_12069,N_12491);
and U12714 (N_12714,N_12376,N_12181);
and U12715 (N_12715,N_12300,N_12094);
or U12716 (N_12716,N_12352,N_12283);
nand U12717 (N_12717,N_12326,N_12399);
and U12718 (N_12718,N_12292,N_12422);
nand U12719 (N_12719,N_12059,N_12388);
xnor U12720 (N_12720,N_12461,N_12341);
and U12721 (N_12721,N_12163,N_12270);
nand U12722 (N_12722,N_12350,N_12022);
xnor U12723 (N_12723,N_12129,N_12021);
xor U12724 (N_12724,N_12011,N_12430);
nand U12725 (N_12725,N_12104,N_12286);
xor U12726 (N_12726,N_12246,N_12498);
nor U12727 (N_12727,N_12381,N_12028);
nand U12728 (N_12728,N_12473,N_12153);
nor U12729 (N_12729,N_12408,N_12318);
nor U12730 (N_12730,N_12130,N_12409);
xnor U12731 (N_12731,N_12460,N_12052);
xnor U12732 (N_12732,N_12044,N_12123);
nor U12733 (N_12733,N_12196,N_12396);
or U12734 (N_12734,N_12138,N_12344);
nor U12735 (N_12735,N_12249,N_12037);
or U12736 (N_12736,N_12310,N_12265);
xor U12737 (N_12737,N_12150,N_12057);
and U12738 (N_12738,N_12187,N_12390);
and U12739 (N_12739,N_12124,N_12389);
xor U12740 (N_12740,N_12343,N_12077);
nand U12741 (N_12741,N_12185,N_12436);
nand U12742 (N_12742,N_12013,N_12253);
and U12743 (N_12743,N_12054,N_12417);
nor U12744 (N_12744,N_12243,N_12095);
or U12745 (N_12745,N_12439,N_12050);
xnor U12746 (N_12746,N_12322,N_12429);
or U12747 (N_12747,N_12340,N_12009);
nand U12748 (N_12748,N_12240,N_12457);
and U12749 (N_12749,N_12236,N_12487);
nor U12750 (N_12750,N_12213,N_12373);
and U12751 (N_12751,N_12039,N_12497);
xnor U12752 (N_12752,N_12290,N_12344);
nor U12753 (N_12753,N_12151,N_12455);
and U12754 (N_12754,N_12371,N_12165);
and U12755 (N_12755,N_12182,N_12130);
xor U12756 (N_12756,N_12487,N_12335);
and U12757 (N_12757,N_12092,N_12196);
nor U12758 (N_12758,N_12221,N_12105);
nand U12759 (N_12759,N_12261,N_12244);
nand U12760 (N_12760,N_12115,N_12022);
nand U12761 (N_12761,N_12093,N_12011);
nand U12762 (N_12762,N_12179,N_12283);
nor U12763 (N_12763,N_12337,N_12273);
nor U12764 (N_12764,N_12356,N_12077);
nor U12765 (N_12765,N_12412,N_12011);
nor U12766 (N_12766,N_12386,N_12137);
xor U12767 (N_12767,N_12002,N_12349);
nor U12768 (N_12768,N_12470,N_12129);
xnor U12769 (N_12769,N_12273,N_12285);
nor U12770 (N_12770,N_12324,N_12269);
nor U12771 (N_12771,N_12274,N_12311);
nor U12772 (N_12772,N_12051,N_12389);
xnor U12773 (N_12773,N_12471,N_12096);
xnor U12774 (N_12774,N_12421,N_12060);
or U12775 (N_12775,N_12125,N_12351);
xor U12776 (N_12776,N_12188,N_12133);
or U12777 (N_12777,N_12322,N_12068);
or U12778 (N_12778,N_12212,N_12344);
and U12779 (N_12779,N_12339,N_12110);
nor U12780 (N_12780,N_12219,N_12178);
xnor U12781 (N_12781,N_12116,N_12365);
xnor U12782 (N_12782,N_12318,N_12370);
and U12783 (N_12783,N_12101,N_12035);
nand U12784 (N_12784,N_12442,N_12045);
xnor U12785 (N_12785,N_12362,N_12156);
or U12786 (N_12786,N_12141,N_12407);
nor U12787 (N_12787,N_12213,N_12232);
nor U12788 (N_12788,N_12402,N_12097);
or U12789 (N_12789,N_12137,N_12159);
xnor U12790 (N_12790,N_12218,N_12055);
nor U12791 (N_12791,N_12099,N_12331);
or U12792 (N_12792,N_12377,N_12132);
and U12793 (N_12793,N_12201,N_12247);
nand U12794 (N_12794,N_12022,N_12436);
and U12795 (N_12795,N_12067,N_12131);
nand U12796 (N_12796,N_12115,N_12271);
or U12797 (N_12797,N_12099,N_12219);
xor U12798 (N_12798,N_12165,N_12000);
or U12799 (N_12799,N_12473,N_12305);
and U12800 (N_12800,N_12039,N_12131);
or U12801 (N_12801,N_12014,N_12423);
xor U12802 (N_12802,N_12357,N_12115);
xnor U12803 (N_12803,N_12208,N_12098);
or U12804 (N_12804,N_12418,N_12040);
nand U12805 (N_12805,N_12405,N_12031);
nor U12806 (N_12806,N_12488,N_12295);
and U12807 (N_12807,N_12056,N_12489);
and U12808 (N_12808,N_12315,N_12062);
and U12809 (N_12809,N_12106,N_12164);
or U12810 (N_12810,N_12269,N_12406);
and U12811 (N_12811,N_12079,N_12258);
xor U12812 (N_12812,N_12012,N_12300);
and U12813 (N_12813,N_12048,N_12151);
and U12814 (N_12814,N_12200,N_12118);
nand U12815 (N_12815,N_12195,N_12354);
xnor U12816 (N_12816,N_12272,N_12447);
xnor U12817 (N_12817,N_12070,N_12198);
and U12818 (N_12818,N_12054,N_12372);
nand U12819 (N_12819,N_12365,N_12357);
or U12820 (N_12820,N_12335,N_12046);
xnor U12821 (N_12821,N_12485,N_12386);
nand U12822 (N_12822,N_12006,N_12482);
or U12823 (N_12823,N_12077,N_12100);
or U12824 (N_12824,N_12385,N_12433);
nand U12825 (N_12825,N_12378,N_12102);
and U12826 (N_12826,N_12429,N_12455);
or U12827 (N_12827,N_12108,N_12308);
or U12828 (N_12828,N_12118,N_12306);
and U12829 (N_12829,N_12238,N_12058);
nand U12830 (N_12830,N_12094,N_12329);
nor U12831 (N_12831,N_12290,N_12164);
nand U12832 (N_12832,N_12290,N_12001);
and U12833 (N_12833,N_12332,N_12030);
xor U12834 (N_12834,N_12479,N_12397);
nand U12835 (N_12835,N_12369,N_12083);
xor U12836 (N_12836,N_12173,N_12322);
nor U12837 (N_12837,N_12493,N_12481);
xnor U12838 (N_12838,N_12355,N_12046);
and U12839 (N_12839,N_12180,N_12149);
nor U12840 (N_12840,N_12295,N_12127);
or U12841 (N_12841,N_12066,N_12166);
nand U12842 (N_12842,N_12346,N_12126);
and U12843 (N_12843,N_12154,N_12244);
or U12844 (N_12844,N_12098,N_12073);
nor U12845 (N_12845,N_12386,N_12254);
nor U12846 (N_12846,N_12409,N_12087);
or U12847 (N_12847,N_12495,N_12153);
nor U12848 (N_12848,N_12189,N_12081);
xor U12849 (N_12849,N_12223,N_12313);
nor U12850 (N_12850,N_12214,N_12184);
and U12851 (N_12851,N_12005,N_12415);
xnor U12852 (N_12852,N_12329,N_12398);
and U12853 (N_12853,N_12051,N_12397);
nor U12854 (N_12854,N_12339,N_12200);
or U12855 (N_12855,N_12238,N_12207);
and U12856 (N_12856,N_12153,N_12302);
and U12857 (N_12857,N_12114,N_12041);
nor U12858 (N_12858,N_12379,N_12218);
or U12859 (N_12859,N_12395,N_12340);
nand U12860 (N_12860,N_12006,N_12315);
or U12861 (N_12861,N_12100,N_12465);
or U12862 (N_12862,N_12053,N_12461);
nand U12863 (N_12863,N_12021,N_12451);
xor U12864 (N_12864,N_12099,N_12334);
nor U12865 (N_12865,N_12359,N_12079);
or U12866 (N_12866,N_12084,N_12025);
and U12867 (N_12867,N_12285,N_12145);
or U12868 (N_12868,N_12107,N_12456);
or U12869 (N_12869,N_12161,N_12085);
nand U12870 (N_12870,N_12494,N_12134);
nor U12871 (N_12871,N_12161,N_12066);
nor U12872 (N_12872,N_12263,N_12037);
xor U12873 (N_12873,N_12387,N_12196);
and U12874 (N_12874,N_12428,N_12388);
nor U12875 (N_12875,N_12122,N_12398);
nor U12876 (N_12876,N_12213,N_12491);
nand U12877 (N_12877,N_12063,N_12470);
nand U12878 (N_12878,N_12111,N_12190);
nand U12879 (N_12879,N_12447,N_12327);
and U12880 (N_12880,N_12445,N_12032);
xor U12881 (N_12881,N_12083,N_12096);
xnor U12882 (N_12882,N_12109,N_12319);
nor U12883 (N_12883,N_12467,N_12056);
nand U12884 (N_12884,N_12395,N_12167);
and U12885 (N_12885,N_12116,N_12179);
nor U12886 (N_12886,N_12247,N_12213);
nor U12887 (N_12887,N_12051,N_12327);
or U12888 (N_12888,N_12282,N_12445);
and U12889 (N_12889,N_12357,N_12382);
nand U12890 (N_12890,N_12272,N_12219);
and U12891 (N_12891,N_12170,N_12048);
and U12892 (N_12892,N_12005,N_12166);
and U12893 (N_12893,N_12471,N_12354);
and U12894 (N_12894,N_12193,N_12188);
and U12895 (N_12895,N_12025,N_12217);
nand U12896 (N_12896,N_12250,N_12340);
nand U12897 (N_12897,N_12406,N_12264);
nor U12898 (N_12898,N_12196,N_12119);
nor U12899 (N_12899,N_12247,N_12263);
nor U12900 (N_12900,N_12337,N_12049);
or U12901 (N_12901,N_12424,N_12409);
xnor U12902 (N_12902,N_12145,N_12294);
or U12903 (N_12903,N_12409,N_12447);
and U12904 (N_12904,N_12254,N_12143);
nor U12905 (N_12905,N_12387,N_12310);
nor U12906 (N_12906,N_12359,N_12415);
and U12907 (N_12907,N_12424,N_12139);
or U12908 (N_12908,N_12466,N_12181);
nand U12909 (N_12909,N_12233,N_12364);
or U12910 (N_12910,N_12380,N_12423);
xnor U12911 (N_12911,N_12295,N_12399);
nand U12912 (N_12912,N_12033,N_12353);
and U12913 (N_12913,N_12274,N_12455);
nand U12914 (N_12914,N_12005,N_12386);
and U12915 (N_12915,N_12095,N_12258);
xor U12916 (N_12916,N_12328,N_12112);
nand U12917 (N_12917,N_12422,N_12262);
nand U12918 (N_12918,N_12136,N_12499);
nand U12919 (N_12919,N_12373,N_12044);
nor U12920 (N_12920,N_12231,N_12087);
nor U12921 (N_12921,N_12083,N_12062);
or U12922 (N_12922,N_12483,N_12418);
and U12923 (N_12923,N_12005,N_12436);
or U12924 (N_12924,N_12220,N_12306);
nor U12925 (N_12925,N_12213,N_12318);
nand U12926 (N_12926,N_12189,N_12186);
nor U12927 (N_12927,N_12261,N_12056);
xor U12928 (N_12928,N_12061,N_12257);
and U12929 (N_12929,N_12348,N_12159);
nor U12930 (N_12930,N_12396,N_12003);
or U12931 (N_12931,N_12390,N_12389);
xor U12932 (N_12932,N_12149,N_12148);
or U12933 (N_12933,N_12344,N_12403);
or U12934 (N_12934,N_12221,N_12055);
and U12935 (N_12935,N_12133,N_12306);
nand U12936 (N_12936,N_12226,N_12447);
or U12937 (N_12937,N_12098,N_12296);
nor U12938 (N_12938,N_12277,N_12492);
nor U12939 (N_12939,N_12246,N_12040);
nor U12940 (N_12940,N_12211,N_12391);
xnor U12941 (N_12941,N_12123,N_12041);
nor U12942 (N_12942,N_12230,N_12193);
and U12943 (N_12943,N_12380,N_12063);
and U12944 (N_12944,N_12304,N_12354);
nor U12945 (N_12945,N_12008,N_12316);
xnor U12946 (N_12946,N_12018,N_12219);
or U12947 (N_12947,N_12052,N_12226);
nand U12948 (N_12948,N_12071,N_12485);
nand U12949 (N_12949,N_12064,N_12444);
and U12950 (N_12950,N_12050,N_12311);
and U12951 (N_12951,N_12244,N_12307);
nor U12952 (N_12952,N_12121,N_12394);
nand U12953 (N_12953,N_12048,N_12037);
nor U12954 (N_12954,N_12386,N_12294);
or U12955 (N_12955,N_12256,N_12189);
nor U12956 (N_12956,N_12196,N_12030);
xor U12957 (N_12957,N_12045,N_12283);
nand U12958 (N_12958,N_12460,N_12394);
nand U12959 (N_12959,N_12411,N_12027);
xnor U12960 (N_12960,N_12331,N_12069);
nor U12961 (N_12961,N_12209,N_12162);
nor U12962 (N_12962,N_12486,N_12187);
nor U12963 (N_12963,N_12162,N_12233);
xor U12964 (N_12964,N_12416,N_12345);
xor U12965 (N_12965,N_12016,N_12339);
nor U12966 (N_12966,N_12491,N_12338);
nand U12967 (N_12967,N_12266,N_12032);
and U12968 (N_12968,N_12205,N_12183);
nand U12969 (N_12969,N_12213,N_12107);
and U12970 (N_12970,N_12332,N_12267);
xnor U12971 (N_12971,N_12078,N_12390);
nor U12972 (N_12972,N_12353,N_12137);
nand U12973 (N_12973,N_12317,N_12115);
or U12974 (N_12974,N_12404,N_12395);
and U12975 (N_12975,N_12069,N_12043);
xnor U12976 (N_12976,N_12345,N_12374);
or U12977 (N_12977,N_12270,N_12306);
xor U12978 (N_12978,N_12211,N_12128);
nor U12979 (N_12979,N_12317,N_12061);
and U12980 (N_12980,N_12337,N_12335);
nand U12981 (N_12981,N_12170,N_12216);
nor U12982 (N_12982,N_12494,N_12182);
or U12983 (N_12983,N_12029,N_12460);
nor U12984 (N_12984,N_12418,N_12220);
nor U12985 (N_12985,N_12082,N_12387);
nand U12986 (N_12986,N_12362,N_12435);
xnor U12987 (N_12987,N_12355,N_12161);
nor U12988 (N_12988,N_12342,N_12199);
nand U12989 (N_12989,N_12006,N_12139);
nand U12990 (N_12990,N_12071,N_12038);
nor U12991 (N_12991,N_12108,N_12358);
xor U12992 (N_12992,N_12174,N_12106);
nand U12993 (N_12993,N_12250,N_12327);
or U12994 (N_12994,N_12155,N_12091);
or U12995 (N_12995,N_12132,N_12250);
nand U12996 (N_12996,N_12299,N_12357);
nor U12997 (N_12997,N_12269,N_12055);
nand U12998 (N_12998,N_12046,N_12180);
or U12999 (N_12999,N_12043,N_12137);
nor U13000 (N_13000,N_12512,N_12606);
xor U13001 (N_13001,N_12833,N_12838);
xnor U13002 (N_13002,N_12585,N_12636);
xnor U13003 (N_13003,N_12962,N_12748);
xnor U13004 (N_13004,N_12506,N_12642);
or U13005 (N_13005,N_12968,N_12873);
nand U13006 (N_13006,N_12563,N_12657);
nor U13007 (N_13007,N_12683,N_12567);
xor U13008 (N_13008,N_12956,N_12644);
xor U13009 (N_13009,N_12519,N_12868);
or U13010 (N_13010,N_12888,N_12869);
nor U13011 (N_13011,N_12635,N_12861);
xor U13012 (N_13012,N_12762,N_12942);
xor U13013 (N_13013,N_12536,N_12661);
nor U13014 (N_13014,N_12617,N_12784);
xor U13015 (N_13015,N_12953,N_12676);
or U13016 (N_13016,N_12907,N_12716);
nor U13017 (N_13017,N_12863,N_12745);
nand U13018 (N_13018,N_12930,N_12874);
nand U13019 (N_13019,N_12774,N_12997);
nand U13020 (N_13020,N_12562,N_12847);
xor U13021 (N_13021,N_12523,N_12651);
nand U13022 (N_13022,N_12742,N_12602);
nand U13023 (N_13023,N_12925,N_12828);
nand U13024 (N_13024,N_12990,N_12744);
nor U13025 (N_13025,N_12928,N_12500);
nand U13026 (N_13026,N_12998,N_12949);
nand U13027 (N_13027,N_12741,N_12731);
or U13028 (N_13028,N_12937,N_12668);
nor U13029 (N_13029,N_12913,N_12779);
xor U13030 (N_13030,N_12950,N_12595);
or U13031 (N_13031,N_12687,N_12896);
and U13032 (N_13032,N_12502,N_12673);
or U13033 (N_13033,N_12877,N_12872);
nor U13034 (N_13034,N_12870,N_12836);
nand U13035 (N_13035,N_12556,N_12507);
and U13036 (N_13036,N_12715,N_12920);
nor U13037 (N_13037,N_12705,N_12750);
or U13038 (N_13038,N_12826,N_12540);
nor U13039 (N_13039,N_12631,N_12797);
nor U13040 (N_13040,N_12926,N_12577);
or U13041 (N_13041,N_12856,N_12952);
nor U13042 (N_13042,N_12575,N_12746);
or U13043 (N_13043,N_12692,N_12627);
xnor U13044 (N_13044,N_12591,N_12660);
nand U13045 (N_13045,N_12646,N_12876);
nand U13046 (N_13046,N_12558,N_12701);
or U13047 (N_13047,N_12560,N_12520);
and U13048 (N_13048,N_12600,N_12882);
nor U13049 (N_13049,N_12948,N_12807);
xnor U13050 (N_13050,N_12666,N_12695);
or U13051 (N_13051,N_12800,N_12781);
xor U13052 (N_13052,N_12840,N_12685);
nor U13053 (N_13053,N_12813,N_12670);
or U13054 (N_13054,N_12770,N_12794);
or U13055 (N_13055,N_12923,N_12945);
or U13056 (N_13056,N_12915,N_12572);
nand U13057 (N_13057,N_12772,N_12921);
xnor U13058 (N_13058,N_12663,N_12897);
nor U13059 (N_13059,N_12712,N_12706);
and U13060 (N_13060,N_12700,N_12974);
nor U13061 (N_13061,N_12973,N_12835);
nor U13062 (N_13062,N_12552,N_12658);
or U13063 (N_13063,N_12656,N_12529);
or U13064 (N_13064,N_12851,N_12761);
nand U13065 (N_13065,N_12621,N_12751);
nor U13066 (N_13066,N_12539,N_12980);
or U13067 (N_13067,N_12778,N_12736);
and U13068 (N_13068,N_12576,N_12830);
nor U13069 (N_13069,N_12822,N_12559);
or U13070 (N_13070,N_12738,N_12739);
and U13071 (N_13071,N_12879,N_12769);
nand U13072 (N_13072,N_12853,N_12790);
xnor U13073 (N_13073,N_12679,N_12903);
nor U13074 (N_13074,N_12932,N_12553);
xor U13075 (N_13075,N_12721,N_12777);
and U13076 (N_13076,N_12538,N_12796);
or U13077 (N_13077,N_12773,N_12598);
nor U13078 (N_13078,N_12625,N_12672);
nor U13079 (N_13079,N_12812,N_12682);
nand U13080 (N_13080,N_12688,N_12846);
nor U13081 (N_13081,N_12987,N_12768);
and U13082 (N_13082,N_12588,N_12501);
or U13083 (N_13083,N_12880,N_12837);
nand U13084 (N_13084,N_12541,N_12983);
nand U13085 (N_13085,N_12916,N_12671);
xnor U13086 (N_13086,N_12816,N_12509);
nor U13087 (N_13087,N_12629,N_12940);
and U13088 (N_13088,N_12589,N_12609);
or U13089 (N_13089,N_12811,N_12714);
xnor U13090 (N_13090,N_12544,N_12664);
and U13091 (N_13091,N_12568,N_12722);
or U13092 (N_13092,N_12537,N_12817);
or U13093 (N_13093,N_12678,N_12970);
and U13094 (N_13094,N_12845,N_12723);
nor U13095 (N_13095,N_12887,N_12667);
nor U13096 (N_13096,N_12883,N_12735);
and U13097 (N_13097,N_12809,N_12599);
nor U13098 (N_13098,N_12675,N_12571);
xor U13099 (N_13099,N_12546,N_12699);
nand U13100 (N_13100,N_12910,N_12999);
and U13101 (N_13101,N_12641,N_12788);
and U13102 (N_13102,N_12726,N_12960);
nor U13103 (N_13103,N_12659,N_12728);
xor U13104 (N_13104,N_12614,N_12711);
or U13105 (N_13105,N_12704,N_12972);
nor U13106 (N_13106,N_12593,N_12531);
nor U13107 (N_13107,N_12775,N_12943);
nor U13108 (N_13108,N_12977,N_12582);
xor U13109 (N_13109,N_12993,N_12724);
or U13110 (N_13110,N_12505,N_12867);
and U13111 (N_13111,N_12801,N_12765);
or U13112 (N_13112,N_12933,N_12766);
xor U13113 (N_13113,N_12628,N_12843);
nor U13114 (N_13114,N_12527,N_12815);
nor U13115 (N_13115,N_12583,N_12782);
or U13116 (N_13116,N_12607,N_12601);
and U13117 (N_13117,N_12908,N_12548);
and U13118 (N_13118,N_12992,N_12767);
nor U13119 (N_13119,N_12821,N_12639);
nor U13120 (N_13120,N_12899,N_12680);
nor U13121 (N_13121,N_12611,N_12653);
or U13122 (N_13122,N_12717,N_12669);
or U13123 (N_13123,N_12691,N_12957);
nor U13124 (N_13124,N_12946,N_12608);
and U13125 (N_13125,N_12982,N_12924);
xor U13126 (N_13126,N_12787,N_12587);
xnor U13127 (N_13127,N_12793,N_12820);
or U13128 (N_13128,N_12708,N_12941);
xnor U13129 (N_13129,N_12834,N_12650);
nand U13130 (N_13130,N_12814,N_12752);
and U13131 (N_13131,N_12984,N_12892);
nor U13132 (N_13132,N_12978,N_12802);
and U13133 (N_13133,N_12578,N_12524);
xor U13134 (N_13134,N_12737,N_12719);
xnor U13135 (N_13135,N_12976,N_12624);
nand U13136 (N_13136,N_12569,N_12818);
or U13137 (N_13137,N_12864,N_12677);
nor U13138 (N_13138,N_12652,N_12565);
nand U13139 (N_13139,N_12909,N_12596);
xor U13140 (N_13140,N_12967,N_12862);
xor U13141 (N_13141,N_12694,N_12917);
nand U13142 (N_13142,N_12969,N_12854);
xnor U13143 (N_13143,N_12645,N_12686);
or U13144 (N_13144,N_12939,N_12698);
and U13145 (N_13145,N_12532,N_12819);
or U13146 (N_13146,N_12994,N_12935);
or U13147 (N_13147,N_12702,N_12791);
nand U13148 (N_13148,N_12806,N_12757);
xnor U13149 (N_13149,N_12848,N_12919);
or U13150 (N_13150,N_12780,N_12630);
nor U13151 (N_13151,N_12798,N_12570);
nor U13152 (N_13152,N_12755,N_12743);
xor U13153 (N_13153,N_12612,N_12959);
or U13154 (N_13154,N_12740,N_12514);
nor U13155 (N_13155,N_12966,N_12912);
xnor U13156 (N_13156,N_12718,N_12906);
and U13157 (N_13157,N_12991,N_12852);
xnor U13158 (N_13158,N_12931,N_12513);
nor U13159 (N_13159,N_12754,N_12508);
and U13160 (N_13160,N_12725,N_12844);
or U13161 (N_13161,N_12886,N_12535);
nor U13162 (N_13162,N_12561,N_12799);
xnor U13163 (N_13163,N_12965,N_12996);
nand U13164 (N_13164,N_12733,N_12597);
xnor U13165 (N_13165,N_12517,N_12549);
nor U13166 (N_13166,N_12647,N_12890);
or U13167 (N_13167,N_12989,N_12613);
nor U13168 (N_13168,N_12518,N_12929);
or U13169 (N_13169,N_12626,N_12665);
nor U13170 (N_13170,N_12895,N_12654);
or U13171 (N_13171,N_12902,N_12808);
and U13172 (N_13172,N_12860,N_12640);
xor U13173 (N_13173,N_12753,N_12842);
nand U13174 (N_13174,N_12789,N_12900);
xnor U13175 (N_13175,N_12979,N_12875);
and U13176 (N_13176,N_12901,N_12958);
xnor U13177 (N_13177,N_12771,N_12841);
xnor U13178 (N_13178,N_12734,N_12881);
nor U13179 (N_13179,N_12696,N_12516);
and U13180 (N_13180,N_12971,N_12655);
nor U13181 (N_13181,N_12605,N_12995);
nor U13182 (N_13182,N_12824,N_12526);
or U13183 (N_13183,N_12622,N_12894);
and U13184 (N_13184,N_12573,N_12580);
nor U13185 (N_13185,N_12690,N_12574);
nor U13186 (N_13186,N_12710,N_12555);
or U13187 (N_13187,N_12893,N_12947);
xnor U13188 (N_13188,N_12891,N_12805);
or U13189 (N_13189,N_12551,N_12525);
or U13190 (N_13190,N_12649,N_12689);
or U13191 (N_13191,N_12975,N_12986);
nand U13192 (N_13192,N_12963,N_12633);
or U13193 (N_13193,N_12693,N_12581);
nor U13194 (N_13194,N_12922,N_12785);
and U13195 (N_13195,N_12648,N_12638);
xor U13196 (N_13196,N_12503,N_12889);
and U13197 (N_13197,N_12988,N_12604);
nor U13198 (N_13198,N_12730,N_12759);
and U13199 (N_13199,N_12510,N_12985);
nand U13200 (N_13200,N_12878,N_12713);
xor U13201 (N_13201,N_12911,N_12623);
and U13202 (N_13202,N_12758,N_12885);
or U13203 (N_13203,N_12584,N_12566);
xnor U13204 (N_13204,N_12783,N_12884);
or U13205 (N_13205,N_12547,N_12827);
nand U13206 (N_13206,N_12756,N_12603);
nand U13207 (N_13207,N_12620,N_12825);
or U13208 (N_13208,N_12550,N_12951);
nand U13209 (N_13209,N_12803,N_12955);
and U13210 (N_13210,N_12610,N_12934);
xnor U13211 (N_13211,N_12961,N_12554);
xnor U13212 (N_13212,N_12936,N_12729);
xor U13213 (N_13213,N_12964,N_12839);
and U13214 (N_13214,N_12810,N_12760);
or U13215 (N_13215,N_12594,N_12720);
nor U13216 (N_13216,N_12564,N_12674);
nand U13217 (N_13217,N_12545,N_12522);
nor U13218 (N_13218,N_12857,N_12684);
nand U13219 (N_13219,N_12749,N_12709);
xor U13220 (N_13220,N_12776,N_12681);
and U13221 (N_13221,N_12981,N_12707);
and U13222 (N_13222,N_12634,N_12764);
nor U13223 (N_13223,N_12747,N_12521);
nand U13224 (N_13224,N_12533,N_12543);
and U13225 (N_13225,N_12865,N_12831);
and U13226 (N_13226,N_12795,N_12542);
and U13227 (N_13227,N_12590,N_12832);
or U13228 (N_13228,N_12662,N_12823);
xnor U13229 (N_13229,N_12859,N_12850);
nand U13230 (N_13230,N_12511,N_12858);
nand U13231 (N_13231,N_12905,N_12927);
nor U13232 (N_13232,N_12938,N_12618);
xor U13233 (N_13233,N_12849,N_12528);
and U13234 (N_13234,N_12643,N_12703);
nor U13235 (N_13235,N_12727,N_12866);
or U13236 (N_13236,N_12557,N_12616);
or U13237 (N_13237,N_12619,N_12898);
nor U13238 (N_13238,N_12855,N_12792);
nand U13239 (N_13239,N_12786,N_12871);
and U13240 (N_13240,N_12918,N_12904);
and U13241 (N_13241,N_12763,N_12579);
and U13242 (N_13242,N_12530,N_12592);
and U13243 (N_13243,N_12586,N_12615);
nor U13244 (N_13244,N_12632,N_12534);
nand U13245 (N_13245,N_12515,N_12697);
or U13246 (N_13246,N_12804,N_12504);
xor U13247 (N_13247,N_12954,N_12637);
nor U13248 (N_13248,N_12829,N_12732);
and U13249 (N_13249,N_12944,N_12914);
or U13250 (N_13250,N_12630,N_12516);
nor U13251 (N_13251,N_12981,N_12608);
nand U13252 (N_13252,N_12747,N_12580);
or U13253 (N_13253,N_12526,N_12537);
xnor U13254 (N_13254,N_12717,N_12541);
nand U13255 (N_13255,N_12819,N_12802);
nor U13256 (N_13256,N_12712,N_12918);
or U13257 (N_13257,N_12568,N_12747);
nor U13258 (N_13258,N_12599,N_12965);
nor U13259 (N_13259,N_12880,N_12795);
nand U13260 (N_13260,N_12735,N_12742);
nor U13261 (N_13261,N_12758,N_12764);
nand U13262 (N_13262,N_12749,N_12623);
or U13263 (N_13263,N_12945,N_12637);
nor U13264 (N_13264,N_12826,N_12505);
nand U13265 (N_13265,N_12669,N_12877);
xnor U13266 (N_13266,N_12974,N_12928);
and U13267 (N_13267,N_12555,N_12643);
and U13268 (N_13268,N_12572,N_12999);
or U13269 (N_13269,N_12568,N_12977);
and U13270 (N_13270,N_12830,N_12826);
xor U13271 (N_13271,N_12780,N_12799);
nand U13272 (N_13272,N_12539,N_12830);
and U13273 (N_13273,N_12536,N_12833);
nand U13274 (N_13274,N_12664,N_12915);
nand U13275 (N_13275,N_12857,N_12760);
and U13276 (N_13276,N_12979,N_12687);
nand U13277 (N_13277,N_12703,N_12888);
nor U13278 (N_13278,N_12755,N_12837);
and U13279 (N_13279,N_12632,N_12744);
xnor U13280 (N_13280,N_12816,N_12869);
nor U13281 (N_13281,N_12518,N_12573);
nand U13282 (N_13282,N_12675,N_12760);
nand U13283 (N_13283,N_12838,N_12585);
nor U13284 (N_13284,N_12710,N_12509);
nor U13285 (N_13285,N_12767,N_12717);
xor U13286 (N_13286,N_12803,N_12736);
nand U13287 (N_13287,N_12585,N_12981);
and U13288 (N_13288,N_12888,N_12555);
or U13289 (N_13289,N_12712,N_12936);
or U13290 (N_13290,N_12548,N_12672);
nor U13291 (N_13291,N_12500,N_12760);
nor U13292 (N_13292,N_12742,N_12979);
xor U13293 (N_13293,N_12795,N_12755);
xnor U13294 (N_13294,N_12775,N_12814);
nor U13295 (N_13295,N_12757,N_12663);
xnor U13296 (N_13296,N_12645,N_12542);
nand U13297 (N_13297,N_12759,N_12800);
nand U13298 (N_13298,N_12887,N_12923);
or U13299 (N_13299,N_12714,N_12998);
nor U13300 (N_13300,N_12997,N_12764);
or U13301 (N_13301,N_12721,N_12660);
nand U13302 (N_13302,N_12749,N_12565);
nor U13303 (N_13303,N_12933,N_12539);
nor U13304 (N_13304,N_12902,N_12787);
and U13305 (N_13305,N_12695,N_12776);
or U13306 (N_13306,N_12989,N_12905);
nand U13307 (N_13307,N_12591,N_12846);
nor U13308 (N_13308,N_12603,N_12788);
or U13309 (N_13309,N_12988,N_12827);
xnor U13310 (N_13310,N_12842,N_12919);
xnor U13311 (N_13311,N_12987,N_12716);
nand U13312 (N_13312,N_12787,N_12783);
nor U13313 (N_13313,N_12566,N_12669);
or U13314 (N_13314,N_12749,N_12515);
xnor U13315 (N_13315,N_12542,N_12643);
and U13316 (N_13316,N_12960,N_12657);
or U13317 (N_13317,N_12941,N_12848);
nor U13318 (N_13318,N_12749,N_12555);
or U13319 (N_13319,N_12869,N_12703);
or U13320 (N_13320,N_12691,N_12774);
xor U13321 (N_13321,N_12507,N_12937);
nand U13322 (N_13322,N_12566,N_12796);
nand U13323 (N_13323,N_12853,N_12669);
xnor U13324 (N_13324,N_12996,N_12841);
nor U13325 (N_13325,N_12824,N_12558);
nand U13326 (N_13326,N_12554,N_12894);
nand U13327 (N_13327,N_12511,N_12811);
nor U13328 (N_13328,N_12945,N_12639);
nand U13329 (N_13329,N_12969,N_12561);
nand U13330 (N_13330,N_12601,N_12910);
or U13331 (N_13331,N_12887,N_12730);
nor U13332 (N_13332,N_12986,N_12873);
xnor U13333 (N_13333,N_12613,N_12637);
nor U13334 (N_13334,N_12503,N_12902);
nand U13335 (N_13335,N_12985,N_12723);
nand U13336 (N_13336,N_12947,N_12635);
and U13337 (N_13337,N_12777,N_12698);
xor U13338 (N_13338,N_12598,N_12957);
and U13339 (N_13339,N_12679,N_12793);
and U13340 (N_13340,N_12750,N_12538);
xor U13341 (N_13341,N_12768,N_12951);
and U13342 (N_13342,N_12581,N_12950);
nand U13343 (N_13343,N_12505,N_12984);
nor U13344 (N_13344,N_12765,N_12750);
nor U13345 (N_13345,N_12741,N_12806);
or U13346 (N_13346,N_12644,N_12604);
and U13347 (N_13347,N_12670,N_12916);
and U13348 (N_13348,N_12937,N_12838);
or U13349 (N_13349,N_12763,N_12557);
or U13350 (N_13350,N_12679,N_12563);
and U13351 (N_13351,N_12954,N_12663);
and U13352 (N_13352,N_12848,N_12999);
nor U13353 (N_13353,N_12842,N_12856);
or U13354 (N_13354,N_12863,N_12980);
or U13355 (N_13355,N_12553,N_12851);
and U13356 (N_13356,N_12971,N_12524);
nor U13357 (N_13357,N_12651,N_12531);
nand U13358 (N_13358,N_12654,N_12975);
nor U13359 (N_13359,N_12734,N_12682);
or U13360 (N_13360,N_12853,N_12572);
nor U13361 (N_13361,N_12715,N_12821);
xnor U13362 (N_13362,N_12554,N_12690);
xor U13363 (N_13363,N_12745,N_12668);
nand U13364 (N_13364,N_12837,N_12879);
nand U13365 (N_13365,N_12509,N_12753);
nor U13366 (N_13366,N_12736,N_12536);
xor U13367 (N_13367,N_12671,N_12894);
xor U13368 (N_13368,N_12523,N_12659);
xnor U13369 (N_13369,N_12646,N_12530);
and U13370 (N_13370,N_12625,N_12859);
nand U13371 (N_13371,N_12726,N_12885);
nor U13372 (N_13372,N_12637,N_12755);
nand U13373 (N_13373,N_12980,N_12932);
or U13374 (N_13374,N_12611,N_12754);
nand U13375 (N_13375,N_12609,N_12784);
nand U13376 (N_13376,N_12668,N_12897);
nor U13377 (N_13377,N_12893,N_12748);
nor U13378 (N_13378,N_12614,N_12933);
nand U13379 (N_13379,N_12725,N_12838);
or U13380 (N_13380,N_12531,N_12772);
and U13381 (N_13381,N_12721,N_12538);
nor U13382 (N_13382,N_12956,N_12877);
or U13383 (N_13383,N_12933,N_12719);
nor U13384 (N_13384,N_12805,N_12542);
xor U13385 (N_13385,N_12724,N_12903);
or U13386 (N_13386,N_12514,N_12610);
or U13387 (N_13387,N_12908,N_12824);
xnor U13388 (N_13388,N_12947,N_12529);
nand U13389 (N_13389,N_12941,N_12545);
or U13390 (N_13390,N_12887,N_12761);
nand U13391 (N_13391,N_12745,N_12716);
or U13392 (N_13392,N_12717,N_12718);
nand U13393 (N_13393,N_12828,N_12780);
and U13394 (N_13394,N_12768,N_12802);
nand U13395 (N_13395,N_12538,N_12665);
xor U13396 (N_13396,N_12927,N_12951);
or U13397 (N_13397,N_12867,N_12554);
xor U13398 (N_13398,N_12865,N_12875);
and U13399 (N_13399,N_12701,N_12681);
nor U13400 (N_13400,N_12806,N_12994);
xnor U13401 (N_13401,N_12690,N_12928);
and U13402 (N_13402,N_12877,N_12986);
xnor U13403 (N_13403,N_12653,N_12619);
nand U13404 (N_13404,N_12527,N_12660);
xnor U13405 (N_13405,N_12939,N_12744);
xnor U13406 (N_13406,N_12943,N_12944);
xor U13407 (N_13407,N_12786,N_12591);
and U13408 (N_13408,N_12598,N_12568);
or U13409 (N_13409,N_12575,N_12665);
nor U13410 (N_13410,N_12779,N_12930);
or U13411 (N_13411,N_12620,N_12580);
xor U13412 (N_13412,N_12695,N_12620);
nand U13413 (N_13413,N_12561,N_12876);
nand U13414 (N_13414,N_12778,N_12657);
xnor U13415 (N_13415,N_12930,N_12802);
nor U13416 (N_13416,N_12967,N_12816);
or U13417 (N_13417,N_12753,N_12687);
nand U13418 (N_13418,N_12625,N_12777);
and U13419 (N_13419,N_12536,N_12850);
nand U13420 (N_13420,N_12778,N_12814);
nand U13421 (N_13421,N_12507,N_12631);
and U13422 (N_13422,N_12996,N_12508);
nand U13423 (N_13423,N_12801,N_12512);
nand U13424 (N_13424,N_12597,N_12963);
nand U13425 (N_13425,N_12962,N_12707);
nor U13426 (N_13426,N_12652,N_12558);
or U13427 (N_13427,N_12535,N_12658);
and U13428 (N_13428,N_12737,N_12988);
or U13429 (N_13429,N_12960,N_12654);
nor U13430 (N_13430,N_12849,N_12988);
nor U13431 (N_13431,N_12558,N_12948);
nor U13432 (N_13432,N_12748,N_12885);
nand U13433 (N_13433,N_12968,N_12836);
or U13434 (N_13434,N_12508,N_12726);
xnor U13435 (N_13435,N_12884,N_12532);
nand U13436 (N_13436,N_12825,N_12686);
nor U13437 (N_13437,N_12793,N_12663);
and U13438 (N_13438,N_12517,N_12777);
nand U13439 (N_13439,N_12987,N_12811);
nand U13440 (N_13440,N_12818,N_12504);
nand U13441 (N_13441,N_12646,N_12989);
xnor U13442 (N_13442,N_12670,N_12778);
xnor U13443 (N_13443,N_12819,N_12797);
nand U13444 (N_13444,N_12885,N_12859);
xor U13445 (N_13445,N_12590,N_12575);
xor U13446 (N_13446,N_12682,N_12980);
nor U13447 (N_13447,N_12758,N_12975);
and U13448 (N_13448,N_12815,N_12736);
nand U13449 (N_13449,N_12986,N_12965);
and U13450 (N_13450,N_12913,N_12744);
or U13451 (N_13451,N_12621,N_12916);
nand U13452 (N_13452,N_12533,N_12981);
and U13453 (N_13453,N_12548,N_12570);
and U13454 (N_13454,N_12792,N_12996);
nand U13455 (N_13455,N_12964,N_12891);
or U13456 (N_13456,N_12896,N_12541);
xnor U13457 (N_13457,N_12899,N_12853);
xor U13458 (N_13458,N_12952,N_12901);
xnor U13459 (N_13459,N_12517,N_12866);
and U13460 (N_13460,N_12807,N_12518);
xnor U13461 (N_13461,N_12586,N_12678);
xnor U13462 (N_13462,N_12835,N_12613);
and U13463 (N_13463,N_12791,N_12795);
xnor U13464 (N_13464,N_12820,N_12632);
or U13465 (N_13465,N_12751,N_12970);
nor U13466 (N_13466,N_12693,N_12803);
nor U13467 (N_13467,N_12797,N_12874);
and U13468 (N_13468,N_12721,N_12510);
nand U13469 (N_13469,N_12623,N_12819);
nor U13470 (N_13470,N_12679,N_12996);
and U13471 (N_13471,N_12568,N_12832);
nor U13472 (N_13472,N_12941,N_12923);
and U13473 (N_13473,N_12756,N_12682);
and U13474 (N_13474,N_12517,N_12703);
nor U13475 (N_13475,N_12760,N_12742);
and U13476 (N_13476,N_12678,N_12573);
nor U13477 (N_13477,N_12625,N_12603);
and U13478 (N_13478,N_12654,N_12540);
or U13479 (N_13479,N_12503,N_12642);
nor U13480 (N_13480,N_12764,N_12984);
nand U13481 (N_13481,N_12554,N_12825);
nor U13482 (N_13482,N_12928,N_12577);
and U13483 (N_13483,N_12902,N_12708);
nor U13484 (N_13484,N_12584,N_12823);
xor U13485 (N_13485,N_12912,N_12929);
and U13486 (N_13486,N_12799,N_12503);
nand U13487 (N_13487,N_12703,N_12788);
or U13488 (N_13488,N_12752,N_12858);
nand U13489 (N_13489,N_12854,N_12741);
or U13490 (N_13490,N_12552,N_12794);
and U13491 (N_13491,N_12836,N_12509);
or U13492 (N_13492,N_12916,N_12586);
xnor U13493 (N_13493,N_12620,N_12880);
and U13494 (N_13494,N_12939,N_12981);
nand U13495 (N_13495,N_12827,N_12956);
and U13496 (N_13496,N_12844,N_12515);
nand U13497 (N_13497,N_12517,N_12988);
nor U13498 (N_13498,N_12953,N_12913);
xnor U13499 (N_13499,N_12841,N_12797);
and U13500 (N_13500,N_13469,N_13154);
or U13501 (N_13501,N_13377,N_13046);
and U13502 (N_13502,N_13270,N_13347);
xnor U13503 (N_13503,N_13379,N_13261);
or U13504 (N_13504,N_13262,N_13300);
nand U13505 (N_13505,N_13039,N_13441);
nand U13506 (N_13506,N_13415,N_13194);
nand U13507 (N_13507,N_13081,N_13443);
nand U13508 (N_13508,N_13278,N_13173);
or U13509 (N_13509,N_13165,N_13127);
nand U13510 (N_13510,N_13301,N_13299);
nand U13511 (N_13511,N_13069,N_13392);
nor U13512 (N_13512,N_13130,N_13372);
nand U13513 (N_13513,N_13017,N_13411);
and U13514 (N_13514,N_13287,N_13420);
and U13515 (N_13515,N_13326,N_13015);
xor U13516 (N_13516,N_13158,N_13308);
nor U13517 (N_13517,N_13471,N_13280);
xnor U13518 (N_13518,N_13244,N_13119);
nand U13519 (N_13519,N_13283,N_13362);
and U13520 (N_13520,N_13075,N_13160);
nor U13521 (N_13521,N_13272,N_13322);
xnor U13522 (N_13522,N_13329,N_13034);
nor U13523 (N_13523,N_13185,N_13448);
xor U13524 (N_13524,N_13198,N_13213);
or U13525 (N_13525,N_13000,N_13037);
and U13526 (N_13526,N_13401,N_13204);
or U13527 (N_13527,N_13098,N_13397);
nor U13528 (N_13528,N_13170,N_13120);
xnor U13529 (N_13529,N_13445,N_13211);
nor U13530 (N_13530,N_13217,N_13096);
or U13531 (N_13531,N_13063,N_13020);
and U13532 (N_13532,N_13489,N_13054);
or U13533 (N_13533,N_13361,N_13205);
or U13534 (N_13534,N_13241,N_13385);
nand U13535 (N_13535,N_13146,N_13395);
xnor U13536 (N_13536,N_13365,N_13375);
and U13537 (N_13537,N_13378,N_13302);
nor U13538 (N_13538,N_13121,N_13239);
nand U13539 (N_13539,N_13223,N_13394);
nor U13540 (N_13540,N_13051,N_13011);
nand U13541 (N_13541,N_13203,N_13042);
or U13542 (N_13542,N_13148,N_13417);
or U13543 (N_13543,N_13414,N_13188);
nand U13544 (N_13544,N_13257,N_13114);
nor U13545 (N_13545,N_13087,N_13164);
xor U13546 (N_13546,N_13221,N_13058);
and U13547 (N_13547,N_13277,N_13467);
xnor U13548 (N_13548,N_13491,N_13080);
nand U13549 (N_13549,N_13136,N_13009);
nand U13550 (N_13550,N_13040,N_13274);
and U13551 (N_13551,N_13167,N_13123);
and U13552 (N_13552,N_13210,N_13376);
nand U13553 (N_13553,N_13332,N_13142);
nor U13554 (N_13554,N_13413,N_13144);
or U13555 (N_13555,N_13052,N_13012);
or U13556 (N_13556,N_13355,N_13271);
nand U13557 (N_13557,N_13357,N_13468);
or U13558 (N_13558,N_13187,N_13321);
nand U13559 (N_13559,N_13110,N_13026);
nand U13560 (N_13560,N_13062,N_13024);
or U13561 (N_13561,N_13073,N_13228);
or U13562 (N_13562,N_13151,N_13340);
nand U13563 (N_13563,N_13032,N_13422);
nor U13564 (N_13564,N_13006,N_13168);
xor U13565 (N_13565,N_13045,N_13427);
and U13566 (N_13566,N_13499,N_13192);
or U13567 (N_13567,N_13202,N_13072);
xnor U13568 (N_13568,N_13309,N_13150);
or U13569 (N_13569,N_13330,N_13156);
nor U13570 (N_13570,N_13313,N_13227);
or U13571 (N_13571,N_13050,N_13434);
nand U13572 (N_13572,N_13225,N_13311);
and U13573 (N_13573,N_13430,N_13090);
nor U13574 (N_13574,N_13129,N_13193);
or U13575 (N_13575,N_13003,N_13494);
nor U13576 (N_13576,N_13249,N_13460);
and U13577 (N_13577,N_13248,N_13028);
or U13578 (N_13578,N_13266,N_13320);
or U13579 (N_13579,N_13498,N_13306);
nand U13580 (N_13580,N_13482,N_13097);
or U13581 (N_13581,N_13426,N_13078);
nor U13582 (N_13582,N_13483,N_13140);
or U13583 (N_13583,N_13317,N_13153);
and U13584 (N_13584,N_13104,N_13013);
or U13585 (N_13585,N_13327,N_13292);
and U13586 (N_13586,N_13182,N_13041);
xor U13587 (N_13587,N_13149,N_13477);
or U13588 (N_13588,N_13388,N_13288);
or U13589 (N_13589,N_13297,N_13386);
or U13590 (N_13590,N_13094,N_13316);
xor U13591 (N_13591,N_13370,N_13111);
xnor U13592 (N_13592,N_13126,N_13195);
and U13593 (N_13593,N_13246,N_13304);
or U13594 (N_13594,N_13022,N_13323);
nor U13595 (N_13595,N_13486,N_13102);
xnor U13596 (N_13596,N_13218,N_13450);
nand U13597 (N_13597,N_13183,N_13189);
xnor U13598 (N_13598,N_13291,N_13492);
nor U13599 (N_13599,N_13474,N_13137);
nand U13600 (N_13600,N_13059,N_13172);
xor U13601 (N_13601,N_13439,N_13359);
nor U13602 (N_13602,N_13157,N_13001);
nand U13603 (N_13603,N_13402,N_13064);
or U13604 (N_13604,N_13125,N_13033);
or U13605 (N_13605,N_13263,N_13023);
nor U13606 (N_13606,N_13393,N_13464);
or U13607 (N_13607,N_13475,N_13255);
and U13608 (N_13608,N_13267,N_13077);
nand U13609 (N_13609,N_13235,N_13101);
nand U13610 (N_13610,N_13074,N_13162);
xnor U13611 (N_13611,N_13207,N_13497);
nand U13612 (N_13612,N_13452,N_13258);
nand U13613 (N_13613,N_13435,N_13438);
xnor U13614 (N_13614,N_13368,N_13407);
nor U13615 (N_13615,N_13197,N_13147);
xnor U13616 (N_13616,N_13008,N_13175);
nand U13617 (N_13617,N_13229,N_13232);
or U13618 (N_13618,N_13337,N_13016);
nand U13619 (N_13619,N_13408,N_13374);
and U13620 (N_13620,N_13495,N_13134);
or U13621 (N_13621,N_13243,N_13065);
nor U13622 (N_13622,N_13208,N_13479);
nand U13623 (N_13623,N_13002,N_13079);
and U13624 (N_13624,N_13476,N_13382);
or U13625 (N_13625,N_13222,N_13206);
and U13626 (N_13626,N_13176,N_13447);
or U13627 (N_13627,N_13336,N_13462);
xnor U13628 (N_13628,N_13354,N_13472);
or U13629 (N_13629,N_13036,N_13250);
or U13630 (N_13630,N_13117,N_13141);
nor U13631 (N_13631,N_13163,N_13356);
or U13632 (N_13632,N_13294,N_13133);
xnor U13633 (N_13633,N_13366,N_13350);
nor U13634 (N_13634,N_13084,N_13252);
nor U13635 (N_13635,N_13029,N_13296);
or U13636 (N_13636,N_13328,N_13406);
nor U13637 (N_13637,N_13285,N_13343);
and U13638 (N_13638,N_13043,N_13436);
or U13639 (N_13639,N_13412,N_13092);
nor U13640 (N_13640,N_13314,N_13289);
nand U13641 (N_13641,N_13181,N_13038);
nor U13642 (N_13642,N_13410,N_13259);
xor U13643 (N_13643,N_13014,N_13201);
or U13644 (N_13644,N_13260,N_13174);
xnor U13645 (N_13645,N_13371,N_13461);
and U13646 (N_13646,N_13053,N_13115);
and U13647 (N_13647,N_13100,N_13488);
xnor U13648 (N_13648,N_13113,N_13135);
and U13649 (N_13649,N_13238,N_13103);
nand U13650 (N_13650,N_13214,N_13122);
xnor U13651 (N_13651,N_13109,N_13403);
or U13652 (N_13652,N_13021,N_13303);
xor U13653 (N_13653,N_13066,N_13358);
xor U13654 (N_13654,N_13390,N_13421);
or U13655 (N_13655,N_13247,N_13236);
xnor U13656 (N_13656,N_13132,N_13216);
xnor U13657 (N_13657,N_13295,N_13493);
or U13658 (N_13658,N_13047,N_13480);
or U13659 (N_13659,N_13226,N_13035);
nand U13660 (N_13660,N_13025,N_13196);
and U13661 (N_13661,N_13444,N_13440);
nor U13662 (N_13662,N_13335,N_13433);
or U13663 (N_13663,N_13049,N_13107);
or U13664 (N_13664,N_13305,N_13245);
nand U13665 (N_13665,N_13166,N_13349);
and U13666 (N_13666,N_13384,N_13105);
or U13667 (N_13667,N_13383,N_13070);
nor U13668 (N_13668,N_13325,N_13082);
or U13669 (N_13669,N_13404,N_13083);
nand U13670 (N_13670,N_13018,N_13419);
xnor U13671 (N_13671,N_13190,N_13224);
or U13672 (N_13672,N_13298,N_13030);
nand U13673 (N_13673,N_13389,N_13031);
xor U13674 (N_13674,N_13286,N_13199);
and U13675 (N_13675,N_13484,N_13055);
and U13676 (N_13676,N_13345,N_13209);
or U13677 (N_13677,N_13152,N_13449);
or U13678 (N_13678,N_13446,N_13145);
xor U13679 (N_13679,N_13416,N_13071);
xnor U13680 (N_13680,N_13380,N_13454);
nor U13681 (N_13681,N_13004,N_13180);
or U13682 (N_13682,N_13159,N_13124);
xnor U13683 (N_13683,N_13233,N_13429);
or U13684 (N_13684,N_13085,N_13060);
or U13685 (N_13685,N_13352,N_13234);
nand U13686 (N_13686,N_13307,N_13086);
or U13687 (N_13687,N_13056,N_13019);
nand U13688 (N_13688,N_13089,N_13418);
nor U13689 (N_13689,N_13179,N_13273);
nor U13690 (N_13690,N_13437,N_13400);
or U13691 (N_13691,N_13398,N_13219);
or U13692 (N_13692,N_13342,N_13333);
or U13693 (N_13693,N_13138,N_13459);
and U13694 (N_13694,N_13409,N_13353);
nor U13695 (N_13695,N_13470,N_13131);
or U13696 (N_13696,N_13455,N_13282);
nand U13697 (N_13697,N_13473,N_13256);
and U13698 (N_13698,N_13184,N_13360);
or U13699 (N_13699,N_13399,N_13155);
and U13700 (N_13700,N_13265,N_13453);
and U13701 (N_13701,N_13027,N_13010);
nand U13702 (N_13702,N_13344,N_13112);
or U13703 (N_13703,N_13485,N_13348);
or U13704 (N_13704,N_13161,N_13191);
xnor U13705 (N_13705,N_13318,N_13281);
nor U13706 (N_13706,N_13212,N_13143);
and U13707 (N_13707,N_13373,N_13088);
and U13708 (N_13708,N_13108,N_13310);
and U13709 (N_13709,N_13331,N_13240);
xor U13710 (N_13710,N_13431,N_13334);
nand U13711 (N_13711,N_13095,N_13005);
xor U13712 (N_13712,N_13478,N_13369);
xnor U13713 (N_13713,N_13458,N_13496);
nor U13714 (N_13714,N_13405,N_13118);
xnor U13715 (N_13715,N_13215,N_13425);
and U13716 (N_13716,N_13293,N_13091);
nand U13717 (N_13717,N_13057,N_13044);
and U13718 (N_13718,N_13319,N_13264);
or U13719 (N_13719,N_13456,N_13481);
and U13720 (N_13720,N_13284,N_13381);
or U13721 (N_13721,N_13346,N_13387);
or U13722 (N_13722,N_13169,N_13007);
nand U13723 (N_13723,N_13128,N_13254);
nand U13724 (N_13724,N_13457,N_13432);
nand U13725 (N_13725,N_13424,N_13116);
and U13726 (N_13726,N_13339,N_13178);
xnor U13727 (N_13727,N_13338,N_13099);
and U13728 (N_13728,N_13442,N_13093);
or U13729 (N_13729,N_13220,N_13171);
xor U13730 (N_13730,N_13487,N_13279);
and U13731 (N_13731,N_13061,N_13048);
nor U13732 (N_13732,N_13364,N_13341);
nor U13733 (N_13733,N_13231,N_13466);
nand U13734 (N_13734,N_13428,N_13275);
nand U13735 (N_13735,N_13423,N_13391);
nand U13736 (N_13736,N_13067,N_13139);
and U13737 (N_13737,N_13242,N_13315);
nand U13738 (N_13738,N_13076,N_13312);
nand U13739 (N_13739,N_13269,N_13200);
or U13740 (N_13740,N_13367,N_13351);
xnor U13741 (N_13741,N_13230,N_13363);
nand U13742 (N_13742,N_13463,N_13106);
xnor U13743 (N_13743,N_13276,N_13451);
nor U13744 (N_13744,N_13268,N_13490);
xor U13745 (N_13745,N_13253,N_13396);
xor U13746 (N_13746,N_13237,N_13290);
or U13747 (N_13747,N_13186,N_13177);
xor U13748 (N_13748,N_13324,N_13465);
or U13749 (N_13749,N_13251,N_13068);
or U13750 (N_13750,N_13456,N_13430);
xnor U13751 (N_13751,N_13449,N_13046);
and U13752 (N_13752,N_13363,N_13441);
nor U13753 (N_13753,N_13055,N_13246);
nor U13754 (N_13754,N_13162,N_13464);
and U13755 (N_13755,N_13251,N_13299);
or U13756 (N_13756,N_13461,N_13329);
nand U13757 (N_13757,N_13169,N_13277);
nor U13758 (N_13758,N_13444,N_13290);
nand U13759 (N_13759,N_13135,N_13262);
or U13760 (N_13760,N_13421,N_13408);
xor U13761 (N_13761,N_13157,N_13011);
xor U13762 (N_13762,N_13254,N_13073);
xnor U13763 (N_13763,N_13094,N_13013);
or U13764 (N_13764,N_13479,N_13392);
xor U13765 (N_13765,N_13424,N_13441);
and U13766 (N_13766,N_13158,N_13402);
or U13767 (N_13767,N_13066,N_13114);
nand U13768 (N_13768,N_13354,N_13022);
or U13769 (N_13769,N_13392,N_13061);
nor U13770 (N_13770,N_13408,N_13250);
or U13771 (N_13771,N_13119,N_13019);
nor U13772 (N_13772,N_13216,N_13297);
or U13773 (N_13773,N_13053,N_13253);
nor U13774 (N_13774,N_13296,N_13243);
and U13775 (N_13775,N_13010,N_13151);
and U13776 (N_13776,N_13058,N_13472);
nand U13777 (N_13777,N_13488,N_13239);
xor U13778 (N_13778,N_13183,N_13488);
nand U13779 (N_13779,N_13255,N_13043);
and U13780 (N_13780,N_13407,N_13431);
nor U13781 (N_13781,N_13196,N_13417);
or U13782 (N_13782,N_13400,N_13017);
nor U13783 (N_13783,N_13037,N_13052);
and U13784 (N_13784,N_13198,N_13439);
nor U13785 (N_13785,N_13356,N_13121);
nand U13786 (N_13786,N_13092,N_13049);
or U13787 (N_13787,N_13340,N_13403);
and U13788 (N_13788,N_13389,N_13493);
nand U13789 (N_13789,N_13429,N_13486);
or U13790 (N_13790,N_13301,N_13168);
nand U13791 (N_13791,N_13218,N_13464);
xnor U13792 (N_13792,N_13435,N_13462);
and U13793 (N_13793,N_13168,N_13442);
xor U13794 (N_13794,N_13157,N_13164);
or U13795 (N_13795,N_13006,N_13399);
or U13796 (N_13796,N_13249,N_13239);
nand U13797 (N_13797,N_13109,N_13370);
nand U13798 (N_13798,N_13021,N_13350);
or U13799 (N_13799,N_13311,N_13249);
nand U13800 (N_13800,N_13112,N_13473);
xor U13801 (N_13801,N_13480,N_13361);
xnor U13802 (N_13802,N_13422,N_13350);
nor U13803 (N_13803,N_13116,N_13451);
nor U13804 (N_13804,N_13268,N_13176);
or U13805 (N_13805,N_13222,N_13112);
nand U13806 (N_13806,N_13150,N_13230);
nand U13807 (N_13807,N_13400,N_13109);
nand U13808 (N_13808,N_13470,N_13402);
nand U13809 (N_13809,N_13028,N_13427);
nand U13810 (N_13810,N_13171,N_13325);
or U13811 (N_13811,N_13445,N_13168);
nor U13812 (N_13812,N_13236,N_13444);
and U13813 (N_13813,N_13201,N_13465);
nor U13814 (N_13814,N_13016,N_13475);
nor U13815 (N_13815,N_13416,N_13260);
or U13816 (N_13816,N_13435,N_13009);
xnor U13817 (N_13817,N_13175,N_13017);
or U13818 (N_13818,N_13408,N_13228);
xor U13819 (N_13819,N_13096,N_13357);
nor U13820 (N_13820,N_13219,N_13183);
nand U13821 (N_13821,N_13005,N_13373);
and U13822 (N_13822,N_13187,N_13003);
nor U13823 (N_13823,N_13383,N_13431);
nor U13824 (N_13824,N_13420,N_13371);
and U13825 (N_13825,N_13428,N_13348);
xor U13826 (N_13826,N_13419,N_13459);
nand U13827 (N_13827,N_13297,N_13015);
xor U13828 (N_13828,N_13372,N_13217);
or U13829 (N_13829,N_13211,N_13133);
and U13830 (N_13830,N_13311,N_13247);
nor U13831 (N_13831,N_13134,N_13082);
nand U13832 (N_13832,N_13472,N_13482);
or U13833 (N_13833,N_13155,N_13225);
nand U13834 (N_13834,N_13355,N_13225);
nor U13835 (N_13835,N_13123,N_13233);
nand U13836 (N_13836,N_13190,N_13369);
and U13837 (N_13837,N_13146,N_13149);
and U13838 (N_13838,N_13255,N_13445);
or U13839 (N_13839,N_13488,N_13075);
nand U13840 (N_13840,N_13461,N_13307);
xnor U13841 (N_13841,N_13031,N_13349);
nor U13842 (N_13842,N_13046,N_13206);
xnor U13843 (N_13843,N_13407,N_13104);
or U13844 (N_13844,N_13326,N_13143);
and U13845 (N_13845,N_13348,N_13433);
or U13846 (N_13846,N_13184,N_13237);
and U13847 (N_13847,N_13476,N_13375);
nand U13848 (N_13848,N_13436,N_13420);
nor U13849 (N_13849,N_13263,N_13068);
nor U13850 (N_13850,N_13348,N_13080);
xnor U13851 (N_13851,N_13100,N_13069);
or U13852 (N_13852,N_13027,N_13273);
or U13853 (N_13853,N_13007,N_13285);
xnor U13854 (N_13854,N_13424,N_13466);
or U13855 (N_13855,N_13258,N_13370);
and U13856 (N_13856,N_13190,N_13020);
nand U13857 (N_13857,N_13343,N_13062);
nand U13858 (N_13858,N_13182,N_13270);
nand U13859 (N_13859,N_13119,N_13000);
xnor U13860 (N_13860,N_13012,N_13345);
nand U13861 (N_13861,N_13030,N_13410);
xnor U13862 (N_13862,N_13435,N_13432);
xor U13863 (N_13863,N_13205,N_13419);
or U13864 (N_13864,N_13089,N_13163);
and U13865 (N_13865,N_13165,N_13238);
nand U13866 (N_13866,N_13036,N_13478);
or U13867 (N_13867,N_13255,N_13112);
nor U13868 (N_13868,N_13044,N_13484);
xnor U13869 (N_13869,N_13433,N_13399);
nor U13870 (N_13870,N_13324,N_13105);
nand U13871 (N_13871,N_13480,N_13487);
or U13872 (N_13872,N_13187,N_13150);
nand U13873 (N_13873,N_13341,N_13308);
nand U13874 (N_13874,N_13432,N_13344);
nor U13875 (N_13875,N_13086,N_13432);
xor U13876 (N_13876,N_13003,N_13104);
or U13877 (N_13877,N_13278,N_13280);
or U13878 (N_13878,N_13058,N_13290);
nor U13879 (N_13879,N_13099,N_13023);
or U13880 (N_13880,N_13485,N_13465);
xor U13881 (N_13881,N_13000,N_13079);
nor U13882 (N_13882,N_13173,N_13027);
and U13883 (N_13883,N_13309,N_13273);
or U13884 (N_13884,N_13388,N_13073);
and U13885 (N_13885,N_13276,N_13438);
or U13886 (N_13886,N_13359,N_13390);
nand U13887 (N_13887,N_13136,N_13245);
nand U13888 (N_13888,N_13414,N_13497);
xor U13889 (N_13889,N_13260,N_13240);
nand U13890 (N_13890,N_13252,N_13428);
and U13891 (N_13891,N_13460,N_13430);
and U13892 (N_13892,N_13033,N_13344);
xnor U13893 (N_13893,N_13152,N_13213);
xor U13894 (N_13894,N_13434,N_13391);
and U13895 (N_13895,N_13393,N_13235);
and U13896 (N_13896,N_13377,N_13419);
nor U13897 (N_13897,N_13429,N_13226);
or U13898 (N_13898,N_13168,N_13026);
and U13899 (N_13899,N_13223,N_13262);
nor U13900 (N_13900,N_13449,N_13007);
xor U13901 (N_13901,N_13009,N_13002);
nor U13902 (N_13902,N_13177,N_13220);
nor U13903 (N_13903,N_13438,N_13215);
nor U13904 (N_13904,N_13061,N_13264);
or U13905 (N_13905,N_13273,N_13209);
nand U13906 (N_13906,N_13467,N_13102);
nor U13907 (N_13907,N_13201,N_13089);
nor U13908 (N_13908,N_13405,N_13467);
nor U13909 (N_13909,N_13439,N_13440);
nor U13910 (N_13910,N_13122,N_13455);
and U13911 (N_13911,N_13089,N_13289);
nand U13912 (N_13912,N_13039,N_13412);
or U13913 (N_13913,N_13088,N_13380);
or U13914 (N_13914,N_13467,N_13236);
and U13915 (N_13915,N_13239,N_13093);
xor U13916 (N_13916,N_13165,N_13093);
nand U13917 (N_13917,N_13020,N_13314);
or U13918 (N_13918,N_13493,N_13274);
nor U13919 (N_13919,N_13331,N_13204);
or U13920 (N_13920,N_13308,N_13402);
nor U13921 (N_13921,N_13074,N_13181);
xnor U13922 (N_13922,N_13163,N_13263);
xor U13923 (N_13923,N_13128,N_13235);
xor U13924 (N_13924,N_13136,N_13023);
xnor U13925 (N_13925,N_13462,N_13316);
and U13926 (N_13926,N_13344,N_13298);
and U13927 (N_13927,N_13140,N_13348);
nand U13928 (N_13928,N_13153,N_13354);
nand U13929 (N_13929,N_13226,N_13128);
nor U13930 (N_13930,N_13321,N_13129);
nand U13931 (N_13931,N_13041,N_13045);
xor U13932 (N_13932,N_13130,N_13172);
xnor U13933 (N_13933,N_13081,N_13120);
or U13934 (N_13934,N_13272,N_13467);
nor U13935 (N_13935,N_13017,N_13470);
xnor U13936 (N_13936,N_13358,N_13371);
or U13937 (N_13937,N_13264,N_13374);
or U13938 (N_13938,N_13413,N_13233);
xor U13939 (N_13939,N_13175,N_13312);
or U13940 (N_13940,N_13429,N_13485);
xor U13941 (N_13941,N_13227,N_13277);
nor U13942 (N_13942,N_13013,N_13311);
nand U13943 (N_13943,N_13161,N_13277);
or U13944 (N_13944,N_13160,N_13142);
xnor U13945 (N_13945,N_13157,N_13124);
xnor U13946 (N_13946,N_13220,N_13019);
and U13947 (N_13947,N_13301,N_13497);
nor U13948 (N_13948,N_13219,N_13121);
xnor U13949 (N_13949,N_13360,N_13399);
xor U13950 (N_13950,N_13310,N_13490);
xor U13951 (N_13951,N_13122,N_13452);
and U13952 (N_13952,N_13294,N_13223);
xnor U13953 (N_13953,N_13313,N_13068);
xor U13954 (N_13954,N_13225,N_13451);
nor U13955 (N_13955,N_13222,N_13444);
and U13956 (N_13956,N_13028,N_13205);
nor U13957 (N_13957,N_13211,N_13210);
xnor U13958 (N_13958,N_13175,N_13154);
xor U13959 (N_13959,N_13322,N_13176);
nand U13960 (N_13960,N_13106,N_13416);
or U13961 (N_13961,N_13246,N_13331);
nand U13962 (N_13962,N_13348,N_13440);
and U13963 (N_13963,N_13417,N_13094);
or U13964 (N_13964,N_13278,N_13260);
nand U13965 (N_13965,N_13473,N_13494);
and U13966 (N_13966,N_13460,N_13104);
xor U13967 (N_13967,N_13340,N_13376);
nand U13968 (N_13968,N_13443,N_13328);
and U13969 (N_13969,N_13045,N_13334);
and U13970 (N_13970,N_13466,N_13167);
nor U13971 (N_13971,N_13080,N_13363);
nor U13972 (N_13972,N_13122,N_13082);
or U13973 (N_13973,N_13024,N_13159);
nor U13974 (N_13974,N_13142,N_13141);
xor U13975 (N_13975,N_13212,N_13100);
and U13976 (N_13976,N_13408,N_13156);
xnor U13977 (N_13977,N_13464,N_13244);
nand U13978 (N_13978,N_13067,N_13443);
and U13979 (N_13979,N_13034,N_13023);
or U13980 (N_13980,N_13036,N_13430);
and U13981 (N_13981,N_13419,N_13431);
and U13982 (N_13982,N_13197,N_13472);
nor U13983 (N_13983,N_13030,N_13272);
xor U13984 (N_13984,N_13056,N_13199);
nand U13985 (N_13985,N_13385,N_13001);
or U13986 (N_13986,N_13404,N_13461);
nor U13987 (N_13987,N_13463,N_13018);
or U13988 (N_13988,N_13270,N_13058);
nor U13989 (N_13989,N_13223,N_13292);
and U13990 (N_13990,N_13349,N_13477);
or U13991 (N_13991,N_13394,N_13229);
xor U13992 (N_13992,N_13034,N_13160);
and U13993 (N_13993,N_13305,N_13384);
or U13994 (N_13994,N_13243,N_13121);
nor U13995 (N_13995,N_13385,N_13494);
nand U13996 (N_13996,N_13359,N_13459);
xor U13997 (N_13997,N_13282,N_13484);
nor U13998 (N_13998,N_13386,N_13104);
nor U13999 (N_13999,N_13038,N_13379);
and U14000 (N_14000,N_13852,N_13857);
or U14001 (N_14001,N_13821,N_13928);
nand U14002 (N_14002,N_13822,N_13794);
or U14003 (N_14003,N_13882,N_13741);
xnor U14004 (N_14004,N_13909,N_13649);
and U14005 (N_14005,N_13527,N_13792);
and U14006 (N_14006,N_13769,N_13534);
nor U14007 (N_14007,N_13674,N_13910);
nor U14008 (N_14008,N_13580,N_13807);
nand U14009 (N_14009,N_13962,N_13633);
xor U14010 (N_14010,N_13772,N_13914);
xor U14011 (N_14011,N_13791,N_13758);
or U14012 (N_14012,N_13903,N_13627);
nand U14013 (N_14013,N_13537,N_13713);
nand U14014 (N_14014,N_13767,N_13912);
nor U14015 (N_14015,N_13593,N_13734);
or U14016 (N_14016,N_13707,N_13724);
nand U14017 (N_14017,N_13886,N_13860);
xnor U14018 (N_14018,N_13943,N_13679);
or U14019 (N_14019,N_13582,N_13748);
xor U14020 (N_14020,N_13991,N_13884);
nor U14021 (N_14021,N_13826,N_13782);
and U14022 (N_14022,N_13690,N_13892);
or U14023 (N_14023,N_13677,N_13836);
nand U14024 (N_14024,N_13916,N_13917);
nand U14025 (N_14025,N_13825,N_13997);
or U14026 (N_14026,N_13517,N_13875);
xor U14027 (N_14027,N_13592,N_13558);
and U14028 (N_14028,N_13549,N_13541);
or U14029 (N_14029,N_13745,N_13648);
and U14030 (N_14030,N_13625,N_13617);
or U14031 (N_14031,N_13802,N_13557);
nor U14032 (N_14032,N_13766,N_13819);
nor U14033 (N_14033,N_13781,N_13979);
nand U14034 (N_14034,N_13835,N_13828);
xor U14035 (N_14035,N_13737,N_13650);
xor U14036 (N_14036,N_13984,N_13656);
or U14037 (N_14037,N_13880,N_13711);
nand U14038 (N_14038,N_13765,N_13507);
nand U14039 (N_14039,N_13803,N_13978);
nor U14040 (N_14040,N_13850,N_13531);
nand U14041 (N_14041,N_13876,N_13809);
or U14042 (N_14042,N_13501,N_13851);
and U14043 (N_14043,N_13591,N_13746);
and U14044 (N_14044,N_13614,N_13578);
nor U14045 (N_14045,N_13568,N_13814);
or U14046 (N_14046,N_13637,N_13998);
and U14047 (N_14047,N_13702,N_13575);
xnor U14048 (N_14048,N_13606,N_13581);
or U14049 (N_14049,N_13899,N_13529);
or U14050 (N_14050,N_13840,N_13936);
and U14051 (N_14051,N_13981,N_13958);
xor U14052 (N_14052,N_13584,N_13671);
nand U14053 (N_14053,N_13595,N_13925);
nand U14054 (N_14054,N_13990,N_13740);
or U14055 (N_14055,N_13780,N_13691);
and U14056 (N_14056,N_13793,N_13594);
xor U14057 (N_14057,N_13621,N_13921);
nor U14058 (N_14058,N_13629,N_13654);
nor U14059 (N_14059,N_13863,N_13866);
or U14060 (N_14060,N_13783,N_13618);
or U14061 (N_14061,N_13682,N_13735);
or U14062 (N_14062,N_13518,N_13833);
xor U14063 (N_14063,N_13996,N_13983);
nor U14064 (N_14064,N_13804,N_13881);
and U14065 (N_14065,N_13732,N_13940);
and U14066 (N_14066,N_13834,N_13567);
and U14067 (N_14067,N_13846,N_13779);
nor U14068 (N_14068,N_13898,N_13911);
xnor U14069 (N_14069,N_13811,N_13893);
nor U14070 (N_14070,N_13684,N_13873);
nor U14071 (N_14071,N_13610,N_13604);
nor U14072 (N_14072,N_13513,N_13564);
and U14073 (N_14073,N_13569,N_13700);
nand U14074 (N_14074,N_13915,N_13571);
xor U14075 (N_14075,N_13546,N_13738);
xor U14076 (N_14076,N_13858,N_13708);
and U14077 (N_14077,N_13718,N_13602);
or U14078 (N_14078,N_13750,N_13951);
nand U14079 (N_14079,N_13542,N_13528);
nor U14080 (N_14080,N_13658,N_13651);
or U14081 (N_14081,N_13784,N_13986);
and U14082 (N_14082,N_13511,N_13913);
xnor U14083 (N_14083,N_13747,N_13731);
and U14084 (N_14084,N_13956,N_13955);
xor U14085 (N_14085,N_13776,N_13773);
nand U14086 (N_14086,N_13670,N_13506);
and U14087 (N_14087,N_13799,N_13611);
nor U14088 (N_14088,N_13945,N_13757);
nand U14089 (N_14089,N_13641,N_13742);
nor U14090 (N_14090,N_13959,N_13775);
xnor U14091 (N_14091,N_13848,N_13743);
xor U14092 (N_14092,N_13504,N_13714);
xor U14093 (N_14093,N_13817,N_13721);
nand U14094 (N_14094,N_13644,N_13967);
and U14095 (N_14095,N_13662,N_13798);
xor U14096 (N_14096,N_13622,N_13993);
nand U14097 (N_14097,N_13631,N_13706);
xnor U14098 (N_14098,N_13638,N_13918);
xor U14099 (N_14099,N_13572,N_13992);
and U14100 (N_14100,N_13869,N_13597);
nand U14101 (N_14101,N_13647,N_13520);
xnor U14102 (N_14102,N_13503,N_13583);
xor U14103 (N_14103,N_13722,N_13980);
or U14104 (N_14104,N_13535,N_13946);
nor U14105 (N_14105,N_13608,N_13853);
nand U14106 (N_14106,N_13500,N_13639);
or U14107 (N_14107,N_13812,N_13620);
xnor U14108 (N_14108,N_13862,N_13890);
and U14109 (N_14109,N_13904,N_13539);
nor U14110 (N_14110,N_13847,N_13566);
and U14111 (N_14111,N_13538,N_13760);
xor U14112 (N_14112,N_13512,N_13665);
nor U14113 (N_14113,N_13554,N_13556);
nand U14114 (N_14114,N_13628,N_13762);
xor U14115 (N_14115,N_13710,N_13642);
xnor U14116 (N_14116,N_13994,N_13640);
and U14117 (N_14117,N_13953,N_13926);
nand U14118 (N_14118,N_13870,N_13563);
nor U14119 (N_14119,N_13896,N_13970);
nor U14120 (N_14120,N_13502,N_13759);
xnor U14121 (N_14121,N_13877,N_13788);
xnor U14122 (N_14122,N_13570,N_13543);
nand U14123 (N_14123,N_13676,N_13806);
xor U14124 (N_14124,N_13771,N_13823);
or U14125 (N_14125,N_13897,N_13523);
nor U14126 (N_14126,N_13599,N_13891);
and U14127 (N_14127,N_13709,N_13589);
or U14128 (N_14128,N_13626,N_13839);
nor U14129 (N_14129,N_13600,N_13895);
and U14130 (N_14130,N_13934,N_13712);
nand U14131 (N_14131,N_13590,N_13579);
nor U14132 (N_14132,N_13685,N_13944);
nor U14133 (N_14133,N_13937,N_13521);
nand U14134 (N_14134,N_13635,N_13723);
or U14135 (N_14135,N_13831,N_13971);
nand U14136 (N_14136,N_13824,N_13808);
nand U14137 (N_14137,N_13795,N_13796);
nand U14138 (N_14138,N_13588,N_13668);
and U14139 (N_14139,N_13923,N_13948);
and U14140 (N_14140,N_13837,N_13969);
nor U14141 (N_14141,N_13989,N_13612);
or U14142 (N_14142,N_13797,N_13536);
nor U14143 (N_14143,N_13548,N_13716);
nor U14144 (N_14144,N_13954,N_13615);
and U14145 (N_14145,N_13550,N_13975);
or U14146 (N_14146,N_13603,N_13753);
or U14147 (N_14147,N_13973,N_13829);
xor U14148 (N_14148,N_13867,N_13623);
and U14149 (N_14149,N_13810,N_13695);
nor U14150 (N_14150,N_13646,N_13778);
nand U14151 (N_14151,N_13949,N_13704);
nor U14152 (N_14152,N_13774,N_13841);
xor U14153 (N_14153,N_13634,N_13960);
xnor U14154 (N_14154,N_13878,N_13920);
xnor U14155 (N_14155,N_13785,N_13692);
or U14156 (N_14156,N_13843,N_13609);
nand U14157 (N_14157,N_13703,N_13976);
and U14158 (N_14158,N_13883,N_13607);
xor U14159 (N_14159,N_13889,N_13560);
nor U14160 (N_14160,N_13551,N_13968);
or U14161 (N_14161,N_13687,N_13942);
nand U14162 (N_14162,N_13729,N_13522);
xnor U14163 (N_14163,N_13761,N_13756);
nor U14164 (N_14164,N_13616,N_13935);
xor U14165 (N_14165,N_13813,N_13770);
nand U14166 (N_14166,N_13929,N_13552);
nand U14167 (N_14167,N_13533,N_13701);
or U14168 (N_14168,N_13559,N_13856);
nand U14169 (N_14169,N_13645,N_13950);
xnor U14170 (N_14170,N_13601,N_13947);
xor U14171 (N_14171,N_13966,N_13624);
and U14172 (N_14172,N_13699,N_13686);
xnor U14173 (N_14173,N_13669,N_13982);
and U14174 (N_14174,N_13664,N_13816);
nand U14175 (N_14175,N_13505,N_13939);
nor U14176 (N_14176,N_13906,N_13855);
or U14177 (N_14177,N_13977,N_13754);
xnor U14178 (N_14178,N_13832,N_13885);
and U14179 (N_14179,N_13919,N_13540);
and U14180 (N_14180,N_13547,N_13844);
or U14181 (N_14181,N_13988,N_13900);
xor U14182 (N_14182,N_13508,N_13787);
or U14183 (N_14183,N_13598,N_13660);
xnor U14184 (N_14184,N_13827,N_13657);
nand U14185 (N_14185,N_13815,N_13667);
or U14186 (N_14186,N_13931,N_13586);
nand U14187 (N_14187,N_13861,N_13525);
nand U14188 (N_14188,N_13805,N_13530);
or U14189 (N_14189,N_13965,N_13727);
xor U14190 (N_14190,N_13698,N_13532);
nor U14191 (N_14191,N_13924,N_13818);
nand U14192 (N_14192,N_13952,N_13874);
nor U14193 (N_14193,N_13561,N_13719);
xor U14194 (N_14194,N_13694,N_13613);
and U14195 (N_14195,N_13974,N_13894);
or U14196 (N_14196,N_13587,N_13605);
xor U14197 (N_14197,N_13764,N_13820);
and U14198 (N_14198,N_13736,N_13673);
nor U14199 (N_14199,N_13545,N_13653);
and U14200 (N_14200,N_13689,N_13562);
nor U14201 (N_14201,N_13553,N_13619);
xnor U14202 (N_14202,N_13985,N_13663);
xnor U14203 (N_14203,N_13672,N_13879);
nor U14204 (N_14204,N_13661,N_13596);
xnor U14205 (N_14205,N_13509,N_13927);
and U14206 (N_14206,N_13715,N_13696);
nor U14207 (N_14207,N_13720,N_13872);
and U14208 (N_14208,N_13871,N_13938);
nor U14209 (N_14209,N_13845,N_13865);
and U14210 (N_14210,N_13749,N_13730);
and U14211 (N_14211,N_13995,N_13972);
or U14212 (N_14212,N_13519,N_13887);
or U14213 (N_14213,N_13680,N_13728);
nor U14214 (N_14214,N_13632,N_13864);
and U14215 (N_14215,N_13739,N_13963);
xnor U14216 (N_14216,N_13726,N_13801);
nor U14217 (N_14217,N_13905,N_13655);
and U14218 (N_14218,N_13941,N_13636);
xor U14219 (N_14219,N_13901,N_13777);
or U14220 (N_14220,N_13678,N_13544);
xor U14221 (N_14221,N_13987,N_13842);
and U14222 (N_14222,N_13688,N_13515);
xor U14223 (N_14223,N_13859,N_13683);
nor U14224 (N_14224,N_13514,N_13681);
nand U14225 (N_14225,N_13725,N_13577);
and U14226 (N_14226,N_13675,N_13565);
nor U14227 (N_14227,N_13717,N_13922);
nor U14228 (N_14228,N_13907,N_13576);
nor U14229 (N_14229,N_13933,N_13800);
nand U14230 (N_14230,N_13744,N_13902);
and U14231 (N_14231,N_13930,N_13652);
and U14232 (N_14232,N_13733,N_13961);
nor U14233 (N_14233,N_13957,N_13830);
xor U14234 (N_14234,N_13516,N_13630);
nor U14235 (N_14235,N_13555,N_13752);
nand U14236 (N_14236,N_13755,N_13666);
or U14237 (N_14237,N_13697,N_13585);
or U14238 (N_14238,N_13789,N_13693);
xnor U14239 (N_14239,N_13868,N_13574);
and U14240 (N_14240,N_13888,N_13526);
and U14241 (N_14241,N_13838,N_13524);
nand U14242 (N_14242,N_13659,N_13999);
or U14243 (N_14243,N_13964,N_13786);
xnor U14244 (N_14244,N_13510,N_13705);
xor U14245 (N_14245,N_13854,N_13751);
and U14246 (N_14246,N_13763,N_13573);
and U14247 (N_14247,N_13849,N_13908);
nor U14248 (N_14248,N_13790,N_13643);
nand U14249 (N_14249,N_13768,N_13932);
or U14250 (N_14250,N_13857,N_13848);
nor U14251 (N_14251,N_13997,N_13876);
nand U14252 (N_14252,N_13723,N_13532);
or U14253 (N_14253,N_13521,N_13700);
xor U14254 (N_14254,N_13737,N_13661);
or U14255 (N_14255,N_13715,N_13778);
nor U14256 (N_14256,N_13775,N_13887);
nand U14257 (N_14257,N_13728,N_13665);
and U14258 (N_14258,N_13823,N_13810);
nor U14259 (N_14259,N_13525,N_13624);
and U14260 (N_14260,N_13777,N_13749);
and U14261 (N_14261,N_13598,N_13800);
nor U14262 (N_14262,N_13602,N_13955);
xnor U14263 (N_14263,N_13580,N_13749);
and U14264 (N_14264,N_13596,N_13532);
xnor U14265 (N_14265,N_13550,N_13920);
and U14266 (N_14266,N_13882,N_13683);
nand U14267 (N_14267,N_13552,N_13652);
nand U14268 (N_14268,N_13809,N_13774);
xnor U14269 (N_14269,N_13644,N_13694);
xor U14270 (N_14270,N_13622,N_13679);
xnor U14271 (N_14271,N_13678,N_13860);
nor U14272 (N_14272,N_13664,N_13899);
xor U14273 (N_14273,N_13769,N_13668);
nand U14274 (N_14274,N_13817,N_13590);
nand U14275 (N_14275,N_13746,N_13796);
and U14276 (N_14276,N_13626,N_13765);
or U14277 (N_14277,N_13986,N_13957);
xor U14278 (N_14278,N_13786,N_13843);
nor U14279 (N_14279,N_13643,N_13588);
or U14280 (N_14280,N_13868,N_13557);
and U14281 (N_14281,N_13725,N_13825);
nand U14282 (N_14282,N_13840,N_13501);
and U14283 (N_14283,N_13817,N_13560);
and U14284 (N_14284,N_13801,N_13903);
nor U14285 (N_14285,N_13720,N_13601);
xor U14286 (N_14286,N_13938,N_13759);
nor U14287 (N_14287,N_13828,N_13678);
nand U14288 (N_14288,N_13563,N_13799);
and U14289 (N_14289,N_13989,N_13824);
nand U14290 (N_14290,N_13852,N_13970);
nand U14291 (N_14291,N_13995,N_13646);
or U14292 (N_14292,N_13998,N_13716);
or U14293 (N_14293,N_13813,N_13779);
nand U14294 (N_14294,N_13835,N_13673);
nand U14295 (N_14295,N_13794,N_13587);
xor U14296 (N_14296,N_13511,N_13559);
nand U14297 (N_14297,N_13638,N_13850);
nor U14298 (N_14298,N_13804,N_13556);
nand U14299 (N_14299,N_13756,N_13679);
xnor U14300 (N_14300,N_13977,N_13813);
nor U14301 (N_14301,N_13861,N_13674);
nand U14302 (N_14302,N_13771,N_13840);
xnor U14303 (N_14303,N_13978,N_13699);
xor U14304 (N_14304,N_13771,N_13835);
nand U14305 (N_14305,N_13610,N_13935);
xor U14306 (N_14306,N_13850,N_13923);
xor U14307 (N_14307,N_13598,N_13521);
xnor U14308 (N_14308,N_13944,N_13686);
or U14309 (N_14309,N_13810,N_13619);
xnor U14310 (N_14310,N_13608,N_13914);
and U14311 (N_14311,N_13611,N_13723);
xor U14312 (N_14312,N_13711,N_13598);
or U14313 (N_14313,N_13842,N_13983);
and U14314 (N_14314,N_13851,N_13882);
and U14315 (N_14315,N_13762,N_13728);
or U14316 (N_14316,N_13834,N_13551);
and U14317 (N_14317,N_13860,N_13851);
nor U14318 (N_14318,N_13577,N_13557);
and U14319 (N_14319,N_13657,N_13940);
nor U14320 (N_14320,N_13910,N_13800);
or U14321 (N_14321,N_13530,N_13942);
nor U14322 (N_14322,N_13943,N_13993);
and U14323 (N_14323,N_13890,N_13762);
or U14324 (N_14324,N_13895,N_13682);
and U14325 (N_14325,N_13547,N_13592);
nor U14326 (N_14326,N_13674,N_13683);
or U14327 (N_14327,N_13657,N_13809);
nand U14328 (N_14328,N_13541,N_13785);
nor U14329 (N_14329,N_13602,N_13972);
nor U14330 (N_14330,N_13523,N_13975);
xor U14331 (N_14331,N_13511,N_13783);
or U14332 (N_14332,N_13921,N_13506);
nor U14333 (N_14333,N_13829,N_13917);
nor U14334 (N_14334,N_13726,N_13683);
nand U14335 (N_14335,N_13838,N_13931);
nor U14336 (N_14336,N_13829,N_13831);
nor U14337 (N_14337,N_13574,N_13786);
xor U14338 (N_14338,N_13576,N_13838);
nor U14339 (N_14339,N_13978,N_13749);
nand U14340 (N_14340,N_13923,N_13849);
or U14341 (N_14341,N_13908,N_13501);
and U14342 (N_14342,N_13841,N_13847);
nor U14343 (N_14343,N_13529,N_13567);
nand U14344 (N_14344,N_13512,N_13757);
nor U14345 (N_14345,N_13706,N_13780);
nand U14346 (N_14346,N_13582,N_13728);
nand U14347 (N_14347,N_13542,N_13533);
xor U14348 (N_14348,N_13756,N_13759);
and U14349 (N_14349,N_13818,N_13515);
nor U14350 (N_14350,N_13852,N_13767);
nor U14351 (N_14351,N_13923,N_13965);
nand U14352 (N_14352,N_13916,N_13886);
and U14353 (N_14353,N_13509,N_13528);
xor U14354 (N_14354,N_13728,N_13890);
or U14355 (N_14355,N_13655,N_13962);
and U14356 (N_14356,N_13659,N_13975);
or U14357 (N_14357,N_13779,N_13856);
nor U14358 (N_14358,N_13793,N_13790);
or U14359 (N_14359,N_13621,N_13613);
nand U14360 (N_14360,N_13778,N_13558);
and U14361 (N_14361,N_13930,N_13910);
nor U14362 (N_14362,N_13902,N_13689);
and U14363 (N_14363,N_13709,N_13816);
and U14364 (N_14364,N_13826,N_13566);
xor U14365 (N_14365,N_13768,N_13960);
or U14366 (N_14366,N_13755,N_13649);
nand U14367 (N_14367,N_13780,N_13897);
xor U14368 (N_14368,N_13705,N_13903);
or U14369 (N_14369,N_13595,N_13661);
nor U14370 (N_14370,N_13978,N_13622);
or U14371 (N_14371,N_13885,N_13867);
nor U14372 (N_14372,N_13670,N_13981);
and U14373 (N_14373,N_13574,N_13784);
and U14374 (N_14374,N_13701,N_13924);
xor U14375 (N_14375,N_13575,N_13964);
nor U14376 (N_14376,N_13619,N_13840);
or U14377 (N_14377,N_13616,N_13947);
and U14378 (N_14378,N_13631,N_13633);
nor U14379 (N_14379,N_13741,N_13525);
or U14380 (N_14380,N_13815,N_13537);
nor U14381 (N_14381,N_13703,N_13796);
or U14382 (N_14382,N_13805,N_13829);
nor U14383 (N_14383,N_13880,N_13949);
nor U14384 (N_14384,N_13756,N_13832);
or U14385 (N_14385,N_13886,N_13707);
nand U14386 (N_14386,N_13648,N_13787);
or U14387 (N_14387,N_13692,N_13676);
xnor U14388 (N_14388,N_13773,N_13813);
or U14389 (N_14389,N_13651,N_13953);
and U14390 (N_14390,N_13844,N_13542);
nand U14391 (N_14391,N_13810,N_13545);
or U14392 (N_14392,N_13601,N_13844);
nand U14393 (N_14393,N_13632,N_13878);
xnor U14394 (N_14394,N_13834,N_13736);
nand U14395 (N_14395,N_13639,N_13534);
and U14396 (N_14396,N_13944,N_13752);
nor U14397 (N_14397,N_13986,N_13910);
or U14398 (N_14398,N_13899,N_13773);
or U14399 (N_14399,N_13828,N_13543);
xor U14400 (N_14400,N_13681,N_13925);
or U14401 (N_14401,N_13539,N_13981);
nand U14402 (N_14402,N_13720,N_13873);
or U14403 (N_14403,N_13815,N_13694);
or U14404 (N_14404,N_13979,N_13597);
nor U14405 (N_14405,N_13621,N_13916);
or U14406 (N_14406,N_13696,N_13886);
nand U14407 (N_14407,N_13987,N_13592);
nand U14408 (N_14408,N_13649,N_13904);
xnor U14409 (N_14409,N_13834,N_13980);
or U14410 (N_14410,N_13966,N_13925);
or U14411 (N_14411,N_13570,N_13926);
nor U14412 (N_14412,N_13508,N_13851);
and U14413 (N_14413,N_13692,N_13674);
nor U14414 (N_14414,N_13771,N_13939);
nor U14415 (N_14415,N_13559,N_13892);
or U14416 (N_14416,N_13572,N_13615);
and U14417 (N_14417,N_13582,N_13782);
xor U14418 (N_14418,N_13738,N_13787);
nand U14419 (N_14419,N_13619,N_13998);
nor U14420 (N_14420,N_13929,N_13766);
xor U14421 (N_14421,N_13946,N_13883);
xor U14422 (N_14422,N_13961,N_13589);
or U14423 (N_14423,N_13725,N_13777);
nand U14424 (N_14424,N_13899,N_13802);
nand U14425 (N_14425,N_13822,N_13855);
and U14426 (N_14426,N_13717,N_13798);
nor U14427 (N_14427,N_13593,N_13653);
nand U14428 (N_14428,N_13903,N_13879);
or U14429 (N_14429,N_13510,N_13694);
nor U14430 (N_14430,N_13857,N_13733);
nand U14431 (N_14431,N_13652,N_13601);
and U14432 (N_14432,N_13557,N_13702);
or U14433 (N_14433,N_13794,N_13577);
xnor U14434 (N_14434,N_13805,N_13662);
nand U14435 (N_14435,N_13825,N_13685);
and U14436 (N_14436,N_13618,N_13539);
nor U14437 (N_14437,N_13925,N_13910);
or U14438 (N_14438,N_13814,N_13850);
or U14439 (N_14439,N_13559,N_13579);
and U14440 (N_14440,N_13844,N_13564);
and U14441 (N_14441,N_13898,N_13729);
nand U14442 (N_14442,N_13844,N_13586);
and U14443 (N_14443,N_13726,N_13687);
and U14444 (N_14444,N_13918,N_13957);
or U14445 (N_14445,N_13675,N_13516);
and U14446 (N_14446,N_13780,N_13645);
or U14447 (N_14447,N_13547,N_13687);
nor U14448 (N_14448,N_13559,N_13846);
nor U14449 (N_14449,N_13928,N_13635);
or U14450 (N_14450,N_13813,N_13888);
nor U14451 (N_14451,N_13715,N_13571);
nor U14452 (N_14452,N_13965,N_13941);
xor U14453 (N_14453,N_13564,N_13841);
or U14454 (N_14454,N_13937,N_13894);
xnor U14455 (N_14455,N_13660,N_13628);
nand U14456 (N_14456,N_13954,N_13721);
or U14457 (N_14457,N_13880,N_13605);
nand U14458 (N_14458,N_13966,N_13692);
nand U14459 (N_14459,N_13758,N_13714);
and U14460 (N_14460,N_13971,N_13965);
xnor U14461 (N_14461,N_13942,N_13922);
nand U14462 (N_14462,N_13616,N_13899);
nand U14463 (N_14463,N_13767,N_13654);
nor U14464 (N_14464,N_13535,N_13511);
nand U14465 (N_14465,N_13798,N_13715);
nor U14466 (N_14466,N_13746,N_13656);
nor U14467 (N_14467,N_13605,N_13792);
nor U14468 (N_14468,N_13675,N_13689);
and U14469 (N_14469,N_13901,N_13944);
xor U14470 (N_14470,N_13871,N_13889);
or U14471 (N_14471,N_13976,N_13994);
nor U14472 (N_14472,N_13785,N_13557);
xor U14473 (N_14473,N_13759,N_13977);
nor U14474 (N_14474,N_13640,N_13917);
nand U14475 (N_14475,N_13551,N_13988);
xor U14476 (N_14476,N_13613,N_13660);
nand U14477 (N_14477,N_13878,N_13993);
xnor U14478 (N_14478,N_13839,N_13857);
nand U14479 (N_14479,N_13673,N_13606);
or U14480 (N_14480,N_13709,N_13559);
or U14481 (N_14481,N_13602,N_13692);
xnor U14482 (N_14482,N_13687,N_13858);
nor U14483 (N_14483,N_13530,N_13659);
nor U14484 (N_14484,N_13663,N_13791);
xor U14485 (N_14485,N_13842,N_13953);
xor U14486 (N_14486,N_13949,N_13521);
nor U14487 (N_14487,N_13979,N_13547);
nand U14488 (N_14488,N_13707,N_13687);
nor U14489 (N_14489,N_13861,N_13967);
or U14490 (N_14490,N_13717,N_13800);
nand U14491 (N_14491,N_13693,N_13663);
nor U14492 (N_14492,N_13961,N_13714);
xnor U14493 (N_14493,N_13758,N_13952);
and U14494 (N_14494,N_13792,N_13703);
nor U14495 (N_14495,N_13535,N_13821);
nor U14496 (N_14496,N_13925,N_13796);
or U14497 (N_14497,N_13676,N_13825);
nand U14498 (N_14498,N_13887,N_13928);
nand U14499 (N_14499,N_13994,N_13879);
nor U14500 (N_14500,N_14032,N_14073);
and U14501 (N_14501,N_14445,N_14457);
xnor U14502 (N_14502,N_14115,N_14409);
and U14503 (N_14503,N_14475,N_14487);
nor U14504 (N_14504,N_14103,N_14489);
nor U14505 (N_14505,N_14144,N_14141);
or U14506 (N_14506,N_14434,N_14237);
xor U14507 (N_14507,N_14345,N_14432);
nand U14508 (N_14508,N_14278,N_14132);
xnor U14509 (N_14509,N_14203,N_14366);
nand U14510 (N_14510,N_14136,N_14480);
nor U14511 (N_14511,N_14180,N_14482);
nand U14512 (N_14512,N_14394,N_14182);
xor U14513 (N_14513,N_14191,N_14208);
nor U14514 (N_14514,N_14173,N_14396);
and U14515 (N_14515,N_14397,N_14114);
and U14516 (N_14516,N_14378,N_14327);
and U14517 (N_14517,N_14294,N_14137);
nand U14518 (N_14518,N_14427,N_14408);
nor U14519 (N_14519,N_14304,N_14062);
nand U14520 (N_14520,N_14443,N_14054);
nor U14521 (N_14521,N_14213,N_14298);
and U14522 (N_14522,N_14012,N_14185);
xnor U14523 (N_14523,N_14346,N_14264);
and U14524 (N_14524,N_14448,N_14223);
xor U14525 (N_14525,N_14485,N_14099);
and U14526 (N_14526,N_14260,N_14483);
or U14527 (N_14527,N_14258,N_14139);
xnor U14528 (N_14528,N_14041,N_14051);
or U14529 (N_14529,N_14133,N_14222);
and U14530 (N_14530,N_14497,N_14187);
xor U14531 (N_14531,N_14216,N_14053);
xor U14532 (N_14532,N_14022,N_14492);
nor U14533 (N_14533,N_14117,N_14018);
and U14534 (N_14534,N_14287,N_14416);
nand U14535 (N_14535,N_14240,N_14247);
or U14536 (N_14536,N_14209,N_14046);
or U14537 (N_14537,N_14406,N_14233);
or U14538 (N_14538,N_14077,N_14130);
nand U14539 (N_14539,N_14232,N_14342);
nor U14540 (N_14540,N_14498,N_14276);
xnor U14541 (N_14541,N_14079,N_14039);
and U14542 (N_14542,N_14323,N_14150);
nor U14543 (N_14543,N_14035,N_14403);
or U14544 (N_14544,N_14261,N_14273);
xnor U14545 (N_14545,N_14331,N_14083);
xnor U14546 (N_14546,N_14085,N_14411);
nor U14547 (N_14547,N_14248,N_14379);
and U14548 (N_14548,N_14277,N_14013);
xnor U14549 (N_14549,N_14428,N_14110);
nand U14550 (N_14550,N_14239,N_14329);
and U14551 (N_14551,N_14354,N_14338);
nand U14552 (N_14552,N_14072,N_14412);
nor U14553 (N_14553,N_14337,N_14069);
nor U14554 (N_14554,N_14436,N_14148);
xor U14555 (N_14555,N_14259,N_14332);
and U14556 (N_14556,N_14145,N_14206);
nand U14557 (N_14557,N_14280,N_14179);
nand U14558 (N_14558,N_14372,N_14330);
nand U14559 (N_14559,N_14005,N_14373);
xor U14560 (N_14560,N_14156,N_14387);
nand U14561 (N_14561,N_14101,N_14066);
and U14562 (N_14562,N_14356,N_14135);
or U14563 (N_14563,N_14279,N_14349);
or U14564 (N_14564,N_14300,N_14336);
and U14565 (N_14565,N_14462,N_14149);
nor U14566 (N_14566,N_14036,N_14420);
and U14567 (N_14567,N_14441,N_14493);
nand U14568 (N_14568,N_14451,N_14292);
nand U14569 (N_14569,N_14322,N_14033);
or U14570 (N_14570,N_14168,N_14490);
xor U14571 (N_14571,N_14082,N_14104);
or U14572 (N_14572,N_14312,N_14228);
or U14573 (N_14573,N_14272,N_14175);
xnor U14574 (N_14574,N_14319,N_14418);
nand U14575 (N_14575,N_14170,N_14158);
and U14576 (N_14576,N_14028,N_14153);
nor U14577 (N_14577,N_14391,N_14167);
nor U14578 (N_14578,N_14020,N_14204);
nor U14579 (N_14579,N_14186,N_14318);
and U14580 (N_14580,N_14442,N_14154);
and U14581 (N_14581,N_14320,N_14477);
xor U14582 (N_14582,N_14352,N_14328);
xor U14583 (N_14583,N_14383,N_14389);
xnor U14584 (N_14584,N_14146,N_14159);
nand U14585 (N_14585,N_14230,N_14019);
and U14586 (N_14586,N_14461,N_14061);
or U14587 (N_14587,N_14108,N_14042);
nand U14588 (N_14588,N_14450,N_14290);
or U14589 (N_14589,N_14266,N_14365);
xnor U14590 (N_14590,N_14118,N_14227);
xnor U14591 (N_14591,N_14382,N_14404);
nand U14592 (N_14592,N_14375,N_14121);
nand U14593 (N_14593,N_14415,N_14275);
nand U14594 (N_14594,N_14456,N_14333);
or U14595 (N_14595,N_14089,N_14106);
nand U14596 (N_14596,N_14023,N_14267);
or U14597 (N_14597,N_14401,N_14058);
nand U14598 (N_14598,N_14025,N_14122);
xor U14599 (N_14599,N_14355,N_14009);
and U14600 (N_14600,N_14026,N_14245);
xnor U14601 (N_14601,N_14359,N_14430);
and U14602 (N_14602,N_14126,N_14344);
and U14603 (N_14603,N_14008,N_14016);
and U14604 (N_14604,N_14268,N_14164);
or U14605 (N_14605,N_14453,N_14309);
nand U14606 (N_14606,N_14116,N_14090);
xor U14607 (N_14607,N_14285,N_14241);
or U14608 (N_14608,N_14221,N_14057);
nor U14609 (N_14609,N_14444,N_14274);
nor U14610 (N_14610,N_14015,N_14097);
nor U14611 (N_14611,N_14071,N_14440);
and U14612 (N_14612,N_14219,N_14363);
and U14613 (N_14613,N_14157,N_14447);
xor U14614 (N_14614,N_14211,N_14281);
nor U14615 (N_14615,N_14107,N_14194);
nand U14616 (N_14616,N_14488,N_14439);
xor U14617 (N_14617,N_14305,N_14496);
and U14618 (N_14618,N_14068,N_14120);
and U14619 (N_14619,N_14056,N_14065);
nor U14620 (N_14620,N_14392,N_14289);
nor U14621 (N_14621,N_14459,N_14183);
nor U14622 (N_14622,N_14004,N_14293);
or U14623 (N_14623,N_14399,N_14417);
nor U14624 (N_14624,N_14205,N_14324);
and U14625 (N_14625,N_14210,N_14377);
xnor U14626 (N_14626,N_14295,N_14088);
xnor U14627 (N_14627,N_14226,N_14348);
and U14628 (N_14628,N_14311,N_14171);
or U14629 (N_14629,N_14047,N_14236);
nor U14630 (N_14630,N_14464,N_14184);
and U14631 (N_14631,N_14161,N_14251);
xor U14632 (N_14632,N_14469,N_14043);
and U14633 (N_14633,N_14086,N_14421);
xor U14634 (N_14634,N_14124,N_14393);
xor U14635 (N_14635,N_14384,N_14131);
nor U14636 (N_14636,N_14301,N_14165);
or U14637 (N_14637,N_14339,N_14362);
xnor U14638 (N_14638,N_14231,N_14003);
xor U14639 (N_14639,N_14080,N_14014);
and U14640 (N_14640,N_14081,N_14147);
nand U14641 (N_14641,N_14413,N_14370);
and U14642 (N_14642,N_14040,N_14472);
or U14643 (N_14643,N_14095,N_14166);
nor U14644 (N_14644,N_14437,N_14067);
xor U14645 (N_14645,N_14163,N_14119);
xor U14646 (N_14646,N_14407,N_14495);
nand U14647 (N_14647,N_14325,N_14458);
and U14648 (N_14648,N_14064,N_14162);
or U14649 (N_14649,N_14010,N_14225);
or U14650 (N_14650,N_14195,N_14128);
and U14651 (N_14651,N_14050,N_14102);
and U14652 (N_14652,N_14474,N_14201);
xnor U14653 (N_14653,N_14055,N_14253);
nor U14654 (N_14654,N_14315,N_14151);
nand U14655 (N_14655,N_14484,N_14123);
and U14656 (N_14656,N_14405,N_14341);
nor U14657 (N_14657,N_14246,N_14140);
or U14658 (N_14658,N_14358,N_14006);
nor U14659 (N_14659,N_14143,N_14059);
xnor U14660 (N_14660,N_14419,N_14129);
and U14661 (N_14661,N_14021,N_14265);
nand U14662 (N_14662,N_14321,N_14215);
nor U14663 (N_14663,N_14220,N_14244);
nand U14664 (N_14664,N_14172,N_14369);
xor U14665 (N_14665,N_14371,N_14011);
and U14666 (N_14666,N_14017,N_14217);
and U14667 (N_14667,N_14207,N_14282);
or U14668 (N_14668,N_14092,N_14075);
or U14669 (N_14669,N_14096,N_14486);
xor U14670 (N_14670,N_14422,N_14270);
or U14671 (N_14671,N_14060,N_14283);
xor U14672 (N_14672,N_14463,N_14299);
nor U14673 (N_14673,N_14192,N_14316);
or U14674 (N_14674,N_14198,N_14449);
xnor U14675 (N_14675,N_14094,N_14024);
nand U14676 (N_14676,N_14127,N_14381);
or U14677 (N_14677,N_14313,N_14202);
and U14678 (N_14678,N_14465,N_14380);
or U14679 (N_14679,N_14138,N_14303);
or U14680 (N_14680,N_14160,N_14196);
xor U14681 (N_14681,N_14374,N_14335);
and U14682 (N_14682,N_14425,N_14402);
xor U14683 (N_14683,N_14218,N_14471);
nand U14684 (N_14684,N_14269,N_14134);
nor U14685 (N_14685,N_14476,N_14034);
and U14686 (N_14686,N_14314,N_14200);
nor U14687 (N_14687,N_14340,N_14390);
nand U14688 (N_14688,N_14193,N_14386);
nor U14689 (N_14689,N_14093,N_14357);
xnor U14690 (N_14690,N_14286,N_14031);
nor U14691 (N_14691,N_14385,N_14262);
nor U14692 (N_14692,N_14360,N_14169);
and U14693 (N_14693,N_14326,N_14350);
nand U14694 (N_14694,N_14038,N_14306);
nor U14695 (N_14695,N_14255,N_14334);
nand U14696 (N_14696,N_14431,N_14070);
xnor U14697 (N_14697,N_14291,N_14181);
nor U14698 (N_14698,N_14347,N_14078);
and U14699 (N_14699,N_14473,N_14466);
nand U14700 (N_14700,N_14087,N_14027);
xnor U14701 (N_14701,N_14296,N_14214);
or U14702 (N_14702,N_14176,N_14470);
or U14703 (N_14703,N_14398,N_14455);
or U14704 (N_14704,N_14361,N_14368);
and U14705 (N_14705,N_14307,N_14177);
nor U14706 (N_14706,N_14111,N_14410);
and U14707 (N_14707,N_14109,N_14364);
or U14708 (N_14708,N_14438,N_14100);
and U14709 (N_14709,N_14098,N_14481);
nor U14710 (N_14710,N_14142,N_14288);
xnor U14711 (N_14711,N_14367,N_14284);
or U14712 (N_14712,N_14007,N_14271);
xor U14713 (N_14713,N_14242,N_14343);
xor U14714 (N_14714,N_14435,N_14076);
nor U14715 (N_14715,N_14388,N_14001);
and U14716 (N_14716,N_14091,N_14235);
xnor U14717 (N_14717,N_14454,N_14249);
nand U14718 (N_14718,N_14063,N_14030);
or U14719 (N_14719,N_14254,N_14468);
nand U14720 (N_14720,N_14308,N_14234);
nand U14721 (N_14721,N_14446,N_14460);
xor U14722 (N_14722,N_14224,N_14174);
or U14723 (N_14723,N_14229,N_14238);
and U14724 (N_14724,N_14494,N_14044);
or U14725 (N_14725,N_14048,N_14189);
or U14726 (N_14726,N_14049,N_14029);
nor U14727 (N_14727,N_14152,N_14155);
nand U14728 (N_14728,N_14433,N_14297);
nor U14729 (N_14729,N_14353,N_14252);
nor U14730 (N_14730,N_14000,N_14400);
nor U14731 (N_14731,N_14478,N_14467);
nand U14732 (N_14732,N_14074,N_14105);
nand U14733 (N_14733,N_14256,N_14112);
and U14734 (N_14734,N_14479,N_14424);
nand U14735 (N_14735,N_14499,N_14250);
or U14736 (N_14736,N_14212,N_14310);
and U14737 (N_14737,N_14113,N_14423);
or U14738 (N_14738,N_14084,N_14190);
xnor U14739 (N_14739,N_14351,N_14197);
and U14740 (N_14740,N_14243,N_14178);
and U14741 (N_14741,N_14302,N_14037);
nor U14742 (N_14742,N_14452,N_14199);
nand U14743 (N_14743,N_14376,N_14414);
nand U14744 (N_14744,N_14125,N_14395);
or U14745 (N_14745,N_14263,N_14257);
nand U14746 (N_14746,N_14491,N_14045);
and U14747 (N_14747,N_14426,N_14052);
or U14748 (N_14748,N_14188,N_14002);
or U14749 (N_14749,N_14317,N_14429);
and U14750 (N_14750,N_14043,N_14247);
xor U14751 (N_14751,N_14283,N_14372);
and U14752 (N_14752,N_14065,N_14329);
xnor U14753 (N_14753,N_14450,N_14313);
nor U14754 (N_14754,N_14192,N_14113);
nand U14755 (N_14755,N_14455,N_14355);
xnor U14756 (N_14756,N_14045,N_14157);
and U14757 (N_14757,N_14164,N_14257);
nor U14758 (N_14758,N_14380,N_14201);
or U14759 (N_14759,N_14047,N_14088);
xnor U14760 (N_14760,N_14405,N_14217);
and U14761 (N_14761,N_14372,N_14438);
xnor U14762 (N_14762,N_14177,N_14329);
xnor U14763 (N_14763,N_14132,N_14335);
or U14764 (N_14764,N_14379,N_14255);
nor U14765 (N_14765,N_14116,N_14479);
xor U14766 (N_14766,N_14024,N_14459);
nand U14767 (N_14767,N_14076,N_14129);
or U14768 (N_14768,N_14497,N_14242);
xor U14769 (N_14769,N_14174,N_14089);
or U14770 (N_14770,N_14180,N_14037);
or U14771 (N_14771,N_14434,N_14177);
nand U14772 (N_14772,N_14289,N_14040);
or U14773 (N_14773,N_14204,N_14178);
and U14774 (N_14774,N_14291,N_14240);
nor U14775 (N_14775,N_14477,N_14380);
xnor U14776 (N_14776,N_14011,N_14001);
and U14777 (N_14777,N_14070,N_14191);
nor U14778 (N_14778,N_14458,N_14172);
and U14779 (N_14779,N_14267,N_14397);
and U14780 (N_14780,N_14211,N_14135);
or U14781 (N_14781,N_14235,N_14164);
nor U14782 (N_14782,N_14295,N_14261);
nand U14783 (N_14783,N_14464,N_14374);
and U14784 (N_14784,N_14291,N_14405);
nor U14785 (N_14785,N_14341,N_14151);
xor U14786 (N_14786,N_14062,N_14200);
or U14787 (N_14787,N_14243,N_14210);
xnor U14788 (N_14788,N_14371,N_14384);
and U14789 (N_14789,N_14477,N_14126);
xor U14790 (N_14790,N_14277,N_14420);
nand U14791 (N_14791,N_14437,N_14280);
or U14792 (N_14792,N_14270,N_14447);
nand U14793 (N_14793,N_14345,N_14319);
nor U14794 (N_14794,N_14242,N_14069);
nor U14795 (N_14795,N_14462,N_14233);
nand U14796 (N_14796,N_14065,N_14077);
nand U14797 (N_14797,N_14148,N_14371);
xnor U14798 (N_14798,N_14109,N_14067);
nor U14799 (N_14799,N_14098,N_14135);
xnor U14800 (N_14800,N_14250,N_14485);
nand U14801 (N_14801,N_14204,N_14430);
and U14802 (N_14802,N_14326,N_14183);
nor U14803 (N_14803,N_14241,N_14238);
nor U14804 (N_14804,N_14472,N_14315);
or U14805 (N_14805,N_14072,N_14404);
xor U14806 (N_14806,N_14198,N_14188);
nand U14807 (N_14807,N_14447,N_14295);
nor U14808 (N_14808,N_14221,N_14327);
nand U14809 (N_14809,N_14218,N_14206);
xnor U14810 (N_14810,N_14131,N_14121);
and U14811 (N_14811,N_14472,N_14388);
nand U14812 (N_14812,N_14492,N_14193);
or U14813 (N_14813,N_14411,N_14103);
or U14814 (N_14814,N_14293,N_14285);
and U14815 (N_14815,N_14494,N_14188);
xor U14816 (N_14816,N_14265,N_14284);
or U14817 (N_14817,N_14006,N_14457);
xor U14818 (N_14818,N_14191,N_14085);
nor U14819 (N_14819,N_14364,N_14041);
nand U14820 (N_14820,N_14450,N_14410);
nand U14821 (N_14821,N_14370,N_14421);
or U14822 (N_14822,N_14191,N_14287);
or U14823 (N_14823,N_14002,N_14102);
nand U14824 (N_14824,N_14227,N_14103);
or U14825 (N_14825,N_14035,N_14014);
nor U14826 (N_14826,N_14412,N_14263);
nand U14827 (N_14827,N_14484,N_14349);
nor U14828 (N_14828,N_14216,N_14496);
or U14829 (N_14829,N_14164,N_14204);
or U14830 (N_14830,N_14302,N_14443);
nand U14831 (N_14831,N_14215,N_14019);
xnor U14832 (N_14832,N_14420,N_14331);
and U14833 (N_14833,N_14261,N_14447);
and U14834 (N_14834,N_14097,N_14379);
or U14835 (N_14835,N_14219,N_14483);
nor U14836 (N_14836,N_14372,N_14479);
nor U14837 (N_14837,N_14125,N_14209);
nand U14838 (N_14838,N_14483,N_14330);
xnor U14839 (N_14839,N_14296,N_14309);
nand U14840 (N_14840,N_14393,N_14088);
nor U14841 (N_14841,N_14276,N_14176);
or U14842 (N_14842,N_14411,N_14266);
nor U14843 (N_14843,N_14183,N_14422);
or U14844 (N_14844,N_14354,N_14286);
nand U14845 (N_14845,N_14490,N_14341);
nor U14846 (N_14846,N_14245,N_14331);
xor U14847 (N_14847,N_14124,N_14403);
or U14848 (N_14848,N_14259,N_14441);
or U14849 (N_14849,N_14177,N_14052);
and U14850 (N_14850,N_14326,N_14491);
nand U14851 (N_14851,N_14444,N_14099);
xor U14852 (N_14852,N_14289,N_14198);
and U14853 (N_14853,N_14308,N_14198);
nand U14854 (N_14854,N_14023,N_14075);
or U14855 (N_14855,N_14063,N_14026);
nand U14856 (N_14856,N_14149,N_14152);
nand U14857 (N_14857,N_14056,N_14314);
nor U14858 (N_14858,N_14062,N_14330);
nand U14859 (N_14859,N_14210,N_14356);
nor U14860 (N_14860,N_14212,N_14267);
and U14861 (N_14861,N_14390,N_14362);
or U14862 (N_14862,N_14348,N_14349);
nand U14863 (N_14863,N_14011,N_14462);
xor U14864 (N_14864,N_14301,N_14396);
nor U14865 (N_14865,N_14083,N_14299);
nor U14866 (N_14866,N_14293,N_14046);
nand U14867 (N_14867,N_14393,N_14397);
nand U14868 (N_14868,N_14167,N_14320);
nor U14869 (N_14869,N_14009,N_14335);
and U14870 (N_14870,N_14022,N_14293);
nand U14871 (N_14871,N_14005,N_14037);
nand U14872 (N_14872,N_14483,N_14018);
xor U14873 (N_14873,N_14391,N_14221);
nor U14874 (N_14874,N_14007,N_14265);
and U14875 (N_14875,N_14000,N_14249);
nand U14876 (N_14876,N_14425,N_14050);
and U14877 (N_14877,N_14032,N_14150);
and U14878 (N_14878,N_14364,N_14071);
xnor U14879 (N_14879,N_14098,N_14386);
xnor U14880 (N_14880,N_14133,N_14143);
nand U14881 (N_14881,N_14083,N_14128);
nand U14882 (N_14882,N_14406,N_14184);
nor U14883 (N_14883,N_14077,N_14474);
or U14884 (N_14884,N_14397,N_14222);
xnor U14885 (N_14885,N_14168,N_14408);
and U14886 (N_14886,N_14239,N_14264);
and U14887 (N_14887,N_14298,N_14455);
nand U14888 (N_14888,N_14374,N_14107);
nand U14889 (N_14889,N_14325,N_14056);
and U14890 (N_14890,N_14427,N_14215);
nand U14891 (N_14891,N_14295,N_14132);
or U14892 (N_14892,N_14018,N_14390);
or U14893 (N_14893,N_14476,N_14247);
or U14894 (N_14894,N_14315,N_14277);
and U14895 (N_14895,N_14168,N_14092);
xor U14896 (N_14896,N_14375,N_14152);
or U14897 (N_14897,N_14298,N_14429);
nand U14898 (N_14898,N_14497,N_14256);
and U14899 (N_14899,N_14197,N_14232);
and U14900 (N_14900,N_14084,N_14027);
nor U14901 (N_14901,N_14430,N_14147);
and U14902 (N_14902,N_14300,N_14326);
xnor U14903 (N_14903,N_14311,N_14391);
nand U14904 (N_14904,N_14468,N_14152);
nand U14905 (N_14905,N_14241,N_14491);
and U14906 (N_14906,N_14083,N_14017);
xnor U14907 (N_14907,N_14096,N_14126);
nand U14908 (N_14908,N_14053,N_14143);
xor U14909 (N_14909,N_14473,N_14089);
and U14910 (N_14910,N_14435,N_14142);
xor U14911 (N_14911,N_14349,N_14055);
xnor U14912 (N_14912,N_14241,N_14358);
nand U14913 (N_14913,N_14369,N_14448);
nor U14914 (N_14914,N_14163,N_14203);
nor U14915 (N_14915,N_14049,N_14214);
nand U14916 (N_14916,N_14052,N_14204);
xnor U14917 (N_14917,N_14027,N_14294);
or U14918 (N_14918,N_14271,N_14027);
nor U14919 (N_14919,N_14475,N_14230);
or U14920 (N_14920,N_14259,N_14132);
and U14921 (N_14921,N_14372,N_14249);
nand U14922 (N_14922,N_14108,N_14461);
or U14923 (N_14923,N_14399,N_14019);
or U14924 (N_14924,N_14152,N_14313);
and U14925 (N_14925,N_14453,N_14361);
nor U14926 (N_14926,N_14435,N_14487);
nand U14927 (N_14927,N_14231,N_14472);
xnor U14928 (N_14928,N_14021,N_14273);
or U14929 (N_14929,N_14195,N_14141);
or U14930 (N_14930,N_14005,N_14315);
and U14931 (N_14931,N_14407,N_14224);
xor U14932 (N_14932,N_14363,N_14126);
xnor U14933 (N_14933,N_14091,N_14208);
nor U14934 (N_14934,N_14123,N_14363);
nand U14935 (N_14935,N_14262,N_14216);
nor U14936 (N_14936,N_14065,N_14255);
nand U14937 (N_14937,N_14137,N_14306);
nand U14938 (N_14938,N_14111,N_14331);
and U14939 (N_14939,N_14146,N_14387);
nor U14940 (N_14940,N_14214,N_14410);
xor U14941 (N_14941,N_14309,N_14086);
nand U14942 (N_14942,N_14018,N_14206);
nand U14943 (N_14943,N_14089,N_14263);
xnor U14944 (N_14944,N_14314,N_14048);
nand U14945 (N_14945,N_14386,N_14474);
nor U14946 (N_14946,N_14304,N_14450);
nor U14947 (N_14947,N_14061,N_14328);
and U14948 (N_14948,N_14169,N_14282);
or U14949 (N_14949,N_14314,N_14404);
or U14950 (N_14950,N_14485,N_14420);
nor U14951 (N_14951,N_14386,N_14017);
or U14952 (N_14952,N_14414,N_14477);
and U14953 (N_14953,N_14325,N_14480);
nand U14954 (N_14954,N_14222,N_14453);
xnor U14955 (N_14955,N_14082,N_14419);
xor U14956 (N_14956,N_14277,N_14279);
or U14957 (N_14957,N_14147,N_14309);
nand U14958 (N_14958,N_14332,N_14264);
or U14959 (N_14959,N_14226,N_14416);
nor U14960 (N_14960,N_14287,N_14462);
nand U14961 (N_14961,N_14411,N_14174);
nand U14962 (N_14962,N_14408,N_14036);
xnor U14963 (N_14963,N_14232,N_14340);
or U14964 (N_14964,N_14336,N_14467);
or U14965 (N_14965,N_14289,N_14429);
and U14966 (N_14966,N_14174,N_14441);
nor U14967 (N_14967,N_14342,N_14222);
or U14968 (N_14968,N_14446,N_14392);
nand U14969 (N_14969,N_14292,N_14042);
nor U14970 (N_14970,N_14484,N_14010);
and U14971 (N_14971,N_14190,N_14496);
nor U14972 (N_14972,N_14343,N_14272);
and U14973 (N_14973,N_14255,N_14151);
nor U14974 (N_14974,N_14219,N_14067);
or U14975 (N_14975,N_14167,N_14053);
xnor U14976 (N_14976,N_14211,N_14186);
nand U14977 (N_14977,N_14186,N_14051);
or U14978 (N_14978,N_14104,N_14195);
xnor U14979 (N_14979,N_14017,N_14279);
or U14980 (N_14980,N_14345,N_14362);
or U14981 (N_14981,N_14439,N_14121);
and U14982 (N_14982,N_14367,N_14094);
or U14983 (N_14983,N_14319,N_14474);
xnor U14984 (N_14984,N_14088,N_14006);
nor U14985 (N_14985,N_14324,N_14464);
nand U14986 (N_14986,N_14094,N_14362);
nand U14987 (N_14987,N_14387,N_14410);
or U14988 (N_14988,N_14462,N_14217);
nand U14989 (N_14989,N_14239,N_14419);
xor U14990 (N_14990,N_14252,N_14089);
xor U14991 (N_14991,N_14154,N_14040);
nor U14992 (N_14992,N_14004,N_14491);
nor U14993 (N_14993,N_14194,N_14172);
xnor U14994 (N_14994,N_14431,N_14071);
and U14995 (N_14995,N_14426,N_14308);
nor U14996 (N_14996,N_14258,N_14375);
or U14997 (N_14997,N_14108,N_14250);
or U14998 (N_14998,N_14182,N_14071);
nand U14999 (N_14999,N_14204,N_14100);
nand U15000 (N_15000,N_14652,N_14785);
or U15001 (N_15001,N_14943,N_14853);
xor U15002 (N_15002,N_14631,N_14535);
nand U15003 (N_15003,N_14957,N_14705);
nor U15004 (N_15004,N_14677,N_14735);
nand U15005 (N_15005,N_14789,N_14638);
nor U15006 (N_15006,N_14841,N_14547);
and U15007 (N_15007,N_14592,N_14665);
xnor U15008 (N_15008,N_14920,N_14738);
and U15009 (N_15009,N_14594,N_14828);
or U15010 (N_15010,N_14784,N_14777);
nand U15011 (N_15011,N_14668,N_14800);
nand U15012 (N_15012,N_14575,N_14848);
or U15013 (N_15013,N_14513,N_14769);
xnor U15014 (N_15014,N_14707,N_14565);
nand U15015 (N_15015,N_14952,N_14823);
or U15016 (N_15016,N_14775,N_14561);
nor U15017 (N_15017,N_14704,N_14948);
xor U15018 (N_15018,N_14545,N_14574);
nand U15019 (N_15019,N_14696,N_14980);
xor U15020 (N_15020,N_14583,N_14622);
and U15021 (N_15021,N_14995,N_14596);
or U15022 (N_15022,N_14601,N_14693);
nand U15023 (N_15023,N_14660,N_14960);
nand U15024 (N_15024,N_14883,N_14718);
and U15025 (N_15025,N_14849,N_14699);
nand U15026 (N_15026,N_14826,N_14947);
and U15027 (N_15027,N_14959,N_14517);
xor U15028 (N_15028,N_14658,N_14835);
or U15029 (N_15029,N_14595,N_14781);
nand U15030 (N_15030,N_14931,N_14940);
and U15031 (N_15031,N_14743,N_14540);
xnor U15032 (N_15032,N_14766,N_14905);
or U15033 (N_15033,N_14512,N_14926);
or U15034 (N_15034,N_14793,N_14556);
or U15035 (N_15035,N_14861,N_14670);
nand U15036 (N_15036,N_14589,N_14749);
xnor U15037 (N_15037,N_14951,N_14701);
xor U15038 (N_15038,N_14974,N_14962);
xor U15039 (N_15039,N_14868,N_14520);
nor U15040 (N_15040,N_14662,N_14822);
nor U15041 (N_15041,N_14770,N_14754);
or U15042 (N_15042,N_14998,N_14579);
and U15043 (N_15043,N_14802,N_14756);
and U15044 (N_15044,N_14993,N_14873);
xor U15045 (N_15045,N_14879,N_14702);
and U15046 (N_15046,N_14772,N_14641);
and U15047 (N_15047,N_14695,N_14809);
and U15048 (N_15048,N_14676,N_14916);
nand U15049 (N_15049,N_14903,N_14613);
nand U15050 (N_15050,N_14503,N_14944);
xnor U15051 (N_15051,N_14642,N_14746);
xor U15052 (N_15052,N_14570,N_14939);
xnor U15053 (N_15053,N_14724,N_14663);
nor U15054 (N_15054,N_14888,N_14634);
or U15055 (N_15055,N_14831,N_14630);
and U15056 (N_15056,N_14914,N_14618);
and U15057 (N_15057,N_14913,N_14633);
xor U15058 (N_15058,N_14605,N_14505);
xor U15059 (N_15059,N_14874,N_14902);
nor U15060 (N_15060,N_14682,N_14846);
xor U15061 (N_15061,N_14640,N_14965);
nor U15062 (N_15062,N_14946,N_14813);
or U15063 (N_15063,N_14655,N_14921);
xor U15064 (N_15064,N_14697,N_14564);
nand U15065 (N_15065,N_14824,N_14533);
nand U15066 (N_15066,N_14741,N_14686);
xor U15067 (N_15067,N_14563,N_14719);
xor U15068 (N_15068,N_14967,N_14576);
xor U15069 (N_15069,N_14804,N_14996);
xor U15070 (N_15070,N_14657,N_14982);
or U15071 (N_15071,N_14562,N_14765);
nand U15072 (N_15072,N_14710,N_14681);
and U15073 (N_15073,N_14790,N_14593);
and U15074 (N_15074,N_14643,N_14830);
nand U15075 (N_15075,N_14786,N_14977);
or U15076 (N_15076,N_14591,N_14821);
and U15077 (N_15077,N_14684,N_14907);
or U15078 (N_15078,N_14552,N_14623);
and U15079 (N_15079,N_14884,N_14852);
or U15080 (N_15080,N_14997,N_14541);
nand U15081 (N_15081,N_14698,N_14610);
or U15082 (N_15082,N_14598,N_14581);
nand U15083 (N_15083,N_14530,N_14508);
xnor U15084 (N_15084,N_14843,N_14712);
nor U15085 (N_15085,N_14742,N_14901);
nand U15086 (N_15086,N_14838,N_14787);
xnor U15087 (N_15087,N_14871,N_14891);
nor U15088 (N_15088,N_14968,N_14609);
nor U15089 (N_15089,N_14569,N_14555);
or U15090 (N_15090,N_14788,N_14827);
and U15091 (N_15091,N_14644,N_14970);
nor U15092 (N_15092,N_14893,N_14619);
or U15093 (N_15093,N_14900,N_14971);
or U15094 (N_15094,N_14854,N_14509);
xnor U15095 (N_15095,N_14524,N_14715);
nand U15096 (N_15096,N_14616,N_14934);
or U15097 (N_15097,N_14966,N_14600);
and U15098 (N_15098,N_14910,N_14653);
nand U15099 (N_15099,N_14981,N_14805);
or U15100 (N_15100,N_14727,N_14878);
and U15101 (N_15101,N_14812,N_14526);
nand U15102 (N_15102,N_14708,N_14627);
or U15103 (N_15103,N_14674,N_14506);
or U15104 (N_15104,N_14529,N_14932);
xor U15105 (N_15105,N_14956,N_14961);
nand U15106 (N_15106,N_14799,N_14829);
or U15107 (N_15107,N_14645,N_14776);
nand U15108 (N_15108,N_14647,N_14625);
nor U15109 (N_15109,N_14502,N_14978);
and U15110 (N_15110,N_14604,N_14732);
xor U15111 (N_15111,N_14842,N_14935);
nor U15112 (N_15112,N_14679,N_14716);
or U15113 (N_15113,N_14837,N_14811);
nand U15114 (N_15114,N_14882,N_14937);
and U15115 (N_15115,N_14689,N_14528);
and U15116 (N_15116,N_14534,N_14791);
nor U15117 (N_15117,N_14985,N_14938);
xnor U15118 (N_15118,N_14761,N_14872);
nand U15119 (N_15119,N_14875,N_14651);
nand U15120 (N_15120,N_14906,N_14758);
nor U15121 (N_15121,N_14990,N_14845);
nand U15122 (N_15122,N_14771,N_14796);
and U15123 (N_15123,N_14709,N_14825);
nor U15124 (N_15124,N_14975,N_14685);
or U15125 (N_15125,N_14514,N_14984);
or U15126 (N_15126,N_14515,N_14654);
xor U15127 (N_15127,N_14930,N_14726);
or U15128 (N_15128,N_14673,N_14737);
nor U15129 (N_15129,N_14942,N_14582);
and U15130 (N_15130,N_14539,N_14700);
nand U15131 (N_15131,N_14904,N_14869);
nor U15132 (N_15132,N_14887,N_14923);
nand U15133 (N_15133,N_14611,N_14850);
nand U15134 (N_15134,N_14714,N_14606);
and U15135 (N_15135,N_14646,N_14991);
and U15136 (N_15136,N_14972,N_14553);
xnor U15137 (N_15137,N_14692,N_14624);
nor U15138 (N_15138,N_14894,N_14566);
or U15139 (N_15139,N_14747,N_14860);
and U15140 (N_15140,N_14744,N_14635);
nand U15141 (N_15141,N_14585,N_14818);
nand U15142 (N_15142,N_14885,N_14554);
and U15143 (N_15143,N_14759,N_14936);
nor U15144 (N_15144,N_14723,N_14763);
xnor U15145 (N_15145,N_14537,N_14892);
nor U15146 (N_15146,N_14858,N_14527);
nand U15147 (N_15147,N_14953,N_14865);
nor U15148 (N_15148,N_14602,N_14917);
xor U15149 (N_15149,N_14637,N_14855);
or U15150 (N_15150,N_14798,N_14748);
xor U15151 (N_15151,N_14706,N_14745);
nand U15152 (N_15152,N_14750,N_14820);
nand U15153 (N_15153,N_14507,N_14736);
nor U15154 (N_15154,N_14740,N_14979);
xor U15155 (N_15155,N_14896,N_14927);
nand U15156 (N_15156,N_14797,N_14794);
or U15157 (N_15157,N_14510,N_14546);
nand U15158 (N_15158,N_14832,N_14929);
or U15159 (N_15159,N_14801,N_14661);
nand U15160 (N_15160,N_14973,N_14538);
xor U15161 (N_15161,N_14964,N_14728);
and U15162 (N_15162,N_14857,N_14558);
and U15163 (N_15163,N_14525,N_14833);
or U15164 (N_15164,N_14739,N_14544);
nor U15165 (N_15165,N_14992,N_14816);
nand U15166 (N_15166,N_14880,N_14925);
or U15167 (N_15167,N_14950,N_14612);
nand U15168 (N_15168,N_14667,N_14721);
nand U15169 (N_15169,N_14963,N_14792);
nand U15170 (N_15170,N_14577,N_14683);
xnor U15171 (N_15171,N_14680,N_14753);
and U15172 (N_15172,N_14751,N_14919);
nand U15173 (N_15173,N_14599,N_14994);
xnor U15174 (N_15174,N_14877,N_14863);
or U15175 (N_15175,N_14649,N_14531);
nand U15176 (N_15176,N_14779,N_14572);
nand U15177 (N_15177,N_14620,N_14840);
xor U15178 (N_15178,N_14608,N_14976);
nor U15179 (N_15179,N_14899,N_14851);
xor U15180 (N_15180,N_14767,N_14958);
and U15181 (N_15181,N_14725,N_14607);
nand U15182 (N_15182,N_14729,N_14519);
xor U15183 (N_15183,N_14983,N_14690);
nand U15184 (N_15184,N_14722,N_14551);
or U15185 (N_15185,N_14881,N_14752);
xor U15186 (N_15186,N_14780,N_14819);
or U15187 (N_15187,N_14889,N_14941);
nor U15188 (N_15188,N_14694,N_14839);
xor U15189 (N_15189,N_14500,N_14678);
and U15190 (N_15190,N_14542,N_14870);
and U15191 (N_15191,N_14656,N_14867);
or U15192 (N_15192,N_14803,N_14617);
xnor U15193 (N_15193,N_14669,N_14518);
and U15194 (N_15194,N_14588,N_14999);
or U15195 (N_15195,N_14650,N_14626);
or U15196 (N_15196,N_14762,N_14560);
and U15197 (N_15197,N_14720,N_14734);
nand U15198 (N_15198,N_14757,N_14774);
nor U15199 (N_15199,N_14664,N_14717);
and U15200 (N_15200,N_14549,N_14671);
xor U15201 (N_15201,N_14504,N_14987);
nand U15202 (N_15202,N_14532,N_14989);
xnor U15203 (N_15203,N_14814,N_14703);
nor U15204 (N_15204,N_14621,N_14688);
nor U15205 (N_15205,N_14543,N_14639);
nand U15206 (N_15206,N_14856,N_14586);
and U15207 (N_15207,N_14807,N_14578);
or U15208 (N_15208,N_14876,N_14988);
and U15209 (N_15209,N_14886,N_14628);
xor U15210 (N_15210,N_14928,N_14768);
and U15211 (N_15211,N_14580,N_14636);
nor U15212 (N_15212,N_14864,N_14522);
nor U15213 (N_15213,N_14969,N_14713);
and U15214 (N_15214,N_14687,N_14986);
nor U15215 (N_15215,N_14590,N_14922);
and U15216 (N_15216,N_14632,N_14711);
and U15217 (N_15217,N_14773,N_14815);
nor U15218 (N_15218,N_14795,N_14890);
xnor U15219 (N_15219,N_14949,N_14844);
xor U15220 (N_15220,N_14516,N_14659);
and U15221 (N_15221,N_14523,N_14808);
nand U15222 (N_15222,N_14918,N_14666);
nor U15223 (N_15223,N_14755,N_14862);
nor U15224 (N_15224,N_14836,N_14782);
nor U15225 (N_15225,N_14760,N_14675);
nand U15226 (N_15226,N_14730,N_14648);
xnor U15227 (N_15227,N_14817,N_14568);
or U15228 (N_15228,N_14603,N_14629);
nand U15229 (N_15229,N_14909,N_14898);
nand U15230 (N_15230,N_14615,N_14955);
nand U15231 (N_15231,N_14806,N_14933);
or U15232 (N_15232,N_14521,N_14672);
nand U15233 (N_15233,N_14536,N_14614);
xnor U15234 (N_15234,N_14908,N_14810);
nand U15235 (N_15235,N_14691,N_14567);
nand U15236 (N_15236,N_14847,N_14733);
nand U15237 (N_15237,N_14778,N_14866);
xnor U15238 (N_15238,N_14783,N_14550);
or U15239 (N_15239,N_14557,N_14511);
or U15240 (N_15240,N_14731,N_14834);
and U15241 (N_15241,N_14912,N_14915);
nor U15242 (N_15242,N_14895,N_14945);
and U15243 (N_15243,N_14597,N_14573);
nand U15244 (N_15244,N_14571,N_14587);
nand U15245 (N_15245,N_14548,N_14954);
and U15246 (N_15246,N_14911,N_14859);
or U15247 (N_15247,N_14897,N_14559);
or U15248 (N_15248,N_14501,N_14764);
nand U15249 (N_15249,N_14924,N_14584);
nor U15250 (N_15250,N_14556,N_14740);
xor U15251 (N_15251,N_14567,N_14991);
and U15252 (N_15252,N_14715,N_14749);
xnor U15253 (N_15253,N_14684,N_14652);
xnor U15254 (N_15254,N_14598,N_14645);
xnor U15255 (N_15255,N_14757,N_14965);
and U15256 (N_15256,N_14738,N_14983);
or U15257 (N_15257,N_14793,N_14560);
nor U15258 (N_15258,N_14891,N_14829);
xor U15259 (N_15259,N_14730,N_14812);
nor U15260 (N_15260,N_14981,N_14776);
nand U15261 (N_15261,N_14925,N_14863);
and U15262 (N_15262,N_14840,N_14781);
nand U15263 (N_15263,N_14818,N_14842);
nor U15264 (N_15264,N_14835,N_14768);
xor U15265 (N_15265,N_14592,N_14800);
nand U15266 (N_15266,N_14530,N_14607);
nor U15267 (N_15267,N_14806,N_14567);
and U15268 (N_15268,N_14667,N_14625);
xor U15269 (N_15269,N_14731,N_14940);
or U15270 (N_15270,N_14732,N_14871);
or U15271 (N_15271,N_14859,N_14639);
or U15272 (N_15272,N_14599,N_14578);
nor U15273 (N_15273,N_14905,N_14564);
xor U15274 (N_15274,N_14976,N_14632);
nor U15275 (N_15275,N_14738,N_14630);
or U15276 (N_15276,N_14690,N_14854);
nand U15277 (N_15277,N_14575,N_14977);
or U15278 (N_15278,N_14564,N_14616);
nor U15279 (N_15279,N_14701,N_14942);
and U15280 (N_15280,N_14818,N_14534);
nand U15281 (N_15281,N_14887,N_14662);
and U15282 (N_15282,N_14814,N_14860);
nor U15283 (N_15283,N_14914,N_14663);
and U15284 (N_15284,N_14859,N_14700);
nand U15285 (N_15285,N_14958,N_14792);
and U15286 (N_15286,N_14757,N_14787);
or U15287 (N_15287,N_14551,N_14622);
and U15288 (N_15288,N_14837,N_14600);
nand U15289 (N_15289,N_14526,N_14975);
or U15290 (N_15290,N_14896,N_14799);
nand U15291 (N_15291,N_14696,N_14765);
nand U15292 (N_15292,N_14797,N_14635);
or U15293 (N_15293,N_14557,N_14859);
xnor U15294 (N_15294,N_14578,N_14583);
nand U15295 (N_15295,N_14951,N_14915);
nand U15296 (N_15296,N_14789,N_14767);
and U15297 (N_15297,N_14555,N_14510);
and U15298 (N_15298,N_14524,N_14701);
xnor U15299 (N_15299,N_14589,N_14653);
and U15300 (N_15300,N_14937,N_14863);
nand U15301 (N_15301,N_14538,N_14779);
nor U15302 (N_15302,N_14874,N_14900);
xnor U15303 (N_15303,N_14625,N_14650);
and U15304 (N_15304,N_14680,N_14630);
xnor U15305 (N_15305,N_14670,N_14613);
or U15306 (N_15306,N_14694,N_14908);
and U15307 (N_15307,N_14786,N_14903);
or U15308 (N_15308,N_14776,N_14504);
nand U15309 (N_15309,N_14807,N_14792);
and U15310 (N_15310,N_14742,N_14970);
xnor U15311 (N_15311,N_14931,N_14884);
xor U15312 (N_15312,N_14988,N_14526);
nor U15313 (N_15313,N_14582,N_14777);
and U15314 (N_15314,N_14720,N_14861);
nor U15315 (N_15315,N_14791,N_14971);
nor U15316 (N_15316,N_14807,N_14919);
nor U15317 (N_15317,N_14500,N_14666);
xnor U15318 (N_15318,N_14828,N_14630);
nand U15319 (N_15319,N_14742,N_14814);
or U15320 (N_15320,N_14700,N_14780);
xor U15321 (N_15321,N_14752,N_14910);
nand U15322 (N_15322,N_14681,N_14962);
xnor U15323 (N_15323,N_14594,N_14638);
nor U15324 (N_15324,N_14924,N_14755);
xnor U15325 (N_15325,N_14860,N_14831);
and U15326 (N_15326,N_14769,N_14565);
and U15327 (N_15327,N_14680,N_14702);
or U15328 (N_15328,N_14835,N_14885);
nor U15329 (N_15329,N_14824,N_14610);
or U15330 (N_15330,N_14594,N_14537);
or U15331 (N_15331,N_14712,N_14946);
nor U15332 (N_15332,N_14870,N_14558);
xor U15333 (N_15333,N_14763,N_14919);
nand U15334 (N_15334,N_14936,N_14809);
xnor U15335 (N_15335,N_14873,N_14702);
xor U15336 (N_15336,N_14527,N_14885);
or U15337 (N_15337,N_14603,N_14812);
nor U15338 (N_15338,N_14997,N_14565);
xnor U15339 (N_15339,N_14841,N_14712);
nor U15340 (N_15340,N_14972,N_14674);
xnor U15341 (N_15341,N_14716,N_14750);
nand U15342 (N_15342,N_14510,N_14807);
nand U15343 (N_15343,N_14699,N_14926);
xnor U15344 (N_15344,N_14695,N_14988);
nor U15345 (N_15345,N_14701,N_14617);
or U15346 (N_15346,N_14831,N_14512);
xor U15347 (N_15347,N_14797,N_14713);
and U15348 (N_15348,N_14584,N_14556);
and U15349 (N_15349,N_14867,N_14577);
and U15350 (N_15350,N_14730,N_14500);
nor U15351 (N_15351,N_14663,N_14814);
and U15352 (N_15352,N_14645,N_14918);
xnor U15353 (N_15353,N_14753,N_14808);
nand U15354 (N_15354,N_14904,N_14631);
and U15355 (N_15355,N_14806,N_14896);
nand U15356 (N_15356,N_14861,N_14793);
nand U15357 (N_15357,N_14641,N_14619);
nor U15358 (N_15358,N_14948,N_14537);
xor U15359 (N_15359,N_14776,N_14951);
nor U15360 (N_15360,N_14508,N_14879);
xor U15361 (N_15361,N_14941,N_14872);
nor U15362 (N_15362,N_14938,N_14780);
xor U15363 (N_15363,N_14669,N_14923);
xnor U15364 (N_15364,N_14844,N_14544);
or U15365 (N_15365,N_14978,N_14547);
xnor U15366 (N_15366,N_14701,N_14916);
xnor U15367 (N_15367,N_14665,N_14772);
nor U15368 (N_15368,N_14924,N_14919);
nor U15369 (N_15369,N_14863,N_14769);
or U15370 (N_15370,N_14604,N_14898);
xor U15371 (N_15371,N_14944,N_14634);
or U15372 (N_15372,N_14991,N_14928);
nand U15373 (N_15373,N_14706,N_14879);
nand U15374 (N_15374,N_14780,N_14967);
xor U15375 (N_15375,N_14620,N_14993);
xor U15376 (N_15376,N_14576,N_14715);
nor U15377 (N_15377,N_14622,N_14868);
and U15378 (N_15378,N_14918,N_14565);
and U15379 (N_15379,N_14949,N_14989);
and U15380 (N_15380,N_14782,N_14835);
or U15381 (N_15381,N_14709,N_14814);
nor U15382 (N_15382,N_14999,N_14512);
xor U15383 (N_15383,N_14908,N_14571);
nand U15384 (N_15384,N_14916,N_14956);
nor U15385 (N_15385,N_14693,N_14618);
and U15386 (N_15386,N_14798,N_14673);
or U15387 (N_15387,N_14723,N_14634);
xor U15388 (N_15388,N_14551,N_14626);
xor U15389 (N_15389,N_14786,N_14919);
nor U15390 (N_15390,N_14901,N_14948);
nor U15391 (N_15391,N_14788,N_14592);
nor U15392 (N_15392,N_14785,N_14748);
or U15393 (N_15393,N_14737,N_14860);
and U15394 (N_15394,N_14948,N_14871);
or U15395 (N_15395,N_14949,N_14944);
xnor U15396 (N_15396,N_14622,N_14539);
nor U15397 (N_15397,N_14545,N_14880);
nand U15398 (N_15398,N_14763,N_14953);
nand U15399 (N_15399,N_14613,N_14789);
nor U15400 (N_15400,N_14946,N_14819);
nor U15401 (N_15401,N_14640,N_14943);
or U15402 (N_15402,N_14731,N_14723);
nand U15403 (N_15403,N_14882,N_14572);
xnor U15404 (N_15404,N_14639,N_14946);
nor U15405 (N_15405,N_14760,N_14788);
and U15406 (N_15406,N_14747,N_14763);
xnor U15407 (N_15407,N_14605,N_14810);
xnor U15408 (N_15408,N_14714,N_14506);
nand U15409 (N_15409,N_14662,N_14935);
nor U15410 (N_15410,N_14969,N_14872);
or U15411 (N_15411,N_14852,N_14795);
or U15412 (N_15412,N_14665,N_14510);
nor U15413 (N_15413,N_14720,N_14664);
nor U15414 (N_15414,N_14645,N_14538);
nand U15415 (N_15415,N_14745,N_14609);
xor U15416 (N_15416,N_14625,N_14934);
nand U15417 (N_15417,N_14631,N_14967);
or U15418 (N_15418,N_14519,N_14734);
nor U15419 (N_15419,N_14777,N_14900);
or U15420 (N_15420,N_14912,N_14995);
nor U15421 (N_15421,N_14533,N_14765);
nor U15422 (N_15422,N_14814,N_14506);
nand U15423 (N_15423,N_14946,N_14648);
nand U15424 (N_15424,N_14617,N_14577);
nand U15425 (N_15425,N_14733,N_14986);
xor U15426 (N_15426,N_14996,N_14852);
or U15427 (N_15427,N_14716,N_14904);
nor U15428 (N_15428,N_14797,N_14936);
or U15429 (N_15429,N_14940,N_14849);
or U15430 (N_15430,N_14575,N_14503);
or U15431 (N_15431,N_14869,N_14834);
and U15432 (N_15432,N_14569,N_14733);
and U15433 (N_15433,N_14910,N_14644);
and U15434 (N_15434,N_14986,N_14511);
xor U15435 (N_15435,N_14501,N_14782);
or U15436 (N_15436,N_14831,N_14741);
xnor U15437 (N_15437,N_14836,N_14997);
or U15438 (N_15438,N_14970,N_14874);
and U15439 (N_15439,N_14947,N_14979);
nor U15440 (N_15440,N_14859,N_14783);
nor U15441 (N_15441,N_14852,N_14791);
nor U15442 (N_15442,N_14645,N_14859);
and U15443 (N_15443,N_14579,N_14626);
and U15444 (N_15444,N_14857,N_14716);
or U15445 (N_15445,N_14943,N_14895);
or U15446 (N_15446,N_14918,N_14816);
and U15447 (N_15447,N_14536,N_14860);
xor U15448 (N_15448,N_14529,N_14952);
nand U15449 (N_15449,N_14876,N_14903);
xnor U15450 (N_15450,N_14977,N_14626);
or U15451 (N_15451,N_14967,N_14696);
and U15452 (N_15452,N_14652,N_14808);
xnor U15453 (N_15453,N_14808,N_14530);
nand U15454 (N_15454,N_14662,N_14624);
xnor U15455 (N_15455,N_14679,N_14576);
nor U15456 (N_15456,N_14607,N_14641);
or U15457 (N_15457,N_14975,N_14809);
xor U15458 (N_15458,N_14721,N_14502);
or U15459 (N_15459,N_14579,N_14549);
xnor U15460 (N_15460,N_14574,N_14923);
nor U15461 (N_15461,N_14985,N_14719);
nor U15462 (N_15462,N_14833,N_14565);
xnor U15463 (N_15463,N_14692,N_14836);
and U15464 (N_15464,N_14743,N_14931);
xor U15465 (N_15465,N_14755,N_14639);
nand U15466 (N_15466,N_14927,N_14903);
nand U15467 (N_15467,N_14953,N_14527);
xnor U15468 (N_15468,N_14507,N_14806);
nand U15469 (N_15469,N_14864,N_14800);
or U15470 (N_15470,N_14532,N_14669);
and U15471 (N_15471,N_14513,N_14727);
nor U15472 (N_15472,N_14525,N_14590);
nor U15473 (N_15473,N_14873,N_14870);
nand U15474 (N_15474,N_14756,N_14924);
or U15475 (N_15475,N_14669,N_14776);
and U15476 (N_15476,N_14803,N_14698);
and U15477 (N_15477,N_14637,N_14563);
and U15478 (N_15478,N_14790,N_14679);
nor U15479 (N_15479,N_14784,N_14713);
xnor U15480 (N_15480,N_14695,N_14880);
nor U15481 (N_15481,N_14606,N_14849);
or U15482 (N_15482,N_14811,N_14859);
and U15483 (N_15483,N_14855,N_14682);
or U15484 (N_15484,N_14568,N_14831);
or U15485 (N_15485,N_14819,N_14537);
nor U15486 (N_15486,N_14784,N_14907);
xor U15487 (N_15487,N_14659,N_14756);
xnor U15488 (N_15488,N_14816,N_14985);
nor U15489 (N_15489,N_14993,N_14626);
or U15490 (N_15490,N_14893,N_14767);
xor U15491 (N_15491,N_14820,N_14931);
or U15492 (N_15492,N_14670,N_14671);
and U15493 (N_15493,N_14978,N_14578);
and U15494 (N_15494,N_14840,N_14652);
and U15495 (N_15495,N_14962,N_14960);
xor U15496 (N_15496,N_14679,N_14683);
nand U15497 (N_15497,N_14582,N_14837);
or U15498 (N_15498,N_14890,N_14792);
or U15499 (N_15499,N_14796,N_14516);
or U15500 (N_15500,N_15371,N_15083);
nand U15501 (N_15501,N_15067,N_15193);
and U15502 (N_15502,N_15435,N_15120);
xnor U15503 (N_15503,N_15122,N_15298);
or U15504 (N_15504,N_15150,N_15463);
nand U15505 (N_15505,N_15235,N_15064);
xor U15506 (N_15506,N_15207,N_15455);
and U15507 (N_15507,N_15114,N_15495);
nor U15508 (N_15508,N_15348,N_15284);
nor U15509 (N_15509,N_15351,N_15256);
and U15510 (N_15510,N_15418,N_15221);
nor U15511 (N_15511,N_15299,N_15010);
and U15512 (N_15512,N_15433,N_15198);
or U15513 (N_15513,N_15432,N_15084);
nor U15514 (N_15514,N_15292,N_15452);
or U15515 (N_15515,N_15118,N_15102);
nor U15516 (N_15516,N_15394,N_15416);
and U15517 (N_15517,N_15361,N_15440);
nand U15518 (N_15518,N_15191,N_15303);
xor U15519 (N_15519,N_15031,N_15008);
and U15520 (N_15520,N_15183,N_15203);
and U15521 (N_15521,N_15473,N_15308);
and U15522 (N_15522,N_15058,N_15134);
xnor U15523 (N_15523,N_15174,N_15264);
nor U15524 (N_15524,N_15341,N_15386);
or U15525 (N_15525,N_15240,N_15328);
nand U15526 (N_15526,N_15421,N_15148);
or U15527 (N_15527,N_15033,N_15229);
or U15528 (N_15528,N_15089,N_15285);
nand U15529 (N_15529,N_15375,N_15125);
and U15530 (N_15530,N_15252,N_15334);
nor U15531 (N_15531,N_15242,N_15490);
nor U15532 (N_15532,N_15076,N_15331);
or U15533 (N_15533,N_15412,N_15434);
nor U15534 (N_15534,N_15278,N_15407);
or U15535 (N_15535,N_15071,N_15402);
nor U15536 (N_15536,N_15069,N_15306);
or U15537 (N_15537,N_15222,N_15411);
and U15538 (N_15538,N_15271,N_15365);
and U15539 (N_15539,N_15097,N_15037);
xnor U15540 (N_15540,N_15018,N_15263);
nand U15541 (N_15541,N_15146,N_15488);
or U15542 (N_15542,N_15484,N_15214);
nor U15543 (N_15543,N_15498,N_15236);
or U15544 (N_15544,N_15325,N_15115);
nor U15545 (N_15545,N_15181,N_15180);
and U15546 (N_15546,N_15246,N_15200);
xor U15547 (N_15547,N_15281,N_15024);
or U15548 (N_15548,N_15251,N_15056);
xor U15549 (N_15549,N_15289,N_15270);
xor U15550 (N_15550,N_15036,N_15227);
nor U15551 (N_15551,N_15354,N_15238);
nor U15552 (N_15552,N_15483,N_15225);
nand U15553 (N_15553,N_15158,N_15448);
or U15554 (N_15554,N_15176,N_15192);
and U15555 (N_15555,N_15439,N_15109);
or U15556 (N_15556,N_15063,N_15294);
and U15557 (N_15557,N_15123,N_15279);
nor U15558 (N_15558,N_15224,N_15378);
nand U15559 (N_15559,N_15492,N_15074);
or U15560 (N_15560,N_15335,N_15197);
and U15561 (N_15561,N_15035,N_15136);
and U15562 (N_15562,N_15380,N_15346);
nor U15563 (N_15563,N_15232,N_15201);
nor U15564 (N_15564,N_15454,N_15314);
xor U15565 (N_15565,N_15326,N_15040);
xnor U15566 (N_15566,N_15305,N_15245);
and U15567 (N_15567,N_15291,N_15369);
or U15568 (N_15568,N_15268,N_15065);
nand U15569 (N_15569,N_15356,N_15430);
nand U15570 (N_15570,N_15272,N_15112);
and U15571 (N_15571,N_15169,N_15237);
nor U15572 (N_15572,N_15121,N_15179);
nand U15573 (N_15573,N_15493,N_15469);
nand U15574 (N_15574,N_15485,N_15382);
xor U15575 (N_15575,N_15182,N_15247);
xor U15576 (N_15576,N_15423,N_15137);
and U15577 (N_15577,N_15352,N_15442);
nor U15578 (N_15578,N_15302,N_15480);
or U15579 (N_15579,N_15093,N_15135);
xor U15580 (N_15580,N_15399,N_15154);
xnor U15581 (N_15581,N_15189,N_15164);
and U15582 (N_15582,N_15139,N_15280);
nor U15583 (N_15583,N_15397,N_15385);
and U15584 (N_15584,N_15188,N_15377);
and U15585 (N_15585,N_15171,N_15190);
nand U15586 (N_15586,N_15228,N_15419);
or U15587 (N_15587,N_15357,N_15470);
nand U15588 (N_15588,N_15427,N_15390);
xnor U15589 (N_15589,N_15286,N_15262);
and U15590 (N_15590,N_15384,N_15417);
xnor U15591 (N_15591,N_15482,N_15195);
nor U15592 (N_15592,N_15401,N_15087);
nor U15593 (N_15593,N_15081,N_15007);
xnor U15594 (N_15594,N_15259,N_15185);
or U15595 (N_15595,N_15358,N_15467);
nor U15596 (N_15596,N_15428,N_15460);
nor U15597 (N_15597,N_15248,N_15124);
and U15598 (N_15598,N_15218,N_15049);
and U15599 (N_15599,N_15300,N_15145);
or U15600 (N_15600,N_15457,N_15301);
nand U15601 (N_15601,N_15364,N_15458);
nor U15602 (N_15602,N_15426,N_15233);
and U15603 (N_15603,N_15316,N_15349);
and U15604 (N_15604,N_15355,N_15175);
xor U15605 (N_15605,N_15039,N_15451);
nor U15606 (N_15606,N_15277,N_15094);
and U15607 (N_15607,N_15073,N_15297);
xnor U15608 (N_15608,N_15389,N_15046);
or U15609 (N_15609,N_15312,N_15274);
nand U15610 (N_15610,N_15143,N_15099);
xor U15611 (N_15611,N_15051,N_15167);
and U15612 (N_15612,N_15163,N_15019);
or U15613 (N_15613,N_15126,N_15425);
nor U15614 (N_15614,N_15443,N_15045);
xor U15615 (N_15615,N_15186,N_15108);
nor U15616 (N_15616,N_15249,N_15383);
nor U15617 (N_15617,N_15015,N_15424);
xnor U15618 (N_15618,N_15138,N_15017);
and U15619 (N_15619,N_15350,N_15372);
nand U15620 (N_15620,N_15172,N_15059);
or U15621 (N_15621,N_15370,N_15116);
nand U15622 (N_15622,N_15293,N_15324);
nor U15623 (N_15623,N_15220,N_15464);
and U15624 (N_15624,N_15333,N_15343);
nand U15625 (N_15625,N_15034,N_15156);
and U15626 (N_15626,N_15133,N_15003);
or U15627 (N_15627,N_15408,N_15494);
and U15628 (N_15628,N_15206,N_15004);
nand U15629 (N_15629,N_15211,N_15320);
and U15630 (N_15630,N_15290,N_15438);
nand U15631 (N_15631,N_15436,N_15340);
nor U15632 (N_15632,N_15475,N_15344);
nor U15633 (N_15633,N_15155,N_15012);
nor U15634 (N_15634,N_15431,N_15110);
and U15635 (N_15635,N_15250,N_15422);
or U15636 (N_15636,N_15053,N_15239);
nor U15637 (N_15637,N_15132,N_15404);
nand U15638 (N_15638,N_15038,N_15379);
or U15639 (N_15639,N_15068,N_15491);
and U15640 (N_15640,N_15234,N_15338);
nor U15641 (N_15641,N_15282,N_15362);
nor U15642 (N_15642,N_15477,N_15128);
xor U15643 (N_15643,N_15456,N_15311);
or U15644 (N_15644,N_15323,N_15090);
nor U15645 (N_15645,N_15461,N_15168);
nand U15646 (N_15646,N_15437,N_15170);
or U15647 (N_15647,N_15360,N_15013);
nand U15648 (N_15648,N_15409,N_15029);
xnor U15649 (N_15649,N_15450,N_15481);
nor U15650 (N_15650,N_15449,N_15213);
nand U15651 (N_15651,N_15178,N_15459);
or U15652 (N_15652,N_15414,N_15104);
or U15653 (N_15653,N_15107,N_15050);
and U15654 (N_15654,N_15131,N_15283);
and U15655 (N_15655,N_15288,N_15208);
xor U15656 (N_15656,N_15088,N_15337);
xnor U15657 (N_15657,N_15273,N_15368);
nor U15658 (N_15658,N_15266,N_15149);
xor U15659 (N_15659,N_15339,N_15471);
or U15660 (N_15660,N_15079,N_15210);
and U15661 (N_15661,N_15387,N_15048);
xor U15662 (N_15662,N_15223,N_15359);
nor U15663 (N_15663,N_15243,N_15381);
nand U15664 (N_15664,N_15219,N_15057);
xnor U15665 (N_15665,N_15159,N_15441);
nand U15666 (N_15666,N_15275,N_15101);
and U15667 (N_15667,N_15287,N_15147);
nand U15668 (N_15668,N_15129,N_15474);
nor U15669 (N_15669,N_15212,N_15011);
nor U15670 (N_15670,N_15295,N_15028);
xor U15671 (N_15671,N_15130,N_15447);
or U15672 (N_15672,N_15465,N_15199);
and U15673 (N_15673,N_15400,N_15006);
nor U15674 (N_15674,N_15230,N_15119);
xor U15675 (N_15675,N_15085,N_15444);
and U15676 (N_15676,N_15307,N_15269);
xnor U15677 (N_15677,N_15496,N_15086);
nand U15678 (N_15678,N_15042,N_15153);
and U15679 (N_15679,N_15023,N_15032);
nand U15680 (N_15680,N_15244,N_15226);
and U15681 (N_15681,N_15462,N_15165);
nand U15682 (N_15682,N_15100,N_15141);
xor U15683 (N_15683,N_15255,N_15080);
xnor U15684 (N_15684,N_15009,N_15241);
nand U15685 (N_15685,N_15318,N_15096);
or U15686 (N_15686,N_15000,N_15055);
nand U15687 (N_15687,N_15070,N_15257);
or U15688 (N_15688,N_15160,N_15332);
nor U15689 (N_15689,N_15497,N_15091);
or U15690 (N_15690,N_15113,N_15415);
nor U15691 (N_15691,N_15140,N_15472);
xor U15692 (N_15692,N_15253,N_15342);
nand U15693 (N_15693,N_15265,N_15258);
and U15694 (N_15694,N_15478,N_15105);
xor U15695 (N_15695,N_15077,N_15161);
and U15696 (N_15696,N_15187,N_15173);
nand U15697 (N_15697,N_15044,N_15376);
or U15698 (N_15698,N_15276,N_15157);
nor U15699 (N_15699,N_15106,N_15398);
nand U15700 (N_15700,N_15202,N_15062);
or U15701 (N_15701,N_15005,N_15022);
nand U15702 (N_15702,N_15142,N_15061);
and U15703 (N_15703,N_15296,N_15321);
nand U15704 (N_15704,N_15209,N_15066);
and U15705 (N_15705,N_15047,N_15392);
and U15706 (N_15706,N_15001,N_15016);
nor U15707 (N_15707,N_15054,N_15489);
nor U15708 (N_15708,N_15103,N_15111);
nor U15709 (N_15709,N_15027,N_15078);
xnor U15710 (N_15710,N_15313,N_15393);
and U15711 (N_15711,N_15014,N_15327);
or U15712 (N_15712,N_15487,N_15002);
nand U15713 (N_15713,N_15373,N_15304);
or U15714 (N_15714,N_15479,N_15025);
or U15715 (N_15715,N_15310,N_15374);
nand U15716 (N_15716,N_15216,N_15486);
or U15717 (N_15717,N_15072,N_15184);
xor U15718 (N_15718,N_15353,N_15152);
nor U15719 (N_15719,N_15117,N_15410);
nor U15720 (N_15720,N_15468,N_15254);
xor U15721 (N_15721,N_15367,N_15260);
nor U15722 (N_15722,N_15466,N_15127);
or U15723 (N_15723,N_15231,N_15363);
nor U15724 (N_15724,N_15151,N_15043);
nor U15725 (N_15725,N_15261,N_15420);
nor U15726 (N_15726,N_15405,N_15177);
or U15727 (N_15727,N_15082,N_15413);
nand U15728 (N_15728,N_15453,N_15396);
xor U15729 (N_15729,N_15336,N_15330);
nand U15730 (N_15730,N_15391,N_15205);
or U15731 (N_15731,N_15446,N_15204);
nor U15732 (N_15732,N_15144,N_15092);
nand U15733 (N_15733,N_15315,N_15026);
and U15734 (N_15734,N_15403,N_15309);
or U15735 (N_15735,N_15021,N_15060);
nand U15736 (N_15736,N_15388,N_15041);
nand U15737 (N_15737,N_15196,N_15217);
nor U15738 (N_15738,N_15030,N_15395);
nor U15739 (N_15739,N_15347,N_15162);
and U15740 (N_15740,N_15166,N_15052);
xnor U15741 (N_15741,N_15267,N_15319);
or U15742 (N_15742,N_15215,N_15406);
nand U15743 (N_15743,N_15322,N_15075);
and U15744 (N_15744,N_15095,N_15345);
and U15745 (N_15745,N_15317,N_15020);
nand U15746 (N_15746,N_15499,N_15329);
xnor U15747 (N_15747,N_15445,N_15476);
xor U15748 (N_15748,N_15366,N_15429);
nor U15749 (N_15749,N_15098,N_15194);
nand U15750 (N_15750,N_15060,N_15455);
and U15751 (N_15751,N_15139,N_15430);
and U15752 (N_15752,N_15268,N_15105);
and U15753 (N_15753,N_15066,N_15071);
nand U15754 (N_15754,N_15461,N_15245);
xnor U15755 (N_15755,N_15233,N_15139);
nor U15756 (N_15756,N_15221,N_15381);
or U15757 (N_15757,N_15061,N_15015);
or U15758 (N_15758,N_15378,N_15300);
nand U15759 (N_15759,N_15232,N_15325);
nor U15760 (N_15760,N_15283,N_15380);
nor U15761 (N_15761,N_15168,N_15442);
xor U15762 (N_15762,N_15167,N_15043);
or U15763 (N_15763,N_15053,N_15134);
nand U15764 (N_15764,N_15052,N_15026);
xnor U15765 (N_15765,N_15341,N_15224);
and U15766 (N_15766,N_15150,N_15304);
nor U15767 (N_15767,N_15259,N_15455);
xnor U15768 (N_15768,N_15284,N_15394);
nor U15769 (N_15769,N_15362,N_15004);
nand U15770 (N_15770,N_15469,N_15082);
nor U15771 (N_15771,N_15258,N_15374);
xor U15772 (N_15772,N_15400,N_15143);
xnor U15773 (N_15773,N_15107,N_15317);
and U15774 (N_15774,N_15093,N_15103);
nor U15775 (N_15775,N_15404,N_15219);
nand U15776 (N_15776,N_15292,N_15164);
nor U15777 (N_15777,N_15343,N_15195);
and U15778 (N_15778,N_15428,N_15398);
nand U15779 (N_15779,N_15106,N_15418);
and U15780 (N_15780,N_15268,N_15312);
nand U15781 (N_15781,N_15082,N_15149);
xnor U15782 (N_15782,N_15016,N_15029);
xor U15783 (N_15783,N_15418,N_15388);
and U15784 (N_15784,N_15131,N_15323);
or U15785 (N_15785,N_15218,N_15166);
xnor U15786 (N_15786,N_15059,N_15408);
xor U15787 (N_15787,N_15450,N_15390);
xnor U15788 (N_15788,N_15192,N_15338);
nor U15789 (N_15789,N_15324,N_15411);
xnor U15790 (N_15790,N_15280,N_15174);
nor U15791 (N_15791,N_15346,N_15104);
and U15792 (N_15792,N_15146,N_15255);
xor U15793 (N_15793,N_15361,N_15272);
nand U15794 (N_15794,N_15441,N_15029);
xnor U15795 (N_15795,N_15023,N_15210);
nand U15796 (N_15796,N_15354,N_15424);
or U15797 (N_15797,N_15471,N_15076);
nor U15798 (N_15798,N_15110,N_15160);
nand U15799 (N_15799,N_15415,N_15370);
xor U15800 (N_15800,N_15294,N_15360);
and U15801 (N_15801,N_15486,N_15407);
nor U15802 (N_15802,N_15331,N_15470);
xor U15803 (N_15803,N_15228,N_15183);
nand U15804 (N_15804,N_15327,N_15323);
or U15805 (N_15805,N_15073,N_15377);
or U15806 (N_15806,N_15141,N_15020);
xnor U15807 (N_15807,N_15485,N_15489);
and U15808 (N_15808,N_15295,N_15240);
nor U15809 (N_15809,N_15226,N_15121);
and U15810 (N_15810,N_15243,N_15097);
xor U15811 (N_15811,N_15171,N_15325);
xnor U15812 (N_15812,N_15087,N_15460);
or U15813 (N_15813,N_15485,N_15263);
or U15814 (N_15814,N_15318,N_15061);
and U15815 (N_15815,N_15459,N_15274);
nand U15816 (N_15816,N_15188,N_15157);
xor U15817 (N_15817,N_15144,N_15395);
and U15818 (N_15818,N_15363,N_15177);
nor U15819 (N_15819,N_15387,N_15193);
or U15820 (N_15820,N_15378,N_15178);
nand U15821 (N_15821,N_15477,N_15120);
nand U15822 (N_15822,N_15373,N_15270);
and U15823 (N_15823,N_15056,N_15133);
and U15824 (N_15824,N_15240,N_15429);
xnor U15825 (N_15825,N_15045,N_15272);
xor U15826 (N_15826,N_15491,N_15128);
and U15827 (N_15827,N_15309,N_15360);
nand U15828 (N_15828,N_15211,N_15318);
and U15829 (N_15829,N_15026,N_15247);
nor U15830 (N_15830,N_15465,N_15421);
and U15831 (N_15831,N_15469,N_15369);
or U15832 (N_15832,N_15056,N_15332);
or U15833 (N_15833,N_15199,N_15247);
nand U15834 (N_15834,N_15304,N_15360);
nor U15835 (N_15835,N_15471,N_15095);
nand U15836 (N_15836,N_15290,N_15143);
or U15837 (N_15837,N_15056,N_15173);
and U15838 (N_15838,N_15075,N_15233);
xnor U15839 (N_15839,N_15112,N_15337);
nor U15840 (N_15840,N_15251,N_15032);
and U15841 (N_15841,N_15198,N_15237);
nand U15842 (N_15842,N_15380,N_15059);
nor U15843 (N_15843,N_15046,N_15243);
nand U15844 (N_15844,N_15254,N_15034);
nor U15845 (N_15845,N_15421,N_15011);
xnor U15846 (N_15846,N_15365,N_15182);
nand U15847 (N_15847,N_15219,N_15024);
nor U15848 (N_15848,N_15217,N_15153);
and U15849 (N_15849,N_15003,N_15138);
nand U15850 (N_15850,N_15109,N_15280);
or U15851 (N_15851,N_15158,N_15427);
nand U15852 (N_15852,N_15225,N_15005);
nand U15853 (N_15853,N_15194,N_15062);
nor U15854 (N_15854,N_15231,N_15335);
or U15855 (N_15855,N_15106,N_15448);
and U15856 (N_15856,N_15290,N_15217);
xor U15857 (N_15857,N_15253,N_15116);
nand U15858 (N_15858,N_15312,N_15497);
and U15859 (N_15859,N_15295,N_15400);
nand U15860 (N_15860,N_15003,N_15011);
nor U15861 (N_15861,N_15226,N_15416);
nor U15862 (N_15862,N_15267,N_15228);
and U15863 (N_15863,N_15257,N_15303);
nor U15864 (N_15864,N_15110,N_15452);
xnor U15865 (N_15865,N_15134,N_15014);
nor U15866 (N_15866,N_15427,N_15063);
and U15867 (N_15867,N_15227,N_15137);
nand U15868 (N_15868,N_15416,N_15108);
and U15869 (N_15869,N_15147,N_15490);
or U15870 (N_15870,N_15448,N_15401);
nor U15871 (N_15871,N_15278,N_15266);
or U15872 (N_15872,N_15066,N_15163);
and U15873 (N_15873,N_15409,N_15226);
xnor U15874 (N_15874,N_15032,N_15339);
or U15875 (N_15875,N_15260,N_15124);
xnor U15876 (N_15876,N_15407,N_15245);
xor U15877 (N_15877,N_15185,N_15178);
nand U15878 (N_15878,N_15218,N_15351);
or U15879 (N_15879,N_15175,N_15193);
xor U15880 (N_15880,N_15026,N_15212);
nand U15881 (N_15881,N_15371,N_15183);
or U15882 (N_15882,N_15240,N_15109);
xnor U15883 (N_15883,N_15307,N_15163);
nand U15884 (N_15884,N_15037,N_15301);
xor U15885 (N_15885,N_15057,N_15226);
and U15886 (N_15886,N_15460,N_15158);
or U15887 (N_15887,N_15488,N_15396);
and U15888 (N_15888,N_15051,N_15038);
nor U15889 (N_15889,N_15097,N_15425);
or U15890 (N_15890,N_15263,N_15193);
xor U15891 (N_15891,N_15049,N_15499);
nor U15892 (N_15892,N_15298,N_15389);
or U15893 (N_15893,N_15260,N_15170);
nor U15894 (N_15894,N_15012,N_15087);
xor U15895 (N_15895,N_15339,N_15016);
or U15896 (N_15896,N_15035,N_15330);
xor U15897 (N_15897,N_15132,N_15193);
or U15898 (N_15898,N_15169,N_15426);
xnor U15899 (N_15899,N_15298,N_15402);
or U15900 (N_15900,N_15474,N_15233);
nor U15901 (N_15901,N_15201,N_15342);
nand U15902 (N_15902,N_15234,N_15496);
nand U15903 (N_15903,N_15466,N_15378);
nand U15904 (N_15904,N_15198,N_15488);
xnor U15905 (N_15905,N_15341,N_15452);
nand U15906 (N_15906,N_15460,N_15122);
and U15907 (N_15907,N_15332,N_15275);
or U15908 (N_15908,N_15005,N_15034);
nand U15909 (N_15909,N_15064,N_15088);
or U15910 (N_15910,N_15164,N_15428);
nor U15911 (N_15911,N_15190,N_15455);
nand U15912 (N_15912,N_15344,N_15425);
nor U15913 (N_15913,N_15470,N_15309);
or U15914 (N_15914,N_15345,N_15209);
and U15915 (N_15915,N_15168,N_15444);
nand U15916 (N_15916,N_15113,N_15026);
nand U15917 (N_15917,N_15430,N_15148);
and U15918 (N_15918,N_15309,N_15450);
and U15919 (N_15919,N_15036,N_15098);
nor U15920 (N_15920,N_15434,N_15353);
and U15921 (N_15921,N_15313,N_15089);
and U15922 (N_15922,N_15115,N_15085);
or U15923 (N_15923,N_15244,N_15228);
nand U15924 (N_15924,N_15420,N_15054);
or U15925 (N_15925,N_15485,N_15414);
nor U15926 (N_15926,N_15371,N_15286);
nor U15927 (N_15927,N_15476,N_15064);
nor U15928 (N_15928,N_15001,N_15043);
and U15929 (N_15929,N_15414,N_15177);
or U15930 (N_15930,N_15490,N_15222);
xor U15931 (N_15931,N_15382,N_15057);
or U15932 (N_15932,N_15092,N_15277);
nand U15933 (N_15933,N_15014,N_15185);
or U15934 (N_15934,N_15398,N_15309);
nor U15935 (N_15935,N_15435,N_15335);
and U15936 (N_15936,N_15109,N_15231);
or U15937 (N_15937,N_15380,N_15444);
nand U15938 (N_15938,N_15450,N_15488);
nor U15939 (N_15939,N_15025,N_15136);
or U15940 (N_15940,N_15022,N_15118);
nand U15941 (N_15941,N_15122,N_15474);
xnor U15942 (N_15942,N_15204,N_15073);
nor U15943 (N_15943,N_15251,N_15222);
and U15944 (N_15944,N_15354,N_15097);
xnor U15945 (N_15945,N_15007,N_15311);
nor U15946 (N_15946,N_15314,N_15276);
nand U15947 (N_15947,N_15031,N_15225);
or U15948 (N_15948,N_15008,N_15252);
nand U15949 (N_15949,N_15062,N_15014);
xnor U15950 (N_15950,N_15493,N_15266);
xnor U15951 (N_15951,N_15265,N_15309);
nand U15952 (N_15952,N_15358,N_15468);
or U15953 (N_15953,N_15084,N_15031);
and U15954 (N_15954,N_15360,N_15242);
and U15955 (N_15955,N_15453,N_15128);
or U15956 (N_15956,N_15070,N_15355);
nor U15957 (N_15957,N_15248,N_15080);
and U15958 (N_15958,N_15076,N_15097);
nor U15959 (N_15959,N_15201,N_15025);
and U15960 (N_15960,N_15341,N_15052);
xnor U15961 (N_15961,N_15195,N_15381);
nand U15962 (N_15962,N_15354,N_15463);
nor U15963 (N_15963,N_15368,N_15025);
nor U15964 (N_15964,N_15090,N_15179);
xnor U15965 (N_15965,N_15146,N_15329);
xnor U15966 (N_15966,N_15495,N_15299);
nor U15967 (N_15967,N_15080,N_15346);
or U15968 (N_15968,N_15017,N_15364);
nand U15969 (N_15969,N_15286,N_15405);
nor U15970 (N_15970,N_15366,N_15229);
xor U15971 (N_15971,N_15354,N_15262);
or U15972 (N_15972,N_15331,N_15349);
and U15973 (N_15973,N_15240,N_15470);
nor U15974 (N_15974,N_15454,N_15316);
xnor U15975 (N_15975,N_15461,N_15449);
xnor U15976 (N_15976,N_15247,N_15054);
xnor U15977 (N_15977,N_15003,N_15453);
nor U15978 (N_15978,N_15062,N_15347);
and U15979 (N_15979,N_15097,N_15230);
xor U15980 (N_15980,N_15062,N_15017);
xnor U15981 (N_15981,N_15109,N_15328);
nand U15982 (N_15982,N_15096,N_15093);
nor U15983 (N_15983,N_15001,N_15473);
nor U15984 (N_15984,N_15086,N_15165);
xor U15985 (N_15985,N_15151,N_15078);
and U15986 (N_15986,N_15192,N_15296);
nor U15987 (N_15987,N_15120,N_15025);
and U15988 (N_15988,N_15227,N_15344);
and U15989 (N_15989,N_15351,N_15490);
and U15990 (N_15990,N_15281,N_15020);
xnor U15991 (N_15991,N_15245,N_15292);
and U15992 (N_15992,N_15443,N_15363);
and U15993 (N_15993,N_15323,N_15281);
and U15994 (N_15994,N_15301,N_15466);
and U15995 (N_15995,N_15375,N_15470);
nor U15996 (N_15996,N_15250,N_15235);
nand U15997 (N_15997,N_15139,N_15100);
nor U15998 (N_15998,N_15085,N_15015);
and U15999 (N_15999,N_15195,N_15213);
nor U16000 (N_16000,N_15767,N_15559);
nand U16001 (N_16001,N_15697,N_15549);
and U16002 (N_16002,N_15797,N_15635);
or U16003 (N_16003,N_15796,N_15793);
or U16004 (N_16004,N_15546,N_15870);
xnor U16005 (N_16005,N_15712,N_15867);
or U16006 (N_16006,N_15953,N_15917);
xor U16007 (N_16007,N_15863,N_15667);
xor U16008 (N_16008,N_15560,N_15788);
and U16009 (N_16009,N_15829,N_15900);
xnor U16010 (N_16010,N_15789,N_15852);
nand U16011 (N_16011,N_15865,N_15899);
nor U16012 (N_16012,N_15534,N_15731);
and U16013 (N_16013,N_15531,N_15755);
or U16014 (N_16014,N_15980,N_15759);
nand U16015 (N_16015,N_15520,N_15934);
and U16016 (N_16016,N_15817,N_15701);
nand U16017 (N_16017,N_15624,N_15949);
nor U16018 (N_16018,N_15637,N_15842);
and U16019 (N_16019,N_15683,N_15725);
and U16020 (N_16020,N_15555,N_15685);
nand U16021 (N_16021,N_15969,N_15943);
nand U16022 (N_16022,N_15566,N_15897);
nand U16023 (N_16023,N_15726,N_15678);
nand U16024 (N_16024,N_15567,N_15875);
nor U16025 (N_16025,N_15909,N_15910);
nand U16026 (N_16026,N_15643,N_15680);
or U16027 (N_16027,N_15630,N_15884);
or U16028 (N_16028,N_15634,N_15664);
nand U16029 (N_16029,N_15979,N_15923);
or U16030 (N_16030,N_15981,N_15577);
and U16031 (N_16031,N_15606,N_15602);
or U16032 (N_16032,N_15978,N_15754);
xnor U16033 (N_16033,N_15690,N_15764);
nor U16034 (N_16034,N_15654,N_15992);
xor U16035 (N_16035,N_15727,N_15787);
or U16036 (N_16036,N_15735,N_15500);
and U16037 (N_16037,N_15578,N_15580);
and U16038 (N_16038,N_15887,N_15948);
and U16039 (N_16039,N_15583,N_15785);
xnor U16040 (N_16040,N_15803,N_15786);
or U16041 (N_16041,N_15752,N_15618);
nand U16042 (N_16042,N_15914,N_15839);
nor U16043 (N_16043,N_15509,N_15891);
and U16044 (N_16044,N_15812,N_15896);
and U16045 (N_16045,N_15514,N_15898);
or U16046 (N_16046,N_15539,N_15811);
nor U16047 (N_16047,N_15561,N_15874);
or U16048 (N_16048,N_15950,N_15719);
or U16049 (N_16049,N_15807,N_15882);
xnor U16050 (N_16050,N_15951,N_15822);
xor U16051 (N_16051,N_15682,N_15614);
nand U16052 (N_16052,N_15536,N_15699);
nor U16053 (N_16053,N_15600,N_15704);
and U16054 (N_16054,N_15595,N_15573);
or U16055 (N_16055,N_15584,N_15652);
or U16056 (N_16056,N_15629,N_15835);
or U16057 (N_16057,N_15821,N_15706);
nand U16058 (N_16058,N_15657,N_15982);
and U16059 (N_16059,N_15927,N_15962);
nand U16060 (N_16060,N_15763,N_15651);
or U16061 (N_16061,N_15713,N_15504);
nor U16062 (N_16062,N_15838,N_15579);
or U16063 (N_16063,N_15593,N_15881);
and U16064 (N_16064,N_15804,N_15502);
nand U16065 (N_16065,N_15644,N_15505);
xor U16066 (N_16066,N_15547,N_15963);
nand U16067 (N_16067,N_15708,N_15562);
or U16068 (N_16068,N_15771,N_15700);
nand U16069 (N_16069,N_15773,N_15922);
nor U16070 (N_16070,N_15711,N_15626);
and U16071 (N_16071,N_15907,N_15931);
or U16072 (N_16072,N_15503,N_15601);
or U16073 (N_16073,N_15935,N_15599);
xnor U16074 (N_16074,N_15762,N_15660);
nand U16075 (N_16075,N_15622,N_15843);
xnor U16076 (N_16076,N_15993,N_15864);
or U16077 (N_16077,N_15598,N_15707);
nand U16078 (N_16078,N_15823,N_15830);
nand U16079 (N_16079,N_15656,N_15510);
or U16080 (N_16080,N_15723,N_15929);
and U16081 (N_16081,N_15799,N_15750);
nor U16082 (N_16082,N_15686,N_15553);
and U16083 (N_16083,N_15627,N_15798);
xor U16084 (N_16084,N_15977,N_15638);
and U16085 (N_16085,N_15776,N_15973);
and U16086 (N_16086,N_15543,N_15591);
xor U16087 (N_16087,N_15937,N_15659);
and U16088 (N_16088,N_15537,N_15738);
nor U16089 (N_16089,N_15563,N_15904);
or U16090 (N_16090,N_15508,N_15649);
nor U16091 (N_16091,N_15702,N_15903);
and U16092 (N_16092,N_15524,N_15818);
xnor U16093 (N_16093,N_15715,N_15901);
xnor U16094 (N_16094,N_15691,N_15942);
nand U16095 (N_16095,N_15826,N_15589);
nand U16096 (N_16096,N_15941,N_15768);
nand U16097 (N_16097,N_15888,N_15571);
and U16098 (N_16098,N_15609,N_15769);
xor U16099 (N_16099,N_15815,N_15631);
xor U16100 (N_16100,N_15710,N_15885);
xor U16101 (N_16101,N_15564,N_15880);
or U16102 (N_16102,N_15603,N_15517);
or U16103 (N_16103,N_15961,N_15889);
nand U16104 (N_16104,N_15512,N_15971);
nand U16105 (N_16105,N_15997,N_15800);
and U16106 (N_16106,N_15548,N_15860);
or U16107 (N_16107,N_15717,N_15501);
or U16108 (N_16108,N_15625,N_15744);
or U16109 (N_16109,N_15959,N_15586);
or U16110 (N_16110,N_15938,N_15545);
and U16111 (N_16111,N_15783,N_15827);
and U16112 (N_16112,N_15613,N_15871);
nor U16113 (N_16113,N_15930,N_15868);
nand U16114 (N_16114,N_15572,N_15607);
xnor U16115 (N_16115,N_15779,N_15684);
nor U16116 (N_16116,N_15666,N_15845);
and U16117 (N_16117,N_15639,N_15676);
and U16118 (N_16118,N_15729,N_15756);
and U16119 (N_16119,N_15877,N_15530);
nor U16120 (N_16120,N_15990,N_15968);
nor U16121 (N_16121,N_15615,N_15551);
nand U16122 (N_16122,N_15521,N_15540);
or U16123 (N_16123,N_15648,N_15912);
xor U16124 (N_16124,N_15742,N_15714);
nor U16125 (N_16125,N_15612,N_15801);
and U16126 (N_16126,N_15958,N_15989);
nor U16127 (N_16127,N_15529,N_15940);
or U16128 (N_16128,N_15920,N_15525);
and U16129 (N_16129,N_15831,N_15532);
nand U16130 (N_16130,N_15728,N_15585);
and U16131 (N_16131,N_15890,N_15999);
or U16132 (N_16132,N_15740,N_15633);
or U16133 (N_16133,N_15858,N_15819);
or U16134 (N_16134,N_15926,N_15777);
and U16135 (N_16135,N_15693,N_15895);
nor U16136 (N_16136,N_15956,N_15516);
xor U16137 (N_16137,N_15970,N_15522);
nand U16138 (N_16138,N_15965,N_15720);
nor U16139 (N_16139,N_15513,N_15939);
or U16140 (N_16140,N_15533,N_15879);
nand U16141 (N_16141,N_15734,N_15669);
or U16142 (N_16142,N_15733,N_15840);
nor U16143 (N_16143,N_15741,N_15778);
nor U16144 (N_16144,N_15991,N_15743);
nand U16145 (N_16145,N_15645,N_15919);
xor U16146 (N_16146,N_15640,N_15967);
nand U16147 (N_16147,N_15974,N_15966);
nor U16148 (N_16148,N_15668,N_15574);
nand U16149 (N_16149,N_15689,N_15642);
nor U16150 (N_16150,N_15590,N_15558);
nor U16151 (N_16151,N_15780,N_15761);
and U16152 (N_16152,N_15611,N_15745);
xnor U16153 (N_16153,N_15957,N_15915);
or U16154 (N_16154,N_15790,N_15805);
xnor U16155 (N_16155,N_15753,N_15565);
or U16156 (N_16156,N_15834,N_15619);
or U16157 (N_16157,N_15985,N_15809);
nor U16158 (N_16158,N_15673,N_15954);
nand U16159 (N_16159,N_15983,N_15996);
or U16160 (N_16160,N_15594,N_15677);
xor U16161 (N_16161,N_15632,N_15932);
or U16162 (N_16162,N_15984,N_15636);
nor U16163 (N_16163,N_15749,N_15810);
nor U16164 (N_16164,N_15802,N_15808);
or U16165 (N_16165,N_15556,N_15646);
or U16166 (N_16166,N_15587,N_15975);
nand U16167 (N_16167,N_15760,N_15674);
xnor U16168 (N_16168,N_15916,N_15894);
xnor U16169 (N_16169,N_15908,N_15675);
or U16170 (N_16170,N_15732,N_15861);
xor U16171 (N_16171,N_15698,N_15765);
and U16172 (N_16172,N_15592,N_15883);
nor U16173 (N_16173,N_15964,N_15672);
nor U16174 (N_16174,N_15866,N_15972);
xor U16175 (N_16175,N_15862,N_15557);
xor U16176 (N_16176,N_15925,N_15730);
nor U16177 (N_16177,N_15621,N_15737);
nand U16178 (N_16178,N_15581,N_15703);
nand U16179 (N_16179,N_15628,N_15550);
xnor U16180 (N_16180,N_15570,N_15976);
nand U16181 (N_16181,N_15608,N_15945);
and U16182 (N_16182,N_15813,N_15687);
and U16183 (N_16183,N_15705,N_15960);
or U16184 (N_16184,N_15846,N_15825);
and U16185 (N_16185,N_15575,N_15832);
nand U16186 (N_16186,N_15854,N_15662);
nand U16187 (N_16187,N_15671,N_15952);
and U16188 (N_16188,N_15588,N_15528);
or U16189 (N_16189,N_15766,N_15526);
xor U16190 (N_16190,N_15853,N_15775);
xor U16191 (N_16191,N_15869,N_15650);
xnor U16192 (N_16192,N_15616,N_15928);
xor U16193 (N_16193,N_15507,N_15892);
or U16194 (N_16194,N_15987,N_15658);
nor U16195 (N_16195,N_15653,N_15568);
xnor U16196 (N_16196,N_15806,N_15781);
or U16197 (N_16197,N_15506,N_15721);
nor U16198 (N_16198,N_15936,N_15511);
nor U16199 (N_16199,N_15855,N_15918);
nand U16200 (N_16200,N_15541,N_15688);
nand U16201 (N_16201,N_15610,N_15770);
nor U16202 (N_16202,N_15569,N_15748);
nor U16203 (N_16203,N_15774,N_15924);
and U16204 (N_16204,N_15523,N_15515);
nand U16205 (N_16205,N_15527,N_15946);
or U16206 (N_16206,N_15828,N_15623);
xor U16207 (N_16207,N_15955,N_15998);
and U16208 (N_16208,N_15859,N_15542);
and U16209 (N_16209,N_15739,N_15850);
or U16210 (N_16210,N_15836,N_15772);
xnor U16211 (N_16211,N_15988,N_15906);
nor U16212 (N_16212,N_15670,N_15824);
xnor U16213 (N_16213,N_15718,N_15538);
xnor U16214 (N_16214,N_15794,N_15597);
nor U16215 (N_16215,N_15605,N_15554);
nor U16216 (N_16216,N_15679,N_15784);
xor U16217 (N_16217,N_15814,N_15747);
nor U16218 (N_16218,N_15886,N_15893);
or U16219 (N_16219,N_15944,N_15736);
and U16220 (N_16220,N_15617,N_15655);
and U16221 (N_16221,N_15872,N_15841);
xnor U16222 (N_16222,N_15694,N_15552);
or U16223 (N_16223,N_15795,N_15816);
nand U16224 (N_16224,N_15851,N_15751);
nand U16225 (N_16225,N_15758,N_15724);
or U16226 (N_16226,N_15878,N_15921);
or U16227 (N_16227,N_15692,N_15856);
nor U16228 (N_16228,N_15722,N_15620);
nand U16229 (N_16229,N_15604,N_15518);
nor U16230 (N_16230,N_15994,N_15596);
nor U16231 (N_16231,N_15986,N_15844);
and U16232 (N_16232,N_15576,N_15820);
and U16233 (N_16233,N_15791,N_15933);
and U16234 (N_16234,N_15913,N_15848);
and U16235 (N_16235,N_15695,N_15995);
or U16236 (N_16236,N_15905,N_15947);
and U16237 (N_16237,N_15681,N_15911);
or U16238 (N_16238,N_15716,N_15876);
and U16239 (N_16239,N_15661,N_15544);
nor U16240 (N_16240,N_15873,N_15647);
nand U16241 (N_16241,N_15746,N_15641);
and U16242 (N_16242,N_15833,N_15857);
or U16243 (N_16243,N_15849,N_15902);
and U16244 (N_16244,N_15582,N_15519);
nor U16245 (N_16245,N_15535,N_15847);
or U16246 (N_16246,N_15709,N_15757);
nor U16247 (N_16247,N_15696,N_15665);
nand U16248 (N_16248,N_15782,N_15837);
nor U16249 (N_16249,N_15663,N_15792);
nand U16250 (N_16250,N_15516,N_15645);
and U16251 (N_16251,N_15505,N_15645);
and U16252 (N_16252,N_15958,N_15612);
xor U16253 (N_16253,N_15910,N_15555);
xnor U16254 (N_16254,N_15724,N_15590);
nand U16255 (N_16255,N_15947,N_15704);
xor U16256 (N_16256,N_15873,N_15845);
xor U16257 (N_16257,N_15530,N_15562);
xor U16258 (N_16258,N_15704,N_15879);
nand U16259 (N_16259,N_15859,N_15738);
xnor U16260 (N_16260,N_15524,N_15768);
or U16261 (N_16261,N_15871,N_15783);
and U16262 (N_16262,N_15622,N_15526);
and U16263 (N_16263,N_15686,N_15569);
xnor U16264 (N_16264,N_15839,N_15881);
nand U16265 (N_16265,N_15754,N_15663);
nand U16266 (N_16266,N_15704,N_15597);
nand U16267 (N_16267,N_15959,N_15811);
or U16268 (N_16268,N_15826,N_15984);
and U16269 (N_16269,N_15934,N_15874);
or U16270 (N_16270,N_15934,N_15748);
nand U16271 (N_16271,N_15520,N_15623);
and U16272 (N_16272,N_15832,N_15769);
and U16273 (N_16273,N_15947,N_15537);
or U16274 (N_16274,N_15575,N_15586);
nand U16275 (N_16275,N_15511,N_15759);
and U16276 (N_16276,N_15888,N_15992);
or U16277 (N_16277,N_15880,N_15842);
or U16278 (N_16278,N_15539,N_15566);
nor U16279 (N_16279,N_15566,N_15786);
nand U16280 (N_16280,N_15949,N_15607);
nand U16281 (N_16281,N_15931,N_15791);
or U16282 (N_16282,N_15677,N_15997);
xnor U16283 (N_16283,N_15700,N_15991);
nand U16284 (N_16284,N_15615,N_15709);
or U16285 (N_16285,N_15742,N_15536);
nor U16286 (N_16286,N_15837,N_15776);
xor U16287 (N_16287,N_15566,N_15698);
nor U16288 (N_16288,N_15651,N_15882);
xor U16289 (N_16289,N_15657,N_15738);
nand U16290 (N_16290,N_15531,N_15919);
nor U16291 (N_16291,N_15682,N_15822);
and U16292 (N_16292,N_15833,N_15787);
or U16293 (N_16293,N_15828,N_15619);
nand U16294 (N_16294,N_15503,N_15578);
and U16295 (N_16295,N_15580,N_15717);
xnor U16296 (N_16296,N_15778,N_15791);
and U16297 (N_16297,N_15557,N_15967);
nand U16298 (N_16298,N_15820,N_15732);
xnor U16299 (N_16299,N_15924,N_15772);
nor U16300 (N_16300,N_15551,N_15824);
nand U16301 (N_16301,N_15842,N_15536);
or U16302 (N_16302,N_15780,N_15611);
or U16303 (N_16303,N_15784,N_15937);
xnor U16304 (N_16304,N_15648,N_15942);
nand U16305 (N_16305,N_15509,N_15964);
nand U16306 (N_16306,N_15687,N_15501);
nor U16307 (N_16307,N_15671,N_15555);
and U16308 (N_16308,N_15954,N_15519);
nor U16309 (N_16309,N_15734,N_15772);
xnor U16310 (N_16310,N_15527,N_15788);
nand U16311 (N_16311,N_15834,N_15815);
nor U16312 (N_16312,N_15555,N_15646);
nor U16313 (N_16313,N_15524,N_15570);
xnor U16314 (N_16314,N_15809,N_15779);
and U16315 (N_16315,N_15898,N_15761);
or U16316 (N_16316,N_15572,N_15863);
nand U16317 (N_16317,N_15903,N_15916);
and U16318 (N_16318,N_15935,N_15849);
or U16319 (N_16319,N_15749,N_15864);
xor U16320 (N_16320,N_15503,N_15689);
nor U16321 (N_16321,N_15935,N_15604);
or U16322 (N_16322,N_15735,N_15942);
and U16323 (N_16323,N_15919,N_15848);
nand U16324 (N_16324,N_15704,N_15965);
nor U16325 (N_16325,N_15607,N_15627);
and U16326 (N_16326,N_15921,N_15692);
and U16327 (N_16327,N_15819,N_15992);
nand U16328 (N_16328,N_15705,N_15663);
or U16329 (N_16329,N_15757,N_15863);
nor U16330 (N_16330,N_15757,N_15539);
xnor U16331 (N_16331,N_15806,N_15870);
nor U16332 (N_16332,N_15637,N_15568);
xor U16333 (N_16333,N_15803,N_15714);
nor U16334 (N_16334,N_15801,N_15946);
xor U16335 (N_16335,N_15823,N_15680);
or U16336 (N_16336,N_15884,N_15511);
nand U16337 (N_16337,N_15782,N_15952);
nand U16338 (N_16338,N_15720,N_15897);
nand U16339 (N_16339,N_15748,N_15549);
nand U16340 (N_16340,N_15919,N_15561);
nand U16341 (N_16341,N_15915,N_15805);
and U16342 (N_16342,N_15739,N_15918);
or U16343 (N_16343,N_15735,N_15608);
nand U16344 (N_16344,N_15776,N_15939);
nand U16345 (N_16345,N_15523,N_15647);
and U16346 (N_16346,N_15618,N_15946);
nor U16347 (N_16347,N_15639,N_15625);
and U16348 (N_16348,N_15650,N_15896);
xnor U16349 (N_16349,N_15793,N_15654);
or U16350 (N_16350,N_15654,N_15911);
and U16351 (N_16351,N_15576,N_15734);
or U16352 (N_16352,N_15663,N_15601);
nand U16353 (N_16353,N_15710,N_15893);
nor U16354 (N_16354,N_15885,N_15629);
or U16355 (N_16355,N_15652,N_15643);
and U16356 (N_16356,N_15711,N_15982);
nand U16357 (N_16357,N_15609,N_15838);
and U16358 (N_16358,N_15844,N_15696);
xnor U16359 (N_16359,N_15522,N_15503);
nor U16360 (N_16360,N_15851,N_15973);
or U16361 (N_16361,N_15878,N_15939);
and U16362 (N_16362,N_15599,N_15616);
or U16363 (N_16363,N_15654,N_15789);
or U16364 (N_16364,N_15837,N_15685);
nor U16365 (N_16365,N_15874,N_15808);
and U16366 (N_16366,N_15546,N_15811);
xnor U16367 (N_16367,N_15999,N_15764);
nor U16368 (N_16368,N_15837,N_15638);
nor U16369 (N_16369,N_15715,N_15553);
and U16370 (N_16370,N_15962,N_15831);
xnor U16371 (N_16371,N_15775,N_15646);
nor U16372 (N_16372,N_15925,N_15881);
or U16373 (N_16373,N_15916,N_15755);
or U16374 (N_16374,N_15630,N_15646);
xnor U16375 (N_16375,N_15870,N_15820);
xnor U16376 (N_16376,N_15945,N_15780);
and U16377 (N_16377,N_15720,N_15550);
xor U16378 (N_16378,N_15645,N_15989);
xnor U16379 (N_16379,N_15560,N_15935);
or U16380 (N_16380,N_15508,N_15651);
nor U16381 (N_16381,N_15934,N_15974);
and U16382 (N_16382,N_15606,N_15932);
nand U16383 (N_16383,N_15956,N_15635);
or U16384 (N_16384,N_15781,N_15593);
and U16385 (N_16385,N_15553,N_15687);
nand U16386 (N_16386,N_15856,N_15589);
xnor U16387 (N_16387,N_15816,N_15764);
or U16388 (N_16388,N_15630,N_15716);
and U16389 (N_16389,N_15928,N_15611);
or U16390 (N_16390,N_15814,N_15535);
and U16391 (N_16391,N_15703,N_15719);
and U16392 (N_16392,N_15617,N_15804);
nand U16393 (N_16393,N_15935,N_15728);
or U16394 (N_16394,N_15971,N_15804);
nor U16395 (N_16395,N_15984,N_15749);
and U16396 (N_16396,N_15713,N_15746);
or U16397 (N_16397,N_15891,N_15860);
nor U16398 (N_16398,N_15775,N_15694);
nand U16399 (N_16399,N_15832,N_15595);
nand U16400 (N_16400,N_15719,N_15798);
nand U16401 (N_16401,N_15636,N_15665);
xnor U16402 (N_16402,N_15841,N_15720);
nand U16403 (N_16403,N_15975,N_15577);
nor U16404 (N_16404,N_15586,N_15625);
or U16405 (N_16405,N_15679,N_15528);
or U16406 (N_16406,N_15790,N_15964);
or U16407 (N_16407,N_15684,N_15850);
or U16408 (N_16408,N_15882,N_15635);
nand U16409 (N_16409,N_15853,N_15661);
and U16410 (N_16410,N_15505,N_15782);
or U16411 (N_16411,N_15656,N_15604);
nand U16412 (N_16412,N_15927,N_15817);
nand U16413 (N_16413,N_15807,N_15852);
nand U16414 (N_16414,N_15766,N_15551);
nand U16415 (N_16415,N_15971,N_15536);
xnor U16416 (N_16416,N_15959,N_15687);
xnor U16417 (N_16417,N_15823,N_15886);
nor U16418 (N_16418,N_15972,N_15909);
or U16419 (N_16419,N_15944,N_15641);
and U16420 (N_16420,N_15956,N_15824);
or U16421 (N_16421,N_15547,N_15942);
xor U16422 (N_16422,N_15753,N_15773);
nand U16423 (N_16423,N_15826,N_15510);
nor U16424 (N_16424,N_15860,N_15877);
and U16425 (N_16425,N_15845,N_15650);
nor U16426 (N_16426,N_15934,N_15702);
nand U16427 (N_16427,N_15821,N_15652);
nand U16428 (N_16428,N_15585,N_15853);
nand U16429 (N_16429,N_15977,N_15996);
xor U16430 (N_16430,N_15626,N_15712);
nor U16431 (N_16431,N_15749,N_15585);
xor U16432 (N_16432,N_15970,N_15580);
or U16433 (N_16433,N_15661,N_15760);
or U16434 (N_16434,N_15574,N_15501);
nand U16435 (N_16435,N_15943,N_15653);
nand U16436 (N_16436,N_15895,N_15890);
nor U16437 (N_16437,N_15840,N_15716);
nor U16438 (N_16438,N_15660,N_15836);
nor U16439 (N_16439,N_15587,N_15847);
or U16440 (N_16440,N_15993,N_15969);
or U16441 (N_16441,N_15752,N_15651);
or U16442 (N_16442,N_15630,N_15765);
and U16443 (N_16443,N_15819,N_15738);
and U16444 (N_16444,N_15920,N_15638);
nor U16445 (N_16445,N_15538,N_15836);
xnor U16446 (N_16446,N_15754,N_15588);
nand U16447 (N_16447,N_15957,N_15992);
xnor U16448 (N_16448,N_15560,N_15565);
xor U16449 (N_16449,N_15746,N_15984);
nand U16450 (N_16450,N_15526,N_15643);
or U16451 (N_16451,N_15777,N_15932);
nor U16452 (N_16452,N_15550,N_15574);
nor U16453 (N_16453,N_15614,N_15687);
nand U16454 (N_16454,N_15767,N_15519);
nand U16455 (N_16455,N_15560,N_15763);
and U16456 (N_16456,N_15940,N_15911);
nand U16457 (N_16457,N_15749,N_15887);
or U16458 (N_16458,N_15688,N_15748);
nand U16459 (N_16459,N_15954,N_15600);
xnor U16460 (N_16460,N_15832,N_15638);
nor U16461 (N_16461,N_15999,N_15705);
nand U16462 (N_16462,N_15852,N_15871);
nor U16463 (N_16463,N_15598,N_15640);
nor U16464 (N_16464,N_15920,N_15886);
or U16465 (N_16465,N_15774,N_15917);
nand U16466 (N_16466,N_15629,N_15740);
xor U16467 (N_16467,N_15534,N_15512);
nand U16468 (N_16468,N_15636,N_15842);
nand U16469 (N_16469,N_15575,N_15648);
xnor U16470 (N_16470,N_15521,N_15956);
and U16471 (N_16471,N_15935,N_15899);
nor U16472 (N_16472,N_15525,N_15658);
and U16473 (N_16473,N_15670,N_15676);
nand U16474 (N_16474,N_15876,N_15632);
or U16475 (N_16475,N_15664,N_15577);
xnor U16476 (N_16476,N_15502,N_15795);
nor U16477 (N_16477,N_15871,N_15959);
xor U16478 (N_16478,N_15751,N_15757);
nor U16479 (N_16479,N_15982,N_15766);
or U16480 (N_16480,N_15659,N_15800);
and U16481 (N_16481,N_15803,N_15690);
xnor U16482 (N_16482,N_15981,N_15623);
xor U16483 (N_16483,N_15915,N_15563);
and U16484 (N_16484,N_15779,N_15752);
xnor U16485 (N_16485,N_15519,N_15621);
nor U16486 (N_16486,N_15722,N_15962);
xor U16487 (N_16487,N_15556,N_15914);
nor U16488 (N_16488,N_15878,N_15877);
nand U16489 (N_16489,N_15730,N_15773);
or U16490 (N_16490,N_15850,N_15854);
or U16491 (N_16491,N_15946,N_15624);
or U16492 (N_16492,N_15505,N_15620);
or U16493 (N_16493,N_15577,N_15570);
nand U16494 (N_16494,N_15803,N_15596);
nor U16495 (N_16495,N_15771,N_15948);
or U16496 (N_16496,N_15992,N_15980);
nand U16497 (N_16497,N_15653,N_15888);
and U16498 (N_16498,N_15825,N_15939);
or U16499 (N_16499,N_15694,N_15982);
xnor U16500 (N_16500,N_16389,N_16430);
xnor U16501 (N_16501,N_16441,N_16210);
xor U16502 (N_16502,N_16369,N_16480);
nand U16503 (N_16503,N_16300,N_16481);
nor U16504 (N_16504,N_16173,N_16415);
or U16505 (N_16505,N_16404,N_16340);
nor U16506 (N_16506,N_16221,N_16489);
nor U16507 (N_16507,N_16485,N_16090);
or U16508 (N_16508,N_16324,N_16263);
xnor U16509 (N_16509,N_16107,N_16474);
xor U16510 (N_16510,N_16412,N_16342);
xor U16511 (N_16511,N_16432,N_16003);
nor U16512 (N_16512,N_16343,N_16346);
or U16513 (N_16513,N_16436,N_16361);
xnor U16514 (N_16514,N_16152,N_16017);
and U16515 (N_16515,N_16319,N_16241);
xnor U16516 (N_16516,N_16349,N_16227);
xor U16517 (N_16517,N_16116,N_16309);
xor U16518 (N_16518,N_16449,N_16467);
nor U16519 (N_16519,N_16077,N_16357);
nor U16520 (N_16520,N_16479,N_16167);
nand U16521 (N_16521,N_16125,N_16022);
nor U16522 (N_16522,N_16081,N_16180);
xnor U16523 (N_16523,N_16089,N_16420);
nor U16524 (N_16524,N_16040,N_16136);
xnor U16525 (N_16525,N_16265,N_16229);
nor U16526 (N_16526,N_16371,N_16155);
and U16527 (N_16527,N_16145,N_16146);
or U16528 (N_16528,N_16179,N_16454);
nand U16529 (N_16529,N_16071,N_16395);
nand U16530 (N_16530,N_16416,N_16028);
or U16531 (N_16531,N_16405,N_16445);
or U16532 (N_16532,N_16228,N_16399);
xnor U16533 (N_16533,N_16050,N_16095);
nand U16534 (N_16534,N_16446,N_16096);
nor U16535 (N_16535,N_16392,N_16382);
or U16536 (N_16536,N_16491,N_16115);
nand U16537 (N_16537,N_16242,N_16197);
xnor U16538 (N_16538,N_16352,N_16220);
nor U16539 (N_16539,N_16165,N_16086);
nor U16540 (N_16540,N_16147,N_16315);
xnor U16541 (N_16541,N_16196,N_16048);
nand U16542 (N_16542,N_16259,N_16010);
nor U16543 (N_16543,N_16118,N_16287);
nand U16544 (N_16544,N_16200,N_16294);
xor U16545 (N_16545,N_16053,N_16251);
nand U16546 (N_16546,N_16187,N_16381);
nor U16547 (N_16547,N_16433,N_16260);
nor U16548 (N_16548,N_16137,N_16288);
nor U16549 (N_16549,N_16439,N_16326);
nand U16550 (N_16550,N_16380,N_16109);
nor U16551 (N_16551,N_16103,N_16411);
and U16552 (N_16552,N_16066,N_16317);
nor U16553 (N_16553,N_16043,N_16143);
xnor U16554 (N_16554,N_16331,N_16170);
or U16555 (N_16555,N_16398,N_16466);
or U16556 (N_16556,N_16005,N_16183);
nor U16557 (N_16557,N_16188,N_16281);
or U16558 (N_16558,N_16226,N_16217);
nand U16559 (N_16559,N_16201,N_16079);
xor U16560 (N_16560,N_16144,N_16225);
nand U16561 (N_16561,N_16280,N_16164);
or U16562 (N_16562,N_16174,N_16422);
nor U16563 (N_16563,N_16247,N_16435);
nand U16564 (N_16564,N_16482,N_16025);
nor U16565 (N_16565,N_16007,N_16269);
xor U16566 (N_16566,N_16330,N_16451);
nor U16567 (N_16567,N_16410,N_16341);
nor U16568 (N_16568,N_16087,N_16402);
xor U16569 (N_16569,N_16127,N_16224);
xor U16570 (N_16570,N_16396,N_16014);
or U16571 (N_16571,N_16388,N_16397);
nor U16572 (N_16572,N_16458,N_16236);
and U16573 (N_16573,N_16356,N_16496);
nor U16574 (N_16574,N_16246,N_16299);
or U16575 (N_16575,N_16046,N_16002);
and U16576 (N_16576,N_16336,N_16009);
nor U16577 (N_16577,N_16133,N_16069);
xor U16578 (N_16578,N_16243,N_16169);
and U16579 (N_16579,N_16273,N_16293);
nand U16580 (N_16580,N_16407,N_16215);
or U16581 (N_16581,N_16178,N_16334);
xor U16582 (N_16582,N_16000,N_16438);
nor U16583 (N_16583,N_16120,N_16083);
xnor U16584 (N_16584,N_16368,N_16148);
and U16585 (N_16585,N_16181,N_16099);
or U16586 (N_16586,N_16364,N_16151);
and U16587 (N_16587,N_16131,N_16117);
or U16588 (N_16588,N_16354,N_16321);
xnor U16589 (N_16589,N_16031,N_16168);
nand U16590 (N_16590,N_16427,N_16456);
nand U16591 (N_16591,N_16237,N_16037);
or U16592 (N_16592,N_16161,N_16261);
and U16593 (N_16593,N_16256,N_16461);
nor U16594 (N_16594,N_16462,N_16338);
nor U16595 (N_16595,N_16141,N_16272);
nand U16596 (N_16596,N_16473,N_16457);
or U16597 (N_16597,N_16268,N_16463);
and U16598 (N_16598,N_16061,N_16047);
or U16599 (N_16599,N_16013,N_16312);
nor U16600 (N_16600,N_16082,N_16440);
and U16601 (N_16601,N_16302,N_16355);
xnor U16602 (N_16602,N_16498,N_16153);
nor U16603 (N_16603,N_16067,N_16245);
xor U16604 (N_16604,N_16497,N_16162);
and U16605 (N_16605,N_16091,N_16267);
and U16606 (N_16606,N_16375,N_16023);
and U16607 (N_16607,N_16301,N_16163);
and U16608 (N_16608,N_16175,N_16073);
xor U16609 (N_16609,N_16348,N_16222);
and U16610 (N_16610,N_16234,N_16328);
or U16611 (N_16611,N_16006,N_16214);
and U16612 (N_16612,N_16353,N_16278);
xor U16613 (N_16613,N_16475,N_16076);
xnor U16614 (N_16614,N_16306,N_16100);
xnor U16615 (N_16615,N_16374,N_16401);
nor U16616 (N_16616,N_16036,N_16184);
nand U16617 (N_16617,N_16359,N_16376);
nor U16618 (N_16618,N_16094,N_16360);
nand U16619 (N_16619,N_16329,N_16282);
and U16620 (N_16620,N_16279,N_16051);
or U16621 (N_16621,N_16012,N_16239);
and U16622 (N_16622,N_16080,N_16121);
nand U16623 (N_16623,N_16041,N_16024);
nor U16624 (N_16624,N_16139,N_16045);
xnor U16625 (N_16625,N_16414,N_16085);
xnor U16626 (N_16626,N_16327,N_16286);
and U16627 (N_16627,N_16114,N_16365);
or U16628 (N_16628,N_16140,N_16104);
nand U16629 (N_16629,N_16166,N_16142);
nor U16630 (N_16630,N_16377,N_16158);
or U16631 (N_16631,N_16437,N_16105);
or U16632 (N_16632,N_16408,N_16390);
and U16633 (N_16633,N_16413,N_16060);
xnor U16634 (N_16634,N_16035,N_16049);
or U16635 (N_16635,N_16470,N_16264);
nor U16636 (N_16636,N_16387,N_16492);
xor U16637 (N_16637,N_16004,N_16460);
or U16638 (N_16638,N_16064,N_16347);
or U16639 (N_16639,N_16313,N_16084);
nor U16640 (N_16640,N_16394,N_16134);
nor U16641 (N_16641,N_16350,N_16176);
or U16642 (N_16642,N_16464,N_16283);
and U16643 (N_16643,N_16289,N_16274);
or U16644 (N_16644,N_16171,N_16172);
nor U16645 (N_16645,N_16235,N_16443);
nand U16646 (N_16646,N_16240,N_16213);
xnor U16647 (N_16647,N_16029,N_16385);
xnor U16648 (N_16648,N_16033,N_16212);
xnor U16649 (N_16649,N_16123,N_16409);
nor U16650 (N_16650,N_16448,N_16257);
or U16651 (N_16651,N_16465,N_16270);
and U16652 (N_16652,N_16275,N_16198);
nor U16653 (N_16653,N_16042,N_16021);
or U16654 (N_16654,N_16008,N_16001);
xor U16655 (N_16655,N_16128,N_16230);
or U16656 (N_16656,N_16478,N_16032);
nand U16657 (N_16657,N_16304,N_16499);
and U16658 (N_16658,N_16054,N_16450);
nand U16659 (N_16659,N_16106,N_16493);
xor U16660 (N_16660,N_16039,N_16078);
and U16661 (N_16661,N_16316,N_16159);
or U16662 (N_16662,N_16044,N_16386);
or U16663 (N_16663,N_16255,N_16216);
nor U16664 (N_16664,N_16252,N_16026);
and U16665 (N_16665,N_16421,N_16110);
or U16666 (N_16666,N_16129,N_16303);
and U16667 (N_16667,N_16373,N_16455);
nor U16668 (N_16668,N_16190,N_16219);
or U16669 (N_16669,N_16132,N_16488);
nor U16670 (N_16670,N_16384,N_16469);
nand U16671 (N_16671,N_16232,N_16108);
xnor U16672 (N_16672,N_16160,N_16185);
xnor U16673 (N_16673,N_16249,N_16248);
xnor U16674 (N_16674,N_16442,N_16490);
nor U16675 (N_16675,N_16202,N_16298);
nor U16676 (N_16676,N_16192,N_16231);
or U16677 (N_16677,N_16059,N_16322);
or U16678 (N_16678,N_16055,N_16447);
and U16679 (N_16679,N_16471,N_16101);
nor U16680 (N_16680,N_16418,N_16258);
or U16681 (N_16681,N_16182,N_16494);
or U16682 (N_16682,N_16378,N_16149);
and U16683 (N_16683,N_16250,N_16351);
nor U16684 (N_16684,N_16223,N_16135);
xnor U16685 (N_16685,N_16305,N_16487);
nand U16686 (N_16686,N_16130,N_16484);
or U16687 (N_16687,N_16211,N_16391);
or U16688 (N_16688,N_16379,N_16011);
nor U16689 (N_16689,N_16204,N_16431);
nor U16690 (N_16690,N_16034,N_16472);
and U16691 (N_16691,N_16126,N_16266);
and U16692 (N_16692,N_16072,N_16428);
or U16693 (N_16693,N_16363,N_16285);
nor U16694 (N_16694,N_16199,N_16156);
nor U16695 (N_16695,N_16367,N_16195);
and U16696 (N_16696,N_16030,N_16238);
xnor U16697 (N_16697,N_16150,N_16307);
nand U16698 (N_16698,N_16208,N_16310);
nor U16699 (N_16699,N_16370,N_16070);
or U16700 (N_16700,N_16119,N_16335);
xor U16701 (N_16701,N_16308,N_16097);
nand U16702 (N_16702,N_16253,N_16189);
or U16703 (N_16703,N_16452,N_16345);
xor U16704 (N_16704,N_16209,N_16292);
and U16705 (N_16705,N_16019,N_16358);
or U16706 (N_16706,N_16052,N_16337);
or U16707 (N_16707,N_16093,N_16102);
or U16708 (N_16708,N_16332,N_16291);
and U16709 (N_16709,N_16468,N_16383);
xor U16710 (N_16710,N_16020,N_16157);
nor U16711 (N_16711,N_16425,N_16018);
nand U16712 (N_16712,N_16297,N_16057);
nor U16713 (N_16713,N_16074,N_16339);
xnor U16714 (N_16714,N_16276,N_16459);
xnor U16715 (N_16715,N_16333,N_16362);
nand U16716 (N_16716,N_16068,N_16434);
and U16717 (N_16717,N_16177,N_16138);
or U16718 (N_16718,N_16088,N_16063);
or U16719 (N_16719,N_16112,N_16206);
or U16720 (N_16720,N_16400,N_16277);
nor U16721 (N_16721,N_16403,N_16098);
xnor U16722 (N_16722,N_16495,N_16122);
and U16723 (N_16723,N_16062,N_16244);
xor U16724 (N_16724,N_16483,N_16477);
and U16725 (N_16725,N_16296,N_16417);
or U16726 (N_16726,N_16191,N_16344);
or U16727 (N_16727,N_16424,N_16193);
xor U16728 (N_16728,N_16426,N_16205);
nor U16729 (N_16729,N_16262,N_16453);
nor U16730 (N_16730,N_16124,N_16393);
nor U16731 (N_16731,N_16372,N_16366);
xnor U16732 (N_16732,N_16423,N_16444);
and U16733 (N_16733,N_16311,N_16320);
and U16734 (N_16734,N_16486,N_16284);
xor U16735 (N_16735,N_16254,N_16154);
xnor U16736 (N_16736,N_16075,N_16186);
nand U16737 (N_16737,N_16271,N_16323);
and U16738 (N_16738,N_16113,N_16092);
nor U16739 (N_16739,N_16419,N_16207);
nand U16740 (N_16740,N_16203,N_16065);
nand U16741 (N_16741,N_16015,N_16290);
nor U16742 (N_16742,N_16476,N_16056);
and U16743 (N_16743,N_16058,N_16325);
nand U16744 (N_16744,N_16016,N_16218);
nand U16745 (N_16745,N_16027,N_16429);
nand U16746 (N_16746,N_16295,N_16194);
xor U16747 (N_16747,N_16314,N_16111);
and U16748 (N_16748,N_16038,N_16233);
nor U16749 (N_16749,N_16318,N_16406);
and U16750 (N_16750,N_16150,N_16126);
nand U16751 (N_16751,N_16373,N_16480);
nor U16752 (N_16752,N_16082,N_16408);
nor U16753 (N_16753,N_16195,N_16144);
nor U16754 (N_16754,N_16342,N_16032);
and U16755 (N_16755,N_16408,N_16315);
nor U16756 (N_16756,N_16235,N_16156);
or U16757 (N_16757,N_16416,N_16084);
and U16758 (N_16758,N_16379,N_16258);
nand U16759 (N_16759,N_16429,N_16253);
nor U16760 (N_16760,N_16241,N_16221);
nand U16761 (N_16761,N_16371,N_16007);
nand U16762 (N_16762,N_16293,N_16244);
and U16763 (N_16763,N_16427,N_16031);
xnor U16764 (N_16764,N_16316,N_16489);
nor U16765 (N_16765,N_16428,N_16379);
or U16766 (N_16766,N_16343,N_16069);
and U16767 (N_16767,N_16458,N_16043);
nand U16768 (N_16768,N_16145,N_16020);
nor U16769 (N_16769,N_16356,N_16123);
nand U16770 (N_16770,N_16425,N_16328);
nor U16771 (N_16771,N_16190,N_16406);
nor U16772 (N_16772,N_16262,N_16448);
or U16773 (N_16773,N_16013,N_16198);
nand U16774 (N_16774,N_16477,N_16219);
nor U16775 (N_16775,N_16256,N_16050);
nor U16776 (N_16776,N_16277,N_16245);
xnor U16777 (N_16777,N_16415,N_16175);
nand U16778 (N_16778,N_16406,N_16343);
xnor U16779 (N_16779,N_16166,N_16203);
and U16780 (N_16780,N_16499,N_16257);
xnor U16781 (N_16781,N_16383,N_16035);
or U16782 (N_16782,N_16167,N_16295);
nand U16783 (N_16783,N_16139,N_16382);
xor U16784 (N_16784,N_16434,N_16197);
and U16785 (N_16785,N_16492,N_16049);
xnor U16786 (N_16786,N_16299,N_16032);
nor U16787 (N_16787,N_16158,N_16441);
xnor U16788 (N_16788,N_16058,N_16168);
nor U16789 (N_16789,N_16497,N_16283);
nor U16790 (N_16790,N_16173,N_16024);
and U16791 (N_16791,N_16423,N_16234);
nand U16792 (N_16792,N_16163,N_16018);
nor U16793 (N_16793,N_16152,N_16149);
or U16794 (N_16794,N_16236,N_16321);
xor U16795 (N_16795,N_16057,N_16463);
xor U16796 (N_16796,N_16446,N_16202);
nand U16797 (N_16797,N_16305,N_16244);
or U16798 (N_16798,N_16262,N_16477);
nand U16799 (N_16799,N_16106,N_16213);
xor U16800 (N_16800,N_16446,N_16135);
xnor U16801 (N_16801,N_16344,N_16069);
nor U16802 (N_16802,N_16428,N_16488);
xor U16803 (N_16803,N_16327,N_16267);
and U16804 (N_16804,N_16440,N_16406);
or U16805 (N_16805,N_16123,N_16087);
nor U16806 (N_16806,N_16118,N_16047);
xor U16807 (N_16807,N_16069,N_16332);
xor U16808 (N_16808,N_16395,N_16119);
xor U16809 (N_16809,N_16310,N_16043);
nand U16810 (N_16810,N_16211,N_16354);
nor U16811 (N_16811,N_16109,N_16100);
and U16812 (N_16812,N_16409,N_16072);
and U16813 (N_16813,N_16083,N_16256);
or U16814 (N_16814,N_16151,N_16478);
nor U16815 (N_16815,N_16013,N_16103);
and U16816 (N_16816,N_16237,N_16095);
nor U16817 (N_16817,N_16470,N_16156);
xor U16818 (N_16818,N_16104,N_16250);
or U16819 (N_16819,N_16130,N_16165);
nor U16820 (N_16820,N_16467,N_16259);
xor U16821 (N_16821,N_16075,N_16145);
nand U16822 (N_16822,N_16410,N_16021);
nand U16823 (N_16823,N_16341,N_16253);
or U16824 (N_16824,N_16233,N_16095);
nor U16825 (N_16825,N_16341,N_16477);
and U16826 (N_16826,N_16492,N_16264);
nand U16827 (N_16827,N_16145,N_16003);
or U16828 (N_16828,N_16159,N_16023);
nor U16829 (N_16829,N_16251,N_16097);
nor U16830 (N_16830,N_16490,N_16010);
nor U16831 (N_16831,N_16455,N_16041);
nor U16832 (N_16832,N_16215,N_16314);
xnor U16833 (N_16833,N_16481,N_16362);
xor U16834 (N_16834,N_16389,N_16359);
or U16835 (N_16835,N_16444,N_16202);
nor U16836 (N_16836,N_16075,N_16313);
nand U16837 (N_16837,N_16167,N_16401);
nand U16838 (N_16838,N_16005,N_16045);
xor U16839 (N_16839,N_16001,N_16004);
nor U16840 (N_16840,N_16144,N_16193);
nand U16841 (N_16841,N_16329,N_16378);
nand U16842 (N_16842,N_16256,N_16005);
xnor U16843 (N_16843,N_16496,N_16146);
nor U16844 (N_16844,N_16308,N_16325);
xor U16845 (N_16845,N_16013,N_16179);
and U16846 (N_16846,N_16490,N_16102);
xnor U16847 (N_16847,N_16160,N_16371);
nand U16848 (N_16848,N_16135,N_16326);
xor U16849 (N_16849,N_16083,N_16302);
nor U16850 (N_16850,N_16084,N_16194);
nor U16851 (N_16851,N_16018,N_16000);
nand U16852 (N_16852,N_16245,N_16031);
xor U16853 (N_16853,N_16027,N_16166);
nand U16854 (N_16854,N_16290,N_16310);
and U16855 (N_16855,N_16271,N_16054);
nor U16856 (N_16856,N_16036,N_16074);
and U16857 (N_16857,N_16240,N_16480);
or U16858 (N_16858,N_16463,N_16301);
nor U16859 (N_16859,N_16031,N_16280);
nor U16860 (N_16860,N_16443,N_16108);
and U16861 (N_16861,N_16200,N_16446);
and U16862 (N_16862,N_16422,N_16315);
and U16863 (N_16863,N_16382,N_16279);
and U16864 (N_16864,N_16455,N_16487);
or U16865 (N_16865,N_16253,N_16254);
and U16866 (N_16866,N_16214,N_16163);
nand U16867 (N_16867,N_16406,N_16381);
and U16868 (N_16868,N_16367,N_16075);
and U16869 (N_16869,N_16336,N_16059);
and U16870 (N_16870,N_16320,N_16023);
nand U16871 (N_16871,N_16292,N_16483);
nor U16872 (N_16872,N_16089,N_16406);
and U16873 (N_16873,N_16247,N_16324);
and U16874 (N_16874,N_16221,N_16112);
nand U16875 (N_16875,N_16246,N_16285);
xor U16876 (N_16876,N_16092,N_16268);
xor U16877 (N_16877,N_16288,N_16073);
nand U16878 (N_16878,N_16271,N_16484);
nand U16879 (N_16879,N_16282,N_16161);
nor U16880 (N_16880,N_16344,N_16182);
nor U16881 (N_16881,N_16167,N_16303);
nand U16882 (N_16882,N_16055,N_16410);
or U16883 (N_16883,N_16264,N_16086);
or U16884 (N_16884,N_16373,N_16017);
or U16885 (N_16885,N_16394,N_16340);
and U16886 (N_16886,N_16138,N_16253);
nand U16887 (N_16887,N_16039,N_16458);
or U16888 (N_16888,N_16251,N_16433);
or U16889 (N_16889,N_16434,N_16151);
nor U16890 (N_16890,N_16056,N_16309);
nor U16891 (N_16891,N_16491,N_16221);
and U16892 (N_16892,N_16289,N_16193);
and U16893 (N_16893,N_16140,N_16323);
and U16894 (N_16894,N_16215,N_16354);
xor U16895 (N_16895,N_16166,N_16371);
and U16896 (N_16896,N_16247,N_16126);
nor U16897 (N_16897,N_16290,N_16002);
nand U16898 (N_16898,N_16359,N_16204);
or U16899 (N_16899,N_16245,N_16066);
and U16900 (N_16900,N_16300,N_16397);
xnor U16901 (N_16901,N_16209,N_16380);
nor U16902 (N_16902,N_16329,N_16012);
nor U16903 (N_16903,N_16074,N_16451);
nand U16904 (N_16904,N_16074,N_16203);
nand U16905 (N_16905,N_16201,N_16164);
and U16906 (N_16906,N_16142,N_16481);
xor U16907 (N_16907,N_16404,N_16011);
or U16908 (N_16908,N_16476,N_16416);
and U16909 (N_16909,N_16374,N_16246);
nor U16910 (N_16910,N_16291,N_16386);
or U16911 (N_16911,N_16214,N_16397);
and U16912 (N_16912,N_16391,N_16461);
xnor U16913 (N_16913,N_16117,N_16045);
or U16914 (N_16914,N_16138,N_16093);
xnor U16915 (N_16915,N_16268,N_16300);
xor U16916 (N_16916,N_16456,N_16271);
nand U16917 (N_16917,N_16239,N_16071);
nor U16918 (N_16918,N_16179,N_16074);
or U16919 (N_16919,N_16111,N_16437);
nor U16920 (N_16920,N_16034,N_16032);
or U16921 (N_16921,N_16111,N_16272);
xnor U16922 (N_16922,N_16365,N_16157);
nand U16923 (N_16923,N_16341,N_16011);
xnor U16924 (N_16924,N_16218,N_16126);
xor U16925 (N_16925,N_16366,N_16210);
or U16926 (N_16926,N_16423,N_16392);
or U16927 (N_16927,N_16065,N_16288);
or U16928 (N_16928,N_16274,N_16295);
nand U16929 (N_16929,N_16004,N_16316);
or U16930 (N_16930,N_16067,N_16463);
and U16931 (N_16931,N_16416,N_16183);
or U16932 (N_16932,N_16436,N_16086);
and U16933 (N_16933,N_16243,N_16009);
and U16934 (N_16934,N_16319,N_16268);
or U16935 (N_16935,N_16477,N_16368);
nand U16936 (N_16936,N_16164,N_16112);
nor U16937 (N_16937,N_16066,N_16210);
nand U16938 (N_16938,N_16423,N_16224);
nor U16939 (N_16939,N_16492,N_16287);
or U16940 (N_16940,N_16389,N_16049);
nand U16941 (N_16941,N_16250,N_16258);
nand U16942 (N_16942,N_16167,N_16247);
nand U16943 (N_16943,N_16363,N_16343);
or U16944 (N_16944,N_16341,N_16089);
nand U16945 (N_16945,N_16151,N_16173);
or U16946 (N_16946,N_16380,N_16107);
nand U16947 (N_16947,N_16203,N_16128);
nor U16948 (N_16948,N_16304,N_16316);
xnor U16949 (N_16949,N_16198,N_16426);
and U16950 (N_16950,N_16088,N_16131);
xnor U16951 (N_16951,N_16199,N_16044);
xnor U16952 (N_16952,N_16291,N_16277);
nand U16953 (N_16953,N_16367,N_16435);
xnor U16954 (N_16954,N_16463,N_16113);
and U16955 (N_16955,N_16418,N_16246);
nor U16956 (N_16956,N_16112,N_16472);
nor U16957 (N_16957,N_16262,N_16114);
nor U16958 (N_16958,N_16152,N_16027);
xnor U16959 (N_16959,N_16224,N_16274);
nor U16960 (N_16960,N_16052,N_16227);
xnor U16961 (N_16961,N_16497,N_16351);
nor U16962 (N_16962,N_16155,N_16499);
nand U16963 (N_16963,N_16340,N_16315);
nand U16964 (N_16964,N_16095,N_16117);
nand U16965 (N_16965,N_16314,N_16076);
and U16966 (N_16966,N_16173,N_16340);
xnor U16967 (N_16967,N_16417,N_16020);
xor U16968 (N_16968,N_16395,N_16323);
nand U16969 (N_16969,N_16134,N_16276);
and U16970 (N_16970,N_16265,N_16081);
xor U16971 (N_16971,N_16404,N_16048);
or U16972 (N_16972,N_16206,N_16060);
nand U16973 (N_16973,N_16010,N_16466);
or U16974 (N_16974,N_16070,N_16407);
nor U16975 (N_16975,N_16318,N_16139);
or U16976 (N_16976,N_16438,N_16324);
nand U16977 (N_16977,N_16379,N_16176);
or U16978 (N_16978,N_16359,N_16207);
or U16979 (N_16979,N_16115,N_16341);
nor U16980 (N_16980,N_16148,N_16132);
or U16981 (N_16981,N_16359,N_16394);
nor U16982 (N_16982,N_16474,N_16477);
nor U16983 (N_16983,N_16051,N_16103);
nor U16984 (N_16984,N_16427,N_16017);
and U16985 (N_16985,N_16243,N_16139);
nor U16986 (N_16986,N_16200,N_16010);
xor U16987 (N_16987,N_16018,N_16344);
nand U16988 (N_16988,N_16201,N_16323);
or U16989 (N_16989,N_16327,N_16219);
nor U16990 (N_16990,N_16452,N_16149);
xor U16991 (N_16991,N_16354,N_16157);
or U16992 (N_16992,N_16480,N_16328);
or U16993 (N_16993,N_16131,N_16135);
or U16994 (N_16994,N_16417,N_16307);
xor U16995 (N_16995,N_16104,N_16109);
xnor U16996 (N_16996,N_16140,N_16219);
xnor U16997 (N_16997,N_16380,N_16409);
and U16998 (N_16998,N_16161,N_16336);
xnor U16999 (N_16999,N_16093,N_16370);
nor U17000 (N_17000,N_16564,N_16754);
and U17001 (N_17001,N_16607,N_16656);
and U17002 (N_17002,N_16994,N_16649);
nand U17003 (N_17003,N_16655,N_16912);
nor U17004 (N_17004,N_16904,N_16888);
xor U17005 (N_17005,N_16843,N_16879);
nor U17006 (N_17006,N_16702,N_16622);
nor U17007 (N_17007,N_16560,N_16943);
and U17008 (N_17008,N_16821,N_16990);
and U17009 (N_17009,N_16529,N_16871);
nor U17010 (N_17010,N_16900,N_16988);
nand U17011 (N_17011,N_16926,N_16619);
xor U17012 (N_17012,N_16909,N_16767);
nand U17013 (N_17013,N_16770,N_16945);
and U17014 (N_17014,N_16750,N_16877);
nor U17015 (N_17015,N_16747,N_16922);
xnor U17016 (N_17016,N_16615,N_16598);
nor U17017 (N_17017,N_16586,N_16882);
or U17018 (N_17018,N_16813,N_16708);
nand U17019 (N_17019,N_16520,N_16844);
nand U17020 (N_17020,N_16938,N_16775);
nand U17021 (N_17021,N_16704,N_16925);
xor U17022 (N_17022,N_16881,N_16939);
or U17023 (N_17023,N_16531,N_16614);
and U17024 (N_17024,N_16631,N_16974);
xor U17025 (N_17025,N_16737,N_16793);
nand U17026 (N_17026,N_16846,N_16908);
nand U17027 (N_17027,N_16661,N_16823);
nor U17028 (N_17028,N_16694,N_16911);
xor U17029 (N_17029,N_16583,N_16508);
nand U17030 (N_17030,N_16804,N_16735);
xnor U17031 (N_17031,N_16637,N_16776);
nor U17032 (N_17032,N_16645,N_16812);
nand U17033 (N_17033,N_16517,N_16957);
xor U17034 (N_17034,N_16733,N_16653);
xnor U17035 (N_17035,N_16646,N_16968);
xor U17036 (N_17036,N_16633,N_16800);
nor U17037 (N_17037,N_16684,N_16907);
xor U17038 (N_17038,N_16755,N_16666);
and U17039 (N_17039,N_16601,N_16841);
nand U17040 (N_17040,N_16621,N_16618);
nand U17041 (N_17041,N_16967,N_16713);
nor U17042 (N_17042,N_16566,N_16616);
nand U17043 (N_17043,N_16721,N_16978);
or U17044 (N_17044,N_16758,N_16732);
nor U17045 (N_17045,N_16654,N_16710);
and U17046 (N_17046,N_16950,N_16580);
nand U17047 (N_17047,N_16946,N_16860);
xnor U17048 (N_17048,N_16830,N_16986);
nand U17049 (N_17049,N_16647,N_16878);
or U17050 (N_17050,N_16715,N_16759);
and U17051 (N_17051,N_16839,N_16515);
or U17052 (N_17052,N_16769,N_16525);
nor U17053 (N_17053,N_16546,N_16667);
or U17054 (N_17054,N_16507,N_16849);
nand U17055 (N_17055,N_16783,N_16917);
xor U17056 (N_17056,N_16940,N_16850);
nand U17057 (N_17057,N_16673,N_16924);
and U17058 (N_17058,N_16691,N_16728);
nor U17059 (N_17059,N_16724,N_16902);
xnor U17060 (N_17060,N_16640,N_16863);
nor U17061 (N_17061,N_16548,N_16698);
nor U17062 (N_17062,N_16824,N_16512);
nand U17063 (N_17063,N_16829,N_16976);
xnor U17064 (N_17064,N_16751,N_16991);
nand U17065 (N_17065,N_16772,N_16901);
nor U17066 (N_17066,N_16719,N_16869);
and U17067 (N_17067,N_16858,N_16791);
or U17068 (N_17068,N_16592,N_16636);
or U17069 (N_17069,N_16962,N_16969);
and U17070 (N_17070,N_16827,N_16742);
nand U17071 (N_17071,N_16762,N_16630);
xnor U17072 (N_17072,N_16979,N_16574);
nor U17073 (N_17073,N_16761,N_16953);
or U17074 (N_17074,N_16500,N_16789);
and U17075 (N_17075,N_16628,N_16689);
or U17076 (N_17076,N_16572,N_16778);
nor U17077 (N_17077,N_16868,N_16952);
nor U17078 (N_17078,N_16563,N_16683);
xnor U17079 (N_17079,N_16893,N_16537);
and U17080 (N_17080,N_16519,N_16748);
and U17081 (N_17081,N_16916,N_16632);
or U17082 (N_17082,N_16584,N_16588);
nor U17083 (N_17083,N_16623,N_16932);
or U17084 (N_17084,N_16716,N_16831);
xnor U17085 (N_17085,N_16502,N_16725);
nand U17086 (N_17086,N_16826,N_16717);
or U17087 (N_17087,N_16852,N_16526);
xor U17088 (N_17088,N_16806,N_16650);
nand U17089 (N_17089,N_16641,N_16987);
xnor U17090 (N_17090,N_16738,N_16652);
and U17091 (N_17091,N_16712,N_16971);
nand U17092 (N_17092,N_16861,N_16982);
xnor U17093 (N_17093,N_16921,N_16859);
nand U17094 (N_17094,N_16534,N_16948);
nand U17095 (N_17095,N_16707,N_16746);
nand U17096 (N_17096,N_16509,N_16550);
nand U17097 (N_17097,N_16533,N_16568);
xor U17098 (N_17098,N_16571,N_16782);
or U17099 (N_17099,N_16808,N_16536);
or U17100 (N_17100,N_16595,N_16892);
nor U17101 (N_17101,N_16577,N_16788);
or U17102 (N_17102,N_16599,N_16954);
xnor U17103 (N_17103,N_16884,N_16856);
nor U17104 (N_17104,N_16543,N_16559);
or U17105 (N_17105,N_16608,N_16591);
nand U17106 (N_17106,N_16851,N_16765);
nor U17107 (N_17107,N_16933,N_16557);
or U17108 (N_17108,N_16573,N_16729);
xor U17109 (N_17109,N_16690,N_16873);
nor U17110 (N_17110,N_16828,N_16795);
xnor U17111 (N_17111,N_16749,N_16722);
nor U17112 (N_17112,N_16874,N_16555);
xnor U17113 (N_17113,N_16740,N_16842);
or U17114 (N_17114,N_16699,N_16915);
xor U17115 (N_17115,N_16886,N_16743);
xnor U17116 (N_17116,N_16705,N_16671);
xor U17117 (N_17117,N_16644,N_16910);
or U17118 (N_17118,N_16518,N_16984);
and U17119 (N_17119,N_16538,N_16549);
or U17120 (N_17120,N_16567,N_16668);
or U17121 (N_17121,N_16613,N_16585);
and U17122 (N_17122,N_16697,N_16956);
nor U17123 (N_17123,N_16565,N_16899);
or U17124 (N_17124,N_16961,N_16777);
nor U17125 (N_17125,N_16927,N_16784);
and U17126 (N_17126,N_16966,N_16973);
xnor U17127 (N_17127,N_16674,N_16611);
xnor U17128 (N_17128,N_16532,N_16540);
nand U17129 (N_17129,N_16739,N_16744);
and U17130 (N_17130,N_16541,N_16745);
xnor U17131 (N_17131,N_16706,N_16686);
and U17132 (N_17132,N_16685,N_16773);
nor U17133 (N_17133,N_16731,N_16524);
xor U17134 (N_17134,N_16894,N_16810);
and U17135 (N_17135,N_16896,N_16937);
or U17136 (N_17136,N_16928,N_16678);
nand U17137 (N_17137,N_16734,N_16503);
or U17138 (N_17138,N_16709,N_16799);
and U17139 (N_17139,N_16620,N_16774);
and U17140 (N_17140,N_16781,N_16651);
nor U17141 (N_17141,N_16752,N_16594);
or U17142 (N_17142,N_16576,N_16934);
xor U17143 (N_17143,N_16642,N_16786);
xnor U17144 (N_17144,N_16960,N_16870);
or U17145 (N_17145,N_16687,N_16589);
nor U17146 (N_17146,N_16547,N_16511);
xnor U17147 (N_17147,N_16883,N_16897);
nor U17148 (N_17148,N_16836,N_16539);
xnor U17149 (N_17149,N_16720,N_16914);
nand U17150 (N_17150,N_16885,N_16581);
or U17151 (N_17151,N_16544,N_16692);
and U17152 (N_17152,N_16889,N_16562);
and U17153 (N_17153,N_16918,N_16913);
nor U17154 (N_17154,N_16999,N_16768);
nand U17155 (N_17155,N_16835,N_16787);
nor U17156 (N_17156,N_16514,N_16792);
nor U17157 (N_17157,N_16756,N_16741);
and U17158 (N_17158,N_16553,N_16609);
nor U17159 (N_17159,N_16981,N_16880);
and U17160 (N_17160,N_16834,N_16854);
nor U17161 (N_17161,N_16951,N_16643);
nand U17162 (N_17162,N_16985,N_16955);
or U17163 (N_17163,N_16794,N_16865);
or U17164 (N_17164,N_16510,N_16963);
nor U17165 (N_17165,N_16809,N_16818);
xnor U17166 (N_17166,N_16504,N_16838);
and U17167 (N_17167,N_16605,N_16680);
xor U17168 (N_17168,N_16663,N_16887);
xnor U17169 (N_17169,N_16848,N_16675);
xor U17170 (N_17170,N_16891,N_16993);
nor U17171 (N_17171,N_16554,N_16949);
xnor U17172 (N_17172,N_16992,N_16528);
nor U17173 (N_17173,N_16664,N_16657);
xor U17174 (N_17174,N_16895,N_16872);
or U17175 (N_17175,N_16972,N_16682);
xnor U17176 (N_17176,N_16558,N_16864);
xor U17177 (N_17177,N_16505,N_16530);
or U17178 (N_17178,N_16561,N_16989);
nand U17179 (N_17179,N_16796,N_16638);
xnor U17180 (N_17180,N_16736,N_16857);
xnor U17181 (N_17181,N_16906,N_16771);
nand U17182 (N_17182,N_16730,N_16764);
or U17183 (N_17183,N_16941,N_16822);
nand U17184 (N_17184,N_16617,N_16814);
nor U17185 (N_17185,N_16662,N_16820);
or U17186 (N_17186,N_16660,N_16714);
or U17187 (N_17187,N_16805,N_16701);
and U17188 (N_17188,N_16875,N_16596);
xor U17189 (N_17189,N_16629,N_16898);
xnor U17190 (N_17190,N_16876,N_16819);
and U17191 (N_17191,N_16501,N_16527);
or U17192 (N_17192,N_16693,N_16696);
or U17193 (N_17193,N_16626,N_16610);
or U17194 (N_17194,N_16634,N_16700);
xnor U17195 (N_17195,N_16658,N_16837);
nor U17196 (N_17196,N_16965,N_16582);
nor U17197 (N_17197,N_16718,N_16801);
or U17198 (N_17198,N_16726,N_16997);
or U17199 (N_17199,N_16817,N_16723);
or U17200 (N_17200,N_16923,N_16513);
or U17201 (N_17201,N_16798,N_16867);
and U17202 (N_17202,N_16995,N_16944);
xor U17203 (N_17203,N_16807,N_16688);
nor U17204 (N_17204,N_16803,N_16523);
nand U17205 (N_17205,N_16604,N_16845);
xnor U17206 (N_17206,N_16996,N_16711);
xor U17207 (N_17207,N_16551,N_16569);
and U17208 (N_17208,N_16975,N_16606);
xnor U17209 (N_17209,N_16625,N_16603);
or U17210 (N_17210,N_16600,N_16590);
nor U17211 (N_17211,N_16942,N_16624);
or U17212 (N_17212,N_16905,N_16797);
nand U17213 (N_17213,N_16983,N_16766);
nor U17214 (N_17214,N_16677,N_16847);
nor U17215 (N_17215,N_16935,N_16556);
nand U17216 (N_17216,N_16627,N_16840);
nor U17217 (N_17217,N_16665,N_16780);
or U17218 (N_17218,N_16866,N_16575);
or U17219 (N_17219,N_16931,N_16597);
and U17220 (N_17220,N_16579,N_16679);
nand U17221 (N_17221,N_16832,N_16648);
xnor U17222 (N_17222,N_16676,N_16672);
nor U17223 (N_17223,N_16980,N_16578);
or U17224 (N_17224,N_16958,N_16587);
nand U17225 (N_17225,N_16964,N_16760);
or U17226 (N_17226,N_16753,N_16790);
nor U17227 (N_17227,N_16903,N_16816);
or U17228 (N_17228,N_16602,N_16542);
xnor U17229 (N_17229,N_16785,N_16612);
xnor U17230 (N_17230,N_16890,N_16855);
or U17231 (N_17231,N_16535,N_16977);
and U17232 (N_17232,N_16833,N_16635);
or U17233 (N_17233,N_16670,N_16936);
xor U17234 (N_17234,N_16521,N_16802);
nor U17235 (N_17235,N_16763,N_16919);
nor U17236 (N_17236,N_16970,N_16727);
nor U17237 (N_17237,N_16669,N_16779);
and U17238 (N_17238,N_16703,N_16681);
and U17239 (N_17239,N_16659,N_16930);
and U17240 (N_17240,N_16639,N_16998);
and U17241 (N_17241,N_16920,N_16929);
xor U17242 (N_17242,N_16947,N_16757);
nand U17243 (N_17243,N_16545,N_16815);
or U17244 (N_17244,N_16853,N_16862);
nor U17245 (N_17245,N_16552,N_16593);
or U17246 (N_17246,N_16811,N_16506);
or U17247 (N_17247,N_16695,N_16570);
or U17248 (N_17248,N_16959,N_16522);
nand U17249 (N_17249,N_16516,N_16825);
and U17250 (N_17250,N_16919,N_16762);
and U17251 (N_17251,N_16682,N_16694);
or U17252 (N_17252,N_16923,N_16762);
or U17253 (N_17253,N_16635,N_16849);
or U17254 (N_17254,N_16501,N_16863);
or U17255 (N_17255,N_16918,N_16621);
nand U17256 (N_17256,N_16663,N_16899);
nand U17257 (N_17257,N_16983,N_16513);
or U17258 (N_17258,N_16519,N_16948);
xnor U17259 (N_17259,N_16654,N_16863);
nor U17260 (N_17260,N_16808,N_16607);
nor U17261 (N_17261,N_16765,N_16803);
or U17262 (N_17262,N_16621,N_16527);
and U17263 (N_17263,N_16525,N_16858);
nor U17264 (N_17264,N_16553,N_16946);
and U17265 (N_17265,N_16837,N_16736);
xnor U17266 (N_17266,N_16796,N_16514);
or U17267 (N_17267,N_16696,N_16850);
or U17268 (N_17268,N_16624,N_16881);
nor U17269 (N_17269,N_16657,N_16865);
or U17270 (N_17270,N_16762,N_16578);
nor U17271 (N_17271,N_16740,N_16961);
xnor U17272 (N_17272,N_16677,N_16588);
and U17273 (N_17273,N_16507,N_16902);
or U17274 (N_17274,N_16542,N_16639);
nor U17275 (N_17275,N_16756,N_16763);
xnor U17276 (N_17276,N_16740,N_16918);
nand U17277 (N_17277,N_16522,N_16845);
nor U17278 (N_17278,N_16990,N_16977);
and U17279 (N_17279,N_16780,N_16551);
or U17280 (N_17280,N_16617,N_16552);
and U17281 (N_17281,N_16658,N_16894);
and U17282 (N_17282,N_16909,N_16879);
and U17283 (N_17283,N_16706,N_16566);
xnor U17284 (N_17284,N_16932,N_16565);
xor U17285 (N_17285,N_16921,N_16799);
xor U17286 (N_17286,N_16934,N_16693);
and U17287 (N_17287,N_16967,N_16568);
or U17288 (N_17288,N_16506,N_16771);
nand U17289 (N_17289,N_16740,N_16883);
xor U17290 (N_17290,N_16595,N_16851);
nand U17291 (N_17291,N_16560,N_16732);
nor U17292 (N_17292,N_16624,N_16616);
xnor U17293 (N_17293,N_16541,N_16632);
xnor U17294 (N_17294,N_16680,N_16837);
xnor U17295 (N_17295,N_16833,N_16670);
or U17296 (N_17296,N_16727,N_16770);
nand U17297 (N_17297,N_16577,N_16800);
nand U17298 (N_17298,N_16801,N_16620);
nor U17299 (N_17299,N_16840,N_16911);
or U17300 (N_17300,N_16528,N_16936);
and U17301 (N_17301,N_16941,N_16840);
xnor U17302 (N_17302,N_16802,N_16582);
nor U17303 (N_17303,N_16897,N_16778);
nand U17304 (N_17304,N_16707,N_16861);
nand U17305 (N_17305,N_16877,N_16572);
xor U17306 (N_17306,N_16750,N_16983);
xor U17307 (N_17307,N_16935,N_16517);
xnor U17308 (N_17308,N_16508,N_16870);
nand U17309 (N_17309,N_16834,N_16662);
xor U17310 (N_17310,N_16788,N_16796);
or U17311 (N_17311,N_16690,N_16819);
and U17312 (N_17312,N_16572,N_16619);
nor U17313 (N_17313,N_16885,N_16698);
nand U17314 (N_17314,N_16621,N_16533);
or U17315 (N_17315,N_16536,N_16878);
and U17316 (N_17316,N_16553,N_16971);
or U17317 (N_17317,N_16752,N_16707);
xor U17318 (N_17318,N_16877,N_16960);
xor U17319 (N_17319,N_16672,N_16651);
nor U17320 (N_17320,N_16502,N_16887);
xnor U17321 (N_17321,N_16923,N_16580);
nand U17322 (N_17322,N_16924,N_16821);
nand U17323 (N_17323,N_16899,N_16500);
xnor U17324 (N_17324,N_16568,N_16609);
nor U17325 (N_17325,N_16836,N_16977);
nand U17326 (N_17326,N_16876,N_16674);
xnor U17327 (N_17327,N_16626,N_16785);
xor U17328 (N_17328,N_16658,N_16538);
xnor U17329 (N_17329,N_16782,N_16935);
or U17330 (N_17330,N_16848,N_16918);
xor U17331 (N_17331,N_16674,N_16545);
nor U17332 (N_17332,N_16590,N_16946);
xnor U17333 (N_17333,N_16709,N_16995);
nand U17334 (N_17334,N_16557,N_16705);
xor U17335 (N_17335,N_16822,N_16759);
and U17336 (N_17336,N_16519,N_16570);
nand U17337 (N_17337,N_16503,N_16696);
and U17338 (N_17338,N_16887,N_16630);
nor U17339 (N_17339,N_16603,N_16802);
nor U17340 (N_17340,N_16931,N_16646);
or U17341 (N_17341,N_16616,N_16966);
and U17342 (N_17342,N_16746,N_16684);
and U17343 (N_17343,N_16671,N_16676);
or U17344 (N_17344,N_16613,N_16614);
nand U17345 (N_17345,N_16514,N_16616);
nand U17346 (N_17346,N_16828,N_16996);
and U17347 (N_17347,N_16819,N_16803);
and U17348 (N_17348,N_16673,N_16972);
nor U17349 (N_17349,N_16830,N_16870);
nor U17350 (N_17350,N_16924,N_16965);
nor U17351 (N_17351,N_16746,N_16802);
nand U17352 (N_17352,N_16903,N_16579);
and U17353 (N_17353,N_16786,N_16832);
nor U17354 (N_17354,N_16670,N_16909);
nand U17355 (N_17355,N_16617,N_16743);
nor U17356 (N_17356,N_16601,N_16970);
nor U17357 (N_17357,N_16953,N_16807);
or U17358 (N_17358,N_16525,N_16842);
nand U17359 (N_17359,N_16842,N_16775);
nor U17360 (N_17360,N_16591,N_16996);
or U17361 (N_17361,N_16997,N_16993);
xor U17362 (N_17362,N_16852,N_16610);
xor U17363 (N_17363,N_16770,N_16707);
and U17364 (N_17364,N_16610,N_16865);
xor U17365 (N_17365,N_16677,N_16729);
nor U17366 (N_17366,N_16729,N_16759);
nand U17367 (N_17367,N_16631,N_16965);
and U17368 (N_17368,N_16735,N_16914);
nor U17369 (N_17369,N_16925,N_16511);
or U17370 (N_17370,N_16897,N_16594);
xnor U17371 (N_17371,N_16918,N_16648);
nor U17372 (N_17372,N_16771,N_16987);
nand U17373 (N_17373,N_16802,N_16767);
or U17374 (N_17374,N_16732,N_16642);
and U17375 (N_17375,N_16548,N_16950);
xnor U17376 (N_17376,N_16848,N_16905);
nand U17377 (N_17377,N_16557,N_16531);
nand U17378 (N_17378,N_16925,N_16836);
or U17379 (N_17379,N_16698,N_16874);
nor U17380 (N_17380,N_16928,N_16813);
and U17381 (N_17381,N_16961,N_16706);
or U17382 (N_17382,N_16526,N_16755);
and U17383 (N_17383,N_16602,N_16851);
and U17384 (N_17384,N_16869,N_16923);
xor U17385 (N_17385,N_16708,N_16882);
xor U17386 (N_17386,N_16704,N_16632);
nand U17387 (N_17387,N_16557,N_16981);
and U17388 (N_17388,N_16983,N_16825);
and U17389 (N_17389,N_16528,N_16543);
or U17390 (N_17390,N_16681,N_16818);
xnor U17391 (N_17391,N_16573,N_16683);
and U17392 (N_17392,N_16662,N_16579);
or U17393 (N_17393,N_16813,N_16992);
nor U17394 (N_17394,N_16540,N_16712);
or U17395 (N_17395,N_16647,N_16810);
nor U17396 (N_17396,N_16582,N_16670);
xnor U17397 (N_17397,N_16707,N_16641);
nor U17398 (N_17398,N_16663,N_16655);
or U17399 (N_17399,N_16627,N_16887);
nor U17400 (N_17400,N_16977,N_16500);
nor U17401 (N_17401,N_16828,N_16503);
and U17402 (N_17402,N_16500,N_16609);
xnor U17403 (N_17403,N_16850,N_16915);
xnor U17404 (N_17404,N_16751,N_16900);
nor U17405 (N_17405,N_16600,N_16787);
xnor U17406 (N_17406,N_16605,N_16774);
nor U17407 (N_17407,N_16558,N_16797);
nor U17408 (N_17408,N_16678,N_16851);
and U17409 (N_17409,N_16987,N_16745);
nand U17410 (N_17410,N_16834,N_16850);
nand U17411 (N_17411,N_16615,N_16683);
xor U17412 (N_17412,N_16909,N_16934);
nor U17413 (N_17413,N_16836,N_16893);
or U17414 (N_17414,N_16814,N_16588);
nand U17415 (N_17415,N_16523,N_16878);
nor U17416 (N_17416,N_16631,N_16755);
nand U17417 (N_17417,N_16947,N_16815);
and U17418 (N_17418,N_16650,N_16864);
or U17419 (N_17419,N_16992,N_16943);
and U17420 (N_17420,N_16851,N_16500);
nand U17421 (N_17421,N_16875,N_16635);
xnor U17422 (N_17422,N_16981,N_16798);
nand U17423 (N_17423,N_16643,N_16627);
and U17424 (N_17424,N_16906,N_16504);
and U17425 (N_17425,N_16775,N_16774);
and U17426 (N_17426,N_16633,N_16897);
xor U17427 (N_17427,N_16906,N_16958);
xnor U17428 (N_17428,N_16707,N_16665);
nand U17429 (N_17429,N_16861,N_16751);
xor U17430 (N_17430,N_16949,N_16781);
nor U17431 (N_17431,N_16798,N_16668);
nor U17432 (N_17432,N_16971,N_16741);
nand U17433 (N_17433,N_16517,N_16663);
nand U17434 (N_17434,N_16720,N_16856);
nor U17435 (N_17435,N_16894,N_16518);
or U17436 (N_17436,N_16830,N_16596);
nor U17437 (N_17437,N_16589,N_16594);
nor U17438 (N_17438,N_16882,N_16627);
nand U17439 (N_17439,N_16610,N_16589);
or U17440 (N_17440,N_16692,N_16735);
nand U17441 (N_17441,N_16941,N_16693);
nand U17442 (N_17442,N_16580,N_16875);
and U17443 (N_17443,N_16831,N_16907);
and U17444 (N_17444,N_16815,N_16779);
nor U17445 (N_17445,N_16985,N_16979);
nand U17446 (N_17446,N_16742,N_16569);
and U17447 (N_17447,N_16667,N_16849);
nor U17448 (N_17448,N_16950,N_16626);
or U17449 (N_17449,N_16825,N_16958);
or U17450 (N_17450,N_16860,N_16760);
nor U17451 (N_17451,N_16742,N_16692);
or U17452 (N_17452,N_16831,N_16525);
or U17453 (N_17453,N_16603,N_16757);
nor U17454 (N_17454,N_16806,N_16888);
and U17455 (N_17455,N_16630,N_16639);
and U17456 (N_17456,N_16809,N_16887);
xnor U17457 (N_17457,N_16668,N_16941);
and U17458 (N_17458,N_16936,N_16865);
xnor U17459 (N_17459,N_16653,N_16907);
nand U17460 (N_17460,N_16835,N_16850);
nand U17461 (N_17461,N_16667,N_16820);
or U17462 (N_17462,N_16545,N_16667);
xnor U17463 (N_17463,N_16585,N_16761);
nand U17464 (N_17464,N_16595,N_16920);
nor U17465 (N_17465,N_16811,N_16747);
xor U17466 (N_17466,N_16709,N_16981);
nor U17467 (N_17467,N_16548,N_16533);
nor U17468 (N_17468,N_16547,N_16926);
nor U17469 (N_17469,N_16692,N_16922);
or U17470 (N_17470,N_16971,N_16729);
and U17471 (N_17471,N_16751,N_16740);
nand U17472 (N_17472,N_16848,N_16964);
and U17473 (N_17473,N_16926,N_16684);
nor U17474 (N_17474,N_16808,N_16876);
nand U17475 (N_17475,N_16847,N_16800);
and U17476 (N_17476,N_16736,N_16685);
xnor U17477 (N_17477,N_16769,N_16694);
xor U17478 (N_17478,N_16601,N_16736);
and U17479 (N_17479,N_16711,N_16951);
or U17480 (N_17480,N_16876,N_16729);
nor U17481 (N_17481,N_16758,N_16547);
and U17482 (N_17482,N_16568,N_16660);
nand U17483 (N_17483,N_16588,N_16766);
and U17484 (N_17484,N_16743,N_16727);
nand U17485 (N_17485,N_16675,N_16764);
and U17486 (N_17486,N_16991,N_16711);
or U17487 (N_17487,N_16507,N_16623);
xor U17488 (N_17488,N_16671,N_16654);
xnor U17489 (N_17489,N_16589,N_16547);
xor U17490 (N_17490,N_16525,N_16533);
or U17491 (N_17491,N_16517,N_16721);
nand U17492 (N_17492,N_16944,N_16558);
xor U17493 (N_17493,N_16750,N_16841);
xor U17494 (N_17494,N_16683,N_16689);
nor U17495 (N_17495,N_16708,N_16666);
or U17496 (N_17496,N_16973,N_16536);
nor U17497 (N_17497,N_16765,N_16503);
or U17498 (N_17498,N_16897,N_16651);
nand U17499 (N_17499,N_16591,N_16612);
xnor U17500 (N_17500,N_17184,N_17476);
nand U17501 (N_17501,N_17088,N_17411);
or U17502 (N_17502,N_17094,N_17404);
nor U17503 (N_17503,N_17067,N_17024);
and U17504 (N_17504,N_17402,N_17459);
nor U17505 (N_17505,N_17393,N_17110);
xnor U17506 (N_17506,N_17019,N_17320);
and U17507 (N_17507,N_17185,N_17062);
or U17508 (N_17508,N_17315,N_17342);
xnor U17509 (N_17509,N_17008,N_17415);
nand U17510 (N_17510,N_17131,N_17498);
nand U17511 (N_17511,N_17302,N_17198);
nand U17512 (N_17512,N_17406,N_17297);
nand U17513 (N_17513,N_17061,N_17467);
nor U17514 (N_17514,N_17075,N_17105);
nand U17515 (N_17515,N_17041,N_17479);
xor U17516 (N_17516,N_17109,N_17176);
xor U17517 (N_17517,N_17432,N_17240);
nand U17518 (N_17518,N_17304,N_17214);
nand U17519 (N_17519,N_17123,N_17038);
and U17520 (N_17520,N_17349,N_17051);
nor U17521 (N_17521,N_17407,N_17048);
or U17522 (N_17522,N_17028,N_17483);
and U17523 (N_17523,N_17171,N_17063);
nor U17524 (N_17524,N_17283,N_17260);
or U17525 (N_17525,N_17485,N_17301);
nand U17526 (N_17526,N_17225,N_17080);
nor U17527 (N_17527,N_17356,N_17375);
xor U17528 (N_17528,N_17420,N_17231);
xnor U17529 (N_17529,N_17336,N_17433);
xnor U17530 (N_17530,N_17492,N_17368);
nand U17531 (N_17531,N_17427,N_17023);
nand U17532 (N_17532,N_17258,N_17195);
or U17533 (N_17533,N_17106,N_17285);
or U17534 (N_17534,N_17348,N_17142);
nor U17535 (N_17535,N_17376,N_17371);
nor U17536 (N_17536,N_17448,N_17352);
nand U17537 (N_17537,N_17263,N_17175);
or U17538 (N_17538,N_17280,N_17272);
and U17539 (N_17539,N_17383,N_17042);
nor U17540 (N_17540,N_17317,N_17345);
nand U17541 (N_17541,N_17437,N_17238);
nor U17542 (N_17542,N_17457,N_17463);
nor U17543 (N_17543,N_17187,N_17084);
xor U17544 (N_17544,N_17212,N_17453);
xnor U17545 (N_17545,N_17021,N_17097);
and U17546 (N_17546,N_17425,N_17070);
and U17547 (N_17547,N_17226,N_17354);
nor U17548 (N_17548,N_17441,N_17318);
xor U17549 (N_17549,N_17452,N_17409);
and U17550 (N_17550,N_17087,N_17188);
or U17551 (N_17551,N_17194,N_17493);
xnor U17552 (N_17552,N_17093,N_17341);
and U17553 (N_17553,N_17365,N_17209);
or U17554 (N_17554,N_17189,N_17273);
xor U17555 (N_17555,N_17099,N_17363);
and U17556 (N_17556,N_17073,N_17327);
nand U17557 (N_17557,N_17149,N_17165);
nand U17558 (N_17558,N_17282,N_17193);
and U17559 (N_17559,N_17090,N_17435);
or U17560 (N_17560,N_17034,N_17169);
xnor U17561 (N_17561,N_17174,N_17361);
nor U17562 (N_17562,N_17092,N_17072);
or U17563 (N_17563,N_17036,N_17192);
nor U17564 (N_17564,N_17478,N_17446);
nand U17565 (N_17565,N_17253,N_17166);
nor U17566 (N_17566,N_17265,N_17221);
xnor U17567 (N_17567,N_17381,N_17489);
nor U17568 (N_17568,N_17410,N_17074);
nor U17569 (N_17569,N_17141,N_17360);
xor U17570 (N_17570,N_17306,N_17333);
nand U17571 (N_17571,N_17113,N_17119);
xor U17572 (N_17572,N_17292,N_17029);
nor U17573 (N_17573,N_17451,N_17482);
nand U17574 (N_17574,N_17136,N_17199);
nor U17575 (N_17575,N_17264,N_17138);
nor U17576 (N_17576,N_17328,N_17178);
xor U17577 (N_17577,N_17422,N_17372);
and U17578 (N_17578,N_17224,N_17126);
xnor U17579 (N_17579,N_17152,N_17268);
nor U17580 (N_17580,N_17112,N_17168);
xnor U17581 (N_17581,N_17431,N_17229);
nor U17582 (N_17582,N_17191,N_17103);
and U17583 (N_17583,N_17267,N_17274);
nand U17584 (N_17584,N_17252,N_17429);
or U17585 (N_17585,N_17116,N_17346);
and U17586 (N_17586,N_17098,N_17071);
nor U17587 (N_17587,N_17440,N_17130);
nand U17588 (N_17588,N_17227,N_17471);
nand U17589 (N_17589,N_17456,N_17366);
nor U17590 (N_17590,N_17426,N_17173);
or U17591 (N_17591,N_17484,N_17408);
nand U17592 (N_17592,N_17220,N_17147);
xnor U17593 (N_17593,N_17089,N_17197);
xnor U17594 (N_17594,N_17167,N_17319);
nor U17595 (N_17595,N_17044,N_17270);
nand U17596 (N_17596,N_17052,N_17186);
xnor U17597 (N_17597,N_17039,N_17118);
or U17598 (N_17598,N_17158,N_17462);
xor U17599 (N_17599,N_17077,N_17412);
nor U17600 (N_17600,N_17473,N_17190);
nand U17601 (N_17601,N_17201,N_17248);
and U17602 (N_17602,N_17434,N_17066);
or U17603 (N_17603,N_17182,N_17357);
and U17604 (N_17604,N_17490,N_17059);
or U17605 (N_17605,N_17004,N_17083);
nand U17606 (N_17606,N_17058,N_17329);
nand U17607 (N_17607,N_17373,N_17466);
and U17608 (N_17608,N_17207,N_17386);
and U17609 (N_17609,N_17046,N_17278);
or U17610 (N_17610,N_17219,N_17316);
xor U17611 (N_17611,N_17447,N_17284);
nor U17612 (N_17612,N_17218,N_17403);
nand U17613 (N_17613,N_17475,N_17277);
nand U17614 (N_17614,N_17276,N_17464);
nand U17615 (N_17615,N_17413,N_17388);
nand U17616 (N_17616,N_17443,N_17144);
xnor U17617 (N_17617,N_17480,N_17430);
or U17618 (N_17618,N_17369,N_17279);
xnor U17619 (N_17619,N_17120,N_17100);
or U17620 (N_17620,N_17455,N_17170);
and U17621 (N_17621,N_17379,N_17016);
or U17622 (N_17622,N_17013,N_17358);
nor U17623 (N_17623,N_17380,N_17472);
and U17624 (N_17624,N_17204,N_17442);
nand U17625 (N_17625,N_17146,N_17115);
and U17626 (N_17626,N_17295,N_17001);
or U17627 (N_17627,N_17307,N_17164);
or U17628 (N_17628,N_17281,N_17132);
and U17629 (N_17629,N_17450,N_17206);
or U17630 (N_17630,N_17076,N_17153);
xnor U17631 (N_17631,N_17481,N_17065);
and U17632 (N_17632,N_17086,N_17154);
and U17633 (N_17633,N_17156,N_17326);
nand U17634 (N_17634,N_17495,N_17296);
nand U17635 (N_17635,N_17261,N_17037);
and U17636 (N_17636,N_17256,N_17230);
or U17637 (N_17637,N_17344,N_17102);
and U17638 (N_17638,N_17311,N_17101);
nand U17639 (N_17639,N_17057,N_17196);
nand U17640 (N_17640,N_17382,N_17215);
xnor U17641 (N_17641,N_17047,N_17445);
xor U17642 (N_17642,N_17117,N_17324);
nor U17643 (N_17643,N_17275,N_17069);
nor U17644 (N_17644,N_17235,N_17305);
or U17645 (N_17645,N_17499,N_17043);
or U17646 (N_17646,N_17418,N_17374);
nand U17647 (N_17647,N_17249,N_17309);
or U17648 (N_17648,N_17449,N_17269);
nor U17649 (N_17649,N_17290,N_17335);
xnor U17650 (N_17650,N_17211,N_17321);
nor U17651 (N_17651,N_17308,N_17397);
xor U17652 (N_17652,N_17461,N_17122);
nor U17653 (N_17653,N_17351,N_17387);
nor U17654 (N_17654,N_17331,N_17181);
nor U17655 (N_17655,N_17245,N_17232);
nand U17656 (N_17656,N_17162,N_17392);
or U17657 (N_17657,N_17129,N_17355);
xnor U17658 (N_17658,N_17428,N_17385);
and U17659 (N_17659,N_17012,N_17334);
nor U17660 (N_17660,N_17384,N_17310);
or U17661 (N_17661,N_17257,N_17423);
and U17662 (N_17662,N_17108,N_17068);
or U17663 (N_17663,N_17179,N_17026);
or U17664 (N_17664,N_17064,N_17312);
xnor U17665 (N_17665,N_17469,N_17213);
and U17666 (N_17666,N_17203,N_17395);
or U17667 (N_17667,N_17255,N_17151);
nor U17668 (N_17668,N_17010,N_17243);
nor U17669 (N_17669,N_17314,N_17400);
nand U17670 (N_17670,N_17242,N_17298);
or U17671 (N_17671,N_17079,N_17018);
and U17672 (N_17672,N_17056,N_17474);
xnor U17673 (N_17673,N_17091,N_17286);
nand U17674 (N_17674,N_17496,N_17107);
or U17675 (N_17675,N_17009,N_17332);
xnor U17676 (N_17676,N_17303,N_17095);
nor U17677 (N_17677,N_17262,N_17398);
nand U17678 (N_17678,N_17007,N_17159);
nand U17679 (N_17679,N_17160,N_17085);
and U17680 (N_17680,N_17337,N_17200);
xnor U17681 (N_17681,N_17172,N_17055);
nor U17682 (N_17682,N_17439,N_17133);
nand U17683 (N_17683,N_17054,N_17128);
nand U17684 (N_17684,N_17180,N_17208);
and U17685 (N_17685,N_17497,N_17414);
nand U17686 (N_17686,N_17293,N_17148);
nand U17687 (N_17687,N_17460,N_17032);
xor U17688 (N_17688,N_17033,N_17027);
xor U17689 (N_17689,N_17458,N_17210);
xor U17690 (N_17690,N_17259,N_17003);
or U17691 (N_17691,N_17322,N_17340);
nand U17692 (N_17692,N_17299,N_17313);
nand U17693 (N_17693,N_17150,N_17177);
or U17694 (N_17694,N_17416,N_17294);
or U17695 (N_17695,N_17217,N_17394);
and U17696 (N_17696,N_17078,N_17205);
and U17697 (N_17697,N_17081,N_17396);
and U17698 (N_17698,N_17417,N_17005);
nor U17699 (N_17699,N_17271,N_17236);
nand U17700 (N_17700,N_17370,N_17202);
or U17701 (N_17701,N_17390,N_17163);
and U17702 (N_17702,N_17244,N_17246);
or U17703 (N_17703,N_17020,N_17121);
and U17704 (N_17704,N_17488,N_17127);
nand U17705 (N_17705,N_17135,N_17389);
xor U17706 (N_17706,N_17082,N_17161);
and U17707 (N_17707,N_17000,N_17454);
nor U17708 (N_17708,N_17323,N_17233);
or U17709 (N_17709,N_17002,N_17014);
nor U17710 (N_17710,N_17364,N_17125);
xnor U17711 (N_17711,N_17401,N_17143);
nand U17712 (N_17712,N_17251,N_17343);
or U17713 (N_17713,N_17223,N_17011);
xor U17714 (N_17714,N_17300,N_17239);
nand U17715 (N_17715,N_17053,N_17487);
or U17716 (N_17716,N_17140,N_17134);
nand U17717 (N_17717,N_17419,N_17362);
nand U17718 (N_17718,N_17287,N_17139);
nor U17719 (N_17719,N_17250,N_17111);
and U17720 (N_17720,N_17241,N_17438);
and U17721 (N_17721,N_17157,N_17338);
or U17722 (N_17722,N_17228,N_17006);
and U17723 (N_17723,N_17124,N_17145);
or U17724 (N_17724,N_17040,N_17470);
or U17725 (N_17725,N_17050,N_17216);
or U17726 (N_17726,N_17266,N_17378);
nand U17727 (N_17727,N_17494,N_17291);
and U17728 (N_17728,N_17234,N_17137);
and U17729 (N_17729,N_17289,N_17025);
or U17730 (N_17730,N_17237,N_17350);
and U17731 (N_17731,N_17468,N_17030);
xor U17732 (N_17732,N_17391,N_17015);
or U17733 (N_17733,N_17254,N_17424);
or U17734 (N_17734,N_17405,N_17104);
nor U17735 (N_17735,N_17486,N_17330);
and U17736 (N_17736,N_17288,N_17222);
xor U17737 (N_17737,N_17049,N_17477);
nand U17738 (N_17738,N_17022,N_17377);
nand U17739 (N_17739,N_17347,N_17421);
and U17740 (N_17740,N_17399,N_17096);
nor U17741 (N_17741,N_17114,N_17017);
nor U17742 (N_17742,N_17031,N_17325);
and U17743 (N_17743,N_17359,N_17367);
and U17744 (N_17744,N_17060,N_17183);
nor U17745 (N_17745,N_17247,N_17436);
and U17746 (N_17746,N_17465,N_17353);
nor U17747 (N_17747,N_17444,N_17491);
nand U17748 (N_17748,N_17035,N_17045);
nand U17749 (N_17749,N_17339,N_17155);
and U17750 (N_17750,N_17357,N_17179);
nor U17751 (N_17751,N_17143,N_17389);
xnor U17752 (N_17752,N_17341,N_17026);
or U17753 (N_17753,N_17032,N_17325);
nor U17754 (N_17754,N_17172,N_17179);
or U17755 (N_17755,N_17118,N_17069);
nor U17756 (N_17756,N_17417,N_17196);
nor U17757 (N_17757,N_17337,N_17142);
nor U17758 (N_17758,N_17206,N_17435);
nand U17759 (N_17759,N_17357,N_17194);
and U17760 (N_17760,N_17406,N_17186);
or U17761 (N_17761,N_17061,N_17402);
xor U17762 (N_17762,N_17110,N_17132);
nand U17763 (N_17763,N_17233,N_17444);
and U17764 (N_17764,N_17045,N_17268);
and U17765 (N_17765,N_17236,N_17028);
xor U17766 (N_17766,N_17228,N_17017);
or U17767 (N_17767,N_17266,N_17385);
and U17768 (N_17768,N_17059,N_17243);
nor U17769 (N_17769,N_17161,N_17222);
and U17770 (N_17770,N_17248,N_17218);
xor U17771 (N_17771,N_17407,N_17197);
nor U17772 (N_17772,N_17219,N_17040);
nor U17773 (N_17773,N_17031,N_17243);
xnor U17774 (N_17774,N_17009,N_17293);
or U17775 (N_17775,N_17057,N_17377);
and U17776 (N_17776,N_17302,N_17148);
nor U17777 (N_17777,N_17290,N_17408);
nor U17778 (N_17778,N_17014,N_17075);
or U17779 (N_17779,N_17190,N_17409);
and U17780 (N_17780,N_17364,N_17068);
xnor U17781 (N_17781,N_17009,N_17071);
or U17782 (N_17782,N_17047,N_17335);
or U17783 (N_17783,N_17438,N_17207);
nor U17784 (N_17784,N_17039,N_17162);
xnor U17785 (N_17785,N_17098,N_17315);
or U17786 (N_17786,N_17047,N_17242);
xnor U17787 (N_17787,N_17284,N_17300);
xnor U17788 (N_17788,N_17050,N_17204);
xnor U17789 (N_17789,N_17468,N_17049);
nand U17790 (N_17790,N_17187,N_17274);
nand U17791 (N_17791,N_17250,N_17134);
nor U17792 (N_17792,N_17069,N_17053);
or U17793 (N_17793,N_17114,N_17447);
and U17794 (N_17794,N_17220,N_17106);
and U17795 (N_17795,N_17035,N_17443);
and U17796 (N_17796,N_17131,N_17438);
or U17797 (N_17797,N_17009,N_17498);
and U17798 (N_17798,N_17241,N_17369);
and U17799 (N_17799,N_17386,N_17000);
and U17800 (N_17800,N_17150,N_17038);
and U17801 (N_17801,N_17001,N_17179);
xnor U17802 (N_17802,N_17400,N_17197);
xor U17803 (N_17803,N_17163,N_17374);
nor U17804 (N_17804,N_17263,N_17359);
nand U17805 (N_17805,N_17026,N_17171);
xor U17806 (N_17806,N_17261,N_17307);
nor U17807 (N_17807,N_17310,N_17458);
nand U17808 (N_17808,N_17398,N_17052);
or U17809 (N_17809,N_17229,N_17414);
nor U17810 (N_17810,N_17194,N_17149);
xor U17811 (N_17811,N_17382,N_17267);
nor U17812 (N_17812,N_17039,N_17403);
nor U17813 (N_17813,N_17046,N_17360);
nand U17814 (N_17814,N_17434,N_17225);
nand U17815 (N_17815,N_17197,N_17298);
xnor U17816 (N_17816,N_17392,N_17134);
xnor U17817 (N_17817,N_17226,N_17278);
and U17818 (N_17818,N_17320,N_17285);
or U17819 (N_17819,N_17002,N_17334);
or U17820 (N_17820,N_17322,N_17475);
nand U17821 (N_17821,N_17020,N_17075);
nor U17822 (N_17822,N_17058,N_17245);
or U17823 (N_17823,N_17359,N_17048);
nor U17824 (N_17824,N_17280,N_17487);
xnor U17825 (N_17825,N_17070,N_17203);
xnor U17826 (N_17826,N_17146,N_17333);
nand U17827 (N_17827,N_17042,N_17084);
xnor U17828 (N_17828,N_17238,N_17488);
nand U17829 (N_17829,N_17070,N_17211);
nor U17830 (N_17830,N_17227,N_17195);
and U17831 (N_17831,N_17130,N_17052);
nor U17832 (N_17832,N_17276,N_17330);
or U17833 (N_17833,N_17181,N_17343);
nor U17834 (N_17834,N_17349,N_17209);
and U17835 (N_17835,N_17332,N_17192);
nand U17836 (N_17836,N_17358,N_17188);
or U17837 (N_17837,N_17234,N_17014);
nand U17838 (N_17838,N_17228,N_17149);
and U17839 (N_17839,N_17033,N_17301);
nand U17840 (N_17840,N_17196,N_17177);
nand U17841 (N_17841,N_17156,N_17039);
nor U17842 (N_17842,N_17242,N_17156);
or U17843 (N_17843,N_17043,N_17331);
or U17844 (N_17844,N_17058,N_17421);
and U17845 (N_17845,N_17166,N_17358);
or U17846 (N_17846,N_17273,N_17007);
or U17847 (N_17847,N_17282,N_17172);
nand U17848 (N_17848,N_17133,N_17076);
nor U17849 (N_17849,N_17419,N_17263);
nor U17850 (N_17850,N_17236,N_17115);
nand U17851 (N_17851,N_17422,N_17086);
and U17852 (N_17852,N_17333,N_17401);
nor U17853 (N_17853,N_17315,N_17101);
xor U17854 (N_17854,N_17460,N_17461);
nand U17855 (N_17855,N_17267,N_17291);
or U17856 (N_17856,N_17236,N_17466);
nor U17857 (N_17857,N_17278,N_17213);
or U17858 (N_17858,N_17262,N_17324);
nor U17859 (N_17859,N_17221,N_17012);
nor U17860 (N_17860,N_17127,N_17374);
xor U17861 (N_17861,N_17098,N_17263);
xnor U17862 (N_17862,N_17153,N_17088);
or U17863 (N_17863,N_17226,N_17088);
xor U17864 (N_17864,N_17357,N_17006);
xor U17865 (N_17865,N_17268,N_17289);
nor U17866 (N_17866,N_17094,N_17307);
and U17867 (N_17867,N_17324,N_17161);
and U17868 (N_17868,N_17068,N_17398);
or U17869 (N_17869,N_17405,N_17460);
or U17870 (N_17870,N_17209,N_17269);
nor U17871 (N_17871,N_17221,N_17241);
nand U17872 (N_17872,N_17374,N_17100);
or U17873 (N_17873,N_17175,N_17093);
or U17874 (N_17874,N_17090,N_17485);
nor U17875 (N_17875,N_17372,N_17384);
nor U17876 (N_17876,N_17414,N_17359);
xnor U17877 (N_17877,N_17007,N_17024);
xnor U17878 (N_17878,N_17315,N_17133);
nand U17879 (N_17879,N_17304,N_17067);
or U17880 (N_17880,N_17174,N_17393);
nand U17881 (N_17881,N_17148,N_17082);
and U17882 (N_17882,N_17373,N_17280);
or U17883 (N_17883,N_17044,N_17492);
nor U17884 (N_17884,N_17137,N_17426);
and U17885 (N_17885,N_17492,N_17082);
or U17886 (N_17886,N_17402,N_17091);
xor U17887 (N_17887,N_17449,N_17073);
nor U17888 (N_17888,N_17148,N_17344);
nand U17889 (N_17889,N_17116,N_17198);
nor U17890 (N_17890,N_17158,N_17460);
nor U17891 (N_17891,N_17013,N_17285);
xnor U17892 (N_17892,N_17110,N_17168);
nand U17893 (N_17893,N_17436,N_17498);
and U17894 (N_17894,N_17429,N_17025);
nor U17895 (N_17895,N_17234,N_17495);
nand U17896 (N_17896,N_17238,N_17323);
or U17897 (N_17897,N_17357,N_17302);
or U17898 (N_17898,N_17042,N_17416);
xnor U17899 (N_17899,N_17472,N_17095);
and U17900 (N_17900,N_17334,N_17323);
or U17901 (N_17901,N_17142,N_17005);
xor U17902 (N_17902,N_17275,N_17003);
xnor U17903 (N_17903,N_17473,N_17404);
nor U17904 (N_17904,N_17439,N_17465);
and U17905 (N_17905,N_17064,N_17458);
nand U17906 (N_17906,N_17374,N_17424);
nor U17907 (N_17907,N_17368,N_17479);
nand U17908 (N_17908,N_17007,N_17148);
nand U17909 (N_17909,N_17162,N_17359);
nor U17910 (N_17910,N_17283,N_17011);
xor U17911 (N_17911,N_17124,N_17348);
nor U17912 (N_17912,N_17484,N_17273);
or U17913 (N_17913,N_17105,N_17182);
nand U17914 (N_17914,N_17203,N_17044);
and U17915 (N_17915,N_17002,N_17465);
or U17916 (N_17916,N_17377,N_17386);
and U17917 (N_17917,N_17422,N_17382);
nor U17918 (N_17918,N_17114,N_17146);
nor U17919 (N_17919,N_17383,N_17210);
xor U17920 (N_17920,N_17316,N_17393);
and U17921 (N_17921,N_17111,N_17112);
and U17922 (N_17922,N_17364,N_17196);
nand U17923 (N_17923,N_17254,N_17395);
nor U17924 (N_17924,N_17475,N_17011);
xor U17925 (N_17925,N_17192,N_17414);
xor U17926 (N_17926,N_17239,N_17211);
xor U17927 (N_17927,N_17294,N_17481);
or U17928 (N_17928,N_17466,N_17083);
or U17929 (N_17929,N_17363,N_17428);
or U17930 (N_17930,N_17104,N_17023);
xor U17931 (N_17931,N_17452,N_17008);
nor U17932 (N_17932,N_17118,N_17062);
nand U17933 (N_17933,N_17206,N_17428);
or U17934 (N_17934,N_17272,N_17269);
xor U17935 (N_17935,N_17423,N_17343);
or U17936 (N_17936,N_17159,N_17371);
xor U17937 (N_17937,N_17363,N_17392);
nand U17938 (N_17938,N_17211,N_17241);
nand U17939 (N_17939,N_17098,N_17130);
nand U17940 (N_17940,N_17319,N_17386);
nand U17941 (N_17941,N_17331,N_17382);
nor U17942 (N_17942,N_17287,N_17261);
or U17943 (N_17943,N_17336,N_17218);
xnor U17944 (N_17944,N_17093,N_17411);
or U17945 (N_17945,N_17016,N_17097);
and U17946 (N_17946,N_17279,N_17285);
or U17947 (N_17947,N_17086,N_17072);
xor U17948 (N_17948,N_17021,N_17014);
nand U17949 (N_17949,N_17448,N_17288);
xor U17950 (N_17950,N_17125,N_17099);
xnor U17951 (N_17951,N_17242,N_17111);
nor U17952 (N_17952,N_17383,N_17469);
xor U17953 (N_17953,N_17228,N_17336);
nor U17954 (N_17954,N_17451,N_17342);
and U17955 (N_17955,N_17492,N_17397);
nand U17956 (N_17956,N_17244,N_17093);
or U17957 (N_17957,N_17264,N_17265);
and U17958 (N_17958,N_17022,N_17001);
nor U17959 (N_17959,N_17010,N_17078);
xnor U17960 (N_17960,N_17410,N_17222);
nand U17961 (N_17961,N_17020,N_17488);
xnor U17962 (N_17962,N_17405,N_17373);
and U17963 (N_17963,N_17111,N_17181);
nand U17964 (N_17964,N_17282,N_17289);
or U17965 (N_17965,N_17037,N_17182);
and U17966 (N_17966,N_17393,N_17053);
nand U17967 (N_17967,N_17242,N_17163);
and U17968 (N_17968,N_17166,N_17093);
nor U17969 (N_17969,N_17265,N_17328);
xnor U17970 (N_17970,N_17143,N_17317);
or U17971 (N_17971,N_17287,N_17114);
nand U17972 (N_17972,N_17486,N_17033);
and U17973 (N_17973,N_17241,N_17417);
xnor U17974 (N_17974,N_17053,N_17300);
or U17975 (N_17975,N_17159,N_17312);
nor U17976 (N_17976,N_17233,N_17131);
nand U17977 (N_17977,N_17159,N_17221);
nor U17978 (N_17978,N_17252,N_17027);
nand U17979 (N_17979,N_17216,N_17242);
xor U17980 (N_17980,N_17191,N_17387);
nand U17981 (N_17981,N_17193,N_17214);
or U17982 (N_17982,N_17036,N_17253);
xor U17983 (N_17983,N_17086,N_17467);
and U17984 (N_17984,N_17038,N_17195);
nand U17985 (N_17985,N_17103,N_17015);
or U17986 (N_17986,N_17331,N_17413);
or U17987 (N_17987,N_17258,N_17131);
or U17988 (N_17988,N_17055,N_17059);
nor U17989 (N_17989,N_17340,N_17153);
nand U17990 (N_17990,N_17360,N_17100);
nand U17991 (N_17991,N_17356,N_17188);
nor U17992 (N_17992,N_17118,N_17303);
or U17993 (N_17993,N_17293,N_17227);
nor U17994 (N_17994,N_17262,N_17034);
or U17995 (N_17995,N_17143,N_17466);
nand U17996 (N_17996,N_17134,N_17229);
nor U17997 (N_17997,N_17492,N_17096);
or U17998 (N_17998,N_17061,N_17062);
xor U17999 (N_17999,N_17130,N_17107);
xnor U18000 (N_18000,N_17853,N_17925);
and U18001 (N_18001,N_17604,N_17780);
and U18002 (N_18002,N_17718,N_17987);
or U18003 (N_18003,N_17740,N_17803);
xor U18004 (N_18004,N_17659,N_17969);
and U18005 (N_18005,N_17896,N_17614);
nor U18006 (N_18006,N_17817,N_17993);
nor U18007 (N_18007,N_17598,N_17952);
or U18008 (N_18008,N_17919,N_17643);
and U18009 (N_18009,N_17678,N_17544);
nand U18010 (N_18010,N_17961,N_17635);
or U18011 (N_18011,N_17512,N_17907);
nand U18012 (N_18012,N_17697,N_17707);
and U18013 (N_18013,N_17564,N_17885);
and U18014 (N_18014,N_17912,N_17596);
nand U18015 (N_18015,N_17641,N_17540);
xor U18016 (N_18016,N_17599,N_17752);
nand U18017 (N_18017,N_17537,N_17768);
xnor U18018 (N_18018,N_17877,N_17534);
or U18019 (N_18019,N_17954,N_17837);
xnor U18020 (N_18020,N_17711,N_17523);
and U18021 (N_18021,N_17839,N_17840);
and U18022 (N_18022,N_17737,N_17557);
or U18023 (N_18023,N_17589,N_17791);
nor U18024 (N_18024,N_17778,N_17661);
or U18025 (N_18025,N_17953,N_17744);
and U18026 (N_18026,N_17600,N_17841);
nand U18027 (N_18027,N_17974,N_17730);
and U18028 (N_18028,N_17522,N_17668);
nor U18029 (N_18029,N_17725,N_17995);
or U18030 (N_18030,N_17623,N_17856);
nor U18031 (N_18031,N_17767,N_17874);
and U18032 (N_18032,N_17642,N_17597);
xor U18033 (N_18033,N_17875,N_17982);
or U18034 (N_18034,N_17656,N_17543);
nor U18035 (N_18035,N_17942,N_17784);
nand U18036 (N_18036,N_17763,N_17850);
xnor U18037 (N_18037,N_17601,N_17801);
nor U18038 (N_18038,N_17572,N_17943);
nor U18039 (N_18039,N_17783,N_17647);
nor U18040 (N_18040,N_17858,N_17750);
and U18041 (N_18041,N_17658,N_17886);
nor U18042 (N_18042,N_17944,N_17525);
xor U18043 (N_18043,N_17805,N_17680);
or U18044 (N_18044,N_17923,N_17503);
and U18045 (N_18045,N_17786,N_17696);
and U18046 (N_18046,N_17665,N_17866);
and U18047 (N_18047,N_17619,N_17533);
nand U18048 (N_18048,N_17980,N_17552);
or U18049 (N_18049,N_17712,N_17613);
and U18050 (N_18050,N_17899,N_17547);
nand U18051 (N_18051,N_17646,N_17683);
nand U18052 (N_18052,N_17810,N_17594);
or U18053 (N_18053,N_17922,N_17908);
or U18054 (N_18054,N_17688,N_17500);
or U18055 (N_18055,N_17566,N_17978);
or U18056 (N_18056,N_17797,N_17950);
nor U18057 (N_18057,N_17951,N_17505);
nand U18058 (N_18058,N_17719,N_17675);
nor U18059 (N_18059,N_17649,N_17935);
nand U18060 (N_18060,N_17981,N_17798);
nand U18061 (N_18061,N_17677,N_17959);
xor U18062 (N_18062,N_17838,N_17531);
nand U18063 (N_18063,N_17667,N_17548);
nand U18064 (N_18064,N_17824,N_17945);
nand U18065 (N_18065,N_17804,N_17782);
nand U18066 (N_18066,N_17749,N_17536);
and U18067 (N_18067,N_17618,N_17616);
nand U18068 (N_18068,N_17869,N_17507);
xor U18069 (N_18069,N_17990,N_17622);
and U18070 (N_18070,N_17878,N_17873);
and U18071 (N_18071,N_17577,N_17754);
nor U18072 (N_18072,N_17852,N_17814);
or U18073 (N_18073,N_17829,N_17705);
nor U18074 (N_18074,N_17765,N_17602);
xnor U18075 (N_18075,N_17893,N_17862);
nor U18076 (N_18076,N_17631,N_17693);
nor U18077 (N_18077,N_17881,N_17578);
nor U18078 (N_18078,N_17930,N_17563);
and U18079 (N_18079,N_17895,N_17773);
or U18080 (N_18080,N_17679,N_17836);
and U18081 (N_18081,N_17813,N_17884);
xnor U18082 (N_18082,N_17913,N_17670);
and U18083 (N_18083,N_17800,N_17511);
xor U18084 (N_18084,N_17528,N_17891);
nor U18085 (N_18085,N_17920,N_17686);
nand U18086 (N_18086,N_17615,N_17867);
or U18087 (N_18087,N_17892,N_17807);
xnor U18088 (N_18088,N_17915,N_17519);
and U18089 (N_18089,N_17603,N_17651);
or U18090 (N_18090,N_17702,N_17992);
or U18091 (N_18091,N_17558,N_17710);
nor U18092 (N_18092,N_17785,N_17876);
nor U18093 (N_18093,N_17671,N_17593);
nand U18094 (N_18094,N_17806,N_17632);
xnor U18095 (N_18095,N_17729,N_17743);
xnor U18096 (N_18096,N_17762,N_17723);
or U18097 (N_18097,N_17742,N_17538);
nand U18098 (N_18098,N_17976,N_17914);
and U18099 (N_18099,N_17666,N_17588);
nor U18100 (N_18100,N_17595,N_17772);
xnor U18101 (N_18101,N_17720,N_17608);
xor U18102 (N_18102,N_17989,N_17764);
and U18103 (N_18103,N_17706,N_17660);
or U18104 (N_18104,N_17859,N_17606);
and U18105 (N_18105,N_17605,N_17916);
and U18106 (N_18106,N_17554,N_17997);
xor U18107 (N_18107,N_17849,N_17934);
and U18108 (N_18108,N_17940,N_17819);
nand U18109 (N_18109,N_17633,N_17747);
and U18110 (N_18110,N_17575,N_17518);
xor U18111 (N_18111,N_17714,N_17818);
and U18112 (N_18112,N_17816,N_17621);
nand U18113 (N_18113,N_17956,N_17777);
xor U18114 (N_18114,N_17774,N_17610);
nor U18115 (N_18115,N_17701,N_17713);
and U18116 (N_18116,N_17921,N_17863);
and U18117 (N_18117,N_17584,N_17590);
xnor U18118 (N_18118,N_17520,N_17811);
and U18119 (N_18119,N_17898,N_17626);
xor U18120 (N_18120,N_17830,N_17929);
nor U18121 (N_18121,N_17662,N_17581);
nand U18122 (N_18122,N_17851,N_17553);
nand U18123 (N_18123,N_17684,N_17620);
nand U18124 (N_18124,N_17574,N_17761);
nor U18125 (N_18125,N_17627,N_17527);
nand U18126 (N_18126,N_17648,N_17900);
and U18127 (N_18127,N_17630,N_17735);
nand U18128 (N_18128,N_17928,N_17909);
nand U18129 (N_18129,N_17789,N_17689);
or U18130 (N_18130,N_17732,N_17793);
nand U18131 (N_18131,N_17924,N_17906);
or U18132 (N_18132,N_17695,N_17672);
nand U18133 (N_18133,N_17530,N_17741);
or U18134 (N_18134,N_17650,N_17551);
xor U18135 (N_18135,N_17794,N_17644);
xor U18136 (N_18136,N_17988,N_17673);
nand U18137 (N_18137,N_17510,N_17694);
and U18138 (N_18138,N_17733,N_17625);
or U18139 (N_18139,N_17999,N_17766);
xor U18140 (N_18140,N_17795,N_17539);
nand U18141 (N_18141,N_17911,N_17901);
nor U18142 (N_18142,N_17526,N_17687);
xnor U18143 (N_18143,N_17700,N_17790);
nand U18144 (N_18144,N_17704,N_17991);
nor U18145 (N_18145,N_17939,N_17550);
xnor U18146 (N_18146,N_17573,N_17815);
and U18147 (N_18147,N_17502,N_17796);
nand U18148 (N_18148,N_17822,N_17624);
and U18149 (N_18149,N_17760,N_17638);
nor U18150 (N_18150,N_17775,N_17826);
or U18151 (N_18151,N_17835,N_17676);
or U18152 (N_18152,N_17515,N_17521);
nand U18153 (N_18153,N_17889,N_17664);
xor U18154 (N_18154,N_17965,N_17975);
or U18155 (N_18155,N_17580,N_17998);
nand U18156 (N_18156,N_17709,N_17871);
nor U18157 (N_18157,N_17726,N_17971);
xnor U18158 (N_18158,N_17986,N_17514);
nor U18159 (N_18159,N_17788,N_17917);
nand U18160 (N_18160,N_17792,N_17758);
and U18161 (N_18161,N_17946,N_17504);
or U18162 (N_18162,N_17821,N_17808);
or U18163 (N_18163,N_17966,N_17846);
nand U18164 (N_18164,N_17745,N_17739);
and U18165 (N_18165,N_17565,N_17787);
xnor U18166 (N_18166,N_17653,N_17727);
or U18167 (N_18167,N_17654,N_17827);
and U18168 (N_18168,N_17634,N_17517);
and U18169 (N_18169,N_17967,N_17870);
and U18170 (N_18170,N_17825,N_17972);
or U18171 (N_18171,N_17560,N_17532);
xor U18172 (N_18172,N_17834,N_17663);
nor U18173 (N_18173,N_17591,N_17576);
nand U18174 (N_18174,N_17949,N_17958);
nand U18175 (N_18175,N_17582,N_17716);
or U18176 (N_18176,N_17910,N_17535);
nor U18177 (N_18177,N_17887,N_17880);
nand U18178 (N_18178,N_17570,N_17569);
or U18179 (N_18179,N_17562,N_17857);
xnor U18180 (N_18180,N_17657,N_17984);
nor U18181 (N_18181,N_17546,N_17931);
nand U18182 (N_18182,N_17579,N_17549);
nor U18183 (N_18183,N_17926,N_17844);
and U18184 (N_18184,N_17894,N_17905);
xnor U18185 (N_18185,N_17541,N_17831);
nand U18186 (N_18186,N_17904,N_17524);
nand U18187 (N_18187,N_17639,N_17506);
nor U18188 (N_18188,N_17755,N_17759);
and U18189 (N_18189,N_17842,N_17607);
nand U18190 (N_18190,N_17865,N_17698);
or U18191 (N_18191,N_17985,N_17757);
nand U18192 (N_18192,N_17513,N_17724);
nand U18193 (N_18193,N_17864,N_17937);
xor U18194 (N_18194,N_17746,N_17854);
nand U18195 (N_18195,N_17902,N_17996);
xor U18196 (N_18196,N_17652,N_17820);
nand U18197 (N_18197,N_17681,N_17964);
nor U18198 (N_18198,N_17731,N_17957);
nor U18199 (N_18199,N_17722,N_17751);
nor U18200 (N_18200,N_17936,N_17776);
nor U18201 (N_18201,N_17941,N_17612);
nand U18202 (N_18202,N_17636,N_17708);
nor U18203 (N_18203,N_17640,N_17611);
xor U18204 (N_18204,N_17674,N_17833);
and U18205 (N_18205,N_17609,N_17888);
or U18206 (N_18206,N_17559,N_17756);
xnor U18207 (N_18207,N_17699,N_17948);
xor U18208 (N_18208,N_17529,N_17872);
or U18209 (N_18209,N_17586,N_17637);
and U18210 (N_18210,N_17848,N_17545);
nand U18211 (N_18211,N_17861,N_17715);
or U18212 (N_18212,N_17736,N_17728);
or U18213 (N_18213,N_17933,N_17703);
xor U18214 (N_18214,N_17960,N_17682);
nor U18215 (N_18215,N_17883,N_17721);
and U18216 (N_18216,N_17781,N_17809);
nor U18217 (N_18217,N_17962,N_17583);
and U18218 (N_18218,N_17955,N_17977);
nand U18219 (N_18219,N_17812,N_17973);
or U18220 (N_18220,N_17903,N_17645);
xnor U18221 (N_18221,N_17868,N_17947);
nor U18222 (N_18222,N_17556,N_17769);
and U18223 (N_18223,N_17979,N_17685);
nand U18224 (N_18224,N_17617,N_17832);
xnor U18225 (N_18225,N_17779,N_17802);
xor U18226 (N_18226,N_17629,N_17845);
nor U18227 (N_18227,N_17748,N_17897);
nand U18228 (N_18228,N_17669,N_17555);
and U18229 (N_18229,N_17994,N_17717);
and U18230 (N_18230,N_17932,N_17542);
or U18231 (N_18231,N_17799,N_17860);
nand U18232 (N_18232,N_17501,N_17567);
nand U18233 (N_18233,N_17738,N_17753);
xor U18234 (N_18234,N_17568,N_17509);
xnor U18235 (N_18235,N_17879,N_17734);
and U18236 (N_18236,N_17938,N_17561);
nor U18237 (N_18237,N_17585,N_17970);
nand U18238 (N_18238,N_17628,N_17968);
and U18239 (N_18239,N_17508,N_17847);
nand U18240 (N_18240,N_17927,N_17770);
xor U18241 (N_18241,N_17691,N_17828);
and U18242 (N_18242,N_17571,N_17963);
nand U18243 (N_18243,N_17890,N_17655);
or U18244 (N_18244,N_17823,N_17587);
nor U18245 (N_18245,N_17690,N_17516);
or U18246 (N_18246,N_17843,N_17983);
nor U18247 (N_18247,N_17918,N_17882);
nor U18248 (N_18248,N_17855,N_17692);
or U18249 (N_18249,N_17771,N_17592);
or U18250 (N_18250,N_17986,N_17922);
nor U18251 (N_18251,N_17978,N_17786);
or U18252 (N_18252,N_17609,N_17647);
and U18253 (N_18253,N_17647,N_17545);
and U18254 (N_18254,N_17686,N_17698);
xnor U18255 (N_18255,N_17925,N_17914);
and U18256 (N_18256,N_17666,N_17612);
or U18257 (N_18257,N_17707,N_17590);
xor U18258 (N_18258,N_17982,N_17996);
and U18259 (N_18259,N_17886,N_17783);
or U18260 (N_18260,N_17650,N_17778);
or U18261 (N_18261,N_17639,N_17995);
nand U18262 (N_18262,N_17834,N_17753);
xor U18263 (N_18263,N_17566,N_17792);
nor U18264 (N_18264,N_17986,N_17990);
nor U18265 (N_18265,N_17500,N_17722);
or U18266 (N_18266,N_17791,N_17886);
and U18267 (N_18267,N_17621,N_17735);
nand U18268 (N_18268,N_17888,N_17859);
xnor U18269 (N_18269,N_17509,N_17901);
or U18270 (N_18270,N_17981,N_17891);
nand U18271 (N_18271,N_17957,N_17670);
nand U18272 (N_18272,N_17742,N_17899);
nor U18273 (N_18273,N_17767,N_17745);
or U18274 (N_18274,N_17695,N_17654);
or U18275 (N_18275,N_17726,N_17534);
nand U18276 (N_18276,N_17657,N_17512);
nand U18277 (N_18277,N_17610,N_17779);
or U18278 (N_18278,N_17564,N_17784);
xor U18279 (N_18279,N_17722,N_17777);
nor U18280 (N_18280,N_17567,N_17648);
or U18281 (N_18281,N_17698,N_17893);
and U18282 (N_18282,N_17515,N_17765);
and U18283 (N_18283,N_17721,N_17501);
nand U18284 (N_18284,N_17972,N_17841);
and U18285 (N_18285,N_17781,N_17709);
xor U18286 (N_18286,N_17578,N_17878);
and U18287 (N_18287,N_17971,N_17981);
and U18288 (N_18288,N_17870,N_17696);
and U18289 (N_18289,N_17786,N_17573);
nor U18290 (N_18290,N_17608,N_17565);
xnor U18291 (N_18291,N_17920,N_17872);
nor U18292 (N_18292,N_17799,N_17763);
nand U18293 (N_18293,N_17828,N_17728);
xnor U18294 (N_18294,N_17515,N_17668);
xor U18295 (N_18295,N_17747,N_17906);
or U18296 (N_18296,N_17992,N_17558);
or U18297 (N_18297,N_17743,N_17876);
or U18298 (N_18298,N_17532,N_17828);
or U18299 (N_18299,N_17533,N_17632);
nand U18300 (N_18300,N_17838,N_17965);
xor U18301 (N_18301,N_17576,N_17522);
or U18302 (N_18302,N_17995,N_17547);
nand U18303 (N_18303,N_17909,N_17535);
or U18304 (N_18304,N_17529,N_17804);
or U18305 (N_18305,N_17500,N_17879);
and U18306 (N_18306,N_17970,N_17539);
or U18307 (N_18307,N_17539,N_17936);
xor U18308 (N_18308,N_17987,N_17697);
and U18309 (N_18309,N_17982,N_17603);
and U18310 (N_18310,N_17750,N_17623);
xnor U18311 (N_18311,N_17841,N_17879);
nand U18312 (N_18312,N_17748,N_17673);
xnor U18313 (N_18313,N_17652,N_17684);
or U18314 (N_18314,N_17567,N_17919);
nand U18315 (N_18315,N_17973,N_17703);
nand U18316 (N_18316,N_17519,N_17526);
and U18317 (N_18317,N_17729,N_17823);
or U18318 (N_18318,N_17722,N_17615);
xnor U18319 (N_18319,N_17813,N_17534);
xnor U18320 (N_18320,N_17815,N_17830);
nor U18321 (N_18321,N_17681,N_17736);
or U18322 (N_18322,N_17962,N_17714);
xor U18323 (N_18323,N_17697,N_17618);
or U18324 (N_18324,N_17726,N_17688);
and U18325 (N_18325,N_17634,N_17912);
nand U18326 (N_18326,N_17972,N_17828);
and U18327 (N_18327,N_17970,N_17671);
and U18328 (N_18328,N_17511,N_17978);
xor U18329 (N_18329,N_17646,N_17919);
xnor U18330 (N_18330,N_17546,N_17683);
and U18331 (N_18331,N_17816,N_17917);
and U18332 (N_18332,N_17919,N_17767);
nor U18333 (N_18333,N_17770,N_17565);
nor U18334 (N_18334,N_17588,N_17783);
nor U18335 (N_18335,N_17799,N_17834);
xor U18336 (N_18336,N_17743,N_17773);
and U18337 (N_18337,N_17516,N_17907);
and U18338 (N_18338,N_17676,N_17565);
nor U18339 (N_18339,N_17630,N_17539);
or U18340 (N_18340,N_17581,N_17718);
or U18341 (N_18341,N_17745,N_17990);
xnor U18342 (N_18342,N_17778,N_17826);
nor U18343 (N_18343,N_17995,N_17663);
nand U18344 (N_18344,N_17890,N_17805);
nor U18345 (N_18345,N_17921,N_17636);
or U18346 (N_18346,N_17827,N_17778);
xor U18347 (N_18347,N_17835,N_17532);
and U18348 (N_18348,N_17768,N_17642);
nor U18349 (N_18349,N_17690,N_17528);
or U18350 (N_18350,N_17831,N_17867);
and U18351 (N_18351,N_17982,N_17991);
xnor U18352 (N_18352,N_17629,N_17919);
xnor U18353 (N_18353,N_17855,N_17557);
nor U18354 (N_18354,N_17872,N_17770);
xnor U18355 (N_18355,N_17927,N_17996);
or U18356 (N_18356,N_17927,N_17966);
or U18357 (N_18357,N_17883,N_17601);
and U18358 (N_18358,N_17726,N_17887);
and U18359 (N_18359,N_17528,N_17799);
or U18360 (N_18360,N_17564,N_17873);
or U18361 (N_18361,N_17899,N_17975);
or U18362 (N_18362,N_17540,N_17505);
nand U18363 (N_18363,N_17506,N_17805);
xnor U18364 (N_18364,N_17630,N_17804);
nor U18365 (N_18365,N_17597,N_17681);
nand U18366 (N_18366,N_17963,N_17895);
xnor U18367 (N_18367,N_17856,N_17513);
xnor U18368 (N_18368,N_17771,N_17956);
nor U18369 (N_18369,N_17863,N_17681);
and U18370 (N_18370,N_17807,N_17616);
xnor U18371 (N_18371,N_17638,N_17627);
or U18372 (N_18372,N_17704,N_17827);
nand U18373 (N_18373,N_17518,N_17729);
or U18374 (N_18374,N_17842,N_17533);
and U18375 (N_18375,N_17994,N_17522);
or U18376 (N_18376,N_17853,N_17793);
or U18377 (N_18377,N_17814,N_17561);
nor U18378 (N_18378,N_17994,N_17846);
nor U18379 (N_18379,N_17832,N_17695);
nand U18380 (N_18380,N_17527,N_17730);
xor U18381 (N_18381,N_17773,N_17794);
and U18382 (N_18382,N_17627,N_17508);
or U18383 (N_18383,N_17767,N_17669);
xor U18384 (N_18384,N_17520,N_17706);
xor U18385 (N_18385,N_17629,N_17756);
nor U18386 (N_18386,N_17549,N_17903);
or U18387 (N_18387,N_17600,N_17787);
nor U18388 (N_18388,N_17617,N_17817);
nand U18389 (N_18389,N_17758,N_17615);
nand U18390 (N_18390,N_17736,N_17962);
nand U18391 (N_18391,N_17932,N_17547);
xnor U18392 (N_18392,N_17879,N_17872);
nor U18393 (N_18393,N_17676,N_17875);
nand U18394 (N_18394,N_17598,N_17918);
xnor U18395 (N_18395,N_17589,N_17518);
nand U18396 (N_18396,N_17666,N_17551);
and U18397 (N_18397,N_17794,N_17590);
nand U18398 (N_18398,N_17575,N_17975);
nor U18399 (N_18399,N_17749,N_17932);
or U18400 (N_18400,N_17695,N_17702);
xnor U18401 (N_18401,N_17642,N_17666);
or U18402 (N_18402,N_17910,N_17816);
or U18403 (N_18403,N_17694,N_17763);
and U18404 (N_18404,N_17714,N_17802);
and U18405 (N_18405,N_17999,N_17907);
xor U18406 (N_18406,N_17507,N_17885);
nand U18407 (N_18407,N_17644,N_17831);
xor U18408 (N_18408,N_17501,N_17857);
xnor U18409 (N_18409,N_17851,N_17823);
and U18410 (N_18410,N_17598,N_17618);
xnor U18411 (N_18411,N_17767,N_17613);
nor U18412 (N_18412,N_17827,N_17939);
xnor U18413 (N_18413,N_17682,N_17735);
or U18414 (N_18414,N_17591,N_17987);
nor U18415 (N_18415,N_17612,N_17712);
xnor U18416 (N_18416,N_17961,N_17670);
and U18417 (N_18417,N_17846,N_17507);
or U18418 (N_18418,N_17715,N_17708);
nor U18419 (N_18419,N_17714,N_17879);
nand U18420 (N_18420,N_17641,N_17589);
or U18421 (N_18421,N_17854,N_17864);
xor U18422 (N_18422,N_17797,N_17850);
and U18423 (N_18423,N_17960,N_17731);
xnor U18424 (N_18424,N_17519,N_17695);
xor U18425 (N_18425,N_17963,N_17906);
xnor U18426 (N_18426,N_17833,N_17720);
xor U18427 (N_18427,N_17937,N_17760);
xnor U18428 (N_18428,N_17824,N_17978);
nand U18429 (N_18429,N_17955,N_17575);
nor U18430 (N_18430,N_17500,N_17848);
xnor U18431 (N_18431,N_17553,N_17784);
xnor U18432 (N_18432,N_17792,N_17504);
and U18433 (N_18433,N_17921,N_17994);
or U18434 (N_18434,N_17772,N_17581);
nor U18435 (N_18435,N_17870,N_17800);
or U18436 (N_18436,N_17754,N_17602);
xor U18437 (N_18437,N_17862,N_17822);
xnor U18438 (N_18438,N_17673,N_17578);
xor U18439 (N_18439,N_17811,N_17954);
and U18440 (N_18440,N_17774,N_17746);
nor U18441 (N_18441,N_17951,N_17716);
nand U18442 (N_18442,N_17805,N_17889);
nand U18443 (N_18443,N_17775,N_17787);
and U18444 (N_18444,N_17890,N_17698);
and U18445 (N_18445,N_17721,N_17938);
nand U18446 (N_18446,N_17908,N_17801);
and U18447 (N_18447,N_17549,N_17938);
or U18448 (N_18448,N_17837,N_17842);
nand U18449 (N_18449,N_17730,N_17979);
and U18450 (N_18450,N_17658,N_17879);
xnor U18451 (N_18451,N_17701,N_17779);
nor U18452 (N_18452,N_17636,N_17742);
nor U18453 (N_18453,N_17900,N_17558);
xor U18454 (N_18454,N_17779,N_17899);
or U18455 (N_18455,N_17758,N_17830);
nor U18456 (N_18456,N_17648,N_17587);
nor U18457 (N_18457,N_17805,N_17601);
or U18458 (N_18458,N_17862,N_17948);
and U18459 (N_18459,N_17860,N_17851);
xor U18460 (N_18460,N_17750,N_17635);
xnor U18461 (N_18461,N_17909,N_17876);
or U18462 (N_18462,N_17626,N_17800);
and U18463 (N_18463,N_17505,N_17549);
nand U18464 (N_18464,N_17744,N_17540);
nor U18465 (N_18465,N_17834,N_17747);
xnor U18466 (N_18466,N_17657,N_17741);
xor U18467 (N_18467,N_17754,N_17541);
and U18468 (N_18468,N_17750,N_17856);
nand U18469 (N_18469,N_17950,N_17817);
xor U18470 (N_18470,N_17541,N_17769);
nor U18471 (N_18471,N_17756,N_17788);
nor U18472 (N_18472,N_17616,N_17805);
xnor U18473 (N_18473,N_17902,N_17520);
xor U18474 (N_18474,N_17642,N_17581);
xor U18475 (N_18475,N_17998,N_17563);
and U18476 (N_18476,N_17680,N_17954);
nand U18477 (N_18477,N_17899,N_17957);
nor U18478 (N_18478,N_17714,N_17798);
and U18479 (N_18479,N_17867,N_17516);
nor U18480 (N_18480,N_17550,N_17622);
and U18481 (N_18481,N_17544,N_17530);
xor U18482 (N_18482,N_17703,N_17691);
nor U18483 (N_18483,N_17655,N_17545);
nor U18484 (N_18484,N_17636,N_17561);
nand U18485 (N_18485,N_17542,N_17863);
and U18486 (N_18486,N_17805,N_17988);
and U18487 (N_18487,N_17577,N_17881);
xor U18488 (N_18488,N_17915,N_17698);
or U18489 (N_18489,N_17925,N_17953);
xnor U18490 (N_18490,N_17732,N_17926);
xor U18491 (N_18491,N_17710,N_17722);
nor U18492 (N_18492,N_17523,N_17624);
or U18493 (N_18493,N_17613,N_17756);
xnor U18494 (N_18494,N_17675,N_17918);
xnor U18495 (N_18495,N_17612,N_17972);
nand U18496 (N_18496,N_17504,N_17544);
nand U18497 (N_18497,N_17583,N_17638);
xnor U18498 (N_18498,N_17929,N_17925);
xnor U18499 (N_18499,N_17681,N_17663);
and U18500 (N_18500,N_18291,N_18362);
nand U18501 (N_18501,N_18243,N_18131);
xor U18502 (N_18502,N_18135,N_18448);
nor U18503 (N_18503,N_18493,N_18492);
nor U18504 (N_18504,N_18400,N_18441);
and U18505 (N_18505,N_18123,N_18399);
nand U18506 (N_18506,N_18267,N_18407);
nor U18507 (N_18507,N_18372,N_18459);
nor U18508 (N_18508,N_18042,N_18292);
nor U18509 (N_18509,N_18254,N_18195);
xor U18510 (N_18510,N_18252,N_18197);
or U18511 (N_18511,N_18040,N_18280);
nor U18512 (N_18512,N_18415,N_18025);
xor U18513 (N_18513,N_18029,N_18333);
nand U18514 (N_18514,N_18468,N_18274);
nand U18515 (N_18515,N_18159,N_18289);
nand U18516 (N_18516,N_18421,N_18263);
and U18517 (N_18517,N_18390,N_18442);
and U18518 (N_18518,N_18122,N_18199);
or U18519 (N_18519,N_18181,N_18084);
or U18520 (N_18520,N_18149,N_18455);
nor U18521 (N_18521,N_18337,N_18321);
nor U18522 (N_18522,N_18300,N_18111);
nor U18523 (N_18523,N_18478,N_18107);
or U18524 (N_18524,N_18353,N_18250);
or U18525 (N_18525,N_18093,N_18170);
or U18526 (N_18526,N_18268,N_18313);
xnor U18527 (N_18527,N_18347,N_18085);
xor U18528 (N_18528,N_18124,N_18251);
nor U18529 (N_18529,N_18154,N_18392);
nand U18530 (N_18530,N_18299,N_18298);
and U18531 (N_18531,N_18011,N_18158);
or U18532 (N_18532,N_18435,N_18414);
and U18533 (N_18533,N_18237,N_18189);
or U18534 (N_18534,N_18073,N_18401);
and U18535 (N_18535,N_18219,N_18469);
xor U18536 (N_18536,N_18242,N_18036);
nand U18537 (N_18537,N_18235,N_18050);
nor U18538 (N_18538,N_18222,N_18059);
nor U18539 (N_18539,N_18419,N_18352);
xor U18540 (N_18540,N_18256,N_18008);
and U18541 (N_18541,N_18041,N_18273);
or U18542 (N_18542,N_18006,N_18115);
xnor U18543 (N_18543,N_18003,N_18130);
and U18544 (N_18544,N_18338,N_18460);
nor U18545 (N_18545,N_18413,N_18488);
nor U18546 (N_18546,N_18214,N_18479);
and U18547 (N_18547,N_18015,N_18046);
nor U18548 (N_18548,N_18125,N_18438);
xnor U18549 (N_18549,N_18241,N_18229);
nand U18550 (N_18550,N_18100,N_18369);
or U18551 (N_18551,N_18329,N_18183);
xnor U18552 (N_18552,N_18444,N_18010);
nor U18553 (N_18553,N_18112,N_18301);
nor U18554 (N_18554,N_18339,N_18191);
or U18555 (N_18555,N_18344,N_18016);
nor U18556 (N_18556,N_18490,N_18176);
and U18557 (N_18557,N_18416,N_18496);
xor U18558 (N_18558,N_18173,N_18379);
nor U18559 (N_18559,N_18223,N_18001);
nor U18560 (N_18560,N_18366,N_18216);
nand U18561 (N_18561,N_18266,N_18447);
xor U18562 (N_18562,N_18172,N_18395);
and U18563 (N_18563,N_18230,N_18099);
nand U18564 (N_18564,N_18092,N_18062);
nand U18565 (N_18565,N_18018,N_18087);
nor U18566 (N_18566,N_18169,N_18026);
nor U18567 (N_18567,N_18163,N_18226);
nand U18568 (N_18568,N_18127,N_18168);
nand U18569 (N_18569,N_18198,N_18342);
xnor U18570 (N_18570,N_18367,N_18389);
xnor U18571 (N_18571,N_18343,N_18286);
xor U18572 (N_18572,N_18386,N_18458);
and U18573 (N_18573,N_18307,N_18045);
and U18574 (N_18574,N_18151,N_18283);
or U18575 (N_18575,N_18089,N_18261);
xor U18576 (N_18576,N_18102,N_18248);
xnor U18577 (N_18577,N_18153,N_18128);
nor U18578 (N_18578,N_18175,N_18023);
nor U18579 (N_18579,N_18466,N_18311);
and U18580 (N_18580,N_18494,N_18411);
nand U18581 (N_18581,N_18449,N_18218);
and U18582 (N_18582,N_18306,N_18231);
nor U18583 (N_18583,N_18161,N_18303);
and U18584 (N_18584,N_18262,N_18146);
nand U18585 (N_18585,N_18383,N_18038);
nand U18586 (N_18586,N_18418,N_18208);
nand U18587 (N_18587,N_18020,N_18304);
nand U18588 (N_18588,N_18033,N_18009);
nand U18589 (N_18589,N_18108,N_18326);
nand U18590 (N_18590,N_18247,N_18225);
xnor U18591 (N_18591,N_18368,N_18355);
nand U18592 (N_18592,N_18323,N_18239);
and U18593 (N_18593,N_18270,N_18017);
and U18594 (N_18594,N_18117,N_18082);
or U18595 (N_18595,N_18190,N_18489);
xnor U18596 (N_18596,N_18483,N_18005);
or U18597 (N_18597,N_18004,N_18354);
nand U18598 (N_18598,N_18378,N_18098);
xnor U18599 (N_18599,N_18457,N_18477);
nand U18600 (N_18600,N_18373,N_18302);
xor U18601 (N_18601,N_18287,N_18088);
and U18602 (N_18602,N_18480,N_18473);
or U18603 (N_18603,N_18186,N_18269);
nor U18604 (N_18604,N_18398,N_18325);
or U18605 (N_18605,N_18079,N_18077);
xnor U18606 (N_18606,N_18179,N_18486);
nor U18607 (N_18607,N_18019,N_18155);
xor U18608 (N_18608,N_18257,N_18030);
nand U18609 (N_18609,N_18227,N_18060);
nor U18610 (N_18610,N_18110,N_18057);
or U18611 (N_18611,N_18136,N_18174);
nor U18612 (N_18612,N_18080,N_18491);
xor U18613 (N_18613,N_18114,N_18095);
nor U18614 (N_18614,N_18437,N_18370);
xor U18615 (N_18615,N_18319,N_18232);
or U18616 (N_18616,N_18215,N_18143);
nand U18617 (N_18617,N_18456,N_18061);
and U18618 (N_18618,N_18388,N_18365);
or U18619 (N_18619,N_18461,N_18064);
nand U18620 (N_18620,N_18376,N_18096);
xor U18621 (N_18621,N_18295,N_18201);
xnor U18622 (N_18622,N_18336,N_18361);
xnor U18623 (N_18623,N_18275,N_18000);
and U18624 (N_18624,N_18474,N_18380);
or U18625 (N_18625,N_18467,N_18446);
xnor U18626 (N_18626,N_18265,N_18121);
xnor U18627 (N_18627,N_18065,N_18422);
xor U18628 (N_18628,N_18035,N_18051);
nor U18629 (N_18629,N_18272,N_18258);
or U18630 (N_18630,N_18027,N_18425);
xnor U18631 (N_18631,N_18315,N_18113);
nand U18632 (N_18632,N_18071,N_18211);
nand U18633 (N_18633,N_18053,N_18464);
xnor U18634 (N_18634,N_18316,N_18472);
nand U18635 (N_18635,N_18070,N_18423);
and U18636 (N_18636,N_18068,N_18206);
nor U18637 (N_18637,N_18129,N_18324);
or U18638 (N_18638,N_18207,N_18314);
and U18639 (N_18639,N_18360,N_18412);
nand U18640 (N_18640,N_18346,N_18147);
xor U18641 (N_18641,N_18162,N_18305);
nor U18642 (N_18642,N_18278,N_18148);
nor U18643 (N_18643,N_18094,N_18228);
nor U18644 (N_18644,N_18217,N_18402);
nor U18645 (N_18645,N_18024,N_18054);
or U18646 (N_18646,N_18166,N_18471);
and U18647 (N_18647,N_18312,N_18105);
nor U18648 (N_18648,N_18133,N_18371);
xor U18649 (N_18649,N_18450,N_18103);
nor U18650 (N_18650,N_18439,N_18240);
nor U18651 (N_18651,N_18290,N_18090);
or U18652 (N_18652,N_18164,N_18377);
or U18653 (N_18653,N_18067,N_18043);
and U18654 (N_18654,N_18288,N_18204);
or U18655 (N_18655,N_18072,N_18470);
or U18656 (N_18656,N_18185,N_18357);
nand U18657 (N_18657,N_18202,N_18406);
xor U18658 (N_18658,N_18126,N_18385);
nand U18659 (N_18659,N_18255,N_18285);
xor U18660 (N_18660,N_18205,N_18120);
or U18661 (N_18661,N_18497,N_18382);
xnor U18662 (N_18662,N_18167,N_18409);
nor U18663 (N_18663,N_18487,N_18014);
and U18664 (N_18664,N_18445,N_18182);
nor U18665 (N_18665,N_18284,N_18463);
and U18666 (N_18666,N_18048,N_18203);
xnor U18667 (N_18667,N_18293,N_18495);
xnor U18668 (N_18668,N_18405,N_18152);
xor U18669 (N_18669,N_18451,N_18097);
or U18670 (N_18670,N_18139,N_18074);
xor U18671 (N_18671,N_18200,N_18430);
xor U18672 (N_18672,N_18141,N_18221);
or U18673 (N_18673,N_18341,N_18224);
xor U18674 (N_18674,N_18238,N_18433);
or U18675 (N_18675,N_18453,N_18440);
and U18676 (N_18676,N_18058,N_18156);
or U18677 (N_18677,N_18498,N_18297);
nor U18678 (N_18678,N_18171,N_18335);
or U18679 (N_18679,N_18404,N_18318);
and U18680 (N_18680,N_18101,N_18245);
xnor U18681 (N_18681,N_18233,N_18434);
xnor U18682 (N_18682,N_18187,N_18322);
or U18683 (N_18683,N_18249,N_18462);
nand U18684 (N_18684,N_18063,N_18476);
nor U18685 (N_18685,N_18012,N_18310);
nand U18686 (N_18686,N_18013,N_18188);
and U18687 (N_18687,N_18075,N_18276);
or U18688 (N_18688,N_18056,N_18145);
nand U18689 (N_18689,N_18104,N_18157);
xnor U18690 (N_18690,N_18196,N_18427);
and U18691 (N_18691,N_18140,N_18391);
nand U18692 (N_18692,N_18374,N_18177);
nor U18693 (N_18693,N_18039,N_18320);
and U18694 (N_18694,N_18142,N_18481);
xor U18695 (N_18695,N_18138,N_18209);
or U18696 (N_18696,N_18432,N_18282);
or U18697 (N_18697,N_18150,N_18210);
or U18698 (N_18698,N_18246,N_18119);
and U18699 (N_18699,N_18032,N_18116);
or U18700 (N_18700,N_18118,N_18482);
nand U18701 (N_18701,N_18426,N_18364);
and U18702 (N_18702,N_18420,N_18034);
and U18703 (N_18703,N_18384,N_18331);
nand U18704 (N_18704,N_18271,N_18359);
and U18705 (N_18705,N_18317,N_18475);
or U18706 (N_18706,N_18485,N_18296);
nand U18707 (N_18707,N_18443,N_18334);
xor U18708 (N_18708,N_18363,N_18109);
nor U18709 (N_18709,N_18394,N_18253);
and U18710 (N_18710,N_18264,N_18454);
or U18711 (N_18711,N_18028,N_18328);
nand U18712 (N_18712,N_18031,N_18408);
and U18713 (N_18713,N_18212,N_18387);
or U18714 (N_18714,N_18279,N_18424);
and U18715 (N_18715,N_18259,N_18160);
nor U18716 (N_18716,N_18234,N_18281);
nor U18717 (N_18717,N_18184,N_18137);
xnor U18718 (N_18718,N_18022,N_18260);
nand U18719 (N_18719,N_18358,N_18348);
xnor U18720 (N_18720,N_18351,N_18330);
nor U18721 (N_18721,N_18052,N_18180);
xnor U18722 (N_18722,N_18193,N_18047);
xnor U18723 (N_18723,N_18452,N_18309);
xor U18724 (N_18724,N_18277,N_18132);
nor U18725 (N_18725,N_18244,N_18083);
nor U18726 (N_18726,N_18465,N_18381);
and U18727 (N_18727,N_18499,N_18076);
xor U18728 (N_18728,N_18345,N_18081);
or U18729 (N_18729,N_18066,N_18194);
or U18730 (N_18730,N_18007,N_18213);
nand U18731 (N_18731,N_18192,N_18178);
and U18732 (N_18732,N_18049,N_18021);
and U18733 (N_18733,N_18349,N_18165);
nand U18734 (N_18734,N_18236,N_18078);
nand U18735 (N_18735,N_18332,N_18055);
nor U18736 (N_18736,N_18428,N_18294);
nor U18737 (N_18737,N_18429,N_18410);
nor U18738 (N_18738,N_18484,N_18431);
or U18739 (N_18739,N_18069,N_18002);
or U18740 (N_18740,N_18397,N_18086);
nand U18741 (N_18741,N_18106,N_18340);
and U18742 (N_18742,N_18375,N_18356);
xnor U18743 (N_18743,N_18403,N_18396);
xnor U18744 (N_18744,N_18220,N_18134);
xor U18745 (N_18745,N_18393,N_18144);
nand U18746 (N_18746,N_18417,N_18436);
or U18747 (N_18747,N_18327,N_18037);
nor U18748 (N_18748,N_18044,N_18350);
and U18749 (N_18749,N_18091,N_18308);
nand U18750 (N_18750,N_18217,N_18231);
nand U18751 (N_18751,N_18154,N_18092);
or U18752 (N_18752,N_18404,N_18145);
or U18753 (N_18753,N_18175,N_18336);
and U18754 (N_18754,N_18057,N_18487);
nor U18755 (N_18755,N_18102,N_18448);
nand U18756 (N_18756,N_18145,N_18358);
nand U18757 (N_18757,N_18495,N_18436);
or U18758 (N_18758,N_18389,N_18170);
nor U18759 (N_18759,N_18464,N_18042);
xor U18760 (N_18760,N_18154,N_18231);
xnor U18761 (N_18761,N_18356,N_18430);
and U18762 (N_18762,N_18202,N_18357);
xnor U18763 (N_18763,N_18030,N_18033);
or U18764 (N_18764,N_18141,N_18099);
and U18765 (N_18765,N_18468,N_18226);
xnor U18766 (N_18766,N_18345,N_18055);
nand U18767 (N_18767,N_18494,N_18467);
nand U18768 (N_18768,N_18293,N_18071);
nor U18769 (N_18769,N_18137,N_18439);
and U18770 (N_18770,N_18153,N_18008);
and U18771 (N_18771,N_18359,N_18188);
nand U18772 (N_18772,N_18154,N_18278);
and U18773 (N_18773,N_18492,N_18009);
nor U18774 (N_18774,N_18307,N_18110);
nand U18775 (N_18775,N_18397,N_18003);
nand U18776 (N_18776,N_18170,N_18258);
xor U18777 (N_18777,N_18173,N_18062);
and U18778 (N_18778,N_18164,N_18123);
nor U18779 (N_18779,N_18495,N_18143);
nand U18780 (N_18780,N_18430,N_18082);
nand U18781 (N_18781,N_18142,N_18259);
and U18782 (N_18782,N_18231,N_18219);
nand U18783 (N_18783,N_18232,N_18245);
xor U18784 (N_18784,N_18435,N_18114);
xor U18785 (N_18785,N_18347,N_18172);
nor U18786 (N_18786,N_18191,N_18236);
or U18787 (N_18787,N_18231,N_18148);
nand U18788 (N_18788,N_18017,N_18006);
nor U18789 (N_18789,N_18465,N_18282);
nor U18790 (N_18790,N_18096,N_18020);
xor U18791 (N_18791,N_18153,N_18477);
nor U18792 (N_18792,N_18373,N_18436);
or U18793 (N_18793,N_18375,N_18086);
nor U18794 (N_18794,N_18491,N_18431);
xor U18795 (N_18795,N_18344,N_18059);
nor U18796 (N_18796,N_18422,N_18147);
and U18797 (N_18797,N_18057,N_18406);
xor U18798 (N_18798,N_18025,N_18242);
or U18799 (N_18799,N_18208,N_18062);
and U18800 (N_18800,N_18321,N_18336);
or U18801 (N_18801,N_18245,N_18007);
nand U18802 (N_18802,N_18372,N_18089);
and U18803 (N_18803,N_18304,N_18464);
xor U18804 (N_18804,N_18288,N_18104);
xor U18805 (N_18805,N_18119,N_18174);
nor U18806 (N_18806,N_18306,N_18072);
nand U18807 (N_18807,N_18335,N_18100);
and U18808 (N_18808,N_18006,N_18041);
xor U18809 (N_18809,N_18312,N_18493);
nand U18810 (N_18810,N_18314,N_18076);
and U18811 (N_18811,N_18017,N_18276);
nor U18812 (N_18812,N_18162,N_18112);
or U18813 (N_18813,N_18433,N_18421);
nand U18814 (N_18814,N_18399,N_18388);
nand U18815 (N_18815,N_18141,N_18366);
nand U18816 (N_18816,N_18006,N_18177);
xnor U18817 (N_18817,N_18321,N_18232);
xnor U18818 (N_18818,N_18342,N_18023);
xnor U18819 (N_18819,N_18369,N_18487);
xnor U18820 (N_18820,N_18295,N_18467);
nand U18821 (N_18821,N_18365,N_18333);
nand U18822 (N_18822,N_18060,N_18126);
nand U18823 (N_18823,N_18049,N_18214);
or U18824 (N_18824,N_18459,N_18479);
nor U18825 (N_18825,N_18003,N_18494);
or U18826 (N_18826,N_18048,N_18238);
xor U18827 (N_18827,N_18459,N_18250);
nand U18828 (N_18828,N_18173,N_18467);
nand U18829 (N_18829,N_18210,N_18160);
nor U18830 (N_18830,N_18404,N_18135);
and U18831 (N_18831,N_18444,N_18480);
nand U18832 (N_18832,N_18237,N_18099);
or U18833 (N_18833,N_18366,N_18124);
and U18834 (N_18834,N_18122,N_18074);
xor U18835 (N_18835,N_18298,N_18346);
and U18836 (N_18836,N_18141,N_18071);
nor U18837 (N_18837,N_18013,N_18420);
nor U18838 (N_18838,N_18403,N_18454);
and U18839 (N_18839,N_18091,N_18199);
xnor U18840 (N_18840,N_18023,N_18221);
xnor U18841 (N_18841,N_18411,N_18166);
xnor U18842 (N_18842,N_18139,N_18427);
nand U18843 (N_18843,N_18415,N_18226);
nand U18844 (N_18844,N_18451,N_18391);
and U18845 (N_18845,N_18377,N_18175);
or U18846 (N_18846,N_18076,N_18492);
nor U18847 (N_18847,N_18387,N_18306);
nor U18848 (N_18848,N_18131,N_18438);
xor U18849 (N_18849,N_18488,N_18056);
nand U18850 (N_18850,N_18145,N_18289);
nand U18851 (N_18851,N_18159,N_18359);
nor U18852 (N_18852,N_18396,N_18447);
and U18853 (N_18853,N_18210,N_18173);
nor U18854 (N_18854,N_18032,N_18311);
nand U18855 (N_18855,N_18391,N_18436);
nor U18856 (N_18856,N_18148,N_18386);
nand U18857 (N_18857,N_18208,N_18415);
nor U18858 (N_18858,N_18147,N_18142);
or U18859 (N_18859,N_18112,N_18489);
xnor U18860 (N_18860,N_18339,N_18439);
and U18861 (N_18861,N_18307,N_18220);
nand U18862 (N_18862,N_18256,N_18400);
or U18863 (N_18863,N_18380,N_18247);
xnor U18864 (N_18864,N_18084,N_18010);
and U18865 (N_18865,N_18389,N_18202);
xnor U18866 (N_18866,N_18289,N_18193);
xnor U18867 (N_18867,N_18035,N_18141);
nand U18868 (N_18868,N_18391,N_18110);
and U18869 (N_18869,N_18488,N_18483);
nor U18870 (N_18870,N_18460,N_18089);
xor U18871 (N_18871,N_18331,N_18116);
nand U18872 (N_18872,N_18394,N_18189);
and U18873 (N_18873,N_18481,N_18280);
and U18874 (N_18874,N_18101,N_18113);
and U18875 (N_18875,N_18391,N_18078);
and U18876 (N_18876,N_18497,N_18344);
nand U18877 (N_18877,N_18337,N_18225);
and U18878 (N_18878,N_18002,N_18365);
nand U18879 (N_18879,N_18268,N_18157);
nand U18880 (N_18880,N_18309,N_18030);
nor U18881 (N_18881,N_18237,N_18053);
nand U18882 (N_18882,N_18399,N_18421);
xor U18883 (N_18883,N_18103,N_18451);
and U18884 (N_18884,N_18206,N_18329);
nor U18885 (N_18885,N_18315,N_18203);
xor U18886 (N_18886,N_18208,N_18499);
xnor U18887 (N_18887,N_18209,N_18200);
nor U18888 (N_18888,N_18432,N_18061);
xor U18889 (N_18889,N_18037,N_18340);
xor U18890 (N_18890,N_18132,N_18328);
nor U18891 (N_18891,N_18357,N_18333);
nor U18892 (N_18892,N_18474,N_18240);
and U18893 (N_18893,N_18034,N_18323);
nor U18894 (N_18894,N_18055,N_18297);
and U18895 (N_18895,N_18148,N_18445);
nand U18896 (N_18896,N_18464,N_18237);
xnor U18897 (N_18897,N_18282,N_18330);
xor U18898 (N_18898,N_18253,N_18323);
and U18899 (N_18899,N_18300,N_18000);
xnor U18900 (N_18900,N_18417,N_18188);
xor U18901 (N_18901,N_18348,N_18134);
nand U18902 (N_18902,N_18301,N_18236);
or U18903 (N_18903,N_18019,N_18278);
nor U18904 (N_18904,N_18062,N_18310);
and U18905 (N_18905,N_18007,N_18178);
xor U18906 (N_18906,N_18416,N_18290);
and U18907 (N_18907,N_18329,N_18448);
and U18908 (N_18908,N_18167,N_18050);
and U18909 (N_18909,N_18391,N_18114);
and U18910 (N_18910,N_18103,N_18437);
and U18911 (N_18911,N_18420,N_18439);
xor U18912 (N_18912,N_18030,N_18457);
and U18913 (N_18913,N_18207,N_18013);
or U18914 (N_18914,N_18262,N_18270);
xnor U18915 (N_18915,N_18244,N_18470);
xnor U18916 (N_18916,N_18155,N_18040);
nor U18917 (N_18917,N_18232,N_18268);
and U18918 (N_18918,N_18199,N_18108);
or U18919 (N_18919,N_18045,N_18239);
or U18920 (N_18920,N_18414,N_18467);
or U18921 (N_18921,N_18159,N_18228);
nand U18922 (N_18922,N_18311,N_18203);
and U18923 (N_18923,N_18398,N_18015);
and U18924 (N_18924,N_18464,N_18455);
xor U18925 (N_18925,N_18192,N_18474);
or U18926 (N_18926,N_18071,N_18281);
xor U18927 (N_18927,N_18418,N_18197);
xnor U18928 (N_18928,N_18052,N_18021);
xnor U18929 (N_18929,N_18490,N_18489);
and U18930 (N_18930,N_18417,N_18365);
xor U18931 (N_18931,N_18493,N_18053);
nand U18932 (N_18932,N_18114,N_18468);
xor U18933 (N_18933,N_18387,N_18082);
xnor U18934 (N_18934,N_18470,N_18411);
and U18935 (N_18935,N_18064,N_18279);
or U18936 (N_18936,N_18097,N_18012);
and U18937 (N_18937,N_18142,N_18155);
nor U18938 (N_18938,N_18176,N_18429);
and U18939 (N_18939,N_18176,N_18334);
xor U18940 (N_18940,N_18297,N_18024);
xnor U18941 (N_18941,N_18398,N_18379);
and U18942 (N_18942,N_18318,N_18058);
and U18943 (N_18943,N_18160,N_18258);
and U18944 (N_18944,N_18491,N_18487);
nand U18945 (N_18945,N_18241,N_18130);
and U18946 (N_18946,N_18185,N_18054);
nor U18947 (N_18947,N_18337,N_18309);
nand U18948 (N_18948,N_18237,N_18365);
nor U18949 (N_18949,N_18490,N_18316);
nor U18950 (N_18950,N_18200,N_18429);
or U18951 (N_18951,N_18499,N_18332);
nor U18952 (N_18952,N_18215,N_18141);
xnor U18953 (N_18953,N_18329,N_18170);
and U18954 (N_18954,N_18308,N_18367);
nand U18955 (N_18955,N_18228,N_18497);
or U18956 (N_18956,N_18190,N_18220);
or U18957 (N_18957,N_18166,N_18283);
and U18958 (N_18958,N_18330,N_18398);
or U18959 (N_18959,N_18249,N_18230);
nor U18960 (N_18960,N_18286,N_18271);
xor U18961 (N_18961,N_18280,N_18398);
or U18962 (N_18962,N_18006,N_18363);
or U18963 (N_18963,N_18390,N_18000);
and U18964 (N_18964,N_18359,N_18447);
nor U18965 (N_18965,N_18392,N_18297);
or U18966 (N_18966,N_18269,N_18461);
and U18967 (N_18967,N_18024,N_18338);
nor U18968 (N_18968,N_18109,N_18220);
nor U18969 (N_18969,N_18109,N_18008);
or U18970 (N_18970,N_18091,N_18030);
nor U18971 (N_18971,N_18105,N_18250);
xnor U18972 (N_18972,N_18087,N_18101);
and U18973 (N_18973,N_18247,N_18095);
nor U18974 (N_18974,N_18089,N_18196);
and U18975 (N_18975,N_18389,N_18466);
and U18976 (N_18976,N_18142,N_18207);
or U18977 (N_18977,N_18467,N_18438);
and U18978 (N_18978,N_18454,N_18349);
and U18979 (N_18979,N_18084,N_18443);
xor U18980 (N_18980,N_18369,N_18290);
and U18981 (N_18981,N_18152,N_18176);
and U18982 (N_18982,N_18161,N_18292);
nand U18983 (N_18983,N_18031,N_18377);
and U18984 (N_18984,N_18371,N_18351);
xnor U18985 (N_18985,N_18364,N_18278);
nand U18986 (N_18986,N_18420,N_18309);
nor U18987 (N_18987,N_18013,N_18034);
and U18988 (N_18988,N_18428,N_18467);
and U18989 (N_18989,N_18010,N_18412);
xnor U18990 (N_18990,N_18421,N_18230);
and U18991 (N_18991,N_18339,N_18444);
xor U18992 (N_18992,N_18029,N_18285);
and U18993 (N_18993,N_18335,N_18243);
or U18994 (N_18994,N_18035,N_18335);
or U18995 (N_18995,N_18014,N_18108);
and U18996 (N_18996,N_18483,N_18199);
xnor U18997 (N_18997,N_18064,N_18094);
or U18998 (N_18998,N_18308,N_18056);
or U18999 (N_18999,N_18414,N_18396);
or U19000 (N_19000,N_18645,N_18507);
or U19001 (N_19001,N_18806,N_18933);
nand U19002 (N_19002,N_18849,N_18596);
xnor U19003 (N_19003,N_18535,N_18528);
nor U19004 (N_19004,N_18630,N_18706);
nand U19005 (N_19005,N_18823,N_18710);
or U19006 (N_19006,N_18817,N_18972);
or U19007 (N_19007,N_18796,N_18582);
nor U19008 (N_19008,N_18611,N_18727);
and U19009 (N_19009,N_18649,N_18548);
or U19010 (N_19010,N_18729,N_18916);
nor U19011 (N_19011,N_18731,N_18700);
and U19012 (N_19012,N_18565,N_18624);
nor U19013 (N_19013,N_18835,N_18910);
nand U19014 (N_19014,N_18758,N_18716);
or U19015 (N_19015,N_18604,N_18892);
nor U19016 (N_19016,N_18736,N_18865);
nor U19017 (N_19017,N_18762,N_18693);
nor U19018 (N_19018,N_18973,N_18560);
or U19019 (N_19019,N_18730,N_18629);
nand U19020 (N_19020,N_18574,N_18590);
or U19021 (N_19021,N_18976,N_18905);
nand U19022 (N_19022,N_18821,N_18870);
or U19023 (N_19023,N_18831,N_18673);
nand U19024 (N_19024,N_18967,N_18913);
xnor U19025 (N_19025,N_18832,N_18776);
nand U19026 (N_19026,N_18694,N_18543);
nor U19027 (N_19027,N_18891,N_18887);
nand U19028 (N_19028,N_18778,N_18902);
xnor U19029 (N_19029,N_18552,N_18877);
and U19030 (N_19030,N_18669,N_18707);
nand U19031 (N_19031,N_18920,N_18898);
nor U19032 (N_19032,N_18914,N_18637);
and U19033 (N_19033,N_18826,N_18896);
nand U19034 (N_19034,N_18691,N_18573);
xnor U19035 (N_19035,N_18815,N_18968);
and U19036 (N_19036,N_18740,N_18578);
or U19037 (N_19037,N_18800,N_18512);
nor U19038 (N_19038,N_18789,N_18872);
and U19039 (N_19039,N_18654,N_18718);
nand U19040 (N_19040,N_18948,N_18894);
and U19041 (N_19041,N_18864,N_18955);
or U19042 (N_19042,N_18644,N_18842);
or U19043 (N_19043,N_18575,N_18597);
nor U19044 (N_19044,N_18586,N_18900);
xnor U19045 (N_19045,N_18852,N_18811);
nor U19046 (N_19046,N_18613,N_18585);
nor U19047 (N_19047,N_18745,N_18855);
nand U19048 (N_19048,N_18577,N_18871);
xor U19049 (N_19049,N_18827,N_18873);
or U19050 (N_19050,N_18797,N_18570);
xnor U19051 (N_19051,N_18622,N_18885);
xnor U19052 (N_19052,N_18859,N_18752);
nand U19053 (N_19053,N_18841,N_18840);
or U19054 (N_19054,N_18531,N_18982);
and U19055 (N_19055,N_18805,N_18558);
nor U19056 (N_19056,N_18939,N_18559);
xor U19057 (N_19057,N_18792,N_18812);
or U19058 (N_19058,N_18750,N_18628);
nor U19059 (N_19059,N_18970,N_18862);
or U19060 (N_19060,N_18549,N_18681);
or U19061 (N_19061,N_18818,N_18907);
nor U19062 (N_19062,N_18521,N_18638);
xor U19063 (N_19063,N_18717,N_18500);
nor U19064 (N_19064,N_18991,N_18881);
nand U19065 (N_19065,N_18544,N_18799);
or U19066 (N_19066,N_18663,N_18742);
and U19067 (N_19067,N_18743,N_18860);
or U19068 (N_19068,N_18781,N_18690);
or U19069 (N_19069,N_18779,N_18850);
or U19070 (N_19070,N_18553,N_18834);
nor U19071 (N_19071,N_18788,N_18858);
and U19072 (N_19072,N_18899,N_18770);
xor U19073 (N_19073,N_18768,N_18647);
nand U19074 (N_19074,N_18915,N_18954);
xnor U19075 (N_19075,N_18666,N_18632);
nor U19076 (N_19076,N_18719,N_18616);
or U19077 (N_19077,N_18845,N_18712);
xnor U19078 (N_19078,N_18839,N_18532);
or U19079 (N_19079,N_18748,N_18886);
or U19080 (N_19080,N_18909,N_18904);
nand U19081 (N_19081,N_18912,N_18822);
nand U19082 (N_19082,N_18861,N_18568);
xor U19083 (N_19083,N_18983,N_18966);
nor U19084 (N_19084,N_18600,N_18773);
nand U19085 (N_19085,N_18790,N_18820);
xor U19086 (N_19086,N_18562,N_18828);
nor U19087 (N_19087,N_18659,N_18514);
xor U19088 (N_19088,N_18515,N_18765);
nand U19089 (N_19089,N_18890,N_18678);
nor U19090 (N_19090,N_18656,N_18756);
nand U19091 (N_19091,N_18633,N_18723);
nor U19092 (N_19092,N_18995,N_18876);
nand U19093 (N_19093,N_18988,N_18676);
and U19094 (N_19094,N_18927,N_18592);
nand U19095 (N_19095,N_18520,N_18674);
or U19096 (N_19096,N_18994,N_18889);
nor U19097 (N_19097,N_18935,N_18533);
or U19098 (N_19098,N_18527,N_18506);
nand U19099 (N_19099,N_18696,N_18522);
or U19100 (N_19100,N_18607,N_18567);
xor U19101 (N_19101,N_18857,N_18542);
nor U19102 (N_19102,N_18989,N_18683);
and U19103 (N_19103,N_18614,N_18602);
or U19104 (N_19104,N_18921,N_18657);
and U19105 (N_19105,N_18804,N_18741);
and U19106 (N_19106,N_18516,N_18772);
nand U19107 (N_19107,N_18583,N_18959);
xor U19108 (N_19108,N_18952,N_18829);
and U19109 (N_19109,N_18767,N_18794);
nor U19110 (N_19110,N_18793,N_18941);
and U19111 (N_19111,N_18721,N_18963);
or U19112 (N_19112,N_18884,N_18503);
xor U19113 (N_19113,N_18720,N_18722);
xnor U19114 (N_19114,N_18584,N_18652);
xor U19115 (N_19115,N_18523,N_18878);
or U19116 (N_19116,N_18844,N_18699);
nand U19117 (N_19117,N_18769,N_18687);
and U19118 (N_19118,N_18651,N_18618);
nor U19119 (N_19119,N_18546,N_18711);
nor U19120 (N_19120,N_18668,N_18705);
nor U19121 (N_19121,N_18923,N_18908);
or U19122 (N_19122,N_18650,N_18605);
and U19123 (N_19123,N_18971,N_18809);
xor U19124 (N_19124,N_18938,N_18940);
xnor U19125 (N_19125,N_18919,N_18807);
nand U19126 (N_19126,N_18689,N_18739);
xnor U19127 (N_19127,N_18763,N_18903);
or U19128 (N_19128,N_18934,N_18550);
xor U19129 (N_19129,N_18677,N_18761);
xnor U19130 (N_19130,N_18753,N_18924);
and U19131 (N_19131,N_18709,N_18545);
and U19132 (N_19132,N_18517,N_18942);
nor U19133 (N_19133,N_18996,N_18901);
nor U19134 (N_19134,N_18930,N_18524);
nand U19135 (N_19135,N_18569,N_18813);
nand U19136 (N_19136,N_18639,N_18853);
nor U19137 (N_19137,N_18791,N_18626);
and U19138 (N_19138,N_18897,N_18867);
and U19139 (N_19139,N_18836,N_18642);
and U19140 (N_19140,N_18981,N_18534);
and U19141 (N_19141,N_18974,N_18848);
and U19142 (N_19142,N_18679,N_18610);
xnor U19143 (N_19143,N_18764,N_18888);
nor U19144 (N_19144,N_18843,N_18526);
nand U19145 (N_19145,N_18975,N_18698);
nand U19146 (N_19146,N_18692,N_18958);
or U19147 (N_19147,N_18635,N_18587);
and U19148 (N_19148,N_18634,N_18987);
nand U19149 (N_19149,N_18564,N_18879);
nand U19150 (N_19150,N_18714,N_18738);
or U19151 (N_19151,N_18518,N_18945);
and U19152 (N_19152,N_18874,N_18759);
nor U19153 (N_19153,N_18851,N_18866);
and U19154 (N_19154,N_18755,N_18947);
nand U19155 (N_19155,N_18728,N_18869);
nor U19156 (N_19156,N_18785,N_18598);
or U19157 (N_19157,N_18648,N_18846);
nand U19158 (N_19158,N_18979,N_18803);
nand U19159 (N_19159,N_18715,N_18685);
or U19160 (N_19160,N_18774,N_18675);
nand U19161 (N_19161,N_18906,N_18554);
nor U19162 (N_19162,N_18957,N_18978);
and U19163 (N_19163,N_18641,N_18606);
nor U19164 (N_19164,N_18536,N_18951);
and U19165 (N_19165,N_18833,N_18505);
nand U19166 (N_19166,N_18949,N_18653);
or U19167 (N_19167,N_18928,N_18766);
nor U19168 (N_19168,N_18929,N_18964);
or U19169 (N_19169,N_18992,N_18667);
nor U19170 (N_19170,N_18980,N_18631);
and U19171 (N_19171,N_18501,N_18814);
xor U19172 (N_19172,N_18782,N_18603);
or U19173 (N_19173,N_18737,N_18880);
xnor U19174 (N_19174,N_18786,N_18703);
xnor U19175 (N_19175,N_18619,N_18950);
or U19176 (N_19176,N_18601,N_18985);
nand U19177 (N_19177,N_18581,N_18854);
and U19178 (N_19178,N_18627,N_18608);
or U19179 (N_19179,N_18816,N_18670);
or U19180 (N_19180,N_18724,N_18960);
nor U19181 (N_19181,N_18893,N_18932);
xnor U19182 (N_19182,N_18875,N_18557);
or U19183 (N_19183,N_18882,N_18733);
or U19184 (N_19184,N_18708,N_18922);
nor U19185 (N_19185,N_18771,N_18946);
or U19186 (N_19186,N_18593,N_18795);
nor U19187 (N_19187,N_18686,N_18961);
nand U19188 (N_19188,N_18556,N_18984);
nor U19189 (N_19189,N_18732,N_18688);
nor U19190 (N_19190,N_18625,N_18510);
or U19191 (N_19191,N_18911,N_18615);
nand U19192 (N_19192,N_18682,N_18787);
and U19193 (N_19193,N_18591,N_18956);
and U19194 (N_19194,N_18620,N_18672);
and U19195 (N_19195,N_18671,N_18830);
xnor U19196 (N_19196,N_18918,N_18856);
xnor U19197 (N_19197,N_18965,N_18555);
or U19198 (N_19198,N_18895,N_18917);
nand U19199 (N_19199,N_18749,N_18680);
xnor U19200 (N_19200,N_18810,N_18847);
and U19201 (N_19201,N_18777,N_18986);
nand U19202 (N_19202,N_18697,N_18541);
nor U19203 (N_19203,N_18623,N_18643);
nand U19204 (N_19204,N_18997,N_18513);
xnor U19205 (N_19205,N_18609,N_18931);
xnor U19206 (N_19206,N_18646,N_18746);
and U19207 (N_19207,N_18754,N_18798);
xnor U19208 (N_19208,N_18863,N_18599);
or U19209 (N_19209,N_18735,N_18572);
and U19210 (N_19210,N_18726,N_18519);
or U19211 (N_19211,N_18801,N_18547);
or U19212 (N_19212,N_18713,N_18998);
and U19213 (N_19213,N_18636,N_18757);
nand U19214 (N_19214,N_18775,N_18819);
nor U19215 (N_19215,N_18502,N_18744);
nand U19216 (N_19216,N_18760,N_18538);
nor U19217 (N_19217,N_18808,N_18944);
nand U19218 (N_19218,N_18509,N_18962);
and U19219 (N_19219,N_18655,N_18617);
xor U19220 (N_19220,N_18540,N_18943);
and U19221 (N_19221,N_18612,N_18969);
and U19222 (N_19222,N_18802,N_18508);
or U19223 (N_19223,N_18684,N_18784);
nand U19224 (N_19224,N_18551,N_18621);
or U19225 (N_19225,N_18658,N_18511);
xor U19226 (N_19226,N_18751,N_18594);
xnor U19227 (N_19227,N_18580,N_18576);
and U19228 (N_19228,N_18566,N_18588);
xor U19229 (N_19229,N_18539,N_18595);
xnor U19230 (N_19230,N_18701,N_18504);
and U19231 (N_19231,N_18953,N_18664);
nor U19232 (N_19232,N_18747,N_18925);
nor U19233 (N_19233,N_18640,N_18936);
nor U19234 (N_19234,N_18783,N_18661);
xnor U19235 (N_19235,N_18734,N_18662);
and U19236 (N_19236,N_18937,N_18926);
nand U19237 (N_19237,N_18868,N_18825);
nor U19238 (N_19238,N_18837,N_18702);
or U19239 (N_19239,N_18999,N_18530);
nor U19240 (N_19240,N_18993,N_18589);
nor U19241 (N_19241,N_18561,N_18660);
or U19242 (N_19242,N_18704,N_18571);
or U19243 (N_19243,N_18838,N_18883);
xor U19244 (N_19244,N_18725,N_18579);
or U19245 (N_19245,N_18525,N_18665);
nor U19246 (N_19246,N_18537,N_18780);
nor U19247 (N_19247,N_18563,N_18824);
xor U19248 (N_19248,N_18695,N_18990);
and U19249 (N_19249,N_18529,N_18977);
and U19250 (N_19250,N_18592,N_18666);
nand U19251 (N_19251,N_18719,N_18584);
xnor U19252 (N_19252,N_18698,N_18794);
and U19253 (N_19253,N_18989,N_18503);
nand U19254 (N_19254,N_18921,N_18869);
xor U19255 (N_19255,N_18787,N_18918);
nor U19256 (N_19256,N_18663,N_18575);
and U19257 (N_19257,N_18933,N_18599);
and U19258 (N_19258,N_18656,N_18840);
nor U19259 (N_19259,N_18847,N_18567);
xor U19260 (N_19260,N_18565,N_18838);
nor U19261 (N_19261,N_18919,N_18786);
nand U19262 (N_19262,N_18948,N_18960);
nor U19263 (N_19263,N_18515,N_18917);
xnor U19264 (N_19264,N_18801,N_18925);
nor U19265 (N_19265,N_18953,N_18573);
or U19266 (N_19266,N_18559,N_18556);
or U19267 (N_19267,N_18539,N_18875);
nor U19268 (N_19268,N_18779,N_18910);
or U19269 (N_19269,N_18816,N_18533);
xnor U19270 (N_19270,N_18985,N_18907);
xor U19271 (N_19271,N_18822,N_18836);
nor U19272 (N_19272,N_18736,N_18706);
and U19273 (N_19273,N_18578,N_18662);
xor U19274 (N_19274,N_18518,N_18882);
or U19275 (N_19275,N_18853,N_18925);
xnor U19276 (N_19276,N_18533,N_18866);
nor U19277 (N_19277,N_18580,N_18911);
and U19278 (N_19278,N_18733,N_18735);
xor U19279 (N_19279,N_18947,N_18879);
or U19280 (N_19280,N_18955,N_18865);
xnor U19281 (N_19281,N_18608,N_18625);
nor U19282 (N_19282,N_18516,N_18726);
or U19283 (N_19283,N_18997,N_18854);
or U19284 (N_19284,N_18871,N_18808);
nand U19285 (N_19285,N_18514,N_18923);
or U19286 (N_19286,N_18831,N_18740);
xor U19287 (N_19287,N_18556,N_18652);
xnor U19288 (N_19288,N_18728,N_18847);
or U19289 (N_19289,N_18788,N_18541);
or U19290 (N_19290,N_18976,N_18543);
and U19291 (N_19291,N_18927,N_18643);
or U19292 (N_19292,N_18838,N_18929);
and U19293 (N_19293,N_18900,N_18561);
nor U19294 (N_19294,N_18582,N_18879);
or U19295 (N_19295,N_18621,N_18881);
nand U19296 (N_19296,N_18632,N_18645);
and U19297 (N_19297,N_18558,N_18724);
nand U19298 (N_19298,N_18757,N_18587);
nor U19299 (N_19299,N_18991,N_18703);
nand U19300 (N_19300,N_18828,N_18770);
xor U19301 (N_19301,N_18575,N_18840);
nor U19302 (N_19302,N_18834,N_18732);
xnor U19303 (N_19303,N_18613,N_18853);
nor U19304 (N_19304,N_18829,N_18699);
nand U19305 (N_19305,N_18958,N_18715);
or U19306 (N_19306,N_18556,N_18695);
xnor U19307 (N_19307,N_18843,N_18808);
xor U19308 (N_19308,N_18514,N_18670);
xor U19309 (N_19309,N_18613,N_18975);
nor U19310 (N_19310,N_18966,N_18870);
xnor U19311 (N_19311,N_18994,N_18919);
or U19312 (N_19312,N_18886,N_18710);
or U19313 (N_19313,N_18868,N_18869);
xnor U19314 (N_19314,N_18996,N_18826);
nand U19315 (N_19315,N_18607,N_18851);
or U19316 (N_19316,N_18627,N_18794);
nand U19317 (N_19317,N_18739,N_18966);
or U19318 (N_19318,N_18866,N_18932);
and U19319 (N_19319,N_18918,N_18944);
or U19320 (N_19320,N_18702,N_18622);
or U19321 (N_19321,N_18707,N_18579);
and U19322 (N_19322,N_18894,N_18500);
xnor U19323 (N_19323,N_18764,N_18815);
and U19324 (N_19324,N_18982,N_18822);
or U19325 (N_19325,N_18706,N_18808);
or U19326 (N_19326,N_18970,N_18801);
nand U19327 (N_19327,N_18822,N_18503);
nor U19328 (N_19328,N_18740,N_18802);
nor U19329 (N_19329,N_18918,N_18777);
or U19330 (N_19330,N_18934,N_18873);
and U19331 (N_19331,N_18765,N_18622);
and U19332 (N_19332,N_18914,N_18718);
nor U19333 (N_19333,N_18998,N_18610);
or U19334 (N_19334,N_18789,N_18736);
xor U19335 (N_19335,N_18615,N_18934);
nor U19336 (N_19336,N_18967,N_18523);
and U19337 (N_19337,N_18585,N_18973);
and U19338 (N_19338,N_18870,N_18816);
nand U19339 (N_19339,N_18955,N_18875);
nand U19340 (N_19340,N_18732,N_18712);
or U19341 (N_19341,N_18716,N_18530);
xnor U19342 (N_19342,N_18943,N_18949);
or U19343 (N_19343,N_18834,N_18592);
or U19344 (N_19344,N_18781,N_18589);
or U19345 (N_19345,N_18871,N_18821);
xor U19346 (N_19346,N_18565,N_18564);
nor U19347 (N_19347,N_18537,N_18709);
nor U19348 (N_19348,N_18630,N_18994);
nor U19349 (N_19349,N_18581,N_18993);
nand U19350 (N_19350,N_18537,N_18784);
and U19351 (N_19351,N_18970,N_18650);
xor U19352 (N_19352,N_18882,N_18728);
xnor U19353 (N_19353,N_18822,N_18728);
or U19354 (N_19354,N_18830,N_18589);
and U19355 (N_19355,N_18907,N_18967);
xnor U19356 (N_19356,N_18822,N_18721);
nor U19357 (N_19357,N_18654,N_18831);
or U19358 (N_19358,N_18966,N_18874);
xnor U19359 (N_19359,N_18821,N_18777);
nand U19360 (N_19360,N_18669,N_18934);
nand U19361 (N_19361,N_18577,N_18549);
or U19362 (N_19362,N_18759,N_18668);
or U19363 (N_19363,N_18742,N_18818);
or U19364 (N_19364,N_18802,N_18873);
nand U19365 (N_19365,N_18950,N_18537);
or U19366 (N_19366,N_18719,N_18587);
nand U19367 (N_19367,N_18655,N_18912);
nand U19368 (N_19368,N_18542,N_18652);
nand U19369 (N_19369,N_18659,N_18642);
nor U19370 (N_19370,N_18791,N_18503);
or U19371 (N_19371,N_18757,N_18680);
nand U19372 (N_19372,N_18894,N_18870);
nor U19373 (N_19373,N_18982,N_18661);
nor U19374 (N_19374,N_18753,N_18831);
and U19375 (N_19375,N_18847,N_18521);
and U19376 (N_19376,N_18631,N_18833);
or U19377 (N_19377,N_18829,N_18717);
and U19378 (N_19378,N_18871,N_18772);
or U19379 (N_19379,N_18974,N_18702);
nand U19380 (N_19380,N_18620,N_18575);
nor U19381 (N_19381,N_18895,N_18661);
or U19382 (N_19382,N_18616,N_18888);
nor U19383 (N_19383,N_18859,N_18945);
or U19384 (N_19384,N_18815,N_18849);
and U19385 (N_19385,N_18833,N_18870);
nor U19386 (N_19386,N_18788,N_18954);
or U19387 (N_19387,N_18926,N_18909);
nor U19388 (N_19388,N_18992,N_18782);
nor U19389 (N_19389,N_18595,N_18992);
or U19390 (N_19390,N_18890,N_18739);
and U19391 (N_19391,N_18857,N_18756);
nor U19392 (N_19392,N_18650,N_18528);
nor U19393 (N_19393,N_18576,N_18874);
nor U19394 (N_19394,N_18747,N_18557);
or U19395 (N_19395,N_18648,N_18818);
nor U19396 (N_19396,N_18924,N_18740);
xnor U19397 (N_19397,N_18700,N_18749);
nand U19398 (N_19398,N_18664,N_18901);
nand U19399 (N_19399,N_18572,N_18778);
and U19400 (N_19400,N_18810,N_18842);
nand U19401 (N_19401,N_18949,N_18762);
nor U19402 (N_19402,N_18971,N_18631);
or U19403 (N_19403,N_18586,N_18839);
and U19404 (N_19404,N_18881,N_18558);
or U19405 (N_19405,N_18720,N_18799);
and U19406 (N_19406,N_18589,N_18900);
or U19407 (N_19407,N_18573,N_18975);
and U19408 (N_19408,N_18909,N_18639);
nor U19409 (N_19409,N_18540,N_18897);
or U19410 (N_19410,N_18580,N_18959);
nand U19411 (N_19411,N_18941,N_18746);
nand U19412 (N_19412,N_18965,N_18703);
and U19413 (N_19413,N_18671,N_18654);
or U19414 (N_19414,N_18505,N_18846);
nand U19415 (N_19415,N_18504,N_18600);
and U19416 (N_19416,N_18840,N_18612);
and U19417 (N_19417,N_18603,N_18754);
xnor U19418 (N_19418,N_18522,N_18625);
nand U19419 (N_19419,N_18572,N_18789);
and U19420 (N_19420,N_18724,N_18536);
and U19421 (N_19421,N_18884,N_18587);
nand U19422 (N_19422,N_18687,N_18614);
nor U19423 (N_19423,N_18880,N_18788);
nand U19424 (N_19424,N_18813,N_18929);
or U19425 (N_19425,N_18749,N_18614);
nand U19426 (N_19426,N_18643,N_18522);
and U19427 (N_19427,N_18875,N_18694);
and U19428 (N_19428,N_18704,N_18659);
or U19429 (N_19429,N_18901,N_18663);
xnor U19430 (N_19430,N_18541,N_18591);
xor U19431 (N_19431,N_18559,N_18538);
nor U19432 (N_19432,N_18593,N_18634);
xor U19433 (N_19433,N_18615,N_18868);
and U19434 (N_19434,N_18758,N_18913);
or U19435 (N_19435,N_18612,N_18657);
xor U19436 (N_19436,N_18694,N_18641);
nor U19437 (N_19437,N_18543,N_18912);
and U19438 (N_19438,N_18975,N_18675);
xor U19439 (N_19439,N_18864,N_18558);
nor U19440 (N_19440,N_18959,N_18500);
and U19441 (N_19441,N_18668,N_18849);
nand U19442 (N_19442,N_18715,N_18729);
or U19443 (N_19443,N_18799,N_18636);
or U19444 (N_19444,N_18868,N_18735);
xor U19445 (N_19445,N_18679,N_18860);
xnor U19446 (N_19446,N_18943,N_18944);
and U19447 (N_19447,N_18865,N_18674);
or U19448 (N_19448,N_18626,N_18525);
nand U19449 (N_19449,N_18892,N_18847);
or U19450 (N_19450,N_18722,N_18837);
or U19451 (N_19451,N_18949,N_18687);
or U19452 (N_19452,N_18678,N_18861);
nand U19453 (N_19453,N_18968,N_18840);
nor U19454 (N_19454,N_18626,N_18665);
nand U19455 (N_19455,N_18617,N_18590);
xnor U19456 (N_19456,N_18536,N_18608);
nand U19457 (N_19457,N_18872,N_18817);
and U19458 (N_19458,N_18973,N_18790);
or U19459 (N_19459,N_18531,N_18978);
nand U19460 (N_19460,N_18608,N_18875);
nor U19461 (N_19461,N_18959,N_18951);
or U19462 (N_19462,N_18967,N_18940);
or U19463 (N_19463,N_18762,N_18840);
nor U19464 (N_19464,N_18512,N_18701);
nor U19465 (N_19465,N_18710,N_18963);
and U19466 (N_19466,N_18762,N_18872);
nand U19467 (N_19467,N_18876,N_18848);
nor U19468 (N_19468,N_18866,N_18732);
and U19469 (N_19469,N_18615,N_18558);
and U19470 (N_19470,N_18725,N_18962);
or U19471 (N_19471,N_18724,N_18890);
and U19472 (N_19472,N_18705,N_18925);
nor U19473 (N_19473,N_18878,N_18655);
xnor U19474 (N_19474,N_18793,N_18675);
nand U19475 (N_19475,N_18716,N_18658);
or U19476 (N_19476,N_18543,N_18947);
nor U19477 (N_19477,N_18890,N_18812);
xor U19478 (N_19478,N_18868,N_18907);
or U19479 (N_19479,N_18795,N_18676);
and U19480 (N_19480,N_18893,N_18677);
nand U19481 (N_19481,N_18914,N_18977);
xor U19482 (N_19482,N_18560,N_18896);
or U19483 (N_19483,N_18955,N_18929);
nor U19484 (N_19484,N_18851,N_18645);
nor U19485 (N_19485,N_18512,N_18749);
and U19486 (N_19486,N_18584,N_18947);
nor U19487 (N_19487,N_18709,N_18665);
nor U19488 (N_19488,N_18660,N_18893);
xnor U19489 (N_19489,N_18639,N_18899);
and U19490 (N_19490,N_18701,N_18660);
and U19491 (N_19491,N_18546,N_18833);
or U19492 (N_19492,N_18553,N_18706);
nor U19493 (N_19493,N_18685,N_18792);
and U19494 (N_19494,N_18852,N_18748);
nor U19495 (N_19495,N_18769,N_18897);
nand U19496 (N_19496,N_18895,N_18749);
xnor U19497 (N_19497,N_18967,N_18976);
nand U19498 (N_19498,N_18812,N_18541);
xnor U19499 (N_19499,N_18789,N_18740);
nand U19500 (N_19500,N_19304,N_19418);
nand U19501 (N_19501,N_19423,N_19351);
or U19502 (N_19502,N_19420,N_19051);
and U19503 (N_19503,N_19175,N_19146);
nor U19504 (N_19504,N_19361,N_19435);
and U19505 (N_19505,N_19379,N_19490);
xor U19506 (N_19506,N_19476,N_19133);
and U19507 (N_19507,N_19067,N_19160);
xor U19508 (N_19508,N_19073,N_19303);
xnor U19509 (N_19509,N_19238,N_19348);
nor U19510 (N_19510,N_19168,N_19109);
nor U19511 (N_19511,N_19217,N_19220);
or U19512 (N_19512,N_19413,N_19211);
xor U19513 (N_19513,N_19158,N_19359);
and U19514 (N_19514,N_19330,N_19003);
xnor U19515 (N_19515,N_19154,N_19336);
or U19516 (N_19516,N_19261,N_19322);
and U19517 (N_19517,N_19063,N_19015);
and U19518 (N_19518,N_19159,N_19468);
and U19519 (N_19519,N_19430,N_19077);
xnor U19520 (N_19520,N_19489,N_19444);
xnor U19521 (N_19521,N_19125,N_19378);
nand U19522 (N_19522,N_19108,N_19396);
xor U19523 (N_19523,N_19409,N_19208);
or U19524 (N_19524,N_19149,N_19086);
nand U19525 (N_19525,N_19392,N_19162);
and U19526 (N_19526,N_19122,N_19478);
and U19527 (N_19527,N_19163,N_19152);
and U19528 (N_19528,N_19130,N_19124);
xor U19529 (N_19529,N_19337,N_19453);
and U19530 (N_19530,N_19172,N_19090);
nand U19531 (N_19531,N_19427,N_19150);
or U19532 (N_19532,N_19038,N_19377);
nand U19533 (N_19533,N_19100,N_19284);
xor U19534 (N_19534,N_19030,N_19087);
nor U19535 (N_19535,N_19381,N_19045);
xnor U19536 (N_19536,N_19082,N_19354);
and U19537 (N_19537,N_19400,N_19367);
nor U19538 (N_19538,N_19456,N_19107);
nor U19539 (N_19539,N_19165,N_19137);
xnor U19540 (N_19540,N_19474,N_19389);
and U19541 (N_19541,N_19364,N_19306);
nor U19542 (N_19542,N_19251,N_19385);
xnor U19543 (N_19543,N_19233,N_19411);
or U19544 (N_19544,N_19000,N_19469);
nand U19545 (N_19545,N_19200,N_19243);
or U19546 (N_19546,N_19188,N_19311);
xnor U19547 (N_19547,N_19252,N_19472);
and U19548 (N_19548,N_19282,N_19484);
xnor U19549 (N_19549,N_19041,N_19424);
and U19550 (N_19550,N_19498,N_19157);
xnor U19551 (N_19551,N_19186,N_19260);
xor U19552 (N_19552,N_19017,N_19253);
nand U19553 (N_19553,N_19232,N_19242);
nand U19554 (N_19554,N_19013,N_19237);
xnor U19555 (N_19555,N_19249,N_19245);
nand U19556 (N_19556,N_19450,N_19225);
nor U19557 (N_19557,N_19290,N_19262);
or U19558 (N_19558,N_19401,N_19139);
nand U19559 (N_19559,N_19001,N_19083);
and U19560 (N_19560,N_19278,N_19184);
nand U19561 (N_19561,N_19016,N_19458);
or U19562 (N_19562,N_19452,N_19270);
and U19563 (N_19563,N_19477,N_19023);
nand U19564 (N_19564,N_19391,N_19010);
xor U19565 (N_19565,N_19121,N_19250);
or U19566 (N_19566,N_19374,N_19002);
and U19567 (N_19567,N_19022,N_19328);
or U19568 (N_19568,N_19375,N_19204);
or U19569 (N_19569,N_19174,N_19324);
nand U19570 (N_19570,N_19224,N_19206);
nand U19571 (N_19571,N_19438,N_19214);
and U19572 (N_19572,N_19058,N_19226);
and U19573 (N_19573,N_19425,N_19470);
or U19574 (N_19574,N_19037,N_19187);
nand U19575 (N_19575,N_19399,N_19240);
and U19576 (N_19576,N_19487,N_19296);
nor U19577 (N_19577,N_19321,N_19212);
and U19578 (N_19578,N_19119,N_19235);
or U19579 (N_19579,N_19293,N_19179);
or U19580 (N_19580,N_19177,N_19076);
or U19581 (N_19581,N_19024,N_19061);
and U19582 (N_19582,N_19292,N_19496);
nor U19583 (N_19583,N_19007,N_19471);
and U19584 (N_19584,N_19151,N_19320);
nor U19585 (N_19585,N_19316,N_19056);
and U19586 (N_19586,N_19355,N_19443);
nor U19587 (N_19587,N_19239,N_19228);
nand U19588 (N_19588,N_19035,N_19310);
nor U19589 (N_19589,N_19464,N_19408);
xor U19590 (N_19590,N_19386,N_19466);
nand U19591 (N_19591,N_19429,N_19332);
nand U19592 (N_19592,N_19171,N_19459);
nor U19593 (N_19593,N_19044,N_19368);
nor U19594 (N_19594,N_19446,N_19094);
nor U19595 (N_19595,N_19120,N_19112);
or U19596 (N_19596,N_19205,N_19053);
or U19597 (N_19597,N_19148,N_19315);
and U19598 (N_19598,N_19020,N_19352);
nor U19599 (N_19599,N_19138,N_19365);
and U19600 (N_19600,N_19366,N_19440);
nor U19601 (N_19601,N_19495,N_19027);
or U19602 (N_19602,N_19263,N_19173);
nor U19603 (N_19603,N_19319,N_19380);
nand U19604 (N_19604,N_19092,N_19445);
and U19605 (N_19605,N_19104,N_19405);
xnor U19606 (N_19606,N_19447,N_19300);
xnor U19607 (N_19607,N_19285,N_19074);
nor U19608 (N_19608,N_19054,N_19075);
nand U19609 (N_19609,N_19031,N_19271);
nor U19610 (N_19610,N_19481,N_19195);
or U19611 (N_19611,N_19091,N_19080);
xor U19612 (N_19612,N_19442,N_19126);
nand U19613 (N_19613,N_19140,N_19115);
nand U19614 (N_19614,N_19323,N_19387);
or U19615 (N_19615,N_19064,N_19431);
or U19616 (N_19616,N_19455,N_19236);
or U19617 (N_19617,N_19181,N_19393);
or U19618 (N_19618,N_19089,N_19416);
nand U19619 (N_19619,N_19190,N_19096);
nor U19620 (N_19620,N_19347,N_19118);
or U19621 (N_19621,N_19215,N_19398);
and U19622 (N_19622,N_19488,N_19299);
or U19623 (N_19623,N_19098,N_19461);
and U19624 (N_19624,N_19196,N_19185);
or U19625 (N_19625,N_19014,N_19065);
or U19626 (N_19626,N_19264,N_19275);
or U19627 (N_19627,N_19417,N_19426);
nor U19628 (N_19628,N_19071,N_19277);
xnor U19629 (N_19629,N_19167,N_19265);
nor U19630 (N_19630,N_19032,N_19259);
nand U19631 (N_19631,N_19371,N_19410);
nor U19632 (N_19632,N_19170,N_19213);
xor U19633 (N_19633,N_19216,N_19349);
xor U19634 (N_19634,N_19297,N_19201);
or U19635 (N_19635,N_19345,N_19166);
and U19636 (N_19636,N_19189,N_19403);
nand U19637 (N_19637,N_19331,N_19338);
nor U19638 (N_19638,N_19329,N_19273);
xor U19639 (N_19639,N_19407,N_19207);
and U19640 (N_19640,N_19388,N_19372);
xor U19641 (N_19641,N_19286,N_19369);
and U19642 (N_19642,N_19376,N_19419);
nand U19643 (N_19643,N_19356,N_19218);
nor U19644 (N_19644,N_19143,N_19111);
xnor U19645 (N_19645,N_19008,N_19103);
or U19646 (N_19646,N_19467,N_19040);
nand U19647 (N_19647,N_19287,N_19117);
nand U19648 (N_19648,N_19258,N_19390);
xor U19649 (N_19649,N_19192,N_19301);
and U19650 (N_19650,N_19101,N_19072);
nor U19651 (N_19651,N_19383,N_19004);
nand U19652 (N_19652,N_19169,N_19473);
xnor U19653 (N_19653,N_19436,N_19475);
and U19654 (N_19654,N_19033,N_19019);
nor U19655 (N_19655,N_19088,N_19341);
nand U19656 (N_19656,N_19194,N_19132);
nor U19657 (N_19657,N_19312,N_19123);
xor U19658 (N_19658,N_19486,N_19268);
nand U19659 (N_19659,N_19248,N_19210);
and U19660 (N_19660,N_19283,N_19437);
xor U19661 (N_19661,N_19081,N_19256);
xor U19662 (N_19662,N_19281,N_19317);
nor U19663 (N_19663,N_19449,N_19079);
xnor U19664 (N_19664,N_19362,N_19421);
xor U19665 (N_19665,N_19127,N_19334);
nand U19666 (N_19666,N_19448,N_19463);
nand U19667 (N_19667,N_19183,N_19145);
and U19668 (N_19668,N_19113,N_19497);
and U19669 (N_19669,N_19156,N_19428);
nor U19670 (N_19670,N_19343,N_19397);
nand U19671 (N_19671,N_19018,N_19454);
xnor U19672 (N_19672,N_19493,N_19485);
nor U19673 (N_19673,N_19241,N_19360);
xnor U19674 (N_19674,N_19147,N_19274);
xor U19675 (N_19675,N_19255,N_19223);
xnor U19676 (N_19676,N_19026,N_19085);
xor U19677 (N_19677,N_19093,N_19342);
or U19678 (N_19678,N_19494,N_19234);
nand U19679 (N_19679,N_19070,N_19247);
and U19680 (N_19680,N_19460,N_19178);
nand U19681 (N_19681,N_19308,N_19221);
nand U19682 (N_19682,N_19483,N_19307);
nand U19683 (N_19683,N_19350,N_19394);
nand U19684 (N_19684,N_19357,N_19344);
nor U19685 (N_19685,N_19084,N_19095);
nor U19686 (N_19686,N_19021,N_19314);
nand U19687 (N_19687,N_19006,N_19062);
nand U19688 (N_19688,N_19294,N_19289);
xnor U19689 (N_19689,N_19049,N_19042);
nand U19690 (N_19690,N_19333,N_19462);
nor U19691 (N_19691,N_19193,N_19039);
or U19692 (N_19692,N_19298,N_19465);
and U19693 (N_19693,N_19370,N_19059);
nand U19694 (N_19694,N_19227,N_19036);
nor U19695 (N_19695,N_19231,N_19395);
nor U19696 (N_19696,N_19128,N_19219);
and U19697 (N_19697,N_19164,N_19102);
xor U19698 (N_19698,N_19346,N_19025);
and U19699 (N_19699,N_19131,N_19499);
nor U19700 (N_19700,N_19028,N_19129);
nand U19701 (N_19701,N_19327,N_19142);
nor U19702 (N_19702,N_19155,N_19309);
xor U19703 (N_19703,N_19302,N_19011);
and U19704 (N_19704,N_19029,N_19406);
xor U19705 (N_19705,N_19373,N_19402);
nor U19706 (N_19706,N_19441,N_19340);
and U19707 (N_19707,N_19055,N_19222);
and U19708 (N_19708,N_19313,N_19105);
xnor U19709 (N_19709,N_19339,N_19116);
or U19710 (N_19710,N_19491,N_19305);
xor U19711 (N_19711,N_19451,N_19203);
and U19712 (N_19712,N_19057,N_19229);
or U19713 (N_19713,N_19078,N_19097);
and U19714 (N_19714,N_19197,N_19335);
nand U19715 (N_19715,N_19230,N_19295);
or U19716 (N_19716,N_19353,N_19439);
nand U19717 (N_19717,N_19246,N_19069);
nor U19718 (N_19718,N_19060,N_19280);
and U19719 (N_19719,N_19363,N_19318);
and U19720 (N_19720,N_19209,N_19276);
xnor U19721 (N_19721,N_19291,N_19176);
or U19722 (N_19722,N_19202,N_19161);
and U19723 (N_19723,N_19043,N_19034);
nand U19724 (N_19724,N_19144,N_19432);
xnor U19725 (N_19725,N_19012,N_19180);
nor U19726 (N_19726,N_19480,N_19272);
nor U19727 (N_19727,N_19048,N_19279);
or U19728 (N_19728,N_19457,N_19136);
nand U19729 (N_19729,N_19254,N_19182);
xnor U19730 (N_19730,N_19047,N_19482);
nor U19731 (N_19731,N_19135,N_19191);
and U19732 (N_19732,N_19153,N_19244);
nand U19733 (N_19733,N_19269,N_19099);
nor U19734 (N_19734,N_19325,N_19492);
nand U19735 (N_19735,N_19412,N_19052);
xor U19736 (N_19736,N_19415,N_19066);
nor U19737 (N_19737,N_19358,N_19134);
xor U19738 (N_19738,N_19434,N_19106);
nor U19739 (N_19739,N_19199,N_19009);
and U19740 (N_19740,N_19198,N_19422);
and U19741 (N_19741,N_19288,N_19068);
and U19742 (N_19742,N_19384,N_19433);
nand U19743 (N_19743,N_19326,N_19050);
nand U19744 (N_19744,N_19257,N_19404);
nand U19745 (N_19745,N_19141,N_19266);
nand U19746 (N_19746,N_19479,N_19382);
and U19747 (N_19747,N_19046,N_19267);
or U19748 (N_19748,N_19005,N_19114);
nand U19749 (N_19749,N_19110,N_19414);
nand U19750 (N_19750,N_19174,N_19386);
nand U19751 (N_19751,N_19328,N_19130);
and U19752 (N_19752,N_19204,N_19350);
nor U19753 (N_19753,N_19393,N_19412);
nor U19754 (N_19754,N_19001,N_19141);
and U19755 (N_19755,N_19148,N_19078);
and U19756 (N_19756,N_19091,N_19321);
or U19757 (N_19757,N_19186,N_19350);
xor U19758 (N_19758,N_19368,N_19326);
nor U19759 (N_19759,N_19008,N_19360);
nand U19760 (N_19760,N_19111,N_19109);
nand U19761 (N_19761,N_19033,N_19440);
xnor U19762 (N_19762,N_19251,N_19190);
or U19763 (N_19763,N_19433,N_19270);
or U19764 (N_19764,N_19371,N_19320);
or U19765 (N_19765,N_19117,N_19251);
or U19766 (N_19766,N_19239,N_19419);
nor U19767 (N_19767,N_19091,N_19456);
nor U19768 (N_19768,N_19186,N_19322);
nand U19769 (N_19769,N_19082,N_19033);
nor U19770 (N_19770,N_19041,N_19073);
xor U19771 (N_19771,N_19269,N_19139);
xor U19772 (N_19772,N_19156,N_19413);
and U19773 (N_19773,N_19161,N_19235);
nor U19774 (N_19774,N_19243,N_19169);
or U19775 (N_19775,N_19428,N_19005);
xor U19776 (N_19776,N_19484,N_19232);
xor U19777 (N_19777,N_19017,N_19222);
or U19778 (N_19778,N_19239,N_19221);
nor U19779 (N_19779,N_19222,N_19271);
and U19780 (N_19780,N_19299,N_19205);
xnor U19781 (N_19781,N_19159,N_19190);
or U19782 (N_19782,N_19060,N_19307);
nand U19783 (N_19783,N_19145,N_19217);
xnor U19784 (N_19784,N_19058,N_19010);
or U19785 (N_19785,N_19128,N_19112);
or U19786 (N_19786,N_19093,N_19204);
xnor U19787 (N_19787,N_19038,N_19262);
xnor U19788 (N_19788,N_19198,N_19236);
nor U19789 (N_19789,N_19382,N_19187);
xnor U19790 (N_19790,N_19031,N_19070);
xor U19791 (N_19791,N_19249,N_19149);
nand U19792 (N_19792,N_19117,N_19260);
or U19793 (N_19793,N_19397,N_19434);
xnor U19794 (N_19794,N_19090,N_19485);
or U19795 (N_19795,N_19399,N_19441);
nand U19796 (N_19796,N_19324,N_19213);
and U19797 (N_19797,N_19314,N_19410);
and U19798 (N_19798,N_19419,N_19195);
and U19799 (N_19799,N_19066,N_19296);
and U19800 (N_19800,N_19274,N_19396);
nand U19801 (N_19801,N_19163,N_19336);
xor U19802 (N_19802,N_19428,N_19112);
nor U19803 (N_19803,N_19053,N_19375);
or U19804 (N_19804,N_19472,N_19192);
and U19805 (N_19805,N_19205,N_19203);
or U19806 (N_19806,N_19146,N_19346);
xor U19807 (N_19807,N_19078,N_19114);
nor U19808 (N_19808,N_19147,N_19325);
nor U19809 (N_19809,N_19328,N_19371);
nand U19810 (N_19810,N_19010,N_19118);
xnor U19811 (N_19811,N_19214,N_19263);
nand U19812 (N_19812,N_19209,N_19359);
xnor U19813 (N_19813,N_19489,N_19185);
and U19814 (N_19814,N_19353,N_19100);
or U19815 (N_19815,N_19400,N_19068);
nor U19816 (N_19816,N_19404,N_19494);
nand U19817 (N_19817,N_19231,N_19084);
and U19818 (N_19818,N_19107,N_19231);
xnor U19819 (N_19819,N_19133,N_19220);
or U19820 (N_19820,N_19466,N_19305);
and U19821 (N_19821,N_19165,N_19139);
nand U19822 (N_19822,N_19007,N_19206);
nor U19823 (N_19823,N_19211,N_19395);
or U19824 (N_19824,N_19056,N_19135);
and U19825 (N_19825,N_19365,N_19493);
or U19826 (N_19826,N_19151,N_19190);
xnor U19827 (N_19827,N_19016,N_19047);
xnor U19828 (N_19828,N_19443,N_19440);
and U19829 (N_19829,N_19374,N_19388);
nand U19830 (N_19830,N_19274,N_19123);
nor U19831 (N_19831,N_19129,N_19428);
xor U19832 (N_19832,N_19447,N_19423);
xor U19833 (N_19833,N_19277,N_19283);
or U19834 (N_19834,N_19359,N_19306);
xnor U19835 (N_19835,N_19438,N_19090);
and U19836 (N_19836,N_19288,N_19092);
nand U19837 (N_19837,N_19154,N_19351);
and U19838 (N_19838,N_19473,N_19262);
nand U19839 (N_19839,N_19037,N_19460);
xor U19840 (N_19840,N_19220,N_19409);
and U19841 (N_19841,N_19309,N_19327);
nand U19842 (N_19842,N_19439,N_19429);
nor U19843 (N_19843,N_19083,N_19063);
nor U19844 (N_19844,N_19328,N_19332);
and U19845 (N_19845,N_19245,N_19044);
nor U19846 (N_19846,N_19352,N_19219);
or U19847 (N_19847,N_19134,N_19437);
nand U19848 (N_19848,N_19022,N_19476);
xnor U19849 (N_19849,N_19295,N_19449);
nand U19850 (N_19850,N_19416,N_19311);
nor U19851 (N_19851,N_19199,N_19192);
or U19852 (N_19852,N_19134,N_19359);
or U19853 (N_19853,N_19110,N_19281);
nand U19854 (N_19854,N_19055,N_19127);
xnor U19855 (N_19855,N_19373,N_19050);
and U19856 (N_19856,N_19353,N_19267);
xor U19857 (N_19857,N_19139,N_19454);
or U19858 (N_19858,N_19335,N_19044);
xnor U19859 (N_19859,N_19406,N_19271);
xnor U19860 (N_19860,N_19289,N_19435);
and U19861 (N_19861,N_19257,N_19338);
and U19862 (N_19862,N_19142,N_19002);
xor U19863 (N_19863,N_19372,N_19001);
and U19864 (N_19864,N_19087,N_19179);
and U19865 (N_19865,N_19269,N_19073);
or U19866 (N_19866,N_19017,N_19433);
nor U19867 (N_19867,N_19122,N_19306);
nand U19868 (N_19868,N_19332,N_19041);
xor U19869 (N_19869,N_19189,N_19106);
and U19870 (N_19870,N_19273,N_19069);
nor U19871 (N_19871,N_19387,N_19123);
and U19872 (N_19872,N_19074,N_19171);
or U19873 (N_19873,N_19308,N_19313);
xnor U19874 (N_19874,N_19464,N_19355);
xor U19875 (N_19875,N_19362,N_19436);
xnor U19876 (N_19876,N_19449,N_19249);
nand U19877 (N_19877,N_19366,N_19495);
xnor U19878 (N_19878,N_19219,N_19046);
and U19879 (N_19879,N_19076,N_19059);
xnor U19880 (N_19880,N_19235,N_19443);
or U19881 (N_19881,N_19234,N_19211);
nand U19882 (N_19882,N_19366,N_19352);
nand U19883 (N_19883,N_19310,N_19111);
and U19884 (N_19884,N_19456,N_19352);
nor U19885 (N_19885,N_19306,N_19455);
and U19886 (N_19886,N_19328,N_19285);
nor U19887 (N_19887,N_19243,N_19390);
or U19888 (N_19888,N_19477,N_19396);
and U19889 (N_19889,N_19463,N_19323);
and U19890 (N_19890,N_19027,N_19385);
and U19891 (N_19891,N_19258,N_19459);
nand U19892 (N_19892,N_19125,N_19228);
nand U19893 (N_19893,N_19470,N_19403);
and U19894 (N_19894,N_19019,N_19444);
or U19895 (N_19895,N_19063,N_19109);
xnor U19896 (N_19896,N_19028,N_19194);
xnor U19897 (N_19897,N_19449,N_19425);
and U19898 (N_19898,N_19321,N_19332);
or U19899 (N_19899,N_19085,N_19342);
and U19900 (N_19900,N_19312,N_19298);
nor U19901 (N_19901,N_19405,N_19362);
or U19902 (N_19902,N_19421,N_19316);
xnor U19903 (N_19903,N_19412,N_19104);
and U19904 (N_19904,N_19383,N_19216);
nand U19905 (N_19905,N_19300,N_19118);
nor U19906 (N_19906,N_19212,N_19364);
nand U19907 (N_19907,N_19438,N_19180);
nor U19908 (N_19908,N_19035,N_19375);
nand U19909 (N_19909,N_19222,N_19163);
nor U19910 (N_19910,N_19419,N_19478);
nor U19911 (N_19911,N_19331,N_19166);
nand U19912 (N_19912,N_19398,N_19450);
and U19913 (N_19913,N_19078,N_19153);
nand U19914 (N_19914,N_19326,N_19415);
nand U19915 (N_19915,N_19022,N_19075);
xnor U19916 (N_19916,N_19051,N_19264);
nor U19917 (N_19917,N_19230,N_19276);
or U19918 (N_19918,N_19142,N_19140);
xnor U19919 (N_19919,N_19245,N_19419);
nor U19920 (N_19920,N_19254,N_19349);
or U19921 (N_19921,N_19279,N_19087);
and U19922 (N_19922,N_19391,N_19092);
or U19923 (N_19923,N_19391,N_19085);
or U19924 (N_19924,N_19214,N_19067);
nor U19925 (N_19925,N_19047,N_19379);
or U19926 (N_19926,N_19286,N_19245);
xor U19927 (N_19927,N_19424,N_19097);
nand U19928 (N_19928,N_19027,N_19209);
xnor U19929 (N_19929,N_19267,N_19059);
nor U19930 (N_19930,N_19183,N_19441);
xor U19931 (N_19931,N_19007,N_19234);
nand U19932 (N_19932,N_19389,N_19158);
nand U19933 (N_19933,N_19142,N_19440);
nor U19934 (N_19934,N_19229,N_19004);
and U19935 (N_19935,N_19251,N_19150);
nand U19936 (N_19936,N_19195,N_19434);
and U19937 (N_19937,N_19148,N_19292);
or U19938 (N_19938,N_19021,N_19389);
or U19939 (N_19939,N_19477,N_19147);
or U19940 (N_19940,N_19385,N_19154);
nor U19941 (N_19941,N_19248,N_19284);
nand U19942 (N_19942,N_19066,N_19129);
xor U19943 (N_19943,N_19202,N_19182);
or U19944 (N_19944,N_19023,N_19216);
xnor U19945 (N_19945,N_19221,N_19178);
and U19946 (N_19946,N_19432,N_19009);
xnor U19947 (N_19947,N_19211,N_19032);
nor U19948 (N_19948,N_19131,N_19410);
and U19949 (N_19949,N_19200,N_19448);
nor U19950 (N_19950,N_19237,N_19134);
nand U19951 (N_19951,N_19281,N_19183);
or U19952 (N_19952,N_19259,N_19463);
nor U19953 (N_19953,N_19315,N_19373);
nand U19954 (N_19954,N_19361,N_19430);
and U19955 (N_19955,N_19082,N_19336);
or U19956 (N_19956,N_19412,N_19077);
and U19957 (N_19957,N_19221,N_19123);
or U19958 (N_19958,N_19214,N_19237);
xor U19959 (N_19959,N_19446,N_19104);
xor U19960 (N_19960,N_19232,N_19288);
or U19961 (N_19961,N_19479,N_19034);
and U19962 (N_19962,N_19184,N_19320);
or U19963 (N_19963,N_19480,N_19419);
nor U19964 (N_19964,N_19354,N_19264);
nand U19965 (N_19965,N_19085,N_19321);
xnor U19966 (N_19966,N_19130,N_19044);
or U19967 (N_19967,N_19382,N_19039);
nand U19968 (N_19968,N_19236,N_19051);
and U19969 (N_19969,N_19059,N_19212);
nor U19970 (N_19970,N_19460,N_19107);
xor U19971 (N_19971,N_19481,N_19163);
nand U19972 (N_19972,N_19029,N_19231);
nor U19973 (N_19973,N_19405,N_19005);
xnor U19974 (N_19974,N_19308,N_19068);
xor U19975 (N_19975,N_19417,N_19018);
xnor U19976 (N_19976,N_19497,N_19237);
and U19977 (N_19977,N_19127,N_19237);
xor U19978 (N_19978,N_19480,N_19218);
nor U19979 (N_19979,N_19140,N_19453);
xnor U19980 (N_19980,N_19241,N_19497);
and U19981 (N_19981,N_19493,N_19092);
or U19982 (N_19982,N_19256,N_19195);
and U19983 (N_19983,N_19195,N_19013);
nor U19984 (N_19984,N_19349,N_19110);
nand U19985 (N_19985,N_19023,N_19083);
and U19986 (N_19986,N_19045,N_19356);
xnor U19987 (N_19987,N_19073,N_19082);
nor U19988 (N_19988,N_19322,N_19199);
and U19989 (N_19989,N_19259,N_19392);
or U19990 (N_19990,N_19273,N_19117);
xnor U19991 (N_19991,N_19459,N_19096);
xor U19992 (N_19992,N_19090,N_19138);
nand U19993 (N_19993,N_19296,N_19123);
nand U19994 (N_19994,N_19082,N_19134);
or U19995 (N_19995,N_19234,N_19330);
or U19996 (N_19996,N_19228,N_19077);
nor U19997 (N_19997,N_19089,N_19494);
and U19998 (N_19998,N_19069,N_19376);
and U19999 (N_19999,N_19088,N_19297);
and U20000 (N_20000,N_19555,N_19658);
xnor U20001 (N_20001,N_19630,N_19774);
and U20002 (N_20002,N_19900,N_19510);
xnor U20003 (N_20003,N_19515,N_19558);
or U20004 (N_20004,N_19699,N_19566);
nand U20005 (N_20005,N_19870,N_19969);
nand U20006 (N_20006,N_19990,N_19679);
or U20007 (N_20007,N_19924,N_19741);
xnor U20008 (N_20008,N_19604,N_19633);
xor U20009 (N_20009,N_19749,N_19761);
nand U20010 (N_20010,N_19542,N_19512);
nand U20011 (N_20011,N_19675,N_19597);
or U20012 (N_20012,N_19618,N_19746);
and U20013 (N_20013,N_19583,N_19757);
nand U20014 (N_20014,N_19948,N_19937);
or U20015 (N_20015,N_19502,N_19765);
nor U20016 (N_20016,N_19895,N_19753);
nand U20017 (N_20017,N_19918,N_19603);
nor U20018 (N_20018,N_19958,N_19607);
xor U20019 (N_20019,N_19686,N_19609);
or U20020 (N_20020,N_19876,N_19816);
nand U20021 (N_20021,N_19561,N_19782);
nand U20022 (N_20022,N_19581,N_19522);
nor U20023 (N_20023,N_19513,N_19683);
or U20024 (N_20024,N_19756,N_19552);
and U20025 (N_20025,N_19664,N_19790);
nand U20026 (N_20026,N_19810,N_19826);
nor U20027 (N_20027,N_19734,N_19562);
xnor U20028 (N_20028,N_19942,N_19696);
nor U20029 (N_20029,N_19639,N_19856);
or U20030 (N_20030,N_19579,N_19845);
or U20031 (N_20031,N_19649,N_19963);
or U20032 (N_20032,N_19913,N_19935);
nand U20033 (N_20033,N_19614,N_19640);
nand U20034 (N_20034,N_19500,N_19925);
nor U20035 (N_20035,N_19844,N_19612);
or U20036 (N_20036,N_19673,N_19668);
nand U20037 (N_20037,N_19724,N_19674);
and U20038 (N_20038,N_19939,N_19827);
nor U20039 (N_20039,N_19831,N_19771);
xor U20040 (N_20040,N_19571,N_19824);
nand U20041 (N_20041,N_19687,N_19634);
or U20042 (N_20042,N_19823,N_19751);
or U20043 (N_20043,N_19800,N_19892);
nor U20044 (N_20044,N_19930,N_19898);
nand U20045 (N_20045,N_19791,N_19954);
nor U20046 (N_20046,N_19569,N_19672);
or U20047 (N_20047,N_19884,N_19815);
xnor U20048 (N_20048,N_19952,N_19706);
nand U20049 (N_20049,N_19722,N_19999);
and U20050 (N_20050,N_19694,N_19803);
nor U20051 (N_20051,N_19835,N_19795);
and U20052 (N_20052,N_19850,N_19528);
or U20053 (N_20053,N_19965,N_19615);
nand U20054 (N_20054,N_19654,N_19773);
nand U20055 (N_20055,N_19585,N_19540);
xor U20056 (N_20056,N_19716,N_19986);
xor U20057 (N_20057,N_19855,N_19647);
and U20058 (N_20058,N_19915,N_19933);
xor U20059 (N_20059,N_19828,N_19886);
or U20060 (N_20060,N_19802,N_19692);
nand U20061 (N_20061,N_19594,N_19878);
nand U20062 (N_20062,N_19703,N_19707);
nand U20063 (N_20063,N_19993,N_19830);
xnor U20064 (N_20064,N_19872,N_19956);
nand U20065 (N_20065,N_19610,N_19841);
nor U20066 (N_20066,N_19588,N_19992);
xnor U20067 (N_20067,N_19789,N_19521);
and U20068 (N_20068,N_19702,N_19662);
xor U20069 (N_20069,N_19661,N_19742);
and U20070 (N_20070,N_19573,N_19723);
xor U20071 (N_20071,N_19953,N_19605);
xnor U20072 (N_20072,N_19635,N_19794);
and U20073 (N_20073,N_19887,N_19981);
and U20074 (N_20074,N_19893,N_19919);
nor U20075 (N_20075,N_19681,N_19508);
nand U20076 (N_20076,N_19584,N_19978);
or U20077 (N_20077,N_19690,N_19866);
nor U20078 (N_20078,N_19621,N_19667);
or U20079 (N_20079,N_19917,N_19677);
or U20080 (N_20080,N_19665,N_19806);
nand U20081 (N_20081,N_19975,N_19813);
nand U20082 (N_20082,N_19670,N_19541);
or U20083 (N_20083,N_19931,N_19808);
nor U20084 (N_20084,N_19807,N_19736);
xnor U20085 (N_20085,N_19567,N_19595);
xor U20086 (N_20086,N_19962,N_19851);
nand U20087 (N_20087,N_19908,N_19708);
xor U20088 (N_20088,N_19998,N_19971);
nor U20089 (N_20089,N_19941,N_19889);
xnor U20090 (N_20090,N_19783,N_19559);
nor U20091 (N_20091,N_19564,N_19503);
or U20092 (N_20092,N_19881,N_19821);
nand U20093 (N_20093,N_19580,N_19611);
or U20094 (N_20094,N_19758,N_19682);
nor U20095 (N_20095,N_19625,N_19775);
or U20096 (N_20096,N_19593,N_19904);
nor U20097 (N_20097,N_19711,N_19947);
and U20098 (N_20098,N_19617,N_19590);
xor U20099 (N_20099,N_19659,N_19720);
nor U20100 (N_20100,N_19620,N_19713);
nor U20101 (N_20101,N_19680,N_19781);
nor U20102 (N_20102,N_19899,N_19518);
xor U20103 (N_20103,N_19530,N_19606);
nor U20104 (N_20104,N_19601,N_19766);
or U20105 (N_20105,N_19767,N_19860);
or U20106 (N_20106,N_19853,N_19959);
nand U20107 (N_20107,N_19875,N_19576);
and U20108 (N_20108,N_19764,N_19636);
xnor U20109 (N_20109,N_19575,N_19516);
nor U20110 (N_20110,N_19743,N_19747);
or U20111 (N_20111,N_19652,N_19712);
or U20112 (N_20112,N_19921,N_19587);
nor U20113 (N_20113,N_19685,N_19849);
xnor U20114 (N_20114,N_19988,N_19506);
nor U20115 (N_20115,N_19565,N_19907);
or U20116 (N_20116,N_19519,N_19832);
or U20117 (N_20117,N_19560,N_19922);
xnor U20118 (N_20118,N_19987,N_19535);
or U20119 (N_20119,N_19750,N_19985);
nor U20120 (N_20120,N_19619,N_19780);
xnor U20121 (N_20121,N_19678,N_19883);
or U20122 (N_20122,N_19996,N_19622);
nor U20123 (N_20123,N_19834,N_19950);
and U20124 (N_20124,N_19762,N_19650);
or U20125 (N_20125,N_19691,N_19777);
nand U20126 (N_20126,N_19745,N_19570);
or U20127 (N_20127,N_19859,N_19563);
nand U20128 (N_20128,N_19727,N_19877);
or U20129 (N_20129,N_19890,N_19920);
and U20130 (N_20130,N_19602,N_19550);
and U20131 (N_20131,N_19738,N_19863);
nor U20132 (N_20132,N_19509,N_19531);
xnor U20133 (N_20133,N_19995,N_19906);
and U20134 (N_20134,N_19546,N_19578);
xor U20135 (N_20135,N_19772,N_19949);
nor U20136 (N_20136,N_19505,N_19770);
nand U20137 (N_20137,N_19582,N_19520);
or U20138 (N_20138,N_19936,N_19905);
xnor U20139 (N_20139,N_19754,N_19852);
xor U20140 (N_20140,N_19651,N_19538);
xor U20141 (N_20141,N_19637,N_19785);
or U20142 (N_20142,N_19547,N_19655);
nand U20143 (N_20143,N_19600,N_19669);
or U20144 (N_20144,N_19778,N_19974);
xor U20145 (N_20145,N_19534,N_19966);
xnor U20146 (N_20146,N_19577,N_19737);
and U20147 (N_20147,N_19833,N_19693);
or U20148 (N_20148,N_19689,N_19786);
or U20149 (N_20149,N_19631,N_19556);
and U20150 (N_20150,N_19728,N_19858);
nand U20151 (N_20151,N_19784,N_19896);
and U20152 (N_20152,N_19970,N_19874);
xnor U20153 (N_20153,N_19861,N_19836);
and U20154 (N_20154,N_19788,N_19549);
xnor U20155 (N_20155,N_19589,N_19525);
nand U20156 (N_20156,N_19968,N_19574);
xnor U20157 (N_20157,N_19721,N_19846);
nand U20158 (N_20158,N_19543,N_19997);
nand U20159 (N_20159,N_19792,N_19646);
xor U20160 (N_20160,N_19539,N_19752);
nor U20161 (N_20161,N_19916,N_19725);
nor U20162 (N_20162,N_19873,N_19901);
or U20163 (N_20163,N_19591,N_19980);
xnor U20164 (N_20164,N_19553,N_19596);
nor U20165 (N_20165,N_19729,N_19864);
and U20166 (N_20166,N_19599,N_19710);
or U20167 (N_20167,N_19812,N_19982);
xnor U20168 (N_20168,N_19944,N_19857);
nand U20169 (N_20169,N_19991,N_19551);
xor U20170 (N_20170,N_19511,N_19926);
xnor U20171 (N_20171,N_19989,N_19548);
or U20172 (N_20172,N_19760,N_19840);
and U20173 (N_20173,N_19695,N_19776);
and U20174 (N_20174,N_19748,N_19645);
xor U20175 (N_20175,N_19641,N_19927);
nand U20176 (N_20176,N_19811,N_19608);
and U20177 (N_20177,N_19865,N_19653);
xnor U20178 (N_20178,N_19701,N_19504);
and U20179 (N_20179,N_19718,N_19914);
or U20180 (N_20180,N_19739,N_19976);
nor U20181 (N_20181,N_19979,N_19964);
or U20182 (N_20182,N_19799,N_19871);
or U20183 (N_20183,N_19967,N_19663);
nor U20184 (N_20184,N_19938,N_19533);
nand U20185 (N_20185,N_19961,N_19838);
or U20186 (N_20186,N_19726,N_19912);
xor U20187 (N_20187,N_19869,N_19973);
and U20188 (N_20188,N_19787,N_19638);
and U20189 (N_20189,N_19526,N_19544);
xnor U20190 (N_20190,N_19829,N_19793);
and U20191 (N_20191,N_19660,N_19598);
or U20192 (N_20192,N_19983,N_19805);
xnor U20193 (N_20193,N_19769,N_19527);
nor U20194 (N_20194,N_19885,N_19848);
nor U20195 (N_20195,N_19759,N_19984);
nor U20196 (N_20196,N_19523,N_19779);
and U20197 (N_20197,N_19820,N_19592);
or U20198 (N_20198,N_19940,N_19545);
nor U20199 (N_20199,N_19717,N_19529);
nand U20200 (N_20200,N_19897,N_19888);
nor U20201 (N_20201,N_19819,N_19801);
nor U20202 (N_20202,N_19891,N_19700);
nor U20203 (N_20203,N_19629,N_19797);
nor U20204 (N_20204,N_19903,N_19644);
or U20205 (N_20205,N_19839,N_19972);
nand U20206 (N_20206,N_19524,N_19735);
nor U20207 (N_20207,N_19656,N_19643);
nor U20208 (N_20208,N_19854,N_19568);
or U20209 (N_20209,N_19809,N_19843);
nor U20210 (N_20210,N_19697,N_19847);
or U20211 (N_20211,N_19945,N_19946);
nand U20212 (N_20212,N_19514,N_19837);
or U20213 (N_20213,N_19626,N_19796);
nor U20214 (N_20214,N_19902,N_19817);
nor U20215 (N_20215,N_19740,N_19744);
nor U20216 (N_20216,N_19763,N_19755);
nor U20217 (N_20217,N_19671,N_19501);
xor U20218 (N_20218,N_19880,N_19537);
nor U20219 (N_20219,N_19825,N_19732);
or U20220 (N_20220,N_19911,N_19532);
or U20221 (N_20221,N_19704,N_19731);
nor U20222 (N_20222,N_19715,N_19623);
and U20223 (N_20223,N_19632,N_19804);
or U20224 (N_20224,N_19624,N_19932);
xor U20225 (N_20225,N_19733,N_19557);
or U20226 (N_20226,N_19648,N_19867);
xnor U20227 (N_20227,N_19714,N_19798);
nand U20228 (N_20228,N_19955,N_19507);
nand U20229 (N_20229,N_19684,N_19822);
xor U20230 (N_20230,N_19616,N_19960);
or U20231 (N_20231,N_19642,N_19862);
nand U20232 (N_20232,N_19666,N_19928);
or U20233 (N_20233,N_19676,N_19768);
and U20234 (N_20234,N_19613,N_19657);
nor U20235 (N_20235,N_19627,N_19536);
and U20236 (N_20236,N_19814,N_19882);
nor U20237 (N_20237,N_19951,N_19923);
and U20238 (N_20238,N_19943,N_19709);
nor U20239 (N_20239,N_19818,N_19719);
nor U20240 (N_20240,N_19909,N_19698);
nor U20241 (N_20241,N_19994,N_19628);
and U20242 (N_20242,N_19879,N_19572);
nor U20243 (N_20243,N_19730,N_19934);
xor U20244 (N_20244,N_19929,N_19554);
or U20245 (N_20245,N_19688,N_19894);
nor U20246 (N_20246,N_19868,N_19957);
or U20247 (N_20247,N_19586,N_19842);
nand U20248 (N_20248,N_19977,N_19910);
xnor U20249 (N_20249,N_19517,N_19705);
nand U20250 (N_20250,N_19846,N_19810);
or U20251 (N_20251,N_19616,N_19886);
or U20252 (N_20252,N_19860,N_19771);
or U20253 (N_20253,N_19532,N_19725);
nor U20254 (N_20254,N_19718,N_19907);
xor U20255 (N_20255,N_19639,N_19876);
xor U20256 (N_20256,N_19704,N_19612);
nand U20257 (N_20257,N_19553,N_19976);
or U20258 (N_20258,N_19908,N_19868);
nand U20259 (N_20259,N_19867,N_19798);
xor U20260 (N_20260,N_19711,N_19894);
nand U20261 (N_20261,N_19948,N_19812);
nand U20262 (N_20262,N_19785,N_19600);
nor U20263 (N_20263,N_19750,N_19697);
and U20264 (N_20264,N_19930,N_19824);
or U20265 (N_20265,N_19631,N_19592);
xnor U20266 (N_20266,N_19955,N_19775);
nor U20267 (N_20267,N_19573,N_19949);
and U20268 (N_20268,N_19670,N_19695);
and U20269 (N_20269,N_19889,N_19632);
xor U20270 (N_20270,N_19623,N_19838);
or U20271 (N_20271,N_19958,N_19737);
and U20272 (N_20272,N_19657,N_19999);
nand U20273 (N_20273,N_19516,N_19932);
and U20274 (N_20274,N_19618,N_19693);
or U20275 (N_20275,N_19688,N_19596);
nor U20276 (N_20276,N_19867,N_19742);
and U20277 (N_20277,N_19892,N_19699);
nand U20278 (N_20278,N_19842,N_19641);
and U20279 (N_20279,N_19737,N_19769);
nor U20280 (N_20280,N_19920,N_19765);
nand U20281 (N_20281,N_19655,N_19806);
xnor U20282 (N_20282,N_19818,N_19558);
or U20283 (N_20283,N_19996,N_19593);
nor U20284 (N_20284,N_19603,N_19678);
nor U20285 (N_20285,N_19777,N_19811);
xor U20286 (N_20286,N_19688,N_19733);
nand U20287 (N_20287,N_19876,N_19720);
and U20288 (N_20288,N_19999,N_19918);
or U20289 (N_20289,N_19583,N_19740);
or U20290 (N_20290,N_19857,N_19647);
and U20291 (N_20291,N_19972,N_19587);
or U20292 (N_20292,N_19653,N_19674);
nand U20293 (N_20293,N_19527,N_19584);
nor U20294 (N_20294,N_19778,N_19588);
and U20295 (N_20295,N_19890,N_19621);
nand U20296 (N_20296,N_19758,N_19756);
and U20297 (N_20297,N_19626,N_19739);
and U20298 (N_20298,N_19678,N_19634);
and U20299 (N_20299,N_19528,N_19697);
or U20300 (N_20300,N_19681,N_19988);
nor U20301 (N_20301,N_19934,N_19601);
and U20302 (N_20302,N_19829,N_19624);
or U20303 (N_20303,N_19987,N_19985);
xnor U20304 (N_20304,N_19523,N_19539);
nor U20305 (N_20305,N_19583,N_19575);
xnor U20306 (N_20306,N_19581,N_19768);
or U20307 (N_20307,N_19740,N_19838);
nand U20308 (N_20308,N_19699,N_19818);
nand U20309 (N_20309,N_19655,N_19573);
nor U20310 (N_20310,N_19550,N_19957);
or U20311 (N_20311,N_19929,N_19586);
and U20312 (N_20312,N_19998,N_19974);
or U20313 (N_20313,N_19992,N_19829);
nand U20314 (N_20314,N_19958,N_19576);
nand U20315 (N_20315,N_19831,N_19884);
and U20316 (N_20316,N_19900,N_19598);
and U20317 (N_20317,N_19893,N_19733);
and U20318 (N_20318,N_19619,N_19752);
xnor U20319 (N_20319,N_19827,N_19910);
or U20320 (N_20320,N_19929,N_19823);
or U20321 (N_20321,N_19719,N_19648);
nor U20322 (N_20322,N_19873,N_19806);
or U20323 (N_20323,N_19652,N_19623);
and U20324 (N_20324,N_19864,N_19818);
and U20325 (N_20325,N_19543,N_19502);
nand U20326 (N_20326,N_19735,N_19743);
xor U20327 (N_20327,N_19693,N_19538);
nor U20328 (N_20328,N_19819,N_19628);
and U20329 (N_20329,N_19732,N_19713);
xor U20330 (N_20330,N_19531,N_19666);
and U20331 (N_20331,N_19869,N_19676);
nor U20332 (N_20332,N_19713,N_19625);
or U20333 (N_20333,N_19515,N_19666);
or U20334 (N_20334,N_19703,N_19616);
nor U20335 (N_20335,N_19717,N_19898);
nor U20336 (N_20336,N_19687,N_19798);
and U20337 (N_20337,N_19827,N_19991);
or U20338 (N_20338,N_19530,N_19894);
or U20339 (N_20339,N_19835,N_19975);
nor U20340 (N_20340,N_19523,N_19559);
xor U20341 (N_20341,N_19664,N_19805);
xnor U20342 (N_20342,N_19761,N_19600);
nand U20343 (N_20343,N_19756,N_19731);
nor U20344 (N_20344,N_19851,N_19773);
xor U20345 (N_20345,N_19843,N_19874);
nand U20346 (N_20346,N_19751,N_19876);
xnor U20347 (N_20347,N_19705,N_19831);
or U20348 (N_20348,N_19987,N_19588);
nand U20349 (N_20349,N_19913,N_19857);
nand U20350 (N_20350,N_19869,N_19590);
nor U20351 (N_20351,N_19961,N_19765);
or U20352 (N_20352,N_19828,N_19965);
xnor U20353 (N_20353,N_19543,N_19984);
and U20354 (N_20354,N_19601,N_19562);
and U20355 (N_20355,N_19851,N_19933);
nand U20356 (N_20356,N_19667,N_19536);
xor U20357 (N_20357,N_19706,N_19755);
nor U20358 (N_20358,N_19800,N_19934);
and U20359 (N_20359,N_19815,N_19963);
nand U20360 (N_20360,N_19577,N_19592);
nand U20361 (N_20361,N_19803,N_19823);
and U20362 (N_20362,N_19965,N_19609);
xor U20363 (N_20363,N_19879,N_19570);
nor U20364 (N_20364,N_19658,N_19624);
or U20365 (N_20365,N_19890,N_19580);
or U20366 (N_20366,N_19632,N_19626);
nor U20367 (N_20367,N_19594,N_19559);
and U20368 (N_20368,N_19848,N_19738);
nand U20369 (N_20369,N_19877,N_19606);
xor U20370 (N_20370,N_19877,N_19664);
or U20371 (N_20371,N_19613,N_19829);
nor U20372 (N_20372,N_19918,N_19835);
or U20373 (N_20373,N_19937,N_19729);
xor U20374 (N_20374,N_19707,N_19701);
nor U20375 (N_20375,N_19847,N_19855);
nor U20376 (N_20376,N_19911,N_19750);
nand U20377 (N_20377,N_19836,N_19920);
and U20378 (N_20378,N_19795,N_19770);
and U20379 (N_20379,N_19957,N_19753);
and U20380 (N_20380,N_19916,N_19630);
nand U20381 (N_20381,N_19630,N_19767);
nand U20382 (N_20382,N_19822,N_19610);
xnor U20383 (N_20383,N_19521,N_19540);
nor U20384 (N_20384,N_19562,N_19521);
xor U20385 (N_20385,N_19947,N_19928);
or U20386 (N_20386,N_19788,N_19583);
or U20387 (N_20387,N_19520,N_19984);
xnor U20388 (N_20388,N_19835,N_19787);
or U20389 (N_20389,N_19706,N_19631);
xor U20390 (N_20390,N_19708,N_19646);
or U20391 (N_20391,N_19864,N_19920);
and U20392 (N_20392,N_19675,N_19559);
and U20393 (N_20393,N_19793,N_19671);
or U20394 (N_20394,N_19658,N_19841);
xor U20395 (N_20395,N_19951,N_19617);
xor U20396 (N_20396,N_19742,N_19941);
nand U20397 (N_20397,N_19741,N_19842);
nor U20398 (N_20398,N_19635,N_19608);
nand U20399 (N_20399,N_19780,N_19800);
nor U20400 (N_20400,N_19785,N_19596);
or U20401 (N_20401,N_19952,N_19982);
xor U20402 (N_20402,N_19943,N_19854);
and U20403 (N_20403,N_19591,N_19842);
nor U20404 (N_20404,N_19877,N_19941);
and U20405 (N_20405,N_19521,N_19671);
xor U20406 (N_20406,N_19651,N_19825);
and U20407 (N_20407,N_19788,N_19574);
nand U20408 (N_20408,N_19854,N_19919);
nand U20409 (N_20409,N_19856,N_19996);
and U20410 (N_20410,N_19773,N_19970);
nor U20411 (N_20411,N_19956,N_19771);
and U20412 (N_20412,N_19936,N_19747);
and U20413 (N_20413,N_19795,N_19896);
nor U20414 (N_20414,N_19579,N_19831);
xnor U20415 (N_20415,N_19867,N_19691);
nand U20416 (N_20416,N_19907,N_19542);
and U20417 (N_20417,N_19832,N_19610);
nor U20418 (N_20418,N_19837,N_19613);
and U20419 (N_20419,N_19875,N_19547);
and U20420 (N_20420,N_19757,N_19988);
nand U20421 (N_20421,N_19973,N_19573);
or U20422 (N_20422,N_19605,N_19603);
nor U20423 (N_20423,N_19979,N_19995);
and U20424 (N_20424,N_19848,N_19901);
xor U20425 (N_20425,N_19606,N_19950);
xor U20426 (N_20426,N_19907,N_19990);
nor U20427 (N_20427,N_19815,N_19540);
xor U20428 (N_20428,N_19535,N_19820);
xor U20429 (N_20429,N_19565,N_19820);
xor U20430 (N_20430,N_19986,N_19588);
nand U20431 (N_20431,N_19840,N_19624);
and U20432 (N_20432,N_19501,N_19540);
nand U20433 (N_20433,N_19540,N_19871);
and U20434 (N_20434,N_19505,N_19610);
or U20435 (N_20435,N_19893,N_19885);
nor U20436 (N_20436,N_19536,N_19748);
and U20437 (N_20437,N_19683,N_19582);
nor U20438 (N_20438,N_19750,N_19964);
or U20439 (N_20439,N_19586,N_19505);
or U20440 (N_20440,N_19918,N_19799);
and U20441 (N_20441,N_19533,N_19727);
nor U20442 (N_20442,N_19979,N_19800);
nand U20443 (N_20443,N_19540,N_19849);
nor U20444 (N_20444,N_19689,N_19683);
and U20445 (N_20445,N_19596,N_19915);
nand U20446 (N_20446,N_19888,N_19946);
nand U20447 (N_20447,N_19696,N_19628);
and U20448 (N_20448,N_19500,N_19570);
nand U20449 (N_20449,N_19928,N_19883);
and U20450 (N_20450,N_19837,N_19806);
nand U20451 (N_20451,N_19852,N_19616);
or U20452 (N_20452,N_19508,N_19587);
and U20453 (N_20453,N_19759,N_19646);
nor U20454 (N_20454,N_19643,N_19548);
nor U20455 (N_20455,N_19912,N_19572);
nor U20456 (N_20456,N_19872,N_19733);
nor U20457 (N_20457,N_19874,N_19688);
xnor U20458 (N_20458,N_19781,N_19837);
nor U20459 (N_20459,N_19883,N_19988);
nand U20460 (N_20460,N_19589,N_19558);
and U20461 (N_20461,N_19867,N_19598);
nand U20462 (N_20462,N_19566,N_19676);
or U20463 (N_20463,N_19705,N_19569);
nand U20464 (N_20464,N_19606,N_19632);
or U20465 (N_20465,N_19993,N_19669);
xnor U20466 (N_20466,N_19794,N_19762);
nor U20467 (N_20467,N_19695,N_19951);
xor U20468 (N_20468,N_19539,N_19806);
nor U20469 (N_20469,N_19561,N_19612);
nor U20470 (N_20470,N_19988,N_19668);
and U20471 (N_20471,N_19705,N_19590);
or U20472 (N_20472,N_19923,N_19514);
nand U20473 (N_20473,N_19740,N_19876);
nand U20474 (N_20474,N_19507,N_19930);
nand U20475 (N_20475,N_19997,N_19676);
nand U20476 (N_20476,N_19869,N_19749);
xor U20477 (N_20477,N_19824,N_19543);
or U20478 (N_20478,N_19946,N_19700);
nand U20479 (N_20479,N_19558,N_19741);
nand U20480 (N_20480,N_19757,N_19531);
or U20481 (N_20481,N_19533,N_19531);
xor U20482 (N_20482,N_19580,N_19660);
or U20483 (N_20483,N_19560,N_19847);
and U20484 (N_20484,N_19849,N_19844);
and U20485 (N_20485,N_19530,N_19923);
xnor U20486 (N_20486,N_19917,N_19597);
nor U20487 (N_20487,N_19695,N_19983);
nor U20488 (N_20488,N_19518,N_19858);
xnor U20489 (N_20489,N_19862,N_19711);
nand U20490 (N_20490,N_19633,N_19513);
nor U20491 (N_20491,N_19622,N_19692);
and U20492 (N_20492,N_19507,N_19555);
xnor U20493 (N_20493,N_19646,N_19805);
and U20494 (N_20494,N_19709,N_19673);
or U20495 (N_20495,N_19705,N_19969);
or U20496 (N_20496,N_19597,N_19515);
or U20497 (N_20497,N_19939,N_19517);
xor U20498 (N_20498,N_19878,N_19551);
nor U20499 (N_20499,N_19939,N_19679);
or U20500 (N_20500,N_20287,N_20099);
xnor U20501 (N_20501,N_20059,N_20441);
or U20502 (N_20502,N_20114,N_20104);
or U20503 (N_20503,N_20466,N_20291);
xnor U20504 (N_20504,N_20437,N_20179);
xor U20505 (N_20505,N_20455,N_20365);
nand U20506 (N_20506,N_20393,N_20141);
nor U20507 (N_20507,N_20159,N_20269);
nor U20508 (N_20508,N_20226,N_20169);
or U20509 (N_20509,N_20336,N_20371);
and U20510 (N_20510,N_20003,N_20325);
nand U20511 (N_20511,N_20115,N_20354);
nand U20512 (N_20512,N_20264,N_20407);
or U20513 (N_20513,N_20488,N_20357);
nand U20514 (N_20514,N_20000,N_20185);
nand U20515 (N_20515,N_20487,N_20001);
xor U20516 (N_20516,N_20014,N_20206);
nand U20517 (N_20517,N_20318,N_20465);
nand U20518 (N_20518,N_20058,N_20095);
or U20519 (N_20519,N_20043,N_20424);
and U20520 (N_20520,N_20372,N_20327);
xnor U20521 (N_20521,N_20235,N_20148);
nor U20522 (N_20522,N_20335,N_20237);
or U20523 (N_20523,N_20121,N_20499);
nor U20524 (N_20524,N_20019,N_20244);
xor U20525 (N_20525,N_20385,N_20219);
or U20526 (N_20526,N_20435,N_20026);
or U20527 (N_20527,N_20170,N_20038);
nor U20528 (N_20528,N_20176,N_20066);
nand U20529 (N_20529,N_20078,N_20012);
xor U20530 (N_20530,N_20129,N_20163);
xor U20531 (N_20531,N_20476,N_20212);
or U20532 (N_20532,N_20109,N_20173);
and U20533 (N_20533,N_20032,N_20098);
nand U20534 (N_20534,N_20234,N_20259);
xnor U20535 (N_20535,N_20306,N_20414);
nor U20536 (N_20536,N_20168,N_20120);
or U20537 (N_20537,N_20057,N_20417);
nor U20538 (N_20538,N_20086,N_20343);
xnor U20539 (N_20539,N_20134,N_20381);
or U20540 (N_20540,N_20440,N_20101);
or U20541 (N_20541,N_20268,N_20194);
or U20542 (N_20542,N_20198,N_20221);
nand U20543 (N_20543,N_20353,N_20274);
and U20544 (N_20544,N_20425,N_20421);
nor U20545 (N_20545,N_20412,N_20410);
or U20546 (N_20546,N_20482,N_20184);
xor U20547 (N_20547,N_20303,N_20160);
nor U20548 (N_20548,N_20413,N_20047);
and U20549 (N_20549,N_20061,N_20054);
xnor U20550 (N_20550,N_20345,N_20279);
xnor U20551 (N_20551,N_20239,N_20124);
nand U20552 (N_20552,N_20228,N_20128);
and U20553 (N_20553,N_20192,N_20069);
nor U20554 (N_20554,N_20207,N_20278);
nand U20555 (N_20555,N_20085,N_20055);
xor U20556 (N_20556,N_20052,N_20215);
nor U20557 (N_20557,N_20208,N_20131);
or U20558 (N_20558,N_20222,N_20415);
nand U20559 (N_20559,N_20007,N_20009);
and U20560 (N_20560,N_20399,N_20039);
xor U20561 (N_20561,N_20387,N_20458);
nor U20562 (N_20562,N_20250,N_20351);
xor U20563 (N_20563,N_20213,N_20356);
xnor U20564 (N_20564,N_20094,N_20119);
or U20565 (N_20565,N_20472,N_20113);
xnor U20566 (N_20566,N_20147,N_20401);
xor U20567 (N_20567,N_20097,N_20355);
nor U20568 (N_20568,N_20132,N_20041);
nand U20569 (N_20569,N_20186,N_20090);
nand U20570 (N_20570,N_20460,N_20200);
or U20571 (N_20571,N_20161,N_20311);
and U20572 (N_20572,N_20375,N_20408);
nor U20573 (N_20573,N_20158,N_20008);
nor U20574 (N_20574,N_20349,N_20048);
nand U20575 (N_20575,N_20233,N_20155);
or U20576 (N_20576,N_20252,N_20304);
and U20577 (N_20577,N_20439,N_20056);
and U20578 (N_20578,N_20175,N_20493);
and U20579 (N_20579,N_20416,N_20309);
xnor U20580 (N_20580,N_20072,N_20263);
or U20581 (N_20581,N_20367,N_20073);
xnor U20582 (N_20582,N_20396,N_20293);
or U20583 (N_20583,N_20108,N_20151);
and U20584 (N_20584,N_20145,N_20117);
or U20585 (N_20585,N_20266,N_20400);
nor U20586 (N_20586,N_20203,N_20130);
or U20587 (N_20587,N_20436,N_20299);
and U20588 (N_20588,N_20395,N_20316);
nand U20589 (N_20589,N_20199,N_20190);
and U20590 (N_20590,N_20352,N_20285);
and U20591 (N_20591,N_20204,N_20020);
nand U20592 (N_20592,N_20388,N_20404);
nor U20593 (N_20593,N_20459,N_20081);
nor U20594 (N_20594,N_20143,N_20380);
nor U20595 (N_20595,N_20305,N_20050);
or U20596 (N_20596,N_20005,N_20374);
nand U20597 (N_20597,N_20489,N_20286);
nand U20598 (N_20598,N_20178,N_20107);
and U20599 (N_20599,N_20432,N_20247);
xor U20600 (N_20600,N_20284,N_20331);
and U20601 (N_20601,N_20112,N_20110);
xor U20602 (N_20602,N_20308,N_20260);
and U20603 (N_20603,N_20373,N_20321);
nand U20604 (N_20604,N_20338,N_20033);
or U20605 (N_20605,N_20002,N_20150);
xnor U20606 (N_20606,N_20497,N_20246);
or U20607 (N_20607,N_20288,N_20491);
nand U20608 (N_20608,N_20411,N_20063);
xor U20609 (N_20609,N_20133,N_20093);
xnor U20610 (N_20610,N_20368,N_20049);
nor U20611 (N_20611,N_20486,N_20232);
and U20612 (N_20612,N_20358,N_20273);
xnor U20613 (N_20613,N_20453,N_20270);
and U20614 (N_20614,N_20477,N_20138);
and U20615 (N_20615,N_20210,N_20422);
nor U20616 (N_20616,N_20484,N_20485);
xnor U20617 (N_20617,N_20146,N_20323);
nand U20618 (N_20618,N_20347,N_20167);
nor U20619 (N_20619,N_20181,N_20378);
and U20620 (N_20620,N_20156,N_20241);
or U20621 (N_20621,N_20340,N_20201);
nor U20622 (N_20622,N_20433,N_20088);
nand U20623 (N_20623,N_20272,N_20289);
xor U20624 (N_20624,N_20363,N_20330);
nand U20625 (N_20625,N_20251,N_20312);
and U20626 (N_20626,N_20123,N_20454);
nor U20627 (N_20627,N_20322,N_20195);
and U20628 (N_20628,N_20125,N_20282);
nand U20629 (N_20629,N_20403,N_20448);
xor U20630 (N_20630,N_20220,N_20447);
xor U20631 (N_20631,N_20070,N_20202);
nand U20632 (N_20632,N_20089,N_20255);
and U20633 (N_20633,N_20297,N_20036);
xor U20634 (N_20634,N_20467,N_20080);
xnor U20635 (N_20635,N_20314,N_20051);
nand U20636 (N_20636,N_20024,N_20118);
or U20637 (N_20637,N_20258,N_20328);
nand U20638 (N_20638,N_20209,N_20267);
nor U20639 (N_20639,N_20361,N_20025);
nand U20640 (N_20640,N_20294,N_20397);
or U20641 (N_20641,N_20077,N_20341);
nand U20642 (N_20642,N_20083,N_20382);
nor U20643 (N_20643,N_20225,N_20344);
nor U20644 (N_20644,N_20450,N_20139);
and U20645 (N_20645,N_20253,N_20182);
and U20646 (N_20646,N_20216,N_20479);
and U20647 (N_20647,N_20394,N_20122);
and U20648 (N_20648,N_20362,N_20045);
nand U20649 (N_20649,N_20197,N_20423);
nor U20650 (N_20650,N_20494,N_20295);
nor U20651 (N_20651,N_20370,N_20172);
nand U20652 (N_20652,N_20281,N_20075);
nand U20653 (N_20653,N_20383,N_20135);
nand U20654 (N_20654,N_20214,N_20030);
xor U20655 (N_20655,N_20339,N_20006);
and U20656 (N_20656,N_20392,N_20230);
nor U20657 (N_20657,N_20369,N_20496);
and U20658 (N_20658,N_20062,N_20211);
and U20659 (N_20659,N_20153,N_20154);
xnor U20660 (N_20660,N_20256,N_20449);
xnor U20661 (N_20661,N_20060,N_20067);
or U20662 (N_20662,N_20010,N_20189);
or U20663 (N_20663,N_20096,N_20438);
xnor U20664 (N_20664,N_20142,N_20348);
xnor U20665 (N_20665,N_20034,N_20224);
nand U20666 (N_20666,N_20102,N_20280);
xnor U20667 (N_20667,N_20434,N_20171);
or U20668 (N_20668,N_20475,N_20042);
or U20669 (N_20669,N_20461,N_20027);
and U20670 (N_20670,N_20324,N_20428);
nand U20671 (N_20671,N_20326,N_20205);
and U20672 (N_20672,N_20366,N_20164);
or U20673 (N_20673,N_20473,N_20180);
and U20674 (N_20674,N_20332,N_20064);
and U20675 (N_20675,N_20329,N_20087);
nand U20676 (N_20676,N_20126,N_20457);
and U20677 (N_20677,N_20405,N_20290);
nor U20678 (N_20678,N_20333,N_20334);
xnor U20679 (N_20679,N_20152,N_20053);
or U20680 (N_20680,N_20307,N_20227);
xor U20681 (N_20681,N_20337,N_20359);
or U20682 (N_20682,N_20320,N_20031);
and U20683 (N_20683,N_20243,N_20013);
nor U20684 (N_20684,N_20174,N_20071);
xnor U20685 (N_20685,N_20470,N_20011);
nor U20686 (N_20686,N_20111,N_20229);
xnor U20687 (N_20687,N_20183,N_20218);
nor U20688 (N_20688,N_20409,N_20379);
or U20689 (N_20689,N_20313,N_20445);
or U20690 (N_20690,N_20474,N_20376);
xnor U20691 (N_20691,N_20296,N_20495);
or U20692 (N_20692,N_20028,N_20136);
and U20693 (N_20693,N_20217,N_20350);
xnor U20694 (N_20694,N_20074,N_20100);
and U20695 (N_20695,N_20490,N_20157);
nand U20696 (N_20696,N_20044,N_20301);
xor U20697 (N_20697,N_20018,N_20223);
nor U20698 (N_20698,N_20236,N_20106);
and U20699 (N_20699,N_20193,N_20364);
nor U20700 (N_20700,N_20127,N_20406);
and U20701 (N_20701,N_20137,N_20426);
xor U20702 (N_20702,N_20319,N_20248);
and U20703 (N_20703,N_20022,N_20261);
xor U20704 (N_20704,N_20249,N_20276);
or U20705 (N_20705,N_20238,N_20177);
and U20706 (N_20706,N_20079,N_20300);
or U20707 (N_20707,N_20016,N_20389);
or U20708 (N_20708,N_20188,N_20462);
or U20709 (N_20709,N_20076,N_20469);
nand U20710 (N_20710,N_20166,N_20398);
or U20711 (N_20711,N_20464,N_20046);
or U20712 (N_20712,N_20084,N_20283);
or U20713 (N_20713,N_20430,N_20390);
xor U20714 (N_20714,N_20443,N_20035);
xnor U20715 (N_20715,N_20446,N_20360);
and U20716 (N_20716,N_20342,N_20480);
nor U20717 (N_20717,N_20242,N_20015);
nand U20718 (N_20718,N_20140,N_20481);
or U20719 (N_20719,N_20292,N_20029);
nand U20720 (N_20720,N_20245,N_20254);
xor U20721 (N_20721,N_20240,N_20471);
nand U20722 (N_20722,N_20040,N_20105);
nand U20723 (N_20723,N_20191,N_20420);
nor U20724 (N_20724,N_20265,N_20456);
or U20725 (N_20725,N_20451,N_20262);
xor U20726 (N_20726,N_20231,N_20429);
nor U20727 (N_20727,N_20442,N_20092);
and U20728 (N_20728,N_20452,N_20196);
xor U20729 (N_20729,N_20298,N_20021);
and U20730 (N_20730,N_20431,N_20144);
nor U20731 (N_20731,N_20427,N_20483);
or U20732 (N_20732,N_20498,N_20384);
xnor U20733 (N_20733,N_20257,N_20346);
nand U20734 (N_20734,N_20004,N_20103);
xor U20735 (N_20735,N_20277,N_20386);
or U20736 (N_20736,N_20317,N_20418);
or U20737 (N_20737,N_20017,N_20065);
and U20738 (N_20738,N_20444,N_20037);
and U20739 (N_20739,N_20275,N_20419);
nand U20740 (N_20740,N_20162,N_20468);
and U20741 (N_20741,N_20082,N_20302);
nand U20742 (N_20742,N_20165,N_20463);
nor U20743 (N_20743,N_20402,N_20091);
or U20744 (N_20744,N_20149,N_20116);
nor U20745 (N_20745,N_20492,N_20271);
xor U20746 (N_20746,N_20377,N_20068);
xnor U20747 (N_20747,N_20315,N_20478);
nand U20748 (N_20748,N_20187,N_20391);
xnor U20749 (N_20749,N_20023,N_20310);
xnor U20750 (N_20750,N_20360,N_20052);
nand U20751 (N_20751,N_20082,N_20209);
nand U20752 (N_20752,N_20401,N_20013);
or U20753 (N_20753,N_20112,N_20121);
or U20754 (N_20754,N_20232,N_20326);
xnor U20755 (N_20755,N_20290,N_20168);
xnor U20756 (N_20756,N_20310,N_20022);
xor U20757 (N_20757,N_20380,N_20027);
nand U20758 (N_20758,N_20431,N_20100);
nor U20759 (N_20759,N_20392,N_20087);
nand U20760 (N_20760,N_20385,N_20435);
nand U20761 (N_20761,N_20347,N_20331);
nand U20762 (N_20762,N_20463,N_20150);
nor U20763 (N_20763,N_20116,N_20348);
or U20764 (N_20764,N_20401,N_20406);
nand U20765 (N_20765,N_20217,N_20486);
or U20766 (N_20766,N_20460,N_20097);
xor U20767 (N_20767,N_20076,N_20280);
or U20768 (N_20768,N_20027,N_20292);
and U20769 (N_20769,N_20135,N_20140);
xnor U20770 (N_20770,N_20479,N_20245);
nor U20771 (N_20771,N_20164,N_20424);
xnor U20772 (N_20772,N_20247,N_20100);
or U20773 (N_20773,N_20236,N_20289);
and U20774 (N_20774,N_20247,N_20358);
or U20775 (N_20775,N_20481,N_20289);
xor U20776 (N_20776,N_20483,N_20226);
or U20777 (N_20777,N_20049,N_20401);
or U20778 (N_20778,N_20482,N_20164);
or U20779 (N_20779,N_20011,N_20147);
or U20780 (N_20780,N_20289,N_20119);
nand U20781 (N_20781,N_20343,N_20344);
xnor U20782 (N_20782,N_20092,N_20025);
or U20783 (N_20783,N_20175,N_20212);
and U20784 (N_20784,N_20042,N_20195);
nor U20785 (N_20785,N_20103,N_20085);
xor U20786 (N_20786,N_20471,N_20483);
nand U20787 (N_20787,N_20424,N_20031);
or U20788 (N_20788,N_20202,N_20151);
and U20789 (N_20789,N_20013,N_20496);
nand U20790 (N_20790,N_20344,N_20444);
xnor U20791 (N_20791,N_20380,N_20100);
xor U20792 (N_20792,N_20236,N_20024);
and U20793 (N_20793,N_20245,N_20426);
and U20794 (N_20794,N_20345,N_20312);
nand U20795 (N_20795,N_20262,N_20333);
or U20796 (N_20796,N_20445,N_20479);
or U20797 (N_20797,N_20249,N_20058);
nor U20798 (N_20798,N_20380,N_20279);
nand U20799 (N_20799,N_20174,N_20224);
xnor U20800 (N_20800,N_20139,N_20231);
xnor U20801 (N_20801,N_20116,N_20029);
xor U20802 (N_20802,N_20486,N_20214);
xor U20803 (N_20803,N_20172,N_20236);
nand U20804 (N_20804,N_20005,N_20187);
xnor U20805 (N_20805,N_20467,N_20233);
nand U20806 (N_20806,N_20218,N_20352);
or U20807 (N_20807,N_20012,N_20171);
nand U20808 (N_20808,N_20453,N_20273);
nor U20809 (N_20809,N_20067,N_20132);
xor U20810 (N_20810,N_20028,N_20492);
nand U20811 (N_20811,N_20499,N_20470);
xnor U20812 (N_20812,N_20335,N_20229);
nand U20813 (N_20813,N_20200,N_20269);
nand U20814 (N_20814,N_20058,N_20240);
or U20815 (N_20815,N_20131,N_20145);
xor U20816 (N_20816,N_20134,N_20429);
xnor U20817 (N_20817,N_20460,N_20204);
and U20818 (N_20818,N_20034,N_20447);
xor U20819 (N_20819,N_20475,N_20441);
nor U20820 (N_20820,N_20085,N_20346);
nand U20821 (N_20821,N_20426,N_20311);
nand U20822 (N_20822,N_20169,N_20490);
and U20823 (N_20823,N_20147,N_20425);
and U20824 (N_20824,N_20108,N_20043);
nand U20825 (N_20825,N_20329,N_20077);
or U20826 (N_20826,N_20273,N_20080);
nand U20827 (N_20827,N_20005,N_20062);
nor U20828 (N_20828,N_20388,N_20246);
nand U20829 (N_20829,N_20413,N_20360);
or U20830 (N_20830,N_20404,N_20041);
nor U20831 (N_20831,N_20177,N_20192);
or U20832 (N_20832,N_20445,N_20265);
nor U20833 (N_20833,N_20208,N_20099);
xnor U20834 (N_20834,N_20140,N_20007);
xor U20835 (N_20835,N_20451,N_20364);
xnor U20836 (N_20836,N_20297,N_20366);
nor U20837 (N_20837,N_20061,N_20297);
nor U20838 (N_20838,N_20017,N_20022);
or U20839 (N_20839,N_20034,N_20302);
nand U20840 (N_20840,N_20251,N_20314);
xor U20841 (N_20841,N_20181,N_20396);
nand U20842 (N_20842,N_20210,N_20190);
or U20843 (N_20843,N_20345,N_20407);
nor U20844 (N_20844,N_20316,N_20088);
nor U20845 (N_20845,N_20453,N_20004);
and U20846 (N_20846,N_20468,N_20412);
nor U20847 (N_20847,N_20136,N_20073);
and U20848 (N_20848,N_20203,N_20371);
nor U20849 (N_20849,N_20144,N_20445);
or U20850 (N_20850,N_20448,N_20204);
nor U20851 (N_20851,N_20223,N_20284);
and U20852 (N_20852,N_20395,N_20189);
nand U20853 (N_20853,N_20197,N_20149);
nand U20854 (N_20854,N_20071,N_20074);
and U20855 (N_20855,N_20433,N_20234);
or U20856 (N_20856,N_20045,N_20154);
xor U20857 (N_20857,N_20044,N_20395);
and U20858 (N_20858,N_20429,N_20117);
and U20859 (N_20859,N_20228,N_20304);
nand U20860 (N_20860,N_20429,N_20490);
nand U20861 (N_20861,N_20145,N_20103);
or U20862 (N_20862,N_20391,N_20156);
and U20863 (N_20863,N_20400,N_20307);
xnor U20864 (N_20864,N_20355,N_20012);
xnor U20865 (N_20865,N_20211,N_20233);
nand U20866 (N_20866,N_20174,N_20054);
nand U20867 (N_20867,N_20336,N_20497);
xor U20868 (N_20868,N_20020,N_20349);
nand U20869 (N_20869,N_20325,N_20490);
and U20870 (N_20870,N_20321,N_20161);
and U20871 (N_20871,N_20141,N_20033);
and U20872 (N_20872,N_20416,N_20168);
xor U20873 (N_20873,N_20298,N_20433);
or U20874 (N_20874,N_20323,N_20248);
or U20875 (N_20875,N_20099,N_20082);
and U20876 (N_20876,N_20412,N_20382);
nand U20877 (N_20877,N_20045,N_20125);
and U20878 (N_20878,N_20052,N_20129);
or U20879 (N_20879,N_20491,N_20369);
nand U20880 (N_20880,N_20459,N_20432);
nand U20881 (N_20881,N_20055,N_20417);
nor U20882 (N_20882,N_20297,N_20403);
xnor U20883 (N_20883,N_20245,N_20017);
nand U20884 (N_20884,N_20242,N_20220);
nand U20885 (N_20885,N_20045,N_20040);
nor U20886 (N_20886,N_20142,N_20147);
nand U20887 (N_20887,N_20057,N_20028);
and U20888 (N_20888,N_20342,N_20217);
or U20889 (N_20889,N_20059,N_20231);
and U20890 (N_20890,N_20243,N_20114);
nor U20891 (N_20891,N_20044,N_20116);
nor U20892 (N_20892,N_20014,N_20204);
xnor U20893 (N_20893,N_20428,N_20220);
xnor U20894 (N_20894,N_20266,N_20175);
xor U20895 (N_20895,N_20467,N_20235);
xor U20896 (N_20896,N_20474,N_20211);
or U20897 (N_20897,N_20068,N_20049);
or U20898 (N_20898,N_20219,N_20427);
nor U20899 (N_20899,N_20413,N_20486);
and U20900 (N_20900,N_20126,N_20480);
nand U20901 (N_20901,N_20346,N_20433);
or U20902 (N_20902,N_20000,N_20157);
or U20903 (N_20903,N_20494,N_20387);
nand U20904 (N_20904,N_20112,N_20408);
or U20905 (N_20905,N_20171,N_20444);
xor U20906 (N_20906,N_20047,N_20184);
and U20907 (N_20907,N_20476,N_20141);
or U20908 (N_20908,N_20297,N_20029);
nor U20909 (N_20909,N_20042,N_20000);
or U20910 (N_20910,N_20480,N_20344);
and U20911 (N_20911,N_20284,N_20161);
xor U20912 (N_20912,N_20279,N_20334);
or U20913 (N_20913,N_20000,N_20365);
nor U20914 (N_20914,N_20408,N_20345);
or U20915 (N_20915,N_20118,N_20367);
xor U20916 (N_20916,N_20294,N_20367);
xor U20917 (N_20917,N_20360,N_20194);
nor U20918 (N_20918,N_20207,N_20044);
xnor U20919 (N_20919,N_20208,N_20181);
nor U20920 (N_20920,N_20015,N_20445);
nor U20921 (N_20921,N_20443,N_20020);
or U20922 (N_20922,N_20158,N_20405);
and U20923 (N_20923,N_20274,N_20086);
nor U20924 (N_20924,N_20495,N_20351);
nand U20925 (N_20925,N_20384,N_20197);
or U20926 (N_20926,N_20428,N_20486);
nor U20927 (N_20927,N_20323,N_20091);
nand U20928 (N_20928,N_20413,N_20292);
or U20929 (N_20929,N_20313,N_20368);
xor U20930 (N_20930,N_20226,N_20216);
and U20931 (N_20931,N_20129,N_20485);
or U20932 (N_20932,N_20037,N_20119);
nor U20933 (N_20933,N_20492,N_20197);
nand U20934 (N_20934,N_20271,N_20048);
nor U20935 (N_20935,N_20427,N_20279);
nand U20936 (N_20936,N_20161,N_20328);
or U20937 (N_20937,N_20004,N_20447);
or U20938 (N_20938,N_20068,N_20194);
nor U20939 (N_20939,N_20053,N_20344);
or U20940 (N_20940,N_20472,N_20269);
or U20941 (N_20941,N_20446,N_20244);
nor U20942 (N_20942,N_20241,N_20440);
or U20943 (N_20943,N_20077,N_20255);
and U20944 (N_20944,N_20416,N_20066);
or U20945 (N_20945,N_20050,N_20319);
nand U20946 (N_20946,N_20434,N_20428);
nor U20947 (N_20947,N_20152,N_20484);
xnor U20948 (N_20948,N_20412,N_20023);
or U20949 (N_20949,N_20348,N_20266);
and U20950 (N_20950,N_20241,N_20006);
and U20951 (N_20951,N_20002,N_20134);
nor U20952 (N_20952,N_20068,N_20015);
and U20953 (N_20953,N_20498,N_20460);
nor U20954 (N_20954,N_20048,N_20337);
nand U20955 (N_20955,N_20343,N_20208);
and U20956 (N_20956,N_20198,N_20056);
nor U20957 (N_20957,N_20422,N_20145);
nor U20958 (N_20958,N_20392,N_20455);
and U20959 (N_20959,N_20186,N_20107);
xnor U20960 (N_20960,N_20011,N_20092);
and U20961 (N_20961,N_20490,N_20329);
and U20962 (N_20962,N_20050,N_20061);
xor U20963 (N_20963,N_20089,N_20159);
and U20964 (N_20964,N_20354,N_20233);
xor U20965 (N_20965,N_20467,N_20066);
nand U20966 (N_20966,N_20280,N_20032);
xnor U20967 (N_20967,N_20486,N_20446);
and U20968 (N_20968,N_20014,N_20047);
nor U20969 (N_20969,N_20311,N_20057);
nand U20970 (N_20970,N_20365,N_20267);
nand U20971 (N_20971,N_20128,N_20458);
xnor U20972 (N_20972,N_20086,N_20377);
nor U20973 (N_20973,N_20002,N_20144);
xor U20974 (N_20974,N_20485,N_20034);
or U20975 (N_20975,N_20309,N_20490);
nor U20976 (N_20976,N_20077,N_20229);
xnor U20977 (N_20977,N_20324,N_20196);
nand U20978 (N_20978,N_20447,N_20231);
or U20979 (N_20979,N_20075,N_20449);
and U20980 (N_20980,N_20279,N_20213);
or U20981 (N_20981,N_20245,N_20383);
or U20982 (N_20982,N_20334,N_20253);
xnor U20983 (N_20983,N_20365,N_20178);
xnor U20984 (N_20984,N_20452,N_20082);
nor U20985 (N_20985,N_20071,N_20440);
nor U20986 (N_20986,N_20171,N_20069);
or U20987 (N_20987,N_20313,N_20488);
or U20988 (N_20988,N_20002,N_20242);
nand U20989 (N_20989,N_20327,N_20494);
or U20990 (N_20990,N_20368,N_20083);
nor U20991 (N_20991,N_20340,N_20100);
nand U20992 (N_20992,N_20220,N_20120);
nor U20993 (N_20993,N_20221,N_20240);
or U20994 (N_20994,N_20104,N_20428);
nor U20995 (N_20995,N_20443,N_20347);
nor U20996 (N_20996,N_20129,N_20355);
xnor U20997 (N_20997,N_20494,N_20191);
nor U20998 (N_20998,N_20495,N_20475);
or U20999 (N_20999,N_20043,N_20050);
or U21000 (N_21000,N_20820,N_20702);
and U21001 (N_21001,N_20832,N_20667);
xor U21002 (N_21002,N_20552,N_20573);
nor U21003 (N_21003,N_20612,N_20668);
or U21004 (N_21004,N_20676,N_20823);
or U21005 (N_21005,N_20590,N_20642);
nor U21006 (N_21006,N_20703,N_20587);
xnor U21007 (N_21007,N_20885,N_20530);
nor U21008 (N_21008,N_20718,N_20829);
or U21009 (N_21009,N_20792,N_20958);
or U21010 (N_21010,N_20911,N_20834);
and U21011 (N_21011,N_20582,N_20806);
nand U21012 (N_21012,N_20564,N_20881);
and U21013 (N_21013,N_20910,N_20981);
nor U21014 (N_21014,N_20729,N_20571);
and U21015 (N_21015,N_20923,N_20796);
and U21016 (N_21016,N_20860,N_20560);
and U21017 (N_21017,N_20713,N_20887);
nand U21018 (N_21018,N_20840,N_20535);
or U21019 (N_21019,N_20558,N_20515);
nand U21020 (N_21020,N_20540,N_20528);
or U21021 (N_21021,N_20782,N_20960);
nor U21022 (N_21022,N_20996,N_20882);
nand U21023 (N_21023,N_20733,N_20949);
or U21024 (N_21024,N_20870,N_20610);
nor U21025 (N_21025,N_20943,N_20915);
or U21026 (N_21026,N_20921,N_20811);
nand U21027 (N_21027,N_20987,N_20767);
nor U21028 (N_21028,N_20762,N_20594);
and U21029 (N_21029,N_20504,N_20867);
nand U21030 (N_21030,N_20719,N_20776);
xnor U21031 (N_21031,N_20717,N_20576);
and U21032 (N_21032,N_20722,N_20939);
and U21033 (N_21033,N_20875,N_20744);
or U21034 (N_21034,N_20848,N_20505);
and U21035 (N_21035,N_20751,N_20933);
xnor U21036 (N_21036,N_20974,N_20685);
nor U21037 (N_21037,N_20740,N_20756);
nand U21038 (N_21038,N_20924,N_20636);
and U21039 (N_21039,N_20514,N_20798);
or U21040 (N_21040,N_20565,N_20866);
and U21041 (N_21041,N_20544,N_20682);
and U21042 (N_21042,N_20659,N_20691);
nor U21043 (N_21043,N_20853,N_20844);
nor U21044 (N_21044,N_20927,N_20764);
nor U21045 (N_21045,N_20695,N_20510);
nor U21046 (N_21046,N_20584,N_20634);
nor U21047 (N_21047,N_20539,N_20783);
nor U21048 (N_21048,N_20519,N_20613);
or U21049 (N_21049,N_20543,N_20684);
xnor U21050 (N_21050,N_20680,N_20726);
or U21051 (N_21051,N_20581,N_20843);
and U21052 (N_21052,N_20556,N_20794);
nor U21053 (N_21053,N_20900,N_20517);
or U21054 (N_21054,N_20561,N_20553);
and U21055 (N_21055,N_20889,N_20688);
or U21056 (N_21056,N_20800,N_20706);
nor U21057 (N_21057,N_20745,N_20502);
nor U21058 (N_21058,N_20847,N_20654);
nor U21059 (N_21059,N_20503,N_20616);
and U21060 (N_21060,N_20966,N_20932);
nor U21061 (N_21061,N_20896,N_20942);
xor U21062 (N_21062,N_20777,N_20748);
and U21063 (N_21063,N_20550,N_20940);
xor U21064 (N_21064,N_20786,N_20652);
nor U21065 (N_21065,N_20724,N_20791);
or U21066 (N_21066,N_20577,N_20611);
nand U21067 (N_21067,N_20670,N_20524);
nor U21068 (N_21068,N_20961,N_20934);
xnor U21069 (N_21069,N_20700,N_20529);
nor U21070 (N_21070,N_20708,N_20772);
nor U21071 (N_21071,N_20959,N_20557);
xor U21072 (N_21072,N_20980,N_20880);
nor U21073 (N_21073,N_20647,N_20648);
or U21074 (N_21074,N_20818,N_20809);
nor U21075 (N_21075,N_20917,N_20998);
xor U21076 (N_21076,N_20973,N_20775);
and U21077 (N_21077,N_20780,N_20689);
nor U21078 (N_21078,N_20597,N_20827);
nor U21079 (N_21079,N_20928,N_20984);
or U21080 (N_21080,N_20570,N_20603);
and U21081 (N_21081,N_20891,N_20549);
xor U21082 (N_21082,N_20629,N_20954);
and U21083 (N_21083,N_20578,N_20817);
and U21084 (N_21084,N_20737,N_20930);
and U21085 (N_21085,N_20975,N_20588);
nand U21086 (N_21086,N_20845,N_20812);
xnor U21087 (N_21087,N_20707,N_20825);
xor U21088 (N_21088,N_20938,N_20563);
xor U21089 (N_21089,N_20660,N_20819);
and U21090 (N_21090,N_20732,N_20761);
nor U21091 (N_21091,N_20861,N_20895);
nand U21092 (N_21092,N_20931,N_20534);
xnor U21093 (N_21093,N_20909,N_20686);
nand U21094 (N_21094,N_20763,N_20626);
xor U21095 (N_21095,N_20950,N_20525);
nor U21096 (N_21096,N_20669,N_20991);
nor U21097 (N_21097,N_20888,N_20547);
and U21098 (N_21098,N_20674,N_20639);
xor U21099 (N_21099,N_20567,N_20901);
xor U21100 (N_21100,N_20822,N_20752);
or U21101 (N_21101,N_20913,N_20720);
and U21102 (N_21102,N_20985,N_20769);
nand U21103 (N_21103,N_20551,N_20758);
nand U21104 (N_21104,N_20992,N_20747);
xor U21105 (N_21105,N_20768,N_20908);
nand U21106 (N_21106,N_20646,N_20856);
nor U21107 (N_21107,N_20741,N_20953);
nand U21108 (N_21108,N_20739,N_20678);
and U21109 (N_21109,N_20677,N_20993);
nor U21110 (N_21110,N_20835,N_20671);
nand U21111 (N_21111,N_20562,N_20692);
nand U21112 (N_21112,N_20661,N_20651);
xnor U21113 (N_21113,N_20941,N_20605);
nand U21114 (N_21114,N_20989,N_20983);
xor U21115 (N_21115,N_20650,N_20546);
or U21116 (N_21116,N_20750,N_20868);
or U21117 (N_21117,N_20548,N_20977);
and U21118 (N_21118,N_20716,N_20501);
nand U21119 (N_21119,N_20805,N_20833);
xnor U21120 (N_21120,N_20830,N_20795);
or U21121 (N_21121,N_20693,N_20814);
xor U21122 (N_21122,N_20754,N_20978);
xnor U21123 (N_21123,N_20766,N_20971);
nand U21124 (N_21124,N_20628,N_20645);
nand U21125 (N_21125,N_20615,N_20995);
and U21126 (N_21126,N_20884,N_20904);
and U21127 (N_21127,N_20536,N_20937);
and U21128 (N_21128,N_20710,N_20893);
nand U21129 (N_21129,N_20638,N_20583);
xnor U21130 (N_21130,N_20999,N_20559);
and U21131 (N_21131,N_20585,N_20625);
or U21132 (N_21132,N_20600,N_20963);
xor U21133 (N_21133,N_20789,N_20533);
xnor U21134 (N_21134,N_20962,N_20922);
or U21135 (N_21135,N_20877,N_20527);
and U21136 (N_21136,N_20824,N_20619);
nand U21137 (N_21137,N_20618,N_20951);
nor U21138 (N_21138,N_20586,N_20500);
or U21139 (N_21139,N_20666,N_20735);
and U21140 (N_21140,N_20774,N_20836);
or U21141 (N_21141,N_20779,N_20749);
or U21142 (N_21142,N_20579,N_20627);
and U21143 (N_21143,N_20906,N_20596);
nand U21144 (N_21144,N_20518,N_20759);
and U21145 (N_21145,N_20698,N_20972);
and U21146 (N_21146,N_20863,N_20591);
nand U21147 (N_21147,N_20513,N_20694);
and U21148 (N_21148,N_20755,N_20969);
xor U21149 (N_21149,N_20742,N_20935);
nand U21150 (N_21150,N_20714,N_20599);
nand U21151 (N_21151,N_20801,N_20890);
and U21152 (N_21152,N_20810,N_20738);
nor U21153 (N_21153,N_20701,N_20925);
and U21154 (N_21154,N_20662,N_20944);
xnor U21155 (N_21155,N_20859,N_20555);
or U21156 (N_21156,N_20920,N_20771);
or U21157 (N_21157,N_20602,N_20512);
or U21158 (N_21158,N_20675,N_20526);
xor U21159 (N_21159,N_20631,N_20862);
and U21160 (N_21160,N_20797,N_20569);
nand U21161 (N_21161,N_20690,N_20699);
xor U21162 (N_21162,N_20821,N_20839);
nand U21163 (N_21163,N_20873,N_20545);
and U21164 (N_21164,N_20886,N_20879);
or U21165 (N_21165,N_20872,N_20606);
xor U21166 (N_21166,N_20947,N_20624);
nand U21167 (N_21167,N_20926,N_20687);
xnor U21168 (N_21168,N_20620,N_20704);
and U21169 (N_21169,N_20593,N_20968);
and U21170 (N_21170,N_20948,N_20865);
nor U21171 (N_21171,N_20637,N_20657);
nor U21172 (N_21172,N_20842,N_20617);
or U21173 (N_21173,N_20673,N_20878);
and U21174 (N_21174,N_20816,N_20815);
nand U21175 (N_21175,N_20640,N_20967);
nor U21176 (N_21176,N_20936,N_20976);
and U21177 (N_21177,N_20516,N_20955);
and U21178 (N_21178,N_20725,N_20956);
xnor U21179 (N_21179,N_20918,N_20574);
nor U21180 (N_21180,N_20965,N_20994);
nor U21181 (N_21181,N_20541,N_20858);
or U21182 (N_21182,N_20731,N_20508);
or U21183 (N_21183,N_20964,N_20635);
nand U21184 (N_21184,N_20907,N_20898);
nor U21185 (N_21185,N_20849,N_20990);
xor U21186 (N_21186,N_20630,N_20988);
xor U21187 (N_21187,N_20787,N_20532);
nor U21188 (N_21188,N_20793,N_20734);
and U21189 (N_21189,N_20538,N_20655);
or U21190 (N_21190,N_20892,N_20773);
or U21191 (N_21191,N_20641,N_20765);
xor U21192 (N_21192,N_20572,N_20899);
or U21193 (N_21193,N_20643,N_20770);
and U21194 (N_21194,N_20753,N_20658);
nor U21195 (N_21195,N_20608,N_20633);
or U21196 (N_21196,N_20997,N_20785);
xnor U21197 (N_21197,N_20663,N_20912);
nor U21198 (N_21198,N_20905,N_20679);
nor U21199 (N_21199,N_20903,N_20803);
nand U21200 (N_21200,N_20592,N_20531);
xor U21201 (N_21201,N_20813,N_20757);
nor U21202 (N_21202,N_20982,N_20857);
or U21203 (N_21203,N_20623,N_20598);
nand U21204 (N_21204,N_20851,N_20715);
nor U21205 (N_21205,N_20871,N_20568);
or U21206 (N_21206,N_20644,N_20575);
and U21207 (N_21207,N_20683,N_20723);
nor U21208 (N_21208,N_20522,N_20916);
xor U21209 (N_21209,N_20506,N_20945);
xor U21210 (N_21210,N_20696,N_20607);
xor U21211 (N_21211,N_20622,N_20952);
nor U21212 (N_21212,N_20802,N_20838);
and U21213 (N_21213,N_20601,N_20846);
xnor U21214 (N_21214,N_20957,N_20509);
nand U21215 (N_21215,N_20697,N_20537);
nand U21216 (N_21216,N_20790,N_20784);
nor U21217 (N_21217,N_20746,N_20799);
nor U21218 (N_21218,N_20902,N_20743);
and U21219 (N_21219,N_20681,N_20781);
or U21220 (N_21220,N_20869,N_20542);
nand U21221 (N_21221,N_20664,N_20826);
xnor U21222 (N_21222,N_20946,N_20807);
nand U21223 (N_21223,N_20854,N_20589);
and U21224 (N_21224,N_20523,N_20711);
and U21225 (N_21225,N_20855,N_20841);
nor U21226 (N_21226,N_20709,N_20614);
or U21227 (N_21227,N_20864,N_20831);
or U21228 (N_21228,N_20665,N_20788);
xor U21229 (N_21229,N_20604,N_20979);
xor U21230 (N_21230,N_20566,N_20609);
xor U21231 (N_21231,N_20914,N_20621);
and U21232 (N_21232,N_20850,N_20736);
xor U21233 (N_21233,N_20728,N_20554);
or U21234 (N_21234,N_20894,N_20649);
nand U21235 (N_21235,N_20520,N_20595);
nand U21236 (N_21236,N_20760,N_20511);
nor U21237 (N_21237,N_20653,N_20874);
or U21238 (N_21238,N_20580,N_20852);
and U21239 (N_21239,N_20876,N_20632);
nand U21240 (N_21240,N_20883,N_20778);
and U21241 (N_21241,N_20804,N_20970);
nor U21242 (N_21242,N_20727,N_20837);
and U21243 (N_21243,N_20919,N_20721);
or U21244 (N_21244,N_20897,N_20705);
xnor U21245 (N_21245,N_20521,N_20808);
or U21246 (N_21246,N_20986,N_20828);
nor U21247 (N_21247,N_20656,N_20730);
and U21248 (N_21248,N_20712,N_20672);
and U21249 (N_21249,N_20507,N_20929);
nor U21250 (N_21250,N_20583,N_20615);
or U21251 (N_21251,N_20942,N_20817);
nor U21252 (N_21252,N_20890,N_20657);
nor U21253 (N_21253,N_20993,N_20894);
or U21254 (N_21254,N_20800,N_20911);
xor U21255 (N_21255,N_20991,N_20900);
nand U21256 (N_21256,N_20562,N_20508);
nand U21257 (N_21257,N_20898,N_20561);
nor U21258 (N_21258,N_20666,N_20751);
or U21259 (N_21259,N_20688,N_20626);
nand U21260 (N_21260,N_20539,N_20829);
nand U21261 (N_21261,N_20657,N_20844);
or U21262 (N_21262,N_20723,N_20524);
and U21263 (N_21263,N_20609,N_20832);
nor U21264 (N_21264,N_20830,N_20857);
nand U21265 (N_21265,N_20727,N_20783);
nor U21266 (N_21266,N_20620,N_20664);
or U21267 (N_21267,N_20958,N_20950);
or U21268 (N_21268,N_20758,N_20642);
nor U21269 (N_21269,N_20845,N_20991);
xor U21270 (N_21270,N_20733,N_20778);
nor U21271 (N_21271,N_20727,N_20771);
and U21272 (N_21272,N_20536,N_20587);
or U21273 (N_21273,N_20686,N_20768);
nand U21274 (N_21274,N_20897,N_20677);
and U21275 (N_21275,N_20951,N_20966);
nor U21276 (N_21276,N_20933,N_20899);
nor U21277 (N_21277,N_20815,N_20741);
xnor U21278 (N_21278,N_20978,N_20866);
nor U21279 (N_21279,N_20592,N_20664);
or U21280 (N_21280,N_20614,N_20559);
nor U21281 (N_21281,N_20656,N_20718);
nand U21282 (N_21282,N_20952,N_20977);
or U21283 (N_21283,N_20982,N_20540);
and U21284 (N_21284,N_20576,N_20530);
nand U21285 (N_21285,N_20974,N_20761);
or U21286 (N_21286,N_20523,N_20988);
nand U21287 (N_21287,N_20564,N_20519);
and U21288 (N_21288,N_20782,N_20976);
and U21289 (N_21289,N_20973,N_20992);
and U21290 (N_21290,N_20628,N_20966);
and U21291 (N_21291,N_20749,N_20665);
or U21292 (N_21292,N_20547,N_20520);
or U21293 (N_21293,N_20821,N_20604);
or U21294 (N_21294,N_20695,N_20823);
and U21295 (N_21295,N_20521,N_20740);
or U21296 (N_21296,N_20837,N_20907);
xnor U21297 (N_21297,N_20997,N_20706);
xnor U21298 (N_21298,N_20908,N_20625);
and U21299 (N_21299,N_20552,N_20904);
nor U21300 (N_21300,N_20604,N_20686);
or U21301 (N_21301,N_20501,N_20896);
nor U21302 (N_21302,N_20508,N_20846);
nor U21303 (N_21303,N_20538,N_20531);
and U21304 (N_21304,N_20838,N_20616);
and U21305 (N_21305,N_20984,N_20842);
nand U21306 (N_21306,N_20890,N_20924);
xor U21307 (N_21307,N_20531,N_20946);
and U21308 (N_21308,N_20930,N_20647);
and U21309 (N_21309,N_20740,N_20866);
nor U21310 (N_21310,N_20627,N_20860);
xor U21311 (N_21311,N_20819,N_20767);
or U21312 (N_21312,N_20522,N_20672);
or U21313 (N_21313,N_20958,N_20544);
or U21314 (N_21314,N_20912,N_20805);
nor U21315 (N_21315,N_20545,N_20711);
nand U21316 (N_21316,N_20750,N_20595);
nand U21317 (N_21317,N_20751,N_20848);
and U21318 (N_21318,N_20536,N_20893);
nor U21319 (N_21319,N_20676,N_20884);
or U21320 (N_21320,N_20612,N_20989);
and U21321 (N_21321,N_20798,N_20711);
nor U21322 (N_21322,N_20530,N_20712);
xor U21323 (N_21323,N_20904,N_20776);
nor U21324 (N_21324,N_20716,N_20900);
or U21325 (N_21325,N_20681,N_20669);
nor U21326 (N_21326,N_20814,N_20765);
nor U21327 (N_21327,N_20800,N_20536);
nor U21328 (N_21328,N_20534,N_20643);
or U21329 (N_21329,N_20871,N_20954);
nor U21330 (N_21330,N_20717,N_20769);
nand U21331 (N_21331,N_20841,N_20885);
nand U21332 (N_21332,N_20700,N_20944);
and U21333 (N_21333,N_20645,N_20782);
xor U21334 (N_21334,N_20966,N_20871);
xor U21335 (N_21335,N_20591,N_20664);
nor U21336 (N_21336,N_20830,N_20704);
or U21337 (N_21337,N_20520,N_20728);
nor U21338 (N_21338,N_20748,N_20659);
nand U21339 (N_21339,N_20541,N_20705);
or U21340 (N_21340,N_20711,N_20563);
nor U21341 (N_21341,N_20565,N_20708);
and U21342 (N_21342,N_20635,N_20936);
nand U21343 (N_21343,N_20815,N_20631);
or U21344 (N_21344,N_20739,N_20687);
and U21345 (N_21345,N_20867,N_20645);
xor U21346 (N_21346,N_20924,N_20888);
and U21347 (N_21347,N_20870,N_20811);
nand U21348 (N_21348,N_20672,N_20597);
or U21349 (N_21349,N_20763,N_20771);
or U21350 (N_21350,N_20748,N_20788);
or U21351 (N_21351,N_20860,N_20924);
and U21352 (N_21352,N_20657,N_20629);
nor U21353 (N_21353,N_20664,N_20989);
and U21354 (N_21354,N_20726,N_20614);
nand U21355 (N_21355,N_20526,N_20558);
xnor U21356 (N_21356,N_20547,N_20903);
xor U21357 (N_21357,N_20754,N_20980);
or U21358 (N_21358,N_20896,N_20770);
nand U21359 (N_21359,N_20911,N_20914);
or U21360 (N_21360,N_20929,N_20990);
nand U21361 (N_21361,N_20615,N_20682);
nor U21362 (N_21362,N_20756,N_20927);
xor U21363 (N_21363,N_20994,N_20648);
nor U21364 (N_21364,N_20530,N_20628);
or U21365 (N_21365,N_20974,N_20810);
and U21366 (N_21366,N_20742,N_20535);
nor U21367 (N_21367,N_20622,N_20919);
xor U21368 (N_21368,N_20807,N_20673);
and U21369 (N_21369,N_20822,N_20885);
nor U21370 (N_21370,N_20500,N_20561);
nand U21371 (N_21371,N_20594,N_20788);
nor U21372 (N_21372,N_20707,N_20963);
nor U21373 (N_21373,N_20505,N_20937);
or U21374 (N_21374,N_20615,N_20525);
and U21375 (N_21375,N_20949,N_20938);
or U21376 (N_21376,N_20965,N_20525);
xor U21377 (N_21377,N_20701,N_20883);
and U21378 (N_21378,N_20942,N_20635);
xnor U21379 (N_21379,N_20675,N_20656);
and U21380 (N_21380,N_20617,N_20603);
xor U21381 (N_21381,N_20819,N_20624);
xor U21382 (N_21382,N_20847,N_20968);
xnor U21383 (N_21383,N_20646,N_20515);
nand U21384 (N_21384,N_20639,N_20768);
and U21385 (N_21385,N_20752,N_20919);
xnor U21386 (N_21386,N_20638,N_20991);
nand U21387 (N_21387,N_20802,N_20886);
and U21388 (N_21388,N_20855,N_20837);
nand U21389 (N_21389,N_20923,N_20701);
and U21390 (N_21390,N_20772,N_20868);
and U21391 (N_21391,N_20966,N_20552);
and U21392 (N_21392,N_20773,N_20950);
nor U21393 (N_21393,N_20641,N_20595);
and U21394 (N_21394,N_20565,N_20567);
nand U21395 (N_21395,N_20672,N_20778);
xnor U21396 (N_21396,N_20758,N_20797);
nand U21397 (N_21397,N_20670,N_20712);
and U21398 (N_21398,N_20617,N_20580);
and U21399 (N_21399,N_20969,N_20771);
and U21400 (N_21400,N_20831,N_20777);
and U21401 (N_21401,N_20618,N_20957);
or U21402 (N_21402,N_20804,N_20952);
nand U21403 (N_21403,N_20659,N_20605);
nand U21404 (N_21404,N_20695,N_20888);
nor U21405 (N_21405,N_20796,N_20743);
nor U21406 (N_21406,N_20667,N_20790);
xor U21407 (N_21407,N_20732,N_20651);
and U21408 (N_21408,N_20596,N_20905);
or U21409 (N_21409,N_20820,N_20947);
or U21410 (N_21410,N_20970,N_20555);
and U21411 (N_21411,N_20515,N_20858);
and U21412 (N_21412,N_20562,N_20718);
and U21413 (N_21413,N_20730,N_20625);
and U21414 (N_21414,N_20611,N_20636);
nor U21415 (N_21415,N_20854,N_20920);
nor U21416 (N_21416,N_20864,N_20896);
nor U21417 (N_21417,N_20686,N_20644);
and U21418 (N_21418,N_20617,N_20777);
and U21419 (N_21419,N_20910,N_20682);
and U21420 (N_21420,N_20510,N_20702);
or U21421 (N_21421,N_20592,N_20860);
xnor U21422 (N_21422,N_20555,N_20763);
nand U21423 (N_21423,N_20744,N_20502);
xnor U21424 (N_21424,N_20567,N_20643);
or U21425 (N_21425,N_20978,N_20727);
nor U21426 (N_21426,N_20967,N_20995);
and U21427 (N_21427,N_20843,N_20813);
and U21428 (N_21428,N_20789,N_20664);
and U21429 (N_21429,N_20903,N_20644);
or U21430 (N_21430,N_20585,N_20736);
nor U21431 (N_21431,N_20912,N_20851);
nand U21432 (N_21432,N_20935,N_20606);
nor U21433 (N_21433,N_20597,N_20828);
xnor U21434 (N_21434,N_20983,N_20778);
or U21435 (N_21435,N_20648,N_20891);
or U21436 (N_21436,N_20506,N_20835);
or U21437 (N_21437,N_20702,N_20663);
xor U21438 (N_21438,N_20546,N_20694);
nor U21439 (N_21439,N_20623,N_20574);
and U21440 (N_21440,N_20525,N_20686);
xnor U21441 (N_21441,N_20655,N_20571);
nand U21442 (N_21442,N_20886,N_20953);
xor U21443 (N_21443,N_20943,N_20954);
xor U21444 (N_21444,N_20568,N_20962);
nor U21445 (N_21445,N_20526,N_20630);
and U21446 (N_21446,N_20640,N_20662);
and U21447 (N_21447,N_20939,N_20754);
xor U21448 (N_21448,N_20762,N_20723);
nor U21449 (N_21449,N_20554,N_20656);
and U21450 (N_21450,N_20581,N_20572);
or U21451 (N_21451,N_20735,N_20589);
and U21452 (N_21452,N_20515,N_20992);
xnor U21453 (N_21453,N_20747,N_20776);
nand U21454 (N_21454,N_20920,N_20847);
xor U21455 (N_21455,N_20623,N_20800);
nor U21456 (N_21456,N_20928,N_20587);
and U21457 (N_21457,N_20942,N_20570);
nor U21458 (N_21458,N_20555,N_20994);
nor U21459 (N_21459,N_20956,N_20586);
xnor U21460 (N_21460,N_20626,N_20610);
xnor U21461 (N_21461,N_20826,N_20790);
nand U21462 (N_21462,N_20791,N_20579);
nor U21463 (N_21463,N_20702,N_20530);
nand U21464 (N_21464,N_20522,N_20561);
or U21465 (N_21465,N_20608,N_20738);
nor U21466 (N_21466,N_20675,N_20613);
nand U21467 (N_21467,N_20660,N_20636);
or U21468 (N_21468,N_20731,N_20714);
nor U21469 (N_21469,N_20961,N_20818);
nor U21470 (N_21470,N_20960,N_20952);
nand U21471 (N_21471,N_20872,N_20724);
nand U21472 (N_21472,N_20507,N_20828);
xnor U21473 (N_21473,N_20996,N_20873);
nand U21474 (N_21474,N_20893,N_20897);
and U21475 (N_21475,N_20772,N_20637);
xor U21476 (N_21476,N_20919,N_20688);
nor U21477 (N_21477,N_20502,N_20625);
or U21478 (N_21478,N_20637,N_20977);
nand U21479 (N_21479,N_20779,N_20505);
nor U21480 (N_21480,N_20621,N_20733);
and U21481 (N_21481,N_20556,N_20636);
or U21482 (N_21482,N_20623,N_20839);
nand U21483 (N_21483,N_20890,N_20848);
or U21484 (N_21484,N_20837,N_20591);
and U21485 (N_21485,N_20501,N_20986);
nand U21486 (N_21486,N_20623,N_20856);
and U21487 (N_21487,N_20566,N_20552);
or U21488 (N_21488,N_20952,N_20519);
xnor U21489 (N_21489,N_20560,N_20916);
and U21490 (N_21490,N_20702,N_20658);
and U21491 (N_21491,N_20751,N_20877);
xor U21492 (N_21492,N_20753,N_20725);
xor U21493 (N_21493,N_20884,N_20885);
or U21494 (N_21494,N_20735,N_20900);
nand U21495 (N_21495,N_20997,N_20592);
and U21496 (N_21496,N_20809,N_20882);
and U21497 (N_21497,N_20732,N_20542);
or U21498 (N_21498,N_20641,N_20913);
nand U21499 (N_21499,N_20840,N_20760);
xor U21500 (N_21500,N_21193,N_21369);
or U21501 (N_21501,N_21482,N_21064);
xnor U21502 (N_21502,N_21428,N_21246);
and U21503 (N_21503,N_21441,N_21200);
or U21504 (N_21504,N_21387,N_21418);
and U21505 (N_21505,N_21271,N_21244);
nor U21506 (N_21506,N_21232,N_21431);
nor U21507 (N_21507,N_21166,N_21410);
or U21508 (N_21508,N_21459,N_21274);
xor U21509 (N_21509,N_21411,N_21006);
xnor U21510 (N_21510,N_21372,N_21336);
xnor U21511 (N_21511,N_21165,N_21107);
and U21512 (N_21512,N_21305,N_21043);
and U21513 (N_21513,N_21367,N_21124);
or U21514 (N_21514,N_21360,N_21098);
or U21515 (N_21515,N_21404,N_21498);
and U21516 (N_21516,N_21474,N_21283);
nand U21517 (N_21517,N_21121,N_21061);
xor U21518 (N_21518,N_21446,N_21344);
or U21519 (N_21519,N_21077,N_21249);
or U21520 (N_21520,N_21310,N_21088);
xnor U21521 (N_21521,N_21148,N_21079);
or U21522 (N_21522,N_21081,N_21172);
nor U21523 (N_21523,N_21253,N_21044);
and U21524 (N_21524,N_21201,N_21300);
nand U21525 (N_21525,N_21227,N_21101);
and U21526 (N_21526,N_21256,N_21025);
nand U21527 (N_21527,N_21097,N_21291);
and U21528 (N_21528,N_21213,N_21119);
or U21529 (N_21529,N_21037,N_21421);
and U21530 (N_21530,N_21219,N_21013);
or U21531 (N_21531,N_21465,N_21447);
or U21532 (N_21532,N_21481,N_21018);
or U21533 (N_21533,N_21318,N_21074);
nor U21534 (N_21534,N_21399,N_21270);
or U21535 (N_21535,N_21178,N_21438);
and U21536 (N_21536,N_21021,N_21080);
nand U21537 (N_21537,N_21276,N_21339);
or U21538 (N_21538,N_21192,N_21290);
or U21539 (N_21539,N_21440,N_21126);
nor U21540 (N_21540,N_21089,N_21324);
or U21541 (N_21541,N_21164,N_21345);
nand U21542 (N_21542,N_21480,N_21221);
and U21543 (N_21543,N_21112,N_21231);
nor U21544 (N_21544,N_21083,N_21194);
xnor U21545 (N_21545,N_21365,N_21398);
or U21546 (N_21546,N_21199,N_21279);
nand U21547 (N_21547,N_21351,N_21479);
and U21548 (N_21548,N_21304,N_21241);
or U21549 (N_21549,N_21058,N_21214);
nor U21550 (N_21550,N_21278,N_21461);
xnor U21551 (N_21551,N_21175,N_21051);
nor U21552 (N_21552,N_21314,N_21316);
and U21553 (N_21553,N_21469,N_21054);
or U21554 (N_21554,N_21180,N_21347);
xnor U21555 (N_21555,N_21208,N_21104);
or U21556 (N_21556,N_21093,N_21209);
nand U21557 (N_21557,N_21229,N_21266);
xnor U21558 (N_21558,N_21460,N_21202);
or U21559 (N_21559,N_21417,N_21471);
xor U21560 (N_21560,N_21235,N_21243);
nand U21561 (N_21561,N_21153,N_21149);
or U21562 (N_21562,N_21182,N_21176);
and U21563 (N_21563,N_21495,N_21204);
nand U21564 (N_21564,N_21497,N_21046);
nand U21565 (N_21565,N_21008,N_21250);
or U21566 (N_21566,N_21301,N_21419);
nor U21567 (N_21567,N_21400,N_21135);
xnor U21568 (N_21568,N_21273,N_21415);
nor U21569 (N_21569,N_21371,N_21009);
xor U21570 (N_21570,N_21167,N_21335);
nor U21571 (N_21571,N_21319,N_21434);
or U21572 (N_21572,N_21147,N_21174);
nor U21573 (N_21573,N_21412,N_21113);
nand U21574 (N_21574,N_21352,N_21285);
nand U21575 (N_21575,N_21189,N_21233);
nand U21576 (N_21576,N_21389,N_21303);
and U21577 (N_21577,N_21409,N_21102);
nand U21578 (N_21578,N_21420,N_21312);
nor U21579 (N_21579,N_21267,N_21143);
nor U21580 (N_21580,N_21252,N_21185);
or U21581 (N_21581,N_21217,N_21125);
xor U21582 (N_21582,N_21466,N_21364);
nor U21583 (N_21583,N_21075,N_21368);
and U21584 (N_21584,N_21152,N_21132);
nor U21585 (N_21585,N_21222,N_21131);
and U21586 (N_21586,N_21425,N_21163);
xor U21587 (N_21587,N_21133,N_21378);
nor U21588 (N_21588,N_21401,N_21067);
and U21589 (N_21589,N_21216,N_21491);
and U21590 (N_21590,N_21255,N_21001);
or U21591 (N_21591,N_21297,N_21071);
nor U21592 (N_21592,N_21159,N_21040);
nand U21593 (N_21593,N_21122,N_21085);
or U21594 (N_21594,N_21464,N_21045);
xor U21595 (N_21595,N_21026,N_21141);
or U21596 (N_21596,N_21109,N_21263);
xor U21597 (N_21597,N_21057,N_21358);
and U21598 (N_21598,N_21269,N_21332);
or U21599 (N_21599,N_21490,N_21186);
nand U21600 (N_21600,N_21309,N_21184);
or U21601 (N_21601,N_21333,N_21343);
nor U21602 (N_21602,N_21385,N_21203);
and U21603 (N_21603,N_21116,N_21029);
nand U21604 (N_21604,N_21313,N_21003);
nand U21605 (N_21605,N_21477,N_21388);
or U21606 (N_21606,N_21099,N_21151);
xor U21607 (N_21607,N_21111,N_21160);
nor U21608 (N_21608,N_21416,N_21448);
nand U21609 (N_21609,N_21090,N_21258);
or U21610 (N_21610,N_21036,N_21238);
or U21611 (N_21611,N_21407,N_21329);
xor U21612 (N_21612,N_21082,N_21120);
xnor U21613 (N_21613,N_21393,N_21257);
or U21614 (N_21614,N_21261,N_21210);
nor U21615 (N_21615,N_21170,N_21042);
nor U21616 (N_21616,N_21472,N_21445);
and U21617 (N_21617,N_21287,N_21264);
xor U21618 (N_21618,N_21158,N_21414);
nand U21619 (N_21619,N_21228,N_21442);
nor U21620 (N_21620,N_21038,N_21259);
xnor U21621 (N_21621,N_21103,N_21195);
and U21622 (N_21622,N_21405,N_21296);
and U21623 (N_21623,N_21475,N_21374);
nor U21624 (N_21624,N_21327,N_21390);
nand U21625 (N_21625,N_21179,N_21130);
or U21626 (N_21626,N_21322,N_21295);
xnor U21627 (N_21627,N_21069,N_21062);
xnor U21628 (N_21628,N_21260,N_21034);
and U21629 (N_21629,N_21177,N_21338);
xnor U21630 (N_21630,N_21114,N_21489);
nor U21631 (N_21631,N_21355,N_21108);
or U21632 (N_21632,N_21155,N_21383);
or U21633 (N_21633,N_21022,N_21137);
and U21634 (N_21634,N_21357,N_21380);
or U21635 (N_21635,N_21427,N_21325);
nand U21636 (N_21636,N_21342,N_21242);
nand U21637 (N_21637,N_21262,N_21236);
nor U21638 (N_21638,N_21348,N_21424);
and U21639 (N_21639,N_21039,N_21053);
nand U21640 (N_21640,N_21012,N_21019);
xnor U21641 (N_21641,N_21394,N_21451);
xnor U21642 (N_21642,N_21437,N_21072);
xor U21643 (N_21643,N_21092,N_21328);
nand U21644 (N_21644,N_21488,N_21140);
or U21645 (N_21645,N_21454,N_21105);
or U21646 (N_21646,N_21220,N_21494);
and U21647 (N_21647,N_21485,N_21286);
and U21648 (N_21648,N_21065,N_21031);
or U21649 (N_21649,N_21207,N_21307);
xnor U21650 (N_21650,N_21323,N_21033);
or U21651 (N_21651,N_21188,N_21017);
or U21652 (N_21652,N_21002,N_21063);
nand U21653 (N_21653,N_21359,N_21168);
or U21654 (N_21654,N_21123,N_21430);
xnor U21655 (N_21655,N_21396,N_21076);
xor U21656 (N_21656,N_21373,N_21483);
and U21657 (N_21657,N_21408,N_21473);
or U21658 (N_21658,N_21066,N_21321);
and U21659 (N_21659,N_21384,N_21115);
or U21660 (N_21660,N_21056,N_21138);
or U21661 (N_21661,N_21049,N_21086);
nand U21662 (N_21662,N_21280,N_21306);
nor U21663 (N_21663,N_21190,N_21311);
xnor U21664 (N_21664,N_21499,N_21302);
xnor U21665 (N_21665,N_21350,N_21361);
nor U21666 (N_21666,N_21239,N_21059);
nand U21667 (N_21667,N_21395,N_21432);
or U21668 (N_21668,N_21308,N_21289);
nor U21669 (N_21669,N_21268,N_21376);
nand U21670 (N_21670,N_21128,N_21183);
nor U21671 (N_21671,N_21020,N_21218);
nand U21672 (N_21672,N_21173,N_21106);
xor U21673 (N_21673,N_21024,N_21462);
and U21674 (N_21674,N_21030,N_21340);
or U21675 (N_21675,N_21320,N_21456);
and U21676 (N_21676,N_21248,N_21382);
nand U21677 (N_21677,N_21237,N_21055);
and U21678 (N_21678,N_21377,N_21047);
nand U21679 (N_21679,N_21455,N_21370);
or U21680 (N_21680,N_21452,N_21337);
and U21681 (N_21681,N_21288,N_21134);
and U21682 (N_21682,N_21487,N_21486);
nor U21683 (N_21683,N_21027,N_21315);
nor U21684 (N_21684,N_21225,N_21215);
nor U21685 (N_21685,N_21245,N_21096);
or U21686 (N_21686,N_21095,N_21145);
nand U21687 (N_21687,N_21197,N_21161);
nor U21688 (N_21688,N_21035,N_21413);
nor U21689 (N_21689,N_21292,N_21354);
nand U21690 (N_21690,N_21453,N_21362);
or U21691 (N_21691,N_21277,N_21230);
or U21692 (N_21692,N_21349,N_21060);
or U21693 (N_21693,N_21010,N_21251);
xor U21694 (N_21694,N_21272,N_21493);
nand U21695 (N_21695,N_21478,N_21187);
xor U21696 (N_21696,N_21224,N_21041);
nand U21697 (N_21697,N_21299,N_21144);
nand U21698 (N_21698,N_21100,N_21223);
and U21699 (N_21699,N_21444,N_21356);
nor U21700 (N_21700,N_21023,N_21363);
or U21701 (N_21701,N_21381,N_21391);
or U21702 (N_21702,N_21423,N_21139);
nand U21703 (N_21703,N_21330,N_21275);
nand U21704 (N_21704,N_21136,N_21375);
or U21705 (N_21705,N_21129,N_21331);
nand U21706 (N_21706,N_21169,N_21484);
nand U21707 (N_21707,N_21171,N_21265);
xnor U21708 (N_21708,N_21293,N_21386);
nand U21709 (N_21709,N_21403,N_21181);
nor U21710 (N_21710,N_21467,N_21005);
or U21711 (N_21711,N_21298,N_21439);
xor U21712 (N_21712,N_21247,N_21028);
or U21713 (N_21713,N_21191,N_21048);
or U21714 (N_21714,N_21435,N_21118);
nor U21715 (N_21715,N_21450,N_21294);
or U21716 (N_21716,N_21234,N_21470);
nor U21717 (N_21717,N_21196,N_21226);
and U21718 (N_21718,N_21087,N_21254);
nand U21719 (N_21719,N_21392,N_21433);
and U21720 (N_21720,N_21281,N_21284);
nand U21721 (N_21721,N_21476,N_21422);
nor U21722 (N_21722,N_21084,N_21206);
and U21723 (N_21723,N_21334,N_21492);
xnor U21724 (N_21724,N_21016,N_21240);
nand U21725 (N_21725,N_21007,N_21015);
or U21726 (N_21726,N_21463,N_21496);
xnor U21727 (N_21727,N_21156,N_21142);
or U21728 (N_21728,N_21117,N_21426);
nand U21729 (N_21729,N_21154,N_21406);
nand U21730 (N_21730,N_21379,N_21458);
and U21731 (N_21731,N_21162,N_21032);
nand U21732 (N_21732,N_21317,N_21150);
nand U21733 (N_21733,N_21198,N_21004);
and U21734 (N_21734,N_21070,N_21436);
or U21735 (N_21735,N_21211,N_21011);
or U21736 (N_21736,N_21212,N_21353);
or U21737 (N_21737,N_21341,N_21468);
xor U21738 (N_21738,N_21366,N_21157);
xnor U21739 (N_21739,N_21346,N_21073);
nor U21740 (N_21740,N_21127,N_21052);
xor U21741 (N_21741,N_21146,N_21110);
nor U21742 (N_21742,N_21429,N_21091);
or U21743 (N_21743,N_21457,N_21449);
nor U21744 (N_21744,N_21326,N_21014);
or U21745 (N_21745,N_21205,N_21050);
and U21746 (N_21746,N_21402,N_21068);
or U21747 (N_21747,N_21397,N_21094);
and U21748 (N_21748,N_21000,N_21282);
nand U21749 (N_21749,N_21443,N_21078);
xnor U21750 (N_21750,N_21267,N_21258);
nand U21751 (N_21751,N_21419,N_21410);
nor U21752 (N_21752,N_21118,N_21483);
or U21753 (N_21753,N_21216,N_21104);
or U21754 (N_21754,N_21237,N_21053);
and U21755 (N_21755,N_21020,N_21101);
nand U21756 (N_21756,N_21312,N_21267);
or U21757 (N_21757,N_21046,N_21217);
or U21758 (N_21758,N_21117,N_21458);
and U21759 (N_21759,N_21204,N_21000);
nor U21760 (N_21760,N_21109,N_21375);
nand U21761 (N_21761,N_21414,N_21167);
nor U21762 (N_21762,N_21073,N_21471);
nor U21763 (N_21763,N_21389,N_21447);
or U21764 (N_21764,N_21152,N_21016);
or U21765 (N_21765,N_21223,N_21278);
nor U21766 (N_21766,N_21398,N_21011);
or U21767 (N_21767,N_21107,N_21172);
nand U21768 (N_21768,N_21396,N_21186);
nand U21769 (N_21769,N_21433,N_21355);
xor U21770 (N_21770,N_21091,N_21299);
and U21771 (N_21771,N_21037,N_21134);
nand U21772 (N_21772,N_21064,N_21104);
nand U21773 (N_21773,N_21453,N_21103);
and U21774 (N_21774,N_21118,N_21253);
or U21775 (N_21775,N_21442,N_21164);
xor U21776 (N_21776,N_21396,N_21333);
or U21777 (N_21777,N_21094,N_21475);
and U21778 (N_21778,N_21248,N_21106);
xor U21779 (N_21779,N_21045,N_21447);
nand U21780 (N_21780,N_21169,N_21476);
nand U21781 (N_21781,N_21305,N_21194);
xnor U21782 (N_21782,N_21195,N_21006);
and U21783 (N_21783,N_21276,N_21423);
nor U21784 (N_21784,N_21287,N_21459);
and U21785 (N_21785,N_21212,N_21333);
or U21786 (N_21786,N_21376,N_21142);
or U21787 (N_21787,N_21489,N_21192);
nand U21788 (N_21788,N_21215,N_21344);
or U21789 (N_21789,N_21476,N_21036);
nand U21790 (N_21790,N_21094,N_21324);
xor U21791 (N_21791,N_21376,N_21176);
nor U21792 (N_21792,N_21055,N_21028);
nand U21793 (N_21793,N_21371,N_21220);
nand U21794 (N_21794,N_21396,N_21249);
and U21795 (N_21795,N_21496,N_21423);
nand U21796 (N_21796,N_21047,N_21231);
and U21797 (N_21797,N_21474,N_21319);
xnor U21798 (N_21798,N_21499,N_21355);
nor U21799 (N_21799,N_21153,N_21283);
and U21800 (N_21800,N_21401,N_21374);
and U21801 (N_21801,N_21055,N_21454);
nor U21802 (N_21802,N_21220,N_21242);
and U21803 (N_21803,N_21220,N_21235);
nor U21804 (N_21804,N_21278,N_21346);
xor U21805 (N_21805,N_21117,N_21457);
nand U21806 (N_21806,N_21347,N_21161);
and U21807 (N_21807,N_21062,N_21306);
or U21808 (N_21808,N_21256,N_21334);
and U21809 (N_21809,N_21294,N_21311);
or U21810 (N_21810,N_21169,N_21238);
nor U21811 (N_21811,N_21354,N_21272);
or U21812 (N_21812,N_21345,N_21209);
and U21813 (N_21813,N_21219,N_21289);
nor U21814 (N_21814,N_21010,N_21482);
nand U21815 (N_21815,N_21328,N_21172);
and U21816 (N_21816,N_21038,N_21125);
or U21817 (N_21817,N_21443,N_21495);
xor U21818 (N_21818,N_21329,N_21008);
nor U21819 (N_21819,N_21468,N_21101);
and U21820 (N_21820,N_21091,N_21011);
xnor U21821 (N_21821,N_21229,N_21013);
xor U21822 (N_21822,N_21255,N_21288);
or U21823 (N_21823,N_21444,N_21167);
xor U21824 (N_21824,N_21298,N_21357);
or U21825 (N_21825,N_21073,N_21495);
and U21826 (N_21826,N_21330,N_21268);
nand U21827 (N_21827,N_21151,N_21196);
xnor U21828 (N_21828,N_21188,N_21176);
nand U21829 (N_21829,N_21100,N_21374);
or U21830 (N_21830,N_21032,N_21474);
nor U21831 (N_21831,N_21428,N_21066);
and U21832 (N_21832,N_21495,N_21141);
and U21833 (N_21833,N_21252,N_21389);
xnor U21834 (N_21834,N_21135,N_21495);
and U21835 (N_21835,N_21332,N_21461);
or U21836 (N_21836,N_21336,N_21468);
xnor U21837 (N_21837,N_21399,N_21219);
or U21838 (N_21838,N_21264,N_21084);
xor U21839 (N_21839,N_21363,N_21020);
nor U21840 (N_21840,N_21314,N_21094);
and U21841 (N_21841,N_21476,N_21410);
xnor U21842 (N_21842,N_21031,N_21378);
or U21843 (N_21843,N_21291,N_21438);
or U21844 (N_21844,N_21346,N_21340);
nor U21845 (N_21845,N_21443,N_21478);
and U21846 (N_21846,N_21371,N_21016);
nand U21847 (N_21847,N_21442,N_21317);
nand U21848 (N_21848,N_21182,N_21031);
xor U21849 (N_21849,N_21216,N_21463);
or U21850 (N_21850,N_21090,N_21335);
and U21851 (N_21851,N_21410,N_21423);
xor U21852 (N_21852,N_21176,N_21331);
nand U21853 (N_21853,N_21394,N_21224);
nor U21854 (N_21854,N_21382,N_21433);
nand U21855 (N_21855,N_21194,N_21036);
and U21856 (N_21856,N_21424,N_21263);
or U21857 (N_21857,N_21471,N_21124);
xnor U21858 (N_21858,N_21495,N_21416);
xnor U21859 (N_21859,N_21365,N_21143);
or U21860 (N_21860,N_21470,N_21162);
or U21861 (N_21861,N_21094,N_21494);
and U21862 (N_21862,N_21173,N_21466);
nand U21863 (N_21863,N_21264,N_21459);
nand U21864 (N_21864,N_21148,N_21258);
xnor U21865 (N_21865,N_21235,N_21314);
xor U21866 (N_21866,N_21175,N_21371);
nor U21867 (N_21867,N_21493,N_21228);
and U21868 (N_21868,N_21029,N_21300);
nor U21869 (N_21869,N_21172,N_21269);
xor U21870 (N_21870,N_21451,N_21121);
and U21871 (N_21871,N_21438,N_21135);
or U21872 (N_21872,N_21256,N_21410);
xor U21873 (N_21873,N_21047,N_21064);
or U21874 (N_21874,N_21383,N_21180);
and U21875 (N_21875,N_21255,N_21400);
xnor U21876 (N_21876,N_21358,N_21144);
and U21877 (N_21877,N_21154,N_21116);
nand U21878 (N_21878,N_21274,N_21152);
nor U21879 (N_21879,N_21387,N_21198);
xor U21880 (N_21880,N_21312,N_21355);
nand U21881 (N_21881,N_21228,N_21073);
nand U21882 (N_21882,N_21112,N_21046);
nor U21883 (N_21883,N_21313,N_21449);
or U21884 (N_21884,N_21011,N_21323);
xnor U21885 (N_21885,N_21133,N_21325);
and U21886 (N_21886,N_21194,N_21210);
and U21887 (N_21887,N_21210,N_21158);
nand U21888 (N_21888,N_21384,N_21257);
or U21889 (N_21889,N_21260,N_21332);
xnor U21890 (N_21890,N_21425,N_21330);
xor U21891 (N_21891,N_21129,N_21157);
and U21892 (N_21892,N_21335,N_21422);
or U21893 (N_21893,N_21396,N_21175);
and U21894 (N_21894,N_21437,N_21156);
xor U21895 (N_21895,N_21208,N_21195);
xnor U21896 (N_21896,N_21355,N_21223);
xor U21897 (N_21897,N_21308,N_21463);
xnor U21898 (N_21898,N_21247,N_21211);
nor U21899 (N_21899,N_21232,N_21100);
nand U21900 (N_21900,N_21439,N_21106);
xnor U21901 (N_21901,N_21134,N_21435);
nor U21902 (N_21902,N_21156,N_21411);
and U21903 (N_21903,N_21117,N_21464);
or U21904 (N_21904,N_21473,N_21293);
nand U21905 (N_21905,N_21140,N_21025);
nand U21906 (N_21906,N_21268,N_21185);
nor U21907 (N_21907,N_21324,N_21485);
and U21908 (N_21908,N_21097,N_21410);
nor U21909 (N_21909,N_21402,N_21431);
or U21910 (N_21910,N_21149,N_21269);
and U21911 (N_21911,N_21136,N_21290);
nor U21912 (N_21912,N_21459,N_21135);
or U21913 (N_21913,N_21189,N_21125);
nor U21914 (N_21914,N_21217,N_21110);
or U21915 (N_21915,N_21056,N_21195);
and U21916 (N_21916,N_21212,N_21032);
and U21917 (N_21917,N_21218,N_21066);
nand U21918 (N_21918,N_21198,N_21161);
nand U21919 (N_21919,N_21234,N_21182);
xor U21920 (N_21920,N_21202,N_21062);
or U21921 (N_21921,N_21014,N_21478);
and U21922 (N_21922,N_21497,N_21296);
nand U21923 (N_21923,N_21156,N_21388);
xnor U21924 (N_21924,N_21163,N_21033);
or U21925 (N_21925,N_21273,N_21143);
nand U21926 (N_21926,N_21042,N_21244);
xor U21927 (N_21927,N_21285,N_21181);
and U21928 (N_21928,N_21311,N_21411);
and U21929 (N_21929,N_21497,N_21368);
and U21930 (N_21930,N_21012,N_21161);
nand U21931 (N_21931,N_21406,N_21282);
or U21932 (N_21932,N_21432,N_21115);
and U21933 (N_21933,N_21381,N_21093);
nand U21934 (N_21934,N_21086,N_21343);
and U21935 (N_21935,N_21111,N_21356);
nand U21936 (N_21936,N_21104,N_21085);
xor U21937 (N_21937,N_21367,N_21279);
xor U21938 (N_21938,N_21345,N_21347);
xor U21939 (N_21939,N_21004,N_21421);
nand U21940 (N_21940,N_21013,N_21155);
nand U21941 (N_21941,N_21401,N_21052);
nand U21942 (N_21942,N_21397,N_21479);
or U21943 (N_21943,N_21356,N_21218);
and U21944 (N_21944,N_21465,N_21033);
xnor U21945 (N_21945,N_21052,N_21496);
nor U21946 (N_21946,N_21458,N_21098);
or U21947 (N_21947,N_21383,N_21367);
and U21948 (N_21948,N_21496,N_21007);
and U21949 (N_21949,N_21418,N_21261);
xnor U21950 (N_21950,N_21228,N_21431);
nand U21951 (N_21951,N_21247,N_21185);
xor U21952 (N_21952,N_21275,N_21220);
or U21953 (N_21953,N_21283,N_21400);
and U21954 (N_21954,N_21411,N_21396);
or U21955 (N_21955,N_21499,N_21427);
and U21956 (N_21956,N_21132,N_21202);
xnor U21957 (N_21957,N_21375,N_21288);
and U21958 (N_21958,N_21458,N_21229);
and U21959 (N_21959,N_21402,N_21123);
xnor U21960 (N_21960,N_21378,N_21059);
or U21961 (N_21961,N_21193,N_21474);
or U21962 (N_21962,N_21372,N_21448);
and U21963 (N_21963,N_21094,N_21139);
nand U21964 (N_21964,N_21188,N_21077);
or U21965 (N_21965,N_21131,N_21087);
nand U21966 (N_21966,N_21272,N_21494);
xor U21967 (N_21967,N_21211,N_21009);
or U21968 (N_21968,N_21427,N_21068);
and U21969 (N_21969,N_21097,N_21276);
nand U21970 (N_21970,N_21073,N_21132);
or U21971 (N_21971,N_21038,N_21417);
nand U21972 (N_21972,N_21260,N_21061);
nand U21973 (N_21973,N_21304,N_21412);
nor U21974 (N_21974,N_21139,N_21436);
and U21975 (N_21975,N_21244,N_21297);
nand U21976 (N_21976,N_21406,N_21091);
and U21977 (N_21977,N_21066,N_21405);
and U21978 (N_21978,N_21347,N_21327);
xor U21979 (N_21979,N_21236,N_21089);
or U21980 (N_21980,N_21415,N_21287);
xor U21981 (N_21981,N_21011,N_21039);
or U21982 (N_21982,N_21358,N_21449);
nor U21983 (N_21983,N_21142,N_21141);
nor U21984 (N_21984,N_21277,N_21461);
nand U21985 (N_21985,N_21180,N_21095);
nand U21986 (N_21986,N_21275,N_21313);
nor U21987 (N_21987,N_21158,N_21047);
nand U21988 (N_21988,N_21347,N_21391);
nor U21989 (N_21989,N_21270,N_21088);
nor U21990 (N_21990,N_21337,N_21048);
nand U21991 (N_21991,N_21209,N_21151);
nor U21992 (N_21992,N_21059,N_21264);
or U21993 (N_21993,N_21288,N_21164);
and U21994 (N_21994,N_21101,N_21416);
xnor U21995 (N_21995,N_21031,N_21227);
nor U21996 (N_21996,N_21261,N_21111);
or U21997 (N_21997,N_21311,N_21142);
or U21998 (N_21998,N_21128,N_21263);
nor U21999 (N_21999,N_21147,N_21296);
nor U22000 (N_22000,N_21571,N_21956);
or U22001 (N_22001,N_21867,N_21868);
and U22002 (N_22002,N_21902,N_21653);
and U22003 (N_22003,N_21930,N_21924);
nor U22004 (N_22004,N_21741,N_21961);
and U22005 (N_22005,N_21797,N_21853);
nor U22006 (N_22006,N_21903,N_21700);
or U22007 (N_22007,N_21918,N_21845);
xnor U22008 (N_22008,N_21752,N_21732);
and U22009 (N_22009,N_21911,N_21955);
nand U22010 (N_22010,N_21729,N_21507);
and U22011 (N_22011,N_21977,N_21767);
nand U22012 (N_22012,N_21830,N_21884);
nand U22013 (N_22013,N_21703,N_21739);
or U22014 (N_22014,N_21899,N_21530);
xnor U22015 (N_22015,N_21652,N_21801);
and U22016 (N_22016,N_21621,N_21985);
and U22017 (N_22017,N_21788,N_21622);
xnor U22018 (N_22018,N_21642,N_21861);
nor U22019 (N_22019,N_21774,N_21560);
or U22020 (N_22020,N_21919,N_21921);
xnor U22021 (N_22021,N_21516,N_21886);
nand U22022 (N_22022,N_21912,N_21909);
or U22023 (N_22023,N_21719,N_21879);
nand U22024 (N_22024,N_21541,N_21689);
or U22025 (N_22025,N_21633,N_21900);
nor U22026 (N_22026,N_21979,N_21790);
or U22027 (N_22027,N_21957,N_21959);
xnor U22028 (N_22028,N_21614,N_21908);
or U22029 (N_22029,N_21818,N_21596);
and U22030 (N_22030,N_21546,N_21746);
xnor U22031 (N_22031,N_21984,N_21595);
nand U22032 (N_22032,N_21567,N_21603);
or U22033 (N_22033,N_21514,N_21898);
xnor U22034 (N_22034,N_21615,N_21625);
and U22035 (N_22035,N_21855,N_21577);
nand U22036 (N_22036,N_21630,N_21964);
nor U22037 (N_22037,N_21618,N_21883);
or U22038 (N_22038,N_21510,N_21518);
or U22039 (N_22039,N_21815,N_21755);
nor U22040 (N_22040,N_21584,N_21535);
nand U22041 (N_22041,N_21948,N_21509);
xor U22042 (N_22042,N_21929,N_21681);
xor U22043 (N_22043,N_21869,N_21728);
and U22044 (N_22044,N_21931,N_21655);
nand U22045 (N_22045,N_21798,N_21722);
or U22046 (N_22046,N_21573,N_21547);
nor U22047 (N_22047,N_21654,N_21940);
and U22048 (N_22048,N_21593,N_21831);
or U22049 (N_22049,N_21662,N_21785);
xor U22050 (N_22050,N_21678,N_21795);
nand U22051 (N_22051,N_21937,N_21674);
xnor U22052 (N_22052,N_21970,N_21742);
or U22053 (N_22053,N_21705,N_21713);
or U22054 (N_22054,N_21607,N_21968);
nand U22055 (N_22055,N_21664,N_21865);
and U22056 (N_22056,N_21646,N_21528);
nand U22057 (N_22057,N_21980,N_21562);
or U22058 (N_22058,N_21834,N_21843);
and U22059 (N_22059,N_21694,N_21574);
or U22060 (N_22060,N_21859,N_21780);
xnor U22061 (N_22061,N_21572,N_21597);
xnor U22062 (N_22062,N_21822,N_21692);
nand U22063 (N_22063,N_21975,N_21794);
and U22064 (N_22064,N_21896,N_21872);
or U22065 (N_22065,N_21952,N_21650);
nor U22066 (N_22066,N_21522,N_21992);
nor U22067 (N_22067,N_21950,N_21561);
nand U22068 (N_22068,N_21675,N_21928);
xnor U22069 (N_22069,N_21922,N_21761);
xor U22070 (N_22070,N_21871,N_21768);
nor U22071 (N_22071,N_21738,N_21698);
xor U22072 (N_22072,N_21876,N_21540);
and U22073 (N_22073,N_21582,N_21832);
nor U22074 (N_22074,N_21878,N_21640);
nor U22075 (N_22075,N_21925,N_21580);
nor U22076 (N_22076,N_21566,N_21661);
or U22077 (N_22077,N_21537,N_21519);
or U22078 (N_22078,N_21745,N_21691);
nor U22079 (N_22079,N_21555,N_21723);
and U22080 (N_22080,N_21808,N_21823);
nand U22081 (N_22081,N_21944,N_21881);
nor U22082 (N_22082,N_21647,N_21627);
and U22083 (N_22083,N_21586,N_21846);
or U22084 (N_22084,N_21943,N_21734);
and U22085 (N_22085,N_21799,N_21617);
nor U22086 (N_22086,N_21576,N_21524);
nand U22087 (N_22087,N_21765,N_21628);
nor U22088 (N_22088,N_21508,N_21666);
and U22089 (N_22089,N_21776,N_21987);
xor U22090 (N_22090,N_21836,N_21549);
xnor U22091 (N_22091,N_21915,N_21778);
nor U22092 (N_22092,N_21683,N_21641);
nor U22093 (N_22093,N_21564,N_21726);
or U22094 (N_22094,N_21880,N_21704);
or U22095 (N_22095,N_21707,N_21578);
nand U22096 (N_22096,N_21753,N_21645);
xnor U22097 (N_22097,N_21663,N_21671);
nand U22098 (N_22098,N_21803,N_21757);
nor U22099 (N_22099,N_21721,N_21552);
or U22100 (N_22100,N_21973,N_21766);
nor U22101 (N_22101,N_21825,N_21706);
xor U22102 (N_22102,N_21833,N_21720);
xnor U22103 (N_22103,N_21751,N_21620);
nand U22104 (N_22104,N_21747,N_21838);
nand U22105 (N_22105,N_21748,N_21553);
and U22106 (N_22106,N_21532,N_21544);
or U22107 (N_22107,N_21762,N_21737);
or U22108 (N_22108,N_21856,N_21775);
and U22109 (N_22109,N_21502,N_21520);
nor U22110 (N_22110,N_21895,N_21543);
xnor U22111 (N_22111,N_21538,N_21864);
or U22112 (N_22112,N_21995,N_21835);
or U22113 (N_22113,N_21634,N_21512);
nand U22114 (N_22114,N_21804,N_21974);
xor U22115 (N_22115,N_21682,N_21668);
nand U22116 (N_22116,N_21816,N_21550);
xor U22117 (N_22117,N_21810,N_21998);
or U22118 (N_22118,N_21887,N_21939);
or U22119 (N_22119,N_21960,N_21826);
xor U22120 (N_22120,N_21852,N_21500);
or U22121 (N_22121,N_21882,N_21923);
nand U22122 (N_22122,N_21904,N_21981);
or U22123 (N_22123,N_21773,N_21787);
or U22124 (N_22124,N_21701,N_21945);
xor U22125 (N_22125,N_21539,N_21972);
xor U22126 (N_22126,N_21659,N_21536);
nand U22127 (N_22127,N_21885,N_21559);
nand U22128 (N_22128,N_21933,N_21688);
and U22129 (N_22129,N_21932,N_21901);
and U22130 (N_22130,N_21534,N_21781);
nand U22131 (N_22131,N_21714,N_21840);
nand U22132 (N_22132,N_21828,N_21807);
nand U22133 (N_22133,N_21623,N_21809);
nor U22134 (N_22134,N_21632,N_21744);
xor U22135 (N_22135,N_21942,N_21926);
or U22136 (N_22136,N_21862,N_21783);
and U22137 (N_22137,N_21989,N_21777);
or U22138 (N_22138,N_21568,N_21731);
and U22139 (N_22139,N_21545,N_21847);
nor U22140 (N_22140,N_21583,N_21697);
xnor U22141 (N_22141,N_21565,N_21504);
xnor U22142 (N_22142,N_21938,N_21690);
xnor U22143 (N_22143,N_21730,N_21651);
xnor U22144 (N_22144,N_21563,N_21609);
and U22145 (N_22145,N_21616,N_21824);
xnor U22146 (N_22146,N_21837,N_21905);
and U22147 (N_22147,N_21758,N_21660);
or U22148 (N_22148,N_21643,N_21786);
and U22149 (N_22149,N_21699,N_21637);
and U22150 (N_22150,N_21849,N_21672);
xor U22151 (N_22151,N_21947,N_21990);
and U22152 (N_22152,N_21844,N_21892);
and U22153 (N_22153,N_21941,N_21986);
nor U22154 (N_22154,N_21715,N_21910);
xnor U22155 (N_22155,N_21648,N_21749);
nor U22156 (N_22156,N_21554,N_21695);
nand U22157 (N_22157,N_21588,N_21743);
or U22158 (N_22158,N_21604,N_21754);
or U22159 (N_22159,N_21579,N_21649);
xnor U22160 (N_22160,N_21687,N_21548);
or U22161 (N_22161,N_21907,N_21624);
xor U22162 (N_22162,N_21971,N_21954);
nand U22163 (N_22163,N_21599,N_21870);
nand U22164 (N_22164,N_21501,N_21812);
nor U22165 (N_22165,N_21521,N_21820);
nor U22166 (N_22166,N_21764,N_21791);
nor U22167 (N_22167,N_21811,N_21740);
xor U22168 (N_22168,N_21866,N_21965);
nand U22169 (N_22169,N_21779,N_21890);
or U22170 (N_22170,N_21893,N_21736);
and U22171 (N_22171,N_21605,N_21877);
xnor U22172 (N_22172,N_21503,N_21644);
or U22173 (N_22173,N_21934,N_21897);
and U22174 (N_22174,N_21669,N_21684);
or U22175 (N_22175,N_21805,N_21978);
nor U22176 (N_22176,N_21817,N_21608);
and U22177 (N_22177,N_21724,N_21581);
or U22178 (N_22178,N_21993,N_21750);
xor U22179 (N_22179,N_21629,N_21613);
xor U22180 (N_22180,N_21712,N_21966);
nand U22181 (N_22181,N_21569,N_21531);
and U22182 (N_22182,N_21917,N_21829);
nand U22183 (N_22183,N_21601,N_21958);
or U22184 (N_22184,N_21557,N_21770);
nor U22185 (N_22185,N_21927,N_21611);
nand U22186 (N_22186,N_21874,N_21889);
nand U22187 (N_22187,N_21710,N_21575);
or U22188 (N_22188,N_21725,N_21665);
nand U22189 (N_22189,N_21556,N_21619);
and U22190 (N_22190,N_21850,N_21696);
or U22191 (N_22191,N_21914,N_21991);
or U22192 (N_22192,N_21793,N_21686);
or U22193 (N_22193,N_21967,N_21983);
nand U22194 (N_22194,N_21506,N_21551);
nor U22195 (N_22195,N_21888,N_21594);
or U22196 (N_22196,N_21685,N_21670);
or U22197 (N_22197,N_21821,N_21631);
xor U22198 (N_22198,N_21784,N_21673);
nor U22199 (N_22199,N_21589,N_21936);
nor U22200 (N_22200,N_21760,N_21570);
and U22201 (N_22201,N_21679,N_21800);
nor U22202 (N_22202,N_21657,N_21935);
nor U22203 (N_22203,N_21946,N_21529);
nor U22204 (N_22204,N_21677,N_21598);
xnor U22205 (N_22205,N_21511,N_21558);
or U22206 (N_22206,N_21848,N_21708);
xnor U22207 (N_22207,N_21515,N_21875);
nor U22208 (N_22208,N_21894,N_21638);
or U22209 (N_22209,N_21612,N_21819);
xor U22210 (N_22210,N_21842,N_21769);
nand U22211 (N_22211,N_21996,N_21735);
nor U22212 (N_22212,N_21802,N_21827);
nand U22213 (N_22213,N_21709,N_21658);
and U22214 (N_22214,N_21860,N_21839);
and U22215 (N_22215,N_21756,N_21587);
xnor U22216 (N_22216,N_21988,N_21727);
and U22217 (N_22217,N_21527,N_21851);
and U22218 (N_22218,N_21676,N_21976);
xnor U22219 (N_22219,N_21763,N_21667);
nor U22220 (N_22220,N_21717,N_21982);
or U22221 (N_22221,N_21772,N_21792);
nor U22222 (N_22222,N_21916,N_21639);
and U22223 (N_22223,N_21542,N_21814);
or U22224 (N_22224,N_21963,N_21857);
nor U22225 (N_22225,N_21994,N_21863);
or U22226 (N_22226,N_21525,N_21962);
nor U22227 (N_22227,N_21759,N_21523);
and U22228 (N_22228,N_21891,N_21841);
xnor U22229 (N_22229,N_21969,N_21920);
xnor U22230 (N_22230,N_21610,N_21693);
and U22231 (N_22231,N_21636,N_21873);
or U22232 (N_22232,N_21606,N_21999);
nor U22233 (N_22233,N_21602,N_21906);
or U22234 (N_22234,N_21656,N_21951);
or U22235 (N_22235,N_21796,N_21813);
xnor U22236 (N_22236,N_21505,N_21953);
or U22237 (N_22237,N_21733,N_21533);
xnor U22238 (N_22238,N_21718,N_21591);
xnor U22239 (N_22239,N_21680,N_21592);
nor U22240 (N_22240,N_21635,N_21997);
nor U22241 (N_22241,N_21854,N_21782);
and U22242 (N_22242,N_21949,N_21711);
or U22243 (N_22243,N_21771,N_21626);
xor U22244 (N_22244,N_21585,N_21513);
xor U22245 (N_22245,N_21517,N_21590);
xnor U22246 (N_22246,N_21716,N_21526);
or U22247 (N_22247,N_21806,N_21858);
and U22248 (N_22248,N_21789,N_21600);
xnor U22249 (N_22249,N_21702,N_21913);
nor U22250 (N_22250,N_21892,N_21767);
nor U22251 (N_22251,N_21785,N_21660);
xnor U22252 (N_22252,N_21924,N_21788);
nand U22253 (N_22253,N_21726,N_21619);
or U22254 (N_22254,N_21618,N_21798);
xor U22255 (N_22255,N_21947,N_21705);
xor U22256 (N_22256,N_21914,N_21669);
nand U22257 (N_22257,N_21939,N_21620);
xnor U22258 (N_22258,N_21717,N_21857);
or U22259 (N_22259,N_21685,N_21500);
and U22260 (N_22260,N_21787,N_21638);
xor U22261 (N_22261,N_21913,N_21741);
xnor U22262 (N_22262,N_21915,N_21683);
and U22263 (N_22263,N_21877,N_21574);
and U22264 (N_22264,N_21919,N_21671);
nor U22265 (N_22265,N_21660,N_21973);
or U22266 (N_22266,N_21786,N_21609);
or U22267 (N_22267,N_21769,N_21682);
nor U22268 (N_22268,N_21949,N_21697);
xor U22269 (N_22269,N_21770,N_21626);
nand U22270 (N_22270,N_21847,N_21966);
or U22271 (N_22271,N_21809,N_21865);
xor U22272 (N_22272,N_21966,N_21982);
nor U22273 (N_22273,N_21999,N_21517);
nand U22274 (N_22274,N_21586,N_21675);
nor U22275 (N_22275,N_21992,N_21781);
or U22276 (N_22276,N_21733,N_21699);
and U22277 (N_22277,N_21958,N_21990);
or U22278 (N_22278,N_21686,N_21803);
or U22279 (N_22279,N_21582,N_21541);
or U22280 (N_22280,N_21966,N_21724);
and U22281 (N_22281,N_21528,N_21759);
or U22282 (N_22282,N_21967,N_21930);
nor U22283 (N_22283,N_21683,N_21839);
nor U22284 (N_22284,N_21620,N_21529);
and U22285 (N_22285,N_21980,N_21773);
nor U22286 (N_22286,N_21961,N_21927);
nor U22287 (N_22287,N_21580,N_21593);
nor U22288 (N_22288,N_21644,N_21714);
or U22289 (N_22289,N_21838,N_21813);
xnor U22290 (N_22290,N_21804,N_21983);
and U22291 (N_22291,N_21535,N_21706);
nor U22292 (N_22292,N_21501,N_21833);
xor U22293 (N_22293,N_21808,N_21810);
xor U22294 (N_22294,N_21647,N_21946);
and U22295 (N_22295,N_21637,N_21647);
and U22296 (N_22296,N_21982,N_21898);
nand U22297 (N_22297,N_21618,N_21533);
or U22298 (N_22298,N_21832,N_21844);
nand U22299 (N_22299,N_21501,N_21690);
xnor U22300 (N_22300,N_21667,N_21658);
nor U22301 (N_22301,N_21662,N_21796);
or U22302 (N_22302,N_21756,N_21534);
or U22303 (N_22303,N_21558,N_21605);
and U22304 (N_22304,N_21939,N_21597);
or U22305 (N_22305,N_21950,N_21761);
or U22306 (N_22306,N_21573,N_21719);
nor U22307 (N_22307,N_21565,N_21765);
or U22308 (N_22308,N_21799,N_21621);
xnor U22309 (N_22309,N_21617,N_21956);
or U22310 (N_22310,N_21615,N_21944);
xnor U22311 (N_22311,N_21829,N_21712);
nor U22312 (N_22312,N_21920,N_21571);
nor U22313 (N_22313,N_21749,N_21669);
or U22314 (N_22314,N_21728,N_21577);
nand U22315 (N_22315,N_21690,N_21506);
nor U22316 (N_22316,N_21822,N_21820);
xnor U22317 (N_22317,N_21669,N_21862);
nand U22318 (N_22318,N_21959,N_21567);
and U22319 (N_22319,N_21877,N_21522);
or U22320 (N_22320,N_21652,N_21841);
xor U22321 (N_22321,N_21827,N_21602);
nor U22322 (N_22322,N_21761,N_21914);
and U22323 (N_22323,N_21986,N_21876);
or U22324 (N_22324,N_21590,N_21557);
nor U22325 (N_22325,N_21518,N_21878);
xnor U22326 (N_22326,N_21667,N_21715);
and U22327 (N_22327,N_21944,N_21865);
or U22328 (N_22328,N_21993,N_21836);
nand U22329 (N_22329,N_21597,N_21920);
nand U22330 (N_22330,N_21900,N_21744);
or U22331 (N_22331,N_21979,N_21917);
or U22332 (N_22332,N_21581,N_21893);
nand U22333 (N_22333,N_21683,N_21503);
xnor U22334 (N_22334,N_21705,N_21913);
or U22335 (N_22335,N_21624,N_21766);
nand U22336 (N_22336,N_21870,N_21927);
nor U22337 (N_22337,N_21825,N_21533);
nand U22338 (N_22338,N_21726,N_21714);
nor U22339 (N_22339,N_21627,N_21663);
nor U22340 (N_22340,N_21850,N_21506);
or U22341 (N_22341,N_21934,N_21851);
and U22342 (N_22342,N_21801,N_21770);
and U22343 (N_22343,N_21784,N_21574);
and U22344 (N_22344,N_21780,N_21503);
and U22345 (N_22345,N_21858,N_21524);
nor U22346 (N_22346,N_21693,N_21799);
xor U22347 (N_22347,N_21673,N_21539);
nor U22348 (N_22348,N_21971,N_21530);
nor U22349 (N_22349,N_21968,N_21869);
or U22350 (N_22350,N_21826,N_21853);
nor U22351 (N_22351,N_21678,N_21707);
nand U22352 (N_22352,N_21948,N_21950);
xor U22353 (N_22353,N_21777,N_21585);
or U22354 (N_22354,N_21502,N_21948);
or U22355 (N_22355,N_21594,N_21818);
xor U22356 (N_22356,N_21890,N_21727);
or U22357 (N_22357,N_21563,N_21733);
or U22358 (N_22358,N_21914,N_21969);
xor U22359 (N_22359,N_21822,N_21589);
or U22360 (N_22360,N_21611,N_21536);
nor U22361 (N_22361,N_21679,N_21880);
and U22362 (N_22362,N_21551,N_21885);
and U22363 (N_22363,N_21677,N_21984);
nor U22364 (N_22364,N_21690,N_21763);
nor U22365 (N_22365,N_21779,N_21861);
nand U22366 (N_22366,N_21712,N_21941);
nand U22367 (N_22367,N_21982,N_21937);
and U22368 (N_22368,N_21514,N_21832);
nor U22369 (N_22369,N_21576,N_21876);
nor U22370 (N_22370,N_21846,N_21771);
and U22371 (N_22371,N_21967,N_21803);
xor U22372 (N_22372,N_21785,N_21515);
and U22373 (N_22373,N_21664,N_21723);
xor U22374 (N_22374,N_21543,N_21909);
and U22375 (N_22375,N_21731,N_21540);
or U22376 (N_22376,N_21972,N_21576);
or U22377 (N_22377,N_21862,N_21615);
and U22378 (N_22378,N_21771,N_21865);
xnor U22379 (N_22379,N_21788,N_21923);
nor U22380 (N_22380,N_21796,N_21672);
or U22381 (N_22381,N_21987,N_21829);
xor U22382 (N_22382,N_21903,N_21711);
nand U22383 (N_22383,N_21602,N_21616);
nor U22384 (N_22384,N_21834,N_21527);
and U22385 (N_22385,N_21698,N_21557);
xnor U22386 (N_22386,N_21897,N_21832);
or U22387 (N_22387,N_21518,N_21786);
xnor U22388 (N_22388,N_21819,N_21930);
nand U22389 (N_22389,N_21855,N_21779);
nor U22390 (N_22390,N_21738,N_21901);
nor U22391 (N_22391,N_21675,N_21940);
or U22392 (N_22392,N_21844,N_21880);
nand U22393 (N_22393,N_21800,N_21697);
nand U22394 (N_22394,N_21620,N_21641);
nand U22395 (N_22395,N_21892,N_21565);
or U22396 (N_22396,N_21683,N_21746);
nor U22397 (N_22397,N_21751,N_21656);
nand U22398 (N_22398,N_21531,N_21573);
nand U22399 (N_22399,N_21591,N_21916);
xor U22400 (N_22400,N_21531,N_21837);
or U22401 (N_22401,N_21769,N_21917);
nor U22402 (N_22402,N_21886,N_21974);
nor U22403 (N_22403,N_21661,N_21905);
or U22404 (N_22404,N_21925,N_21902);
nor U22405 (N_22405,N_21699,N_21969);
and U22406 (N_22406,N_21621,N_21653);
xor U22407 (N_22407,N_21620,N_21516);
and U22408 (N_22408,N_21740,N_21502);
or U22409 (N_22409,N_21547,N_21540);
or U22410 (N_22410,N_21559,N_21763);
and U22411 (N_22411,N_21867,N_21956);
and U22412 (N_22412,N_21615,N_21566);
or U22413 (N_22413,N_21652,N_21839);
xor U22414 (N_22414,N_21560,N_21925);
or U22415 (N_22415,N_21887,N_21504);
nand U22416 (N_22416,N_21501,N_21988);
nand U22417 (N_22417,N_21613,N_21524);
or U22418 (N_22418,N_21869,N_21631);
xnor U22419 (N_22419,N_21735,N_21774);
and U22420 (N_22420,N_21753,N_21781);
or U22421 (N_22421,N_21910,N_21764);
xor U22422 (N_22422,N_21657,N_21999);
and U22423 (N_22423,N_21624,N_21982);
xnor U22424 (N_22424,N_21885,N_21974);
nor U22425 (N_22425,N_21811,N_21581);
nand U22426 (N_22426,N_21786,N_21771);
xor U22427 (N_22427,N_21765,N_21883);
xnor U22428 (N_22428,N_21733,N_21761);
or U22429 (N_22429,N_21976,N_21961);
or U22430 (N_22430,N_21609,N_21993);
nor U22431 (N_22431,N_21504,N_21551);
xor U22432 (N_22432,N_21701,N_21504);
xor U22433 (N_22433,N_21800,N_21686);
or U22434 (N_22434,N_21552,N_21974);
xnor U22435 (N_22435,N_21622,N_21914);
nor U22436 (N_22436,N_21610,N_21703);
and U22437 (N_22437,N_21507,N_21852);
or U22438 (N_22438,N_21909,N_21708);
xor U22439 (N_22439,N_21679,N_21625);
and U22440 (N_22440,N_21765,N_21954);
and U22441 (N_22441,N_21899,N_21679);
xor U22442 (N_22442,N_21853,N_21798);
nor U22443 (N_22443,N_21808,N_21961);
and U22444 (N_22444,N_21619,N_21749);
and U22445 (N_22445,N_21948,N_21872);
nand U22446 (N_22446,N_21976,N_21791);
or U22447 (N_22447,N_21686,N_21890);
and U22448 (N_22448,N_21860,N_21674);
nor U22449 (N_22449,N_21541,N_21540);
or U22450 (N_22450,N_21754,N_21892);
xnor U22451 (N_22451,N_21706,N_21618);
or U22452 (N_22452,N_21860,N_21656);
xor U22453 (N_22453,N_21593,N_21971);
nor U22454 (N_22454,N_21978,N_21919);
nand U22455 (N_22455,N_21984,N_21653);
and U22456 (N_22456,N_21549,N_21916);
or U22457 (N_22457,N_21857,N_21666);
xor U22458 (N_22458,N_21768,N_21880);
and U22459 (N_22459,N_21740,N_21728);
and U22460 (N_22460,N_21791,N_21843);
and U22461 (N_22461,N_21533,N_21969);
xnor U22462 (N_22462,N_21605,N_21848);
xnor U22463 (N_22463,N_21538,N_21513);
and U22464 (N_22464,N_21527,N_21913);
nor U22465 (N_22465,N_21521,N_21909);
or U22466 (N_22466,N_21755,N_21720);
nand U22467 (N_22467,N_21897,N_21681);
nor U22468 (N_22468,N_21556,N_21567);
nand U22469 (N_22469,N_21765,N_21833);
or U22470 (N_22470,N_21768,N_21716);
xnor U22471 (N_22471,N_21702,N_21906);
and U22472 (N_22472,N_21608,N_21923);
xnor U22473 (N_22473,N_21848,N_21809);
nand U22474 (N_22474,N_21788,N_21771);
nand U22475 (N_22475,N_21778,N_21865);
or U22476 (N_22476,N_21730,N_21970);
nand U22477 (N_22477,N_21635,N_21873);
xor U22478 (N_22478,N_21506,N_21717);
and U22479 (N_22479,N_21713,N_21643);
nor U22480 (N_22480,N_21688,N_21769);
nor U22481 (N_22481,N_21987,N_21831);
nor U22482 (N_22482,N_21668,N_21615);
xor U22483 (N_22483,N_21575,N_21685);
and U22484 (N_22484,N_21736,N_21660);
nor U22485 (N_22485,N_21653,N_21767);
nand U22486 (N_22486,N_21842,N_21830);
nand U22487 (N_22487,N_21602,N_21860);
nor U22488 (N_22488,N_21849,N_21679);
nand U22489 (N_22489,N_21592,N_21904);
or U22490 (N_22490,N_21847,N_21721);
or U22491 (N_22491,N_21997,N_21718);
xnor U22492 (N_22492,N_21930,N_21659);
nor U22493 (N_22493,N_21835,N_21722);
nor U22494 (N_22494,N_21531,N_21592);
and U22495 (N_22495,N_21665,N_21615);
nor U22496 (N_22496,N_21731,N_21950);
nand U22497 (N_22497,N_21581,N_21866);
or U22498 (N_22498,N_21600,N_21564);
and U22499 (N_22499,N_21721,N_21930);
or U22500 (N_22500,N_22236,N_22191);
or U22501 (N_22501,N_22472,N_22018);
xnor U22502 (N_22502,N_22494,N_22287);
or U22503 (N_22503,N_22117,N_22224);
or U22504 (N_22504,N_22248,N_22484);
and U22505 (N_22505,N_22405,N_22298);
and U22506 (N_22506,N_22193,N_22458);
xnor U22507 (N_22507,N_22231,N_22065);
nor U22508 (N_22508,N_22032,N_22017);
nand U22509 (N_22509,N_22415,N_22040);
xnor U22510 (N_22510,N_22085,N_22064);
and U22511 (N_22511,N_22079,N_22159);
and U22512 (N_22512,N_22344,N_22100);
or U22513 (N_22513,N_22277,N_22376);
or U22514 (N_22514,N_22206,N_22075);
nor U22515 (N_22515,N_22007,N_22271);
or U22516 (N_22516,N_22073,N_22135);
nand U22517 (N_22517,N_22011,N_22350);
and U22518 (N_22518,N_22255,N_22340);
nor U22519 (N_22519,N_22365,N_22378);
and U22520 (N_22520,N_22414,N_22299);
nand U22521 (N_22521,N_22057,N_22004);
xnor U22522 (N_22522,N_22456,N_22041);
xor U22523 (N_22523,N_22078,N_22264);
xor U22524 (N_22524,N_22269,N_22164);
and U22525 (N_22525,N_22058,N_22323);
nand U22526 (N_22526,N_22253,N_22145);
nor U22527 (N_22527,N_22161,N_22325);
and U22528 (N_22528,N_22156,N_22439);
or U22529 (N_22529,N_22295,N_22094);
nor U22530 (N_22530,N_22015,N_22397);
or U22531 (N_22531,N_22238,N_22374);
or U22532 (N_22532,N_22256,N_22444);
and U22533 (N_22533,N_22211,N_22370);
nand U22534 (N_22534,N_22476,N_22385);
and U22535 (N_22535,N_22357,N_22321);
nor U22536 (N_22536,N_22436,N_22364);
or U22537 (N_22537,N_22251,N_22177);
nand U22538 (N_22538,N_22190,N_22317);
xor U22539 (N_22539,N_22309,N_22022);
xor U22540 (N_22540,N_22339,N_22398);
or U22541 (N_22541,N_22390,N_22074);
or U22542 (N_22542,N_22025,N_22250);
xor U22543 (N_22543,N_22132,N_22194);
and U22544 (N_22544,N_22128,N_22375);
or U22545 (N_22545,N_22146,N_22147);
nand U22546 (N_22546,N_22335,N_22400);
and U22547 (N_22547,N_22380,N_22168);
and U22548 (N_22548,N_22438,N_22288);
or U22549 (N_22549,N_22417,N_22113);
nand U22550 (N_22550,N_22054,N_22282);
xnor U22551 (N_22551,N_22221,N_22105);
or U22552 (N_22552,N_22173,N_22227);
nor U22553 (N_22553,N_22188,N_22123);
and U22554 (N_22554,N_22432,N_22349);
and U22555 (N_22555,N_22242,N_22420);
or U22556 (N_22556,N_22297,N_22047);
xor U22557 (N_22557,N_22216,N_22272);
xor U22558 (N_22558,N_22151,N_22284);
nor U22559 (N_22559,N_22363,N_22412);
or U22560 (N_22560,N_22329,N_22495);
or U22561 (N_22561,N_22419,N_22258);
xnor U22562 (N_22562,N_22210,N_22052);
nor U22563 (N_22563,N_22289,N_22245);
or U22564 (N_22564,N_22394,N_22279);
and U22565 (N_22565,N_22172,N_22174);
nand U22566 (N_22566,N_22071,N_22268);
and U22567 (N_22567,N_22285,N_22209);
xnor U22568 (N_22568,N_22450,N_22372);
nand U22569 (N_22569,N_22232,N_22498);
xnor U22570 (N_22570,N_22154,N_22158);
or U22571 (N_22571,N_22067,N_22008);
nand U22572 (N_22572,N_22430,N_22120);
xnor U22573 (N_22573,N_22097,N_22036);
or U22574 (N_22574,N_22316,N_22477);
nor U22575 (N_22575,N_22028,N_22333);
nand U22576 (N_22576,N_22169,N_22009);
and U22577 (N_22577,N_22000,N_22452);
xnor U22578 (N_22578,N_22114,N_22108);
or U22579 (N_22579,N_22142,N_22343);
nor U22580 (N_22580,N_22387,N_22134);
nor U22581 (N_22581,N_22220,N_22381);
and U22582 (N_22582,N_22042,N_22005);
and U22583 (N_22583,N_22267,N_22384);
nand U22584 (N_22584,N_22373,N_22021);
and U22585 (N_22585,N_22263,N_22468);
nand U22586 (N_22586,N_22010,N_22337);
nand U22587 (N_22587,N_22491,N_22121);
xor U22588 (N_22588,N_22129,N_22424);
nand U22589 (N_22589,N_22334,N_22214);
nor U22590 (N_22590,N_22493,N_22081);
or U22591 (N_22591,N_22001,N_22207);
and U22592 (N_22592,N_22311,N_22240);
xnor U22593 (N_22593,N_22141,N_22422);
nand U22594 (N_22594,N_22237,N_22006);
xor U22595 (N_22595,N_22362,N_22396);
and U22596 (N_22596,N_22192,N_22433);
xnor U22597 (N_22597,N_22171,N_22201);
nor U22598 (N_22598,N_22093,N_22459);
xnor U22599 (N_22599,N_22249,N_22478);
or U22600 (N_22600,N_22087,N_22103);
or U22601 (N_22601,N_22002,N_22109);
xor U22602 (N_22602,N_22356,N_22019);
nand U22603 (N_22603,N_22359,N_22187);
and U22604 (N_22604,N_22170,N_22300);
or U22605 (N_22605,N_22229,N_22106);
or U22606 (N_22606,N_22195,N_22204);
nand U22607 (N_22607,N_22320,N_22104);
and U22608 (N_22608,N_22274,N_22455);
nor U22609 (N_22609,N_22386,N_22425);
and U22610 (N_22610,N_22149,N_22198);
nor U22611 (N_22611,N_22399,N_22395);
nor U22612 (N_22612,N_22180,N_22096);
xor U22613 (N_22613,N_22358,N_22441);
and U22614 (N_22614,N_22199,N_22030);
and U22615 (N_22615,N_22013,N_22163);
xor U22616 (N_22616,N_22102,N_22303);
xor U22617 (N_22617,N_22202,N_22083);
and U22618 (N_22618,N_22377,N_22461);
nor U22619 (N_22619,N_22186,N_22427);
xnor U22620 (N_22620,N_22301,N_22403);
nand U22621 (N_22621,N_22314,N_22341);
or U22622 (N_22622,N_22404,N_22310);
nand U22623 (N_22623,N_22391,N_22080);
and U22624 (N_22624,N_22185,N_22489);
nor U22625 (N_22625,N_22166,N_22487);
or U22626 (N_22626,N_22176,N_22235);
nor U22627 (N_22627,N_22020,N_22345);
nor U22628 (N_22628,N_22184,N_22084);
nor U22629 (N_22629,N_22228,N_22259);
and U22630 (N_22630,N_22247,N_22382);
nand U22631 (N_22631,N_22283,N_22055);
nand U22632 (N_22632,N_22098,N_22127);
or U22633 (N_22633,N_22411,N_22347);
nor U22634 (N_22634,N_22153,N_22012);
or U22635 (N_22635,N_22175,N_22024);
and U22636 (N_22636,N_22150,N_22183);
nand U22637 (N_22637,N_22046,N_22144);
nand U22638 (N_22638,N_22429,N_22077);
and U22639 (N_22639,N_22355,N_22125);
nor U22640 (N_22640,N_22124,N_22203);
nor U22641 (N_22641,N_22312,N_22239);
and U22642 (N_22642,N_22157,N_22082);
nand U22643 (N_22643,N_22070,N_22446);
xnor U22644 (N_22644,N_22291,N_22076);
or U22645 (N_22645,N_22112,N_22016);
nand U22646 (N_22646,N_22490,N_22467);
nand U22647 (N_22647,N_22421,N_22407);
nor U22648 (N_22648,N_22293,N_22483);
nor U22649 (N_22649,N_22039,N_22331);
xnor U22650 (N_22650,N_22034,N_22252);
nand U22651 (N_22651,N_22475,N_22230);
nor U22652 (N_22652,N_22118,N_22482);
nand U22653 (N_22653,N_22029,N_22060);
and U22654 (N_22654,N_22049,N_22217);
xnor U22655 (N_22655,N_22480,N_22089);
and U22656 (N_22656,N_22449,N_22465);
nor U22657 (N_22657,N_22371,N_22069);
and U22658 (N_22658,N_22448,N_22296);
nor U22659 (N_22659,N_22315,N_22426);
and U22660 (N_22660,N_22457,N_22179);
xor U22661 (N_22661,N_22160,N_22326);
or U22662 (N_22662,N_22479,N_22481);
nand U22663 (N_22663,N_22402,N_22416);
or U22664 (N_22664,N_22434,N_22244);
nor U22665 (N_22665,N_22401,N_22338);
nor U22666 (N_22666,N_22393,N_22473);
xor U22667 (N_22667,N_22418,N_22066);
and U22668 (N_22668,N_22212,N_22437);
xor U22669 (N_22669,N_22361,N_22383);
or U22670 (N_22670,N_22027,N_22360);
xor U22671 (N_22671,N_22306,N_22471);
nand U22672 (N_22672,N_22140,N_22409);
xor U22673 (N_22673,N_22023,N_22435);
nand U22674 (N_22674,N_22213,N_22031);
nor U22675 (N_22675,N_22068,N_22290);
or U22676 (N_22676,N_22332,N_22053);
and U22677 (N_22677,N_22178,N_22155);
nor U22678 (N_22678,N_22136,N_22059);
xor U22679 (N_22679,N_22408,N_22095);
or U22680 (N_22680,N_22351,N_22307);
xor U22681 (N_22681,N_22276,N_22318);
nor U22682 (N_22682,N_22225,N_22045);
or U22683 (N_22683,N_22428,N_22138);
or U22684 (N_22684,N_22454,N_22189);
xnor U22685 (N_22685,N_22111,N_22280);
nor U22686 (N_22686,N_22262,N_22092);
nand U22687 (N_22687,N_22392,N_22469);
and U22688 (N_22688,N_22143,N_22302);
nor U22689 (N_22689,N_22099,N_22308);
xor U22690 (N_22690,N_22126,N_22453);
nand U22691 (N_22691,N_22003,N_22130);
nor U22692 (N_22692,N_22026,N_22200);
nor U22693 (N_22693,N_22485,N_22051);
nor U22694 (N_22694,N_22443,N_22165);
nor U22695 (N_22695,N_22197,N_22035);
xnor U22696 (N_22696,N_22014,N_22499);
or U22697 (N_22697,N_22336,N_22257);
nand U22698 (N_22698,N_22223,N_22327);
nor U22699 (N_22699,N_22226,N_22037);
and U22700 (N_22700,N_22261,N_22440);
nor U22701 (N_22701,N_22265,N_22462);
nand U22702 (N_22702,N_22088,N_22451);
nor U22703 (N_22703,N_22460,N_22496);
and U22704 (N_22704,N_22196,N_22294);
and U22705 (N_22705,N_22050,N_22497);
nor U22706 (N_22706,N_22222,N_22474);
nand U22707 (N_22707,N_22354,N_22205);
or U22708 (N_22708,N_22061,N_22445);
and U22709 (N_22709,N_22324,N_22167);
nand U22710 (N_22710,N_22389,N_22208);
and U22711 (N_22711,N_22313,N_22043);
nor U22712 (N_22712,N_22260,N_22218);
nor U22713 (N_22713,N_22246,N_22492);
and U22714 (N_22714,N_22148,N_22342);
nor U22715 (N_22715,N_22278,N_22233);
xor U22716 (N_22716,N_22116,N_22319);
and U22717 (N_22717,N_22072,N_22266);
nor U22718 (N_22718,N_22447,N_22322);
or U22719 (N_22719,N_22431,N_22215);
and U22720 (N_22720,N_22330,N_22466);
and U22721 (N_22721,N_22273,N_22348);
and U22722 (N_22722,N_22056,N_22275);
nor U22723 (N_22723,N_22038,N_22090);
and U22724 (N_22724,N_22423,N_22352);
or U22725 (N_22725,N_22388,N_22486);
nor U22726 (N_22726,N_22181,N_22328);
nor U22727 (N_22727,N_22131,N_22044);
nor U22728 (N_22728,N_22270,N_22346);
nor U22729 (N_22729,N_22488,N_22292);
nand U22730 (N_22730,N_22286,N_22254);
xor U22731 (N_22731,N_22139,N_22368);
and U22732 (N_22732,N_22048,N_22182);
nand U22733 (N_22733,N_22162,N_22367);
nand U22734 (N_22734,N_22406,N_22234);
nand U22735 (N_22735,N_22152,N_22133);
or U22736 (N_22736,N_22219,N_22243);
or U22737 (N_22737,N_22304,N_22463);
and U22738 (N_22738,N_22086,N_22033);
nor U22739 (N_22739,N_22119,N_22410);
and U22740 (N_22740,N_22353,N_22063);
nand U22741 (N_22741,N_22110,N_22241);
nor U22742 (N_22742,N_22062,N_22122);
xnor U22743 (N_22743,N_22464,N_22281);
nor U22744 (N_22744,N_22369,N_22305);
and U22745 (N_22745,N_22115,N_22379);
xnor U22746 (N_22746,N_22413,N_22470);
or U22747 (N_22747,N_22101,N_22366);
xor U22748 (N_22748,N_22442,N_22091);
nand U22749 (N_22749,N_22107,N_22137);
nand U22750 (N_22750,N_22122,N_22073);
xor U22751 (N_22751,N_22398,N_22353);
and U22752 (N_22752,N_22407,N_22322);
xor U22753 (N_22753,N_22070,N_22195);
and U22754 (N_22754,N_22442,N_22469);
nor U22755 (N_22755,N_22206,N_22142);
nand U22756 (N_22756,N_22378,N_22075);
xnor U22757 (N_22757,N_22282,N_22152);
xnor U22758 (N_22758,N_22433,N_22293);
nand U22759 (N_22759,N_22482,N_22351);
and U22760 (N_22760,N_22011,N_22163);
nor U22761 (N_22761,N_22480,N_22420);
or U22762 (N_22762,N_22014,N_22302);
xor U22763 (N_22763,N_22318,N_22058);
nand U22764 (N_22764,N_22418,N_22291);
xor U22765 (N_22765,N_22451,N_22424);
xor U22766 (N_22766,N_22238,N_22000);
nor U22767 (N_22767,N_22307,N_22400);
nor U22768 (N_22768,N_22168,N_22372);
nand U22769 (N_22769,N_22179,N_22027);
nand U22770 (N_22770,N_22162,N_22112);
xor U22771 (N_22771,N_22248,N_22432);
xnor U22772 (N_22772,N_22179,N_22140);
or U22773 (N_22773,N_22407,N_22120);
and U22774 (N_22774,N_22413,N_22017);
or U22775 (N_22775,N_22216,N_22223);
nor U22776 (N_22776,N_22153,N_22245);
nor U22777 (N_22777,N_22412,N_22328);
xor U22778 (N_22778,N_22337,N_22253);
and U22779 (N_22779,N_22091,N_22016);
or U22780 (N_22780,N_22342,N_22274);
and U22781 (N_22781,N_22309,N_22301);
or U22782 (N_22782,N_22105,N_22000);
or U22783 (N_22783,N_22331,N_22014);
xor U22784 (N_22784,N_22096,N_22245);
nand U22785 (N_22785,N_22219,N_22125);
xnor U22786 (N_22786,N_22380,N_22386);
or U22787 (N_22787,N_22475,N_22286);
xor U22788 (N_22788,N_22025,N_22026);
nor U22789 (N_22789,N_22240,N_22152);
or U22790 (N_22790,N_22277,N_22460);
nand U22791 (N_22791,N_22289,N_22302);
xnor U22792 (N_22792,N_22137,N_22226);
and U22793 (N_22793,N_22485,N_22034);
nor U22794 (N_22794,N_22268,N_22189);
nand U22795 (N_22795,N_22325,N_22344);
nor U22796 (N_22796,N_22015,N_22302);
or U22797 (N_22797,N_22073,N_22441);
and U22798 (N_22798,N_22388,N_22050);
and U22799 (N_22799,N_22454,N_22184);
and U22800 (N_22800,N_22148,N_22243);
nor U22801 (N_22801,N_22022,N_22349);
nand U22802 (N_22802,N_22210,N_22220);
and U22803 (N_22803,N_22398,N_22312);
xnor U22804 (N_22804,N_22042,N_22423);
nor U22805 (N_22805,N_22238,N_22285);
and U22806 (N_22806,N_22250,N_22350);
nand U22807 (N_22807,N_22240,N_22156);
xor U22808 (N_22808,N_22093,N_22212);
nand U22809 (N_22809,N_22089,N_22496);
and U22810 (N_22810,N_22103,N_22291);
nor U22811 (N_22811,N_22071,N_22326);
nor U22812 (N_22812,N_22458,N_22276);
and U22813 (N_22813,N_22300,N_22013);
nor U22814 (N_22814,N_22407,N_22194);
nand U22815 (N_22815,N_22453,N_22021);
nor U22816 (N_22816,N_22135,N_22091);
and U22817 (N_22817,N_22379,N_22330);
nor U22818 (N_22818,N_22024,N_22049);
or U22819 (N_22819,N_22304,N_22405);
nor U22820 (N_22820,N_22254,N_22119);
or U22821 (N_22821,N_22025,N_22283);
and U22822 (N_22822,N_22079,N_22190);
nor U22823 (N_22823,N_22012,N_22368);
and U22824 (N_22824,N_22487,N_22421);
nand U22825 (N_22825,N_22355,N_22037);
and U22826 (N_22826,N_22498,N_22477);
nand U22827 (N_22827,N_22357,N_22187);
and U22828 (N_22828,N_22062,N_22015);
nand U22829 (N_22829,N_22366,N_22338);
xnor U22830 (N_22830,N_22006,N_22130);
xor U22831 (N_22831,N_22470,N_22360);
nand U22832 (N_22832,N_22289,N_22356);
xor U22833 (N_22833,N_22091,N_22260);
and U22834 (N_22834,N_22138,N_22324);
nand U22835 (N_22835,N_22296,N_22305);
xnor U22836 (N_22836,N_22343,N_22207);
and U22837 (N_22837,N_22038,N_22011);
nand U22838 (N_22838,N_22189,N_22412);
and U22839 (N_22839,N_22340,N_22086);
nand U22840 (N_22840,N_22411,N_22146);
xor U22841 (N_22841,N_22375,N_22194);
nand U22842 (N_22842,N_22417,N_22069);
nand U22843 (N_22843,N_22473,N_22058);
or U22844 (N_22844,N_22445,N_22178);
xnor U22845 (N_22845,N_22327,N_22288);
xor U22846 (N_22846,N_22040,N_22115);
xnor U22847 (N_22847,N_22363,N_22403);
and U22848 (N_22848,N_22028,N_22087);
nor U22849 (N_22849,N_22394,N_22493);
or U22850 (N_22850,N_22074,N_22114);
nand U22851 (N_22851,N_22412,N_22198);
or U22852 (N_22852,N_22197,N_22103);
and U22853 (N_22853,N_22079,N_22292);
nand U22854 (N_22854,N_22115,N_22158);
nand U22855 (N_22855,N_22240,N_22185);
xnor U22856 (N_22856,N_22012,N_22038);
nor U22857 (N_22857,N_22174,N_22111);
nor U22858 (N_22858,N_22352,N_22269);
nor U22859 (N_22859,N_22324,N_22017);
xor U22860 (N_22860,N_22409,N_22459);
xnor U22861 (N_22861,N_22464,N_22220);
nor U22862 (N_22862,N_22392,N_22312);
xnor U22863 (N_22863,N_22024,N_22195);
and U22864 (N_22864,N_22237,N_22303);
or U22865 (N_22865,N_22091,N_22031);
and U22866 (N_22866,N_22273,N_22387);
xnor U22867 (N_22867,N_22418,N_22407);
and U22868 (N_22868,N_22339,N_22006);
xnor U22869 (N_22869,N_22190,N_22212);
nand U22870 (N_22870,N_22221,N_22248);
or U22871 (N_22871,N_22086,N_22315);
xnor U22872 (N_22872,N_22126,N_22144);
xor U22873 (N_22873,N_22232,N_22357);
or U22874 (N_22874,N_22108,N_22454);
nand U22875 (N_22875,N_22168,N_22155);
nor U22876 (N_22876,N_22327,N_22141);
nand U22877 (N_22877,N_22414,N_22334);
and U22878 (N_22878,N_22008,N_22171);
or U22879 (N_22879,N_22274,N_22436);
or U22880 (N_22880,N_22074,N_22138);
nand U22881 (N_22881,N_22180,N_22366);
nand U22882 (N_22882,N_22469,N_22282);
or U22883 (N_22883,N_22394,N_22287);
nor U22884 (N_22884,N_22144,N_22383);
or U22885 (N_22885,N_22336,N_22032);
or U22886 (N_22886,N_22258,N_22154);
or U22887 (N_22887,N_22164,N_22338);
or U22888 (N_22888,N_22193,N_22034);
or U22889 (N_22889,N_22102,N_22413);
nor U22890 (N_22890,N_22318,N_22168);
nand U22891 (N_22891,N_22213,N_22226);
nor U22892 (N_22892,N_22345,N_22455);
nand U22893 (N_22893,N_22153,N_22260);
nor U22894 (N_22894,N_22128,N_22334);
nor U22895 (N_22895,N_22233,N_22415);
nand U22896 (N_22896,N_22244,N_22392);
xor U22897 (N_22897,N_22429,N_22153);
or U22898 (N_22898,N_22032,N_22174);
and U22899 (N_22899,N_22156,N_22146);
nand U22900 (N_22900,N_22126,N_22267);
or U22901 (N_22901,N_22444,N_22068);
or U22902 (N_22902,N_22346,N_22160);
or U22903 (N_22903,N_22091,N_22456);
nor U22904 (N_22904,N_22071,N_22483);
or U22905 (N_22905,N_22172,N_22102);
nand U22906 (N_22906,N_22403,N_22157);
xnor U22907 (N_22907,N_22178,N_22490);
or U22908 (N_22908,N_22368,N_22437);
and U22909 (N_22909,N_22099,N_22476);
nand U22910 (N_22910,N_22478,N_22329);
or U22911 (N_22911,N_22184,N_22287);
nor U22912 (N_22912,N_22426,N_22128);
nand U22913 (N_22913,N_22137,N_22099);
or U22914 (N_22914,N_22211,N_22169);
xor U22915 (N_22915,N_22251,N_22377);
xnor U22916 (N_22916,N_22366,N_22086);
nand U22917 (N_22917,N_22320,N_22075);
and U22918 (N_22918,N_22415,N_22381);
nand U22919 (N_22919,N_22180,N_22309);
or U22920 (N_22920,N_22204,N_22068);
nor U22921 (N_22921,N_22257,N_22028);
nor U22922 (N_22922,N_22457,N_22335);
or U22923 (N_22923,N_22203,N_22474);
and U22924 (N_22924,N_22429,N_22155);
and U22925 (N_22925,N_22388,N_22125);
nand U22926 (N_22926,N_22348,N_22127);
nand U22927 (N_22927,N_22005,N_22423);
and U22928 (N_22928,N_22429,N_22009);
or U22929 (N_22929,N_22396,N_22077);
and U22930 (N_22930,N_22450,N_22266);
nor U22931 (N_22931,N_22356,N_22137);
or U22932 (N_22932,N_22278,N_22430);
nand U22933 (N_22933,N_22208,N_22221);
and U22934 (N_22934,N_22013,N_22441);
xnor U22935 (N_22935,N_22086,N_22424);
and U22936 (N_22936,N_22443,N_22042);
and U22937 (N_22937,N_22047,N_22013);
nand U22938 (N_22938,N_22425,N_22014);
and U22939 (N_22939,N_22315,N_22457);
nor U22940 (N_22940,N_22307,N_22476);
nor U22941 (N_22941,N_22150,N_22312);
or U22942 (N_22942,N_22106,N_22224);
xnor U22943 (N_22943,N_22183,N_22022);
xor U22944 (N_22944,N_22230,N_22359);
or U22945 (N_22945,N_22396,N_22076);
nand U22946 (N_22946,N_22460,N_22118);
or U22947 (N_22947,N_22401,N_22492);
nor U22948 (N_22948,N_22166,N_22150);
or U22949 (N_22949,N_22112,N_22276);
nand U22950 (N_22950,N_22071,N_22166);
or U22951 (N_22951,N_22374,N_22444);
nor U22952 (N_22952,N_22141,N_22155);
nor U22953 (N_22953,N_22100,N_22389);
xnor U22954 (N_22954,N_22141,N_22221);
nand U22955 (N_22955,N_22430,N_22272);
or U22956 (N_22956,N_22324,N_22258);
nor U22957 (N_22957,N_22449,N_22283);
xor U22958 (N_22958,N_22133,N_22388);
or U22959 (N_22959,N_22257,N_22440);
xnor U22960 (N_22960,N_22049,N_22021);
nand U22961 (N_22961,N_22034,N_22218);
nand U22962 (N_22962,N_22361,N_22394);
or U22963 (N_22963,N_22367,N_22345);
or U22964 (N_22964,N_22285,N_22000);
and U22965 (N_22965,N_22237,N_22219);
or U22966 (N_22966,N_22339,N_22349);
and U22967 (N_22967,N_22059,N_22438);
or U22968 (N_22968,N_22100,N_22433);
xnor U22969 (N_22969,N_22155,N_22418);
or U22970 (N_22970,N_22118,N_22155);
and U22971 (N_22971,N_22447,N_22272);
or U22972 (N_22972,N_22166,N_22291);
and U22973 (N_22973,N_22298,N_22161);
and U22974 (N_22974,N_22079,N_22423);
and U22975 (N_22975,N_22476,N_22203);
nor U22976 (N_22976,N_22407,N_22221);
nand U22977 (N_22977,N_22209,N_22379);
nor U22978 (N_22978,N_22014,N_22241);
and U22979 (N_22979,N_22131,N_22203);
or U22980 (N_22980,N_22121,N_22311);
and U22981 (N_22981,N_22019,N_22355);
and U22982 (N_22982,N_22270,N_22122);
nor U22983 (N_22983,N_22076,N_22455);
xor U22984 (N_22984,N_22400,N_22152);
and U22985 (N_22985,N_22004,N_22145);
xnor U22986 (N_22986,N_22474,N_22338);
nor U22987 (N_22987,N_22304,N_22433);
nor U22988 (N_22988,N_22348,N_22109);
nor U22989 (N_22989,N_22418,N_22013);
xor U22990 (N_22990,N_22217,N_22338);
nor U22991 (N_22991,N_22174,N_22369);
nor U22992 (N_22992,N_22062,N_22434);
xor U22993 (N_22993,N_22149,N_22044);
nand U22994 (N_22994,N_22241,N_22369);
nand U22995 (N_22995,N_22011,N_22255);
nand U22996 (N_22996,N_22317,N_22017);
and U22997 (N_22997,N_22464,N_22240);
and U22998 (N_22998,N_22187,N_22237);
xnor U22999 (N_22999,N_22330,N_22119);
nor U23000 (N_23000,N_22913,N_22888);
nand U23001 (N_23001,N_22535,N_22669);
xor U23002 (N_23002,N_22644,N_22703);
nor U23003 (N_23003,N_22557,N_22765);
nand U23004 (N_23004,N_22991,N_22802);
and U23005 (N_23005,N_22894,N_22912);
nand U23006 (N_23006,N_22590,N_22944);
or U23007 (N_23007,N_22870,N_22635);
nor U23008 (N_23008,N_22562,N_22609);
or U23009 (N_23009,N_22873,N_22769);
and U23010 (N_23010,N_22841,N_22604);
nor U23011 (N_23011,N_22868,N_22937);
xnor U23012 (N_23012,N_22835,N_22903);
and U23013 (N_23013,N_22907,N_22610);
and U23014 (N_23014,N_22757,N_22943);
nor U23015 (N_23015,N_22803,N_22794);
nand U23016 (N_23016,N_22598,N_22645);
and U23017 (N_23017,N_22720,N_22917);
nor U23018 (N_23018,N_22852,N_22756);
or U23019 (N_23019,N_22999,N_22707);
nor U23020 (N_23020,N_22682,N_22534);
xnor U23021 (N_23021,N_22694,N_22824);
or U23022 (N_23022,N_22850,N_22960);
xor U23023 (N_23023,N_22760,N_22602);
and U23024 (N_23024,N_22930,N_22838);
nor U23025 (N_23025,N_22680,N_22654);
nor U23026 (N_23026,N_22821,N_22789);
and U23027 (N_23027,N_22509,N_22513);
or U23028 (N_23028,N_22800,N_22671);
nand U23029 (N_23029,N_22528,N_22660);
and U23030 (N_23030,N_22640,N_22786);
nor U23031 (N_23031,N_22896,N_22507);
and U23032 (N_23032,N_22872,N_22901);
or U23033 (N_23033,N_22674,N_22619);
xor U23034 (N_23034,N_22808,N_22722);
nor U23035 (N_23035,N_22607,N_22844);
and U23036 (N_23036,N_22891,N_22819);
or U23037 (N_23037,N_22993,N_22996);
nor U23038 (N_23038,N_22730,N_22813);
and U23039 (N_23039,N_22822,N_22593);
nand U23040 (N_23040,N_22869,N_22963);
xnor U23041 (N_23041,N_22898,N_22701);
and U23042 (N_23042,N_22630,N_22804);
or U23043 (N_23043,N_22832,N_22867);
and U23044 (N_23044,N_22755,N_22633);
nor U23045 (N_23045,N_22935,N_22727);
and U23046 (N_23046,N_22905,N_22600);
nor U23047 (N_23047,N_22875,N_22828);
and U23048 (N_23048,N_22909,N_22743);
xor U23049 (N_23049,N_22959,N_22721);
or U23050 (N_23050,N_22564,N_22710);
or U23051 (N_23051,N_22693,N_22791);
nor U23052 (N_23052,N_22849,N_22941);
and U23053 (N_23053,N_22878,N_22667);
or U23054 (N_23054,N_22613,N_22874);
xnor U23055 (N_23055,N_22950,N_22541);
nand U23056 (N_23056,N_22723,N_22927);
or U23057 (N_23057,N_22911,N_22677);
or U23058 (N_23058,N_22620,N_22954);
nor U23059 (N_23059,N_22952,N_22639);
or U23060 (N_23060,N_22812,N_22866);
or U23061 (N_23061,N_22759,N_22882);
nor U23062 (N_23062,N_22864,N_22592);
nand U23063 (N_23063,N_22575,N_22711);
and U23064 (N_23064,N_22653,N_22746);
xnor U23065 (N_23065,N_22829,N_22725);
nor U23066 (N_23066,N_22742,N_22517);
or U23067 (N_23067,N_22706,N_22962);
or U23068 (N_23068,N_22751,N_22763);
and U23069 (N_23069,N_22596,N_22801);
nand U23070 (N_23070,N_22544,N_22670);
and U23071 (N_23071,N_22576,N_22735);
and U23072 (N_23072,N_22573,N_22987);
nor U23073 (N_23073,N_22775,N_22974);
or U23074 (N_23074,N_22508,N_22897);
xor U23075 (N_23075,N_22548,N_22732);
xor U23076 (N_23076,N_22688,N_22606);
nand U23077 (N_23077,N_22538,N_22536);
nand U23078 (N_23078,N_22923,N_22940);
and U23079 (N_23079,N_22915,N_22764);
or U23080 (N_23080,N_22846,N_22853);
nand U23081 (N_23081,N_22530,N_22861);
xor U23082 (N_23082,N_22807,N_22704);
nor U23083 (N_23083,N_22776,N_22792);
and U23084 (N_23084,N_22597,N_22785);
nand U23085 (N_23085,N_22699,N_22865);
and U23086 (N_23086,N_22744,N_22692);
xnor U23087 (N_23087,N_22766,N_22972);
nor U23088 (N_23088,N_22880,N_22724);
or U23089 (N_23089,N_22558,N_22877);
nand U23090 (N_23090,N_22885,N_22809);
or U23091 (N_23091,N_22626,N_22545);
nor U23092 (N_23092,N_22529,N_22554);
nor U23093 (N_23093,N_22563,N_22931);
nand U23094 (N_23094,N_22718,N_22936);
or U23095 (N_23095,N_22871,N_22657);
xor U23096 (N_23096,N_22556,N_22787);
or U23097 (N_23097,N_22580,N_22656);
nor U23098 (N_23098,N_22783,N_22551);
nand U23099 (N_23099,N_22729,N_22738);
nor U23100 (N_23100,N_22665,N_22924);
nor U23101 (N_23101,N_22958,N_22647);
and U23102 (N_23102,N_22599,N_22820);
nand U23103 (N_23103,N_22622,N_22797);
xnor U23104 (N_23104,N_22664,N_22964);
or U23105 (N_23105,N_22525,N_22966);
nand U23106 (N_23106,N_22697,N_22568);
nand U23107 (N_23107,N_22876,N_22956);
nor U23108 (N_23108,N_22501,N_22527);
nor U23109 (N_23109,N_22994,N_22526);
and U23110 (N_23110,N_22643,N_22740);
or U23111 (N_23111,N_22511,N_22552);
nor U23112 (N_23112,N_22675,N_22942);
or U23113 (N_23113,N_22632,N_22712);
xnor U23114 (N_23114,N_22949,N_22741);
nor U23115 (N_23115,N_22523,N_22601);
or U23116 (N_23116,N_22906,N_22805);
or U23117 (N_23117,N_22638,N_22934);
nor U23118 (N_23118,N_22773,N_22886);
and U23119 (N_23119,N_22522,N_22839);
and U23120 (N_23120,N_22651,N_22578);
xor U23121 (N_23121,N_22737,N_22843);
nor U23122 (N_23122,N_22831,N_22679);
and U23123 (N_23123,N_22666,N_22771);
nor U23124 (N_23124,N_22796,N_22565);
and U23125 (N_23125,N_22628,N_22709);
and U23126 (N_23126,N_22826,N_22790);
or U23127 (N_23127,N_22524,N_22689);
nor U23128 (N_23128,N_22520,N_22579);
xor U23129 (N_23129,N_22947,N_22559);
and U23130 (N_23130,N_22659,N_22845);
xor U23131 (N_23131,N_22577,N_22793);
and U23132 (N_23132,N_22842,N_22696);
nand U23133 (N_23133,N_22572,N_22982);
xor U23134 (N_23134,N_22505,N_22887);
and U23135 (N_23135,N_22502,N_22646);
nand U23136 (N_23136,N_22811,N_22782);
and U23137 (N_23137,N_22595,N_22662);
or U23138 (N_23138,N_22848,N_22854);
xnor U23139 (N_23139,N_22521,N_22990);
xor U23140 (N_23140,N_22895,N_22862);
xor U23141 (N_23141,N_22761,N_22516);
or U23142 (N_23142,N_22851,N_22733);
nor U23143 (N_23143,N_22946,N_22705);
nor U23144 (N_23144,N_22605,N_22540);
nand U23145 (N_23145,N_22997,N_22980);
and U23146 (N_23146,N_22570,N_22858);
and U23147 (N_23147,N_22961,N_22634);
xnor U23148 (N_23148,N_22648,N_22919);
nor U23149 (N_23149,N_22629,N_22615);
xnor U23150 (N_23150,N_22770,N_22883);
nand U23151 (N_23151,N_22717,N_22546);
nand U23152 (N_23152,N_22532,N_22929);
and U23153 (N_23153,N_22772,N_22779);
xnor U23154 (N_23154,N_22672,N_22921);
nor U23155 (N_23155,N_22621,N_22860);
and U23156 (N_23156,N_22591,N_22784);
xnor U23157 (N_23157,N_22614,N_22547);
nand U23158 (N_23158,N_22661,N_22902);
and U23159 (N_23159,N_22543,N_22938);
xnor U23160 (N_23160,N_22594,N_22992);
and U23161 (N_23161,N_22560,N_22624);
and U23162 (N_23162,N_22676,N_22856);
or U23163 (N_23163,N_22857,N_22700);
and U23164 (N_23164,N_22539,N_22778);
xor U23165 (N_23165,N_22798,N_22537);
xor U23166 (N_23166,N_22975,N_22890);
and U23167 (N_23167,N_22823,N_22714);
xor U23168 (N_23168,N_22518,N_22840);
xor U23169 (N_23169,N_22799,N_22767);
or U23170 (N_23170,N_22566,N_22762);
xor U23171 (N_23171,N_22879,N_22988);
or U23172 (N_23172,N_22588,N_22780);
and U23173 (N_23173,N_22561,N_22636);
or U23174 (N_23174,N_22981,N_22739);
and U23175 (N_23175,N_22702,N_22745);
xnor U23176 (N_23176,N_22863,N_22691);
or U23177 (N_23177,N_22571,N_22795);
xor U23178 (N_23178,N_22503,N_22989);
xor U23179 (N_23179,N_22584,N_22978);
nor U23180 (N_23180,N_22658,N_22892);
or U23181 (N_23181,N_22510,N_22920);
or U23182 (N_23182,N_22618,N_22678);
xor U23183 (N_23183,N_22726,N_22758);
and U23184 (N_23184,N_22833,N_22663);
or U23185 (N_23185,N_22569,N_22983);
or U23186 (N_23186,N_22719,N_22631);
and U23187 (N_23187,N_22922,N_22684);
nand U23188 (N_23188,N_22728,N_22567);
xor U23189 (N_23189,N_22768,N_22582);
nand U23190 (N_23190,N_22918,N_22752);
or U23191 (N_23191,N_22816,N_22847);
nand U23192 (N_23192,N_22973,N_22926);
and U23193 (N_23193,N_22627,N_22555);
or U23194 (N_23194,N_22855,N_22910);
nor U23195 (N_23195,N_22998,N_22683);
xnor U23196 (N_23196,N_22976,N_22749);
nor U23197 (N_23197,N_22617,N_22553);
nor U23198 (N_23198,N_22673,N_22550);
nand U23199 (N_23199,N_22957,N_22754);
and U23200 (N_23200,N_22668,N_22967);
xnor U23201 (N_23201,N_22986,N_22500);
nor U23202 (N_23202,N_22932,N_22916);
xnor U23203 (N_23203,N_22585,N_22933);
nor U23204 (N_23204,N_22977,N_22750);
or U23205 (N_23205,N_22514,N_22837);
nor U23206 (N_23206,N_22899,N_22985);
or U23207 (N_23207,N_22881,N_22731);
nand U23208 (N_23208,N_22806,N_22581);
xor U23209 (N_23209,N_22655,N_22748);
nand U23210 (N_23210,N_22681,N_22531);
xnor U23211 (N_23211,N_22649,N_22815);
xor U23212 (N_23212,N_22995,N_22914);
nand U23213 (N_23213,N_22951,N_22589);
or U23214 (N_23214,N_22512,N_22747);
and U23215 (N_23215,N_22587,N_22788);
xor U23216 (N_23216,N_22641,N_22818);
and U23217 (N_23217,N_22686,N_22519);
nand U23218 (N_23218,N_22965,N_22971);
nor U23219 (N_23219,N_22968,N_22612);
nor U23220 (N_23220,N_22574,N_22928);
nor U23221 (N_23221,N_22939,N_22984);
or U23222 (N_23222,N_22955,N_22970);
and U23223 (N_23223,N_22637,N_22549);
nor U23224 (N_23224,N_22893,N_22908);
and U23225 (N_23225,N_22753,N_22623);
xnor U23226 (N_23226,N_22652,N_22830);
and U23227 (N_23227,N_22781,N_22825);
nand U23228 (N_23228,N_22586,N_22611);
or U23229 (N_23229,N_22969,N_22836);
nor U23230 (N_23230,N_22827,N_22583);
and U23231 (N_23231,N_22810,N_22685);
nor U23232 (N_23232,N_22734,N_22889);
xor U23233 (N_23233,N_22814,N_22736);
or U23234 (N_23234,N_22904,N_22925);
nor U23235 (N_23235,N_22608,N_22650);
or U23236 (N_23236,N_22625,N_22945);
or U23237 (N_23237,N_22504,N_22777);
nand U23238 (N_23238,N_22533,N_22979);
xnor U23239 (N_23239,N_22515,N_22616);
nor U23240 (N_23240,N_22690,N_22884);
nand U23241 (N_23241,N_22687,N_22774);
nor U23242 (N_23242,N_22953,N_22642);
and U23243 (N_23243,N_22834,N_22817);
nor U23244 (N_23244,N_22716,N_22542);
or U23245 (N_23245,N_22713,N_22708);
or U23246 (N_23246,N_22506,N_22698);
xnor U23247 (N_23247,N_22695,N_22948);
or U23248 (N_23248,N_22603,N_22859);
xnor U23249 (N_23249,N_22715,N_22900);
nor U23250 (N_23250,N_22804,N_22863);
nor U23251 (N_23251,N_22747,N_22637);
and U23252 (N_23252,N_22721,N_22771);
and U23253 (N_23253,N_22789,N_22721);
nor U23254 (N_23254,N_22690,N_22863);
and U23255 (N_23255,N_22818,N_22596);
and U23256 (N_23256,N_22778,N_22632);
nor U23257 (N_23257,N_22721,N_22875);
or U23258 (N_23258,N_22844,N_22510);
xnor U23259 (N_23259,N_22782,N_22573);
xor U23260 (N_23260,N_22654,N_22692);
xnor U23261 (N_23261,N_22688,N_22658);
or U23262 (N_23262,N_22664,N_22877);
nor U23263 (N_23263,N_22580,N_22883);
and U23264 (N_23264,N_22833,N_22908);
or U23265 (N_23265,N_22567,N_22644);
nor U23266 (N_23266,N_22542,N_22720);
nand U23267 (N_23267,N_22680,N_22913);
xor U23268 (N_23268,N_22629,N_22892);
nor U23269 (N_23269,N_22742,N_22796);
or U23270 (N_23270,N_22687,N_22981);
and U23271 (N_23271,N_22801,N_22584);
or U23272 (N_23272,N_22867,N_22695);
or U23273 (N_23273,N_22787,N_22958);
and U23274 (N_23274,N_22683,N_22872);
nor U23275 (N_23275,N_22869,N_22591);
xor U23276 (N_23276,N_22810,N_22952);
and U23277 (N_23277,N_22758,N_22607);
and U23278 (N_23278,N_22534,N_22787);
xor U23279 (N_23279,N_22517,N_22671);
nand U23280 (N_23280,N_22615,N_22642);
xnor U23281 (N_23281,N_22604,N_22785);
or U23282 (N_23282,N_22968,N_22572);
or U23283 (N_23283,N_22933,N_22943);
or U23284 (N_23284,N_22614,N_22792);
nand U23285 (N_23285,N_22831,N_22894);
xnor U23286 (N_23286,N_22788,N_22598);
nand U23287 (N_23287,N_22637,N_22684);
nand U23288 (N_23288,N_22706,N_22984);
nand U23289 (N_23289,N_22773,N_22664);
and U23290 (N_23290,N_22776,N_22502);
or U23291 (N_23291,N_22716,N_22645);
xor U23292 (N_23292,N_22532,N_22797);
nor U23293 (N_23293,N_22773,N_22529);
nand U23294 (N_23294,N_22725,N_22797);
xor U23295 (N_23295,N_22879,N_22716);
and U23296 (N_23296,N_22696,N_22959);
or U23297 (N_23297,N_22749,N_22870);
nand U23298 (N_23298,N_22823,N_22750);
xor U23299 (N_23299,N_22960,N_22560);
and U23300 (N_23300,N_22955,N_22841);
xor U23301 (N_23301,N_22666,N_22591);
nand U23302 (N_23302,N_22701,N_22815);
or U23303 (N_23303,N_22889,N_22758);
or U23304 (N_23304,N_22657,N_22631);
nor U23305 (N_23305,N_22505,N_22674);
and U23306 (N_23306,N_22643,N_22937);
and U23307 (N_23307,N_22542,N_22951);
nor U23308 (N_23308,N_22689,N_22538);
xnor U23309 (N_23309,N_22520,N_22721);
nand U23310 (N_23310,N_22512,N_22519);
nor U23311 (N_23311,N_22762,N_22640);
nor U23312 (N_23312,N_22933,N_22716);
nor U23313 (N_23313,N_22773,N_22649);
xor U23314 (N_23314,N_22974,N_22930);
and U23315 (N_23315,N_22816,N_22824);
nand U23316 (N_23316,N_22980,N_22610);
xor U23317 (N_23317,N_22627,N_22726);
or U23318 (N_23318,N_22808,N_22669);
or U23319 (N_23319,N_22817,N_22735);
nor U23320 (N_23320,N_22655,N_22882);
nand U23321 (N_23321,N_22950,N_22981);
nand U23322 (N_23322,N_22658,N_22836);
or U23323 (N_23323,N_22508,N_22994);
nor U23324 (N_23324,N_22605,N_22890);
xnor U23325 (N_23325,N_22968,N_22549);
nor U23326 (N_23326,N_22918,N_22690);
nand U23327 (N_23327,N_22664,N_22780);
xnor U23328 (N_23328,N_22625,N_22803);
nand U23329 (N_23329,N_22684,N_22833);
or U23330 (N_23330,N_22512,N_22633);
nand U23331 (N_23331,N_22732,N_22642);
or U23332 (N_23332,N_22805,N_22758);
nand U23333 (N_23333,N_22965,N_22954);
or U23334 (N_23334,N_22559,N_22578);
nor U23335 (N_23335,N_22886,N_22870);
nand U23336 (N_23336,N_22976,N_22581);
xnor U23337 (N_23337,N_22619,N_22747);
nor U23338 (N_23338,N_22713,N_22955);
xnor U23339 (N_23339,N_22704,N_22531);
nor U23340 (N_23340,N_22967,N_22640);
nand U23341 (N_23341,N_22721,N_22957);
or U23342 (N_23342,N_22532,N_22561);
xnor U23343 (N_23343,N_22506,N_22795);
nor U23344 (N_23344,N_22803,N_22771);
nor U23345 (N_23345,N_22935,N_22717);
xor U23346 (N_23346,N_22842,N_22764);
or U23347 (N_23347,N_22635,N_22958);
or U23348 (N_23348,N_22657,N_22700);
and U23349 (N_23349,N_22641,N_22599);
xnor U23350 (N_23350,N_22718,N_22567);
xor U23351 (N_23351,N_22642,N_22684);
nand U23352 (N_23352,N_22674,N_22891);
xor U23353 (N_23353,N_22763,N_22558);
nand U23354 (N_23354,N_22585,N_22683);
xnor U23355 (N_23355,N_22542,N_22761);
or U23356 (N_23356,N_22524,N_22767);
nor U23357 (N_23357,N_22566,N_22789);
xor U23358 (N_23358,N_22683,N_22917);
xor U23359 (N_23359,N_22783,N_22817);
nor U23360 (N_23360,N_22992,N_22939);
nand U23361 (N_23361,N_22724,N_22531);
nand U23362 (N_23362,N_22854,N_22742);
xnor U23363 (N_23363,N_22542,N_22956);
xor U23364 (N_23364,N_22615,N_22611);
nor U23365 (N_23365,N_22672,N_22908);
nand U23366 (N_23366,N_22841,N_22673);
and U23367 (N_23367,N_22981,N_22799);
nand U23368 (N_23368,N_22789,N_22911);
nor U23369 (N_23369,N_22737,N_22754);
nand U23370 (N_23370,N_22568,N_22769);
and U23371 (N_23371,N_22839,N_22616);
nor U23372 (N_23372,N_22987,N_22739);
or U23373 (N_23373,N_22571,N_22629);
nor U23374 (N_23374,N_22729,N_22612);
xor U23375 (N_23375,N_22557,N_22978);
xor U23376 (N_23376,N_22739,N_22841);
and U23377 (N_23377,N_22983,N_22875);
nand U23378 (N_23378,N_22571,N_22737);
nor U23379 (N_23379,N_22809,N_22649);
nor U23380 (N_23380,N_22736,N_22657);
nand U23381 (N_23381,N_22901,N_22838);
or U23382 (N_23382,N_22744,N_22705);
or U23383 (N_23383,N_22778,N_22606);
and U23384 (N_23384,N_22865,N_22722);
xnor U23385 (N_23385,N_22626,N_22645);
nand U23386 (N_23386,N_22813,N_22704);
and U23387 (N_23387,N_22566,N_22776);
nor U23388 (N_23388,N_22685,N_22537);
or U23389 (N_23389,N_22932,N_22966);
and U23390 (N_23390,N_22833,N_22519);
xnor U23391 (N_23391,N_22829,N_22817);
xnor U23392 (N_23392,N_22804,N_22898);
xor U23393 (N_23393,N_22627,N_22958);
nand U23394 (N_23394,N_22959,N_22917);
xor U23395 (N_23395,N_22770,N_22692);
or U23396 (N_23396,N_22803,N_22802);
nand U23397 (N_23397,N_22891,N_22774);
nor U23398 (N_23398,N_22992,N_22968);
or U23399 (N_23399,N_22643,N_22511);
nand U23400 (N_23400,N_22889,N_22672);
nor U23401 (N_23401,N_22655,N_22692);
nor U23402 (N_23402,N_22912,N_22785);
nand U23403 (N_23403,N_22757,N_22716);
and U23404 (N_23404,N_22637,N_22958);
and U23405 (N_23405,N_22827,N_22804);
nor U23406 (N_23406,N_22566,N_22687);
nand U23407 (N_23407,N_22893,N_22854);
nor U23408 (N_23408,N_22505,N_22675);
nor U23409 (N_23409,N_22640,N_22695);
and U23410 (N_23410,N_22565,N_22547);
xnor U23411 (N_23411,N_22644,N_22641);
nor U23412 (N_23412,N_22798,N_22985);
xnor U23413 (N_23413,N_22956,N_22808);
xnor U23414 (N_23414,N_22747,N_22983);
or U23415 (N_23415,N_22979,N_22791);
or U23416 (N_23416,N_22552,N_22632);
nand U23417 (N_23417,N_22562,N_22584);
or U23418 (N_23418,N_22581,N_22530);
and U23419 (N_23419,N_22922,N_22977);
xnor U23420 (N_23420,N_22694,N_22919);
nor U23421 (N_23421,N_22548,N_22866);
and U23422 (N_23422,N_22640,N_22615);
or U23423 (N_23423,N_22602,N_22671);
nor U23424 (N_23424,N_22530,N_22941);
or U23425 (N_23425,N_22906,N_22821);
and U23426 (N_23426,N_22514,N_22912);
nand U23427 (N_23427,N_22772,N_22801);
xor U23428 (N_23428,N_22570,N_22767);
nor U23429 (N_23429,N_22607,N_22736);
nor U23430 (N_23430,N_22905,N_22842);
nor U23431 (N_23431,N_22601,N_22624);
and U23432 (N_23432,N_22976,N_22895);
nor U23433 (N_23433,N_22864,N_22789);
nor U23434 (N_23434,N_22857,N_22641);
and U23435 (N_23435,N_22631,N_22836);
nor U23436 (N_23436,N_22578,N_22655);
or U23437 (N_23437,N_22792,N_22827);
nor U23438 (N_23438,N_22699,N_22898);
xor U23439 (N_23439,N_22682,N_22522);
nor U23440 (N_23440,N_22957,N_22988);
or U23441 (N_23441,N_22820,N_22509);
and U23442 (N_23442,N_22846,N_22722);
or U23443 (N_23443,N_22661,N_22619);
and U23444 (N_23444,N_22666,N_22958);
xor U23445 (N_23445,N_22825,N_22735);
and U23446 (N_23446,N_22953,N_22727);
nand U23447 (N_23447,N_22793,N_22708);
nor U23448 (N_23448,N_22536,N_22856);
nand U23449 (N_23449,N_22881,N_22539);
nor U23450 (N_23450,N_22989,N_22599);
xor U23451 (N_23451,N_22814,N_22830);
or U23452 (N_23452,N_22642,N_22526);
nand U23453 (N_23453,N_22813,N_22656);
nor U23454 (N_23454,N_22633,N_22521);
and U23455 (N_23455,N_22604,N_22823);
or U23456 (N_23456,N_22657,N_22753);
nor U23457 (N_23457,N_22953,N_22901);
nor U23458 (N_23458,N_22781,N_22549);
and U23459 (N_23459,N_22748,N_22578);
nor U23460 (N_23460,N_22588,N_22911);
xor U23461 (N_23461,N_22614,N_22504);
nor U23462 (N_23462,N_22626,N_22911);
nand U23463 (N_23463,N_22606,N_22785);
nand U23464 (N_23464,N_22808,N_22515);
xnor U23465 (N_23465,N_22692,N_22536);
xor U23466 (N_23466,N_22905,N_22514);
xnor U23467 (N_23467,N_22889,N_22725);
and U23468 (N_23468,N_22541,N_22576);
nor U23469 (N_23469,N_22610,N_22804);
nor U23470 (N_23470,N_22655,N_22757);
or U23471 (N_23471,N_22905,N_22839);
or U23472 (N_23472,N_22755,N_22745);
or U23473 (N_23473,N_22560,N_22761);
and U23474 (N_23474,N_22819,N_22948);
nor U23475 (N_23475,N_22998,N_22574);
nor U23476 (N_23476,N_22882,N_22773);
nor U23477 (N_23477,N_22574,N_22668);
xnor U23478 (N_23478,N_22675,N_22716);
xor U23479 (N_23479,N_22645,N_22908);
xor U23480 (N_23480,N_22938,N_22595);
or U23481 (N_23481,N_22889,N_22575);
xor U23482 (N_23482,N_22826,N_22661);
xnor U23483 (N_23483,N_22914,N_22817);
or U23484 (N_23484,N_22936,N_22697);
and U23485 (N_23485,N_22525,N_22968);
nand U23486 (N_23486,N_22783,N_22723);
or U23487 (N_23487,N_22819,N_22566);
nand U23488 (N_23488,N_22505,N_22834);
nand U23489 (N_23489,N_22833,N_22868);
nand U23490 (N_23490,N_22550,N_22810);
and U23491 (N_23491,N_22801,N_22529);
or U23492 (N_23492,N_22519,N_22943);
xor U23493 (N_23493,N_22985,N_22550);
nor U23494 (N_23494,N_22870,N_22849);
and U23495 (N_23495,N_22914,N_22960);
and U23496 (N_23496,N_22639,N_22868);
or U23497 (N_23497,N_22532,N_22820);
nor U23498 (N_23498,N_22583,N_22767);
nand U23499 (N_23499,N_22721,N_22551);
and U23500 (N_23500,N_23375,N_23158);
xnor U23501 (N_23501,N_23123,N_23367);
or U23502 (N_23502,N_23215,N_23490);
or U23503 (N_23503,N_23454,N_23027);
nor U23504 (N_23504,N_23205,N_23114);
nand U23505 (N_23505,N_23415,N_23406);
nand U23506 (N_23506,N_23004,N_23300);
xnor U23507 (N_23507,N_23301,N_23395);
or U23508 (N_23508,N_23096,N_23348);
nor U23509 (N_23509,N_23154,N_23070);
nand U23510 (N_23510,N_23260,N_23031);
nand U23511 (N_23511,N_23001,N_23339);
nor U23512 (N_23512,N_23410,N_23332);
or U23513 (N_23513,N_23378,N_23151);
xnor U23514 (N_23514,N_23000,N_23443);
nand U23515 (N_23515,N_23069,N_23086);
nor U23516 (N_23516,N_23099,N_23178);
xnor U23517 (N_23517,N_23186,N_23376);
xor U23518 (N_23518,N_23212,N_23209);
xnor U23519 (N_23519,N_23062,N_23015);
xor U23520 (N_23520,N_23308,N_23382);
and U23521 (N_23521,N_23257,N_23373);
nand U23522 (N_23522,N_23456,N_23335);
or U23523 (N_23523,N_23316,N_23038);
and U23524 (N_23524,N_23153,N_23087);
nand U23525 (N_23525,N_23098,N_23133);
nor U23526 (N_23526,N_23168,N_23407);
nand U23527 (N_23527,N_23221,N_23197);
nor U23528 (N_23528,N_23005,N_23105);
and U23529 (N_23529,N_23017,N_23318);
or U23530 (N_23530,N_23253,N_23222);
and U23531 (N_23531,N_23306,N_23262);
or U23532 (N_23532,N_23130,N_23315);
and U23533 (N_23533,N_23052,N_23381);
xnor U23534 (N_23534,N_23055,N_23353);
xor U23535 (N_23535,N_23448,N_23419);
nand U23536 (N_23536,N_23231,N_23311);
nor U23537 (N_23537,N_23374,N_23021);
nand U23538 (N_23538,N_23463,N_23477);
xor U23539 (N_23539,N_23169,N_23446);
nor U23540 (N_23540,N_23405,N_23418);
nand U23541 (N_23541,N_23285,N_23207);
or U23542 (N_23542,N_23343,N_23246);
nor U23543 (N_23543,N_23080,N_23267);
nand U23544 (N_23544,N_23046,N_23408);
and U23545 (N_23545,N_23310,N_23440);
xor U23546 (N_23546,N_23333,N_23493);
nor U23547 (N_23547,N_23251,N_23228);
nor U23548 (N_23548,N_23423,N_23450);
xor U23549 (N_23549,N_23214,N_23165);
and U23550 (N_23550,N_23428,N_23045);
or U23551 (N_23551,N_23459,N_23152);
nand U23552 (N_23552,N_23449,N_23107);
or U23553 (N_23553,N_23307,N_23494);
xnor U23554 (N_23554,N_23377,N_23043);
and U23555 (N_23555,N_23058,N_23003);
or U23556 (N_23556,N_23040,N_23092);
nor U23557 (N_23557,N_23239,N_23095);
or U23558 (N_23558,N_23236,N_23427);
or U23559 (N_23559,N_23111,N_23386);
nand U23560 (N_23560,N_23137,N_23319);
and U23561 (N_23561,N_23030,N_23065);
or U23562 (N_23562,N_23258,N_23366);
nand U23563 (N_23563,N_23163,N_23276);
xor U23564 (N_23564,N_23391,N_23486);
xnor U23565 (N_23565,N_23256,N_23009);
nor U23566 (N_23566,N_23242,N_23094);
xor U23567 (N_23567,N_23324,N_23115);
nand U23568 (N_23568,N_23255,N_23136);
or U23569 (N_23569,N_23141,N_23287);
nor U23570 (N_23570,N_23220,N_23283);
nor U23571 (N_23571,N_23126,N_23201);
nand U23572 (N_23572,N_23400,N_23421);
xnor U23573 (N_23573,N_23061,N_23329);
and U23574 (N_23574,N_23057,N_23438);
xnor U23575 (N_23575,N_23349,N_23259);
and U23576 (N_23576,N_23396,N_23434);
or U23577 (N_23577,N_23128,N_23411);
nand U23578 (N_23578,N_23112,N_23149);
nor U23579 (N_23579,N_23199,N_23489);
nand U23580 (N_23580,N_23179,N_23340);
nand U23581 (N_23581,N_23483,N_23357);
nand U23582 (N_23582,N_23473,N_23398);
and U23583 (N_23583,N_23478,N_23206);
nor U23584 (N_23584,N_23254,N_23089);
or U23585 (N_23585,N_23488,N_23441);
and U23586 (N_23586,N_23060,N_23139);
nor U23587 (N_23587,N_23088,N_23291);
xnor U23588 (N_23588,N_23263,N_23218);
nor U23589 (N_23589,N_23379,N_23394);
nor U23590 (N_23590,N_23225,N_23485);
and U23591 (N_23591,N_23020,N_23232);
or U23592 (N_23592,N_23338,N_23024);
nand U23593 (N_23593,N_23167,N_23193);
nor U23594 (N_23594,N_23350,N_23150);
or U23595 (N_23595,N_23445,N_23413);
xnor U23596 (N_23596,N_23131,N_23326);
nor U23597 (N_23597,N_23144,N_23172);
and U23598 (N_23598,N_23482,N_23320);
and U23599 (N_23599,N_23109,N_23044);
or U23600 (N_23600,N_23387,N_23250);
nor U23601 (N_23601,N_23195,N_23426);
or U23602 (N_23602,N_23281,N_23202);
or U23603 (N_23603,N_23019,N_23497);
and U23604 (N_23604,N_23397,N_23064);
nand U23605 (N_23605,N_23277,N_23425);
nor U23606 (N_23606,N_23476,N_23286);
and U23607 (N_23607,N_23298,N_23016);
xnor U23608 (N_23608,N_23113,N_23292);
nor U23609 (N_23609,N_23295,N_23341);
nor U23610 (N_23610,N_23142,N_23304);
xor U23611 (N_23611,N_23176,N_23330);
and U23612 (N_23612,N_23275,N_23264);
nor U23613 (N_23613,N_23491,N_23191);
or U23614 (N_23614,N_23066,N_23196);
nand U23615 (N_23615,N_23082,N_23104);
nor U23616 (N_23616,N_23235,N_23203);
nor U23617 (N_23617,N_23447,N_23124);
nand U23618 (N_23618,N_23211,N_23177);
nor U23619 (N_23619,N_23480,N_23063);
and U23620 (N_23620,N_23127,N_23466);
or U23621 (N_23621,N_23472,N_23039);
and U23622 (N_23622,N_23302,N_23247);
nand U23623 (N_23623,N_23081,N_23336);
xnor U23624 (N_23624,N_23006,N_23297);
nor U23625 (N_23625,N_23143,N_23420);
xor U23626 (N_23626,N_23075,N_23498);
or U23627 (N_23627,N_23155,N_23078);
or U23628 (N_23628,N_23238,N_23355);
and U23629 (N_23629,N_23369,N_23370);
or U23630 (N_23630,N_23194,N_23180);
nor U23631 (N_23631,N_23125,N_23162);
or U23632 (N_23632,N_23029,N_23455);
or U23633 (N_23633,N_23054,N_23312);
or U23634 (N_23634,N_23189,N_23204);
xor U23635 (N_23635,N_23296,N_23083);
nand U23636 (N_23636,N_23271,N_23467);
or U23637 (N_23637,N_23299,N_23389);
nor U23638 (N_23638,N_23103,N_23412);
or U23639 (N_23639,N_23041,N_23119);
xor U23640 (N_23640,N_23346,N_23118);
or U23641 (N_23641,N_23170,N_23334);
xor U23642 (N_23642,N_23240,N_23101);
xnor U23643 (N_23643,N_23442,N_23337);
nand U23644 (N_23644,N_23331,N_23171);
and U23645 (N_23645,N_23495,N_23437);
nor U23646 (N_23646,N_23272,N_23037);
xnor U23647 (N_23647,N_23404,N_23470);
nor U23648 (N_23648,N_23079,N_23471);
nand U23649 (N_23649,N_23077,N_23223);
nor U23650 (N_23650,N_23280,N_23399);
nand U23651 (N_23651,N_23278,N_23229);
nand U23652 (N_23652,N_23116,N_23475);
and U23653 (N_23653,N_23008,N_23249);
and U23654 (N_23654,N_23159,N_23157);
xnor U23655 (N_23655,N_23460,N_23084);
nor U23656 (N_23656,N_23309,N_23452);
and U23657 (N_23657,N_23313,N_23190);
or U23658 (N_23658,N_23184,N_23388);
and U23659 (N_23659,N_23435,N_23347);
or U23660 (N_23660,N_23213,N_23091);
and U23661 (N_23661,N_23034,N_23085);
xnor U23662 (N_23662,N_23284,N_23166);
xor U23663 (N_23663,N_23457,N_23265);
or U23664 (N_23664,N_23192,N_23245);
xor U23665 (N_23665,N_23068,N_23444);
xor U23666 (N_23666,N_23072,N_23132);
nor U23667 (N_23667,N_23050,N_23289);
nor U23668 (N_23668,N_23416,N_23056);
nor U23669 (N_23669,N_23282,N_23414);
or U23670 (N_23670,N_23268,N_23492);
or U23671 (N_23671,N_23033,N_23042);
nor U23672 (N_23672,N_23013,N_23174);
xor U23673 (N_23673,N_23474,N_23362);
xor U23674 (N_23674,N_23422,N_23110);
and U23675 (N_23675,N_23059,N_23325);
nand U23676 (N_23676,N_23200,N_23499);
xor U23677 (N_23677,N_23048,N_23208);
nand U23678 (N_23678,N_23430,N_23342);
and U23679 (N_23679,N_23351,N_23022);
nor U23680 (N_23680,N_23146,N_23403);
and U23681 (N_23681,N_23007,N_23147);
xnor U23682 (N_23682,N_23481,N_23224);
nand U23683 (N_23683,N_23173,N_23090);
nand U23684 (N_23684,N_23135,N_23252);
or U23685 (N_23685,N_23164,N_23417);
or U23686 (N_23686,N_23294,N_23241);
nor U23687 (N_23687,N_23051,N_23049);
and U23688 (N_23688,N_23036,N_23469);
xor U23689 (N_23689,N_23380,N_23108);
xnor U23690 (N_23690,N_23035,N_23237);
or U23691 (N_23691,N_23279,N_23451);
xor U23692 (N_23692,N_23356,N_23361);
or U23693 (N_23693,N_23359,N_23401);
xor U23694 (N_23694,N_23244,N_23328);
nor U23695 (N_23695,N_23436,N_23288);
nor U23696 (N_23696,N_23145,N_23432);
or U23697 (N_23697,N_23219,N_23138);
xnor U23698 (N_23698,N_23439,N_23269);
or U23699 (N_23699,N_23465,N_23402);
and U23700 (N_23700,N_23243,N_23305);
xnor U23701 (N_23701,N_23161,N_23458);
xor U23702 (N_23702,N_23317,N_23479);
and U23703 (N_23703,N_23273,N_23032);
nand U23704 (N_23704,N_23183,N_23384);
nor U23705 (N_23705,N_23129,N_23274);
or U23706 (N_23706,N_23266,N_23322);
or U23707 (N_23707,N_23230,N_23372);
nand U23708 (N_23708,N_23368,N_23496);
nand U23709 (N_23709,N_23392,N_23363);
nand U23710 (N_23710,N_23217,N_23010);
and U23711 (N_23711,N_23358,N_23484);
nand U23712 (N_23712,N_23431,N_23227);
or U23713 (N_23713,N_23409,N_23453);
or U23714 (N_23714,N_23074,N_23188);
or U23715 (N_23715,N_23424,N_23140);
nor U23716 (N_23716,N_23012,N_23234);
nor U23717 (N_23717,N_23148,N_23100);
and U23718 (N_23718,N_23198,N_23023);
nand U23719 (N_23719,N_23383,N_23393);
nand U23720 (N_23720,N_23429,N_23187);
or U23721 (N_23721,N_23323,N_23216);
or U23722 (N_23722,N_23120,N_23067);
and U23723 (N_23723,N_23026,N_23134);
xor U23724 (N_23724,N_23106,N_23122);
nor U23725 (N_23725,N_23182,N_23156);
nand U23726 (N_23726,N_23160,N_23175);
and U23727 (N_23727,N_23014,N_23365);
xnor U23728 (N_23728,N_23364,N_23210);
nand U23729 (N_23729,N_23102,N_23303);
xor U23730 (N_23730,N_23018,N_23076);
nand U23731 (N_23731,N_23345,N_23028);
xnor U23732 (N_23732,N_23462,N_23433);
and U23733 (N_23733,N_23293,N_23461);
nor U23734 (N_23734,N_23314,N_23047);
nor U23735 (N_23735,N_23464,N_23093);
and U23736 (N_23736,N_23352,N_23097);
nor U23737 (N_23737,N_23321,N_23233);
nand U23738 (N_23738,N_23025,N_23327);
xnor U23739 (N_23739,N_23121,N_23248);
nand U23740 (N_23740,N_23468,N_23073);
and U23741 (N_23741,N_23117,N_23290);
or U23742 (N_23742,N_23053,N_23071);
nand U23743 (N_23743,N_23354,N_23011);
nor U23744 (N_23744,N_23181,N_23226);
and U23745 (N_23745,N_23002,N_23385);
xor U23746 (N_23746,N_23390,N_23344);
nand U23747 (N_23747,N_23270,N_23371);
or U23748 (N_23748,N_23261,N_23487);
or U23749 (N_23749,N_23185,N_23360);
nand U23750 (N_23750,N_23102,N_23259);
xnor U23751 (N_23751,N_23009,N_23476);
nor U23752 (N_23752,N_23485,N_23078);
and U23753 (N_23753,N_23244,N_23431);
or U23754 (N_23754,N_23176,N_23402);
nor U23755 (N_23755,N_23146,N_23224);
and U23756 (N_23756,N_23454,N_23009);
xor U23757 (N_23757,N_23397,N_23352);
nand U23758 (N_23758,N_23265,N_23289);
or U23759 (N_23759,N_23279,N_23251);
xnor U23760 (N_23760,N_23440,N_23174);
or U23761 (N_23761,N_23425,N_23125);
and U23762 (N_23762,N_23229,N_23047);
nor U23763 (N_23763,N_23174,N_23162);
or U23764 (N_23764,N_23378,N_23476);
nor U23765 (N_23765,N_23140,N_23302);
nor U23766 (N_23766,N_23058,N_23005);
xor U23767 (N_23767,N_23087,N_23456);
nand U23768 (N_23768,N_23230,N_23444);
or U23769 (N_23769,N_23205,N_23347);
and U23770 (N_23770,N_23263,N_23208);
nand U23771 (N_23771,N_23316,N_23489);
xnor U23772 (N_23772,N_23120,N_23373);
or U23773 (N_23773,N_23276,N_23145);
and U23774 (N_23774,N_23290,N_23372);
nand U23775 (N_23775,N_23470,N_23347);
or U23776 (N_23776,N_23438,N_23416);
nor U23777 (N_23777,N_23399,N_23111);
xnor U23778 (N_23778,N_23081,N_23400);
xnor U23779 (N_23779,N_23133,N_23011);
nand U23780 (N_23780,N_23477,N_23351);
nand U23781 (N_23781,N_23046,N_23220);
nor U23782 (N_23782,N_23067,N_23397);
nand U23783 (N_23783,N_23168,N_23325);
or U23784 (N_23784,N_23003,N_23138);
nor U23785 (N_23785,N_23482,N_23044);
nand U23786 (N_23786,N_23136,N_23014);
and U23787 (N_23787,N_23311,N_23012);
and U23788 (N_23788,N_23012,N_23293);
or U23789 (N_23789,N_23385,N_23456);
and U23790 (N_23790,N_23168,N_23060);
nand U23791 (N_23791,N_23430,N_23482);
nand U23792 (N_23792,N_23478,N_23027);
nor U23793 (N_23793,N_23080,N_23304);
xor U23794 (N_23794,N_23412,N_23439);
nor U23795 (N_23795,N_23015,N_23186);
xor U23796 (N_23796,N_23055,N_23220);
nand U23797 (N_23797,N_23375,N_23071);
nor U23798 (N_23798,N_23317,N_23382);
nor U23799 (N_23799,N_23245,N_23223);
and U23800 (N_23800,N_23471,N_23264);
nor U23801 (N_23801,N_23206,N_23378);
nor U23802 (N_23802,N_23433,N_23295);
nor U23803 (N_23803,N_23143,N_23182);
or U23804 (N_23804,N_23440,N_23230);
nand U23805 (N_23805,N_23218,N_23426);
and U23806 (N_23806,N_23456,N_23267);
or U23807 (N_23807,N_23147,N_23020);
nor U23808 (N_23808,N_23066,N_23115);
xnor U23809 (N_23809,N_23247,N_23050);
and U23810 (N_23810,N_23313,N_23263);
or U23811 (N_23811,N_23252,N_23343);
and U23812 (N_23812,N_23246,N_23271);
and U23813 (N_23813,N_23189,N_23495);
and U23814 (N_23814,N_23367,N_23192);
nor U23815 (N_23815,N_23363,N_23422);
and U23816 (N_23816,N_23185,N_23498);
nand U23817 (N_23817,N_23115,N_23351);
and U23818 (N_23818,N_23164,N_23177);
xnor U23819 (N_23819,N_23494,N_23427);
nand U23820 (N_23820,N_23130,N_23336);
nand U23821 (N_23821,N_23478,N_23432);
or U23822 (N_23822,N_23344,N_23373);
nand U23823 (N_23823,N_23071,N_23099);
and U23824 (N_23824,N_23140,N_23433);
or U23825 (N_23825,N_23200,N_23008);
nand U23826 (N_23826,N_23010,N_23454);
and U23827 (N_23827,N_23271,N_23122);
or U23828 (N_23828,N_23399,N_23231);
or U23829 (N_23829,N_23471,N_23021);
nand U23830 (N_23830,N_23012,N_23003);
xnor U23831 (N_23831,N_23246,N_23389);
and U23832 (N_23832,N_23398,N_23059);
xnor U23833 (N_23833,N_23102,N_23251);
xnor U23834 (N_23834,N_23437,N_23112);
and U23835 (N_23835,N_23300,N_23062);
and U23836 (N_23836,N_23126,N_23491);
nor U23837 (N_23837,N_23304,N_23360);
xnor U23838 (N_23838,N_23470,N_23153);
or U23839 (N_23839,N_23150,N_23363);
nor U23840 (N_23840,N_23378,N_23451);
and U23841 (N_23841,N_23407,N_23172);
and U23842 (N_23842,N_23246,N_23086);
nand U23843 (N_23843,N_23048,N_23259);
and U23844 (N_23844,N_23165,N_23429);
nor U23845 (N_23845,N_23417,N_23147);
and U23846 (N_23846,N_23472,N_23250);
or U23847 (N_23847,N_23225,N_23496);
and U23848 (N_23848,N_23182,N_23069);
nor U23849 (N_23849,N_23344,N_23430);
nand U23850 (N_23850,N_23489,N_23094);
and U23851 (N_23851,N_23114,N_23373);
xnor U23852 (N_23852,N_23399,N_23367);
xor U23853 (N_23853,N_23446,N_23227);
xnor U23854 (N_23854,N_23457,N_23087);
and U23855 (N_23855,N_23197,N_23207);
or U23856 (N_23856,N_23475,N_23292);
xor U23857 (N_23857,N_23214,N_23406);
xnor U23858 (N_23858,N_23038,N_23460);
nor U23859 (N_23859,N_23442,N_23275);
and U23860 (N_23860,N_23252,N_23140);
xnor U23861 (N_23861,N_23190,N_23098);
nand U23862 (N_23862,N_23044,N_23238);
nand U23863 (N_23863,N_23293,N_23440);
and U23864 (N_23864,N_23181,N_23008);
and U23865 (N_23865,N_23156,N_23463);
nand U23866 (N_23866,N_23491,N_23263);
nand U23867 (N_23867,N_23448,N_23055);
or U23868 (N_23868,N_23202,N_23487);
nand U23869 (N_23869,N_23156,N_23233);
nand U23870 (N_23870,N_23467,N_23190);
xor U23871 (N_23871,N_23408,N_23119);
or U23872 (N_23872,N_23363,N_23215);
nand U23873 (N_23873,N_23490,N_23462);
xor U23874 (N_23874,N_23178,N_23481);
nor U23875 (N_23875,N_23039,N_23363);
nand U23876 (N_23876,N_23453,N_23037);
and U23877 (N_23877,N_23364,N_23121);
or U23878 (N_23878,N_23159,N_23334);
nor U23879 (N_23879,N_23250,N_23188);
nand U23880 (N_23880,N_23109,N_23299);
and U23881 (N_23881,N_23435,N_23453);
xor U23882 (N_23882,N_23253,N_23039);
and U23883 (N_23883,N_23135,N_23098);
xnor U23884 (N_23884,N_23475,N_23387);
xnor U23885 (N_23885,N_23281,N_23430);
nand U23886 (N_23886,N_23445,N_23011);
or U23887 (N_23887,N_23275,N_23355);
or U23888 (N_23888,N_23041,N_23384);
nand U23889 (N_23889,N_23055,N_23293);
and U23890 (N_23890,N_23354,N_23276);
or U23891 (N_23891,N_23432,N_23440);
or U23892 (N_23892,N_23379,N_23438);
and U23893 (N_23893,N_23013,N_23407);
xnor U23894 (N_23894,N_23229,N_23150);
xor U23895 (N_23895,N_23104,N_23097);
nand U23896 (N_23896,N_23233,N_23496);
or U23897 (N_23897,N_23366,N_23264);
nor U23898 (N_23898,N_23380,N_23267);
or U23899 (N_23899,N_23206,N_23058);
or U23900 (N_23900,N_23349,N_23001);
nor U23901 (N_23901,N_23463,N_23240);
nand U23902 (N_23902,N_23296,N_23084);
or U23903 (N_23903,N_23333,N_23267);
xnor U23904 (N_23904,N_23041,N_23117);
nor U23905 (N_23905,N_23429,N_23292);
and U23906 (N_23906,N_23014,N_23225);
xor U23907 (N_23907,N_23360,N_23450);
or U23908 (N_23908,N_23232,N_23143);
nand U23909 (N_23909,N_23404,N_23198);
xor U23910 (N_23910,N_23168,N_23260);
xor U23911 (N_23911,N_23423,N_23287);
xor U23912 (N_23912,N_23124,N_23377);
nand U23913 (N_23913,N_23280,N_23492);
xnor U23914 (N_23914,N_23450,N_23169);
and U23915 (N_23915,N_23064,N_23350);
xnor U23916 (N_23916,N_23321,N_23244);
nor U23917 (N_23917,N_23199,N_23144);
xor U23918 (N_23918,N_23497,N_23371);
and U23919 (N_23919,N_23376,N_23015);
nor U23920 (N_23920,N_23385,N_23312);
nor U23921 (N_23921,N_23205,N_23169);
and U23922 (N_23922,N_23130,N_23028);
nand U23923 (N_23923,N_23284,N_23043);
and U23924 (N_23924,N_23282,N_23388);
nor U23925 (N_23925,N_23376,N_23270);
xnor U23926 (N_23926,N_23316,N_23081);
nor U23927 (N_23927,N_23089,N_23093);
nand U23928 (N_23928,N_23245,N_23202);
nand U23929 (N_23929,N_23082,N_23178);
xor U23930 (N_23930,N_23411,N_23241);
nor U23931 (N_23931,N_23276,N_23443);
nor U23932 (N_23932,N_23060,N_23084);
nand U23933 (N_23933,N_23389,N_23050);
nor U23934 (N_23934,N_23149,N_23003);
or U23935 (N_23935,N_23204,N_23137);
xnor U23936 (N_23936,N_23031,N_23004);
and U23937 (N_23937,N_23377,N_23070);
xor U23938 (N_23938,N_23151,N_23470);
xnor U23939 (N_23939,N_23309,N_23220);
or U23940 (N_23940,N_23340,N_23261);
nand U23941 (N_23941,N_23497,N_23327);
nor U23942 (N_23942,N_23103,N_23359);
xnor U23943 (N_23943,N_23277,N_23046);
nor U23944 (N_23944,N_23312,N_23381);
nor U23945 (N_23945,N_23364,N_23367);
nor U23946 (N_23946,N_23465,N_23042);
nor U23947 (N_23947,N_23377,N_23141);
xnor U23948 (N_23948,N_23426,N_23211);
and U23949 (N_23949,N_23220,N_23290);
nor U23950 (N_23950,N_23270,N_23170);
xor U23951 (N_23951,N_23118,N_23401);
and U23952 (N_23952,N_23351,N_23250);
and U23953 (N_23953,N_23383,N_23402);
nand U23954 (N_23954,N_23068,N_23481);
or U23955 (N_23955,N_23434,N_23153);
xor U23956 (N_23956,N_23173,N_23250);
xor U23957 (N_23957,N_23331,N_23114);
nand U23958 (N_23958,N_23219,N_23178);
xor U23959 (N_23959,N_23014,N_23087);
and U23960 (N_23960,N_23493,N_23426);
or U23961 (N_23961,N_23191,N_23297);
xnor U23962 (N_23962,N_23461,N_23167);
and U23963 (N_23963,N_23018,N_23357);
nand U23964 (N_23964,N_23466,N_23492);
or U23965 (N_23965,N_23107,N_23003);
xnor U23966 (N_23966,N_23301,N_23352);
or U23967 (N_23967,N_23489,N_23125);
xnor U23968 (N_23968,N_23158,N_23238);
nand U23969 (N_23969,N_23259,N_23496);
nor U23970 (N_23970,N_23248,N_23466);
nand U23971 (N_23971,N_23491,N_23314);
nor U23972 (N_23972,N_23397,N_23297);
and U23973 (N_23973,N_23447,N_23139);
nand U23974 (N_23974,N_23491,N_23120);
xor U23975 (N_23975,N_23138,N_23224);
nand U23976 (N_23976,N_23349,N_23368);
or U23977 (N_23977,N_23397,N_23051);
or U23978 (N_23978,N_23296,N_23393);
or U23979 (N_23979,N_23126,N_23046);
and U23980 (N_23980,N_23321,N_23429);
and U23981 (N_23981,N_23003,N_23447);
xor U23982 (N_23982,N_23400,N_23255);
nand U23983 (N_23983,N_23453,N_23036);
and U23984 (N_23984,N_23440,N_23099);
and U23985 (N_23985,N_23059,N_23090);
xnor U23986 (N_23986,N_23013,N_23439);
nand U23987 (N_23987,N_23380,N_23347);
nor U23988 (N_23988,N_23442,N_23313);
or U23989 (N_23989,N_23125,N_23467);
xnor U23990 (N_23990,N_23175,N_23192);
xnor U23991 (N_23991,N_23432,N_23216);
nor U23992 (N_23992,N_23286,N_23151);
or U23993 (N_23993,N_23423,N_23061);
nor U23994 (N_23994,N_23442,N_23362);
xnor U23995 (N_23995,N_23391,N_23426);
nor U23996 (N_23996,N_23156,N_23262);
xor U23997 (N_23997,N_23183,N_23348);
xor U23998 (N_23998,N_23117,N_23101);
xor U23999 (N_23999,N_23484,N_23167);
nor U24000 (N_24000,N_23995,N_23909);
nor U24001 (N_24001,N_23503,N_23877);
xnor U24002 (N_24002,N_23817,N_23810);
nand U24003 (N_24003,N_23752,N_23669);
or U24004 (N_24004,N_23580,N_23574);
xor U24005 (N_24005,N_23692,N_23647);
or U24006 (N_24006,N_23798,N_23983);
nor U24007 (N_24007,N_23620,N_23947);
nand U24008 (N_24008,N_23735,N_23860);
nand U24009 (N_24009,N_23904,N_23611);
or U24010 (N_24010,N_23788,N_23686);
and U24011 (N_24011,N_23906,N_23654);
and U24012 (N_24012,N_23957,N_23601);
or U24013 (N_24013,N_23684,N_23764);
nor U24014 (N_24014,N_23510,N_23949);
nand U24015 (N_24015,N_23790,N_23883);
xor U24016 (N_24016,N_23655,N_23586);
nor U24017 (N_24017,N_23555,N_23713);
xnor U24018 (N_24018,N_23675,N_23805);
nand U24019 (N_24019,N_23688,N_23799);
or U24020 (N_24020,N_23938,N_23832);
nor U24021 (N_24021,N_23859,N_23558);
xnor U24022 (N_24022,N_23702,N_23980);
or U24023 (N_24023,N_23635,N_23722);
nand U24024 (N_24024,N_23596,N_23993);
nor U24025 (N_24025,N_23984,N_23766);
or U24026 (N_24026,N_23756,N_23755);
xnor U24027 (N_24027,N_23780,N_23613);
nor U24028 (N_24028,N_23989,N_23927);
xor U24029 (N_24029,N_23977,N_23819);
nand U24030 (N_24030,N_23824,N_23880);
nor U24031 (N_24031,N_23533,N_23630);
or U24032 (N_24032,N_23678,N_23825);
nor U24033 (N_24033,N_23711,N_23908);
nand U24034 (N_24034,N_23800,N_23600);
or U24035 (N_24035,N_23708,N_23786);
xnor U24036 (N_24036,N_23769,N_23879);
or U24037 (N_24037,N_23840,N_23687);
nor U24038 (N_24038,N_23594,N_23531);
or U24039 (N_24039,N_23916,N_23639);
nand U24040 (N_24040,N_23597,N_23683);
and U24041 (N_24041,N_23863,N_23971);
or U24042 (N_24042,N_23645,N_23759);
or U24043 (N_24043,N_23646,N_23872);
nor U24044 (N_24044,N_23706,N_23595);
or U24045 (N_24045,N_23871,N_23821);
or U24046 (N_24046,N_23760,N_23748);
nand U24047 (N_24047,N_23593,N_23848);
or U24048 (N_24048,N_23865,N_23624);
nor U24049 (N_24049,N_23718,N_23978);
xor U24050 (N_24050,N_23553,N_23910);
nand U24051 (N_24051,N_23925,N_23576);
xor U24052 (N_24052,N_23843,N_23705);
or U24053 (N_24053,N_23912,N_23508);
nor U24054 (N_24054,N_23770,N_23968);
and U24055 (N_24055,N_23578,N_23794);
or U24056 (N_24056,N_23728,N_23552);
or U24057 (N_24057,N_23888,N_23658);
and U24058 (N_24058,N_23785,N_23823);
xnor U24059 (N_24059,N_23773,N_23515);
nand U24060 (N_24060,N_23844,N_23588);
and U24061 (N_24061,N_23621,N_23712);
or U24062 (N_24062,N_23778,N_23583);
and U24063 (N_24063,N_23549,N_23640);
xor U24064 (N_24064,N_23710,N_23884);
xor U24065 (N_24065,N_23610,N_23808);
xor U24066 (N_24066,N_23691,N_23599);
and U24067 (N_24067,N_23672,N_23699);
or U24068 (N_24068,N_23698,N_23648);
or U24069 (N_24069,N_23618,N_23606);
or U24070 (N_24070,N_23579,N_23864);
and U24071 (N_24071,N_23839,N_23592);
and U24072 (N_24072,N_23801,N_23716);
xnor U24073 (N_24073,N_23616,N_23784);
nand U24074 (N_24074,N_23598,N_23941);
xor U24075 (N_24075,N_23582,N_23791);
or U24076 (N_24076,N_23665,N_23589);
xnor U24077 (N_24077,N_23724,N_23584);
xor U24078 (N_24078,N_23822,N_23931);
or U24079 (N_24079,N_23952,N_23902);
or U24080 (N_24080,N_23763,N_23886);
xor U24081 (N_24081,N_23929,N_23750);
xnor U24082 (N_24082,N_23869,N_23890);
and U24083 (N_24083,N_23697,N_23680);
or U24084 (N_24084,N_23967,N_23591);
xor U24085 (N_24085,N_23546,N_23878);
or U24086 (N_24086,N_23913,N_23638);
nand U24087 (N_24087,N_23847,N_23537);
and U24088 (N_24088,N_23551,N_23694);
and U24089 (N_24089,N_23747,N_23700);
and U24090 (N_24090,N_23815,N_23943);
xnor U24091 (N_24091,N_23532,N_23674);
or U24092 (N_24092,N_23723,N_23516);
nand U24093 (N_24093,N_23571,N_23850);
nand U24094 (N_24094,N_23994,N_23731);
nor U24095 (N_24095,N_23568,N_23856);
or U24096 (N_24096,N_23612,N_23525);
and U24097 (N_24097,N_23973,N_23948);
nand U24098 (N_24098,N_23714,N_23746);
nand U24099 (N_24099,N_23758,N_23535);
and U24100 (N_24100,N_23975,N_23566);
nor U24101 (N_24101,N_23849,N_23804);
nor U24102 (N_24102,N_23765,N_23959);
or U24103 (N_24103,N_23667,N_23831);
nand U24104 (N_24104,N_23881,N_23545);
nand U24105 (N_24105,N_23563,N_23542);
and U24106 (N_24106,N_23561,N_23519);
and U24107 (N_24107,N_23905,N_23741);
and U24108 (N_24108,N_23795,N_23936);
nor U24109 (N_24109,N_23603,N_23816);
or U24110 (N_24110,N_23809,N_23744);
or U24111 (N_24111,N_23842,N_23939);
nand U24112 (N_24112,N_23783,N_23547);
nor U24113 (N_24113,N_23608,N_23668);
xnor U24114 (N_24114,N_23991,N_23919);
or U24115 (N_24115,N_23693,N_23853);
and U24116 (N_24116,N_23512,N_23623);
xnor U24117 (N_24117,N_23889,N_23518);
and U24118 (N_24118,N_23565,N_23836);
xor U24119 (N_24119,N_23570,N_23709);
and U24120 (N_24120,N_23845,N_23935);
nand U24121 (N_24121,N_23707,N_23605);
xor U24122 (N_24122,N_23837,N_23619);
nor U24123 (N_24123,N_23528,N_23854);
or U24124 (N_24124,N_23676,N_23664);
nand U24125 (N_24125,N_23671,N_23972);
nor U24126 (N_24126,N_23642,N_23781);
or U24127 (N_24127,N_23614,N_23685);
or U24128 (N_24128,N_23732,N_23660);
nor U24129 (N_24129,N_23999,N_23577);
or U24130 (N_24130,N_23696,N_23942);
xnor U24131 (N_24131,N_23602,N_23895);
nor U24132 (N_24132,N_23920,N_23604);
or U24133 (N_24133,N_23944,N_23524);
nor U24134 (N_24134,N_23922,N_23511);
and U24135 (N_24135,N_23803,N_23868);
or U24136 (N_24136,N_23826,N_23717);
nand U24137 (N_24137,N_23587,N_23885);
xnor U24138 (N_24138,N_23539,N_23634);
xnor U24139 (N_24139,N_23946,N_23981);
or U24140 (N_24140,N_23581,N_23522);
and U24141 (N_24141,N_23726,N_23673);
or U24142 (N_24142,N_23857,N_23911);
nand U24143 (N_24143,N_23923,N_23779);
or U24144 (N_24144,N_23988,N_23966);
nand U24145 (N_24145,N_23813,N_23768);
and U24146 (N_24146,N_23829,N_23990);
xor U24147 (N_24147,N_23926,N_23743);
xnor U24148 (N_24148,N_23641,N_23543);
nor U24149 (N_24149,N_23754,N_23969);
nor U24150 (N_24150,N_23887,N_23562);
and U24151 (N_24151,N_23734,N_23529);
nor U24152 (N_24152,N_23502,N_23745);
xor U24153 (N_24153,N_23721,N_23882);
nand U24154 (N_24154,N_23541,N_23590);
nand U24155 (N_24155,N_23695,N_23500);
nand U24156 (N_24156,N_23974,N_23715);
nand U24157 (N_24157,N_23807,N_23544);
and U24158 (N_24158,N_23749,N_23738);
nand U24159 (N_24159,N_23940,N_23792);
xnor U24160 (N_24160,N_23986,N_23559);
or U24161 (N_24161,N_23762,N_23838);
and U24162 (N_24162,N_23637,N_23960);
or U24163 (N_24163,N_23523,N_23729);
and U24164 (N_24164,N_23666,N_23793);
nand U24165 (N_24165,N_23720,N_23569);
and U24166 (N_24166,N_23841,N_23898);
nand U24167 (N_24167,N_23629,N_23656);
xor U24168 (N_24168,N_23628,N_23852);
nand U24169 (N_24169,N_23753,N_23725);
and U24170 (N_24170,N_23806,N_23733);
nor U24171 (N_24171,N_23985,N_23505);
nand U24172 (N_24172,N_23903,N_23893);
xor U24173 (N_24173,N_23509,N_23631);
or U24174 (N_24174,N_23520,N_23951);
nand U24175 (N_24175,N_23862,N_23540);
xnor U24176 (N_24176,N_23757,N_23771);
and U24177 (N_24177,N_23918,N_23915);
and U24178 (N_24178,N_23573,N_23690);
or U24179 (N_24179,N_23662,N_23987);
xnor U24180 (N_24180,N_23534,N_23742);
or U24181 (N_24181,N_23530,N_23997);
xnor U24182 (N_24182,N_23556,N_23682);
nand U24183 (N_24183,N_23653,N_23955);
nor U24184 (N_24184,N_23567,N_23504);
nand U24185 (N_24185,N_23796,N_23643);
and U24186 (N_24186,N_23736,N_23575);
or U24187 (N_24187,N_23896,N_23970);
nor U24188 (N_24188,N_23644,N_23703);
nor U24189 (N_24189,N_23661,N_23870);
nand U24190 (N_24190,N_23681,N_23617);
nand U24191 (N_24191,N_23874,N_23876);
nor U24192 (N_24192,N_23517,N_23830);
and U24193 (N_24193,N_23834,N_23789);
nor U24194 (N_24194,N_23536,N_23615);
nor U24195 (N_24195,N_23964,N_23979);
or U24196 (N_24196,N_23659,N_23514);
nor U24197 (N_24197,N_23507,N_23907);
nand U24198 (N_24198,N_23689,N_23891);
or U24199 (N_24199,N_23787,N_23636);
xnor U24200 (N_24200,N_23777,N_23740);
nor U24201 (N_24201,N_23892,N_23767);
or U24202 (N_24202,N_23867,N_23812);
nand U24203 (N_24203,N_23751,N_23921);
xnor U24204 (N_24204,N_23833,N_23992);
or U24205 (N_24205,N_23737,N_23627);
nor U24206 (N_24206,N_23739,N_23501);
xnor U24207 (N_24207,N_23866,N_23998);
nand U24208 (N_24208,N_23996,N_23704);
nor U24209 (N_24209,N_23572,N_23560);
and U24210 (N_24210,N_23632,N_23962);
and U24211 (N_24211,N_23719,N_23609);
or U24212 (N_24212,N_23633,N_23622);
nor U24213 (N_24213,N_23963,N_23932);
xnor U24214 (N_24214,N_23965,N_23900);
or U24215 (N_24215,N_23814,N_23585);
or U24216 (N_24216,N_23506,N_23820);
and U24217 (N_24217,N_23554,N_23538);
nor U24218 (N_24218,N_23548,N_23873);
or U24219 (N_24219,N_23651,N_23861);
nor U24220 (N_24220,N_23818,N_23858);
or U24221 (N_24221,N_23652,N_23982);
or U24222 (N_24222,N_23625,N_23901);
nor U24223 (N_24223,N_23782,N_23827);
or U24224 (N_24224,N_23526,N_23924);
nand U24225 (N_24225,N_23550,N_23828);
nor U24226 (N_24226,N_23958,N_23761);
nand U24227 (N_24227,N_23961,N_23701);
nor U24228 (N_24228,N_23626,N_23774);
nor U24229 (N_24229,N_23557,N_23954);
and U24230 (N_24230,N_23727,N_23670);
and U24231 (N_24231,N_23937,N_23802);
and U24232 (N_24232,N_23663,N_23657);
and U24233 (N_24233,N_23933,N_23649);
nor U24234 (N_24234,N_23730,N_23953);
nand U24235 (N_24235,N_23930,N_23797);
or U24236 (N_24236,N_23945,N_23677);
nand U24237 (N_24237,N_23679,N_23917);
nor U24238 (N_24238,N_23835,N_23897);
xor U24239 (N_24239,N_23875,N_23607);
and U24240 (N_24240,N_23650,N_23521);
nor U24241 (N_24241,N_23934,N_23772);
nor U24242 (N_24242,N_23775,N_23564);
nand U24243 (N_24243,N_23513,N_23976);
nor U24244 (N_24244,N_23855,N_23899);
nand U24245 (N_24245,N_23851,N_23776);
nand U24246 (N_24246,N_23914,N_23846);
nor U24247 (N_24247,N_23956,N_23894);
xnor U24248 (N_24248,N_23527,N_23811);
and U24249 (N_24249,N_23928,N_23950);
nor U24250 (N_24250,N_23696,N_23834);
or U24251 (N_24251,N_23962,N_23658);
or U24252 (N_24252,N_23945,N_23693);
nor U24253 (N_24253,N_23666,N_23962);
nand U24254 (N_24254,N_23907,N_23840);
xor U24255 (N_24255,N_23905,N_23938);
nand U24256 (N_24256,N_23794,N_23831);
xor U24257 (N_24257,N_23641,N_23923);
nand U24258 (N_24258,N_23669,N_23517);
nand U24259 (N_24259,N_23714,N_23871);
or U24260 (N_24260,N_23563,N_23503);
and U24261 (N_24261,N_23645,N_23998);
nor U24262 (N_24262,N_23735,N_23909);
xor U24263 (N_24263,N_23591,N_23834);
nand U24264 (N_24264,N_23982,N_23619);
and U24265 (N_24265,N_23847,N_23941);
nor U24266 (N_24266,N_23768,N_23566);
or U24267 (N_24267,N_23540,N_23743);
and U24268 (N_24268,N_23848,N_23581);
nand U24269 (N_24269,N_23573,N_23931);
or U24270 (N_24270,N_23955,N_23734);
nor U24271 (N_24271,N_23971,N_23960);
and U24272 (N_24272,N_23806,N_23711);
or U24273 (N_24273,N_23776,N_23606);
nor U24274 (N_24274,N_23694,N_23935);
or U24275 (N_24275,N_23832,N_23738);
or U24276 (N_24276,N_23545,N_23727);
and U24277 (N_24277,N_23982,N_23931);
nor U24278 (N_24278,N_23947,N_23757);
xnor U24279 (N_24279,N_23588,N_23794);
nand U24280 (N_24280,N_23659,N_23866);
nor U24281 (N_24281,N_23609,N_23805);
nor U24282 (N_24282,N_23580,N_23833);
xor U24283 (N_24283,N_23942,N_23674);
nor U24284 (N_24284,N_23871,N_23989);
xor U24285 (N_24285,N_23788,N_23600);
and U24286 (N_24286,N_23707,N_23757);
and U24287 (N_24287,N_23532,N_23944);
nor U24288 (N_24288,N_23872,N_23679);
nand U24289 (N_24289,N_23552,N_23529);
xnor U24290 (N_24290,N_23744,N_23584);
nand U24291 (N_24291,N_23809,N_23796);
nor U24292 (N_24292,N_23861,N_23742);
and U24293 (N_24293,N_23651,N_23881);
nand U24294 (N_24294,N_23579,N_23924);
or U24295 (N_24295,N_23700,N_23917);
or U24296 (N_24296,N_23514,N_23913);
and U24297 (N_24297,N_23515,N_23885);
nand U24298 (N_24298,N_23928,N_23710);
or U24299 (N_24299,N_23746,N_23782);
nand U24300 (N_24300,N_23726,N_23504);
xor U24301 (N_24301,N_23737,N_23786);
xnor U24302 (N_24302,N_23626,N_23697);
or U24303 (N_24303,N_23904,N_23845);
and U24304 (N_24304,N_23656,N_23975);
xor U24305 (N_24305,N_23840,N_23655);
xor U24306 (N_24306,N_23937,N_23695);
xnor U24307 (N_24307,N_23856,N_23563);
nand U24308 (N_24308,N_23545,N_23944);
and U24309 (N_24309,N_23881,N_23809);
and U24310 (N_24310,N_23611,N_23713);
xor U24311 (N_24311,N_23883,N_23534);
or U24312 (N_24312,N_23714,N_23692);
nor U24313 (N_24313,N_23590,N_23860);
xor U24314 (N_24314,N_23721,N_23640);
nand U24315 (N_24315,N_23995,N_23739);
or U24316 (N_24316,N_23886,N_23887);
xnor U24317 (N_24317,N_23843,N_23820);
nand U24318 (N_24318,N_23851,N_23580);
nand U24319 (N_24319,N_23734,N_23670);
nor U24320 (N_24320,N_23806,N_23877);
nor U24321 (N_24321,N_23793,N_23754);
nor U24322 (N_24322,N_23837,N_23875);
and U24323 (N_24323,N_23726,N_23794);
nand U24324 (N_24324,N_23562,N_23533);
and U24325 (N_24325,N_23878,N_23874);
nor U24326 (N_24326,N_23933,N_23813);
or U24327 (N_24327,N_23610,N_23732);
xnor U24328 (N_24328,N_23538,N_23848);
xor U24329 (N_24329,N_23639,N_23737);
and U24330 (N_24330,N_23728,N_23956);
or U24331 (N_24331,N_23812,N_23927);
or U24332 (N_24332,N_23869,N_23578);
nand U24333 (N_24333,N_23859,N_23810);
nor U24334 (N_24334,N_23615,N_23785);
or U24335 (N_24335,N_23808,N_23717);
xor U24336 (N_24336,N_23552,N_23888);
xor U24337 (N_24337,N_23679,N_23985);
and U24338 (N_24338,N_23679,N_23528);
or U24339 (N_24339,N_23775,N_23710);
or U24340 (N_24340,N_23903,N_23900);
nand U24341 (N_24341,N_23617,N_23726);
nand U24342 (N_24342,N_23926,N_23936);
xor U24343 (N_24343,N_23967,N_23801);
xnor U24344 (N_24344,N_23939,N_23674);
or U24345 (N_24345,N_23979,N_23690);
or U24346 (N_24346,N_23650,N_23762);
nor U24347 (N_24347,N_23513,N_23737);
nor U24348 (N_24348,N_23722,N_23934);
nand U24349 (N_24349,N_23738,N_23513);
nor U24350 (N_24350,N_23883,N_23824);
nand U24351 (N_24351,N_23704,N_23867);
and U24352 (N_24352,N_23901,N_23944);
nor U24353 (N_24353,N_23923,N_23857);
or U24354 (N_24354,N_23757,N_23837);
nand U24355 (N_24355,N_23529,N_23613);
nand U24356 (N_24356,N_23875,N_23533);
or U24357 (N_24357,N_23546,N_23944);
and U24358 (N_24358,N_23664,N_23583);
and U24359 (N_24359,N_23796,N_23805);
nor U24360 (N_24360,N_23659,N_23560);
and U24361 (N_24361,N_23509,N_23823);
nand U24362 (N_24362,N_23866,N_23979);
nand U24363 (N_24363,N_23535,N_23836);
and U24364 (N_24364,N_23876,N_23732);
and U24365 (N_24365,N_23584,N_23518);
nand U24366 (N_24366,N_23850,N_23623);
and U24367 (N_24367,N_23576,N_23537);
nor U24368 (N_24368,N_23904,N_23590);
nor U24369 (N_24369,N_23695,N_23534);
or U24370 (N_24370,N_23509,N_23939);
and U24371 (N_24371,N_23528,N_23664);
and U24372 (N_24372,N_23520,N_23512);
and U24373 (N_24373,N_23929,N_23538);
nor U24374 (N_24374,N_23867,N_23697);
xor U24375 (N_24375,N_23517,N_23589);
nor U24376 (N_24376,N_23778,N_23515);
nand U24377 (N_24377,N_23516,N_23948);
nor U24378 (N_24378,N_23888,N_23905);
xor U24379 (N_24379,N_23696,N_23573);
and U24380 (N_24380,N_23841,N_23735);
nand U24381 (N_24381,N_23770,N_23983);
nand U24382 (N_24382,N_23543,N_23594);
nand U24383 (N_24383,N_23560,N_23612);
nor U24384 (N_24384,N_23916,N_23682);
nor U24385 (N_24385,N_23718,N_23800);
nand U24386 (N_24386,N_23988,N_23509);
nand U24387 (N_24387,N_23810,N_23644);
xor U24388 (N_24388,N_23597,N_23507);
nand U24389 (N_24389,N_23811,N_23714);
or U24390 (N_24390,N_23621,N_23639);
xnor U24391 (N_24391,N_23813,N_23898);
nor U24392 (N_24392,N_23870,N_23873);
nor U24393 (N_24393,N_23905,N_23830);
nand U24394 (N_24394,N_23850,N_23910);
or U24395 (N_24395,N_23604,N_23917);
xnor U24396 (N_24396,N_23795,N_23695);
and U24397 (N_24397,N_23592,N_23791);
nor U24398 (N_24398,N_23618,N_23623);
nor U24399 (N_24399,N_23818,N_23942);
nor U24400 (N_24400,N_23938,N_23943);
and U24401 (N_24401,N_23603,N_23599);
nor U24402 (N_24402,N_23541,N_23964);
nor U24403 (N_24403,N_23692,N_23753);
nor U24404 (N_24404,N_23677,N_23563);
xor U24405 (N_24405,N_23786,N_23640);
nand U24406 (N_24406,N_23639,N_23715);
xnor U24407 (N_24407,N_23634,N_23788);
xor U24408 (N_24408,N_23880,N_23744);
nor U24409 (N_24409,N_23769,N_23774);
nand U24410 (N_24410,N_23629,N_23941);
xnor U24411 (N_24411,N_23687,N_23650);
nor U24412 (N_24412,N_23810,N_23572);
xnor U24413 (N_24413,N_23683,N_23788);
nor U24414 (N_24414,N_23632,N_23583);
xor U24415 (N_24415,N_23675,N_23713);
xnor U24416 (N_24416,N_23962,N_23681);
xnor U24417 (N_24417,N_23719,N_23970);
xor U24418 (N_24418,N_23695,N_23733);
xnor U24419 (N_24419,N_23836,N_23730);
xnor U24420 (N_24420,N_23937,N_23680);
or U24421 (N_24421,N_23776,N_23917);
or U24422 (N_24422,N_23663,N_23642);
nand U24423 (N_24423,N_23678,N_23672);
nor U24424 (N_24424,N_23971,N_23938);
xor U24425 (N_24425,N_23880,N_23909);
nand U24426 (N_24426,N_23849,N_23714);
xor U24427 (N_24427,N_23553,N_23607);
or U24428 (N_24428,N_23752,N_23799);
nand U24429 (N_24429,N_23787,N_23692);
nand U24430 (N_24430,N_23595,N_23840);
xor U24431 (N_24431,N_23513,N_23871);
nand U24432 (N_24432,N_23851,N_23633);
and U24433 (N_24433,N_23589,N_23960);
nor U24434 (N_24434,N_23873,N_23524);
xnor U24435 (N_24435,N_23682,N_23860);
nor U24436 (N_24436,N_23597,N_23986);
nor U24437 (N_24437,N_23871,N_23519);
nor U24438 (N_24438,N_23960,N_23638);
or U24439 (N_24439,N_23889,N_23537);
nor U24440 (N_24440,N_23787,N_23990);
xor U24441 (N_24441,N_23800,N_23590);
nor U24442 (N_24442,N_23952,N_23977);
nor U24443 (N_24443,N_23553,N_23731);
nand U24444 (N_24444,N_23678,N_23831);
or U24445 (N_24445,N_23801,N_23622);
nor U24446 (N_24446,N_23976,N_23631);
and U24447 (N_24447,N_23604,N_23824);
nand U24448 (N_24448,N_23952,N_23626);
nand U24449 (N_24449,N_23603,N_23730);
and U24450 (N_24450,N_23520,N_23946);
and U24451 (N_24451,N_23590,N_23684);
nand U24452 (N_24452,N_23679,N_23526);
or U24453 (N_24453,N_23973,N_23716);
nor U24454 (N_24454,N_23728,N_23844);
xnor U24455 (N_24455,N_23932,N_23629);
nor U24456 (N_24456,N_23836,N_23802);
nand U24457 (N_24457,N_23911,N_23614);
nor U24458 (N_24458,N_23862,N_23950);
or U24459 (N_24459,N_23805,N_23986);
nand U24460 (N_24460,N_23831,N_23872);
or U24461 (N_24461,N_23760,N_23935);
and U24462 (N_24462,N_23722,N_23819);
xor U24463 (N_24463,N_23856,N_23919);
xor U24464 (N_24464,N_23586,N_23833);
and U24465 (N_24465,N_23712,N_23592);
nand U24466 (N_24466,N_23896,N_23673);
nor U24467 (N_24467,N_23877,N_23902);
nor U24468 (N_24468,N_23840,N_23738);
nor U24469 (N_24469,N_23578,N_23693);
nor U24470 (N_24470,N_23810,N_23803);
and U24471 (N_24471,N_23762,N_23727);
xor U24472 (N_24472,N_23639,N_23624);
xor U24473 (N_24473,N_23547,N_23543);
or U24474 (N_24474,N_23655,N_23607);
nor U24475 (N_24475,N_23788,N_23991);
and U24476 (N_24476,N_23508,N_23659);
xnor U24477 (N_24477,N_23598,N_23652);
nor U24478 (N_24478,N_23993,N_23560);
xnor U24479 (N_24479,N_23835,N_23539);
or U24480 (N_24480,N_23641,N_23618);
or U24481 (N_24481,N_23856,N_23747);
and U24482 (N_24482,N_23991,N_23689);
and U24483 (N_24483,N_23966,N_23829);
and U24484 (N_24484,N_23568,N_23722);
nand U24485 (N_24485,N_23709,N_23565);
nand U24486 (N_24486,N_23697,N_23618);
nor U24487 (N_24487,N_23631,N_23597);
nor U24488 (N_24488,N_23897,N_23751);
and U24489 (N_24489,N_23638,N_23808);
nor U24490 (N_24490,N_23788,N_23720);
nor U24491 (N_24491,N_23896,N_23706);
nor U24492 (N_24492,N_23745,N_23984);
and U24493 (N_24493,N_23612,N_23944);
xor U24494 (N_24494,N_23617,N_23955);
and U24495 (N_24495,N_23581,N_23790);
xnor U24496 (N_24496,N_23733,N_23756);
nand U24497 (N_24497,N_23608,N_23524);
or U24498 (N_24498,N_23713,N_23533);
xnor U24499 (N_24499,N_23984,N_23874);
or U24500 (N_24500,N_24228,N_24105);
nand U24501 (N_24501,N_24248,N_24305);
and U24502 (N_24502,N_24344,N_24475);
nand U24503 (N_24503,N_24492,N_24004);
or U24504 (N_24504,N_24289,N_24083);
xnor U24505 (N_24505,N_24015,N_24296);
nor U24506 (N_24506,N_24064,N_24482);
or U24507 (N_24507,N_24002,N_24449);
nand U24508 (N_24508,N_24234,N_24405);
nand U24509 (N_24509,N_24307,N_24298);
xnor U24510 (N_24510,N_24139,N_24461);
xor U24511 (N_24511,N_24195,N_24028);
or U24512 (N_24512,N_24212,N_24050);
nand U24513 (N_24513,N_24210,N_24487);
and U24514 (N_24514,N_24398,N_24164);
nor U24515 (N_24515,N_24090,N_24463);
or U24516 (N_24516,N_24330,N_24432);
nor U24517 (N_24517,N_24394,N_24396);
nand U24518 (N_24518,N_24364,N_24039);
and U24519 (N_24519,N_24081,N_24240);
and U24520 (N_24520,N_24467,N_24230);
nand U24521 (N_24521,N_24437,N_24291);
or U24522 (N_24522,N_24159,N_24172);
and U24523 (N_24523,N_24478,N_24313);
xor U24524 (N_24524,N_24203,N_24054);
nor U24525 (N_24525,N_24088,N_24132);
and U24526 (N_24526,N_24480,N_24158);
and U24527 (N_24527,N_24067,N_24471);
nand U24528 (N_24528,N_24166,N_24079);
and U24529 (N_24529,N_24078,N_24495);
or U24530 (N_24530,N_24429,N_24435);
nor U24531 (N_24531,N_24100,N_24285);
nor U24532 (N_24532,N_24071,N_24318);
xor U24533 (N_24533,N_24268,N_24341);
xor U24534 (N_24534,N_24231,N_24473);
or U24535 (N_24535,N_24315,N_24140);
or U24536 (N_24536,N_24033,N_24409);
or U24537 (N_24537,N_24277,N_24392);
and U24538 (N_24538,N_24499,N_24246);
xor U24539 (N_24539,N_24274,N_24352);
nor U24540 (N_24540,N_24468,N_24456);
nand U24541 (N_24541,N_24312,N_24157);
xor U24542 (N_24542,N_24196,N_24019);
nor U24543 (N_24543,N_24148,N_24102);
nor U24544 (N_24544,N_24010,N_24243);
or U24545 (N_24545,N_24008,N_24339);
and U24546 (N_24546,N_24217,N_24378);
xnor U24547 (N_24547,N_24031,N_24184);
nor U24548 (N_24548,N_24325,N_24163);
or U24549 (N_24549,N_24051,N_24253);
xnor U24550 (N_24550,N_24138,N_24488);
nand U24551 (N_24551,N_24282,N_24410);
xor U24552 (N_24552,N_24142,N_24057);
nor U24553 (N_24553,N_24109,N_24169);
and U24554 (N_24554,N_24145,N_24370);
and U24555 (N_24555,N_24239,N_24023);
xnor U24556 (N_24556,N_24194,N_24007);
and U24557 (N_24557,N_24262,N_24290);
or U24558 (N_24558,N_24306,N_24399);
or U24559 (N_24559,N_24301,N_24238);
and U24560 (N_24560,N_24418,N_24016);
nor U24561 (N_24561,N_24348,N_24146);
and U24562 (N_24562,N_24181,N_24059);
nand U24563 (N_24563,N_24451,N_24186);
or U24564 (N_24564,N_24056,N_24123);
nand U24565 (N_24565,N_24269,N_24481);
xor U24566 (N_24566,N_24401,N_24130);
nor U24567 (N_24567,N_24419,N_24334);
nand U24568 (N_24568,N_24303,N_24252);
nor U24569 (N_24569,N_24490,N_24384);
nand U24570 (N_24570,N_24221,N_24332);
nor U24571 (N_24571,N_24074,N_24044);
nor U24572 (N_24572,N_24249,N_24182);
nor U24573 (N_24573,N_24244,N_24397);
nor U24574 (N_24574,N_24161,N_24095);
nor U24575 (N_24575,N_24052,N_24323);
or U24576 (N_24576,N_24267,N_24092);
and U24577 (N_24577,N_24207,N_24227);
or U24578 (N_24578,N_24460,N_24260);
nor U24579 (N_24579,N_24011,N_24324);
nor U24580 (N_24580,N_24255,N_24155);
and U24581 (N_24581,N_24333,N_24385);
nor U24582 (N_24582,N_24256,N_24204);
nor U24583 (N_24583,N_24417,N_24328);
xor U24584 (N_24584,N_24319,N_24125);
nand U24585 (N_24585,N_24165,N_24286);
or U24586 (N_24586,N_24359,N_24014);
or U24587 (N_24587,N_24005,N_24038);
nand U24588 (N_24588,N_24462,N_24136);
nor U24589 (N_24589,N_24469,N_24474);
xor U24590 (N_24590,N_24251,N_24126);
or U24591 (N_24591,N_24189,N_24201);
xnor U24592 (N_24592,N_24131,N_24073);
or U24593 (N_24593,N_24425,N_24171);
nor U24594 (N_24594,N_24329,N_24342);
nand U24595 (N_24595,N_24128,N_24340);
xor U24596 (N_24596,N_24192,N_24273);
or U24597 (N_24597,N_24021,N_24381);
or U24598 (N_24598,N_24193,N_24173);
nor U24599 (N_24599,N_24127,N_24094);
xor U24600 (N_24600,N_24407,N_24363);
and U24601 (N_24601,N_24302,N_24486);
or U24602 (N_24602,N_24112,N_24066);
xnor U24603 (N_24603,N_24278,N_24477);
nor U24604 (N_24604,N_24426,N_24235);
and U24605 (N_24605,N_24497,N_24436);
and U24606 (N_24606,N_24496,N_24406);
nor U24607 (N_24607,N_24421,N_24135);
xor U24608 (N_24608,N_24368,N_24408);
and U24609 (N_24609,N_24224,N_24216);
nor U24610 (N_24610,N_24391,N_24012);
xnor U24611 (N_24611,N_24080,N_24365);
nor U24612 (N_24612,N_24150,N_24393);
and U24613 (N_24613,N_24226,N_24295);
xor U24614 (N_24614,N_24063,N_24472);
or U24615 (N_24615,N_24009,N_24395);
and U24616 (N_24616,N_24452,N_24220);
nor U24617 (N_24617,N_24156,N_24085);
nor U24618 (N_24618,N_24129,N_24287);
xor U24619 (N_24619,N_24087,N_24353);
nor U24620 (N_24620,N_24089,N_24383);
nand U24621 (N_24621,N_24035,N_24279);
or U24622 (N_24622,N_24376,N_24241);
and U24623 (N_24623,N_24427,N_24206);
nand U24624 (N_24624,N_24036,N_24053);
or U24625 (N_24625,N_24441,N_24320);
nand U24626 (N_24626,N_24065,N_24388);
nor U24627 (N_24627,N_24082,N_24440);
xnor U24628 (N_24628,N_24254,N_24459);
xor U24629 (N_24629,N_24360,N_24366);
and U24630 (N_24630,N_24120,N_24357);
xor U24631 (N_24631,N_24026,N_24069);
xnor U24632 (N_24632,N_24024,N_24450);
nor U24633 (N_24633,N_24293,N_24034);
or U24634 (N_24634,N_24103,N_24420);
and U24635 (N_24635,N_24335,N_24179);
nand U24636 (N_24636,N_24162,N_24355);
nand U24637 (N_24637,N_24219,N_24374);
nand U24638 (N_24638,N_24389,N_24098);
and U24639 (N_24639,N_24237,N_24160);
nor U24640 (N_24640,N_24108,N_24032);
nor U24641 (N_24641,N_24464,N_24077);
nor U24642 (N_24642,N_24134,N_24331);
nand U24643 (N_24643,N_24466,N_24233);
or U24644 (N_24644,N_24387,N_24211);
or U24645 (N_24645,N_24042,N_24356);
xor U24646 (N_24646,N_24321,N_24223);
or U24647 (N_24647,N_24424,N_24358);
xor U24648 (N_24648,N_24245,N_24371);
nand U24649 (N_24649,N_24261,N_24119);
or U24650 (N_24650,N_24154,N_24099);
xnor U24651 (N_24651,N_24174,N_24075);
xor U24652 (N_24652,N_24362,N_24280);
nor U24653 (N_24653,N_24442,N_24045);
and U24654 (N_24654,N_24018,N_24271);
or U24655 (N_24655,N_24197,N_24068);
and U24656 (N_24656,N_24485,N_24188);
nand U24657 (N_24657,N_24354,N_24143);
or U24658 (N_24658,N_24046,N_24465);
nand U24659 (N_24659,N_24185,N_24137);
xnor U24660 (N_24660,N_24297,N_24263);
and U24661 (N_24661,N_24379,N_24281);
nand U24662 (N_24662,N_24151,N_24043);
xor U24663 (N_24663,N_24141,N_24205);
or U24664 (N_24664,N_24022,N_24236);
nor U24665 (N_24665,N_24093,N_24316);
nor U24666 (N_24666,N_24431,N_24122);
and U24667 (N_24667,N_24214,N_24483);
nor U24668 (N_24668,N_24153,N_24444);
xnor U24669 (N_24669,N_24176,N_24218);
or U24670 (N_24670,N_24152,N_24327);
nand U24671 (N_24671,N_24209,N_24190);
or U24672 (N_24672,N_24266,N_24343);
nand U24673 (N_24673,N_24454,N_24402);
nor U24674 (N_24674,N_24367,N_24175);
nor U24675 (N_24675,N_24413,N_24111);
xnor U24676 (N_24676,N_24373,N_24001);
or U24677 (N_24677,N_24041,N_24351);
nor U24678 (N_24678,N_24457,N_24013);
nand U24679 (N_24679,N_24242,N_24178);
or U24680 (N_24680,N_24422,N_24250);
nand U24681 (N_24681,N_24086,N_24037);
xor U24682 (N_24682,N_24114,N_24058);
nand U24683 (N_24683,N_24170,N_24350);
xor U24684 (N_24684,N_24117,N_24491);
nand U24685 (N_24685,N_24439,N_24149);
nand U24686 (N_24686,N_24265,N_24084);
or U24687 (N_24687,N_24489,N_24403);
nor U24688 (N_24688,N_24443,N_24115);
or U24689 (N_24689,N_24415,N_24433);
xnor U24690 (N_24690,N_24498,N_24215);
nor U24691 (N_24691,N_24453,N_24446);
and U24692 (N_24692,N_24110,N_24386);
or U24693 (N_24693,N_24264,N_24101);
nand U24694 (N_24694,N_24347,N_24258);
nor U24695 (N_24695,N_24003,N_24198);
and U24696 (N_24696,N_24275,N_24375);
nand U24697 (N_24697,N_24411,N_24310);
nor U24698 (N_24698,N_24337,N_24445);
nor U24699 (N_24699,N_24308,N_24048);
xor U24700 (N_24700,N_24076,N_24121);
nor U24701 (N_24701,N_24259,N_24199);
or U24702 (N_24702,N_24072,N_24372);
and U24703 (N_24703,N_24030,N_24412);
xor U24704 (N_24704,N_24326,N_24070);
or U24705 (N_24705,N_24232,N_24183);
and U24706 (N_24706,N_24428,N_24345);
nor U24707 (N_24707,N_24147,N_24292);
xor U24708 (N_24708,N_24493,N_24276);
xnor U24709 (N_24709,N_24494,N_24191);
nand U24710 (N_24710,N_24060,N_24314);
xor U24711 (N_24711,N_24447,N_24400);
nor U24712 (N_24712,N_24430,N_24272);
nand U24713 (N_24713,N_24369,N_24270);
nor U24714 (N_24714,N_24202,N_24017);
nor U24715 (N_24715,N_24284,N_24177);
nor U24716 (N_24716,N_24438,N_24187);
and U24717 (N_24717,N_24283,N_24257);
nand U24718 (N_24718,N_24104,N_24479);
and U24719 (N_24719,N_24288,N_24049);
nor U24720 (N_24720,N_24404,N_24096);
nand U24721 (N_24721,N_24213,N_24062);
nand U24722 (N_24722,N_24047,N_24097);
nor U24723 (N_24723,N_24377,N_24029);
nand U24724 (N_24724,N_24336,N_24091);
or U24725 (N_24725,N_24317,N_24113);
nor U24726 (N_24726,N_24448,N_24025);
nand U24727 (N_24727,N_24208,N_24020);
and U24728 (N_24728,N_24349,N_24390);
and U24729 (N_24729,N_24309,N_24470);
nand U24730 (N_24730,N_24455,N_24346);
nand U24731 (N_24731,N_24106,N_24180);
xnor U24732 (N_24732,N_24144,N_24247);
nor U24733 (N_24733,N_24000,N_24055);
xnor U24734 (N_24734,N_24300,N_24040);
nor U24735 (N_24735,N_24225,N_24423);
nand U24736 (N_24736,N_24322,N_24299);
xor U24737 (N_24737,N_24168,N_24107);
and U24738 (N_24738,N_24118,N_24133);
or U24739 (N_24739,N_24294,N_24200);
or U24740 (N_24740,N_24006,N_24458);
or U24741 (N_24741,N_24338,N_24414);
nor U24742 (N_24742,N_24484,N_24361);
xor U24743 (N_24743,N_24061,N_24167);
nor U24744 (N_24744,N_24380,N_24229);
nand U24745 (N_24745,N_24027,N_24222);
or U24746 (N_24746,N_24434,N_24304);
nor U24747 (N_24747,N_24116,N_24416);
or U24748 (N_24748,N_24311,N_24476);
and U24749 (N_24749,N_24382,N_24124);
and U24750 (N_24750,N_24458,N_24137);
xnor U24751 (N_24751,N_24190,N_24322);
and U24752 (N_24752,N_24002,N_24172);
or U24753 (N_24753,N_24273,N_24495);
nor U24754 (N_24754,N_24018,N_24319);
or U24755 (N_24755,N_24129,N_24108);
nor U24756 (N_24756,N_24289,N_24096);
xnor U24757 (N_24757,N_24495,N_24417);
or U24758 (N_24758,N_24004,N_24136);
and U24759 (N_24759,N_24151,N_24448);
nor U24760 (N_24760,N_24298,N_24233);
and U24761 (N_24761,N_24180,N_24307);
or U24762 (N_24762,N_24461,N_24155);
xnor U24763 (N_24763,N_24446,N_24020);
xor U24764 (N_24764,N_24052,N_24324);
nand U24765 (N_24765,N_24074,N_24101);
and U24766 (N_24766,N_24448,N_24313);
nand U24767 (N_24767,N_24492,N_24383);
xnor U24768 (N_24768,N_24429,N_24163);
nor U24769 (N_24769,N_24468,N_24471);
or U24770 (N_24770,N_24357,N_24176);
nor U24771 (N_24771,N_24296,N_24032);
and U24772 (N_24772,N_24386,N_24434);
nor U24773 (N_24773,N_24014,N_24189);
nand U24774 (N_24774,N_24486,N_24207);
nand U24775 (N_24775,N_24472,N_24284);
or U24776 (N_24776,N_24012,N_24218);
or U24777 (N_24777,N_24372,N_24248);
nand U24778 (N_24778,N_24197,N_24492);
xor U24779 (N_24779,N_24494,N_24038);
nor U24780 (N_24780,N_24246,N_24303);
and U24781 (N_24781,N_24152,N_24475);
or U24782 (N_24782,N_24164,N_24439);
and U24783 (N_24783,N_24391,N_24123);
nor U24784 (N_24784,N_24397,N_24366);
xnor U24785 (N_24785,N_24490,N_24460);
xor U24786 (N_24786,N_24160,N_24087);
nand U24787 (N_24787,N_24042,N_24008);
or U24788 (N_24788,N_24102,N_24271);
and U24789 (N_24789,N_24002,N_24398);
and U24790 (N_24790,N_24446,N_24320);
or U24791 (N_24791,N_24142,N_24022);
and U24792 (N_24792,N_24192,N_24356);
nor U24793 (N_24793,N_24492,N_24092);
nor U24794 (N_24794,N_24132,N_24259);
and U24795 (N_24795,N_24451,N_24132);
nand U24796 (N_24796,N_24005,N_24276);
and U24797 (N_24797,N_24383,N_24286);
or U24798 (N_24798,N_24000,N_24492);
and U24799 (N_24799,N_24413,N_24211);
xor U24800 (N_24800,N_24196,N_24322);
xor U24801 (N_24801,N_24472,N_24119);
and U24802 (N_24802,N_24343,N_24224);
or U24803 (N_24803,N_24173,N_24008);
and U24804 (N_24804,N_24444,N_24241);
nor U24805 (N_24805,N_24221,N_24339);
nand U24806 (N_24806,N_24427,N_24183);
nand U24807 (N_24807,N_24293,N_24270);
xnor U24808 (N_24808,N_24224,N_24130);
nor U24809 (N_24809,N_24402,N_24098);
nand U24810 (N_24810,N_24310,N_24020);
nor U24811 (N_24811,N_24318,N_24429);
nor U24812 (N_24812,N_24304,N_24007);
and U24813 (N_24813,N_24104,N_24184);
and U24814 (N_24814,N_24018,N_24341);
nand U24815 (N_24815,N_24050,N_24185);
xor U24816 (N_24816,N_24194,N_24336);
nand U24817 (N_24817,N_24129,N_24256);
xor U24818 (N_24818,N_24479,N_24062);
xor U24819 (N_24819,N_24214,N_24481);
and U24820 (N_24820,N_24238,N_24265);
and U24821 (N_24821,N_24282,N_24125);
nor U24822 (N_24822,N_24354,N_24125);
xnor U24823 (N_24823,N_24080,N_24428);
xor U24824 (N_24824,N_24110,N_24158);
nor U24825 (N_24825,N_24489,N_24110);
nor U24826 (N_24826,N_24491,N_24447);
xor U24827 (N_24827,N_24246,N_24088);
nor U24828 (N_24828,N_24325,N_24045);
xnor U24829 (N_24829,N_24101,N_24024);
or U24830 (N_24830,N_24016,N_24005);
or U24831 (N_24831,N_24140,N_24322);
and U24832 (N_24832,N_24389,N_24007);
or U24833 (N_24833,N_24353,N_24139);
nand U24834 (N_24834,N_24285,N_24184);
and U24835 (N_24835,N_24457,N_24292);
xor U24836 (N_24836,N_24376,N_24143);
nor U24837 (N_24837,N_24353,N_24485);
xnor U24838 (N_24838,N_24361,N_24083);
nor U24839 (N_24839,N_24291,N_24093);
or U24840 (N_24840,N_24475,N_24473);
or U24841 (N_24841,N_24190,N_24307);
and U24842 (N_24842,N_24178,N_24403);
or U24843 (N_24843,N_24231,N_24423);
or U24844 (N_24844,N_24475,N_24138);
or U24845 (N_24845,N_24334,N_24485);
nand U24846 (N_24846,N_24432,N_24418);
nor U24847 (N_24847,N_24403,N_24309);
nor U24848 (N_24848,N_24265,N_24078);
and U24849 (N_24849,N_24442,N_24195);
xnor U24850 (N_24850,N_24156,N_24041);
and U24851 (N_24851,N_24270,N_24411);
nand U24852 (N_24852,N_24300,N_24016);
and U24853 (N_24853,N_24247,N_24183);
or U24854 (N_24854,N_24387,N_24239);
nand U24855 (N_24855,N_24409,N_24170);
and U24856 (N_24856,N_24216,N_24402);
xor U24857 (N_24857,N_24320,N_24127);
or U24858 (N_24858,N_24474,N_24265);
or U24859 (N_24859,N_24029,N_24368);
nor U24860 (N_24860,N_24296,N_24024);
nand U24861 (N_24861,N_24488,N_24369);
nor U24862 (N_24862,N_24479,N_24054);
xnor U24863 (N_24863,N_24166,N_24247);
or U24864 (N_24864,N_24075,N_24235);
nor U24865 (N_24865,N_24214,N_24017);
xnor U24866 (N_24866,N_24417,N_24017);
xor U24867 (N_24867,N_24145,N_24043);
or U24868 (N_24868,N_24074,N_24411);
nor U24869 (N_24869,N_24036,N_24396);
and U24870 (N_24870,N_24321,N_24249);
or U24871 (N_24871,N_24413,N_24170);
xor U24872 (N_24872,N_24456,N_24151);
xnor U24873 (N_24873,N_24496,N_24272);
nor U24874 (N_24874,N_24439,N_24053);
and U24875 (N_24875,N_24260,N_24472);
nor U24876 (N_24876,N_24336,N_24381);
xnor U24877 (N_24877,N_24354,N_24201);
nor U24878 (N_24878,N_24421,N_24110);
xnor U24879 (N_24879,N_24193,N_24273);
nor U24880 (N_24880,N_24382,N_24113);
nor U24881 (N_24881,N_24357,N_24468);
nor U24882 (N_24882,N_24250,N_24390);
nand U24883 (N_24883,N_24197,N_24448);
xor U24884 (N_24884,N_24020,N_24491);
or U24885 (N_24885,N_24474,N_24274);
nand U24886 (N_24886,N_24003,N_24060);
and U24887 (N_24887,N_24342,N_24036);
or U24888 (N_24888,N_24015,N_24378);
nor U24889 (N_24889,N_24268,N_24360);
and U24890 (N_24890,N_24139,N_24429);
or U24891 (N_24891,N_24109,N_24228);
nand U24892 (N_24892,N_24009,N_24102);
nor U24893 (N_24893,N_24148,N_24274);
nor U24894 (N_24894,N_24488,N_24046);
nor U24895 (N_24895,N_24093,N_24438);
xnor U24896 (N_24896,N_24225,N_24030);
nor U24897 (N_24897,N_24293,N_24129);
or U24898 (N_24898,N_24211,N_24050);
and U24899 (N_24899,N_24271,N_24164);
nand U24900 (N_24900,N_24187,N_24411);
nand U24901 (N_24901,N_24467,N_24275);
or U24902 (N_24902,N_24456,N_24077);
and U24903 (N_24903,N_24468,N_24417);
nand U24904 (N_24904,N_24147,N_24057);
nor U24905 (N_24905,N_24073,N_24153);
nor U24906 (N_24906,N_24268,N_24445);
and U24907 (N_24907,N_24295,N_24401);
or U24908 (N_24908,N_24416,N_24445);
nor U24909 (N_24909,N_24118,N_24211);
nor U24910 (N_24910,N_24447,N_24374);
or U24911 (N_24911,N_24064,N_24398);
nor U24912 (N_24912,N_24038,N_24475);
nor U24913 (N_24913,N_24288,N_24261);
xor U24914 (N_24914,N_24393,N_24217);
nor U24915 (N_24915,N_24488,N_24144);
xor U24916 (N_24916,N_24055,N_24413);
and U24917 (N_24917,N_24416,N_24449);
and U24918 (N_24918,N_24250,N_24380);
nand U24919 (N_24919,N_24297,N_24087);
nand U24920 (N_24920,N_24282,N_24316);
nand U24921 (N_24921,N_24102,N_24250);
nand U24922 (N_24922,N_24146,N_24101);
and U24923 (N_24923,N_24459,N_24025);
or U24924 (N_24924,N_24337,N_24334);
nand U24925 (N_24925,N_24413,N_24258);
and U24926 (N_24926,N_24347,N_24252);
nor U24927 (N_24927,N_24474,N_24023);
xnor U24928 (N_24928,N_24386,N_24077);
nor U24929 (N_24929,N_24407,N_24265);
nand U24930 (N_24930,N_24209,N_24404);
xnor U24931 (N_24931,N_24486,N_24494);
nor U24932 (N_24932,N_24245,N_24297);
xnor U24933 (N_24933,N_24138,N_24169);
nor U24934 (N_24934,N_24071,N_24209);
xnor U24935 (N_24935,N_24474,N_24091);
or U24936 (N_24936,N_24261,N_24139);
and U24937 (N_24937,N_24450,N_24422);
nand U24938 (N_24938,N_24425,N_24119);
xnor U24939 (N_24939,N_24231,N_24042);
and U24940 (N_24940,N_24302,N_24218);
nand U24941 (N_24941,N_24424,N_24387);
nor U24942 (N_24942,N_24482,N_24240);
or U24943 (N_24943,N_24102,N_24275);
nor U24944 (N_24944,N_24295,N_24232);
nand U24945 (N_24945,N_24352,N_24289);
nor U24946 (N_24946,N_24165,N_24475);
and U24947 (N_24947,N_24175,N_24473);
or U24948 (N_24948,N_24281,N_24217);
xor U24949 (N_24949,N_24081,N_24219);
xor U24950 (N_24950,N_24443,N_24259);
and U24951 (N_24951,N_24384,N_24296);
xnor U24952 (N_24952,N_24288,N_24100);
nand U24953 (N_24953,N_24003,N_24313);
xor U24954 (N_24954,N_24143,N_24367);
nand U24955 (N_24955,N_24493,N_24042);
nand U24956 (N_24956,N_24164,N_24020);
nand U24957 (N_24957,N_24442,N_24282);
xnor U24958 (N_24958,N_24103,N_24199);
and U24959 (N_24959,N_24036,N_24318);
nand U24960 (N_24960,N_24178,N_24032);
nor U24961 (N_24961,N_24279,N_24139);
xnor U24962 (N_24962,N_24118,N_24288);
xor U24963 (N_24963,N_24462,N_24349);
xnor U24964 (N_24964,N_24361,N_24345);
nor U24965 (N_24965,N_24055,N_24067);
xnor U24966 (N_24966,N_24080,N_24391);
nand U24967 (N_24967,N_24387,N_24277);
and U24968 (N_24968,N_24349,N_24214);
xor U24969 (N_24969,N_24208,N_24474);
nand U24970 (N_24970,N_24363,N_24152);
xnor U24971 (N_24971,N_24124,N_24356);
xnor U24972 (N_24972,N_24224,N_24322);
nor U24973 (N_24973,N_24489,N_24206);
nand U24974 (N_24974,N_24024,N_24473);
and U24975 (N_24975,N_24385,N_24486);
and U24976 (N_24976,N_24138,N_24435);
nand U24977 (N_24977,N_24224,N_24247);
or U24978 (N_24978,N_24093,N_24159);
xor U24979 (N_24979,N_24490,N_24466);
nor U24980 (N_24980,N_24459,N_24084);
or U24981 (N_24981,N_24038,N_24442);
or U24982 (N_24982,N_24289,N_24052);
and U24983 (N_24983,N_24218,N_24321);
or U24984 (N_24984,N_24003,N_24462);
and U24985 (N_24985,N_24440,N_24304);
xor U24986 (N_24986,N_24041,N_24155);
nor U24987 (N_24987,N_24256,N_24429);
nand U24988 (N_24988,N_24093,N_24164);
or U24989 (N_24989,N_24145,N_24498);
or U24990 (N_24990,N_24113,N_24383);
nor U24991 (N_24991,N_24301,N_24068);
nand U24992 (N_24992,N_24097,N_24056);
nor U24993 (N_24993,N_24041,N_24396);
nor U24994 (N_24994,N_24245,N_24181);
and U24995 (N_24995,N_24468,N_24201);
or U24996 (N_24996,N_24271,N_24215);
or U24997 (N_24997,N_24309,N_24236);
xor U24998 (N_24998,N_24368,N_24171);
nor U24999 (N_24999,N_24396,N_24077);
and U25000 (N_25000,N_24751,N_24541);
nor U25001 (N_25001,N_24756,N_24822);
and U25002 (N_25002,N_24949,N_24651);
or U25003 (N_25003,N_24523,N_24576);
or U25004 (N_25004,N_24642,N_24870);
nand U25005 (N_25005,N_24806,N_24851);
and U25006 (N_25006,N_24779,N_24614);
or U25007 (N_25007,N_24901,N_24568);
or U25008 (N_25008,N_24959,N_24531);
xor U25009 (N_25009,N_24625,N_24585);
nor U25010 (N_25010,N_24655,N_24786);
or U25011 (N_25011,N_24704,N_24716);
or U25012 (N_25012,N_24667,N_24686);
and U25013 (N_25013,N_24931,N_24906);
nor U25014 (N_25014,N_24616,N_24634);
nor U25015 (N_25015,N_24998,N_24781);
xor U25016 (N_25016,N_24976,N_24729);
and U25017 (N_25017,N_24963,N_24577);
nor U25018 (N_25018,N_24617,N_24538);
nor U25019 (N_25019,N_24546,N_24774);
or U25020 (N_25020,N_24865,N_24664);
and U25021 (N_25021,N_24883,N_24515);
nor U25022 (N_25022,N_24623,N_24811);
xor U25023 (N_25023,N_24895,N_24773);
nor U25024 (N_25024,N_24837,N_24987);
and U25025 (N_25025,N_24805,N_24532);
and U25026 (N_25026,N_24711,N_24725);
or U25027 (N_25027,N_24993,N_24794);
nand U25028 (N_25028,N_24596,N_24548);
nand U25029 (N_25029,N_24525,N_24519);
and U25030 (N_25030,N_24605,N_24561);
nand U25031 (N_25031,N_24507,N_24710);
or U25032 (N_25032,N_24937,N_24898);
nor U25033 (N_25033,N_24910,N_24875);
or U25034 (N_25034,N_24545,N_24734);
nor U25035 (N_25035,N_24827,N_24738);
or U25036 (N_25036,N_24698,N_24742);
nor U25037 (N_25037,N_24814,N_24957);
nor U25038 (N_25038,N_24662,N_24755);
xor U25039 (N_25039,N_24956,N_24999);
or U25040 (N_25040,N_24619,N_24672);
or U25041 (N_25041,N_24624,N_24852);
nand U25042 (N_25042,N_24534,N_24816);
and U25043 (N_25043,N_24863,N_24592);
or U25044 (N_25044,N_24801,N_24652);
and U25045 (N_25045,N_24650,N_24726);
nor U25046 (N_25046,N_24778,N_24589);
or U25047 (N_25047,N_24992,N_24640);
nor U25048 (N_25048,N_24854,N_24914);
and U25049 (N_25049,N_24946,N_24537);
and U25050 (N_25050,N_24661,N_24749);
nor U25051 (N_25051,N_24722,N_24767);
xnor U25052 (N_25052,N_24760,N_24921);
or U25053 (N_25053,N_24974,N_24830);
xor U25054 (N_25054,N_24657,N_24842);
and U25055 (N_25055,N_24526,N_24952);
or U25056 (N_25056,N_24780,N_24673);
xor U25057 (N_25057,N_24501,N_24691);
nor U25058 (N_25058,N_24653,N_24579);
xor U25059 (N_25059,N_24697,N_24593);
or U25060 (N_25060,N_24804,N_24905);
nor U25061 (N_25061,N_24971,N_24675);
xor U25062 (N_25062,N_24934,N_24550);
xor U25063 (N_25063,N_24911,N_24853);
and U25064 (N_25064,N_24601,N_24542);
xor U25065 (N_25065,N_24636,N_24766);
or U25066 (N_25066,N_24972,N_24693);
or U25067 (N_25067,N_24688,N_24721);
or U25068 (N_25068,N_24648,N_24984);
xnor U25069 (N_25069,N_24939,N_24915);
and U25070 (N_25070,N_24897,N_24833);
and U25071 (N_25071,N_24647,N_24643);
and U25072 (N_25072,N_24754,N_24500);
nor U25073 (N_25073,N_24978,N_24995);
or U25074 (N_25074,N_24654,N_24739);
and U25075 (N_25075,N_24543,N_24613);
xnor U25076 (N_25076,N_24769,N_24689);
and U25077 (N_25077,N_24586,N_24784);
or U25078 (N_25078,N_24802,N_24789);
xor U25079 (N_25079,N_24938,N_24513);
or U25080 (N_25080,N_24890,N_24812);
nand U25081 (N_25081,N_24630,N_24904);
or U25082 (N_25082,N_24790,N_24891);
and U25083 (N_25083,N_24676,N_24819);
or U25084 (N_25084,N_24552,N_24708);
nor U25085 (N_25085,N_24682,N_24565);
nor U25086 (N_25086,N_24571,N_24700);
nand U25087 (N_25087,N_24887,N_24683);
nor U25088 (N_25088,N_24884,N_24713);
nand U25089 (N_25089,N_24813,N_24757);
and U25090 (N_25090,N_24581,N_24793);
and U25091 (N_25091,N_24847,N_24958);
nand U25092 (N_25092,N_24916,N_24936);
nand U25093 (N_25093,N_24509,N_24743);
or U25094 (N_25094,N_24553,N_24626);
nand U25095 (N_25095,N_24680,N_24600);
or U25096 (N_25096,N_24599,N_24867);
nor U25097 (N_25097,N_24718,N_24569);
nand U25098 (N_25098,N_24508,N_24953);
and U25099 (N_25099,N_24788,N_24836);
and U25100 (N_25100,N_24970,N_24889);
nand U25101 (N_25101,N_24748,N_24799);
nand U25102 (N_25102,N_24922,N_24759);
and U25103 (N_25103,N_24843,N_24530);
nor U25104 (N_25104,N_24646,N_24832);
or U25105 (N_25105,N_24763,N_24872);
nand U25106 (N_25106,N_24618,N_24660);
nor U25107 (N_25107,N_24674,N_24849);
nand U25108 (N_25108,N_24896,N_24684);
nand U25109 (N_25109,N_24735,N_24840);
nand U25110 (N_25110,N_24740,N_24797);
nor U25111 (N_25111,N_24539,N_24982);
nand U25112 (N_25112,N_24544,N_24920);
nor U25113 (N_25113,N_24528,N_24703);
or U25114 (N_25114,N_24787,N_24835);
or U25115 (N_25115,N_24514,N_24940);
nor U25116 (N_25116,N_24641,N_24608);
or U25117 (N_25117,N_24947,N_24908);
and U25118 (N_25118,N_24798,N_24583);
xnor U25119 (N_25119,N_24587,N_24732);
xnor U25120 (N_25120,N_24909,N_24925);
xnor U25121 (N_25121,N_24570,N_24838);
nor U25122 (N_25122,N_24558,N_24930);
nor U25123 (N_25123,N_24723,N_24727);
xnor U25124 (N_25124,N_24750,N_24566);
or U25125 (N_25125,N_24628,N_24745);
xnor U25126 (N_25126,N_24562,N_24876);
nor U25127 (N_25127,N_24817,N_24772);
or U25128 (N_25128,N_24609,N_24633);
and U25129 (N_25129,N_24841,N_24997);
nor U25130 (N_25130,N_24955,N_24503);
nand U25131 (N_25131,N_24681,N_24629);
and U25132 (N_25132,N_24965,N_24604);
and U25133 (N_25133,N_24556,N_24728);
nor U25134 (N_25134,N_24928,N_24969);
nor U25135 (N_25135,N_24768,N_24828);
nor U25136 (N_25136,N_24582,N_24714);
nor U25137 (N_25137,N_24900,N_24632);
and U25138 (N_25138,N_24517,N_24815);
nand U25139 (N_25139,N_24961,N_24848);
or U25140 (N_25140,N_24879,N_24511);
xor U25141 (N_25141,N_24856,N_24635);
nor U25142 (N_25142,N_24518,N_24512);
or U25143 (N_25143,N_24510,N_24927);
xor U25144 (N_25144,N_24803,N_24724);
xor U25145 (N_25145,N_24549,N_24719);
nand U25146 (N_25146,N_24758,N_24973);
xnor U25147 (N_25147,N_24873,N_24603);
and U25148 (N_25148,N_24687,N_24899);
and U25149 (N_25149,N_24504,N_24824);
nor U25150 (N_25150,N_24671,N_24575);
nand U25151 (N_25151,N_24845,N_24860);
nand U25152 (N_25152,N_24639,N_24744);
xor U25153 (N_25153,N_24945,N_24560);
xor U25154 (N_25154,N_24871,N_24764);
nand U25155 (N_25155,N_24747,N_24610);
nor U25156 (N_25156,N_24717,N_24882);
xnor U25157 (N_25157,N_24888,N_24730);
or U25158 (N_25158,N_24800,N_24831);
or U25159 (N_25159,N_24598,N_24918);
xnor U25160 (N_25160,N_24886,N_24771);
nor U25161 (N_25161,N_24715,N_24935);
and U25162 (N_25162,N_24706,N_24690);
or U25163 (N_25163,N_24559,N_24712);
nor U25164 (N_25164,N_24810,N_24645);
xor U25165 (N_25165,N_24658,N_24980);
and U25166 (N_25166,N_24590,N_24669);
and U25167 (N_25167,N_24555,N_24505);
and U25168 (N_25168,N_24588,N_24554);
xor U25169 (N_25169,N_24663,N_24753);
or U25170 (N_25170,N_24962,N_24996);
and U25171 (N_25171,N_24795,N_24536);
and U25172 (N_25172,N_24701,N_24903);
xor U25173 (N_25173,N_24994,N_24951);
and U25174 (N_25174,N_24649,N_24933);
nor U25175 (N_25175,N_24866,N_24825);
xnor U25176 (N_25176,N_24943,N_24572);
nand U25177 (N_25177,N_24820,N_24988);
or U25178 (N_25178,N_24869,N_24622);
or U25179 (N_25179,N_24902,N_24941);
xnor U25180 (N_25180,N_24948,N_24907);
nor U25181 (N_25181,N_24737,N_24981);
nor U25182 (N_25182,N_24846,N_24637);
nand U25183 (N_25183,N_24893,N_24777);
or U25184 (N_25184,N_24573,N_24964);
nand U25185 (N_25185,N_24631,N_24540);
nor U25186 (N_25186,N_24783,N_24868);
or U25187 (N_25187,N_24989,N_24923);
or U25188 (N_25188,N_24597,N_24591);
nand U25189 (N_25189,N_24808,N_24775);
and U25190 (N_25190,N_24944,N_24638);
nand U25191 (N_25191,N_24595,N_24954);
nand U25192 (N_25192,N_24821,N_24913);
nor U25193 (N_25193,N_24557,N_24551);
nand U25194 (N_25194,N_24564,N_24521);
and U25195 (N_25195,N_24516,N_24733);
nor U25196 (N_25196,N_24611,N_24834);
or U25197 (N_25197,N_24761,N_24796);
nor U25198 (N_25198,N_24968,N_24859);
nor U25199 (N_25199,N_24983,N_24917);
and U25200 (N_25200,N_24791,N_24929);
or U25201 (N_25201,N_24823,N_24584);
and U25202 (N_25202,N_24885,N_24694);
nor U25203 (N_25203,N_24894,N_24807);
or U25204 (N_25204,N_24874,N_24977);
or U25205 (N_25205,N_24696,N_24967);
nand U25206 (N_25206,N_24979,N_24547);
or U25207 (N_25207,N_24892,N_24644);
nor U25208 (N_25208,N_24861,N_24620);
nand U25209 (N_25209,N_24991,N_24785);
nand U25210 (N_25210,N_24881,N_24912);
and U25211 (N_25211,N_24966,N_24855);
xor U25212 (N_25212,N_24563,N_24776);
xnor U25213 (N_25213,N_24685,N_24522);
nor U25214 (N_25214,N_24878,N_24919);
nand U25215 (N_25215,N_24839,N_24844);
and U25216 (N_25216,N_24765,N_24782);
nor U25217 (N_25217,N_24524,N_24659);
xnor U25218 (N_25218,N_24741,N_24762);
xor U25219 (N_25219,N_24520,N_24770);
and U25220 (N_25220,N_24699,N_24877);
nor U25221 (N_25221,N_24668,N_24677);
xnor U25222 (N_25222,N_24612,N_24932);
and U25223 (N_25223,N_24506,N_24679);
and U25224 (N_25224,N_24527,N_24924);
nand U25225 (N_25225,N_24666,N_24567);
xnor U25226 (N_25226,N_24746,N_24578);
or U25227 (N_25227,N_24720,N_24792);
and U25228 (N_25228,N_24692,N_24574);
or U25229 (N_25229,N_24857,N_24880);
nand U25230 (N_25230,N_24705,N_24594);
and U25231 (N_25231,N_24709,N_24862);
nand U25232 (N_25232,N_24665,N_24809);
or U25233 (N_25233,N_24580,N_24985);
or U25234 (N_25234,N_24926,N_24975);
xor U25235 (N_25235,N_24533,N_24990);
nand U25236 (N_25236,N_24752,N_24670);
and U25237 (N_25237,N_24826,N_24678);
and U25238 (N_25238,N_24621,N_24529);
nor U25239 (N_25239,N_24850,N_24607);
and U25240 (N_25240,N_24864,N_24942);
or U25241 (N_25241,N_24858,N_24736);
or U25242 (N_25242,N_24950,N_24615);
xor U25243 (N_25243,N_24818,N_24960);
xor U25244 (N_25244,N_24986,N_24602);
xor U25245 (N_25245,N_24627,N_24829);
xor U25246 (N_25246,N_24731,N_24656);
or U25247 (N_25247,N_24606,N_24695);
and U25248 (N_25248,N_24702,N_24502);
or U25249 (N_25249,N_24707,N_24535);
nor U25250 (N_25250,N_24553,N_24746);
nand U25251 (N_25251,N_24714,N_24583);
nor U25252 (N_25252,N_24908,N_24918);
and U25253 (N_25253,N_24640,N_24514);
nor U25254 (N_25254,N_24713,N_24614);
and U25255 (N_25255,N_24957,N_24625);
or U25256 (N_25256,N_24841,N_24594);
or U25257 (N_25257,N_24586,N_24622);
nor U25258 (N_25258,N_24501,N_24642);
nand U25259 (N_25259,N_24614,N_24564);
xnor U25260 (N_25260,N_24726,N_24751);
or U25261 (N_25261,N_24688,N_24759);
nor U25262 (N_25262,N_24615,N_24894);
nor U25263 (N_25263,N_24801,N_24765);
or U25264 (N_25264,N_24983,N_24594);
nor U25265 (N_25265,N_24558,N_24536);
nand U25266 (N_25266,N_24999,N_24893);
or U25267 (N_25267,N_24910,N_24644);
xnor U25268 (N_25268,N_24965,N_24807);
xor U25269 (N_25269,N_24738,N_24704);
nand U25270 (N_25270,N_24887,N_24597);
or U25271 (N_25271,N_24854,N_24563);
nor U25272 (N_25272,N_24561,N_24607);
nor U25273 (N_25273,N_24555,N_24717);
or U25274 (N_25274,N_24950,N_24769);
and U25275 (N_25275,N_24592,N_24921);
nor U25276 (N_25276,N_24929,N_24649);
nand U25277 (N_25277,N_24535,N_24710);
and U25278 (N_25278,N_24930,N_24695);
nand U25279 (N_25279,N_24817,N_24653);
nor U25280 (N_25280,N_24747,N_24964);
or U25281 (N_25281,N_24719,N_24792);
nand U25282 (N_25282,N_24530,N_24734);
nor U25283 (N_25283,N_24970,N_24557);
nor U25284 (N_25284,N_24651,N_24761);
or U25285 (N_25285,N_24627,N_24571);
and U25286 (N_25286,N_24571,N_24919);
xnor U25287 (N_25287,N_24785,N_24865);
and U25288 (N_25288,N_24562,N_24507);
nor U25289 (N_25289,N_24838,N_24692);
nor U25290 (N_25290,N_24555,N_24677);
or U25291 (N_25291,N_24692,N_24889);
or U25292 (N_25292,N_24767,N_24616);
or U25293 (N_25293,N_24609,N_24900);
nor U25294 (N_25294,N_24756,N_24786);
or U25295 (N_25295,N_24715,N_24634);
or U25296 (N_25296,N_24683,N_24819);
and U25297 (N_25297,N_24846,N_24766);
or U25298 (N_25298,N_24851,N_24840);
nand U25299 (N_25299,N_24534,N_24586);
and U25300 (N_25300,N_24831,N_24676);
xnor U25301 (N_25301,N_24686,N_24810);
nor U25302 (N_25302,N_24830,N_24958);
nor U25303 (N_25303,N_24918,N_24987);
xnor U25304 (N_25304,N_24650,N_24631);
xor U25305 (N_25305,N_24693,N_24602);
nand U25306 (N_25306,N_24669,N_24605);
and U25307 (N_25307,N_24894,N_24822);
and U25308 (N_25308,N_24667,N_24543);
or U25309 (N_25309,N_24737,N_24841);
and U25310 (N_25310,N_24542,N_24586);
or U25311 (N_25311,N_24859,N_24738);
or U25312 (N_25312,N_24649,N_24625);
nor U25313 (N_25313,N_24527,N_24659);
nor U25314 (N_25314,N_24888,N_24794);
nand U25315 (N_25315,N_24904,N_24697);
and U25316 (N_25316,N_24598,N_24652);
nand U25317 (N_25317,N_24728,N_24983);
nand U25318 (N_25318,N_24783,N_24654);
xnor U25319 (N_25319,N_24788,N_24851);
xnor U25320 (N_25320,N_24918,N_24703);
xnor U25321 (N_25321,N_24964,N_24976);
or U25322 (N_25322,N_24710,N_24929);
nand U25323 (N_25323,N_24839,N_24529);
xor U25324 (N_25324,N_24837,N_24845);
or U25325 (N_25325,N_24735,N_24868);
or U25326 (N_25326,N_24650,N_24565);
xnor U25327 (N_25327,N_24721,N_24866);
xnor U25328 (N_25328,N_24644,N_24890);
and U25329 (N_25329,N_24769,N_24628);
xnor U25330 (N_25330,N_24564,N_24810);
or U25331 (N_25331,N_24569,N_24698);
nand U25332 (N_25332,N_24530,N_24868);
nand U25333 (N_25333,N_24932,N_24789);
xor U25334 (N_25334,N_24816,N_24642);
xnor U25335 (N_25335,N_24788,N_24890);
or U25336 (N_25336,N_24798,N_24546);
nand U25337 (N_25337,N_24919,N_24682);
or U25338 (N_25338,N_24925,N_24876);
xnor U25339 (N_25339,N_24876,N_24773);
xor U25340 (N_25340,N_24810,N_24594);
nand U25341 (N_25341,N_24620,N_24923);
nor U25342 (N_25342,N_24857,N_24697);
and U25343 (N_25343,N_24987,N_24637);
nor U25344 (N_25344,N_24723,N_24775);
nand U25345 (N_25345,N_24704,N_24929);
nor U25346 (N_25346,N_24890,N_24957);
xnor U25347 (N_25347,N_24706,N_24802);
xor U25348 (N_25348,N_24715,N_24651);
xnor U25349 (N_25349,N_24691,N_24564);
and U25350 (N_25350,N_24710,N_24771);
xnor U25351 (N_25351,N_24951,N_24892);
or U25352 (N_25352,N_24537,N_24846);
or U25353 (N_25353,N_24679,N_24890);
xnor U25354 (N_25354,N_24825,N_24787);
nand U25355 (N_25355,N_24888,N_24599);
or U25356 (N_25356,N_24998,N_24894);
nor U25357 (N_25357,N_24603,N_24634);
nor U25358 (N_25358,N_24552,N_24612);
nand U25359 (N_25359,N_24512,N_24819);
xor U25360 (N_25360,N_24698,N_24858);
nand U25361 (N_25361,N_24519,N_24537);
or U25362 (N_25362,N_24777,N_24852);
nor U25363 (N_25363,N_24760,N_24916);
xor U25364 (N_25364,N_24535,N_24681);
xnor U25365 (N_25365,N_24744,N_24812);
and U25366 (N_25366,N_24732,N_24750);
and U25367 (N_25367,N_24842,N_24748);
xnor U25368 (N_25368,N_24817,N_24503);
xnor U25369 (N_25369,N_24897,N_24755);
nand U25370 (N_25370,N_24546,N_24840);
nor U25371 (N_25371,N_24688,N_24587);
xnor U25372 (N_25372,N_24965,N_24693);
nor U25373 (N_25373,N_24750,N_24516);
nor U25374 (N_25374,N_24512,N_24956);
xor U25375 (N_25375,N_24867,N_24712);
or U25376 (N_25376,N_24673,N_24778);
nand U25377 (N_25377,N_24896,N_24657);
and U25378 (N_25378,N_24645,N_24628);
nor U25379 (N_25379,N_24694,N_24904);
nand U25380 (N_25380,N_24959,N_24647);
and U25381 (N_25381,N_24631,N_24576);
and U25382 (N_25382,N_24502,N_24983);
nor U25383 (N_25383,N_24851,N_24855);
or U25384 (N_25384,N_24766,N_24790);
nor U25385 (N_25385,N_24635,N_24983);
and U25386 (N_25386,N_24724,N_24552);
nand U25387 (N_25387,N_24909,N_24783);
nor U25388 (N_25388,N_24617,N_24705);
xor U25389 (N_25389,N_24890,N_24684);
nand U25390 (N_25390,N_24944,N_24879);
nor U25391 (N_25391,N_24684,N_24662);
or U25392 (N_25392,N_24898,N_24669);
nand U25393 (N_25393,N_24644,N_24896);
or U25394 (N_25394,N_24710,N_24635);
and U25395 (N_25395,N_24723,N_24635);
and U25396 (N_25396,N_24611,N_24795);
nand U25397 (N_25397,N_24878,N_24511);
nor U25398 (N_25398,N_24602,N_24847);
and U25399 (N_25399,N_24817,N_24802);
nor U25400 (N_25400,N_24902,N_24759);
nor U25401 (N_25401,N_24553,N_24532);
or U25402 (N_25402,N_24829,N_24915);
nand U25403 (N_25403,N_24614,N_24972);
and U25404 (N_25404,N_24864,N_24700);
nand U25405 (N_25405,N_24630,N_24664);
and U25406 (N_25406,N_24604,N_24761);
nor U25407 (N_25407,N_24626,N_24530);
nor U25408 (N_25408,N_24872,N_24613);
or U25409 (N_25409,N_24552,N_24881);
xor U25410 (N_25410,N_24601,N_24639);
nand U25411 (N_25411,N_24518,N_24966);
xor U25412 (N_25412,N_24587,N_24677);
xor U25413 (N_25413,N_24532,N_24576);
or U25414 (N_25414,N_24577,N_24925);
nor U25415 (N_25415,N_24828,N_24522);
or U25416 (N_25416,N_24664,N_24851);
nor U25417 (N_25417,N_24716,N_24804);
or U25418 (N_25418,N_24756,N_24632);
xor U25419 (N_25419,N_24941,N_24912);
xor U25420 (N_25420,N_24650,N_24632);
and U25421 (N_25421,N_24677,N_24605);
xor U25422 (N_25422,N_24965,N_24930);
and U25423 (N_25423,N_24770,N_24909);
nor U25424 (N_25424,N_24696,N_24847);
and U25425 (N_25425,N_24706,N_24785);
and U25426 (N_25426,N_24670,N_24896);
or U25427 (N_25427,N_24762,N_24617);
and U25428 (N_25428,N_24514,N_24574);
or U25429 (N_25429,N_24579,N_24887);
and U25430 (N_25430,N_24770,N_24808);
xnor U25431 (N_25431,N_24859,N_24964);
and U25432 (N_25432,N_24979,N_24544);
and U25433 (N_25433,N_24654,N_24584);
xnor U25434 (N_25434,N_24843,N_24998);
nor U25435 (N_25435,N_24665,N_24667);
xnor U25436 (N_25436,N_24932,N_24605);
or U25437 (N_25437,N_24536,N_24697);
nor U25438 (N_25438,N_24764,N_24687);
xor U25439 (N_25439,N_24711,N_24656);
nand U25440 (N_25440,N_24794,N_24795);
and U25441 (N_25441,N_24927,N_24638);
or U25442 (N_25442,N_24544,N_24722);
xor U25443 (N_25443,N_24695,N_24814);
nor U25444 (N_25444,N_24976,N_24709);
xor U25445 (N_25445,N_24697,N_24873);
and U25446 (N_25446,N_24516,N_24749);
and U25447 (N_25447,N_24820,N_24913);
nand U25448 (N_25448,N_24843,N_24720);
nor U25449 (N_25449,N_24825,N_24586);
nor U25450 (N_25450,N_24977,N_24750);
and U25451 (N_25451,N_24700,N_24634);
xnor U25452 (N_25452,N_24981,N_24524);
nand U25453 (N_25453,N_24908,N_24624);
nor U25454 (N_25454,N_24980,N_24809);
xnor U25455 (N_25455,N_24912,N_24783);
nand U25456 (N_25456,N_24802,N_24788);
and U25457 (N_25457,N_24855,N_24802);
nand U25458 (N_25458,N_24507,N_24663);
or U25459 (N_25459,N_24731,N_24941);
or U25460 (N_25460,N_24922,N_24757);
and U25461 (N_25461,N_24699,N_24513);
and U25462 (N_25462,N_24584,N_24577);
nor U25463 (N_25463,N_24605,N_24795);
or U25464 (N_25464,N_24706,N_24618);
nand U25465 (N_25465,N_24738,N_24766);
nand U25466 (N_25466,N_24679,N_24955);
and U25467 (N_25467,N_24853,N_24567);
and U25468 (N_25468,N_24559,N_24818);
and U25469 (N_25469,N_24792,N_24917);
nand U25470 (N_25470,N_24794,N_24855);
xnor U25471 (N_25471,N_24756,N_24645);
and U25472 (N_25472,N_24604,N_24546);
nor U25473 (N_25473,N_24619,N_24540);
xor U25474 (N_25474,N_24771,N_24914);
or U25475 (N_25475,N_24795,N_24888);
xnor U25476 (N_25476,N_24612,N_24651);
or U25477 (N_25477,N_24996,N_24610);
or U25478 (N_25478,N_24730,N_24784);
nand U25479 (N_25479,N_24985,N_24930);
and U25480 (N_25480,N_24766,N_24878);
xnor U25481 (N_25481,N_24547,N_24717);
or U25482 (N_25482,N_24664,N_24682);
or U25483 (N_25483,N_24672,N_24748);
nor U25484 (N_25484,N_24697,N_24978);
and U25485 (N_25485,N_24657,N_24886);
xnor U25486 (N_25486,N_24750,N_24700);
and U25487 (N_25487,N_24677,N_24670);
xor U25488 (N_25488,N_24728,N_24833);
xnor U25489 (N_25489,N_24904,N_24773);
or U25490 (N_25490,N_24832,N_24761);
or U25491 (N_25491,N_24586,N_24655);
nor U25492 (N_25492,N_24708,N_24673);
nor U25493 (N_25493,N_24804,N_24895);
or U25494 (N_25494,N_24575,N_24923);
nor U25495 (N_25495,N_24698,N_24692);
xor U25496 (N_25496,N_24691,N_24638);
xor U25497 (N_25497,N_24637,N_24535);
nand U25498 (N_25498,N_24698,N_24804);
xnor U25499 (N_25499,N_24802,N_24931);
nand U25500 (N_25500,N_25300,N_25319);
and U25501 (N_25501,N_25400,N_25361);
or U25502 (N_25502,N_25110,N_25383);
xnor U25503 (N_25503,N_25075,N_25280);
nor U25504 (N_25504,N_25479,N_25342);
or U25505 (N_25505,N_25092,N_25482);
nor U25506 (N_25506,N_25355,N_25381);
nor U25507 (N_25507,N_25083,N_25344);
or U25508 (N_25508,N_25152,N_25149);
nand U25509 (N_25509,N_25397,N_25379);
xor U25510 (N_25510,N_25273,N_25208);
xnor U25511 (N_25511,N_25061,N_25188);
nor U25512 (N_25512,N_25071,N_25475);
or U25513 (N_25513,N_25348,N_25401);
xnor U25514 (N_25514,N_25121,N_25410);
and U25515 (N_25515,N_25298,N_25173);
xor U25516 (N_25516,N_25105,N_25391);
nand U25517 (N_25517,N_25130,N_25021);
and U25518 (N_25518,N_25328,N_25136);
and U25519 (N_25519,N_25299,N_25050);
nand U25520 (N_25520,N_25179,N_25223);
nor U25521 (N_25521,N_25477,N_25154);
or U25522 (N_25522,N_25473,N_25045);
nand U25523 (N_25523,N_25468,N_25100);
xnor U25524 (N_25524,N_25417,N_25111);
or U25525 (N_25525,N_25404,N_25074);
xor U25526 (N_25526,N_25118,N_25093);
nor U25527 (N_25527,N_25043,N_25448);
nand U25528 (N_25528,N_25425,N_25192);
nand U25529 (N_25529,N_25002,N_25187);
nor U25530 (N_25530,N_25023,N_25172);
nand U25531 (N_25531,N_25016,N_25142);
nand U25532 (N_25532,N_25272,N_25339);
nor U25533 (N_25533,N_25215,N_25120);
or U25534 (N_25534,N_25116,N_25466);
and U25535 (N_25535,N_25214,N_25153);
or U25536 (N_25536,N_25139,N_25488);
or U25537 (N_25537,N_25407,N_25119);
and U25538 (N_25538,N_25206,N_25041);
nand U25539 (N_25539,N_25239,N_25426);
and U25540 (N_25540,N_25487,N_25122);
and U25541 (N_25541,N_25305,N_25308);
or U25542 (N_25542,N_25205,N_25375);
nand U25543 (N_25543,N_25324,N_25220);
xnor U25544 (N_25544,N_25064,N_25144);
nand U25545 (N_25545,N_25387,N_25474);
and U25546 (N_25546,N_25157,N_25447);
nand U25547 (N_25547,N_25285,N_25087);
nor U25548 (N_25548,N_25242,N_25186);
nand U25549 (N_25549,N_25351,N_25039);
or U25550 (N_25550,N_25469,N_25015);
nor U25551 (N_25551,N_25465,N_25143);
nor U25552 (N_25552,N_25322,N_25313);
or U25553 (N_25553,N_25180,N_25085);
and U25554 (N_25554,N_25356,N_25040);
or U25555 (N_25555,N_25017,N_25219);
nor U25556 (N_25556,N_25398,N_25390);
and U25557 (N_25557,N_25073,N_25395);
nand U25558 (N_25558,N_25261,N_25104);
and U25559 (N_25559,N_25102,N_25221);
or U25560 (N_25560,N_25252,N_25081);
and U25561 (N_25561,N_25070,N_25115);
and U25562 (N_25562,N_25485,N_25354);
and U25563 (N_25563,N_25294,N_25067);
nand U25564 (N_25564,N_25042,N_25459);
and U25565 (N_25565,N_25218,N_25441);
nor U25566 (N_25566,N_25278,N_25276);
or U25567 (N_25567,N_25183,N_25006);
xor U25568 (N_25568,N_25283,N_25336);
and U25569 (N_25569,N_25007,N_25442);
xnor U25570 (N_25570,N_25090,N_25229);
nor U25571 (N_25571,N_25321,N_25151);
or U25572 (N_25572,N_25225,N_25303);
nor U25573 (N_25573,N_25416,N_25048);
nand U25574 (N_25574,N_25453,N_25134);
and U25575 (N_25575,N_25211,N_25436);
xor U25576 (N_25576,N_25293,N_25484);
xor U25577 (N_25577,N_25297,N_25369);
nor U25578 (N_25578,N_25076,N_25086);
and U25579 (N_25579,N_25445,N_25231);
or U25580 (N_25580,N_25201,N_25125);
nor U25581 (N_25581,N_25177,N_25176);
or U25582 (N_25582,N_25112,N_25147);
and U25583 (N_25583,N_25254,N_25366);
nand U25584 (N_25584,N_25378,N_25020);
xor U25585 (N_25585,N_25146,N_25331);
and U25586 (N_25586,N_25088,N_25068);
xnor U25587 (N_25587,N_25106,N_25318);
and U25588 (N_25588,N_25423,N_25377);
or U25589 (N_25589,N_25051,N_25160);
nor U25590 (N_25590,N_25138,N_25427);
nand U25591 (N_25591,N_25207,N_25341);
and U25592 (N_25592,N_25026,N_25098);
xor U25593 (N_25593,N_25195,N_25198);
nand U25594 (N_25594,N_25103,N_25168);
and U25595 (N_25595,N_25127,N_25367);
or U25596 (N_25596,N_25150,N_25370);
and U25597 (N_25597,N_25237,N_25360);
xnor U25598 (N_25598,N_25182,N_25422);
nand U25599 (N_25599,N_25114,N_25333);
or U25600 (N_25600,N_25253,N_25164);
or U25601 (N_25601,N_25449,N_25108);
and U25602 (N_25602,N_25190,N_25492);
xnor U25603 (N_25603,N_25058,N_25454);
and U25604 (N_25604,N_25162,N_25347);
and U25605 (N_25605,N_25343,N_25265);
and U25606 (N_25606,N_25287,N_25307);
xor U25607 (N_25607,N_25271,N_25413);
or U25608 (N_25608,N_25311,N_25196);
and U25609 (N_25609,N_25458,N_25066);
nor U25610 (N_25610,N_25148,N_25038);
or U25611 (N_25611,N_25433,N_25184);
xnor U25612 (N_25612,N_25428,N_25212);
nand U25613 (N_25613,N_25117,N_25394);
nand U25614 (N_25614,N_25352,N_25245);
nand U25615 (N_25615,N_25099,N_25364);
nand U25616 (N_25616,N_25419,N_25498);
nand U25617 (N_25617,N_25028,N_25135);
and U25618 (N_25618,N_25248,N_25385);
or U25619 (N_25619,N_25250,N_25317);
or U25620 (N_25620,N_25497,N_25132);
nand U25621 (N_25621,N_25174,N_25141);
and U25622 (N_25622,N_25464,N_25382);
nand U25623 (N_25623,N_25240,N_25025);
and U25624 (N_25624,N_25279,N_25386);
and U25625 (N_25625,N_25290,N_25191);
nor U25626 (N_25626,N_25365,N_25249);
xnor U25627 (N_25627,N_25140,N_25315);
nand U25628 (N_25628,N_25084,N_25309);
nand U25629 (N_25629,N_25096,N_25396);
and U25630 (N_25630,N_25037,N_25241);
and U25631 (N_25631,N_25292,N_25197);
or U25632 (N_25632,N_25209,N_25415);
or U25633 (N_25633,N_25437,N_25392);
and U25634 (N_25634,N_25289,N_25480);
xnor U25635 (N_25635,N_25194,N_25049);
or U25636 (N_25636,N_25330,N_25266);
or U25637 (N_25637,N_25463,N_25384);
nand U25638 (N_25638,N_25471,N_25226);
and U25639 (N_25639,N_25010,N_25052);
nor U25640 (N_25640,N_25044,N_25165);
nand U25641 (N_25641,N_25362,N_25430);
or U25642 (N_25642,N_25284,N_25376);
xor U25643 (N_25643,N_25403,N_25003);
nand U25644 (N_25644,N_25349,N_25388);
and U25645 (N_25645,N_25078,N_25286);
xnor U25646 (N_25646,N_25414,N_25189);
nand U25647 (N_25647,N_25457,N_25082);
xor U25648 (N_25648,N_25033,N_25243);
xor U25649 (N_25649,N_25126,N_25418);
or U25650 (N_25650,N_25259,N_25461);
xor U25651 (N_25651,N_25455,N_25036);
and U25652 (N_25652,N_25200,N_25263);
nor U25653 (N_25653,N_25451,N_25235);
nor U25654 (N_25654,N_25199,N_25247);
or U25655 (N_25655,N_25462,N_25296);
or U25656 (N_25656,N_25268,N_25275);
and U25657 (N_25657,N_25432,N_25238);
or U25658 (N_25658,N_25350,N_25424);
nor U25659 (N_25659,N_25251,N_25359);
and U25660 (N_25660,N_25274,N_25137);
xnor U25661 (N_25661,N_25302,N_25363);
xnor U25662 (N_25662,N_25089,N_25000);
nor U25663 (N_25663,N_25486,N_25421);
or U25664 (N_25664,N_25373,N_25203);
xor U25665 (N_25665,N_25167,N_25262);
nand U25666 (N_25666,N_25499,N_25435);
xnor U25667 (N_25667,N_25326,N_25046);
nand U25668 (N_25668,N_25267,N_25411);
or U25669 (N_25669,N_25054,N_25217);
nand U25670 (N_25670,N_25476,N_25264);
nor U25671 (N_25671,N_25222,N_25358);
nor U25672 (N_25672,N_25008,N_25027);
and U25673 (N_25673,N_25438,N_25439);
xor U25674 (N_25674,N_25277,N_25374);
nand U25675 (N_25675,N_25306,N_25101);
nor U25676 (N_25676,N_25059,N_25269);
nand U25677 (N_25677,N_25327,N_25069);
nand U25678 (N_25678,N_25004,N_25490);
nand U25679 (N_25679,N_25060,N_25478);
xnor U25680 (N_25680,N_25014,N_25224);
xor U25681 (N_25681,N_25314,N_25357);
and U25682 (N_25682,N_25193,N_25345);
nor U25683 (N_25683,N_25062,N_25493);
nor U25684 (N_25684,N_25094,N_25178);
or U25685 (N_25685,N_25338,N_25408);
nor U25686 (N_25686,N_25095,N_25019);
or U25687 (N_25687,N_25133,N_25163);
xnor U25688 (N_25688,N_25109,N_25446);
xnor U25689 (N_25689,N_25030,N_25281);
xor U25690 (N_25690,N_25034,N_25443);
nor U25691 (N_25691,N_25452,N_25246);
and U25692 (N_25692,N_25063,N_25258);
and U25693 (N_25693,N_25053,N_25232);
xnor U25694 (N_25694,N_25181,N_25077);
nor U25695 (N_25695,N_25065,N_25057);
nand U25696 (N_25696,N_25399,N_25337);
or U25697 (N_25697,N_25291,N_25009);
nor U25698 (N_25698,N_25234,N_25320);
nor U25699 (N_25699,N_25420,N_25494);
xnor U25700 (N_25700,N_25012,N_25018);
or U25701 (N_25701,N_25123,N_25204);
or U25702 (N_25702,N_25107,N_25216);
nand U25703 (N_25703,N_25483,N_25389);
xnor U25704 (N_25704,N_25213,N_25032);
nand U25705 (N_25705,N_25295,N_25323);
xor U25706 (N_25706,N_25079,N_25495);
or U25707 (N_25707,N_25288,N_25072);
nand U25708 (N_25708,N_25113,N_25334);
or U25709 (N_25709,N_25166,N_25353);
and U25710 (N_25710,N_25155,N_25380);
nand U25711 (N_25711,N_25450,N_25169);
xor U25712 (N_25712,N_25372,N_25244);
xor U25713 (N_25713,N_25227,N_25145);
or U25714 (N_25714,N_25035,N_25256);
and U25715 (N_25715,N_25460,N_25056);
nand U25716 (N_25716,N_25161,N_25047);
xor U25717 (N_25717,N_25124,N_25260);
or U25718 (N_25718,N_25402,N_25282);
nor U25719 (N_25719,N_25175,N_25013);
or U25720 (N_25720,N_25128,N_25312);
and U25721 (N_25721,N_25316,N_25055);
xor U25722 (N_25722,N_25202,N_25431);
or U25723 (N_25723,N_25470,N_25409);
and U25724 (N_25724,N_25301,N_25310);
xnor U25725 (N_25725,N_25210,N_25022);
nor U25726 (N_25726,N_25097,N_25412);
and U25727 (N_25727,N_25257,N_25005);
xor U25728 (N_25728,N_25171,N_25329);
or U25729 (N_25729,N_25158,N_25491);
or U25730 (N_25730,N_25434,N_25346);
or U25731 (N_25731,N_25001,N_25456);
xor U25732 (N_25732,N_25159,N_25325);
or U25733 (N_25733,N_25405,N_25481);
or U25734 (N_25734,N_25371,N_25011);
nor U25735 (N_25735,N_25129,N_25270);
or U25736 (N_25736,N_25185,N_25080);
or U25737 (N_25737,N_25472,N_25406);
xnor U25738 (N_25738,N_25170,N_25496);
and U25739 (N_25739,N_25467,N_25444);
nor U25740 (N_25740,N_25024,N_25340);
or U25741 (N_25741,N_25131,N_25332);
or U25742 (N_25742,N_25091,N_25228);
and U25743 (N_25743,N_25304,N_25031);
nor U25744 (N_25744,N_25429,N_25156);
xnor U25745 (N_25745,N_25393,N_25335);
and U25746 (N_25746,N_25233,N_25230);
xnor U25747 (N_25747,N_25489,N_25440);
or U25748 (N_25748,N_25255,N_25236);
xnor U25749 (N_25749,N_25029,N_25368);
xnor U25750 (N_25750,N_25072,N_25341);
or U25751 (N_25751,N_25105,N_25406);
and U25752 (N_25752,N_25265,N_25133);
and U25753 (N_25753,N_25152,N_25247);
nand U25754 (N_25754,N_25221,N_25472);
nand U25755 (N_25755,N_25323,N_25029);
or U25756 (N_25756,N_25133,N_25478);
nor U25757 (N_25757,N_25249,N_25401);
nor U25758 (N_25758,N_25013,N_25205);
xor U25759 (N_25759,N_25009,N_25011);
nor U25760 (N_25760,N_25026,N_25091);
or U25761 (N_25761,N_25326,N_25343);
nand U25762 (N_25762,N_25331,N_25105);
or U25763 (N_25763,N_25017,N_25311);
nand U25764 (N_25764,N_25130,N_25364);
nand U25765 (N_25765,N_25268,N_25085);
xor U25766 (N_25766,N_25120,N_25393);
and U25767 (N_25767,N_25332,N_25018);
and U25768 (N_25768,N_25285,N_25230);
or U25769 (N_25769,N_25455,N_25320);
xor U25770 (N_25770,N_25220,N_25399);
nand U25771 (N_25771,N_25230,N_25405);
nor U25772 (N_25772,N_25248,N_25240);
and U25773 (N_25773,N_25161,N_25122);
or U25774 (N_25774,N_25128,N_25417);
or U25775 (N_25775,N_25270,N_25278);
nor U25776 (N_25776,N_25466,N_25389);
nor U25777 (N_25777,N_25226,N_25460);
nand U25778 (N_25778,N_25218,N_25181);
and U25779 (N_25779,N_25157,N_25359);
and U25780 (N_25780,N_25021,N_25097);
nand U25781 (N_25781,N_25313,N_25049);
nor U25782 (N_25782,N_25345,N_25160);
or U25783 (N_25783,N_25145,N_25488);
xor U25784 (N_25784,N_25363,N_25084);
or U25785 (N_25785,N_25424,N_25371);
and U25786 (N_25786,N_25477,N_25378);
or U25787 (N_25787,N_25049,N_25102);
nor U25788 (N_25788,N_25184,N_25196);
xor U25789 (N_25789,N_25225,N_25226);
or U25790 (N_25790,N_25310,N_25173);
or U25791 (N_25791,N_25085,N_25024);
and U25792 (N_25792,N_25000,N_25458);
nor U25793 (N_25793,N_25452,N_25462);
and U25794 (N_25794,N_25375,N_25128);
nand U25795 (N_25795,N_25094,N_25261);
xnor U25796 (N_25796,N_25192,N_25393);
xnor U25797 (N_25797,N_25414,N_25394);
and U25798 (N_25798,N_25203,N_25018);
nand U25799 (N_25799,N_25307,N_25251);
or U25800 (N_25800,N_25288,N_25293);
nand U25801 (N_25801,N_25125,N_25495);
or U25802 (N_25802,N_25233,N_25384);
xor U25803 (N_25803,N_25160,N_25469);
nand U25804 (N_25804,N_25448,N_25424);
and U25805 (N_25805,N_25284,N_25087);
nor U25806 (N_25806,N_25200,N_25021);
xnor U25807 (N_25807,N_25240,N_25015);
nand U25808 (N_25808,N_25134,N_25234);
and U25809 (N_25809,N_25172,N_25160);
or U25810 (N_25810,N_25319,N_25462);
and U25811 (N_25811,N_25415,N_25038);
or U25812 (N_25812,N_25083,N_25245);
and U25813 (N_25813,N_25347,N_25066);
and U25814 (N_25814,N_25156,N_25462);
nand U25815 (N_25815,N_25024,N_25483);
and U25816 (N_25816,N_25179,N_25191);
and U25817 (N_25817,N_25333,N_25036);
or U25818 (N_25818,N_25291,N_25408);
and U25819 (N_25819,N_25480,N_25341);
nor U25820 (N_25820,N_25238,N_25208);
nor U25821 (N_25821,N_25462,N_25306);
xnor U25822 (N_25822,N_25410,N_25497);
xnor U25823 (N_25823,N_25390,N_25160);
nand U25824 (N_25824,N_25181,N_25148);
nor U25825 (N_25825,N_25015,N_25065);
or U25826 (N_25826,N_25440,N_25029);
nor U25827 (N_25827,N_25282,N_25433);
xor U25828 (N_25828,N_25424,N_25250);
xor U25829 (N_25829,N_25261,N_25232);
nor U25830 (N_25830,N_25123,N_25328);
and U25831 (N_25831,N_25184,N_25097);
and U25832 (N_25832,N_25397,N_25206);
and U25833 (N_25833,N_25099,N_25085);
nor U25834 (N_25834,N_25128,N_25316);
and U25835 (N_25835,N_25201,N_25196);
or U25836 (N_25836,N_25024,N_25174);
and U25837 (N_25837,N_25376,N_25038);
and U25838 (N_25838,N_25385,N_25233);
nor U25839 (N_25839,N_25493,N_25164);
nor U25840 (N_25840,N_25215,N_25153);
nand U25841 (N_25841,N_25397,N_25146);
nor U25842 (N_25842,N_25147,N_25163);
or U25843 (N_25843,N_25344,N_25207);
nand U25844 (N_25844,N_25356,N_25161);
and U25845 (N_25845,N_25456,N_25283);
xor U25846 (N_25846,N_25341,N_25204);
nor U25847 (N_25847,N_25313,N_25094);
and U25848 (N_25848,N_25493,N_25095);
and U25849 (N_25849,N_25377,N_25470);
or U25850 (N_25850,N_25272,N_25494);
nor U25851 (N_25851,N_25150,N_25144);
or U25852 (N_25852,N_25120,N_25318);
xnor U25853 (N_25853,N_25461,N_25319);
nand U25854 (N_25854,N_25064,N_25345);
nand U25855 (N_25855,N_25460,N_25095);
nor U25856 (N_25856,N_25162,N_25423);
or U25857 (N_25857,N_25183,N_25384);
nor U25858 (N_25858,N_25166,N_25417);
nand U25859 (N_25859,N_25093,N_25368);
or U25860 (N_25860,N_25089,N_25020);
nand U25861 (N_25861,N_25170,N_25027);
xnor U25862 (N_25862,N_25142,N_25371);
nand U25863 (N_25863,N_25040,N_25420);
nor U25864 (N_25864,N_25124,N_25020);
or U25865 (N_25865,N_25498,N_25000);
or U25866 (N_25866,N_25211,N_25006);
nand U25867 (N_25867,N_25213,N_25331);
or U25868 (N_25868,N_25015,N_25448);
nor U25869 (N_25869,N_25053,N_25190);
xor U25870 (N_25870,N_25067,N_25178);
xor U25871 (N_25871,N_25297,N_25251);
nor U25872 (N_25872,N_25123,N_25434);
xor U25873 (N_25873,N_25095,N_25002);
xnor U25874 (N_25874,N_25247,N_25261);
and U25875 (N_25875,N_25186,N_25381);
nor U25876 (N_25876,N_25272,N_25456);
nand U25877 (N_25877,N_25454,N_25047);
nand U25878 (N_25878,N_25499,N_25198);
or U25879 (N_25879,N_25386,N_25463);
or U25880 (N_25880,N_25054,N_25011);
nand U25881 (N_25881,N_25125,N_25263);
nand U25882 (N_25882,N_25170,N_25010);
nand U25883 (N_25883,N_25144,N_25252);
and U25884 (N_25884,N_25450,N_25224);
nand U25885 (N_25885,N_25185,N_25207);
or U25886 (N_25886,N_25294,N_25206);
nand U25887 (N_25887,N_25090,N_25195);
or U25888 (N_25888,N_25087,N_25001);
xor U25889 (N_25889,N_25159,N_25373);
nand U25890 (N_25890,N_25265,N_25104);
and U25891 (N_25891,N_25127,N_25025);
nand U25892 (N_25892,N_25250,N_25311);
nor U25893 (N_25893,N_25363,N_25101);
nor U25894 (N_25894,N_25006,N_25435);
nor U25895 (N_25895,N_25499,N_25448);
nor U25896 (N_25896,N_25499,N_25027);
nand U25897 (N_25897,N_25315,N_25481);
or U25898 (N_25898,N_25081,N_25177);
nor U25899 (N_25899,N_25300,N_25428);
nand U25900 (N_25900,N_25337,N_25049);
xnor U25901 (N_25901,N_25234,N_25155);
and U25902 (N_25902,N_25381,N_25451);
nor U25903 (N_25903,N_25152,N_25456);
nor U25904 (N_25904,N_25070,N_25268);
and U25905 (N_25905,N_25261,N_25160);
xnor U25906 (N_25906,N_25261,N_25240);
nor U25907 (N_25907,N_25078,N_25094);
nor U25908 (N_25908,N_25329,N_25164);
and U25909 (N_25909,N_25169,N_25422);
or U25910 (N_25910,N_25477,N_25128);
nor U25911 (N_25911,N_25141,N_25420);
and U25912 (N_25912,N_25492,N_25478);
xnor U25913 (N_25913,N_25013,N_25471);
or U25914 (N_25914,N_25379,N_25276);
nor U25915 (N_25915,N_25068,N_25220);
and U25916 (N_25916,N_25202,N_25476);
or U25917 (N_25917,N_25354,N_25184);
and U25918 (N_25918,N_25417,N_25310);
xor U25919 (N_25919,N_25279,N_25185);
nor U25920 (N_25920,N_25356,N_25105);
xnor U25921 (N_25921,N_25056,N_25244);
xor U25922 (N_25922,N_25178,N_25351);
xor U25923 (N_25923,N_25018,N_25104);
nor U25924 (N_25924,N_25043,N_25027);
xnor U25925 (N_25925,N_25420,N_25113);
or U25926 (N_25926,N_25489,N_25494);
and U25927 (N_25927,N_25238,N_25040);
xor U25928 (N_25928,N_25332,N_25100);
or U25929 (N_25929,N_25296,N_25198);
xnor U25930 (N_25930,N_25003,N_25293);
xor U25931 (N_25931,N_25058,N_25334);
nand U25932 (N_25932,N_25297,N_25144);
nor U25933 (N_25933,N_25076,N_25299);
nor U25934 (N_25934,N_25207,N_25468);
or U25935 (N_25935,N_25199,N_25417);
or U25936 (N_25936,N_25150,N_25425);
and U25937 (N_25937,N_25174,N_25410);
and U25938 (N_25938,N_25257,N_25353);
nor U25939 (N_25939,N_25213,N_25103);
xor U25940 (N_25940,N_25068,N_25054);
or U25941 (N_25941,N_25320,N_25219);
and U25942 (N_25942,N_25299,N_25276);
nand U25943 (N_25943,N_25045,N_25123);
and U25944 (N_25944,N_25236,N_25240);
and U25945 (N_25945,N_25162,N_25163);
and U25946 (N_25946,N_25467,N_25386);
nor U25947 (N_25947,N_25427,N_25127);
nand U25948 (N_25948,N_25475,N_25277);
nand U25949 (N_25949,N_25378,N_25174);
or U25950 (N_25950,N_25416,N_25334);
nor U25951 (N_25951,N_25357,N_25450);
and U25952 (N_25952,N_25183,N_25484);
xor U25953 (N_25953,N_25200,N_25307);
xnor U25954 (N_25954,N_25105,N_25430);
nand U25955 (N_25955,N_25387,N_25115);
xor U25956 (N_25956,N_25176,N_25381);
and U25957 (N_25957,N_25334,N_25123);
and U25958 (N_25958,N_25420,N_25498);
nand U25959 (N_25959,N_25172,N_25279);
or U25960 (N_25960,N_25419,N_25327);
xor U25961 (N_25961,N_25426,N_25494);
nand U25962 (N_25962,N_25125,N_25497);
nor U25963 (N_25963,N_25235,N_25428);
xor U25964 (N_25964,N_25478,N_25444);
nand U25965 (N_25965,N_25161,N_25083);
nand U25966 (N_25966,N_25284,N_25425);
nor U25967 (N_25967,N_25360,N_25047);
nor U25968 (N_25968,N_25042,N_25410);
or U25969 (N_25969,N_25057,N_25258);
nor U25970 (N_25970,N_25235,N_25206);
nor U25971 (N_25971,N_25255,N_25073);
nand U25972 (N_25972,N_25192,N_25194);
xor U25973 (N_25973,N_25153,N_25365);
nor U25974 (N_25974,N_25100,N_25185);
or U25975 (N_25975,N_25073,N_25210);
nand U25976 (N_25976,N_25406,N_25045);
nor U25977 (N_25977,N_25000,N_25383);
xor U25978 (N_25978,N_25465,N_25402);
xnor U25979 (N_25979,N_25170,N_25476);
nor U25980 (N_25980,N_25466,N_25122);
or U25981 (N_25981,N_25320,N_25490);
nand U25982 (N_25982,N_25009,N_25184);
and U25983 (N_25983,N_25203,N_25128);
xnor U25984 (N_25984,N_25464,N_25352);
and U25985 (N_25985,N_25051,N_25034);
nor U25986 (N_25986,N_25242,N_25166);
nor U25987 (N_25987,N_25402,N_25100);
and U25988 (N_25988,N_25185,N_25343);
and U25989 (N_25989,N_25178,N_25111);
xor U25990 (N_25990,N_25367,N_25140);
and U25991 (N_25991,N_25479,N_25349);
nand U25992 (N_25992,N_25153,N_25101);
or U25993 (N_25993,N_25450,N_25479);
nor U25994 (N_25994,N_25036,N_25011);
and U25995 (N_25995,N_25462,N_25377);
and U25996 (N_25996,N_25328,N_25134);
nor U25997 (N_25997,N_25006,N_25268);
nor U25998 (N_25998,N_25245,N_25096);
nor U25999 (N_25999,N_25359,N_25417);
nor U26000 (N_26000,N_25835,N_25673);
nor U26001 (N_26001,N_25860,N_25740);
nor U26002 (N_26002,N_25664,N_25517);
nor U26003 (N_26003,N_25595,N_25568);
xnor U26004 (N_26004,N_25756,N_25791);
and U26005 (N_26005,N_25563,N_25620);
or U26006 (N_26006,N_25540,N_25840);
nand U26007 (N_26007,N_25799,N_25846);
nor U26008 (N_26008,N_25898,N_25886);
and U26009 (N_26009,N_25985,N_25688);
xnor U26010 (N_26010,N_25739,N_25809);
xnor U26011 (N_26011,N_25694,N_25948);
nor U26012 (N_26012,N_25735,N_25677);
or U26013 (N_26013,N_25807,N_25648);
or U26014 (N_26014,N_25612,N_25858);
xnor U26015 (N_26015,N_25770,N_25854);
xor U26016 (N_26016,N_25779,N_25908);
nand U26017 (N_26017,N_25843,N_25988);
nand U26018 (N_26018,N_25716,N_25700);
nand U26019 (N_26019,N_25682,N_25755);
or U26020 (N_26020,N_25573,N_25668);
nand U26021 (N_26021,N_25610,N_25781);
nand U26022 (N_26022,N_25519,N_25891);
or U26023 (N_26023,N_25530,N_25941);
nor U26024 (N_26024,N_25827,N_25670);
nand U26025 (N_26025,N_25650,N_25982);
and U26026 (N_26026,N_25732,N_25832);
or U26027 (N_26027,N_25798,N_25775);
and U26028 (N_26028,N_25511,N_25584);
and U26029 (N_26029,N_25880,N_25917);
nor U26030 (N_26030,N_25533,N_25606);
nand U26031 (N_26031,N_25872,N_25793);
and U26032 (N_26032,N_25507,N_25868);
xnor U26033 (N_26033,N_25696,N_25580);
nand U26034 (N_26034,N_25713,N_25721);
and U26035 (N_26035,N_25502,N_25587);
nand U26036 (N_26036,N_25959,N_25744);
or U26037 (N_26037,N_25725,N_25548);
nor U26038 (N_26038,N_25776,N_25510);
nor U26039 (N_26039,N_25594,N_25984);
nor U26040 (N_26040,N_25593,N_25869);
or U26041 (N_26041,N_25963,N_25904);
xor U26042 (N_26042,N_25845,N_25741);
xnor U26043 (N_26043,N_25585,N_25557);
and U26044 (N_26044,N_25718,N_25635);
xor U26045 (N_26045,N_25609,N_25778);
or U26046 (N_26046,N_25693,N_25676);
xor U26047 (N_26047,N_25911,N_25802);
or U26048 (N_26048,N_25737,N_25569);
xor U26049 (N_26049,N_25782,N_25634);
xor U26050 (N_26050,N_25893,N_25929);
xor U26051 (N_26051,N_25539,N_25598);
nor U26052 (N_26052,N_25932,N_25754);
or U26053 (N_26053,N_25980,N_25986);
and U26054 (N_26054,N_25976,N_25686);
nand U26055 (N_26055,N_25897,N_25852);
nor U26056 (N_26056,N_25998,N_25611);
and U26057 (N_26057,N_25909,N_25603);
nor U26058 (N_26058,N_25816,N_25863);
and U26059 (N_26059,N_25810,N_25605);
nand U26060 (N_26060,N_25643,N_25652);
and U26061 (N_26061,N_25995,N_25947);
nand U26062 (N_26062,N_25830,N_25766);
nand U26063 (N_26063,N_25964,N_25831);
xor U26064 (N_26064,N_25742,N_25990);
nand U26065 (N_26065,N_25535,N_25637);
or U26066 (N_26066,N_25551,N_25906);
or U26067 (N_26067,N_25687,N_25822);
nand U26068 (N_26068,N_25559,N_25654);
or U26069 (N_26069,N_25850,N_25567);
nand U26070 (N_26070,N_25892,N_25834);
nor U26071 (N_26071,N_25973,N_25921);
xnor U26072 (N_26072,N_25987,N_25758);
xnor U26073 (N_26073,N_25545,N_25707);
nor U26074 (N_26074,N_25797,N_25592);
nand U26075 (N_26075,N_25949,N_25523);
xnor U26076 (N_26076,N_25599,N_25513);
or U26077 (N_26077,N_25547,N_25556);
and U26078 (N_26078,N_25621,N_25727);
and U26079 (N_26079,N_25862,N_25975);
or U26080 (N_26080,N_25820,N_25704);
nor U26081 (N_26081,N_25882,N_25943);
xnor U26082 (N_26082,N_25914,N_25967);
nand U26083 (N_26083,N_25788,N_25812);
nor U26084 (N_26084,N_25814,N_25570);
xnor U26085 (N_26085,N_25660,N_25936);
and U26086 (N_26086,N_25656,N_25583);
and U26087 (N_26087,N_25819,N_25711);
and U26088 (N_26088,N_25581,N_25504);
nor U26089 (N_26089,N_25920,N_25870);
xor U26090 (N_26090,N_25828,N_25544);
xnor U26091 (N_26091,N_25528,N_25708);
nand U26092 (N_26092,N_25780,N_25759);
nor U26093 (N_26093,N_25684,N_25919);
nand U26094 (N_26094,N_25726,N_25743);
and U26095 (N_26095,N_25745,N_25526);
xor U26096 (N_26096,N_25903,N_25918);
nor U26097 (N_26097,N_25794,N_25757);
nor U26098 (N_26098,N_25895,N_25768);
and U26099 (N_26099,N_25763,N_25666);
nand U26100 (N_26100,N_25833,N_25695);
nand U26101 (N_26101,N_25930,N_25717);
nand U26102 (N_26102,N_25628,N_25715);
and U26103 (N_26103,N_25789,N_25894);
nand U26104 (N_26104,N_25508,N_25829);
xnor U26105 (N_26105,N_25887,N_25588);
or U26106 (N_26106,N_25848,N_25590);
nor U26107 (N_26107,N_25997,N_25871);
xnor U26108 (N_26108,N_25912,N_25983);
or U26109 (N_26109,N_25719,N_25579);
nand U26110 (N_26110,N_25974,N_25591);
nor U26111 (N_26111,N_25817,N_25730);
and U26112 (N_26112,N_25578,N_25999);
nor U26113 (N_26113,N_25626,N_25589);
nor U26114 (N_26114,N_25746,N_25646);
and U26115 (N_26115,N_25979,N_25636);
or U26116 (N_26116,N_25572,N_25600);
nor U26117 (N_26117,N_25859,N_25942);
and U26118 (N_26118,N_25857,N_25630);
xor U26119 (N_26119,N_25773,N_25796);
and U26120 (N_26120,N_25981,N_25888);
nand U26121 (N_26121,N_25965,N_25795);
nor U26122 (N_26122,N_25709,N_25762);
or U26123 (N_26123,N_25826,N_25771);
xnor U26124 (N_26124,N_25808,N_25764);
nand U26125 (N_26125,N_25625,N_25607);
nand U26126 (N_26126,N_25501,N_25518);
or U26127 (N_26127,N_25699,N_25790);
nor U26128 (N_26128,N_25777,N_25847);
and U26129 (N_26129,N_25861,N_25978);
nor U26130 (N_26130,N_25885,N_25939);
and U26131 (N_26131,N_25825,N_25516);
or U26132 (N_26132,N_25608,N_25706);
xor U26133 (N_26133,N_25747,N_25968);
and U26134 (N_26134,N_25916,N_25989);
nand U26135 (N_26135,N_25824,N_25627);
nand U26136 (N_26136,N_25541,N_25734);
nor U26137 (N_26137,N_25750,N_25966);
nor U26138 (N_26138,N_25615,N_25549);
nand U26139 (N_26139,N_25783,N_25878);
and U26140 (N_26140,N_25867,N_25616);
xor U26141 (N_26141,N_25554,N_25765);
nor U26142 (N_26142,N_25524,N_25738);
nor U26143 (N_26143,N_25565,N_25881);
or U26144 (N_26144,N_25619,N_25969);
nor U26145 (N_26145,N_25683,N_25604);
and U26146 (N_26146,N_25803,N_25701);
and U26147 (N_26147,N_25576,N_25566);
or U26148 (N_26148,N_25691,N_25937);
or U26149 (N_26149,N_25681,N_25784);
nor U26150 (N_26150,N_25574,N_25586);
xor U26151 (N_26151,N_25955,N_25890);
and U26152 (N_26152,N_25953,N_25512);
nand U26153 (N_26153,N_25582,N_25724);
nor U26154 (N_26154,N_25851,N_25531);
nor U26155 (N_26155,N_25896,N_25875);
or U26156 (N_26156,N_25640,N_25749);
xor U26157 (N_26157,N_25876,N_25503);
xnor U26158 (N_26158,N_25752,N_25924);
xor U26159 (N_26159,N_25927,N_25658);
nor U26160 (N_26160,N_25602,N_25877);
nor U26161 (N_26161,N_25655,N_25651);
and U26162 (N_26162,N_25804,N_25506);
nand U26163 (N_26163,N_25561,N_25690);
nand U26164 (N_26164,N_25913,N_25785);
nand U26165 (N_26165,N_25991,N_25992);
xnor U26166 (N_26166,N_25856,N_25552);
and U26167 (N_26167,N_25613,N_25933);
or U26168 (N_26168,N_25662,N_25546);
or U26169 (N_26169,N_25571,N_25874);
xor U26170 (N_26170,N_25527,N_25994);
nand U26171 (N_26171,N_25761,N_25926);
or U26172 (N_26172,N_25931,N_25962);
nor U26173 (N_26173,N_25672,N_25597);
and U26174 (N_26174,N_25925,N_25748);
nand U26175 (N_26175,N_25884,N_25663);
nand U26176 (N_26176,N_25614,N_25558);
nand U26177 (N_26177,N_25515,N_25902);
or U26178 (N_26178,N_25542,N_25792);
xor U26179 (N_26179,N_25760,N_25639);
nand U26180 (N_26180,N_25769,N_25751);
or U26181 (N_26181,N_25647,N_25883);
nand U26182 (N_26182,N_25534,N_25631);
or U26183 (N_26183,N_25865,N_25813);
nor U26184 (N_26184,N_25720,N_25522);
and U26185 (N_26185,N_25529,N_25899);
xor U26186 (N_26186,N_25946,N_25629);
nor U26187 (N_26187,N_25632,N_25692);
nor U26188 (N_26188,N_25901,N_25514);
and U26189 (N_26189,N_25910,N_25623);
xnor U26190 (N_26190,N_25849,N_25944);
xnor U26191 (N_26191,N_25905,N_25577);
or U26192 (N_26192,N_25786,N_25818);
and U26193 (N_26193,N_25657,N_25772);
nand U26194 (N_26194,N_25520,N_25853);
or U26195 (N_26195,N_25633,N_25705);
and U26196 (N_26196,N_25889,N_25841);
and U26197 (N_26197,N_25806,N_25767);
or U26198 (N_26198,N_25731,N_25564);
nand U26199 (N_26199,N_25642,N_25753);
and U26200 (N_26200,N_25601,N_25938);
or U26201 (N_26201,N_25972,N_25971);
and U26202 (N_26202,N_25675,N_25679);
nor U26203 (N_26203,N_25934,N_25823);
nor U26204 (N_26204,N_25710,N_25500);
nor U26205 (N_26205,N_25935,N_25815);
and U26206 (N_26206,N_25555,N_25970);
xnor U26207 (N_26207,N_25618,N_25509);
and U26208 (N_26208,N_25900,N_25617);
or U26209 (N_26209,N_25532,N_25952);
xnor U26210 (N_26210,N_25907,N_25915);
nand U26211 (N_26211,N_25560,N_25689);
nor U26212 (N_26212,N_25993,N_25838);
nor U26213 (N_26213,N_25956,N_25641);
nand U26214 (N_26214,N_25622,N_25712);
xor U26215 (N_26215,N_25703,N_25958);
nand U26216 (N_26216,N_25698,N_25680);
nor U26217 (N_26217,N_25553,N_25787);
nor U26218 (N_26218,N_25678,N_25821);
nand U26219 (N_26219,N_25575,N_25811);
xor U26220 (N_26220,N_25644,N_25729);
or U26221 (N_26221,N_25665,N_25536);
and U26222 (N_26222,N_25928,N_25645);
nor U26223 (N_26223,N_25844,N_25722);
nor U26224 (N_26224,N_25659,N_25922);
nor U26225 (N_26225,N_25702,N_25805);
nand U26226 (N_26226,N_25638,N_25669);
and U26227 (N_26227,N_25940,N_25550);
nand U26228 (N_26228,N_25774,N_25661);
and U26229 (N_26229,N_25977,N_25951);
nor U26230 (N_26230,N_25537,N_25723);
and U26231 (N_26231,N_25624,N_25697);
nor U26232 (N_26232,N_25923,N_25525);
nor U26233 (N_26233,N_25842,N_25957);
nor U26234 (N_26234,N_25538,N_25837);
xnor U26235 (N_26235,N_25873,N_25653);
nand U26236 (N_26236,N_25801,N_25685);
or U26237 (N_26237,N_25800,N_25596);
nor U26238 (N_26238,N_25714,N_25674);
and U26239 (N_26239,N_25667,N_25954);
and U26240 (N_26240,N_25866,N_25950);
nor U26241 (N_26241,N_25733,N_25736);
or U26242 (N_26242,N_25864,N_25855);
nand U26243 (N_26243,N_25960,N_25996);
nor U26244 (N_26244,N_25879,N_25521);
nor U26245 (N_26245,N_25649,N_25961);
nor U26246 (N_26246,N_25839,N_25543);
nor U26247 (N_26247,N_25945,N_25836);
or U26248 (N_26248,N_25671,N_25505);
nor U26249 (N_26249,N_25728,N_25562);
nand U26250 (N_26250,N_25667,N_25861);
nor U26251 (N_26251,N_25543,N_25727);
nor U26252 (N_26252,N_25923,N_25771);
xor U26253 (N_26253,N_25810,N_25899);
nor U26254 (N_26254,N_25851,N_25738);
nor U26255 (N_26255,N_25521,N_25592);
or U26256 (N_26256,N_25947,N_25513);
xor U26257 (N_26257,N_25641,N_25610);
xnor U26258 (N_26258,N_25841,N_25930);
xor U26259 (N_26259,N_25909,N_25987);
nor U26260 (N_26260,N_25710,N_25613);
nand U26261 (N_26261,N_25651,N_25596);
nor U26262 (N_26262,N_25538,N_25544);
or U26263 (N_26263,N_25897,N_25789);
and U26264 (N_26264,N_25681,N_25986);
or U26265 (N_26265,N_25820,N_25863);
nor U26266 (N_26266,N_25649,N_25730);
nor U26267 (N_26267,N_25554,N_25858);
and U26268 (N_26268,N_25869,N_25611);
and U26269 (N_26269,N_25897,N_25705);
and U26270 (N_26270,N_25775,N_25965);
xor U26271 (N_26271,N_25534,N_25779);
nand U26272 (N_26272,N_25677,N_25944);
or U26273 (N_26273,N_25876,N_25866);
nand U26274 (N_26274,N_25982,N_25816);
or U26275 (N_26275,N_25782,N_25743);
and U26276 (N_26276,N_25875,N_25524);
and U26277 (N_26277,N_25826,N_25912);
nor U26278 (N_26278,N_25929,N_25772);
xnor U26279 (N_26279,N_25609,N_25685);
nor U26280 (N_26280,N_25959,N_25653);
and U26281 (N_26281,N_25858,N_25870);
and U26282 (N_26282,N_25886,N_25644);
and U26283 (N_26283,N_25967,N_25617);
and U26284 (N_26284,N_25915,N_25672);
xnor U26285 (N_26285,N_25614,N_25630);
xor U26286 (N_26286,N_25605,N_25719);
xor U26287 (N_26287,N_25732,N_25594);
nor U26288 (N_26288,N_25849,N_25705);
xor U26289 (N_26289,N_25554,N_25666);
or U26290 (N_26290,N_25934,N_25892);
nor U26291 (N_26291,N_25780,N_25909);
nand U26292 (N_26292,N_25961,N_25563);
or U26293 (N_26293,N_25545,N_25861);
nand U26294 (N_26294,N_25507,N_25760);
nand U26295 (N_26295,N_25912,N_25519);
nand U26296 (N_26296,N_25778,N_25501);
nor U26297 (N_26297,N_25936,N_25908);
nor U26298 (N_26298,N_25729,N_25519);
and U26299 (N_26299,N_25972,N_25687);
or U26300 (N_26300,N_25686,N_25917);
or U26301 (N_26301,N_25696,N_25724);
xor U26302 (N_26302,N_25965,N_25606);
nor U26303 (N_26303,N_25657,N_25706);
and U26304 (N_26304,N_25975,N_25706);
xor U26305 (N_26305,N_25881,N_25818);
xor U26306 (N_26306,N_25974,N_25875);
nor U26307 (N_26307,N_25909,N_25620);
or U26308 (N_26308,N_25741,N_25965);
xor U26309 (N_26309,N_25733,N_25643);
or U26310 (N_26310,N_25677,N_25830);
nor U26311 (N_26311,N_25829,N_25957);
nor U26312 (N_26312,N_25606,N_25647);
nor U26313 (N_26313,N_25836,N_25702);
and U26314 (N_26314,N_25763,N_25600);
xnor U26315 (N_26315,N_25661,N_25531);
or U26316 (N_26316,N_25593,N_25950);
nor U26317 (N_26317,N_25889,N_25506);
xnor U26318 (N_26318,N_25908,N_25764);
nand U26319 (N_26319,N_25571,N_25549);
or U26320 (N_26320,N_25969,N_25753);
nor U26321 (N_26321,N_25599,N_25926);
xnor U26322 (N_26322,N_25715,N_25810);
and U26323 (N_26323,N_25823,N_25717);
and U26324 (N_26324,N_25991,N_25687);
and U26325 (N_26325,N_25782,N_25562);
nor U26326 (N_26326,N_25538,N_25715);
nand U26327 (N_26327,N_25757,N_25784);
xor U26328 (N_26328,N_25680,N_25687);
or U26329 (N_26329,N_25845,N_25533);
xor U26330 (N_26330,N_25849,N_25819);
and U26331 (N_26331,N_25709,N_25914);
or U26332 (N_26332,N_25852,N_25854);
xnor U26333 (N_26333,N_25945,N_25727);
xnor U26334 (N_26334,N_25857,N_25526);
nand U26335 (N_26335,N_25537,N_25755);
nor U26336 (N_26336,N_25753,N_25678);
or U26337 (N_26337,N_25976,N_25560);
nor U26338 (N_26338,N_25622,N_25966);
nor U26339 (N_26339,N_25897,N_25973);
and U26340 (N_26340,N_25611,N_25885);
xnor U26341 (N_26341,N_25648,N_25730);
nor U26342 (N_26342,N_25755,N_25522);
and U26343 (N_26343,N_25649,N_25963);
nand U26344 (N_26344,N_25858,N_25901);
nor U26345 (N_26345,N_25526,N_25750);
nor U26346 (N_26346,N_25842,N_25857);
xor U26347 (N_26347,N_25689,N_25691);
nor U26348 (N_26348,N_25984,N_25530);
and U26349 (N_26349,N_25550,N_25758);
nor U26350 (N_26350,N_25872,N_25779);
or U26351 (N_26351,N_25693,N_25603);
nand U26352 (N_26352,N_25907,N_25821);
xor U26353 (N_26353,N_25556,N_25655);
or U26354 (N_26354,N_25559,N_25545);
or U26355 (N_26355,N_25639,N_25852);
and U26356 (N_26356,N_25632,N_25963);
nand U26357 (N_26357,N_25974,N_25554);
nand U26358 (N_26358,N_25828,N_25604);
or U26359 (N_26359,N_25511,N_25726);
xor U26360 (N_26360,N_25822,N_25694);
or U26361 (N_26361,N_25956,N_25850);
xor U26362 (N_26362,N_25886,N_25511);
and U26363 (N_26363,N_25927,N_25791);
nor U26364 (N_26364,N_25872,N_25531);
nor U26365 (N_26365,N_25630,N_25521);
and U26366 (N_26366,N_25675,N_25704);
or U26367 (N_26367,N_25767,N_25930);
nand U26368 (N_26368,N_25912,N_25977);
or U26369 (N_26369,N_25881,N_25692);
xnor U26370 (N_26370,N_25571,N_25740);
xor U26371 (N_26371,N_25737,N_25697);
nor U26372 (N_26372,N_25885,N_25600);
xnor U26373 (N_26373,N_25789,N_25954);
or U26374 (N_26374,N_25721,N_25522);
xor U26375 (N_26375,N_25508,N_25604);
nor U26376 (N_26376,N_25978,N_25616);
and U26377 (N_26377,N_25981,N_25840);
nor U26378 (N_26378,N_25693,N_25724);
nand U26379 (N_26379,N_25691,N_25891);
nor U26380 (N_26380,N_25618,N_25710);
or U26381 (N_26381,N_25726,N_25561);
xor U26382 (N_26382,N_25694,N_25527);
and U26383 (N_26383,N_25628,N_25927);
xor U26384 (N_26384,N_25934,N_25921);
xor U26385 (N_26385,N_25722,N_25876);
or U26386 (N_26386,N_25931,N_25528);
or U26387 (N_26387,N_25611,N_25999);
and U26388 (N_26388,N_25873,N_25785);
nor U26389 (N_26389,N_25844,N_25551);
or U26390 (N_26390,N_25925,N_25522);
and U26391 (N_26391,N_25919,N_25932);
or U26392 (N_26392,N_25816,N_25701);
nor U26393 (N_26393,N_25935,N_25693);
and U26394 (N_26394,N_25834,N_25887);
xor U26395 (N_26395,N_25821,N_25585);
and U26396 (N_26396,N_25548,N_25984);
xor U26397 (N_26397,N_25636,N_25566);
and U26398 (N_26398,N_25677,N_25734);
and U26399 (N_26399,N_25867,N_25796);
nand U26400 (N_26400,N_25742,N_25521);
nor U26401 (N_26401,N_25705,N_25883);
nor U26402 (N_26402,N_25865,N_25962);
nor U26403 (N_26403,N_25592,N_25626);
and U26404 (N_26404,N_25626,N_25884);
xor U26405 (N_26405,N_25566,N_25648);
xnor U26406 (N_26406,N_25823,N_25822);
xor U26407 (N_26407,N_25811,N_25736);
and U26408 (N_26408,N_25652,N_25588);
or U26409 (N_26409,N_25723,N_25785);
or U26410 (N_26410,N_25745,N_25756);
or U26411 (N_26411,N_25623,N_25568);
xor U26412 (N_26412,N_25672,N_25612);
and U26413 (N_26413,N_25807,N_25703);
and U26414 (N_26414,N_25745,N_25966);
nand U26415 (N_26415,N_25572,N_25503);
nor U26416 (N_26416,N_25803,N_25550);
nand U26417 (N_26417,N_25531,N_25547);
nor U26418 (N_26418,N_25837,N_25812);
nand U26419 (N_26419,N_25893,N_25884);
and U26420 (N_26420,N_25568,N_25922);
nor U26421 (N_26421,N_25599,N_25880);
and U26422 (N_26422,N_25508,N_25699);
nand U26423 (N_26423,N_25954,N_25969);
and U26424 (N_26424,N_25558,N_25666);
or U26425 (N_26425,N_25532,N_25587);
nor U26426 (N_26426,N_25759,N_25577);
nor U26427 (N_26427,N_25637,N_25645);
nor U26428 (N_26428,N_25935,N_25581);
xnor U26429 (N_26429,N_25815,N_25538);
nand U26430 (N_26430,N_25633,N_25765);
nor U26431 (N_26431,N_25544,N_25917);
or U26432 (N_26432,N_25900,N_25758);
and U26433 (N_26433,N_25644,N_25718);
and U26434 (N_26434,N_25986,N_25841);
nand U26435 (N_26435,N_25895,N_25777);
nand U26436 (N_26436,N_25864,N_25704);
and U26437 (N_26437,N_25531,N_25572);
nand U26438 (N_26438,N_25972,N_25869);
nor U26439 (N_26439,N_25747,N_25702);
or U26440 (N_26440,N_25975,N_25685);
or U26441 (N_26441,N_25849,N_25572);
xor U26442 (N_26442,N_25551,N_25678);
and U26443 (N_26443,N_25768,N_25668);
nand U26444 (N_26444,N_25762,N_25877);
and U26445 (N_26445,N_25712,N_25901);
nand U26446 (N_26446,N_25567,N_25655);
or U26447 (N_26447,N_25521,N_25652);
nand U26448 (N_26448,N_25681,N_25977);
or U26449 (N_26449,N_25659,N_25822);
nand U26450 (N_26450,N_25823,N_25722);
nand U26451 (N_26451,N_25515,N_25864);
and U26452 (N_26452,N_25848,N_25779);
nand U26453 (N_26453,N_25716,N_25662);
xor U26454 (N_26454,N_25550,N_25687);
and U26455 (N_26455,N_25613,N_25712);
nor U26456 (N_26456,N_25992,N_25559);
nor U26457 (N_26457,N_25984,N_25931);
nor U26458 (N_26458,N_25743,N_25912);
and U26459 (N_26459,N_25519,N_25910);
nand U26460 (N_26460,N_25952,N_25777);
and U26461 (N_26461,N_25945,N_25967);
nor U26462 (N_26462,N_25665,N_25772);
and U26463 (N_26463,N_25724,N_25702);
xor U26464 (N_26464,N_25539,N_25581);
and U26465 (N_26465,N_25886,N_25769);
nand U26466 (N_26466,N_25804,N_25690);
and U26467 (N_26467,N_25604,N_25869);
nor U26468 (N_26468,N_25687,N_25549);
and U26469 (N_26469,N_25790,N_25573);
xor U26470 (N_26470,N_25938,N_25571);
nand U26471 (N_26471,N_25870,N_25893);
and U26472 (N_26472,N_25504,N_25697);
nor U26473 (N_26473,N_25748,N_25539);
or U26474 (N_26474,N_25555,N_25800);
or U26475 (N_26475,N_25966,N_25984);
and U26476 (N_26476,N_25763,N_25995);
and U26477 (N_26477,N_25676,N_25701);
nand U26478 (N_26478,N_25899,N_25655);
nand U26479 (N_26479,N_25890,N_25900);
and U26480 (N_26480,N_25518,N_25602);
or U26481 (N_26481,N_25998,N_25628);
nand U26482 (N_26482,N_25838,N_25704);
or U26483 (N_26483,N_25846,N_25773);
nor U26484 (N_26484,N_25786,N_25700);
xnor U26485 (N_26485,N_25848,N_25899);
nor U26486 (N_26486,N_25982,N_25778);
nand U26487 (N_26487,N_25920,N_25834);
xor U26488 (N_26488,N_25502,N_25843);
xnor U26489 (N_26489,N_25959,N_25978);
and U26490 (N_26490,N_25994,N_25952);
nor U26491 (N_26491,N_25757,N_25510);
xor U26492 (N_26492,N_25808,N_25594);
xor U26493 (N_26493,N_25678,N_25993);
or U26494 (N_26494,N_25703,N_25616);
nand U26495 (N_26495,N_25564,N_25968);
nor U26496 (N_26496,N_25873,N_25750);
xnor U26497 (N_26497,N_25528,N_25624);
xor U26498 (N_26498,N_25662,N_25773);
or U26499 (N_26499,N_25863,N_25593);
nor U26500 (N_26500,N_26293,N_26169);
and U26501 (N_26501,N_26070,N_26115);
nand U26502 (N_26502,N_26244,N_26069);
xnor U26503 (N_26503,N_26073,N_26288);
and U26504 (N_26504,N_26160,N_26272);
and U26505 (N_26505,N_26313,N_26162);
or U26506 (N_26506,N_26155,N_26248);
xnor U26507 (N_26507,N_26096,N_26241);
or U26508 (N_26508,N_26078,N_26226);
or U26509 (N_26509,N_26132,N_26268);
xnor U26510 (N_26510,N_26189,N_26403);
nand U26511 (N_26511,N_26441,N_26215);
nor U26512 (N_26512,N_26320,N_26006);
or U26513 (N_26513,N_26233,N_26323);
or U26514 (N_26514,N_26190,N_26458);
nand U26515 (N_26515,N_26135,N_26174);
xor U26516 (N_26516,N_26001,N_26129);
and U26517 (N_26517,N_26271,N_26326);
or U26518 (N_26518,N_26407,N_26220);
nand U26519 (N_26519,N_26305,N_26142);
xor U26520 (N_26520,N_26402,N_26116);
or U26521 (N_26521,N_26059,N_26036);
and U26522 (N_26522,N_26089,N_26154);
or U26523 (N_26523,N_26422,N_26367);
or U26524 (N_26524,N_26348,N_26037);
nor U26525 (N_26525,N_26076,N_26253);
and U26526 (N_26526,N_26490,N_26273);
or U26527 (N_26527,N_26020,N_26491);
nand U26528 (N_26528,N_26282,N_26083);
nor U26529 (N_26529,N_26062,N_26318);
nor U26530 (N_26530,N_26368,N_26229);
nor U26531 (N_26531,N_26114,N_26209);
nand U26532 (N_26532,N_26093,N_26499);
nand U26533 (N_26533,N_26476,N_26383);
nor U26534 (N_26534,N_26104,N_26193);
nand U26535 (N_26535,N_26284,N_26445);
and U26536 (N_26536,N_26287,N_26084);
nor U26537 (N_26537,N_26346,N_26314);
and U26538 (N_26538,N_26315,N_26025);
and U26539 (N_26539,N_26497,N_26300);
nor U26540 (N_26540,N_26296,N_26342);
xnor U26541 (N_26541,N_26124,N_26033);
and U26542 (N_26542,N_26003,N_26400);
nor U26543 (N_26543,N_26294,N_26390);
or U26544 (N_26544,N_26236,N_26055);
xor U26545 (N_26545,N_26477,N_26240);
and U26546 (N_26546,N_26332,N_26480);
or U26547 (N_26547,N_26417,N_26136);
xnor U26548 (N_26548,N_26245,N_26186);
xnor U26549 (N_26549,N_26385,N_26043);
or U26550 (N_26550,N_26275,N_26382);
nand U26551 (N_26551,N_26004,N_26398);
or U26552 (N_26552,N_26450,N_26176);
xor U26553 (N_26553,N_26427,N_26374);
and U26554 (N_26554,N_26375,N_26331);
nor U26555 (N_26555,N_26128,N_26479);
and U26556 (N_26556,N_26340,N_26231);
and U26557 (N_26557,N_26052,N_26266);
nor U26558 (N_26558,N_26466,N_26111);
xor U26559 (N_26559,N_26172,N_26386);
xor U26560 (N_26560,N_26097,N_26144);
and U26561 (N_26561,N_26291,N_26322);
xnor U26562 (N_26562,N_26079,N_26222);
nor U26563 (N_26563,N_26436,N_26380);
or U26564 (N_26564,N_26038,N_26041);
nand U26565 (N_26565,N_26311,N_26462);
nor U26566 (N_26566,N_26100,N_26184);
or U26567 (N_26567,N_26121,N_26484);
nand U26568 (N_26568,N_26179,N_26065);
or U26569 (N_26569,N_26439,N_26112);
or U26570 (N_26570,N_26212,N_26373);
nor U26571 (N_26571,N_26355,N_26103);
or U26572 (N_26572,N_26123,N_26082);
and U26573 (N_26573,N_26015,N_26219);
nor U26574 (N_26574,N_26406,N_26396);
or U26575 (N_26575,N_26306,N_26042);
and U26576 (N_26576,N_26252,N_26304);
nor U26577 (N_26577,N_26013,N_26347);
nand U26578 (N_26578,N_26310,N_26363);
and U26579 (N_26579,N_26276,N_26081);
xor U26580 (N_26580,N_26295,N_26392);
or U26581 (N_26581,N_26428,N_26464);
or U26582 (N_26582,N_26443,N_26388);
xnor U26583 (N_26583,N_26319,N_26005);
or U26584 (N_26584,N_26451,N_26000);
xnor U26585 (N_26585,N_26164,N_26026);
nand U26586 (N_26586,N_26357,N_26196);
nor U26587 (N_26587,N_26493,N_26178);
or U26588 (N_26588,N_26413,N_26071);
nand U26589 (N_26589,N_26438,N_26447);
xor U26590 (N_26590,N_26411,N_26085);
or U26591 (N_26591,N_26453,N_26281);
nor U26592 (N_26592,N_26011,N_26257);
nor U26593 (N_26593,N_26418,N_26452);
or U26594 (N_26594,N_26370,N_26412);
and U26595 (N_26595,N_26214,N_26246);
or U26596 (N_26596,N_26143,N_26335);
xor U26597 (N_26597,N_26454,N_26165);
nand U26598 (N_26598,N_26475,N_26469);
nand U26599 (N_26599,N_26200,N_26211);
nor U26600 (N_26600,N_26008,N_26007);
nor U26601 (N_26601,N_26095,N_26456);
and U26602 (N_26602,N_26470,N_26182);
or U26603 (N_26603,N_26039,N_26031);
and U26604 (N_26604,N_26146,N_26205);
xnor U26605 (N_26605,N_26194,N_26343);
nor U26606 (N_26606,N_26433,N_26399);
nand U26607 (N_26607,N_26105,N_26106);
and U26608 (N_26608,N_26483,N_26175);
xnor U26609 (N_26609,N_26309,N_26389);
or U26610 (N_26610,N_26101,N_26159);
or U26611 (N_26611,N_26199,N_26267);
nor U26612 (N_26612,N_26122,N_26012);
nor U26613 (N_26613,N_26045,N_26047);
xnor U26614 (N_26614,N_26364,N_26247);
nor U26615 (N_26615,N_26325,N_26242);
nor U26616 (N_26616,N_26298,N_26206);
or U26617 (N_26617,N_26393,N_26459);
xor U26618 (N_26618,N_26152,N_26110);
and U26619 (N_26619,N_26127,N_26051);
xnor U26620 (N_26620,N_26192,N_26430);
xnor U26621 (N_26621,N_26170,N_26139);
nand U26622 (N_26622,N_26232,N_26197);
nand U26623 (N_26623,N_26260,N_26440);
nand U26624 (N_26624,N_26217,N_26496);
or U26625 (N_26625,N_26054,N_26077);
nor U26626 (N_26626,N_26297,N_26149);
nor U26627 (N_26627,N_26191,N_26088);
or U26628 (N_26628,N_26237,N_26337);
and U26629 (N_26629,N_26307,N_26181);
xor U26630 (N_26630,N_26140,N_26249);
nand U26631 (N_26631,N_26158,N_26460);
xnor U26632 (N_26632,N_26218,N_26327);
nor U26633 (N_26633,N_26448,N_26317);
nor U26634 (N_26634,N_26435,N_26032);
nor U26635 (N_26635,N_26415,N_26457);
nand U26636 (N_26636,N_26075,N_26256);
nand U26637 (N_26637,N_26414,N_26423);
and U26638 (N_26638,N_26324,N_26285);
or U26639 (N_26639,N_26362,N_26163);
nand U26640 (N_26640,N_26254,N_26431);
nor U26641 (N_26641,N_26177,N_26372);
nor U26642 (N_26642,N_26377,N_26424);
nand U26643 (N_26643,N_26056,N_26487);
nor U26644 (N_26644,N_26265,N_26471);
or U26645 (N_26645,N_26345,N_26488);
nor U26646 (N_26646,N_26329,N_26405);
xor U26647 (N_26647,N_26094,N_26230);
and U26648 (N_26648,N_26404,N_26384);
and U26649 (N_26649,N_26019,N_26328);
nand U26650 (N_26650,N_26336,N_26022);
xor U26651 (N_26651,N_26481,N_26270);
xor U26652 (N_26652,N_26072,N_26017);
or U26653 (N_26653,N_26040,N_26303);
nand U26654 (N_26654,N_26126,N_26473);
or U26655 (N_26655,N_26207,N_26187);
xnor U26656 (N_26656,N_26108,N_26419);
or U26657 (N_26657,N_26210,N_26202);
xor U26658 (N_26658,N_26301,N_26223);
xnor U26659 (N_26659,N_26489,N_26379);
or U26660 (N_26660,N_26361,N_26283);
xor U26661 (N_26661,N_26213,N_26321);
or U26662 (N_26662,N_26153,N_26359);
nor U26663 (N_26663,N_26118,N_26201);
nand U26664 (N_26664,N_26173,N_26014);
and U26665 (N_26665,N_26058,N_26208);
nand U26666 (N_26666,N_26482,N_26203);
nand U26667 (N_26667,N_26030,N_26290);
nand U26668 (N_26668,N_26002,N_26292);
or U26669 (N_26669,N_26274,N_26060);
xnor U26670 (N_26670,N_26048,N_26034);
nor U26671 (N_26671,N_26109,N_26349);
xnor U26672 (N_26672,N_26333,N_26107);
and U26673 (N_26673,N_26063,N_26369);
xnor U26674 (N_26674,N_26408,N_26134);
nor U26675 (N_26675,N_26024,N_26302);
nor U26676 (N_26676,N_26010,N_26099);
nand U26677 (N_26677,N_26120,N_26061);
and U26678 (N_26678,N_26044,N_26133);
nor U26679 (N_26679,N_26027,N_26092);
or U26680 (N_26680,N_26365,N_26442);
and U26681 (N_26681,N_26351,N_26021);
xnor U26682 (N_26682,N_26049,N_26366);
nor U26683 (N_26683,N_26494,N_26474);
nand U26684 (N_26684,N_26156,N_26086);
or U26685 (N_26685,N_26279,N_26278);
and U26686 (N_26686,N_26350,N_26147);
and U26687 (N_26687,N_26145,N_26131);
nor U26688 (N_26688,N_26125,N_26018);
xnor U26689 (N_26689,N_26468,N_26251);
and U26690 (N_26690,N_26360,N_26148);
xor U26691 (N_26691,N_26113,N_26334);
and U26692 (N_26692,N_26437,N_26394);
nand U26693 (N_26693,N_26050,N_26035);
nand U26694 (N_26694,N_26016,N_26185);
or U26695 (N_26695,N_26353,N_26472);
nor U26696 (N_26696,N_26498,N_26028);
xnor U26697 (N_26697,N_26261,N_26316);
or U26698 (N_26698,N_26397,N_26239);
and U26699 (N_26699,N_26409,N_26102);
xor U26700 (N_26700,N_26280,N_26166);
nand U26701 (N_26701,N_26444,N_26066);
nand U26702 (N_26702,N_26264,N_26358);
nand U26703 (N_26703,N_26312,N_26255);
or U26704 (N_26704,N_26074,N_26461);
and U26705 (N_26705,N_26080,N_26150);
or U26706 (N_26706,N_26426,N_26420);
and U26707 (N_26707,N_26371,N_26161);
xnor U26708 (N_26708,N_26262,N_26098);
xnor U26709 (N_26709,N_26425,N_26141);
or U26710 (N_26710,N_26263,N_26151);
and U26711 (N_26711,N_26180,N_26221);
nor U26712 (N_26712,N_26167,N_26168);
or U26713 (N_26713,N_26429,N_26455);
and U26714 (N_26714,N_26486,N_26250);
xor U26715 (N_26715,N_26238,N_26376);
xor U26716 (N_26716,N_26090,N_26068);
xnor U26717 (N_26717,N_26138,N_26198);
and U26718 (N_26718,N_26204,N_26228);
and U26719 (N_26719,N_26119,N_26053);
xnor U26720 (N_26720,N_26216,N_26188);
and U26721 (N_26721,N_26378,N_26277);
and U26722 (N_26722,N_26449,N_26354);
nand U26723 (N_26723,N_26338,N_26225);
nor U26724 (N_26724,N_26344,N_26243);
nand U26725 (N_26725,N_26421,N_26286);
nand U26726 (N_26726,N_26416,N_26387);
nand U26727 (N_26727,N_26463,N_26356);
or U26728 (N_26728,N_26046,N_26395);
nand U26729 (N_26729,N_26183,N_26432);
nor U26730 (N_26730,N_26485,N_26299);
nor U26731 (N_26731,N_26308,N_26330);
nand U26732 (N_26732,N_26171,N_26401);
and U26733 (N_26733,N_26434,N_26091);
nand U26734 (N_26734,N_26067,N_26381);
and U26735 (N_26735,N_26391,N_26064);
and U26736 (N_26736,N_26492,N_26057);
nand U26737 (N_26737,N_26341,N_26465);
xor U26738 (N_26738,N_26410,N_26157);
and U26739 (N_26739,N_26446,N_26227);
xor U26740 (N_26740,N_26339,N_26087);
and U26741 (N_26741,N_26130,N_26029);
and U26742 (N_26742,N_26258,N_26195);
and U26743 (N_26743,N_26137,N_26259);
xor U26744 (N_26744,N_26289,N_26009);
xor U26745 (N_26745,N_26023,N_26352);
or U26746 (N_26746,N_26224,N_26478);
xor U26747 (N_26747,N_26235,N_26117);
and U26748 (N_26748,N_26269,N_26495);
and U26749 (N_26749,N_26467,N_26234);
xnor U26750 (N_26750,N_26294,N_26451);
xnor U26751 (N_26751,N_26078,N_26181);
or U26752 (N_26752,N_26277,N_26372);
nand U26753 (N_26753,N_26323,N_26293);
nand U26754 (N_26754,N_26405,N_26038);
nor U26755 (N_26755,N_26341,N_26321);
xnor U26756 (N_26756,N_26119,N_26186);
nor U26757 (N_26757,N_26261,N_26396);
nor U26758 (N_26758,N_26192,N_26132);
and U26759 (N_26759,N_26259,N_26316);
nor U26760 (N_26760,N_26406,N_26487);
xor U26761 (N_26761,N_26346,N_26467);
xor U26762 (N_26762,N_26030,N_26207);
xor U26763 (N_26763,N_26295,N_26133);
xnor U26764 (N_26764,N_26055,N_26121);
and U26765 (N_26765,N_26181,N_26271);
nand U26766 (N_26766,N_26366,N_26224);
xor U26767 (N_26767,N_26246,N_26097);
nor U26768 (N_26768,N_26259,N_26432);
and U26769 (N_26769,N_26410,N_26310);
nor U26770 (N_26770,N_26168,N_26129);
xor U26771 (N_26771,N_26142,N_26313);
nand U26772 (N_26772,N_26177,N_26292);
or U26773 (N_26773,N_26056,N_26163);
and U26774 (N_26774,N_26292,N_26286);
or U26775 (N_26775,N_26279,N_26319);
and U26776 (N_26776,N_26019,N_26464);
nand U26777 (N_26777,N_26182,N_26164);
nand U26778 (N_26778,N_26112,N_26435);
nor U26779 (N_26779,N_26195,N_26055);
nor U26780 (N_26780,N_26044,N_26092);
and U26781 (N_26781,N_26031,N_26428);
and U26782 (N_26782,N_26417,N_26014);
nand U26783 (N_26783,N_26118,N_26176);
nand U26784 (N_26784,N_26231,N_26188);
xor U26785 (N_26785,N_26042,N_26017);
and U26786 (N_26786,N_26284,N_26003);
nor U26787 (N_26787,N_26135,N_26397);
or U26788 (N_26788,N_26118,N_26014);
xnor U26789 (N_26789,N_26072,N_26268);
and U26790 (N_26790,N_26147,N_26273);
xnor U26791 (N_26791,N_26189,N_26181);
and U26792 (N_26792,N_26229,N_26390);
and U26793 (N_26793,N_26263,N_26481);
nor U26794 (N_26794,N_26434,N_26210);
xor U26795 (N_26795,N_26084,N_26225);
nand U26796 (N_26796,N_26131,N_26449);
or U26797 (N_26797,N_26276,N_26466);
nor U26798 (N_26798,N_26493,N_26194);
or U26799 (N_26799,N_26082,N_26491);
nand U26800 (N_26800,N_26107,N_26271);
nor U26801 (N_26801,N_26310,N_26103);
nand U26802 (N_26802,N_26401,N_26178);
nand U26803 (N_26803,N_26157,N_26074);
xnor U26804 (N_26804,N_26331,N_26317);
and U26805 (N_26805,N_26230,N_26111);
nand U26806 (N_26806,N_26042,N_26087);
or U26807 (N_26807,N_26232,N_26042);
nand U26808 (N_26808,N_26485,N_26166);
xor U26809 (N_26809,N_26268,N_26338);
or U26810 (N_26810,N_26256,N_26469);
nand U26811 (N_26811,N_26234,N_26154);
or U26812 (N_26812,N_26224,N_26014);
or U26813 (N_26813,N_26136,N_26071);
and U26814 (N_26814,N_26138,N_26378);
nor U26815 (N_26815,N_26181,N_26485);
nand U26816 (N_26816,N_26072,N_26459);
or U26817 (N_26817,N_26070,N_26143);
xor U26818 (N_26818,N_26036,N_26318);
nand U26819 (N_26819,N_26345,N_26142);
xnor U26820 (N_26820,N_26199,N_26123);
nor U26821 (N_26821,N_26013,N_26401);
nor U26822 (N_26822,N_26438,N_26055);
nor U26823 (N_26823,N_26390,N_26177);
nand U26824 (N_26824,N_26180,N_26059);
xnor U26825 (N_26825,N_26091,N_26160);
and U26826 (N_26826,N_26422,N_26221);
nor U26827 (N_26827,N_26411,N_26100);
or U26828 (N_26828,N_26499,N_26121);
nor U26829 (N_26829,N_26429,N_26110);
xnor U26830 (N_26830,N_26301,N_26169);
nor U26831 (N_26831,N_26368,N_26376);
nand U26832 (N_26832,N_26257,N_26284);
nand U26833 (N_26833,N_26023,N_26119);
xor U26834 (N_26834,N_26397,N_26498);
nor U26835 (N_26835,N_26353,N_26477);
xnor U26836 (N_26836,N_26025,N_26376);
nand U26837 (N_26837,N_26323,N_26065);
xnor U26838 (N_26838,N_26222,N_26192);
nor U26839 (N_26839,N_26398,N_26175);
or U26840 (N_26840,N_26181,N_26041);
or U26841 (N_26841,N_26427,N_26370);
nand U26842 (N_26842,N_26134,N_26173);
and U26843 (N_26843,N_26095,N_26298);
nand U26844 (N_26844,N_26201,N_26274);
nand U26845 (N_26845,N_26235,N_26047);
nand U26846 (N_26846,N_26015,N_26378);
xnor U26847 (N_26847,N_26161,N_26313);
xnor U26848 (N_26848,N_26046,N_26397);
xor U26849 (N_26849,N_26338,N_26134);
nor U26850 (N_26850,N_26077,N_26280);
nor U26851 (N_26851,N_26393,N_26201);
nor U26852 (N_26852,N_26018,N_26460);
xnor U26853 (N_26853,N_26116,N_26127);
nor U26854 (N_26854,N_26433,N_26194);
or U26855 (N_26855,N_26336,N_26205);
nand U26856 (N_26856,N_26166,N_26263);
nand U26857 (N_26857,N_26089,N_26397);
nand U26858 (N_26858,N_26116,N_26381);
nand U26859 (N_26859,N_26228,N_26454);
xnor U26860 (N_26860,N_26460,N_26144);
and U26861 (N_26861,N_26454,N_26118);
or U26862 (N_26862,N_26188,N_26499);
and U26863 (N_26863,N_26128,N_26460);
xnor U26864 (N_26864,N_26303,N_26362);
nand U26865 (N_26865,N_26007,N_26431);
and U26866 (N_26866,N_26098,N_26139);
xnor U26867 (N_26867,N_26000,N_26063);
nor U26868 (N_26868,N_26466,N_26196);
and U26869 (N_26869,N_26157,N_26497);
xor U26870 (N_26870,N_26411,N_26279);
xnor U26871 (N_26871,N_26418,N_26029);
nand U26872 (N_26872,N_26223,N_26020);
xnor U26873 (N_26873,N_26230,N_26197);
xnor U26874 (N_26874,N_26128,N_26459);
and U26875 (N_26875,N_26209,N_26223);
nor U26876 (N_26876,N_26113,N_26258);
or U26877 (N_26877,N_26249,N_26133);
xor U26878 (N_26878,N_26122,N_26298);
and U26879 (N_26879,N_26102,N_26325);
or U26880 (N_26880,N_26248,N_26225);
xor U26881 (N_26881,N_26404,N_26147);
xnor U26882 (N_26882,N_26415,N_26418);
xnor U26883 (N_26883,N_26164,N_26086);
nor U26884 (N_26884,N_26363,N_26178);
and U26885 (N_26885,N_26250,N_26118);
nand U26886 (N_26886,N_26362,N_26078);
xor U26887 (N_26887,N_26278,N_26422);
nor U26888 (N_26888,N_26285,N_26441);
and U26889 (N_26889,N_26110,N_26043);
or U26890 (N_26890,N_26465,N_26405);
nand U26891 (N_26891,N_26094,N_26155);
nand U26892 (N_26892,N_26414,N_26367);
nor U26893 (N_26893,N_26109,N_26388);
nand U26894 (N_26894,N_26291,N_26103);
xor U26895 (N_26895,N_26424,N_26390);
nor U26896 (N_26896,N_26089,N_26437);
or U26897 (N_26897,N_26087,N_26390);
and U26898 (N_26898,N_26289,N_26430);
or U26899 (N_26899,N_26240,N_26281);
nor U26900 (N_26900,N_26126,N_26199);
xnor U26901 (N_26901,N_26059,N_26019);
nor U26902 (N_26902,N_26460,N_26084);
or U26903 (N_26903,N_26066,N_26068);
or U26904 (N_26904,N_26201,N_26442);
and U26905 (N_26905,N_26409,N_26064);
nor U26906 (N_26906,N_26153,N_26130);
nor U26907 (N_26907,N_26482,N_26451);
and U26908 (N_26908,N_26302,N_26432);
nor U26909 (N_26909,N_26476,N_26140);
nor U26910 (N_26910,N_26121,N_26043);
or U26911 (N_26911,N_26222,N_26116);
or U26912 (N_26912,N_26447,N_26289);
and U26913 (N_26913,N_26375,N_26403);
or U26914 (N_26914,N_26321,N_26276);
nand U26915 (N_26915,N_26071,N_26135);
xnor U26916 (N_26916,N_26376,N_26433);
xor U26917 (N_26917,N_26393,N_26142);
xor U26918 (N_26918,N_26046,N_26137);
or U26919 (N_26919,N_26308,N_26297);
or U26920 (N_26920,N_26200,N_26371);
nor U26921 (N_26921,N_26220,N_26041);
xor U26922 (N_26922,N_26332,N_26072);
nand U26923 (N_26923,N_26249,N_26230);
or U26924 (N_26924,N_26057,N_26131);
nor U26925 (N_26925,N_26423,N_26218);
xnor U26926 (N_26926,N_26112,N_26017);
or U26927 (N_26927,N_26122,N_26025);
xor U26928 (N_26928,N_26040,N_26406);
or U26929 (N_26929,N_26131,N_26420);
nand U26930 (N_26930,N_26396,N_26053);
and U26931 (N_26931,N_26230,N_26142);
nor U26932 (N_26932,N_26013,N_26118);
xnor U26933 (N_26933,N_26367,N_26418);
and U26934 (N_26934,N_26497,N_26451);
or U26935 (N_26935,N_26465,N_26468);
or U26936 (N_26936,N_26358,N_26036);
and U26937 (N_26937,N_26258,N_26265);
or U26938 (N_26938,N_26155,N_26047);
or U26939 (N_26939,N_26234,N_26087);
nor U26940 (N_26940,N_26368,N_26289);
xnor U26941 (N_26941,N_26143,N_26003);
nor U26942 (N_26942,N_26129,N_26480);
nor U26943 (N_26943,N_26412,N_26439);
or U26944 (N_26944,N_26154,N_26180);
nand U26945 (N_26945,N_26291,N_26205);
or U26946 (N_26946,N_26299,N_26266);
and U26947 (N_26947,N_26011,N_26119);
xnor U26948 (N_26948,N_26461,N_26062);
or U26949 (N_26949,N_26465,N_26328);
or U26950 (N_26950,N_26102,N_26481);
nor U26951 (N_26951,N_26179,N_26243);
nor U26952 (N_26952,N_26155,N_26070);
xor U26953 (N_26953,N_26375,N_26053);
nor U26954 (N_26954,N_26277,N_26131);
nor U26955 (N_26955,N_26361,N_26428);
nand U26956 (N_26956,N_26217,N_26115);
xor U26957 (N_26957,N_26300,N_26101);
nor U26958 (N_26958,N_26193,N_26095);
or U26959 (N_26959,N_26284,N_26036);
and U26960 (N_26960,N_26386,N_26396);
nand U26961 (N_26961,N_26006,N_26340);
nand U26962 (N_26962,N_26342,N_26469);
and U26963 (N_26963,N_26114,N_26025);
nor U26964 (N_26964,N_26495,N_26182);
nand U26965 (N_26965,N_26227,N_26257);
and U26966 (N_26966,N_26324,N_26416);
nor U26967 (N_26967,N_26456,N_26228);
or U26968 (N_26968,N_26420,N_26031);
nor U26969 (N_26969,N_26322,N_26257);
nand U26970 (N_26970,N_26268,N_26067);
xnor U26971 (N_26971,N_26369,N_26084);
nand U26972 (N_26972,N_26368,N_26137);
nor U26973 (N_26973,N_26337,N_26472);
nor U26974 (N_26974,N_26061,N_26324);
nor U26975 (N_26975,N_26029,N_26181);
or U26976 (N_26976,N_26465,N_26422);
nor U26977 (N_26977,N_26209,N_26145);
or U26978 (N_26978,N_26118,N_26215);
nor U26979 (N_26979,N_26099,N_26108);
or U26980 (N_26980,N_26325,N_26290);
or U26981 (N_26981,N_26096,N_26295);
nand U26982 (N_26982,N_26299,N_26252);
nand U26983 (N_26983,N_26450,N_26442);
and U26984 (N_26984,N_26205,N_26207);
and U26985 (N_26985,N_26242,N_26393);
nor U26986 (N_26986,N_26176,N_26401);
or U26987 (N_26987,N_26161,N_26014);
and U26988 (N_26988,N_26235,N_26318);
nand U26989 (N_26989,N_26481,N_26196);
nand U26990 (N_26990,N_26064,N_26230);
xor U26991 (N_26991,N_26327,N_26421);
or U26992 (N_26992,N_26389,N_26316);
xnor U26993 (N_26993,N_26280,N_26003);
nand U26994 (N_26994,N_26116,N_26434);
or U26995 (N_26995,N_26140,N_26231);
and U26996 (N_26996,N_26216,N_26304);
or U26997 (N_26997,N_26130,N_26497);
xnor U26998 (N_26998,N_26101,N_26037);
xnor U26999 (N_26999,N_26019,N_26007);
nor U27000 (N_27000,N_26584,N_26949);
and U27001 (N_27001,N_26844,N_26527);
nand U27002 (N_27002,N_26580,N_26583);
and U27003 (N_27003,N_26916,N_26587);
nand U27004 (N_27004,N_26504,N_26694);
and U27005 (N_27005,N_26698,N_26720);
xnor U27006 (N_27006,N_26511,N_26625);
nor U27007 (N_27007,N_26843,N_26830);
nand U27008 (N_27008,N_26598,N_26836);
nand U27009 (N_27009,N_26876,N_26682);
xor U27010 (N_27010,N_26701,N_26899);
nor U27011 (N_27011,N_26523,N_26961);
and U27012 (N_27012,N_26880,N_26744);
or U27013 (N_27013,N_26968,N_26706);
nand U27014 (N_27014,N_26870,N_26767);
or U27015 (N_27015,N_26940,N_26660);
nor U27016 (N_27016,N_26631,N_26762);
xnor U27017 (N_27017,N_26704,N_26909);
and U27018 (N_27018,N_26615,N_26972);
or U27019 (N_27019,N_26683,N_26600);
nand U27020 (N_27020,N_26951,N_26655);
and U27021 (N_27021,N_26853,N_26567);
xnor U27022 (N_27022,N_26936,N_26632);
or U27023 (N_27023,N_26877,N_26654);
and U27024 (N_27024,N_26576,N_26715);
xnor U27025 (N_27025,N_26597,N_26620);
xor U27026 (N_27026,N_26593,N_26651);
or U27027 (N_27027,N_26835,N_26540);
or U27028 (N_27028,N_26652,N_26556);
nor U27029 (N_27029,N_26667,N_26759);
nand U27030 (N_27030,N_26933,N_26994);
or U27031 (N_27031,N_26713,N_26719);
or U27032 (N_27032,N_26924,N_26891);
and U27033 (N_27033,N_26849,N_26524);
nand U27034 (N_27034,N_26781,N_26714);
xor U27035 (N_27035,N_26825,N_26648);
xnor U27036 (N_27036,N_26914,N_26551);
and U27037 (N_27037,N_26791,N_26507);
xnor U27038 (N_27038,N_26862,N_26750);
nor U27039 (N_27039,N_26954,N_26989);
or U27040 (N_27040,N_26579,N_26599);
nand U27041 (N_27041,N_26596,N_26778);
and U27042 (N_27042,N_26866,N_26903);
nand U27043 (N_27043,N_26570,N_26971);
xor U27044 (N_27044,N_26976,N_26578);
nor U27045 (N_27045,N_26585,N_26549);
nor U27046 (N_27046,N_26553,N_26889);
nand U27047 (N_27047,N_26646,N_26979);
and U27048 (N_27048,N_26610,N_26887);
xor U27049 (N_27049,N_26595,N_26860);
or U27050 (N_27050,N_26550,N_26911);
xnor U27051 (N_27051,N_26942,N_26670);
nand U27052 (N_27052,N_26733,N_26734);
nand U27053 (N_27053,N_26624,N_26780);
or U27054 (N_27054,N_26514,N_26582);
or U27055 (N_27055,N_26673,N_26766);
nor U27056 (N_27056,N_26884,N_26619);
and U27057 (N_27057,N_26503,N_26737);
or U27058 (N_27058,N_26752,N_26741);
nor U27059 (N_27059,N_26947,N_26749);
nand U27060 (N_27060,N_26806,N_26970);
nand U27061 (N_27061,N_26832,N_26879);
and U27062 (N_27062,N_26533,N_26642);
and U27063 (N_27063,N_26787,N_26952);
or U27064 (N_27064,N_26622,N_26618);
or U27065 (N_27065,N_26802,N_26756);
xnor U27066 (N_27066,N_26816,N_26690);
xnor U27067 (N_27067,N_26929,N_26941);
nand U27068 (N_27068,N_26569,N_26501);
and U27069 (N_27069,N_26639,N_26902);
nand U27070 (N_27070,N_26526,N_26939);
xnor U27071 (N_27071,N_26831,N_26775);
nor U27072 (N_27072,N_26725,N_26606);
xor U27073 (N_27073,N_26882,N_26895);
and U27074 (N_27074,N_26907,N_26681);
nor U27075 (N_27075,N_26934,N_26539);
nand U27076 (N_27076,N_26537,N_26998);
and U27077 (N_27077,N_26819,N_26510);
nor U27078 (N_27078,N_26638,N_26592);
or U27079 (N_27079,N_26705,N_26804);
or U27080 (N_27080,N_26529,N_26918);
and U27081 (N_27081,N_26894,N_26983);
xor U27082 (N_27082,N_26643,N_26717);
xor U27083 (N_27083,N_26740,N_26702);
and U27084 (N_27084,N_26708,N_26530);
nand U27085 (N_27085,N_26852,N_26845);
nor U27086 (N_27086,N_26685,N_26707);
or U27087 (N_27087,N_26535,N_26855);
or U27088 (N_27088,N_26793,N_26957);
xnor U27089 (N_27089,N_26566,N_26938);
and U27090 (N_27090,N_26532,N_26926);
xnor U27091 (N_27091,N_26962,N_26856);
or U27092 (N_27092,N_26621,N_26921);
xor U27093 (N_27093,N_26857,N_26736);
nand U27094 (N_27094,N_26869,N_26650);
nor U27095 (N_27095,N_26603,N_26950);
and U27096 (N_27096,N_26789,N_26878);
nor U27097 (N_27097,N_26888,N_26742);
nor U27098 (N_27098,N_26575,N_26945);
or U27099 (N_27099,N_26900,N_26997);
nand U27100 (N_27100,N_26847,N_26958);
nand U27101 (N_27101,N_26594,N_26564);
nand U27102 (N_27102,N_26520,N_26788);
nand U27103 (N_27103,N_26657,N_26671);
nor U27104 (N_27104,N_26956,N_26565);
nor U27105 (N_27105,N_26774,N_26798);
nand U27106 (N_27106,N_26935,N_26827);
or U27107 (N_27107,N_26906,N_26810);
nand U27108 (N_27108,N_26771,N_26867);
or U27109 (N_27109,N_26712,N_26699);
nand U27110 (N_27110,N_26839,N_26991);
nand U27111 (N_27111,N_26677,N_26851);
xnor U27112 (N_27112,N_26966,N_26848);
nand U27113 (N_27113,N_26754,N_26908);
xnor U27114 (N_27114,N_26591,N_26777);
and U27115 (N_27115,N_26653,N_26769);
nor U27116 (N_27116,N_26546,N_26666);
nand U27117 (N_27117,N_26915,N_26512);
or U27118 (N_27118,N_26534,N_26863);
nand U27119 (N_27119,N_26659,N_26502);
nor U27120 (N_27120,N_26703,N_26809);
or U27121 (N_27121,N_26992,N_26568);
or U27122 (N_27122,N_26732,N_26829);
nand U27123 (N_27123,N_26723,N_26745);
xnor U27124 (N_27124,N_26913,N_26974);
xnor U27125 (N_27125,N_26692,N_26892);
and U27126 (N_27126,N_26996,N_26927);
nor U27127 (N_27127,N_26676,N_26663);
nor U27128 (N_27128,N_26628,N_26896);
and U27129 (N_27129,N_26883,N_26764);
xor U27130 (N_27130,N_26963,N_26710);
or U27131 (N_27131,N_26881,N_26922);
xnor U27132 (N_27132,N_26519,N_26544);
and U27133 (N_27133,N_26917,N_26633);
nand U27134 (N_27134,N_26981,N_26897);
xor U27135 (N_27135,N_26912,N_26545);
or U27136 (N_27136,N_26795,N_26684);
nand U27137 (N_27137,N_26668,N_26875);
nor U27138 (N_27138,N_26617,N_26800);
or U27139 (N_27139,N_26727,N_26796);
or U27140 (N_27140,N_26817,N_26687);
nand U27141 (N_27141,N_26589,N_26538);
and U27142 (N_27142,N_26525,N_26528);
nand U27143 (N_27143,N_26611,N_26604);
nor U27144 (N_27144,N_26608,N_26978);
and U27145 (N_27145,N_26850,N_26794);
nand U27146 (N_27146,N_26944,N_26842);
nand U27147 (N_27147,N_26662,N_26728);
nand U27148 (N_27148,N_26818,N_26669);
nand U27149 (N_27149,N_26772,N_26932);
or U27150 (N_27150,N_26885,N_26811);
and U27151 (N_27151,N_26557,N_26577);
xnor U27152 (N_27152,N_26973,N_26581);
or U27153 (N_27153,N_26661,N_26815);
or U27154 (N_27154,N_26999,N_26697);
xor U27155 (N_27155,N_26572,N_26531);
or U27156 (N_27156,N_26548,N_26980);
nor U27157 (N_27157,N_26872,N_26623);
nand U27158 (N_27158,N_26588,N_26834);
and U27159 (N_27159,N_26898,N_26672);
xor U27160 (N_27160,N_26751,N_26873);
xor U27161 (N_27161,N_26985,N_26874);
or U27162 (N_27162,N_26782,N_26695);
or U27163 (N_27163,N_26964,N_26814);
and U27164 (N_27164,N_26828,N_26923);
nor U27165 (N_27165,N_26743,N_26637);
nand U27166 (N_27166,N_26559,N_26858);
and U27167 (N_27167,N_26987,N_26679);
xnor U27168 (N_27168,N_26641,N_26688);
xor U27169 (N_27169,N_26574,N_26689);
or U27170 (N_27170,N_26948,N_26506);
or U27171 (N_27171,N_26516,N_26861);
or U27172 (N_27172,N_26770,N_26813);
nand U27173 (N_27173,N_26634,N_26711);
or U27174 (N_27174,N_26807,N_26910);
or U27175 (N_27175,N_26696,N_26627);
or U27176 (N_27176,N_26930,N_26645);
xor U27177 (N_27177,N_26724,N_26748);
or U27178 (N_27178,N_26757,N_26602);
or U27179 (N_27179,N_26840,N_26630);
and U27180 (N_27180,N_26808,N_26718);
and U27181 (N_27181,N_26776,N_26833);
or U27182 (N_27182,N_26821,N_26773);
nor U27183 (N_27183,N_26854,N_26784);
nor U27184 (N_27184,N_26955,N_26865);
nor U27185 (N_27185,N_26613,N_26629);
nor U27186 (N_27186,N_26636,N_26779);
xor U27187 (N_27187,N_26904,N_26605);
nand U27188 (N_27188,N_26920,N_26729);
nand U27189 (N_27189,N_26768,N_26590);
and U27190 (N_27190,N_26509,N_26561);
or U27191 (N_27191,N_26508,N_26612);
or U27192 (N_27192,N_26763,N_26977);
or U27193 (N_27193,N_26799,N_26601);
nand U27194 (N_27194,N_26990,N_26626);
and U27195 (N_27195,N_26986,N_26571);
nor U27196 (N_27196,N_26931,N_26988);
and U27197 (N_27197,N_26901,N_26747);
nand U27198 (N_27198,N_26893,N_26649);
nor U27199 (N_27199,N_26755,N_26726);
nor U27200 (N_27200,N_26890,N_26993);
nand U27201 (N_27201,N_26792,N_26586);
nor U27202 (N_27202,N_26868,N_26846);
xor U27203 (N_27203,N_26607,N_26691);
and U27204 (N_27204,N_26946,N_26925);
nor U27205 (N_27205,N_26678,N_26758);
nor U27206 (N_27206,N_26919,N_26826);
nand U27207 (N_27207,N_26822,N_26555);
nand U27208 (N_27208,N_26656,N_26969);
and U27209 (N_27209,N_26790,N_26943);
nand U27210 (N_27210,N_26665,N_26563);
and U27211 (N_27211,N_26554,N_26616);
or U27212 (N_27212,N_26805,N_26693);
nand U27213 (N_27213,N_26675,N_26841);
xnor U27214 (N_27214,N_26786,N_26735);
or U27215 (N_27215,N_26838,N_26647);
nor U27216 (N_27216,N_26765,N_26500);
or U27217 (N_27217,N_26560,N_26982);
xor U27218 (N_27218,N_26552,N_26761);
nand U27219 (N_27219,N_26812,N_26716);
nand U27220 (N_27220,N_26536,N_26515);
xor U27221 (N_27221,N_26753,N_26797);
nor U27222 (N_27222,N_26824,N_26558);
nor U27223 (N_27223,N_26658,N_26859);
and U27224 (N_27224,N_26886,N_26543);
nand U27225 (N_27225,N_26995,N_26785);
xor U27226 (N_27226,N_26739,N_26928);
and U27227 (N_27227,N_26871,N_26521);
xnor U27228 (N_27228,N_26542,N_26905);
or U27229 (N_27229,N_26562,N_26746);
nor U27230 (N_27230,N_26820,N_26573);
nand U27231 (N_27231,N_26823,N_26803);
nand U27232 (N_27232,N_26975,N_26721);
xnor U27233 (N_27233,N_26522,N_26801);
or U27234 (N_27234,N_26738,N_26635);
xnor U27235 (N_27235,N_26686,N_26664);
nor U27236 (N_27236,N_26513,N_26614);
nor U27237 (N_27237,N_26644,N_26864);
and U27238 (N_27238,N_26783,N_26837);
nand U27239 (N_27239,N_26640,N_26731);
and U27240 (N_27240,N_26760,N_26984);
nand U27241 (N_27241,N_26674,N_26953);
nor U27242 (N_27242,N_26967,N_26937);
nor U27243 (N_27243,N_26959,N_26609);
nand U27244 (N_27244,N_26680,N_26518);
nor U27245 (N_27245,N_26505,N_26965);
xor U27246 (N_27246,N_26722,N_26700);
and U27247 (N_27247,N_26709,N_26547);
nor U27248 (N_27248,N_26960,N_26541);
and U27249 (N_27249,N_26517,N_26730);
nor U27250 (N_27250,N_26907,N_26875);
and U27251 (N_27251,N_26546,N_26661);
and U27252 (N_27252,N_26686,N_26614);
and U27253 (N_27253,N_26739,N_26769);
and U27254 (N_27254,N_26566,N_26997);
nor U27255 (N_27255,N_26849,N_26723);
nor U27256 (N_27256,N_26728,N_26918);
nand U27257 (N_27257,N_26856,N_26968);
or U27258 (N_27258,N_26538,N_26679);
and U27259 (N_27259,N_26590,N_26917);
nor U27260 (N_27260,N_26900,N_26993);
xnor U27261 (N_27261,N_26751,N_26810);
nand U27262 (N_27262,N_26575,N_26983);
and U27263 (N_27263,N_26792,N_26734);
nor U27264 (N_27264,N_26709,N_26746);
xor U27265 (N_27265,N_26597,N_26546);
xnor U27266 (N_27266,N_26529,N_26555);
nand U27267 (N_27267,N_26957,N_26608);
nor U27268 (N_27268,N_26668,N_26994);
xnor U27269 (N_27269,N_26894,N_26834);
nand U27270 (N_27270,N_26975,N_26614);
or U27271 (N_27271,N_26515,N_26600);
or U27272 (N_27272,N_26759,N_26569);
or U27273 (N_27273,N_26682,N_26880);
nor U27274 (N_27274,N_26721,N_26723);
xor U27275 (N_27275,N_26943,N_26734);
nor U27276 (N_27276,N_26681,N_26632);
nand U27277 (N_27277,N_26927,N_26783);
nand U27278 (N_27278,N_26892,N_26632);
and U27279 (N_27279,N_26667,N_26869);
xor U27280 (N_27280,N_26797,N_26776);
xnor U27281 (N_27281,N_26614,N_26619);
nor U27282 (N_27282,N_26855,N_26596);
nand U27283 (N_27283,N_26896,N_26953);
and U27284 (N_27284,N_26934,N_26513);
and U27285 (N_27285,N_26771,N_26879);
nor U27286 (N_27286,N_26915,N_26954);
nand U27287 (N_27287,N_26508,N_26733);
nor U27288 (N_27288,N_26881,N_26993);
nand U27289 (N_27289,N_26791,N_26986);
nand U27290 (N_27290,N_26639,N_26855);
nor U27291 (N_27291,N_26614,N_26735);
nand U27292 (N_27292,N_26881,N_26508);
and U27293 (N_27293,N_26706,N_26978);
nor U27294 (N_27294,N_26750,N_26598);
xnor U27295 (N_27295,N_26751,N_26555);
xnor U27296 (N_27296,N_26855,N_26540);
nand U27297 (N_27297,N_26804,N_26723);
nand U27298 (N_27298,N_26971,N_26946);
and U27299 (N_27299,N_26791,N_26503);
xnor U27300 (N_27300,N_26530,N_26680);
and U27301 (N_27301,N_26769,N_26519);
and U27302 (N_27302,N_26966,N_26688);
and U27303 (N_27303,N_26990,N_26982);
nor U27304 (N_27304,N_26911,N_26645);
or U27305 (N_27305,N_26558,N_26878);
xnor U27306 (N_27306,N_26712,N_26543);
or U27307 (N_27307,N_26719,N_26957);
or U27308 (N_27308,N_26691,N_26718);
and U27309 (N_27309,N_26664,N_26916);
or U27310 (N_27310,N_26887,N_26950);
and U27311 (N_27311,N_26521,N_26725);
nand U27312 (N_27312,N_26564,N_26666);
xnor U27313 (N_27313,N_26712,N_26529);
or U27314 (N_27314,N_26616,N_26524);
nor U27315 (N_27315,N_26580,N_26893);
or U27316 (N_27316,N_26687,N_26653);
nand U27317 (N_27317,N_26615,N_26503);
or U27318 (N_27318,N_26932,N_26507);
nand U27319 (N_27319,N_26676,N_26960);
nand U27320 (N_27320,N_26897,N_26618);
nor U27321 (N_27321,N_26595,N_26942);
or U27322 (N_27322,N_26608,N_26744);
nand U27323 (N_27323,N_26696,N_26541);
nand U27324 (N_27324,N_26643,N_26588);
nand U27325 (N_27325,N_26609,N_26774);
nor U27326 (N_27326,N_26742,N_26951);
nand U27327 (N_27327,N_26879,N_26975);
xor U27328 (N_27328,N_26594,N_26788);
xnor U27329 (N_27329,N_26871,N_26995);
or U27330 (N_27330,N_26799,N_26658);
or U27331 (N_27331,N_26762,N_26528);
nand U27332 (N_27332,N_26591,N_26900);
nor U27333 (N_27333,N_26552,N_26643);
nand U27334 (N_27334,N_26516,N_26605);
nor U27335 (N_27335,N_26826,N_26610);
nor U27336 (N_27336,N_26971,N_26718);
or U27337 (N_27337,N_26898,N_26583);
nand U27338 (N_27338,N_26503,N_26892);
and U27339 (N_27339,N_26866,N_26797);
nor U27340 (N_27340,N_26838,N_26959);
nand U27341 (N_27341,N_26951,N_26732);
nand U27342 (N_27342,N_26680,N_26904);
and U27343 (N_27343,N_26668,N_26710);
nor U27344 (N_27344,N_26860,N_26548);
and U27345 (N_27345,N_26510,N_26640);
nor U27346 (N_27346,N_26791,N_26969);
nand U27347 (N_27347,N_26584,N_26874);
xnor U27348 (N_27348,N_26522,N_26605);
nand U27349 (N_27349,N_26642,N_26966);
xor U27350 (N_27350,N_26691,N_26820);
nor U27351 (N_27351,N_26820,N_26517);
xnor U27352 (N_27352,N_26511,N_26779);
xnor U27353 (N_27353,N_26693,N_26631);
xor U27354 (N_27354,N_26600,N_26979);
and U27355 (N_27355,N_26606,N_26790);
nor U27356 (N_27356,N_26546,N_26720);
and U27357 (N_27357,N_26757,N_26831);
or U27358 (N_27358,N_26724,N_26536);
and U27359 (N_27359,N_26548,N_26654);
and U27360 (N_27360,N_26862,N_26641);
or U27361 (N_27361,N_26592,N_26597);
nand U27362 (N_27362,N_26704,N_26902);
xor U27363 (N_27363,N_26702,N_26847);
or U27364 (N_27364,N_26982,N_26958);
or U27365 (N_27365,N_26747,N_26805);
xor U27366 (N_27366,N_26759,N_26954);
xnor U27367 (N_27367,N_26697,N_26963);
and U27368 (N_27368,N_26975,N_26887);
nand U27369 (N_27369,N_26593,N_26897);
or U27370 (N_27370,N_26547,N_26907);
nor U27371 (N_27371,N_26523,N_26857);
nand U27372 (N_27372,N_26899,N_26781);
nor U27373 (N_27373,N_26952,N_26729);
xnor U27374 (N_27374,N_26810,N_26553);
xor U27375 (N_27375,N_26920,N_26748);
nor U27376 (N_27376,N_26850,N_26612);
nor U27377 (N_27377,N_26986,N_26913);
and U27378 (N_27378,N_26677,N_26959);
nand U27379 (N_27379,N_26550,N_26570);
xnor U27380 (N_27380,N_26746,N_26516);
nor U27381 (N_27381,N_26842,N_26527);
xor U27382 (N_27382,N_26781,N_26911);
and U27383 (N_27383,N_26795,N_26578);
or U27384 (N_27384,N_26502,N_26716);
and U27385 (N_27385,N_26609,N_26501);
or U27386 (N_27386,N_26537,N_26970);
nor U27387 (N_27387,N_26673,N_26777);
xor U27388 (N_27388,N_26981,N_26793);
nor U27389 (N_27389,N_26678,N_26887);
nor U27390 (N_27390,N_26826,N_26799);
nand U27391 (N_27391,N_26948,N_26660);
xor U27392 (N_27392,N_26948,N_26899);
nand U27393 (N_27393,N_26767,N_26723);
or U27394 (N_27394,N_26800,N_26551);
or U27395 (N_27395,N_26621,N_26680);
nor U27396 (N_27396,N_26797,N_26734);
and U27397 (N_27397,N_26722,N_26924);
nand U27398 (N_27398,N_26734,N_26774);
xor U27399 (N_27399,N_26597,N_26811);
or U27400 (N_27400,N_26595,N_26907);
nor U27401 (N_27401,N_26725,N_26780);
nand U27402 (N_27402,N_26996,N_26961);
and U27403 (N_27403,N_26838,N_26853);
and U27404 (N_27404,N_26570,N_26948);
or U27405 (N_27405,N_26858,N_26719);
xor U27406 (N_27406,N_26845,N_26669);
nor U27407 (N_27407,N_26671,N_26778);
nor U27408 (N_27408,N_26762,N_26917);
nand U27409 (N_27409,N_26940,N_26995);
xnor U27410 (N_27410,N_26827,N_26741);
nand U27411 (N_27411,N_26619,N_26849);
and U27412 (N_27412,N_26829,N_26804);
nand U27413 (N_27413,N_26605,N_26859);
nand U27414 (N_27414,N_26953,N_26750);
or U27415 (N_27415,N_26845,N_26759);
or U27416 (N_27416,N_26746,N_26976);
xnor U27417 (N_27417,N_26542,N_26539);
nor U27418 (N_27418,N_26513,N_26800);
and U27419 (N_27419,N_26941,N_26588);
or U27420 (N_27420,N_26665,N_26959);
nand U27421 (N_27421,N_26629,N_26955);
nor U27422 (N_27422,N_26724,N_26673);
nand U27423 (N_27423,N_26891,N_26863);
nor U27424 (N_27424,N_26680,N_26910);
nand U27425 (N_27425,N_26897,N_26983);
or U27426 (N_27426,N_26871,N_26620);
nand U27427 (N_27427,N_26910,N_26560);
and U27428 (N_27428,N_26889,N_26814);
xor U27429 (N_27429,N_26746,N_26558);
or U27430 (N_27430,N_26618,N_26829);
and U27431 (N_27431,N_26969,N_26732);
xor U27432 (N_27432,N_26855,N_26942);
xor U27433 (N_27433,N_26724,N_26654);
xnor U27434 (N_27434,N_26886,N_26816);
xnor U27435 (N_27435,N_26684,N_26862);
or U27436 (N_27436,N_26571,N_26889);
or U27437 (N_27437,N_26767,N_26519);
nand U27438 (N_27438,N_26774,N_26754);
xnor U27439 (N_27439,N_26858,N_26780);
xor U27440 (N_27440,N_26573,N_26971);
or U27441 (N_27441,N_26906,N_26654);
nor U27442 (N_27442,N_26544,N_26976);
xor U27443 (N_27443,N_26872,N_26592);
nand U27444 (N_27444,N_26913,N_26969);
nor U27445 (N_27445,N_26635,N_26706);
nor U27446 (N_27446,N_26768,N_26522);
and U27447 (N_27447,N_26612,N_26677);
or U27448 (N_27448,N_26991,N_26533);
nand U27449 (N_27449,N_26780,N_26747);
xor U27450 (N_27450,N_26780,N_26915);
and U27451 (N_27451,N_26866,N_26589);
and U27452 (N_27452,N_26802,N_26553);
or U27453 (N_27453,N_26573,N_26784);
or U27454 (N_27454,N_26918,N_26724);
nand U27455 (N_27455,N_26512,N_26689);
nor U27456 (N_27456,N_26914,N_26722);
or U27457 (N_27457,N_26546,N_26866);
nand U27458 (N_27458,N_26935,N_26540);
nand U27459 (N_27459,N_26559,N_26688);
nor U27460 (N_27460,N_26744,N_26637);
nor U27461 (N_27461,N_26878,N_26713);
xnor U27462 (N_27462,N_26654,N_26549);
and U27463 (N_27463,N_26802,N_26903);
or U27464 (N_27464,N_26602,N_26854);
nand U27465 (N_27465,N_26868,N_26988);
or U27466 (N_27466,N_26573,N_26676);
or U27467 (N_27467,N_26983,N_26961);
and U27468 (N_27468,N_26527,N_26969);
nor U27469 (N_27469,N_26874,N_26578);
xnor U27470 (N_27470,N_26553,N_26869);
or U27471 (N_27471,N_26521,N_26771);
xnor U27472 (N_27472,N_26634,N_26540);
nor U27473 (N_27473,N_26942,N_26840);
nand U27474 (N_27474,N_26923,N_26937);
xnor U27475 (N_27475,N_26986,N_26710);
and U27476 (N_27476,N_26936,N_26658);
and U27477 (N_27477,N_26868,N_26607);
and U27478 (N_27478,N_26852,N_26547);
or U27479 (N_27479,N_26533,N_26798);
xnor U27480 (N_27480,N_26682,N_26910);
and U27481 (N_27481,N_26706,N_26963);
and U27482 (N_27482,N_26858,N_26926);
xnor U27483 (N_27483,N_26955,N_26732);
nand U27484 (N_27484,N_26724,N_26716);
or U27485 (N_27485,N_26899,N_26815);
xor U27486 (N_27486,N_26837,N_26563);
nor U27487 (N_27487,N_26986,N_26985);
and U27488 (N_27488,N_26634,N_26516);
nor U27489 (N_27489,N_26820,N_26808);
and U27490 (N_27490,N_26807,N_26671);
nor U27491 (N_27491,N_26941,N_26760);
nor U27492 (N_27492,N_26757,N_26949);
or U27493 (N_27493,N_26940,N_26689);
nand U27494 (N_27494,N_26782,N_26871);
nand U27495 (N_27495,N_26558,N_26797);
nor U27496 (N_27496,N_26831,N_26538);
or U27497 (N_27497,N_26934,N_26526);
nand U27498 (N_27498,N_26703,N_26804);
nor U27499 (N_27499,N_26835,N_26845);
or U27500 (N_27500,N_27045,N_27241);
nor U27501 (N_27501,N_27176,N_27478);
nand U27502 (N_27502,N_27000,N_27457);
xnor U27503 (N_27503,N_27170,N_27023);
nor U27504 (N_27504,N_27197,N_27008);
or U27505 (N_27505,N_27147,N_27489);
nor U27506 (N_27506,N_27400,N_27096);
xnor U27507 (N_27507,N_27115,N_27180);
nor U27508 (N_27508,N_27325,N_27101);
nand U27509 (N_27509,N_27164,N_27324);
xnor U27510 (N_27510,N_27102,N_27090);
nor U27511 (N_27511,N_27282,N_27066);
or U27512 (N_27512,N_27485,N_27049);
nor U27513 (N_27513,N_27153,N_27472);
xor U27514 (N_27514,N_27309,N_27065);
or U27515 (N_27515,N_27431,N_27021);
xor U27516 (N_27516,N_27301,N_27459);
or U27517 (N_27517,N_27005,N_27482);
xor U27518 (N_27518,N_27006,N_27055);
and U27519 (N_27519,N_27119,N_27015);
nor U27520 (N_27520,N_27320,N_27385);
xnor U27521 (N_27521,N_27022,N_27393);
nand U27522 (N_27522,N_27307,N_27299);
nor U27523 (N_27523,N_27486,N_27037);
nor U27524 (N_27524,N_27283,N_27243);
or U27525 (N_27525,N_27435,N_27098);
or U27526 (N_27526,N_27003,N_27201);
xor U27527 (N_27527,N_27162,N_27268);
xor U27528 (N_27528,N_27257,N_27117);
nand U27529 (N_27529,N_27092,N_27044);
nand U27530 (N_27530,N_27345,N_27134);
or U27531 (N_27531,N_27086,N_27137);
nor U27532 (N_27532,N_27349,N_27246);
or U27533 (N_27533,N_27122,N_27293);
nor U27534 (N_27534,N_27200,N_27326);
nor U27535 (N_27535,N_27218,N_27313);
xor U27536 (N_27536,N_27379,N_27421);
nand U27537 (N_27537,N_27109,N_27468);
and U27538 (N_27538,N_27123,N_27494);
xnor U27539 (N_27539,N_27351,N_27396);
and U27540 (N_27540,N_27208,N_27083);
or U27541 (N_27541,N_27236,N_27451);
and U27542 (N_27542,N_27234,N_27380);
and U27543 (N_27543,N_27461,N_27408);
nand U27544 (N_27544,N_27338,N_27288);
xor U27545 (N_27545,N_27465,N_27254);
nand U27546 (N_27546,N_27437,N_27477);
nor U27547 (N_27547,N_27280,N_27496);
nor U27548 (N_27548,N_27377,N_27108);
xor U27549 (N_27549,N_27375,N_27088);
xnor U27550 (N_27550,N_27394,N_27427);
xnor U27551 (N_27551,N_27429,N_27031);
nor U27552 (N_27552,N_27321,N_27404);
nor U27553 (N_27553,N_27172,N_27253);
and U27554 (N_27554,N_27284,N_27306);
or U27555 (N_27555,N_27185,N_27413);
nand U27556 (N_27556,N_27447,N_27138);
and U27557 (N_27557,N_27228,N_27355);
xor U27558 (N_27558,N_27295,N_27417);
or U27559 (N_27559,N_27312,N_27030);
and U27560 (N_27560,N_27106,N_27329);
nand U27561 (N_27561,N_27418,N_27034);
nor U27562 (N_27562,N_27263,N_27036);
xor U27563 (N_27563,N_27422,N_27047);
xnor U27564 (N_27564,N_27463,N_27099);
xnor U27565 (N_27565,N_27296,N_27395);
or U27566 (N_27566,N_27113,N_27371);
xor U27567 (N_27567,N_27020,N_27124);
and U27568 (N_27568,N_27085,N_27412);
or U27569 (N_27569,N_27432,N_27270);
nor U27570 (N_27570,N_27160,N_27214);
nand U27571 (N_27571,N_27074,N_27084);
nand U27572 (N_27572,N_27439,N_27490);
and U27573 (N_27573,N_27310,N_27484);
and U27574 (N_27574,N_27370,N_27247);
xnor U27575 (N_27575,N_27237,N_27466);
nor U27576 (N_27576,N_27365,N_27029);
xor U27577 (N_27577,N_27093,N_27225);
nor U27578 (N_27578,N_27133,N_27205);
xnor U27579 (N_27579,N_27112,N_27300);
nand U27580 (N_27580,N_27155,N_27195);
xor U27581 (N_27581,N_27464,N_27233);
nor U27582 (N_27582,N_27352,N_27460);
or U27583 (N_27583,N_27317,N_27186);
or U27584 (N_27584,N_27441,N_27054);
nand U27585 (N_27585,N_27043,N_27152);
and U27586 (N_27586,N_27042,N_27358);
and U27587 (N_27587,N_27095,N_27058);
nand U27588 (N_27588,N_27497,N_27311);
xor U27589 (N_27589,N_27278,N_27025);
nand U27590 (N_27590,N_27438,N_27156);
or U27591 (N_27591,N_27190,N_27075);
and U27592 (N_27592,N_27368,N_27245);
xnor U27593 (N_27593,N_27107,N_27322);
nor U27594 (N_27594,N_27266,N_27433);
and U27595 (N_27595,N_27004,N_27056);
and U27596 (N_27596,N_27239,N_27292);
xnor U27597 (N_27597,N_27077,N_27078);
nand U27598 (N_27598,N_27333,N_27327);
nand U27599 (N_27599,N_27420,N_27135);
or U27600 (N_27600,N_27294,N_27181);
xor U27601 (N_27601,N_27399,N_27027);
xor U27602 (N_27602,N_27232,N_27014);
nor U27603 (N_27603,N_27182,N_27040);
nor U27604 (N_27604,N_27011,N_27430);
nor U27605 (N_27605,N_27498,N_27224);
nor U27606 (N_27606,N_27255,N_27059);
nand U27607 (N_27607,N_27426,N_27206);
nand U27608 (N_27608,N_27024,N_27150);
or U27609 (N_27609,N_27127,N_27171);
nand U27610 (N_27610,N_27362,N_27388);
or U27611 (N_27611,N_27428,N_27342);
or U27612 (N_27612,N_27053,N_27364);
or U27613 (N_27613,N_27425,N_27390);
or U27614 (N_27614,N_27258,N_27481);
or U27615 (N_27615,N_27013,N_27244);
nor U27616 (N_27616,N_27252,N_27403);
xor U27617 (N_27617,N_27302,N_27443);
and U27618 (N_27618,N_27374,N_27456);
and U27619 (N_27619,N_27341,N_27248);
nor U27620 (N_27620,N_27082,N_27256);
nand U27621 (N_27621,N_27473,N_27297);
or U27622 (N_27622,N_27340,N_27328);
nor U27623 (N_27623,N_27470,N_27491);
nor U27624 (N_27624,N_27193,N_27046);
nor U27625 (N_27625,N_27479,N_27227);
nand U27626 (N_27626,N_27273,N_27488);
and U27627 (N_27627,N_27018,N_27183);
xor U27628 (N_27628,N_27097,N_27213);
nor U27629 (N_27629,N_27261,N_27226);
nor U27630 (N_27630,N_27409,N_27116);
xor U27631 (N_27631,N_27444,N_27265);
nor U27632 (N_27632,N_27010,N_27149);
or U27633 (N_27633,N_27346,N_27048);
or U27634 (N_27634,N_27363,N_27269);
nor U27635 (N_27635,N_27189,N_27166);
nand U27636 (N_27636,N_27126,N_27033);
nand U27637 (N_27637,N_27383,N_27052);
xnor U27638 (N_27638,N_27279,N_27072);
xnor U27639 (N_27639,N_27209,N_27387);
or U27640 (N_27640,N_27009,N_27114);
or U27641 (N_27641,N_27357,N_27220);
or U27642 (N_27642,N_27323,N_27251);
nand U27643 (N_27643,N_27392,N_27175);
nand U27644 (N_27644,N_27410,N_27452);
xor U27645 (N_27645,N_27262,N_27035);
and U27646 (N_27646,N_27217,N_27071);
or U27647 (N_27647,N_27446,N_27369);
or U27648 (N_27648,N_27305,N_27450);
and U27649 (N_27649,N_27344,N_27148);
or U27650 (N_27650,N_27291,N_27304);
nor U27651 (N_27651,N_27177,N_27240);
nand U27652 (N_27652,N_27129,N_27210);
xnor U27653 (N_27653,N_27499,N_27067);
nor U27654 (N_27654,N_27219,N_27492);
nor U27655 (N_27655,N_27480,N_27070);
nand U27656 (N_27656,N_27064,N_27212);
xor U27657 (N_27657,N_27467,N_27398);
and U27658 (N_27658,N_27314,N_27203);
nand U27659 (N_27659,N_27384,N_27407);
xor U27660 (N_27660,N_27389,N_27125);
or U27661 (N_27661,N_27194,N_27143);
nor U27662 (N_27662,N_27272,N_27289);
xor U27663 (N_27663,N_27332,N_27469);
or U27664 (N_27664,N_27163,N_27386);
nand U27665 (N_27665,N_27416,N_27100);
nand U27666 (N_27666,N_27118,N_27453);
nor U27667 (N_27667,N_27068,N_27196);
and U27668 (N_27668,N_27179,N_27287);
nor U27669 (N_27669,N_27026,N_27360);
nand U27670 (N_27670,N_27128,N_27319);
or U27671 (N_27671,N_27303,N_27264);
and U27672 (N_27672,N_27142,N_27415);
or U27673 (N_27673,N_27238,N_27204);
or U27674 (N_27674,N_27454,N_27120);
or U27675 (N_27675,N_27285,N_27495);
nor U27676 (N_27676,N_27347,N_27381);
or U27677 (N_27677,N_27016,N_27493);
xor U27678 (N_27678,N_27455,N_27373);
nor U27679 (N_27679,N_27073,N_27089);
or U27680 (N_27680,N_27230,N_27343);
nor U27681 (N_27681,N_27187,N_27235);
xor U27682 (N_27682,N_27221,N_27475);
and U27683 (N_27683,N_27121,N_27144);
xor U27684 (N_27684,N_27103,N_27051);
nand U27685 (N_27685,N_27002,N_27315);
xor U27686 (N_27686,N_27242,N_27061);
xor U27687 (N_27687,N_27110,N_27423);
nand U27688 (N_27688,N_27157,N_27174);
nor U27689 (N_27689,N_27382,N_27458);
xnor U27690 (N_27690,N_27216,N_27168);
nor U27691 (N_27691,N_27483,N_27259);
xor U27692 (N_27692,N_27231,N_27376);
nand U27693 (N_27693,N_27361,N_27334);
nor U27694 (N_27694,N_27104,N_27032);
nand U27695 (N_27695,N_27419,N_27378);
or U27696 (N_27696,N_27286,N_27330);
nor U27697 (N_27697,N_27161,N_27146);
nor U27698 (N_27698,N_27350,N_27474);
nor U27699 (N_27699,N_27277,N_27434);
nand U27700 (N_27700,N_27192,N_27339);
xor U27701 (N_27701,N_27308,N_27130);
xnor U27702 (N_27702,N_27318,N_27487);
xnor U27703 (N_27703,N_27159,N_27372);
xor U27704 (N_27704,N_27391,N_27298);
and U27705 (N_27705,N_27359,N_27348);
or U27706 (N_27706,N_27184,N_27424);
nand U27707 (N_27707,N_27202,N_27366);
and U27708 (N_27708,N_27087,N_27215);
or U27709 (N_27709,N_27111,N_27411);
nand U27710 (N_27710,N_27354,N_27198);
xnor U27711 (N_27711,N_27260,N_27145);
and U27712 (N_27712,N_27356,N_27405);
or U27713 (N_27713,N_27276,N_27080);
or U27714 (N_27714,N_27039,N_27076);
or U27715 (N_27715,N_27141,N_27136);
or U27716 (N_27716,N_27471,N_27139);
or U27717 (N_27717,N_27414,N_27316);
and U27718 (N_27718,N_27442,N_27250);
xnor U27719 (N_27719,N_27154,N_27173);
and U27720 (N_27720,N_27207,N_27062);
nand U27721 (N_27721,N_27131,N_27274);
and U27722 (N_27722,N_27038,N_27436);
nor U27723 (N_27723,N_27367,N_27290);
nand U27724 (N_27724,N_27165,N_27140);
or U27725 (N_27725,N_27017,N_27081);
xor U27726 (N_27726,N_27057,N_27397);
xor U27727 (N_27727,N_27222,N_27401);
nor U27728 (N_27728,N_27158,N_27267);
nand U27729 (N_27729,N_27249,N_27335);
or U27730 (N_27730,N_27331,N_27440);
and U27731 (N_27731,N_27105,N_27281);
or U27732 (N_27732,N_27462,N_27275);
or U27733 (N_27733,N_27063,N_27402);
xor U27734 (N_27734,N_27448,N_27336);
nor U27735 (N_27735,N_27079,N_27050);
nor U27736 (N_27736,N_27167,N_27476);
xor U27737 (N_27737,N_27069,N_27169);
nand U27738 (N_27738,N_27094,N_27041);
nor U27739 (N_27739,N_27012,N_27406);
nand U27740 (N_27740,N_27019,N_27229);
xor U27741 (N_27741,N_27353,N_27191);
nor U27742 (N_27742,N_27271,N_27337);
or U27743 (N_27743,N_27132,N_27223);
nand U27744 (N_27744,N_27199,N_27091);
nand U27745 (N_27745,N_27001,N_27178);
nor U27746 (N_27746,N_27007,N_27445);
nor U27747 (N_27747,N_27028,N_27449);
xor U27748 (N_27748,N_27211,N_27188);
nand U27749 (N_27749,N_27151,N_27060);
nor U27750 (N_27750,N_27050,N_27126);
nand U27751 (N_27751,N_27271,N_27303);
or U27752 (N_27752,N_27177,N_27180);
nor U27753 (N_27753,N_27490,N_27195);
and U27754 (N_27754,N_27365,N_27417);
and U27755 (N_27755,N_27470,N_27110);
nor U27756 (N_27756,N_27499,N_27449);
and U27757 (N_27757,N_27244,N_27126);
xor U27758 (N_27758,N_27170,N_27282);
and U27759 (N_27759,N_27053,N_27033);
and U27760 (N_27760,N_27345,N_27076);
or U27761 (N_27761,N_27446,N_27324);
nor U27762 (N_27762,N_27196,N_27351);
or U27763 (N_27763,N_27175,N_27070);
nand U27764 (N_27764,N_27354,N_27158);
nor U27765 (N_27765,N_27180,N_27475);
nor U27766 (N_27766,N_27206,N_27019);
and U27767 (N_27767,N_27018,N_27246);
nand U27768 (N_27768,N_27036,N_27243);
or U27769 (N_27769,N_27187,N_27337);
or U27770 (N_27770,N_27090,N_27478);
xnor U27771 (N_27771,N_27429,N_27239);
nor U27772 (N_27772,N_27178,N_27290);
and U27773 (N_27773,N_27254,N_27347);
nor U27774 (N_27774,N_27494,N_27093);
nand U27775 (N_27775,N_27211,N_27389);
or U27776 (N_27776,N_27129,N_27147);
nand U27777 (N_27777,N_27205,N_27318);
nand U27778 (N_27778,N_27255,N_27039);
and U27779 (N_27779,N_27485,N_27258);
or U27780 (N_27780,N_27445,N_27100);
xnor U27781 (N_27781,N_27143,N_27271);
xnor U27782 (N_27782,N_27283,N_27259);
and U27783 (N_27783,N_27240,N_27057);
nand U27784 (N_27784,N_27001,N_27201);
nor U27785 (N_27785,N_27320,N_27042);
xor U27786 (N_27786,N_27474,N_27249);
or U27787 (N_27787,N_27409,N_27145);
nor U27788 (N_27788,N_27255,N_27271);
or U27789 (N_27789,N_27121,N_27309);
nor U27790 (N_27790,N_27108,N_27398);
xor U27791 (N_27791,N_27494,N_27293);
or U27792 (N_27792,N_27047,N_27221);
nand U27793 (N_27793,N_27081,N_27342);
and U27794 (N_27794,N_27093,N_27180);
nand U27795 (N_27795,N_27140,N_27054);
and U27796 (N_27796,N_27220,N_27039);
and U27797 (N_27797,N_27052,N_27185);
and U27798 (N_27798,N_27204,N_27369);
and U27799 (N_27799,N_27395,N_27431);
nor U27800 (N_27800,N_27214,N_27014);
and U27801 (N_27801,N_27264,N_27283);
and U27802 (N_27802,N_27018,N_27030);
xnor U27803 (N_27803,N_27369,N_27441);
nand U27804 (N_27804,N_27097,N_27285);
or U27805 (N_27805,N_27054,N_27180);
nor U27806 (N_27806,N_27453,N_27046);
and U27807 (N_27807,N_27299,N_27273);
nand U27808 (N_27808,N_27431,N_27285);
xor U27809 (N_27809,N_27209,N_27221);
xor U27810 (N_27810,N_27246,N_27144);
nand U27811 (N_27811,N_27404,N_27082);
xnor U27812 (N_27812,N_27102,N_27027);
and U27813 (N_27813,N_27059,N_27433);
nor U27814 (N_27814,N_27428,N_27193);
or U27815 (N_27815,N_27251,N_27335);
or U27816 (N_27816,N_27237,N_27436);
nor U27817 (N_27817,N_27289,N_27165);
nor U27818 (N_27818,N_27017,N_27421);
nand U27819 (N_27819,N_27407,N_27104);
and U27820 (N_27820,N_27151,N_27232);
nand U27821 (N_27821,N_27103,N_27247);
xnor U27822 (N_27822,N_27056,N_27279);
nor U27823 (N_27823,N_27270,N_27251);
xnor U27824 (N_27824,N_27053,N_27088);
nand U27825 (N_27825,N_27049,N_27327);
nand U27826 (N_27826,N_27058,N_27291);
nor U27827 (N_27827,N_27110,N_27336);
or U27828 (N_27828,N_27009,N_27053);
nand U27829 (N_27829,N_27486,N_27434);
xnor U27830 (N_27830,N_27113,N_27247);
and U27831 (N_27831,N_27226,N_27277);
nand U27832 (N_27832,N_27357,N_27127);
nand U27833 (N_27833,N_27232,N_27214);
nand U27834 (N_27834,N_27382,N_27221);
and U27835 (N_27835,N_27077,N_27133);
and U27836 (N_27836,N_27423,N_27121);
and U27837 (N_27837,N_27091,N_27422);
nand U27838 (N_27838,N_27165,N_27320);
xnor U27839 (N_27839,N_27391,N_27232);
or U27840 (N_27840,N_27007,N_27114);
xor U27841 (N_27841,N_27241,N_27129);
nand U27842 (N_27842,N_27436,N_27014);
xor U27843 (N_27843,N_27222,N_27080);
nand U27844 (N_27844,N_27093,N_27216);
nor U27845 (N_27845,N_27460,N_27073);
and U27846 (N_27846,N_27410,N_27005);
xor U27847 (N_27847,N_27491,N_27112);
xor U27848 (N_27848,N_27069,N_27411);
and U27849 (N_27849,N_27151,N_27283);
nor U27850 (N_27850,N_27443,N_27178);
xnor U27851 (N_27851,N_27372,N_27209);
or U27852 (N_27852,N_27112,N_27381);
or U27853 (N_27853,N_27103,N_27288);
nand U27854 (N_27854,N_27062,N_27230);
xnor U27855 (N_27855,N_27486,N_27010);
nand U27856 (N_27856,N_27291,N_27124);
nand U27857 (N_27857,N_27199,N_27491);
or U27858 (N_27858,N_27188,N_27146);
nor U27859 (N_27859,N_27269,N_27311);
and U27860 (N_27860,N_27177,N_27166);
nor U27861 (N_27861,N_27386,N_27212);
and U27862 (N_27862,N_27043,N_27306);
nor U27863 (N_27863,N_27087,N_27339);
nand U27864 (N_27864,N_27278,N_27352);
nor U27865 (N_27865,N_27399,N_27401);
and U27866 (N_27866,N_27117,N_27431);
and U27867 (N_27867,N_27312,N_27070);
and U27868 (N_27868,N_27331,N_27032);
xnor U27869 (N_27869,N_27253,N_27338);
xor U27870 (N_27870,N_27432,N_27172);
and U27871 (N_27871,N_27404,N_27118);
xnor U27872 (N_27872,N_27335,N_27290);
xnor U27873 (N_27873,N_27127,N_27436);
nor U27874 (N_27874,N_27459,N_27274);
and U27875 (N_27875,N_27169,N_27281);
or U27876 (N_27876,N_27231,N_27473);
or U27877 (N_27877,N_27157,N_27089);
and U27878 (N_27878,N_27309,N_27063);
xor U27879 (N_27879,N_27113,N_27229);
and U27880 (N_27880,N_27332,N_27317);
nor U27881 (N_27881,N_27077,N_27085);
or U27882 (N_27882,N_27155,N_27138);
xnor U27883 (N_27883,N_27476,N_27026);
xor U27884 (N_27884,N_27470,N_27493);
and U27885 (N_27885,N_27229,N_27179);
nand U27886 (N_27886,N_27026,N_27098);
xor U27887 (N_27887,N_27007,N_27373);
nand U27888 (N_27888,N_27215,N_27253);
nor U27889 (N_27889,N_27448,N_27297);
or U27890 (N_27890,N_27298,N_27100);
xor U27891 (N_27891,N_27057,N_27047);
nand U27892 (N_27892,N_27183,N_27121);
or U27893 (N_27893,N_27258,N_27401);
or U27894 (N_27894,N_27262,N_27223);
xor U27895 (N_27895,N_27420,N_27086);
nand U27896 (N_27896,N_27278,N_27010);
and U27897 (N_27897,N_27011,N_27205);
or U27898 (N_27898,N_27405,N_27267);
or U27899 (N_27899,N_27410,N_27279);
nand U27900 (N_27900,N_27078,N_27222);
and U27901 (N_27901,N_27234,N_27092);
xnor U27902 (N_27902,N_27181,N_27220);
or U27903 (N_27903,N_27369,N_27391);
or U27904 (N_27904,N_27045,N_27066);
and U27905 (N_27905,N_27145,N_27216);
and U27906 (N_27906,N_27486,N_27489);
xor U27907 (N_27907,N_27323,N_27131);
xor U27908 (N_27908,N_27128,N_27120);
and U27909 (N_27909,N_27394,N_27291);
or U27910 (N_27910,N_27486,N_27258);
xnor U27911 (N_27911,N_27414,N_27125);
nand U27912 (N_27912,N_27000,N_27281);
nand U27913 (N_27913,N_27306,N_27166);
nor U27914 (N_27914,N_27293,N_27005);
nor U27915 (N_27915,N_27064,N_27238);
nor U27916 (N_27916,N_27268,N_27007);
nor U27917 (N_27917,N_27333,N_27008);
xor U27918 (N_27918,N_27244,N_27023);
nor U27919 (N_27919,N_27057,N_27205);
and U27920 (N_27920,N_27454,N_27313);
nor U27921 (N_27921,N_27235,N_27262);
nor U27922 (N_27922,N_27157,N_27112);
nor U27923 (N_27923,N_27377,N_27219);
nor U27924 (N_27924,N_27060,N_27207);
xor U27925 (N_27925,N_27187,N_27193);
or U27926 (N_27926,N_27001,N_27477);
nand U27927 (N_27927,N_27088,N_27176);
xor U27928 (N_27928,N_27318,N_27321);
xor U27929 (N_27929,N_27245,N_27481);
or U27930 (N_27930,N_27122,N_27101);
or U27931 (N_27931,N_27392,N_27332);
xnor U27932 (N_27932,N_27001,N_27061);
xor U27933 (N_27933,N_27099,N_27136);
nand U27934 (N_27934,N_27257,N_27498);
nand U27935 (N_27935,N_27443,N_27310);
xor U27936 (N_27936,N_27174,N_27263);
xnor U27937 (N_27937,N_27320,N_27172);
nor U27938 (N_27938,N_27121,N_27343);
or U27939 (N_27939,N_27277,N_27435);
or U27940 (N_27940,N_27150,N_27309);
and U27941 (N_27941,N_27444,N_27279);
and U27942 (N_27942,N_27066,N_27027);
nor U27943 (N_27943,N_27291,N_27163);
nor U27944 (N_27944,N_27159,N_27456);
and U27945 (N_27945,N_27146,N_27470);
xor U27946 (N_27946,N_27415,N_27110);
xnor U27947 (N_27947,N_27177,N_27075);
and U27948 (N_27948,N_27196,N_27459);
or U27949 (N_27949,N_27033,N_27054);
xor U27950 (N_27950,N_27011,N_27423);
xnor U27951 (N_27951,N_27458,N_27300);
and U27952 (N_27952,N_27228,N_27193);
nor U27953 (N_27953,N_27446,N_27056);
or U27954 (N_27954,N_27354,N_27327);
nand U27955 (N_27955,N_27172,N_27139);
xnor U27956 (N_27956,N_27038,N_27108);
nand U27957 (N_27957,N_27082,N_27162);
or U27958 (N_27958,N_27493,N_27312);
xor U27959 (N_27959,N_27393,N_27103);
or U27960 (N_27960,N_27245,N_27230);
nor U27961 (N_27961,N_27461,N_27007);
nand U27962 (N_27962,N_27305,N_27141);
nand U27963 (N_27963,N_27026,N_27289);
nand U27964 (N_27964,N_27064,N_27397);
nor U27965 (N_27965,N_27469,N_27367);
or U27966 (N_27966,N_27325,N_27249);
nor U27967 (N_27967,N_27430,N_27150);
nor U27968 (N_27968,N_27114,N_27122);
and U27969 (N_27969,N_27003,N_27158);
xnor U27970 (N_27970,N_27481,N_27330);
nand U27971 (N_27971,N_27297,N_27349);
xnor U27972 (N_27972,N_27397,N_27287);
or U27973 (N_27973,N_27126,N_27172);
nor U27974 (N_27974,N_27265,N_27186);
and U27975 (N_27975,N_27026,N_27433);
nand U27976 (N_27976,N_27243,N_27290);
nor U27977 (N_27977,N_27457,N_27264);
and U27978 (N_27978,N_27207,N_27125);
xor U27979 (N_27979,N_27436,N_27228);
nand U27980 (N_27980,N_27214,N_27288);
and U27981 (N_27981,N_27017,N_27301);
or U27982 (N_27982,N_27493,N_27478);
nor U27983 (N_27983,N_27176,N_27183);
nor U27984 (N_27984,N_27204,N_27074);
nand U27985 (N_27985,N_27287,N_27407);
nor U27986 (N_27986,N_27204,N_27320);
nor U27987 (N_27987,N_27218,N_27449);
nand U27988 (N_27988,N_27246,N_27033);
nand U27989 (N_27989,N_27447,N_27087);
nand U27990 (N_27990,N_27143,N_27356);
nand U27991 (N_27991,N_27290,N_27259);
xor U27992 (N_27992,N_27481,N_27490);
nor U27993 (N_27993,N_27363,N_27292);
xor U27994 (N_27994,N_27056,N_27466);
nor U27995 (N_27995,N_27050,N_27476);
nand U27996 (N_27996,N_27105,N_27439);
and U27997 (N_27997,N_27268,N_27423);
or U27998 (N_27998,N_27392,N_27353);
nor U27999 (N_27999,N_27406,N_27062);
nand U28000 (N_28000,N_27726,N_27712);
or U28001 (N_28001,N_27979,N_27731);
nor U28002 (N_28002,N_27538,N_27813);
nor U28003 (N_28003,N_27877,N_27748);
xnor U28004 (N_28004,N_27986,N_27524);
nand U28005 (N_28005,N_27832,N_27753);
nand U28006 (N_28006,N_27711,N_27937);
and U28007 (N_28007,N_27807,N_27588);
or U28008 (N_28008,N_27963,N_27627);
and U28009 (N_28009,N_27626,N_27826);
or U28010 (N_28010,N_27985,N_27968);
nand U28011 (N_28011,N_27933,N_27722);
nand U28012 (N_28012,N_27769,N_27863);
nand U28013 (N_28013,N_27938,N_27589);
nor U28014 (N_28014,N_27502,N_27660);
or U28015 (N_28015,N_27921,N_27603);
or U28016 (N_28016,N_27892,N_27959);
nand U28017 (N_28017,N_27567,N_27719);
and U28018 (N_28018,N_27874,N_27806);
or U28019 (N_28019,N_27565,N_27971);
or U28020 (N_28020,N_27966,N_27886);
or U28021 (N_28021,N_27695,N_27707);
or U28022 (N_28022,N_27685,N_27773);
nand U28023 (N_28023,N_27500,N_27584);
or U28024 (N_28024,N_27984,N_27827);
nor U28025 (N_28025,N_27727,N_27669);
or U28026 (N_28026,N_27980,N_27704);
nand U28027 (N_28027,N_27868,N_27647);
xnor U28028 (N_28028,N_27612,N_27728);
nor U28029 (N_28029,N_27977,N_27594);
and U28030 (N_28030,N_27583,N_27967);
and U28031 (N_28031,N_27849,N_27530);
and U28032 (N_28032,N_27667,N_27914);
nor U28033 (N_28033,N_27759,N_27574);
and U28034 (N_28034,N_27693,N_27812);
and U28035 (N_28035,N_27746,N_27834);
and U28036 (N_28036,N_27653,N_27640);
nand U28037 (N_28037,N_27998,N_27754);
nor U28038 (N_28038,N_27744,N_27521);
nor U28039 (N_28039,N_27515,N_27687);
nand U28040 (N_28040,N_27549,N_27858);
xor U28041 (N_28041,N_27586,N_27531);
nand U28042 (N_28042,N_27616,N_27720);
nand U28043 (N_28043,N_27663,N_27872);
nand U28044 (N_28044,N_27802,N_27860);
or U28045 (N_28045,N_27790,N_27865);
and U28046 (N_28046,N_27898,N_27657);
nor U28047 (N_28047,N_27717,N_27902);
nand U28048 (N_28048,N_27569,N_27859);
and U28049 (N_28049,N_27996,N_27761);
and U28050 (N_28050,N_27507,N_27792);
xor U28051 (N_28051,N_27679,N_27893);
xor U28052 (N_28052,N_27678,N_27840);
nor U28053 (N_28053,N_27969,N_27879);
nand U28054 (N_28054,N_27970,N_27796);
or U28055 (N_28055,N_27732,N_27781);
nand U28056 (N_28056,N_27501,N_27993);
or U28057 (N_28057,N_27715,N_27899);
xnor U28058 (N_28058,N_27987,N_27536);
nand U28059 (N_28059,N_27808,N_27972);
or U28060 (N_28060,N_27787,N_27511);
xnor U28061 (N_28061,N_27798,N_27836);
nor U28062 (N_28062,N_27825,N_27828);
and U28063 (N_28063,N_27905,N_27694);
xnor U28064 (N_28064,N_27757,N_27648);
nor U28065 (N_28065,N_27528,N_27935);
nor U28066 (N_28066,N_27947,N_27934);
or U28067 (N_28067,N_27570,N_27512);
and U28068 (N_28068,N_27791,N_27949);
or U28069 (N_28069,N_27961,N_27901);
or U28070 (N_28070,N_27591,N_27801);
nor U28071 (N_28071,N_27617,N_27795);
or U28072 (N_28072,N_27862,N_27964);
and U28073 (N_28073,N_27696,N_27821);
and U28074 (N_28074,N_27803,N_27623);
and U28075 (N_28075,N_27700,N_27505);
nor U28076 (N_28076,N_27844,N_27765);
or U28077 (N_28077,N_27846,N_27655);
or U28078 (N_28078,N_27597,N_27764);
xor U28079 (N_28079,N_27742,N_27785);
and U28080 (N_28080,N_27940,N_27881);
nor U28081 (N_28081,N_27670,N_27595);
nor U28082 (N_28082,N_27659,N_27867);
and U28083 (N_28083,N_27558,N_27843);
xor U28084 (N_28084,N_27854,N_27890);
xnor U28085 (N_28085,N_27788,N_27939);
xor U28086 (N_28086,N_27882,N_27776);
xnor U28087 (N_28087,N_27955,N_27572);
nand U28088 (N_28088,N_27811,N_27891);
nor U28089 (N_28089,N_27907,N_27580);
or U28090 (N_28090,N_27800,N_27887);
xor U28091 (N_28091,N_27943,N_27926);
nor U28092 (N_28092,N_27622,N_27629);
and U28093 (N_28093,N_27645,N_27513);
nor U28094 (N_28094,N_27701,N_27504);
and U28095 (N_28095,N_27774,N_27542);
nor U28096 (N_28096,N_27639,N_27824);
and U28097 (N_28097,N_27749,N_27771);
nand U28098 (N_28098,N_27547,N_27637);
nand U28099 (N_28099,N_27672,N_27799);
and U28100 (N_28100,N_27957,N_27852);
nor U28101 (N_28101,N_27573,N_27724);
nand U28102 (N_28102,N_27668,N_27777);
nand U28103 (N_28103,N_27699,N_27503);
nand U28104 (N_28104,N_27631,N_27673);
nand U28105 (N_28105,N_27689,N_27651);
or U28106 (N_28106,N_27999,N_27649);
xor U28107 (N_28107,N_27750,N_27919);
or U28108 (N_28108,N_27534,N_27927);
nor U28109 (N_28109,N_27676,N_27768);
nand U28110 (N_28110,N_27915,N_27628);
nor U28111 (N_28111,N_27516,N_27677);
xor U28112 (N_28112,N_27609,N_27775);
nor U28113 (N_28113,N_27602,N_27793);
or U28114 (N_28114,N_27756,N_27633);
xor U28115 (N_28115,N_27995,N_27822);
nor U28116 (N_28116,N_27838,N_27835);
or U28117 (N_28117,N_27814,N_27973);
and U28118 (N_28118,N_27912,N_27563);
nor U28119 (N_28119,N_27708,N_27621);
and U28120 (N_28120,N_27666,N_27817);
or U28121 (N_28121,N_27948,N_27864);
nor U28122 (N_28122,N_27662,N_27545);
and U28123 (N_28123,N_27888,N_27751);
xnor U28124 (N_28124,N_27686,N_27705);
xnor U28125 (N_28125,N_27730,N_27786);
xnor U28126 (N_28126,N_27615,N_27894);
nor U28127 (N_28127,N_27951,N_27618);
and U28128 (N_28128,N_27850,N_27620);
and U28129 (N_28129,N_27794,N_27716);
and U28130 (N_28130,N_27833,N_27873);
or U28131 (N_28131,N_27925,N_27630);
or U28132 (N_28132,N_27981,N_27982);
nand U28133 (N_28133,N_27758,N_27945);
nand U28134 (N_28134,N_27675,N_27743);
nor U28135 (N_28135,N_27909,N_27723);
and U28136 (N_28136,N_27692,N_27944);
and U28137 (N_28137,N_27889,N_27635);
nand U28138 (N_28138,N_27941,N_27737);
or U28139 (N_28139,N_27527,N_27729);
or U28140 (N_28140,N_27839,N_27555);
nand U28141 (N_28141,N_27548,N_27520);
xor U28142 (N_28142,N_27762,N_27566);
xnor U28143 (N_28143,N_27992,N_27661);
xor U28144 (N_28144,N_27519,N_27604);
and U28145 (N_28145,N_27634,N_27654);
nor U28146 (N_28146,N_27619,N_27975);
and U28147 (N_28147,N_27924,N_27691);
and U28148 (N_28148,N_27568,N_27643);
nand U28149 (N_28149,N_27928,N_27551);
nand U28150 (N_28150,N_27688,N_27805);
or U28151 (N_28151,N_27613,N_27851);
nand U28152 (N_28152,N_27918,N_27823);
nand U28153 (N_28153,N_27958,N_27582);
and U28154 (N_28154,N_27950,N_27857);
nor U28155 (N_28155,N_27564,N_27848);
or U28156 (N_28156,N_27576,N_27978);
and U28157 (N_28157,N_27884,N_27550);
xnor U28158 (N_28158,N_27789,N_27910);
nor U28159 (N_28159,N_27739,N_27514);
xnor U28160 (N_28160,N_27540,N_27638);
or U28161 (N_28161,N_27718,N_27900);
and U28162 (N_28162,N_27554,N_27610);
xnor U28163 (N_28163,N_27606,N_27946);
nand U28164 (N_28164,N_27702,N_27760);
xor U28165 (N_28165,N_27763,N_27713);
nor U28166 (N_28166,N_27681,N_27665);
nand U28167 (N_28167,N_27997,N_27697);
and U28168 (N_28168,N_27797,N_27736);
and U28169 (N_28169,N_27880,N_27952);
nor U28170 (N_28170,N_27674,N_27562);
and U28171 (N_28171,N_27636,N_27991);
xnor U28172 (N_28172,N_27842,N_27656);
xnor U28173 (N_28173,N_27897,N_27988);
and U28174 (N_28174,N_27684,N_27913);
xnor U28175 (N_28175,N_27780,N_27537);
and U28176 (N_28176,N_27923,N_27543);
and U28177 (N_28177,N_27876,N_27600);
or U28178 (N_28178,N_27908,N_27845);
nor U28179 (N_28179,N_27577,N_27772);
nand U28180 (N_28180,N_27587,N_27896);
and U28181 (N_28181,N_27954,N_27810);
or U28182 (N_28182,N_27561,N_27575);
or U28183 (N_28183,N_27733,N_27847);
nor U28184 (N_28184,N_27956,N_27714);
xnor U28185 (N_28185,N_27989,N_27962);
and U28186 (N_28186,N_27624,N_27539);
or U28187 (N_28187,N_27917,N_27818);
and U28188 (N_28188,N_27598,N_27592);
and U28189 (N_28189,N_27556,N_27596);
nand U28190 (N_28190,N_27710,N_27646);
and U28191 (N_28191,N_27599,N_27552);
and U28192 (N_28192,N_27960,N_27916);
nand U28193 (N_28193,N_27607,N_27682);
or U28194 (N_28194,N_27741,N_27906);
nand U28195 (N_28195,N_27837,N_27976);
and U28196 (N_28196,N_27932,N_27931);
or U28197 (N_28197,N_27831,N_27869);
nand U28198 (N_28198,N_27990,N_27571);
or U28199 (N_28199,N_27641,N_27625);
and U28200 (N_28200,N_27652,N_27784);
nand U28201 (N_28201,N_27883,N_27747);
nor U28202 (N_28202,N_27506,N_27875);
nor U28203 (N_28203,N_27841,N_27650);
and U28204 (N_28204,N_27632,N_27541);
nand U28205 (N_28205,N_27767,N_27920);
and U28206 (N_28206,N_27535,N_27930);
nand U28207 (N_28207,N_27809,N_27560);
or U28208 (N_28208,N_27644,N_27829);
nor U28209 (N_28209,N_27664,N_27690);
nor U28210 (N_28210,N_27517,N_27522);
nand U28211 (N_28211,N_27755,N_27614);
nand U28212 (N_28212,N_27861,N_27878);
or U28213 (N_28213,N_27698,N_27819);
and U28214 (N_28214,N_27611,N_27922);
or U28215 (N_28215,N_27853,N_27816);
and U28216 (N_28216,N_27593,N_27903);
and U28217 (N_28217,N_27820,N_27740);
nand U28218 (N_28218,N_27518,N_27706);
xnor U28219 (N_28219,N_27936,N_27745);
and U28220 (N_28220,N_27904,N_27581);
xnor U28221 (N_28221,N_27578,N_27559);
nand U28222 (N_28222,N_27510,N_27871);
or U28223 (N_28223,N_27974,N_27778);
and U28224 (N_28224,N_27709,N_27721);
nor U28225 (N_28225,N_27590,N_27738);
and U28226 (N_28226,N_27782,N_27608);
or U28227 (N_28227,N_27779,N_27752);
xor U28228 (N_28228,N_27532,N_27508);
xor U28229 (N_28229,N_27680,N_27585);
and U28230 (N_28230,N_27725,N_27523);
nor U28231 (N_28231,N_27911,N_27766);
xor U28232 (N_28232,N_27804,N_27703);
nor U28233 (N_28233,N_27642,N_27830);
nor U28234 (N_28234,N_27953,N_27929);
nand U28235 (N_28235,N_27895,N_27942);
or U28236 (N_28236,N_27734,N_27965);
nand U28237 (N_28237,N_27735,N_27815);
and U28238 (N_28238,N_27509,N_27544);
and U28239 (N_28239,N_27579,N_27983);
nor U28240 (N_28240,N_27557,N_27553);
or U28241 (N_28241,N_27855,N_27994);
xnor U28242 (N_28242,N_27526,N_27546);
xor U28243 (N_28243,N_27770,N_27525);
nor U28244 (N_28244,N_27783,N_27605);
nand U28245 (N_28245,N_27856,N_27870);
nor U28246 (N_28246,N_27683,N_27533);
nand U28247 (N_28247,N_27885,N_27529);
nor U28248 (N_28248,N_27866,N_27671);
nand U28249 (N_28249,N_27601,N_27658);
xor U28250 (N_28250,N_27612,N_27583);
or U28251 (N_28251,N_27918,N_27843);
nand U28252 (N_28252,N_27852,N_27765);
and U28253 (N_28253,N_27622,N_27634);
and U28254 (N_28254,N_27839,N_27667);
nand U28255 (N_28255,N_27827,N_27739);
and U28256 (N_28256,N_27531,N_27711);
and U28257 (N_28257,N_27589,N_27730);
xor U28258 (N_28258,N_27577,N_27716);
nand U28259 (N_28259,N_27866,N_27934);
nand U28260 (N_28260,N_27906,N_27799);
or U28261 (N_28261,N_27514,N_27789);
nand U28262 (N_28262,N_27701,N_27885);
nand U28263 (N_28263,N_27811,N_27936);
nand U28264 (N_28264,N_27813,N_27872);
xnor U28265 (N_28265,N_27962,N_27773);
or U28266 (N_28266,N_27622,N_27960);
and U28267 (N_28267,N_27857,N_27881);
and U28268 (N_28268,N_27870,N_27524);
or U28269 (N_28269,N_27924,N_27615);
and U28270 (N_28270,N_27577,N_27945);
xnor U28271 (N_28271,N_27873,N_27918);
nand U28272 (N_28272,N_27965,N_27597);
and U28273 (N_28273,N_27618,N_27724);
and U28274 (N_28274,N_27828,N_27576);
or U28275 (N_28275,N_27998,N_27778);
nor U28276 (N_28276,N_27572,N_27857);
xnor U28277 (N_28277,N_27854,N_27677);
and U28278 (N_28278,N_27842,N_27610);
xnor U28279 (N_28279,N_27650,N_27845);
and U28280 (N_28280,N_27677,N_27765);
and U28281 (N_28281,N_27792,N_27664);
and U28282 (N_28282,N_27822,N_27563);
and U28283 (N_28283,N_27646,N_27919);
nand U28284 (N_28284,N_27610,N_27813);
or U28285 (N_28285,N_27624,N_27515);
and U28286 (N_28286,N_27718,N_27583);
and U28287 (N_28287,N_27649,N_27975);
or U28288 (N_28288,N_27874,N_27748);
xor U28289 (N_28289,N_27801,N_27765);
xnor U28290 (N_28290,N_27947,N_27591);
xor U28291 (N_28291,N_27774,N_27951);
xor U28292 (N_28292,N_27874,N_27711);
nand U28293 (N_28293,N_27714,N_27766);
and U28294 (N_28294,N_27644,N_27607);
or U28295 (N_28295,N_27549,N_27582);
nand U28296 (N_28296,N_27815,N_27821);
nand U28297 (N_28297,N_27829,N_27603);
nor U28298 (N_28298,N_27641,N_27998);
xor U28299 (N_28299,N_27701,N_27625);
nor U28300 (N_28300,N_27659,N_27552);
or U28301 (N_28301,N_27515,N_27878);
nand U28302 (N_28302,N_27803,N_27763);
or U28303 (N_28303,N_27691,N_27693);
nand U28304 (N_28304,N_27613,N_27731);
nand U28305 (N_28305,N_27553,N_27727);
or U28306 (N_28306,N_27623,N_27906);
or U28307 (N_28307,N_27552,N_27688);
and U28308 (N_28308,N_27992,N_27526);
and U28309 (N_28309,N_27721,N_27863);
nand U28310 (N_28310,N_27561,N_27589);
xnor U28311 (N_28311,N_27772,N_27615);
nor U28312 (N_28312,N_27736,N_27894);
nand U28313 (N_28313,N_27809,N_27894);
xnor U28314 (N_28314,N_27708,N_27985);
xor U28315 (N_28315,N_27864,N_27759);
nand U28316 (N_28316,N_27777,N_27569);
and U28317 (N_28317,N_27656,N_27925);
nor U28318 (N_28318,N_27894,N_27996);
nor U28319 (N_28319,N_27536,N_27625);
nor U28320 (N_28320,N_27996,N_27805);
xnor U28321 (N_28321,N_27752,N_27844);
nor U28322 (N_28322,N_27813,N_27567);
or U28323 (N_28323,N_27697,N_27758);
and U28324 (N_28324,N_27876,N_27967);
or U28325 (N_28325,N_27989,N_27937);
or U28326 (N_28326,N_27549,N_27631);
or U28327 (N_28327,N_27691,N_27832);
and U28328 (N_28328,N_27595,N_27593);
nand U28329 (N_28329,N_27856,N_27992);
nor U28330 (N_28330,N_27958,N_27643);
and U28331 (N_28331,N_27555,N_27883);
nand U28332 (N_28332,N_27725,N_27612);
and U28333 (N_28333,N_27843,N_27698);
and U28334 (N_28334,N_27823,N_27855);
nand U28335 (N_28335,N_27819,N_27606);
and U28336 (N_28336,N_27853,N_27765);
xnor U28337 (N_28337,N_27541,N_27664);
and U28338 (N_28338,N_27817,N_27748);
or U28339 (N_28339,N_27796,N_27940);
nand U28340 (N_28340,N_27559,N_27685);
nor U28341 (N_28341,N_27837,N_27706);
nand U28342 (N_28342,N_27700,N_27641);
xor U28343 (N_28343,N_27669,N_27742);
nor U28344 (N_28344,N_27907,N_27617);
nor U28345 (N_28345,N_27572,N_27758);
and U28346 (N_28346,N_27659,N_27769);
nor U28347 (N_28347,N_27648,N_27795);
and U28348 (N_28348,N_27663,N_27949);
xor U28349 (N_28349,N_27725,N_27804);
nor U28350 (N_28350,N_27513,N_27531);
or U28351 (N_28351,N_27664,N_27932);
nor U28352 (N_28352,N_27594,N_27750);
nor U28353 (N_28353,N_27976,N_27693);
and U28354 (N_28354,N_27663,N_27642);
or U28355 (N_28355,N_27605,N_27881);
nand U28356 (N_28356,N_27655,N_27500);
and U28357 (N_28357,N_27817,N_27611);
or U28358 (N_28358,N_27977,N_27898);
or U28359 (N_28359,N_27907,N_27734);
nor U28360 (N_28360,N_27581,N_27998);
xor U28361 (N_28361,N_27897,N_27618);
and U28362 (N_28362,N_27544,N_27946);
nand U28363 (N_28363,N_27932,N_27765);
or U28364 (N_28364,N_27562,N_27586);
or U28365 (N_28365,N_27530,N_27867);
nand U28366 (N_28366,N_27880,N_27786);
or U28367 (N_28367,N_27515,N_27815);
nor U28368 (N_28368,N_27579,N_27968);
nand U28369 (N_28369,N_27852,N_27539);
xnor U28370 (N_28370,N_27887,N_27567);
nand U28371 (N_28371,N_27737,N_27847);
or U28372 (N_28372,N_27627,N_27934);
nor U28373 (N_28373,N_27958,N_27692);
xnor U28374 (N_28374,N_27877,N_27895);
and U28375 (N_28375,N_27832,N_27693);
and U28376 (N_28376,N_27697,N_27815);
nand U28377 (N_28377,N_27863,N_27528);
nor U28378 (N_28378,N_27595,N_27513);
nor U28379 (N_28379,N_27923,N_27772);
and U28380 (N_28380,N_27529,N_27683);
nand U28381 (N_28381,N_27835,N_27623);
xnor U28382 (N_28382,N_27647,N_27577);
and U28383 (N_28383,N_27578,N_27719);
nor U28384 (N_28384,N_27697,N_27848);
nor U28385 (N_28385,N_27718,N_27560);
or U28386 (N_28386,N_27873,N_27692);
nor U28387 (N_28387,N_27652,N_27960);
nor U28388 (N_28388,N_27564,N_27824);
nand U28389 (N_28389,N_27912,N_27974);
xor U28390 (N_28390,N_27690,N_27585);
or U28391 (N_28391,N_27791,N_27536);
nor U28392 (N_28392,N_27719,N_27735);
or U28393 (N_28393,N_27973,N_27853);
and U28394 (N_28394,N_27605,N_27880);
nor U28395 (N_28395,N_27572,N_27842);
xor U28396 (N_28396,N_27812,N_27979);
or U28397 (N_28397,N_27831,N_27545);
or U28398 (N_28398,N_27885,N_27976);
and U28399 (N_28399,N_27807,N_27768);
nor U28400 (N_28400,N_27669,N_27832);
and U28401 (N_28401,N_27771,N_27902);
nor U28402 (N_28402,N_27807,N_27797);
and U28403 (N_28403,N_27988,N_27662);
or U28404 (N_28404,N_27734,N_27951);
xor U28405 (N_28405,N_27621,N_27609);
xnor U28406 (N_28406,N_27852,N_27677);
nor U28407 (N_28407,N_27931,N_27785);
nor U28408 (N_28408,N_27554,N_27561);
or U28409 (N_28409,N_27540,N_27578);
or U28410 (N_28410,N_27896,N_27657);
and U28411 (N_28411,N_27875,N_27899);
nor U28412 (N_28412,N_27687,N_27982);
xnor U28413 (N_28413,N_27938,N_27659);
nand U28414 (N_28414,N_27924,N_27559);
or U28415 (N_28415,N_27715,N_27691);
nand U28416 (N_28416,N_27616,N_27577);
and U28417 (N_28417,N_27872,N_27746);
nor U28418 (N_28418,N_27556,N_27868);
nor U28419 (N_28419,N_27737,N_27985);
or U28420 (N_28420,N_27614,N_27851);
xor U28421 (N_28421,N_27571,N_27785);
xnor U28422 (N_28422,N_27974,N_27502);
or U28423 (N_28423,N_27748,N_27621);
and U28424 (N_28424,N_27815,N_27840);
or U28425 (N_28425,N_27712,N_27930);
or U28426 (N_28426,N_27979,N_27953);
and U28427 (N_28427,N_27834,N_27909);
nor U28428 (N_28428,N_27555,N_27845);
and U28429 (N_28429,N_27986,N_27885);
or U28430 (N_28430,N_27535,N_27936);
nand U28431 (N_28431,N_27862,N_27814);
nor U28432 (N_28432,N_27780,N_27774);
nand U28433 (N_28433,N_27880,N_27556);
or U28434 (N_28434,N_27524,N_27574);
nand U28435 (N_28435,N_27628,N_27600);
xor U28436 (N_28436,N_27956,N_27511);
nand U28437 (N_28437,N_27576,N_27905);
or U28438 (N_28438,N_27543,N_27890);
nor U28439 (N_28439,N_27663,N_27925);
nor U28440 (N_28440,N_27555,N_27801);
nor U28441 (N_28441,N_27971,N_27822);
nand U28442 (N_28442,N_27978,N_27648);
and U28443 (N_28443,N_27508,N_27947);
nand U28444 (N_28444,N_27871,N_27782);
xor U28445 (N_28445,N_27860,N_27997);
nor U28446 (N_28446,N_27541,N_27631);
nand U28447 (N_28447,N_27671,N_27567);
nand U28448 (N_28448,N_27653,N_27865);
and U28449 (N_28449,N_27589,N_27580);
and U28450 (N_28450,N_27880,N_27913);
nor U28451 (N_28451,N_27599,N_27505);
and U28452 (N_28452,N_27534,N_27522);
xor U28453 (N_28453,N_27621,N_27883);
nand U28454 (N_28454,N_27553,N_27874);
and U28455 (N_28455,N_27984,N_27531);
and U28456 (N_28456,N_27583,N_27914);
and U28457 (N_28457,N_27973,N_27695);
xor U28458 (N_28458,N_27975,N_27967);
and U28459 (N_28459,N_27620,N_27723);
and U28460 (N_28460,N_27793,N_27884);
nand U28461 (N_28461,N_27765,N_27710);
xnor U28462 (N_28462,N_27848,N_27546);
nand U28463 (N_28463,N_27844,N_27965);
nand U28464 (N_28464,N_27805,N_27640);
and U28465 (N_28465,N_27990,N_27586);
nand U28466 (N_28466,N_27632,N_27582);
or U28467 (N_28467,N_27995,N_27974);
xnor U28468 (N_28468,N_27862,N_27641);
and U28469 (N_28469,N_27886,N_27968);
nor U28470 (N_28470,N_27827,N_27596);
nand U28471 (N_28471,N_27831,N_27551);
nand U28472 (N_28472,N_27503,N_27518);
nor U28473 (N_28473,N_27814,N_27856);
or U28474 (N_28474,N_27665,N_27810);
nand U28475 (N_28475,N_27982,N_27593);
or U28476 (N_28476,N_27569,N_27998);
nor U28477 (N_28477,N_27505,N_27550);
nor U28478 (N_28478,N_27687,N_27570);
or U28479 (N_28479,N_27975,N_27667);
xor U28480 (N_28480,N_27722,N_27593);
nor U28481 (N_28481,N_27534,N_27621);
and U28482 (N_28482,N_27762,N_27503);
nand U28483 (N_28483,N_27557,N_27649);
and U28484 (N_28484,N_27850,N_27580);
xnor U28485 (N_28485,N_27704,N_27738);
nand U28486 (N_28486,N_27593,N_27876);
or U28487 (N_28487,N_27524,N_27700);
xor U28488 (N_28488,N_27812,N_27769);
xor U28489 (N_28489,N_27601,N_27741);
or U28490 (N_28490,N_27672,N_27946);
nand U28491 (N_28491,N_27635,N_27897);
nand U28492 (N_28492,N_27716,N_27938);
xnor U28493 (N_28493,N_27803,N_27774);
and U28494 (N_28494,N_27891,N_27728);
nand U28495 (N_28495,N_27696,N_27584);
xnor U28496 (N_28496,N_27714,N_27945);
nor U28497 (N_28497,N_27936,N_27729);
nor U28498 (N_28498,N_27706,N_27594);
nor U28499 (N_28499,N_27930,N_27874);
and U28500 (N_28500,N_28366,N_28458);
nor U28501 (N_28501,N_28328,N_28130);
or U28502 (N_28502,N_28396,N_28405);
or U28503 (N_28503,N_28377,N_28023);
nor U28504 (N_28504,N_28210,N_28225);
xnor U28505 (N_28505,N_28250,N_28357);
and U28506 (N_28506,N_28362,N_28232);
xnor U28507 (N_28507,N_28339,N_28176);
and U28508 (N_28508,N_28288,N_28149);
nor U28509 (N_28509,N_28172,N_28404);
and U28510 (N_28510,N_28182,N_28429);
and U28511 (N_28511,N_28363,N_28206);
nand U28512 (N_28512,N_28003,N_28056);
or U28513 (N_28513,N_28469,N_28350);
nand U28514 (N_28514,N_28468,N_28212);
or U28515 (N_28515,N_28355,N_28334);
and U28516 (N_28516,N_28122,N_28416);
and U28517 (N_28517,N_28444,N_28422);
nand U28518 (N_28518,N_28125,N_28072);
nand U28519 (N_28519,N_28139,N_28091);
xnor U28520 (N_28520,N_28138,N_28036);
xnor U28521 (N_28521,N_28092,N_28291);
nor U28522 (N_28522,N_28457,N_28034);
nor U28523 (N_28523,N_28059,N_28345);
xor U28524 (N_28524,N_28046,N_28205);
and U28525 (N_28525,N_28017,N_28244);
or U28526 (N_28526,N_28348,N_28367);
and U28527 (N_28527,N_28266,N_28053);
xnor U28528 (N_28528,N_28443,N_28144);
nand U28529 (N_28529,N_28057,N_28229);
xor U28530 (N_28530,N_28301,N_28491);
or U28531 (N_28531,N_28460,N_28148);
xor U28532 (N_28532,N_28465,N_28425);
xor U28533 (N_28533,N_28493,N_28087);
xor U28534 (N_28534,N_28441,N_28195);
xnor U28535 (N_28535,N_28361,N_28251);
xnor U28536 (N_28536,N_28187,N_28451);
xor U28537 (N_28537,N_28253,N_28019);
and U28538 (N_28538,N_28424,N_28159);
or U28539 (N_28539,N_28329,N_28448);
or U28540 (N_28540,N_28015,N_28461);
or U28541 (N_28541,N_28274,N_28263);
nand U28542 (N_28542,N_28304,N_28342);
xnor U28543 (N_28543,N_28242,N_28446);
nor U28544 (N_28544,N_28267,N_28035);
or U28545 (N_28545,N_28260,N_28038);
or U28546 (N_28546,N_28026,N_28165);
or U28547 (N_28547,N_28074,N_28271);
nand U28548 (N_28548,N_28037,N_28438);
xnor U28549 (N_28549,N_28346,N_28449);
and U28550 (N_28550,N_28347,N_28180);
and U28551 (N_28551,N_28277,N_28049);
nand U28552 (N_28552,N_28373,N_28110);
and U28553 (N_28553,N_28333,N_28143);
nor U28554 (N_28554,N_28005,N_28150);
nand U28555 (N_28555,N_28063,N_28492);
and U28556 (N_28556,N_28399,N_28490);
nand U28557 (N_28557,N_28411,N_28439);
xor U28558 (N_28558,N_28482,N_28137);
xnor U28559 (N_28559,N_28410,N_28322);
or U28560 (N_28560,N_28470,N_28007);
or U28561 (N_28561,N_28295,N_28203);
and U28562 (N_28562,N_28016,N_28314);
nand U28563 (N_28563,N_28331,N_28456);
nor U28564 (N_28564,N_28413,N_28069);
or U28565 (N_28565,N_28066,N_28080);
nor U28566 (N_28566,N_28189,N_28450);
and U28567 (N_28567,N_28484,N_28302);
nor U28568 (N_28568,N_28265,N_28483);
xnor U28569 (N_28569,N_28077,N_28305);
nor U28570 (N_28570,N_28055,N_28094);
xnor U28571 (N_28571,N_28300,N_28221);
nand U28572 (N_28572,N_28129,N_28475);
nand U28573 (N_28573,N_28406,N_28382);
or U28574 (N_28574,N_28147,N_28153);
nor U28575 (N_28575,N_28054,N_28374);
nor U28576 (N_28576,N_28254,N_28039);
and U28577 (N_28577,N_28403,N_28481);
xnor U28578 (N_28578,N_28103,N_28376);
xnor U28579 (N_28579,N_28340,N_28123);
nand U28580 (N_28580,N_28272,N_28409);
nand U28581 (N_28581,N_28359,N_28433);
nor U28582 (N_28582,N_28096,N_28194);
or U28583 (N_28583,N_28351,N_28480);
nor U28584 (N_28584,N_28315,N_28435);
or U28585 (N_28585,N_28257,N_28412);
nand U28586 (N_28586,N_28249,N_28157);
xor U28587 (N_28587,N_28207,N_28160);
xnor U28588 (N_28588,N_28204,N_28168);
and U28589 (N_28589,N_28246,N_28112);
nor U28590 (N_28590,N_28486,N_28218);
or U28591 (N_28591,N_28108,N_28190);
xnor U28592 (N_28592,N_28104,N_28415);
nand U28593 (N_28593,N_28240,N_28175);
and U28594 (N_28594,N_28185,N_28418);
nor U28595 (N_28595,N_28372,N_28061);
xor U28596 (N_28596,N_28178,N_28307);
xnor U28597 (N_28597,N_28447,N_28174);
or U28598 (N_28598,N_28317,N_28417);
and U28599 (N_28599,N_28344,N_28320);
nor U28600 (N_28600,N_28073,N_28052);
nor U28601 (N_28601,N_28261,N_28227);
nand U28602 (N_28602,N_28082,N_28191);
or U28603 (N_28603,N_28264,N_28011);
and U28604 (N_28604,N_28025,N_28485);
xnor U28605 (N_28605,N_28497,N_28256);
nand U28606 (N_28606,N_28236,N_28090);
xnor U28607 (N_28607,N_28088,N_28119);
or U28608 (N_28608,N_28155,N_28131);
and U28609 (N_28609,N_28308,N_28152);
and U28610 (N_28610,N_28336,N_28306);
or U28611 (N_28611,N_28310,N_28196);
xor U28612 (N_28612,N_28161,N_28001);
nand U28613 (N_28613,N_28089,N_28276);
and U28614 (N_28614,N_28476,N_28296);
or U28615 (N_28615,N_28245,N_28022);
nand U28616 (N_28616,N_28170,N_28352);
nand U28617 (N_28617,N_28255,N_28494);
or U28618 (N_28618,N_28006,N_28408);
nand U28619 (N_28619,N_28273,N_28316);
nor U28620 (N_28620,N_28378,N_28107);
xor U28621 (N_28621,N_28084,N_28247);
nand U28622 (N_28622,N_28341,N_28142);
nand U28623 (N_28623,N_28078,N_28040);
nand U28624 (N_28624,N_28379,N_28100);
nor U28625 (N_28625,N_28188,N_28120);
nor U28626 (N_28626,N_28311,N_28325);
and U28627 (N_28627,N_28239,N_28321);
xnor U28628 (N_28628,N_28201,N_28028);
xor U28629 (N_28629,N_28070,N_28437);
and U28630 (N_28630,N_28012,N_28395);
and U28631 (N_28631,N_28224,N_28013);
or U28632 (N_28632,N_28309,N_28156);
nand U28633 (N_28633,N_28293,N_28095);
nand U28634 (N_28634,N_28146,N_28222);
or U28635 (N_28635,N_28427,N_28358);
nand U28636 (N_28636,N_28327,N_28031);
or U28637 (N_28637,N_28420,N_28464);
nand U28638 (N_28638,N_28141,N_28402);
nor U28639 (N_28639,N_28047,N_28114);
nor U28640 (N_28640,N_28101,N_28455);
nand U28641 (N_28641,N_28018,N_28062);
or U28642 (N_28642,N_28285,N_28283);
xnor U28643 (N_28643,N_28216,N_28060);
or U28644 (N_28644,N_28208,N_28145);
and U28645 (N_28645,N_28032,N_28217);
or U28646 (N_28646,N_28428,N_28202);
xnor U28647 (N_28647,N_28097,N_28075);
and U28648 (N_28648,N_28380,N_28466);
and U28649 (N_28649,N_28419,N_28050);
and U28650 (N_28650,N_28223,N_28081);
nand U28651 (N_28651,N_28258,N_28279);
xnor U28652 (N_28652,N_28398,N_28076);
nand U28653 (N_28653,N_28241,N_28126);
or U28654 (N_28654,N_28269,N_28431);
or U28655 (N_28655,N_28198,N_28002);
nor U28656 (N_28656,N_28235,N_28467);
xor U28657 (N_28657,N_28167,N_28337);
or U28658 (N_28658,N_28303,N_28238);
xnor U28659 (N_28659,N_28243,N_28323);
or U28660 (N_28660,N_28388,N_28259);
or U28661 (N_28661,N_28275,N_28248);
nor U28662 (N_28662,N_28299,N_28093);
and U28663 (N_28663,N_28421,N_28099);
or U28664 (N_28664,N_28287,N_28389);
nand U28665 (N_28665,N_28171,N_28237);
nor U28666 (N_28666,N_28163,N_28384);
and U28667 (N_28667,N_28370,N_28332);
or U28668 (N_28668,N_28234,N_28252);
or U28669 (N_28669,N_28445,N_28365);
nor U28670 (N_28670,N_28086,N_28043);
or U28671 (N_28671,N_28330,N_28289);
or U28672 (N_28672,N_28133,N_28098);
nor U28673 (N_28673,N_28083,N_28135);
and U28674 (N_28674,N_28262,N_28354);
and U28675 (N_28675,N_28177,N_28008);
or U28676 (N_28676,N_28312,N_28364);
and U28677 (N_28677,N_28215,N_28181);
and U28678 (N_28678,N_28014,N_28488);
nand U28679 (N_28679,N_28220,N_28192);
nor U28680 (N_28680,N_28349,N_28498);
and U28681 (N_28681,N_28106,N_28113);
nand U28682 (N_28682,N_28109,N_28313);
or U28683 (N_28683,N_28211,N_28284);
or U28684 (N_28684,N_28489,N_28118);
and U28685 (N_28685,N_28381,N_28324);
or U28686 (N_28686,N_28290,N_28209);
nor U28687 (N_28687,N_28029,N_28179);
and U28688 (N_28688,N_28154,N_28064);
nand U28689 (N_28689,N_28392,N_28186);
xnor U28690 (N_28690,N_28294,N_28386);
xnor U28691 (N_28691,N_28027,N_28280);
nand U28692 (N_28692,N_28009,N_28436);
nand U28693 (N_28693,N_28442,N_28479);
and U28694 (N_28694,N_28297,N_28430);
or U28695 (N_28695,N_28200,N_28390);
or U28696 (N_28696,N_28463,N_28230);
and U28697 (N_28697,N_28338,N_28105);
nand U28698 (N_28698,N_28454,N_28117);
xor U28699 (N_28699,N_28400,N_28387);
and U28700 (N_28700,N_28169,N_28000);
or U28701 (N_28701,N_28360,N_28136);
or U28702 (N_28702,N_28426,N_28051);
and U28703 (N_28703,N_28048,N_28414);
or U28704 (N_28704,N_28213,N_28199);
or U28705 (N_28705,N_28472,N_28335);
and U28706 (N_28706,N_28397,N_28487);
xnor U28707 (N_28707,N_28401,N_28292);
nand U28708 (N_28708,N_28343,N_28111);
nand U28709 (N_28709,N_28166,N_28124);
nor U28710 (N_28710,N_28383,N_28116);
and U28711 (N_28711,N_28228,N_28024);
nand U28712 (N_28712,N_28067,N_28044);
or U28713 (N_28713,N_28068,N_28440);
and U28714 (N_28714,N_28151,N_28231);
nor U28715 (N_28715,N_28452,N_28173);
nor U28716 (N_28716,N_28197,N_28102);
and U28717 (N_28717,N_28318,N_28371);
or U28718 (N_28718,N_28393,N_28071);
xnor U28719 (N_28719,N_28164,N_28270);
xor U28720 (N_28720,N_28121,N_28010);
or U28721 (N_28721,N_28375,N_28219);
and U28722 (N_28722,N_28319,N_28085);
nand U28723 (N_28723,N_28158,N_28473);
nand U28724 (N_28724,N_28226,N_28282);
xnor U28725 (N_28725,N_28128,N_28021);
nand U28726 (N_28726,N_28368,N_28042);
and U28727 (N_28727,N_28434,N_28281);
nor U28728 (N_28728,N_28115,N_28033);
nand U28729 (N_28729,N_28471,N_28183);
nand U28730 (N_28730,N_28453,N_28020);
or U28731 (N_28731,N_28079,N_28369);
xnor U28732 (N_28732,N_28030,N_28058);
and U28733 (N_28733,N_28499,N_28268);
xor U28734 (N_28734,N_28134,N_28432);
or U28735 (N_28735,N_28385,N_28423);
nand U28736 (N_28736,N_28474,N_28233);
nor U28737 (N_28737,N_28459,N_28041);
nor U28738 (N_28738,N_28407,N_28478);
or U28739 (N_28739,N_28278,N_28298);
or U28740 (N_28740,N_28065,N_28184);
nand U28741 (N_28741,N_28127,N_28286);
nand U28742 (N_28742,N_28214,N_28495);
and U28743 (N_28743,N_28462,N_28356);
nand U28744 (N_28744,N_28394,N_28326);
xor U28745 (N_28745,N_28004,N_28140);
and U28746 (N_28746,N_28496,N_28353);
nand U28747 (N_28747,N_28045,N_28193);
nor U28748 (N_28748,N_28391,N_28132);
nor U28749 (N_28749,N_28477,N_28162);
nand U28750 (N_28750,N_28347,N_28469);
or U28751 (N_28751,N_28378,N_28218);
nand U28752 (N_28752,N_28423,N_28362);
nand U28753 (N_28753,N_28008,N_28445);
or U28754 (N_28754,N_28498,N_28077);
nor U28755 (N_28755,N_28382,N_28460);
and U28756 (N_28756,N_28206,N_28221);
and U28757 (N_28757,N_28430,N_28229);
nor U28758 (N_28758,N_28063,N_28058);
nor U28759 (N_28759,N_28005,N_28293);
nand U28760 (N_28760,N_28185,N_28170);
nor U28761 (N_28761,N_28035,N_28347);
xor U28762 (N_28762,N_28147,N_28163);
or U28763 (N_28763,N_28437,N_28410);
xor U28764 (N_28764,N_28312,N_28463);
nand U28765 (N_28765,N_28059,N_28018);
nand U28766 (N_28766,N_28373,N_28254);
and U28767 (N_28767,N_28392,N_28071);
nor U28768 (N_28768,N_28389,N_28132);
or U28769 (N_28769,N_28469,N_28034);
or U28770 (N_28770,N_28147,N_28427);
nor U28771 (N_28771,N_28374,N_28164);
or U28772 (N_28772,N_28409,N_28325);
xor U28773 (N_28773,N_28164,N_28051);
xor U28774 (N_28774,N_28312,N_28329);
nand U28775 (N_28775,N_28423,N_28104);
or U28776 (N_28776,N_28275,N_28124);
and U28777 (N_28777,N_28349,N_28187);
xnor U28778 (N_28778,N_28148,N_28015);
xnor U28779 (N_28779,N_28333,N_28418);
or U28780 (N_28780,N_28091,N_28299);
or U28781 (N_28781,N_28275,N_28322);
xnor U28782 (N_28782,N_28449,N_28125);
nand U28783 (N_28783,N_28111,N_28434);
nand U28784 (N_28784,N_28007,N_28241);
or U28785 (N_28785,N_28433,N_28230);
xor U28786 (N_28786,N_28078,N_28212);
xor U28787 (N_28787,N_28345,N_28350);
xnor U28788 (N_28788,N_28374,N_28284);
nand U28789 (N_28789,N_28347,N_28449);
nand U28790 (N_28790,N_28191,N_28283);
nor U28791 (N_28791,N_28045,N_28435);
nand U28792 (N_28792,N_28104,N_28347);
xor U28793 (N_28793,N_28213,N_28230);
xor U28794 (N_28794,N_28171,N_28482);
or U28795 (N_28795,N_28263,N_28260);
xor U28796 (N_28796,N_28488,N_28480);
nand U28797 (N_28797,N_28071,N_28118);
or U28798 (N_28798,N_28152,N_28132);
xor U28799 (N_28799,N_28286,N_28041);
xnor U28800 (N_28800,N_28114,N_28031);
or U28801 (N_28801,N_28390,N_28176);
and U28802 (N_28802,N_28188,N_28074);
or U28803 (N_28803,N_28477,N_28272);
nor U28804 (N_28804,N_28119,N_28251);
nand U28805 (N_28805,N_28427,N_28481);
nor U28806 (N_28806,N_28182,N_28183);
or U28807 (N_28807,N_28300,N_28090);
xnor U28808 (N_28808,N_28339,N_28040);
and U28809 (N_28809,N_28152,N_28241);
nand U28810 (N_28810,N_28173,N_28283);
and U28811 (N_28811,N_28265,N_28144);
or U28812 (N_28812,N_28450,N_28111);
nand U28813 (N_28813,N_28241,N_28276);
xor U28814 (N_28814,N_28204,N_28022);
nand U28815 (N_28815,N_28264,N_28050);
and U28816 (N_28816,N_28311,N_28222);
nor U28817 (N_28817,N_28410,N_28032);
or U28818 (N_28818,N_28268,N_28145);
and U28819 (N_28819,N_28259,N_28323);
xnor U28820 (N_28820,N_28173,N_28414);
nand U28821 (N_28821,N_28320,N_28173);
nor U28822 (N_28822,N_28012,N_28481);
and U28823 (N_28823,N_28482,N_28104);
nand U28824 (N_28824,N_28053,N_28227);
nor U28825 (N_28825,N_28314,N_28083);
xnor U28826 (N_28826,N_28401,N_28284);
nand U28827 (N_28827,N_28285,N_28274);
or U28828 (N_28828,N_28285,N_28223);
nand U28829 (N_28829,N_28116,N_28247);
nor U28830 (N_28830,N_28399,N_28487);
and U28831 (N_28831,N_28316,N_28219);
xor U28832 (N_28832,N_28069,N_28310);
xnor U28833 (N_28833,N_28474,N_28423);
or U28834 (N_28834,N_28447,N_28029);
nand U28835 (N_28835,N_28364,N_28331);
xor U28836 (N_28836,N_28301,N_28360);
or U28837 (N_28837,N_28040,N_28182);
nor U28838 (N_28838,N_28414,N_28074);
or U28839 (N_28839,N_28453,N_28137);
nand U28840 (N_28840,N_28256,N_28112);
and U28841 (N_28841,N_28384,N_28431);
nor U28842 (N_28842,N_28137,N_28237);
and U28843 (N_28843,N_28282,N_28141);
xor U28844 (N_28844,N_28431,N_28018);
nand U28845 (N_28845,N_28159,N_28283);
nand U28846 (N_28846,N_28103,N_28188);
and U28847 (N_28847,N_28307,N_28263);
xor U28848 (N_28848,N_28000,N_28122);
nand U28849 (N_28849,N_28322,N_28177);
or U28850 (N_28850,N_28106,N_28311);
or U28851 (N_28851,N_28279,N_28421);
xnor U28852 (N_28852,N_28106,N_28436);
or U28853 (N_28853,N_28180,N_28373);
and U28854 (N_28854,N_28337,N_28009);
nand U28855 (N_28855,N_28485,N_28035);
nand U28856 (N_28856,N_28205,N_28190);
or U28857 (N_28857,N_28407,N_28291);
and U28858 (N_28858,N_28367,N_28329);
xor U28859 (N_28859,N_28000,N_28316);
or U28860 (N_28860,N_28366,N_28126);
or U28861 (N_28861,N_28367,N_28106);
xnor U28862 (N_28862,N_28168,N_28444);
or U28863 (N_28863,N_28443,N_28021);
nor U28864 (N_28864,N_28099,N_28342);
or U28865 (N_28865,N_28159,N_28117);
xnor U28866 (N_28866,N_28398,N_28164);
nor U28867 (N_28867,N_28090,N_28258);
nor U28868 (N_28868,N_28363,N_28320);
nor U28869 (N_28869,N_28215,N_28107);
nand U28870 (N_28870,N_28257,N_28216);
nand U28871 (N_28871,N_28239,N_28386);
xnor U28872 (N_28872,N_28198,N_28301);
and U28873 (N_28873,N_28462,N_28204);
nor U28874 (N_28874,N_28334,N_28250);
nand U28875 (N_28875,N_28485,N_28203);
and U28876 (N_28876,N_28074,N_28439);
nand U28877 (N_28877,N_28451,N_28337);
and U28878 (N_28878,N_28125,N_28444);
or U28879 (N_28879,N_28021,N_28473);
xor U28880 (N_28880,N_28171,N_28140);
nor U28881 (N_28881,N_28384,N_28117);
nand U28882 (N_28882,N_28083,N_28287);
nand U28883 (N_28883,N_28417,N_28439);
xnor U28884 (N_28884,N_28489,N_28238);
xor U28885 (N_28885,N_28198,N_28022);
xor U28886 (N_28886,N_28106,N_28017);
nand U28887 (N_28887,N_28168,N_28209);
nor U28888 (N_28888,N_28310,N_28353);
nor U28889 (N_28889,N_28169,N_28254);
and U28890 (N_28890,N_28144,N_28210);
xor U28891 (N_28891,N_28418,N_28426);
and U28892 (N_28892,N_28349,N_28290);
nand U28893 (N_28893,N_28150,N_28273);
xnor U28894 (N_28894,N_28300,N_28370);
or U28895 (N_28895,N_28178,N_28079);
xor U28896 (N_28896,N_28259,N_28126);
nor U28897 (N_28897,N_28318,N_28029);
xnor U28898 (N_28898,N_28386,N_28174);
nand U28899 (N_28899,N_28170,N_28436);
and U28900 (N_28900,N_28169,N_28155);
or U28901 (N_28901,N_28430,N_28117);
nand U28902 (N_28902,N_28159,N_28086);
nand U28903 (N_28903,N_28243,N_28086);
xnor U28904 (N_28904,N_28107,N_28495);
or U28905 (N_28905,N_28442,N_28125);
xnor U28906 (N_28906,N_28020,N_28392);
and U28907 (N_28907,N_28081,N_28017);
nor U28908 (N_28908,N_28433,N_28206);
and U28909 (N_28909,N_28109,N_28324);
nand U28910 (N_28910,N_28430,N_28349);
xnor U28911 (N_28911,N_28219,N_28200);
nor U28912 (N_28912,N_28319,N_28492);
or U28913 (N_28913,N_28384,N_28255);
and U28914 (N_28914,N_28348,N_28140);
xor U28915 (N_28915,N_28392,N_28459);
nand U28916 (N_28916,N_28241,N_28210);
nor U28917 (N_28917,N_28406,N_28308);
or U28918 (N_28918,N_28236,N_28148);
or U28919 (N_28919,N_28394,N_28106);
or U28920 (N_28920,N_28270,N_28236);
or U28921 (N_28921,N_28113,N_28029);
xnor U28922 (N_28922,N_28089,N_28463);
xor U28923 (N_28923,N_28446,N_28439);
or U28924 (N_28924,N_28151,N_28306);
xnor U28925 (N_28925,N_28176,N_28452);
and U28926 (N_28926,N_28168,N_28036);
or U28927 (N_28927,N_28377,N_28307);
and U28928 (N_28928,N_28236,N_28056);
nand U28929 (N_28929,N_28470,N_28266);
nand U28930 (N_28930,N_28357,N_28256);
and U28931 (N_28931,N_28321,N_28077);
and U28932 (N_28932,N_28214,N_28151);
xor U28933 (N_28933,N_28297,N_28243);
nor U28934 (N_28934,N_28439,N_28174);
nor U28935 (N_28935,N_28496,N_28435);
nand U28936 (N_28936,N_28225,N_28338);
or U28937 (N_28937,N_28230,N_28424);
or U28938 (N_28938,N_28147,N_28412);
and U28939 (N_28939,N_28014,N_28097);
and U28940 (N_28940,N_28476,N_28217);
nor U28941 (N_28941,N_28460,N_28203);
xor U28942 (N_28942,N_28395,N_28299);
nand U28943 (N_28943,N_28163,N_28465);
nand U28944 (N_28944,N_28333,N_28091);
or U28945 (N_28945,N_28042,N_28209);
nor U28946 (N_28946,N_28415,N_28030);
nand U28947 (N_28947,N_28359,N_28017);
or U28948 (N_28948,N_28250,N_28276);
nor U28949 (N_28949,N_28422,N_28015);
nand U28950 (N_28950,N_28322,N_28476);
xnor U28951 (N_28951,N_28354,N_28010);
xnor U28952 (N_28952,N_28275,N_28414);
nor U28953 (N_28953,N_28246,N_28467);
xor U28954 (N_28954,N_28492,N_28405);
xor U28955 (N_28955,N_28419,N_28253);
nor U28956 (N_28956,N_28485,N_28331);
or U28957 (N_28957,N_28021,N_28107);
nand U28958 (N_28958,N_28166,N_28178);
nand U28959 (N_28959,N_28284,N_28077);
xnor U28960 (N_28960,N_28326,N_28287);
or U28961 (N_28961,N_28267,N_28264);
xor U28962 (N_28962,N_28457,N_28320);
nor U28963 (N_28963,N_28167,N_28115);
xnor U28964 (N_28964,N_28146,N_28118);
nand U28965 (N_28965,N_28439,N_28175);
or U28966 (N_28966,N_28241,N_28309);
nand U28967 (N_28967,N_28242,N_28346);
nor U28968 (N_28968,N_28351,N_28145);
or U28969 (N_28969,N_28032,N_28313);
nor U28970 (N_28970,N_28061,N_28072);
and U28971 (N_28971,N_28189,N_28017);
xnor U28972 (N_28972,N_28495,N_28331);
and U28973 (N_28973,N_28324,N_28148);
or U28974 (N_28974,N_28241,N_28451);
nor U28975 (N_28975,N_28424,N_28360);
nor U28976 (N_28976,N_28185,N_28477);
nand U28977 (N_28977,N_28435,N_28121);
nor U28978 (N_28978,N_28320,N_28042);
xnor U28979 (N_28979,N_28020,N_28224);
xnor U28980 (N_28980,N_28497,N_28299);
and U28981 (N_28981,N_28245,N_28070);
nor U28982 (N_28982,N_28127,N_28470);
or U28983 (N_28983,N_28124,N_28242);
or U28984 (N_28984,N_28062,N_28425);
nand U28985 (N_28985,N_28360,N_28312);
and U28986 (N_28986,N_28194,N_28360);
or U28987 (N_28987,N_28141,N_28296);
and U28988 (N_28988,N_28416,N_28485);
or U28989 (N_28989,N_28442,N_28336);
xor U28990 (N_28990,N_28043,N_28449);
nor U28991 (N_28991,N_28125,N_28496);
nand U28992 (N_28992,N_28268,N_28049);
nor U28993 (N_28993,N_28365,N_28292);
nor U28994 (N_28994,N_28330,N_28294);
xnor U28995 (N_28995,N_28472,N_28180);
and U28996 (N_28996,N_28454,N_28056);
and U28997 (N_28997,N_28371,N_28444);
xor U28998 (N_28998,N_28088,N_28359);
or U28999 (N_28999,N_28316,N_28349);
nor U29000 (N_29000,N_28798,N_28676);
and U29001 (N_29001,N_28892,N_28692);
xor U29002 (N_29002,N_28689,N_28940);
xor U29003 (N_29003,N_28702,N_28558);
xnor U29004 (N_29004,N_28752,N_28618);
nand U29005 (N_29005,N_28761,N_28780);
or U29006 (N_29006,N_28590,N_28991);
nand U29007 (N_29007,N_28994,N_28566);
nor U29008 (N_29008,N_28863,N_28685);
nand U29009 (N_29009,N_28833,N_28652);
nand U29010 (N_29010,N_28866,N_28758);
xor U29011 (N_29011,N_28936,N_28946);
xnor U29012 (N_29012,N_28759,N_28934);
xnor U29013 (N_29013,N_28889,N_28912);
and U29014 (N_29014,N_28903,N_28635);
xor U29015 (N_29015,N_28756,N_28552);
xnor U29016 (N_29016,N_28844,N_28596);
nand U29017 (N_29017,N_28589,N_28536);
and U29018 (N_29018,N_28968,N_28710);
and U29019 (N_29019,N_28620,N_28637);
or U29020 (N_29020,N_28954,N_28703);
or U29021 (N_29021,N_28922,N_28755);
nand U29022 (N_29022,N_28721,N_28645);
nand U29023 (N_29023,N_28656,N_28623);
and U29024 (N_29024,N_28582,N_28714);
nor U29025 (N_29025,N_28932,N_28682);
nor U29026 (N_29026,N_28914,N_28664);
nor U29027 (N_29027,N_28666,N_28701);
xor U29028 (N_29028,N_28654,N_28743);
or U29029 (N_29029,N_28622,N_28830);
xor U29030 (N_29030,N_28665,N_28725);
or U29031 (N_29031,N_28537,N_28799);
nand U29032 (N_29032,N_28748,N_28807);
nor U29033 (N_29033,N_28942,N_28996);
nor U29034 (N_29034,N_28926,N_28823);
or U29035 (N_29035,N_28675,N_28777);
or U29036 (N_29036,N_28723,N_28834);
or U29037 (N_29037,N_28841,N_28984);
and U29038 (N_29038,N_28624,N_28535);
or U29039 (N_29039,N_28684,N_28772);
nor U29040 (N_29040,N_28514,N_28855);
nor U29041 (N_29041,N_28933,N_28771);
and U29042 (N_29042,N_28906,N_28735);
nor U29043 (N_29043,N_28794,N_28547);
or U29044 (N_29044,N_28894,N_28727);
or U29045 (N_29045,N_28680,N_28976);
nor U29046 (N_29046,N_28592,N_28898);
xor U29047 (N_29047,N_28525,N_28929);
nor U29048 (N_29048,N_28893,N_28661);
nand U29049 (N_29049,N_28507,N_28532);
xnor U29050 (N_29050,N_28594,N_28631);
nand U29051 (N_29051,N_28850,N_28765);
xnor U29052 (N_29052,N_28699,N_28712);
nor U29053 (N_29053,N_28557,N_28913);
and U29054 (N_29054,N_28987,N_28901);
and U29055 (N_29055,N_28643,N_28533);
nand U29056 (N_29056,N_28817,N_28647);
xnor U29057 (N_29057,N_28904,N_28585);
and U29058 (N_29058,N_28885,N_28639);
or U29059 (N_29059,N_28587,N_28564);
and U29060 (N_29060,N_28909,N_28825);
xnor U29061 (N_29061,N_28999,N_28878);
or U29062 (N_29062,N_28806,N_28831);
or U29063 (N_29063,N_28730,N_28629);
or U29064 (N_29064,N_28952,N_28767);
or U29065 (N_29065,N_28605,N_28981);
xor U29066 (N_29066,N_28697,N_28642);
and U29067 (N_29067,N_28704,N_28808);
nor U29068 (N_29068,N_28548,N_28625);
nor U29069 (N_29069,N_28917,N_28741);
nand U29070 (N_29070,N_28957,N_28737);
or U29071 (N_29071,N_28916,N_28930);
xor U29072 (N_29072,N_28608,N_28854);
and U29073 (N_29073,N_28503,N_28621);
nor U29074 (N_29074,N_28510,N_28687);
nand U29075 (N_29075,N_28869,N_28876);
or U29076 (N_29076,N_28939,N_28674);
nand U29077 (N_29077,N_28638,N_28811);
and U29078 (N_29078,N_28776,N_28978);
nand U29079 (N_29079,N_28879,N_28857);
and U29080 (N_29080,N_28958,N_28973);
and U29081 (N_29081,N_28745,N_28658);
nor U29082 (N_29082,N_28796,N_28989);
xnor U29083 (N_29083,N_28529,N_28789);
xnor U29084 (N_29084,N_28560,N_28865);
and U29085 (N_29085,N_28667,N_28516);
or U29086 (N_29086,N_28709,N_28500);
xor U29087 (N_29087,N_28531,N_28734);
or U29088 (N_29088,N_28693,N_28905);
or U29089 (N_29089,N_28983,N_28848);
xnor U29090 (N_29090,N_28845,N_28925);
xor U29091 (N_29091,N_28688,N_28574);
xnor U29092 (N_29092,N_28569,N_28736);
xnor U29093 (N_29093,N_28524,N_28839);
nor U29094 (N_29094,N_28706,N_28899);
and U29095 (N_29095,N_28584,N_28657);
nand U29096 (N_29096,N_28813,N_28617);
xor U29097 (N_29097,N_28815,N_28610);
and U29098 (N_29098,N_28801,N_28722);
nor U29099 (N_29099,N_28502,N_28511);
nor U29100 (N_29100,N_28633,N_28570);
xor U29101 (N_29101,N_28953,N_28613);
and U29102 (N_29102,N_28632,N_28578);
and U29103 (N_29103,N_28821,N_28542);
nor U29104 (N_29104,N_28970,N_28985);
or U29105 (N_29105,N_28612,N_28944);
or U29106 (N_29106,N_28543,N_28738);
xnor U29107 (N_29107,N_28782,N_28672);
nor U29108 (N_29108,N_28718,N_28960);
or U29109 (N_29109,N_28711,N_28921);
or U29110 (N_29110,N_28764,N_28897);
xnor U29111 (N_29111,N_28856,N_28522);
and U29112 (N_29112,N_28512,N_28849);
and U29113 (N_29113,N_28828,N_28804);
nor U29114 (N_29114,N_28690,N_28572);
and U29115 (N_29115,N_28923,N_28545);
nand U29116 (N_29116,N_28986,N_28716);
nand U29117 (N_29117,N_28660,N_28877);
xnor U29118 (N_29118,N_28998,N_28551);
and U29119 (N_29119,N_28785,N_28950);
or U29120 (N_29120,N_28843,N_28668);
or U29121 (N_29121,N_28619,N_28746);
nand U29122 (N_29122,N_28762,N_28739);
xor U29123 (N_29123,N_28719,N_28644);
and U29124 (N_29124,N_28949,N_28924);
nor U29125 (N_29125,N_28786,N_28908);
and U29126 (N_29126,N_28681,N_28541);
nand U29127 (N_29127,N_28920,N_28546);
and U29128 (N_29128,N_28663,N_28783);
xor U29129 (N_29129,N_28975,N_28852);
or U29130 (N_29130,N_28744,N_28988);
nor U29131 (N_29131,N_28521,N_28567);
and U29132 (N_29132,N_28683,N_28787);
xor U29133 (N_29133,N_28810,N_28861);
nor U29134 (N_29134,N_28581,N_28513);
nor U29135 (N_29135,N_28951,N_28720);
nand U29136 (N_29136,N_28915,N_28945);
or U29137 (N_29137,N_28995,N_28800);
and U29138 (N_29138,N_28784,N_28880);
or U29139 (N_29139,N_28858,N_28506);
and U29140 (N_29140,N_28943,N_28881);
and U29141 (N_29141,N_28593,N_28606);
or U29142 (N_29142,N_28768,N_28565);
and U29143 (N_29143,N_28760,N_28576);
nand U29144 (N_29144,N_28646,N_28544);
and U29145 (N_29145,N_28947,N_28814);
xor U29146 (N_29146,N_28538,N_28648);
nand U29147 (N_29147,N_28824,N_28829);
and U29148 (N_29148,N_28636,N_28971);
nand U29149 (N_29149,N_28550,N_28846);
and U29150 (N_29150,N_28963,N_28583);
nand U29151 (N_29151,N_28819,N_28747);
or U29152 (N_29152,N_28911,N_28607);
and U29153 (N_29153,N_28563,N_28882);
nand U29154 (N_29154,N_28707,N_28650);
and U29155 (N_29155,N_28937,N_28599);
nor U29156 (N_29156,N_28559,N_28526);
xor U29157 (N_29157,N_28705,N_28571);
or U29158 (N_29158,N_28775,N_28540);
or U29159 (N_29159,N_28790,N_28523);
and U29160 (N_29160,N_28517,N_28867);
nand U29161 (N_29161,N_28895,N_28888);
and U29162 (N_29162,N_28595,N_28980);
xnor U29163 (N_29163,N_28628,N_28910);
nor U29164 (N_29164,N_28669,N_28896);
nor U29165 (N_29165,N_28862,N_28902);
nand U29166 (N_29166,N_28891,N_28577);
nand U29167 (N_29167,N_28508,N_28694);
nand U29168 (N_29168,N_28695,N_28792);
xor U29169 (N_29169,N_28732,N_28842);
and U29170 (N_29170,N_28713,N_28630);
xnor U29171 (N_29171,N_28729,N_28700);
xor U29172 (N_29172,N_28774,N_28769);
or U29173 (N_29173,N_28698,N_28974);
nor U29174 (N_29174,N_28653,N_28634);
xnor U29175 (N_29175,N_28586,N_28555);
nand U29176 (N_29176,N_28860,N_28982);
and U29177 (N_29177,N_28549,N_28561);
nor U29178 (N_29178,N_28686,N_28822);
or U29179 (N_29179,N_28836,N_28626);
nand U29180 (N_29180,N_28853,N_28871);
nand U29181 (N_29181,N_28740,N_28795);
nor U29182 (N_29182,N_28731,N_28805);
nor U29183 (N_29183,N_28875,N_28670);
nand U29184 (N_29184,N_28568,N_28579);
xor U29185 (N_29185,N_28907,N_28931);
and U29186 (N_29186,N_28742,N_28864);
and U29187 (N_29187,N_28791,N_28977);
or U29188 (N_29188,N_28575,N_28553);
nor U29189 (N_29189,N_28649,N_28603);
nand U29190 (N_29190,N_28941,N_28501);
nand U29191 (N_29191,N_28966,N_28874);
nor U29192 (N_29192,N_28770,N_28754);
or U29193 (N_29193,N_28751,N_28997);
or U29194 (N_29194,N_28562,N_28919);
xnor U29195 (N_29195,N_28873,N_28886);
nor U29196 (N_29196,N_28588,N_28655);
nand U29197 (N_29197,N_28859,N_28802);
or U29198 (N_29198,N_28696,N_28509);
nand U29199 (N_29199,N_28827,N_28868);
and U29200 (N_29200,N_28956,N_28763);
xor U29201 (N_29201,N_28900,N_28749);
nor U29202 (N_29202,N_28872,N_28965);
xor U29203 (N_29203,N_28851,N_28673);
nor U29204 (N_29204,N_28964,N_28993);
nor U29205 (N_29205,N_28773,N_28504);
xor U29206 (N_29206,N_28602,N_28961);
nor U29207 (N_29207,N_28962,N_28708);
nand U29208 (N_29208,N_28539,N_28883);
xnor U29209 (N_29209,N_28935,N_28691);
xnor U29210 (N_29210,N_28724,N_28527);
and U29211 (N_29211,N_28928,N_28679);
nand U29212 (N_29212,N_28651,N_28837);
or U29213 (N_29213,N_28591,N_28990);
xor U29214 (N_29214,N_28573,N_28519);
xnor U29215 (N_29215,N_28884,N_28678);
xor U29216 (N_29216,N_28597,N_28580);
nor U29217 (N_29217,N_28816,N_28518);
nor U29218 (N_29218,N_28781,N_28826);
nand U29219 (N_29219,N_28803,N_28659);
xor U29220 (N_29220,N_28955,N_28753);
xor U29221 (N_29221,N_28609,N_28840);
nor U29222 (N_29222,N_28515,N_28887);
nor U29223 (N_29223,N_28979,N_28788);
xnor U29224 (N_29224,N_28554,N_28757);
nor U29225 (N_29225,N_28534,N_28598);
nor U29226 (N_29226,N_28611,N_28556);
or U29227 (N_29227,N_28671,N_28601);
nand U29228 (N_29228,N_28793,N_28938);
or U29229 (N_29229,N_28847,N_28779);
nor U29230 (N_29230,N_28715,N_28520);
and U29231 (N_29231,N_28835,N_28967);
nor U29232 (N_29232,N_28677,N_28838);
xnor U29233 (N_29233,N_28615,N_28766);
and U29234 (N_29234,N_28528,N_28778);
xnor U29235 (N_29235,N_28616,N_28818);
xnor U29236 (N_29236,N_28728,N_28662);
nor U29237 (N_29237,N_28505,N_28832);
xor U29238 (N_29238,N_28797,N_28733);
nand U29239 (N_29239,N_28809,N_28604);
nand U29240 (N_29240,N_28890,N_28948);
nand U29241 (N_29241,N_28972,N_28870);
or U29242 (N_29242,N_28750,N_28640);
xnor U29243 (N_29243,N_28717,N_28627);
or U29244 (N_29244,N_28641,N_28820);
or U29245 (N_29245,N_28812,N_28918);
xnor U29246 (N_29246,N_28600,N_28530);
xnor U29247 (N_29247,N_28969,N_28992);
xnor U29248 (N_29248,N_28927,N_28614);
or U29249 (N_29249,N_28726,N_28959);
nor U29250 (N_29250,N_28840,N_28823);
xnor U29251 (N_29251,N_28900,N_28718);
or U29252 (N_29252,N_28751,N_28636);
nor U29253 (N_29253,N_28695,N_28894);
or U29254 (N_29254,N_28992,N_28652);
or U29255 (N_29255,N_28986,N_28698);
xnor U29256 (N_29256,N_28885,N_28892);
and U29257 (N_29257,N_28853,N_28600);
and U29258 (N_29258,N_28503,N_28631);
or U29259 (N_29259,N_28851,N_28827);
or U29260 (N_29260,N_28686,N_28805);
and U29261 (N_29261,N_28966,N_28547);
xnor U29262 (N_29262,N_28816,N_28511);
or U29263 (N_29263,N_28922,N_28829);
or U29264 (N_29264,N_28507,N_28851);
xnor U29265 (N_29265,N_28922,N_28595);
or U29266 (N_29266,N_28961,N_28995);
nand U29267 (N_29267,N_28585,N_28741);
nand U29268 (N_29268,N_28780,N_28691);
xnor U29269 (N_29269,N_28645,N_28503);
and U29270 (N_29270,N_28702,N_28600);
nor U29271 (N_29271,N_28572,N_28731);
or U29272 (N_29272,N_28741,N_28908);
or U29273 (N_29273,N_28717,N_28897);
nand U29274 (N_29274,N_28606,N_28581);
and U29275 (N_29275,N_28881,N_28502);
and U29276 (N_29276,N_28818,N_28629);
xnor U29277 (N_29277,N_28837,N_28744);
nand U29278 (N_29278,N_28887,N_28963);
xor U29279 (N_29279,N_28730,N_28787);
nand U29280 (N_29280,N_28684,N_28695);
xor U29281 (N_29281,N_28601,N_28865);
and U29282 (N_29282,N_28533,N_28761);
nor U29283 (N_29283,N_28903,N_28502);
nor U29284 (N_29284,N_28924,N_28896);
xor U29285 (N_29285,N_28991,N_28621);
nand U29286 (N_29286,N_28984,N_28666);
and U29287 (N_29287,N_28513,N_28610);
xnor U29288 (N_29288,N_28519,N_28799);
or U29289 (N_29289,N_28525,N_28504);
or U29290 (N_29290,N_28531,N_28797);
nor U29291 (N_29291,N_28529,N_28642);
xor U29292 (N_29292,N_28938,N_28951);
and U29293 (N_29293,N_28785,N_28786);
nand U29294 (N_29294,N_28998,N_28550);
and U29295 (N_29295,N_28579,N_28832);
or U29296 (N_29296,N_28966,N_28800);
or U29297 (N_29297,N_28772,N_28900);
or U29298 (N_29298,N_28666,N_28513);
xor U29299 (N_29299,N_28672,N_28674);
xor U29300 (N_29300,N_28790,N_28953);
and U29301 (N_29301,N_28543,N_28528);
nor U29302 (N_29302,N_28708,N_28673);
xor U29303 (N_29303,N_28818,N_28986);
xor U29304 (N_29304,N_28764,N_28748);
nor U29305 (N_29305,N_28871,N_28617);
or U29306 (N_29306,N_28597,N_28592);
xor U29307 (N_29307,N_28595,N_28864);
xnor U29308 (N_29308,N_28579,N_28513);
nor U29309 (N_29309,N_28695,N_28699);
nor U29310 (N_29310,N_28747,N_28572);
nand U29311 (N_29311,N_28717,N_28866);
nand U29312 (N_29312,N_28684,N_28997);
nor U29313 (N_29313,N_28595,N_28695);
xor U29314 (N_29314,N_28761,N_28723);
xnor U29315 (N_29315,N_28611,N_28783);
or U29316 (N_29316,N_28765,N_28501);
and U29317 (N_29317,N_28937,N_28649);
and U29318 (N_29318,N_28992,N_28918);
xor U29319 (N_29319,N_28977,N_28560);
or U29320 (N_29320,N_28735,N_28519);
xor U29321 (N_29321,N_28927,N_28732);
nor U29322 (N_29322,N_28536,N_28632);
and U29323 (N_29323,N_28544,N_28936);
and U29324 (N_29324,N_28824,N_28674);
xor U29325 (N_29325,N_28903,N_28646);
and U29326 (N_29326,N_28935,N_28531);
or U29327 (N_29327,N_28503,N_28680);
nor U29328 (N_29328,N_28583,N_28750);
nand U29329 (N_29329,N_28578,N_28793);
nand U29330 (N_29330,N_28516,N_28820);
xor U29331 (N_29331,N_28919,N_28889);
xor U29332 (N_29332,N_28991,N_28547);
or U29333 (N_29333,N_28758,N_28844);
nor U29334 (N_29334,N_28657,N_28895);
and U29335 (N_29335,N_28721,N_28806);
and U29336 (N_29336,N_28860,N_28718);
or U29337 (N_29337,N_28954,N_28912);
nand U29338 (N_29338,N_28858,N_28681);
or U29339 (N_29339,N_28773,N_28598);
and U29340 (N_29340,N_28870,N_28609);
nor U29341 (N_29341,N_28984,N_28505);
and U29342 (N_29342,N_28601,N_28550);
nand U29343 (N_29343,N_28923,N_28555);
xor U29344 (N_29344,N_28876,N_28790);
nor U29345 (N_29345,N_28614,N_28917);
nand U29346 (N_29346,N_28738,N_28984);
nor U29347 (N_29347,N_28993,N_28693);
or U29348 (N_29348,N_28921,N_28668);
or U29349 (N_29349,N_28956,N_28756);
nand U29350 (N_29350,N_28884,N_28642);
or U29351 (N_29351,N_28510,N_28714);
nand U29352 (N_29352,N_28658,N_28990);
nor U29353 (N_29353,N_28820,N_28890);
nand U29354 (N_29354,N_28868,N_28568);
or U29355 (N_29355,N_28614,N_28600);
nand U29356 (N_29356,N_28686,N_28556);
and U29357 (N_29357,N_28633,N_28501);
nor U29358 (N_29358,N_28958,N_28658);
nor U29359 (N_29359,N_28906,N_28891);
or U29360 (N_29360,N_28762,N_28574);
xor U29361 (N_29361,N_28853,N_28585);
or U29362 (N_29362,N_28837,N_28958);
and U29363 (N_29363,N_28758,N_28974);
nand U29364 (N_29364,N_28686,N_28559);
or U29365 (N_29365,N_28738,N_28746);
and U29366 (N_29366,N_28855,N_28734);
xor U29367 (N_29367,N_28794,N_28686);
or U29368 (N_29368,N_28708,N_28525);
nand U29369 (N_29369,N_28768,N_28864);
and U29370 (N_29370,N_28817,N_28529);
and U29371 (N_29371,N_28575,N_28658);
xor U29372 (N_29372,N_28553,N_28636);
nor U29373 (N_29373,N_28861,N_28501);
and U29374 (N_29374,N_28966,N_28595);
or U29375 (N_29375,N_28607,N_28588);
nor U29376 (N_29376,N_28819,N_28919);
and U29377 (N_29377,N_28751,N_28968);
nand U29378 (N_29378,N_28947,N_28500);
nand U29379 (N_29379,N_28778,N_28500);
nor U29380 (N_29380,N_28683,N_28996);
xor U29381 (N_29381,N_28737,N_28601);
nor U29382 (N_29382,N_28868,N_28610);
and U29383 (N_29383,N_28561,N_28904);
xnor U29384 (N_29384,N_28975,N_28910);
nand U29385 (N_29385,N_28984,N_28630);
or U29386 (N_29386,N_28850,N_28782);
nor U29387 (N_29387,N_28643,N_28580);
xnor U29388 (N_29388,N_28989,N_28808);
nor U29389 (N_29389,N_28653,N_28559);
nor U29390 (N_29390,N_28561,N_28675);
xnor U29391 (N_29391,N_28731,N_28754);
nand U29392 (N_29392,N_28862,N_28996);
nand U29393 (N_29393,N_28901,N_28905);
and U29394 (N_29394,N_28828,N_28787);
xor U29395 (N_29395,N_28689,N_28692);
nand U29396 (N_29396,N_28707,N_28644);
or U29397 (N_29397,N_28762,N_28867);
and U29398 (N_29398,N_28936,N_28770);
or U29399 (N_29399,N_28755,N_28916);
or U29400 (N_29400,N_28831,N_28581);
and U29401 (N_29401,N_28761,N_28977);
nand U29402 (N_29402,N_28949,N_28950);
and U29403 (N_29403,N_28942,N_28736);
nor U29404 (N_29404,N_28941,N_28758);
or U29405 (N_29405,N_28955,N_28654);
and U29406 (N_29406,N_28740,N_28610);
nand U29407 (N_29407,N_28917,N_28683);
nor U29408 (N_29408,N_28599,N_28528);
nand U29409 (N_29409,N_28591,N_28954);
xor U29410 (N_29410,N_28572,N_28958);
nor U29411 (N_29411,N_28688,N_28520);
xnor U29412 (N_29412,N_28942,N_28801);
nor U29413 (N_29413,N_28512,N_28539);
nor U29414 (N_29414,N_28909,N_28605);
or U29415 (N_29415,N_28934,N_28913);
and U29416 (N_29416,N_28982,N_28576);
or U29417 (N_29417,N_28906,N_28635);
xor U29418 (N_29418,N_28912,N_28862);
nor U29419 (N_29419,N_28720,N_28576);
or U29420 (N_29420,N_28897,N_28607);
or U29421 (N_29421,N_28950,N_28952);
or U29422 (N_29422,N_28772,N_28663);
nor U29423 (N_29423,N_28613,N_28578);
xnor U29424 (N_29424,N_28545,N_28635);
or U29425 (N_29425,N_28542,N_28509);
nor U29426 (N_29426,N_28826,N_28887);
nand U29427 (N_29427,N_28628,N_28561);
or U29428 (N_29428,N_28966,N_28936);
nand U29429 (N_29429,N_28974,N_28670);
or U29430 (N_29430,N_28571,N_28750);
and U29431 (N_29431,N_28985,N_28654);
nor U29432 (N_29432,N_28546,N_28778);
and U29433 (N_29433,N_28513,N_28938);
nand U29434 (N_29434,N_28728,N_28538);
nand U29435 (N_29435,N_28681,N_28811);
xor U29436 (N_29436,N_28755,N_28946);
or U29437 (N_29437,N_28877,N_28581);
nor U29438 (N_29438,N_28896,N_28629);
or U29439 (N_29439,N_28713,N_28837);
nand U29440 (N_29440,N_28897,N_28589);
or U29441 (N_29441,N_28607,N_28643);
xnor U29442 (N_29442,N_28720,N_28979);
nor U29443 (N_29443,N_28564,N_28606);
xor U29444 (N_29444,N_28859,N_28564);
nand U29445 (N_29445,N_28860,N_28587);
xor U29446 (N_29446,N_28872,N_28754);
xor U29447 (N_29447,N_28901,N_28859);
xor U29448 (N_29448,N_28710,N_28955);
and U29449 (N_29449,N_28612,N_28983);
nand U29450 (N_29450,N_28577,N_28684);
xnor U29451 (N_29451,N_28791,N_28699);
nand U29452 (N_29452,N_28801,N_28851);
xnor U29453 (N_29453,N_28861,N_28759);
nand U29454 (N_29454,N_28775,N_28613);
nand U29455 (N_29455,N_28943,N_28891);
or U29456 (N_29456,N_28580,N_28730);
nor U29457 (N_29457,N_28668,N_28648);
xnor U29458 (N_29458,N_28842,N_28746);
xor U29459 (N_29459,N_28905,N_28558);
or U29460 (N_29460,N_28599,N_28722);
and U29461 (N_29461,N_28551,N_28789);
nand U29462 (N_29462,N_28975,N_28651);
nand U29463 (N_29463,N_28772,N_28686);
nor U29464 (N_29464,N_28956,N_28533);
nor U29465 (N_29465,N_28872,N_28760);
nand U29466 (N_29466,N_28908,N_28645);
nand U29467 (N_29467,N_28527,N_28611);
and U29468 (N_29468,N_28931,N_28761);
nor U29469 (N_29469,N_28597,N_28973);
nor U29470 (N_29470,N_28830,N_28760);
and U29471 (N_29471,N_28764,N_28783);
and U29472 (N_29472,N_28951,N_28645);
or U29473 (N_29473,N_28886,N_28808);
or U29474 (N_29474,N_28939,N_28653);
and U29475 (N_29475,N_28693,N_28785);
xor U29476 (N_29476,N_28903,N_28531);
nand U29477 (N_29477,N_28709,N_28809);
nand U29478 (N_29478,N_28721,N_28789);
or U29479 (N_29479,N_28944,N_28644);
or U29480 (N_29480,N_28616,N_28877);
nor U29481 (N_29481,N_28967,N_28670);
or U29482 (N_29482,N_28884,N_28697);
nor U29483 (N_29483,N_28999,N_28615);
nand U29484 (N_29484,N_28966,N_28796);
xnor U29485 (N_29485,N_28969,N_28645);
xor U29486 (N_29486,N_28520,N_28947);
nor U29487 (N_29487,N_28607,N_28669);
nand U29488 (N_29488,N_28696,N_28794);
and U29489 (N_29489,N_28740,N_28826);
xnor U29490 (N_29490,N_28663,N_28738);
nand U29491 (N_29491,N_28519,N_28705);
xnor U29492 (N_29492,N_28667,N_28656);
or U29493 (N_29493,N_28505,N_28553);
nor U29494 (N_29494,N_28572,N_28591);
nand U29495 (N_29495,N_28689,N_28933);
nand U29496 (N_29496,N_28587,N_28505);
xnor U29497 (N_29497,N_28658,N_28956);
or U29498 (N_29498,N_28668,N_28973);
and U29499 (N_29499,N_28642,N_28621);
or U29500 (N_29500,N_29063,N_29092);
nor U29501 (N_29501,N_29334,N_29126);
and U29502 (N_29502,N_29096,N_29255);
or U29503 (N_29503,N_29475,N_29427);
or U29504 (N_29504,N_29261,N_29323);
and U29505 (N_29505,N_29401,N_29499);
xor U29506 (N_29506,N_29129,N_29367);
and U29507 (N_29507,N_29280,N_29433);
nand U29508 (N_29508,N_29268,N_29185);
and U29509 (N_29509,N_29019,N_29359);
xnor U29510 (N_29510,N_29440,N_29013);
nor U29511 (N_29511,N_29179,N_29118);
and U29512 (N_29512,N_29221,N_29465);
and U29513 (N_29513,N_29365,N_29117);
or U29514 (N_29514,N_29027,N_29387);
nand U29515 (N_29515,N_29032,N_29315);
nor U29516 (N_29516,N_29083,N_29138);
xnor U29517 (N_29517,N_29045,N_29296);
nand U29518 (N_29518,N_29362,N_29090);
nor U29519 (N_29519,N_29428,N_29397);
and U29520 (N_29520,N_29243,N_29189);
xnor U29521 (N_29521,N_29214,N_29360);
nor U29522 (N_29522,N_29158,N_29303);
nand U29523 (N_29523,N_29247,N_29064);
xnor U29524 (N_29524,N_29481,N_29017);
or U29525 (N_29525,N_29014,N_29231);
nand U29526 (N_29526,N_29419,N_29077);
xnor U29527 (N_29527,N_29450,N_29207);
xnor U29528 (N_29528,N_29460,N_29383);
nor U29529 (N_29529,N_29327,N_29155);
and U29530 (N_29530,N_29078,N_29445);
nor U29531 (N_29531,N_29060,N_29372);
and U29532 (N_29532,N_29348,N_29108);
nand U29533 (N_29533,N_29277,N_29335);
nand U29534 (N_29534,N_29251,N_29168);
nor U29535 (N_29535,N_29471,N_29270);
and U29536 (N_29536,N_29125,N_29313);
or U29537 (N_29537,N_29209,N_29180);
xor U29538 (N_29538,N_29321,N_29437);
nand U29539 (N_29539,N_29431,N_29235);
nand U29540 (N_29540,N_29099,N_29438);
nand U29541 (N_29541,N_29153,N_29132);
and U29542 (N_29542,N_29402,N_29012);
or U29543 (N_29543,N_29204,N_29072);
or U29544 (N_29544,N_29210,N_29080);
or U29545 (N_29545,N_29049,N_29495);
and U29546 (N_29546,N_29266,N_29197);
nand U29547 (N_29547,N_29020,N_29089);
xor U29548 (N_29548,N_29349,N_29070);
and U29549 (N_29549,N_29140,N_29496);
nor U29550 (N_29550,N_29016,N_29485);
xor U29551 (N_29551,N_29393,N_29224);
nor U29552 (N_29552,N_29202,N_29291);
xnor U29553 (N_29553,N_29187,N_29008);
nor U29554 (N_29554,N_29418,N_29275);
or U29555 (N_29555,N_29037,N_29347);
nor U29556 (N_29556,N_29423,N_29182);
nand U29557 (N_29557,N_29166,N_29497);
xnor U29558 (N_29558,N_29002,N_29144);
nand U29559 (N_29559,N_29074,N_29075);
xor U29560 (N_29560,N_29452,N_29186);
or U29561 (N_29561,N_29382,N_29119);
or U29562 (N_29562,N_29326,N_29410);
and U29563 (N_29563,N_29441,N_29454);
and U29564 (N_29564,N_29007,N_29175);
or U29565 (N_29565,N_29288,N_29171);
xnor U29566 (N_29566,N_29352,N_29458);
or U29567 (N_29567,N_29198,N_29378);
and U29568 (N_29568,N_29264,N_29426);
nor U29569 (N_29569,N_29102,N_29258);
xor U29570 (N_29570,N_29379,N_29273);
nor U29571 (N_29571,N_29361,N_29082);
nor U29572 (N_29572,N_29287,N_29331);
and U29573 (N_29573,N_29476,N_29105);
nand U29574 (N_29574,N_29031,N_29009);
or U29575 (N_29575,N_29226,N_29054);
or U29576 (N_29576,N_29215,N_29399);
nand U29577 (N_29577,N_29374,N_29286);
xor U29578 (N_29578,N_29306,N_29400);
nor U29579 (N_29579,N_29299,N_29162);
or U29580 (N_29580,N_29191,N_29006);
xnor U29581 (N_29581,N_29241,N_29201);
or U29582 (N_29582,N_29176,N_29429);
xnor U29583 (N_29583,N_29223,N_29135);
nor U29584 (N_29584,N_29003,N_29097);
nand U29585 (N_29585,N_29493,N_29203);
nand U29586 (N_29586,N_29114,N_29274);
xnor U29587 (N_29587,N_29259,N_29024);
nor U29588 (N_29588,N_29281,N_29298);
and U29589 (N_29589,N_29130,N_29356);
or U29590 (N_29590,N_29324,N_29469);
nand U29591 (N_29591,N_29085,N_29473);
and U29592 (N_29592,N_29084,N_29041);
and U29593 (N_29593,N_29477,N_29230);
or U29594 (N_29594,N_29283,N_29449);
nand U29595 (N_29595,N_29489,N_29028);
xnor U29596 (N_29596,N_29244,N_29043);
and U29597 (N_29597,N_29328,N_29302);
xor U29598 (N_29598,N_29381,N_29455);
nor U29599 (N_29599,N_29127,N_29375);
nor U29600 (N_29600,N_29464,N_29325);
or U29601 (N_29601,N_29058,N_29222);
or U29602 (N_29602,N_29341,N_29149);
or U29603 (N_29603,N_29373,N_29122);
and U29604 (N_29604,N_29218,N_29079);
xor U29605 (N_29605,N_29121,N_29404);
nor U29606 (N_29606,N_29459,N_29395);
nor U29607 (N_29607,N_29164,N_29447);
nand U29608 (N_29608,N_29232,N_29333);
xor U29609 (N_29609,N_29053,N_29010);
nand U29610 (N_29610,N_29480,N_29157);
xor U29611 (N_29611,N_29068,N_29434);
and U29612 (N_29612,N_29098,N_29040);
and U29613 (N_29613,N_29322,N_29172);
or U29614 (N_29614,N_29297,N_29152);
xnor U29615 (N_29615,N_29319,N_29026);
xnor U29616 (N_29616,N_29474,N_29448);
nand U29617 (N_29617,N_29301,N_29386);
nand U29618 (N_29618,N_29390,N_29021);
nor U29619 (N_29619,N_29173,N_29227);
nand U29620 (N_29620,N_29069,N_29472);
xor U29621 (N_29621,N_29282,N_29409);
nor U29622 (N_29622,N_29432,N_29190);
nand U29623 (N_29623,N_29005,N_29112);
and U29624 (N_29624,N_29256,N_29042);
and U29625 (N_29625,N_29022,N_29442);
or U29626 (N_29626,N_29110,N_29142);
xor U29627 (N_29627,N_29073,N_29370);
or U29628 (N_29628,N_29205,N_29478);
or U29629 (N_29629,N_29174,N_29345);
nor U29630 (N_29630,N_29113,N_29436);
or U29631 (N_29631,N_29358,N_29482);
or U29632 (N_29632,N_29169,N_29394);
or U29633 (N_29633,N_29194,N_29385);
and U29634 (N_29634,N_29057,N_29470);
and U29635 (N_29635,N_29412,N_29444);
nand U29636 (N_29636,N_29290,N_29030);
and U29637 (N_29637,N_29055,N_29029);
xnor U29638 (N_29638,N_29246,N_29211);
nand U29639 (N_29639,N_29200,N_29311);
nand U29640 (N_29640,N_29219,N_29424);
or U29641 (N_29641,N_29364,N_29406);
or U29642 (N_29642,N_29120,N_29093);
nor U29643 (N_29643,N_29184,N_29160);
and U29644 (N_29644,N_29488,N_29177);
xnor U29645 (N_29645,N_29369,N_29192);
nor U29646 (N_29646,N_29217,N_29001);
nand U29647 (N_29647,N_29446,N_29178);
and U29648 (N_29648,N_29307,N_29498);
or U29649 (N_29649,N_29330,N_29047);
nand U29650 (N_29650,N_29229,N_29106);
nor U29651 (N_29651,N_29407,N_29484);
nor U29652 (N_29652,N_29101,N_29237);
xnor U29653 (N_29653,N_29038,N_29220);
xor U29654 (N_29654,N_29025,N_29111);
nand U29655 (N_29655,N_29276,N_29425);
xor U29656 (N_29656,N_29239,N_29159);
xor U29657 (N_29657,N_29076,N_29107);
and U29658 (N_29658,N_29059,N_29254);
nand U29659 (N_29659,N_29467,N_29388);
nand U29660 (N_29660,N_29094,N_29342);
and U29661 (N_29661,N_29167,N_29145);
or U29662 (N_29662,N_29463,N_29018);
nor U29663 (N_29663,N_29318,N_29320);
nand U29664 (N_29664,N_29134,N_29310);
and U29665 (N_29665,N_29353,N_29462);
nor U29666 (N_29666,N_29284,N_29233);
nor U29667 (N_29667,N_29193,N_29116);
or U29668 (N_29668,N_29143,N_29212);
xnor U29669 (N_29669,N_29216,N_29262);
and U29670 (N_29670,N_29257,N_29421);
or U29671 (N_29671,N_29457,N_29236);
nand U29672 (N_29672,N_29461,N_29343);
nand U29673 (N_29673,N_29136,N_29091);
nor U29674 (N_29674,N_29087,N_29163);
or U29675 (N_29675,N_29357,N_29368);
nor U29676 (N_29676,N_29234,N_29420);
nand U29677 (N_29677,N_29346,N_29435);
nor U29678 (N_29678,N_29036,N_29405);
nand U29679 (N_29679,N_29086,N_29295);
nor U29680 (N_29680,N_29071,N_29278);
nand U29681 (N_29681,N_29249,N_29260);
nor U29682 (N_29682,N_29292,N_29067);
nand U29683 (N_29683,N_29062,N_29023);
nand U29684 (N_29684,N_29156,N_29147);
and U29685 (N_29685,N_29430,N_29240);
and U29686 (N_29686,N_29263,N_29034);
xnor U29687 (N_29687,N_29354,N_29033);
xor U29688 (N_29688,N_29199,N_29490);
and U29689 (N_29689,N_29088,N_29004);
nor U29690 (N_29690,N_29265,N_29225);
nand U29691 (N_29691,N_29384,N_29479);
nand U29692 (N_29692,N_29267,N_29300);
nand U29693 (N_29693,N_29046,N_29279);
xor U29694 (N_29694,N_29170,N_29339);
nor U29695 (N_29695,N_29154,N_29051);
xnor U29696 (N_29696,N_29141,N_29269);
xor U29697 (N_29697,N_29165,N_29123);
or U29698 (N_29698,N_29253,N_29248);
xnor U29699 (N_29699,N_29293,N_29188);
and U29700 (N_29700,N_29408,N_29371);
and U29701 (N_29701,N_29439,N_29208);
xor U29702 (N_29702,N_29415,N_29252);
nand U29703 (N_29703,N_29148,N_29308);
nand U29704 (N_29704,N_29414,N_29411);
and U29705 (N_29705,N_29161,N_29242);
xor U29706 (N_29706,N_29355,N_29317);
xor U29707 (N_29707,N_29304,N_29044);
nand U29708 (N_29708,N_29081,N_29312);
nor U29709 (N_29709,N_29039,N_29139);
or U29710 (N_29710,N_29366,N_29494);
and U29711 (N_29711,N_29396,N_29392);
and U29712 (N_29712,N_29453,N_29103);
nor U29713 (N_29713,N_29289,N_29487);
and U29714 (N_29714,N_29468,N_29316);
or U29715 (N_29715,N_29491,N_29422);
or U29716 (N_29716,N_29150,N_29351);
or U29717 (N_29717,N_29413,N_29398);
and U29718 (N_29718,N_29109,N_29451);
nand U29719 (N_29719,N_29492,N_29128);
nor U29720 (N_29720,N_29115,N_29250);
or U29721 (N_29721,N_29104,N_29146);
nor U29722 (N_29722,N_29213,N_29363);
nand U29723 (N_29723,N_29377,N_29337);
xnor U29724 (N_29724,N_29314,N_29151);
nor U29725 (N_29725,N_29066,N_29336);
xor U29726 (N_29726,N_29309,N_29052);
and U29727 (N_29727,N_29271,N_29011);
nand U29728 (N_29728,N_29181,N_29133);
or U29729 (N_29729,N_29035,N_29206);
nand U29730 (N_29730,N_29338,N_29380);
xor U29731 (N_29731,N_29245,N_29389);
xnor U29732 (N_29732,N_29403,N_29272);
xor U29733 (N_29733,N_29305,N_29350);
xor U29734 (N_29734,N_29095,N_29443);
or U29735 (N_29735,N_29332,N_29376);
nand U29736 (N_29736,N_29416,N_29050);
or U29737 (N_29737,N_29456,N_29228);
or U29738 (N_29738,N_29131,N_29056);
nand U29739 (N_29739,N_29285,N_29100);
and U29740 (N_29740,N_29124,N_29483);
or U29741 (N_29741,N_29137,N_29195);
nand U29742 (N_29742,N_29391,N_29466);
xnor U29743 (N_29743,N_29344,N_29196);
nand U29744 (N_29744,N_29015,N_29294);
nor U29745 (N_29745,N_29329,N_29486);
xnor U29746 (N_29746,N_29061,N_29048);
nand U29747 (N_29747,N_29417,N_29000);
nand U29748 (N_29748,N_29238,N_29183);
xor U29749 (N_29749,N_29340,N_29065);
or U29750 (N_29750,N_29141,N_29099);
xnor U29751 (N_29751,N_29038,N_29118);
and U29752 (N_29752,N_29267,N_29093);
nand U29753 (N_29753,N_29374,N_29015);
or U29754 (N_29754,N_29343,N_29399);
nand U29755 (N_29755,N_29211,N_29340);
nand U29756 (N_29756,N_29119,N_29068);
or U29757 (N_29757,N_29009,N_29423);
nor U29758 (N_29758,N_29352,N_29466);
nand U29759 (N_29759,N_29199,N_29408);
and U29760 (N_29760,N_29295,N_29308);
and U29761 (N_29761,N_29032,N_29158);
and U29762 (N_29762,N_29174,N_29352);
nand U29763 (N_29763,N_29312,N_29477);
or U29764 (N_29764,N_29471,N_29329);
xnor U29765 (N_29765,N_29396,N_29301);
xnor U29766 (N_29766,N_29182,N_29245);
or U29767 (N_29767,N_29286,N_29019);
or U29768 (N_29768,N_29320,N_29024);
and U29769 (N_29769,N_29202,N_29433);
nor U29770 (N_29770,N_29294,N_29234);
nor U29771 (N_29771,N_29481,N_29311);
nand U29772 (N_29772,N_29044,N_29402);
xor U29773 (N_29773,N_29352,N_29173);
nand U29774 (N_29774,N_29381,N_29305);
nor U29775 (N_29775,N_29381,N_29198);
xor U29776 (N_29776,N_29257,N_29358);
nor U29777 (N_29777,N_29417,N_29233);
xnor U29778 (N_29778,N_29154,N_29328);
or U29779 (N_29779,N_29251,N_29231);
nand U29780 (N_29780,N_29180,N_29274);
and U29781 (N_29781,N_29103,N_29147);
and U29782 (N_29782,N_29072,N_29094);
nand U29783 (N_29783,N_29349,N_29257);
or U29784 (N_29784,N_29338,N_29284);
or U29785 (N_29785,N_29183,N_29059);
and U29786 (N_29786,N_29350,N_29359);
and U29787 (N_29787,N_29110,N_29434);
or U29788 (N_29788,N_29390,N_29329);
xnor U29789 (N_29789,N_29342,N_29393);
or U29790 (N_29790,N_29110,N_29018);
and U29791 (N_29791,N_29176,N_29320);
nand U29792 (N_29792,N_29199,N_29422);
xor U29793 (N_29793,N_29487,N_29113);
nand U29794 (N_29794,N_29400,N_29283);
nand U29795 (N_29795,N_29447,N_29044);
nor U29796 (N_29796,N_29236,N_29348);
nor U29797 (N_29797,N_29289,N_29152);
and U29798 (N_29798,N_29497,N_29388);
and U29799 (N_29799,N_29473,N_29042);
or U29800 (N_29800,N_29240,N_29248);
or U29801 (N_29801,N_29000,N_29398);
nand U29802 (N_29802,N_29245,N_29263);
nor U29803 (N_29803,N_29266,N_29081);
xnor U29804 (N_29804,N_29037,N_29268);
and U29805 (N_29805,N_29262,N_29325);
nor U29806 (N_29806,N_29327,N_29237);
or U29807 (N_29807,N_29406,N_29271);
nand U29808 (N_29808,N_29015,N_29391);
or U29809 (N_29809,N_29491,N_29210);
nor U29810 (N_29810,N_29378,N_29112);
nor U29811 (N_29811,N_29057,N_29165);
or U29812 (N_29812,N_29303,N_29237);
xor U29813 (N_29813,N_29019,N_29234);
or U29814 (N_29814,N_29451,N_29146);
and U29815 (N_29815,N_29125,N_29389);
nor U29816 (N_29816,N_29394,N_29050);
nand U29817 (N_29817,N_29396,N_29414);
nor U29818 (N_29818,N_29478,N_29082);
nand U29819 (N_29819,N_29370,N_29102);
nand U29820 (N_29820,N_29415,N_29449);
and U29821 (N_29821,N_29286,N_29465);
nor U29822 (N_29822,N_29036,N_29343);
or U29823 (N_29823,N_29071,N_29244);
or U29824 (N_29824,N_29064,N_29348);
and U29825 (N_29825,N_29411,N_29037);
and U29826 (N_29826,N_29130,N_29312);
xor U29827 (N_29827,N_29261,N_29281);
and U29828 (N_29828,N_29339,N_29011);
or U29829 (N_29829,N_29414,N_29234);
xor U29830 (N_29830,N_29093,N_29062);
or U29831 (N_29831,N_29242,N_29120);
xnor U29832 (N_29832,N_29298,N_29249);
xnor U29833 (N_29833,N_29328,N_29411);
xor U29834 (N_29834,N_29331,N_29204);
xnor U29835 (N_29835,N_29383,N_29176);
nor U29836 (N_29836,N_29457,N_29092);
xnor U29837 (N_29837,N_29495,N_29259);
or U29838 (N_29838,N_29276,N_29389);
xnor U29839 (N_29839,N_29147,N_29215);
and U29840 (N_29840,N_29462,N_29147);
nand U29841 (N_29841,N_29370,N_29455);
xnor U29842 (N_29842,N_29234,N_29263);
or U29843 (N_29843,N_29211,N_29147);
xor U29844 (N_29844,N_29118,N_29012);
nand U29845 (N_29845,N_29291,N_29393);
nor U29846 (N_29846,N_29089,N_29409);
nand U29847 (N_29847,N_29249,N_29308);
xor U29848 (N_29848,N_29495,N_29268);
or U29849 (N_29849,N_29062,N_29301);
nor U29850 (N_29850,N_29116,N_29040);
nand U29851 (N_29851,N_29151,N_29446);
and U29852 (N_29852,N_29343,N_29175);
xor U29853 (N_29853,N_29026,N_29272);
nand U29854 (N_29854,N_29481,N_29001);
xnor U29855 (N_29855,N_29491,N_29124);
or U29856 (N_29856,N_29097,N_29182);
nand U29857 (N_29857,N_29428,N_29466);
nand U29858 (N_29858,N_29161,N_29313);
xnor U29859 (N_29859,N_29345,N_29429);
xor U29860 (N_29860,N_29291,N_29383);
and U29861 (N_29861,N_29025,N_29364);
or U29862 (N_29862,N_29330,N_29467);
xor U29863 (N_29863,N_29472,N_29068);
and U29864 (N_29864,N_29439,N_29431);
nor U29865 (N_29865,N_29195,N_29119);
nor U29866 (N_29866,N_29277,N_29455);
or U29867 (N_29867,N_29417,N_29238);
and U29868 (N_29868,N_29123,N_29041);
nand U29869 (N_29869,N_29156,N_29473);
or U29870 (N_29870,N_29281,N_29486);
nor U29871 (N_29871,N_29057,N_29023);
nor U29872 (N_29872,N_29194,N_29166);
nand U29873 (N_29873,N_29335,N_29138);
and U29874 (N_29874,N_29184,N_29264);
nand U29875 (N_29875,N_29017,N_29030);
and U29876 (N_29876,N_29450,N_29202);
or U29877 (N_29877,N_29316,N_29013);
nor U29878 (N_29878,N_29200,N_29073);
and U29879 (N_29879,N_29264,N_29415);
nand U29880 (N_29880,N_29413,N_29346);
or U29881 (N_29881,N_29075,N_29244);
nor U29882 (N_29882,N_29431,N_29171);
and U29883 (N_29883,N_29486,N_29019);
and U29884 (N_29884,N_29034,N_29436);
or U29885 (N_29885,N_29062,N_29438);
xor U29886 (N_29886,N_29114,N_29120);
or U29887 (N_29887,N_29296,N_29220);
nand U29888 (N_29888,N_29037,N_29412);
nor U29889 (N_29889,N_29359,N_29015);
and U29890 (N_29890,N_29184,N_29239);
nand U29891 (N_29891,N_29487,N_29392);
nor U29892 (N_29892,N_29416,N_29118);
or U29893 (N_29893,N_29361,N_29053);
and U29894 (N_29894,N_29115,N_29239);
or U29895 (N_29895,N_29292,N_29353);
and U29896 (N_29896,N_29451,N_29345);
nor U29897 (N_29897,N_29269,N_29271);
nand U29898 (N_29898,N_29496,N_29290);
nor U29899 (N_29899,N_29443,N_29077);
nor U29900 (N_29900,N_29273,N_29184);
nand U29901 (N_29901,N_29080,N_29493);
xor U29902 (N_29902,N_29392,N_29314);
nand U29903 (N_29903,N_29389,N_29072);
or U29904 (N_29904,N_29026,N_29035);
or U29905 (N_29905,N_29109,N_29089);
or U29906 (N_29906,N_29144,N_29028);
and U29907 (N_29907,N_29262,N_29427);
nand U29908 (N_29908,N_29100,N_29106);
xor U29909 (N_29909,N_29177,N_29480);
xor U29910 (N_29910,N_29394,N_29156);
nand U29911 (N_29911,N_29462,N_29276);
xnor U29912 (N_29912,N_29036,N_29305);
or U29913 (N_29913,N_29069,N_29141);
and U29914 (N_29914,N_29146,N_29065);
and U29915 (N_29915,N_29054,N_29182);
xnor U29916 (N_29916,N_29253,N_29182);
and U29917 (N_29917,N_29471,N_29310);
or U29918 (N_29918,N_29138,N_29207);
and U29919 (N_29919,N_29367,N_29227);
or U29920 (N_29920,N_29459,N_29286);
and U29921 (N_29921,N_29059,N_29000);
nand U29922 (N_29922,N_29400,N_29254);
or U29923 (N_29923,N_29130,N_29259);
or U29924 (N_29924,N_29271,N_29049);
xor U29925 (N_29925,N_29199,N_29102);
or U29926 (N_29926,N_29167,N_29147);
and U29927 (N_29927,N_29128,N_29484);
and U29928 (N_29928,N_29329,N_29073);
xor U29929 (N_29929,N_29113,N_29211);
nor U29930 (N_29930,N_29375,N_29443);
nand U29931 (N_29931,N_29443,N_29441);
nor U29932 (N_29932,N_29392,N_29216);
or U29933 (N_29933,N_29158,N_29430);
and U29934 (N_29934,N_29000,N_29474);
nor U29935 (N_29935,N_29380,N_29126);
xor U29936 (N_29936,N_29460,N_29219);
or U29937 (N_29937,N_29321,N_29145);
nand U29938 (N_29938,N_29370,N_29489);
and U29939 (N_29939,N_29286,N_29104);
or U29940 (N_29940,N_29414,N_29225);
nand U29941 (N_29941,N_29367,N_29360);
and U29942 (N_29942,N_29443,N_29384);
nand U29943 (N_29943,N_29398,N_29179);
nand U29944 (N_29944,N_29244,N_29007);
nor U29945 (N_29945,N_29465,N_29236);
xor U29946 (N_29946,N_29073,N_29004);
xor U29947 (N_29947,N_29450,N_29393);
xnor U29948 (N_29948,N_29043,N_29199);
xor U29949 (N_29949,N_29438,N_29382);
xor U29950 (N_29950,N_29330,N_29044);
or U29951 (N_29951,N_29110,N_29112);
xor U29952 (N_29952,N_29389,N_29075);
nand U29953 (N_29953,N_29254,N_29246);
xor U29954 (N_29954,N_29379,N_29045);
nand U29955 (N_29955,N_29311,N_29233);
or U29956 (N_29956,N_29154,N_29029);
xnor U29957 (N_29957,N_29269,N_29390);
nand U29958 (N_29958,N_29393,N_29002);
nand U29959 (N_29959,N_29008,N_29021);
nand U29960 (N_29960,N_29471,N_29100);
xor U29961 (N_29961,N_29056,N_29486);
nand U29962 (N_29962,N_29418,N_29446);
nand U29963 (N_29963,N_29131,N_29391);
nor U29964 (N_29964,N_29106,N_29145);
or U29965 (N_29965,N_29307,N_29021);
or U29966 (N_29966,N_29002,N_29460);
and U29967 (N_29967,N_29130,N_29429);
and U29968 (N_29968,N_29147,N_29023);
and U29969 (N_29969,N_29429,N_29403);
nor U29970 (N_29970,N_29216,N_29052);
xor U29971 (N_29971,N_29279,N_29338);
xor U29972 (N_29972,N_29337,N_29469);
xor U29973 (N_29973,N_29132,N_29125);
xor U29974 (N_29974,N_29340,N_29119);
nor U29975 (N_29975,N_29430,N_29478);
nand U29976 (N_29976,N_29174,N_29097);
nor U29977 (N_29977,N_29132,N_29494);
nand U29978 (N_29978,N_29119,N_29004);
nand U29979 (N_29979,N_29051,N_29212);
or U29980 (N_29980,N_29257,N_29441);
and U29981 (N_29981,N_29266,N_29427);
xor U29982 (N_29982,N_29147,N_29113);
nand U29983 (N_29983,N_29035,N_29316);
and U29984 (N_29984,N_29136,N_29265);
xnor U29985 (N_29985,N_29465,N_29254);
and U29986 (N_29986,N_29304,N_29352);
xor U29987 (N_29987,N_29497,N_29281);
nor U29988 (N_29988,N_29255,N_29044);
or U29989 (N_29989,N_29428,N_29272);
and U29990 (N_29990,N_29272,N_29333);
xor U29991 (N_29991,N_29006,N_29312);
xor U29992 (N_29992,N_29449,N_29448);
nand U29993 (N_29993,N_29320,N_29003);
and U29994 (N_29994,N_29290,N_29316);
nand U29995 (N_29995,N_29134,N_29321);
nand U29996 (N_29996,N_29102,N_29061);
or U29997 (N_29997,N_29209,N_29030);
and U29998 (N_29998,N_29461,N_29339);
nand U29999 (N_29999,N_29354,N_29190);
xnor UO_0 (O_0,N_29738,N_29612);
or UO_1 (O_1,N_29859,N_29535);
nor UO_2 (O_2,N_29803,N_29812);
or UO_3 (O_3,N_29753,N_29751);
nand UO_4 (O_4,N_29972,N_29629);
and UO_5 (O_5,N_29850,N_29977);
or UO_6 (O_6,N_29871,N_29698);
nor UO_7 (O_7,N_29516,N_29996);
and UO_8 (O_8,N_29860,N_29911);
xor UO_9 (O_9,N_29893,N_29684);
xnor UO_10 (O_10,N_29978,N_29964);
nand UO_11 (O_11,N_29584,N_29603);
nor UO_12 (O_12,N_29739,N_29717);
xnor UO_13 (O_13,N_29890,N_29631);
nor UO_14 (O_14,N_29578,N_29961);
nand UO_15 (O_15,N_29575,N_29724);
xnor UO_16 (O_16,N_29904,N_29615);
xor UO_17 (O_17,N_29866,N_29790);
xnor UO_18 (O_18,N_29597,N_29694);
xor UO_19 (O_19,N_29662,N_29951);
nand UO_20 (O_20,N_29679,N_29619);
or UO_21 (O_21,N_29991,N_29976);
nor UO_22 (O_22,N_29586,N_29755);
and UO_23 (O_23,N_29829,N_29855);
nand UO_24 (O_24,N_29593,N_29775);
or UO_25 (O_25,N_29923,N_29922);
and UO_26 (O_26,N_29820,N_29721);
nand UO_27 (O_27,N_29534,N_29811);
xnor UO_28 (O_28,N_29520,N_29943);
xor UO_29 (O_29,N_29680,N_29710);
and UO_30 (O_30,N_29974,N_29806);
or UO_31 (O_31,N_29725,N_29839);
nand UO_32 (O_32,N_29954,N_29639);
xnor UO_33 (O_33,N_29681,N_29748);
nor UO_34 (O_34,N_29645,N_29881);
nor UO_35 (O_35,N_29814,N_29853);
nand UO_36 (O_36,N_29885,N_29572);
nor UO_37 (O_37,N_29825,N_29709);
xor UO_38 (O_38,N_29703,N_29734);
nand UO_39 (O_39,N_29531,N_29979);
and UO_40 (O_40,N_29997,N_29990);
nor UO_41 (O_41,N_29913,N_29826);
or UO_42 (O_42,N_29616,N_29793);
nand UO_43 (O_43,N_29590,N_29513);
nand UO_44 (O_44,N_29816,N_29833);
xor UO_45 (O_45,N_29547,N_29553);
xor UO_46 (O_46,N_29994,N_29944);
xor UO_47 (O_47,N_29765,N_29921);
and UO_48 (O_48,N_29836,N_29595);
nand UO_49 (O_49,N_29875,N_29898);
nor UO_50 (O_50,N_29948,N_29627);
or UO_51 (O_51,N_29569,N_29562);
nand UO_52 (O_52,N_29526,N_29930);
xnor UO_53 (O_53,N_29903,N_29594);
and UO_54 (O_54,N_29503,N_29696);
nor UO_55 (O_55,N_29564,N_29704);
and UO_56 (O_56,N_29604,N_29532);
and UO_57 (O_57,N_29752,N_29788);
nand UO_58 (O_58,N_29744,N_29888);
and UO_59 (O_59,N_29715,N_29641);
nand UO_60 (O_60,N_29942,N_29524);
and UO_61 (O_61,N_29995,N_29999);
nand UO_62 (O_62,N_29637,N_29653);
nor UO_63 (O_63,N_29813,N_29539);
nor UO_64 (O_64,N_29932,N_29673);
xnor UO_65 (O_65,N_29779,N_29889);
and UO_66 (O_66,N_29545,N_29782);
xnor UO_67 (O_67,N_29591,N_29745);
or UO_68 (O_68,N_29953,N_29892);
or UO_69 (O_69,N_29981,N_29567);
or UO_70 (O_70,N_29638,N_29741);
nand UO_71 (O_71,N_29518,N_29769);
and UO_72 (O_72,N_29529,N_29598);
or UO_73 (O_73,N_29664,N_29986);
nand UO_74 (O_74,N_29621,N_29686);
and UO_75 (O_75,N_29588,N_29606);
xnor UO_76 (O_76,N_29540,N_29750);
and UO_77 (O_77,N_29522,N_29632);
xor UO_78 (O_78,N_29613,N_29822);
nor UO_79 (O_79,N_29708,N_29628);
xnor UO_80 (O_80,N_29570,N_29700);
xnor UO_81 (O_81,N_29963,N_29797);
and UO_82 (O_82,N_29667,N_29644);
and UO_83 (O_83,N_29701,N_29506);
nand UO_84 (O_84,N_29969,N_29998);
nor UO_85 (O_85,N_29831,N_29749);
and UO_86 (O_86,N_29537,N_29754);
and UO_87 (O_87,N_29568,N_29800);
and UO_88 (O_88,N_29899,N_29958);
nand UO_89 (O_89,N_29707,N_29589);
xor UO_90 (O_90,N_29926,N_29722);
or UO_91 (O_91,N_29778,N_29602);
or UO_92 (O_92,N_29933,N_29556);
and UO_93 (O_93,N_29884,N_29935);
nor UO_94 (O_94,N_29659,N_29983);
xnor UO_95 (O_95,N_29852,N_29743);
or UO_96 (O_96,N_29576,N_29843);
xor UO_97 (O_97,N_29785,N_29636);
or UO_98 (O_98,N_29729,N_29834);
and UO_99 (O_99,N_29623,N_29924);
xnor UO_100 (O_100,N_29544,N_29620);
xor UO_101 (O_101,N_29920,N_29574);
or UO_102 (O_102,N_29799,N_29716);
nor UO_103 (O_103,N_29863,N_29625);
nor UO_104 (O_104,N_29695,N_29759);
nand UO_105 (O_105,N_29870,N_29756);
nor UO_106 (O_106,N_29542,N_29740);
or UO_107 (O_107,N_29891,N_29557);
or UO_108 (O_108,N_29563,N_29614);
nand UO_109 (O_109,N_29761,N_29960);
nor UO_110 (O_110,N_29856,N_29561);
xor UO_111 (O_111,N_29762,N_29915);
and UO_112 (O_112,N_29808,N_29987);
and UO_113 (O_113,N_29802,N_29925);
or UO_114 (O_114,N_29643,N_29712);
xor UO_115 (O_115,N_29828,N_29505);
nor UO_116 (O_116,N_29661,N_29742);
nand UO_117 (O_117,N_29810,N_29801);
xor UO_118 (O_118,N_29929,N_29730);
or UO_119 (O_119,N_29838,N_29862);
nor UO_120 (O_120,N_29918,N_29946);
or UO_121 (O_121,N_29883,N_29968);
nand UO_122 (O_122,N_29846,N_29872);
or UO_123 (O_123,N_29880,N_29773);
nand UO_124 (O_124,N_29672,N_29767);
and UO_125 (O_125,N_29804,N_29900);
xor UO_126 (O_126,N_29876,N_29959);
nand UO_127 (O_127,N_29879,N_29611);
and UO_128 (O_128,N_29777,N_29720);
or UO_129 (O_129,N_29650,N_29600);
or UO_130 (O_130,N_29549,N_29731);
nor UO_131 (O_131,N_29757,N_29550);
and UO_132 (O_132,N_29624,N_29508);
xnor UO_133 (O_133,N_29992,N_29633);
or UO_134 (O_134,N_29772,N_29560);
xor UO_135 (O_135,N_29548,N_29565);
xnor UO_136 (O_136,N_29798,N_29649);
and UO_137 (O_137,N_29521,N_29842);
or UO_138 (O_138,N_29583,N_29988);
or UO_139 (O_139,N_29919,N_29693);
or UO_140 (O_140,N_29783,N_29657);
or UO_141 (O_141,N_29683,N_29784);
and UO_142 (O_142,N_29723,N_29847);
and UO_143 (O_143,N_29869,N_29766);
nor UO_144 (O_144,N_29546,N_29663);
nor UO_145 (O_145,N_29573,N_29733);
nor UO_146 (O_146,N_29917,N_29993);
xnor UO_147 (O_147,N_29585,N_29536);
nor UO_148 (O_148,N_29732,N_29654);
xor UO_149 (O_149,N_29705,N_29927);
and UO_150 (O_150,N_29760,N_29849);
or UO_151 (O_151,N_29727,N_29566);
or UO_152 (O_152,N_29776,N_29580);
nand UO_153 (O_153,N_29909,N_29551);
and UO_154 (O_154,N_29507,N_29967);
and UO_155 (O_155,N_29677,N_29817);
xor UO_156 (O_156,N_29905,N_29642);
xor UO_157 (O_157,N_29713,N_29651);
xnor UO_158 (O_158,N_29931,N_29897);
and UO_159 (O_159,N_29970,N_29601);
nor UO_160 (O_160,N_29690,N_29941);
nor UO_161 (O_161,N_29940,N_29971);
nand UO_162 (O_162,N_29796,N_29543);
nand UO_163 (O_163,N_29887,N_29910);
and UO_164 (O_164,N_29854,N_29857);
and UO_165 (O_165,N_29945,N_29780);
xnor UO_166 (O_166,N_29596,N_29554);
nand UO_167 (O_167,N_29688,N_29809);
nor UO_168 (O_168,N_29737,N_29552);
nand UO_169 (O_169,N_29824,N_29699);
xnor UO_170 (O_170,N_29607,N_29671);
nor UO_171 (O_171,N_29848,N_29902);
and UO_172 (O_172,N_29500,N_29538);
xnor UO_173 (O_173,N_29858,N_29840);
and UO_174 (O_174,N_29648,N_29874);
xor UO_175 (O_175,N_29984,N_29658);
nor UO_176 (O_176,N_29559,N_29528);
nor UO_177 (O_177,N_29525,N_29794);
or UO_178 (O_178,N_29726,N_29605);
nor UO_179 (O_179,N_29533,N_29830);
or UO_180 (O_180,N_29515,N_29692);
nor UO_181 (O_181,N_29835,N_29938);
nor UO_182 (O_182,N_29711,N_29787);
nor UO_183 (O_183,N_29735,N_29660);
or UO_184 (O_184,N_29936,N_29914);
nand UO_185 (O_185,N_29952,N_29844);
xnor UO_186 (O_186,N_29510,N_29939);
or UO_187 (O_187,N_29666,N_29610);
nand UO_188 (O_188,N_29511,N_29652);
nand UO_189 (O_189,N_29789,N_29702);
nand UO_190 (O_190,N_29882,N_29973);
or UO_191 (O_191,N_29647,N_29581);
nor UO_192 (O_192,N_29655,N_29541);
xnor UO_193 (O_193,N_29937,N_29634);
and UO_194 (O_194,N_29682,N_29719);
nor UO_195 (O_195,N_29530,N_29736);
or UO_196 (O_196,N_29771,N_29763);
or UO_197 (O_197,N_29706,N_29916);
or UO_198 (O_198,N_29504,N_29747);
or UO_199 (O_199,N_29867,N_29956);
and UO_200 (O_200,N_29906,N_29949);
nand UO_201 (O_201,N_29851,N_29622);
or UO_202 (O_202,N_29823,N_29665);
xor UO_203 (O_203,N_29886,N_29608);
nand UO_204 (O_204,N_29630,N_29635);
nand UO_205 (O_205,N_29728,N_29646);
nor UO_206 (O_206,N_29617,N_29555);
and UO_207 (O_207,N_29865,N_29558);
nor UO_208 (O_208,N_29861,N_29901);
and UO_209 (O_209,N_29571,N_29928);
xor UO_210 (O_210,N_29781,N_29656);
and UO_211 (O_211,N_29807,N_29582);
xor UO_212 (O_212,N_29786,N_29895);
nor UO_213 (O_213,N_29966,N_29609);
or UO_214 (O_214,N_29758,N_29519);
or UO_215 (O_215,N_29815,N_29907);
or UO_216 (O_216,N_29845,N_29989);
nor UO_217 (O_217,N_29502,N_29577);
and UO_218 (O_218,N_29687,N_29896);
nor UO_219 (O_219,N_29832,N_29955);
and UO_220 (O_220,N_29821,N_29965);
nor UO_221 (O_221,N_29873,N_29894);
or UO_222 (O_222,N_29805,N_29975);
xnor UO_223 (O_223,N_29509,N_29697);
xor UO_224 (O_224,N_29746,N_29640);
xor UO_225 (O_225,N_29689,N_29795);
nor UO_226 (O_226,N_29770,N_29934);
and UO_227 (O_227,N_29599,N_29587);
and UO_228 (O_228,N_29980,N_29685);
nand UO_229 (O_229,N_29837,N_29517);
xnor UO_230 (O_230,N_29947,N_29676);
or UO_231 (O_231,N_29864,N_29675);
nor UO_232 (O_232,N_29668,N_29878);
and UO_233 (O_233,N_29512,N_29768);
nor UO_234 (O_234,N_29908,N_29982);
nand UO_235 (O_235,N_29669,N_29774);
nand UO_236 (O_236,N_29691,N_29819);
and UO_237 (O_237,N_29670,N_29957);
and UO_238 (O_238,N_29523,N_29592);
nor UO_239 (O_239,N_29618,N_29912);
nor UO_240 (O_240,N_29674,N_29579);
nand UO_241 (O_241,N_29514,N_29718);
or UO_242 (O_242,N_29962,N_29792);
nor UO_243 (O_243,N_29868,N_29791);
and UO_244 (O_244,N_29714,N_29877);
or UO_245 (O_245,N_29678,N_29841);
nand UO_246 (O_246,N_29527,N_29950);
nand UO_247 (O_247,N_29501,N_29827);
nand UO_248 (O_248,N_29626,N_29985);
nand UO_249 (O_249,N_29818,N_29764);
and UO_250 (O_250,N_29902,N_29604);
or UO_251 (O_251,N_29649,N_29608);
nor UO_252 (O_252,N_29932,N_29735);
and UO_253 (O_253,N_29645,N_29764);
and UO_254 (O_254,N_29883,N_29525);
nand UO_255 (O_255,N_29586,N_29742);
nor UO_256 (O_256,N_29954,N_29761);
xor UO_257 (O_257,N_29815,N_29506);
and UO_258 (O_258,N_29738,N_29862);
nor UO_259 (O_259,N_29677,N_29646);
xnor UO_260 (O_260,N_29887,N_29723);
nand UO_261 (O_261,N_29605,N_29937);
xor UO_262 (O_262,N_29568,N_29586);
nand UO_263 (O_263,N_29713,N_29656);
nor UO_264 (O_264,N_29580,N_29623);
or UO_265 (O_265,N_29635,N_29971);
nor UO_266 (O_266,N_29731,N_29696);
xnor UO_267 (O_267,N_29536,N_29957);
nand UO_268 (O_268,N_29900,N_29541);
xor UO_269 (O_269,N_29760,N_29891);
and UO_270 (O_270,N_29568,N_29505);
nor UO_271 (O_271,N_29784,N_29581);
nor UO_272 (O_272,N_29839,N_29643);
nand UO_273 (O_273,N_29959,N_29693);
nor UO_274 (O_274,N_29639,N_29746);
and UO_275 (O_275,N_29840,N_29905);
nand UO_276 (O_276,N_29715,N_29591);
and UO_277 (O_277,N_29980,N_29865);
and UO_278 (O_278,N_29718,N_29722);
nand UO_279 (O_279,N_29828,N_29575);
nor UO_280 (O_280,N_29561,N_29725);
nand UO_281 (O_281,N_29628,N_29507);
or UO_282 (O_282,N_29554,N_29906);
and UO_283 (O_283,N_29932,N_29800);
nor UO_284 (O_284,N_29692,N_29992);
xnor UO_285 (O_285,N_29583,N_29841);
nor UO_286 (O_286,N_29707,N_29772);
and UO_287 (O_287,N_29748,N_29769);
or UO_288 (O_288,N_29872,N_29557);
nand UO_289 (O_289,N_29512,N_29673);
xor UO_290 (O_290,N_29696,N_29558);
nand UO_291 (O_291,N_29701,N_29791);
nand UO_292 (O_292,N_29612,N_29997);
nor UO_293 (O_293,N_29657,N_29951);
nor UO_294 (O_294,N_29978,N_29658);
or UO_295 (O_295,N_29738,N_29570);
xnor UO_296 (O_296,N_29594,N_29576);
xnor UO_297 (O_297,N_29955,N_29526);
or UO_298 (O_298,N_29709,N_29962);
or UO_299 (O_299,N_29800,N_29818);
or UO_300 (O_300,N_29995,N_29680);
and UO_301 (O_301,N_29870,N_29784);
or UO_302 (O_302,N_29645,N_29852);
or UO_303 (O_303,N_29574,N_29562);
or UO_304 (O_304,N_29889,N_29620);
or UO_305 (O_305,N_29675,N_29772);
xnor UO_306 (O_306,N_29617,N_29822);
and UO_307 (O_307,N_29944,N_29777);
and UO_308 (O_308,N_29570,N_29917);
nor UO_309 (O_309,N_29805,N_29501);
nand UO_310 (O_310,N_29969,N_29940);
and UO_311 (O_311,N_29805,N_29766);
xor UO_312 (O_312,N_29565,N_29946);
and UO_313 (O_313,N_29601,N_29583);
xnor UO_314 (O_314,N_29988,N_29510);
nand UO_315 (O_315,N_29734,N_29656);
nand UO_316 (O_316,N_29896,N_29569);
or UO_317 (O_317,N_29911,N_29987);
xor UO_318 (O_318,N_29826,N_29719);
and UO_319 (O_319,N_29962,N_29502);
xor UO_320 (O_320,N_29709,N_29559);
or UO_321 (O_321,N_29989,N_29680);
nor UO_322 (O_322,N_29547,N_29900);
nand UO_323 (O_323,N_29608,N_29615);
and UO_324 (O_324,N_29538,N_29912);
xor UO_325 (O_325,N_29989,N_29816);
nand UO_326 (O_326,N_29522,N_29603);
nand UO_327 (O_327,N_29942,N_29987);
nand UO_328 (O_328,N_29856,N_29833);
nor UO_329 (O_329,N_29673,N_29548);
or UO_330 (O_330,N_29793,N_29661);
and UO_331 (O_331,N_29589,N_29659);
nor UO_332 (O_332,N_29693,N_29988);
and UO_333 (O_333,N_29745,N_29503);
or UO_334 (O_334,N_29818,N_29868);
nor UO_335 (O_335,N_29603,N_29623);
or UO_336 (O_336,N_29845,N_29804);
or UO_337 (O_337,N_29869,N_29684);
and UO_338 (O_338,N_29782,N_29916);
and UO_339 (O_339,N_29525,N_29679);
nand UO_340 (O_340,N_29996,N_29533);
nand UO_341 (O_341,N_29903,N_29564);
and UO_342 (O_342,N_29628,N_29892);
and UO_343 (O_343,N_29752,N_29775);
nand UO_344 (O_344,N_29964,N_29772);
nor UO_345 (O_345,N_29697,N_29520);
or UO_346 (O_346,N_29766,N_29735);
nand UO_347 (O_347,N_29833,N_29947);
or UO_348 (O_348,N_29881,N_29623);
nand UO_349 (O_349,N_29614,N_29689);
nor UO_350 (O_350,N_29732,N_29906);
nor UO_351 (O_351,N_29519,N_29721);
nor UO_352 (O_352,N_29851,N_29893);
nor UO_353 (O_353,N_29903,N_29662);
nor UO_354 (O_354,N_29905,N_29705);
and UO_355 (O_355,N_29698,N_29640);
or UO_356 (O_356,N_29938,N_29608);
or UO_357 (O_357,N_29615,N_29682);
nand UO_358 (O_358,N_29686,N_29891);
nor UO_359 (O_359,N_29501,N_29982);
or UO_360 (O_360,N_29529,N_29577);
xnor UO_361 (O_361,N_29820,N_29780);
and UO_362 (O_362,N_29732,N_29811);
nor UO_363 (O_363,N_29599,N_29768);
and UO_364 (O_364,N_29778,N_29853);
nor UO_365 (O_365,N_29941,N_29893);
and UO_366 (O_366,N_29953,N_29729);
xnor UO_367 (O_367,N_29922,N_29555);
and UO_368 (O_368,N_29878,N_29655);
xor UO_369 (O_369,N_29912,N_29817);
xor UO_370 (O_370,N_29509,N_29850);
nand UO_371 (O_371,N_29512,N_29677);
nor UO_372 (O_372,N_29907,N_29595);
xor UO_373 (O_373,N_29659,N_29666);
and UO_374 (O_374,N_29586,N_29827);
and UO_375 (O_375,N_29934,N_29549);
nand UO_376 (O_376,N_29782,N_29964);
nor UO_377 (O_377,N_29597,N_29791);
and UO_378 (O_378,N_29682,N_29600);
xnor UO_379 (O_379,N_29757,N_29730);
and UO_380 (O_380,N_29917,N_29836);
and UO_381 (O_381,N_29601,N_29895);
or UO_382 (O_382,N_29747,N_29994);
nor UO_383 (O_383,N_29749,N_29861);
nand UO_384 (O_384,N_29903,N_29598);
nor UO_385 (O_385,N_29575,N_29920);
and UO_386 (O_386,N_29976,N_29975);
nand UO_387 (O_387,N_29869,N_29678);
or UO_388 (O_388,N_29905,N_29676);
nand UO_389 (O_389,N_29898,N_29521);
and UO_390 (O_390,N_29570,N_29725);
nor UO_391 (O_391,N_29980,N_29893);
xor UO_392 (O_392,N_29545,N_29761);
or UO_393 (O_393,N_29847,N_29683);
nor UO_394 (O_394,N_29741,N_29955);
or UO_395 (O_395,N_29750,N_29629);
nand UO_396 (O_396,N_29976,N_29759);
or UO_397 (O_397,N_29831,N_29929);
xnor UO_398 (O_398,N_29787,N_29605);
and UO_399 (O_399,N_29788,N_29635);
nor UO_400 (O_400,N_29853,N_29587);
nor UO_401 (O_401,N_29786,N_29834);
nor UO_402 (O_402,N_29838,N_29827);
or UO_403 (O_403,N_29720,N_29585);
xnor UO_404 (O_404,N_29626,N_29566);
or UO_405 (O_405,N_29520,N_29507);
and UO_406 (O_406,N_29967,N_29538);
and UO_407 (O_407,N_29605,N_29656);
and UO_408 (O_408,N_29589,N_29881);
nand UO_409 (O_409,N_29606,N_29825);
xor UO_410 (O_410,N_29668,N_29722);
and UO_411 (O_411,N_29802,N_29526);
or UO_412 (O_412,N_29524,N_29909);
or UO_413 (O_413,N_29753,N_29857);
nor UO_414 (O_414,N_29750,N_29649);
xnor UO_415 (O_415,N_29562,N_29757);
nor UO_416 (O_416,N_29818,N_29849);
and UO_417 (O_417,N_29997,N_29661);
and UO_418 (O_418,N_29900,N_29578);
xnor UO_419 (O_419,N_29835,N_29965);
and UO_420 (O_420,N_29655,N_29925);
or UO_421 (O_421,N_29906,N_29852);
nor UO_422 (O_422,N_29754,N_29784);
and UO_423 (O_423,N_29855,N_29754);
nor UO_424 (O_424,N_29637,N_29509);
or UO_425 (O_425,N_29771,N_29812);
xor UO_426 (O_426,N_29939,N_29734);
nor UO_427 (O_427,N_29889,N_29604);
xor UO_428 (O_428,N_29805,N_29500);
nor UO_429 (O_429,N_29903,N_29707);
nor UO_430 (O_430,N_29812,N_29974);
nand UO_431 (O_431,N_29814,N_29868);
nand UO_432 (O_432,N_29560,N_29960);
xnor UO_433 (O_433,N_29713,N_29703);
and UO_434 (O_434,N_29806,N_29830);
xor UO_435 (O_435,N_29567,N_29646);
and UO_436 (O_436,N_29866,N_29739);
nor UO_437 (O_437,N_29761,N_29924);
nand UO_438 (O_438,N_29845,N_29876);
xnor UO_439 (O_439,N_29591,N_29764);
or UO_440 (O_440,N_29769,N_29742);
nor UO_441 (O_441,N_29824,N_29996);
or UO_442 (O_442,N_29537,N_29651);
nor UO_443 (O_443,N_29909,N_29561);
or UO_444 (O_444,N_29880,N_29804);
xor UO_445 (O_445,N_29536,N_29670);
or UO_446 (O_446,N_29734,N_29615);
xor UO_447 (O_447,N_29714,N_29648);
nor UO_448 (O_448,N_29568,N_29980);
or UO_449 (O_449,N_29559,N_29550);
nand UO_450 (O_450,N_29928,N_29817);
or UO_451 (O_451,N_29623,N_29886);
and UO_452 (O_452,N_29756,N_29999);
and UO_453 (O_453,N_29652,N_29795);
nor UO_454 (O_454,N_29961,N_29968);
nand UO_455 (O_455,N_29753,N_29822);
nor UO_456 (O_456,N_29788,N_29614);
nand UO_457 (O_457,N_29791,N_29710);
nand UO_458 (O_458,N_29965,N_29782);
nor UO_459 (O_459,N_29731,N_29934);
and UO_460 (O_460,N_29652,N_29550);
nand UO_461 (O_461,N_29876,N_29656);
or UO_462 (O_462,N_29520,N_29745);
nand UO_463 (O_463,N_29811,N_29768);
nand UO_464 (O_464,N_29683,N_29712);
xor UO_465 (O_465,N_29565,N_29561);
nand UO_466 (O_466,N_29543,N_29945);
and UO_467 (O_467,N_29739,N_29782);
or UO_468 (O_468,N_29969,N_29606);
nor UO_469 (O_469,N_29971,N_29520);
or UO_470 (O_470,N_29904,N_29651);
or UO_471 (O_471,N_29799,N_29826);
xor UO_472 (O_472,N_29663,N_29852);
nor UO_473 (O_473,N_29791,N_29549);
nor UO_474 (O_474,N_29760,N_29563);
xnor UO_475 (O_475,N_29890,N_29696);
and UO_476 (O_476,N_29805,N_29624);
or UO_477 (O_477,N_29542,N_29888);
xnor UO_478 (O_478,N_29830,N_29579);
xnor UO_479 (O_479,N_29918,N_29929);
xor UO_480 (O_480,N_29760,N_29907);
xnor UO_481 (O_481,N_29693,N_29680);
or UO_482 (O_482,N_29894,N_29816);
or UO_483 (O_483,N_29737,N_29800);
nor UO_484 (O_484,N_29979,N_29724);
and UO_485 (O_485,N_29592,N_29994);
and UO_486 (O_486,N_29686,N_29748);
and UO_487 (O_487,N_29912,N_29710);
and UO_488 (O_488,N_29554,N_29809);
and UO_489 (O_489,N_29731,N_29694);
nand UO_490 (O_490,N_29836,N_29763);
nor UO_491 (O_491,N_29899,N_29799);
and UO_492 (O_492,N_29644,N_29701);
or UO_493 (O_493,N_29810,N_29553);
xor UO_494 (O_494,N_29655,N_29918);
xor UO_495 (O_495,N_29537,N_29509);
or UO_496 (O_496,N_29911,N_29572);
or UO_497 (O_497,N_29823,N_29856);
and UO_498 (O_498,N_29991,N_29995);
or UO_499 (O_499,N_29506,N_29667);
or UO_500 (O_500,N_29540,N_29827);
nor UO_501 (O_501,N_29830,N_29986);
or UO_502 (O_502,N_29626,N_29841);
or UO_503 (O_503,N_29917,N_29587);
nand UO_504 (O_504,N_29706,N_29737);
nor UO_505 (O_505,N_29896,N_29755);
nor UO_506 (O_506,N_29576,N_29619);
nor UO_507 (O_507,N_29533,N_29548);
and UO_508 (O_508,N_29551,N_29722);
or UO_509 (O_509,N_29903,N_29656);
nor UO_510 (O_510,N_29782,N_29659);
xnor UO_511 (O_511,N_29936,N_29548);
and UO_512 (O_512,N_29624,N_29649);
nand UO_513 (O_513,N_29967,N_29614);
or UO_514 (O_514,N_29868,N_29707);
and UO_515 (O_515,N_29638,N_29721);
xor UO_516 (O_516,N_29967,N_29747);
nor UO_517 (O_517,N_29832,N_29693);
xor UO_518 (O_518,N_29822,N_29872);
xor UO_519 (O_519,N_29815,N_29647);
nor UO_520 (O_520,N_29988,N_29509);
nand UO_521 (O_521,N_29956,N_29913);
or UO_522 (O_522,N_29860,N_29802);
and UO_523 (O_523,N_29828,N_29532);
or UO_524 (O_524,N_29848,N_29628);
nand UO_525 (O_525,N_29607,N_29849);
and UO_526 (O_526,N_29737,N_29909);
nand UO_527 (O_527,N_29985,N_29816);
and UO_528 (O_528,N_29596,N_29834);
or UO_529 (O_529,N_29877,N_29809);
and UO_530 (O_530,N_29809,N_29699);
nor UO_531 (O_531,N_29642,N_29544);
or UO_532 (O_532,N_29999,N_29966);
xnor UO_533 (O_533,N_29888,N_29856);
and UO_534 (O_534,N_29552,N_29720);
and UO_535 (O_535,N_29842,N_29861);
and UO_536 (O_536,N_29901,N_29789);
or UO_537 (O_537,N_29527,N_29520);
and UO_538 (O_538,N_29649,N_29659);
and UO_539 (O_539,N_29980,N_29541);
xor UO_540 (O_540,N_29809,N_29701);
and UO_541 (O_541,N_29754,N_29745);
nor UO_542 (O_542,N_29959,N_29841);
or UO_543 (O_543,N_29529,N_29538);
and UO_544 (O_544,N_29898,N_29691);
xnor UO_545 (O_545,N_29585,N_29577);
or UO_546 (O_546,N_29767,N_29560);
or UO_547 (O_547,N_29858,N_29873);
nor UO_548 (O_548,N_29870,N_29982);
nand UO_549 (O_549,N_29513,N_29890);
and UO_550 (O_550,N_29542,N_29664);
nand UO_551 (O_551,N_29541,N_29528);
nand UO_552 (O_552,N_29775,N_29872);
xor UO_553 (O_553,N_29897,N_29695);
nor UO_554 (O_554,N_29559,N_29958);
nor UO_555 (O_555,N_29939,N_29674);
and UO_556 (O_556,N_29821,N_29751);
and UO_557 (O_557,N_29798,N_29913);
nor UO_558 (O_558,N_29857,N_29579);
and UO_559 (O_559,N_29733,N_29816);
and UO_560 (O_560,N_29506,N_29954);
nor UO_561 (O_561,N_29674,N_29827);
or UO_562 (O_562,N_29996,N_29936);
and UO_563 (O_563,N_29735,N_29970);
or UO_564 (O_564,N_29564,N_29716);
nor UO_565 (O_565,N_29956,N_29978);
or UO_566 (O_566,N_29676,N_29833);
and UO_567 (O_567,N_29757,N_29618);
xnor UO_568 (O_568,N_29513,N_29649);
or UO_569 (O_569,N_29636,N_29543);
or UO_570 (O_570,N_29883,N_29542);
or UO_571 (O_571,N_29896,N_29771);
nor UO_572 (O_572,N_29781,N_29597);
or UO_573 (O_573,N_29741,N_29545);
and UO_574 (O_574,N_29565,N_29542);
or UO_575 (O_575,N_29538,N_29949);
xor UO_576 (O_576,N_29924,N_29897);
nor UO_577 (O_577,N_29913,N_29961);
nand UO_578 (O_578,N_29964,N_29928);
xnor UO_579 (O_579,N_29652,N_29924);
and UO_580 (O_580,N_29503,N_29630);
or UO_581 (O_581,N_29711,N_29666);
and UO_582 (O_582,N_29974,N_29961);
and UO_583 (O_583,N_29874,N_29542);
and UO_584 (O_584,N_29721,N_29883);
and UO_585 (O_585,N_29760,N_29740);
nor UO_586 (O_586,N_29760,N_29518);
xnor UO_587 (O_587,N_29633,N_29843);
xnor UO_588 (O_588,N_29684,N_29842);
nand UO_589 (O_589,N_29515,N_29666);
xor UO_590 (O_590,N_29529,N_29699);
and UO_591 (O_591,N_29871,N_29902);
nand UO_592 (O_592,N_29531,N_29866);
nor UO_593 (O_593,N_29728,N_29630);
xnor UO_594 (O_594,N_29627,N_29730);
xnor UO_595 (O_595,N_29650,N_29624);
or UO_596 (O_596,N_29832,N_29605);
nor UO_597 (O_597,N_29625,N_29640);
xor UO_598 (O_598,N_29505,N_29836);
nand UO_599 (O_599,N_29984,N_29635);
and UO_600 (O_600,N_29842,N_29626);
or UO_601 (O_601,N_29879,N_29835);
nand UO_602 (O_602,N_29870,N_29582);
and UO_603 (O_603,N_29648,N_29573);
or UO_604 (O_604,N_29654,N_29934);
nor UO_605 (O_605,N_29695,N_29855);
and UO_606 (O_606,N_29707,N_29693);
nor UO_607 (O_607,N_29646,N_29687);
nand UO_608 (O_608,N_29970,N_29929);
or UO_609 (O_609,N_29852,N_29693);
and UO_610 (O_610,N_29882,N_29674);
and UO_611 (O_611,N_29983,N_29627);
nor UO_612 (O_612,N_29503,N_29856);
or UO_613 (O_613,N_29523,N_29733);
nand UO_614 (O_614,N_29561,N_29504);
xnor UO_615 (O_615,N_29843,N_29734);
xnor UO_616 (O_616,N_29748,N_29994);
or UO_617 (O_617,N_29979,N_29578);
nor UO_618 (O_618,N_29977,N_29997);
and UO_619 (O_619,N_29661,N_29580);
nand UO_620 (O_620,N_29963,N_29599);
or UO_621 (O_621,N_29769,N_29522);
and UO_622 (O_622,N_29712,N_29566);
and UO_623 (O_623,N_29772,N_29562);
and UO_624 (O_624,N_29692,N_29655);
nor UO_625 (O_625,N_29852,N_29887);
or UO_626 (O_626,N_29712,N_29574);
and UO_627 (O_627,N_29791,N_29612);
xnor UO_628 (O_628,N_29987,N_29526);
or UO_629 (O_629,N_29606,N_29754);
nor UO_630 (O_630,N_29939,N_29611);
and UO_631 (O_631,N_29996,N_29508);
xnor UO_632 (O_632,N_29994,N_29685);
xnor UO_633 (O_633,N_29923,N_29624);
or UO_634 (O_634,N_29909,N_29549);
or UO_635 (O_635,N_29895,N_29742);
and UO_636 (O_636,N_29918,N_29826);
and UO_637 (O_637,N_29943,N_29568);
nand UO_638 (O_638,N_29559,N_29749);
nand UO_639 (O_639,N_29674,N_29857);
nand UO_640 (O_640,N_29891,N_29721);
nor UO_641 (O_641,N_29704,N_29688);
nor UO_642 (O_642,N_29644,N_29957);
nand UO_643 (O_643,N_29625,N_29864);
or UO_644 (O_644,N_29693,N_29759);
xor UO_645 (O_645,N_29992,N_29830);
nand UO_646 (O_646,N_29907,N_29773);
xor UO_647 (O_647,N_29522,N_29550);
nor UO_648 (O_648,N_29798,N_29822);
nor UO_649 (O_649,N_29631,N_29521);
nor UO_650 (O_650,N_29652,N_29685);
or UO_651 (O_651,N_29573,N_29767);
nand UO_652 (O_652,N_29607,N_29815);
nand UO_653 (O_653,N_29646,N_29964);
nand UO_654 (O_654,N_29563,N_29698);
and UO_655 (O_655,N_29854,N_29941);
nand UO_656 (O_656,N_29997,N_29664);
and UO_657 (O_657,N_29834,N_29670);
or UO_658 (O_658,N_29679,N_29805);
and UO_659 (O_659,N_29964,N_29599);
and UO_660 (O_660,N_29672,N_29815);
nor UO_661 (O_661,N_29901,N_29628);
and UO_662 (O_662,N_29876,N_29803);
nand UO_663 (O_663,N_29758,N_29676);
nor UO_664 (O_664,N_29729,N_29704);
or UO_665 (O_665,N_29648,N_29632);
nor UO_666 (O_666,N_29935,N_29860);
and UO_667 (O_667,N_29990,N_29778);
xor UO_668 (O_668,N_29687,N_29530);
nand UO_669 (O_669,N_29741,N_29628);
or UO_670 (O_670,N_29707,N_29508);
xor UO_671 (O_671,N_29975,N_29545);
and UO_672 (O_672,N_29733,N_29644);
nor UO_673 (O_673,N_29542,N_29596);
nand UO_674 (O_674,N_29523,N_29723);
nand UO_675 (O_675,N_29718,N_29961);
and UO_676 (O_676,N_29980,N_29660);
nor UO_677 (O_677,N_29990,N_29583);
nor UO_678 (O_678,N_29965,N_29823);
nor UO_679 (O_679,N_29780,N_29543);
or UO_680 (O_680,N_29824,N_29744);
xor UO_681 (O_681,N_29878,N_29829);
nor UO_682 (O_682,N_29803,N_29565);
and UO_683 (O_683,N_29707,N_29530);
and UO_684 (O_684,N_29809,N_29714);
nand UO_685 (O_685,N_29530,N_29905);
nor UO_686 (O_686,N_29712,N_29803);
or UO_687 (O_687,N_29598,N_29741);
nand UO_688 (O_688,N_29533,N_29867);
nand UO_689 (O_689,N_29604,N_29856);
nand UO_690 (O_690,N_29706,N_29871);
nor UO_691 (O_691,N_29999,N_29660);
and UO_692 (O_692,N_29611,N_29536);
and UO_693 (O_693,N_29524,N_29866);
or UO_694 (O_694,N_29742,N_29943);
nand UO_695 (O_695,N_29781,N_29574);
or UO_696 (O_696,N_29647,N_29743);
nor UO_697 (O_697,N_29535,N_29905);
and UO_698 (O_698,N_29707,N_29777);
or UO_699 (O_699,N_29870,N_29783);
or UO_700 (O_700,N_29820,N_29847);
nand UO_701 (O_701,N_29603,N_29920);
nor UO_702 (O_702,N_29921,N_29633);
nor UO_703 (O_703,N_29921,N_29806);
or UO_704 (O_704,N_29860,N_29628);
and UO_705 (O_705,N_29617,N_29663);
nor UO_706 (O_706,N_29681,N_29521);
nor UO_707 (O_707,N_29998,N_29706);
nand UO_708 (O_708,N_29678,N_29705);
and UO_709 (O_709,N_29908,N_29762);
or UO_710 (O_710,N_29897,N_29818);
and UO_711 (O_711,N_29628,N_29872);
or UO_712 (O_712,N_29830,N_29553);
nand UO_713 (O_713,N_29823,N_29895);
nor UO_714 (O_714,N_29714,N_29906);
xnor UO_715 (O_715,N_29637,N_29518);
nor UO_716 (O_716,N_29834,N_29894);
and UO_717 (O_717,N_29679,N_29977);
nor UO_718 (O_718,N_29657,N_29910);
and UO_719 (O_719,N_29539,N_29927);
or UO_720 (O_720,N_29962,N_29536);
nand UO_721 (O_721,N_29849,N_29533);
or UO_722 (O_722,N_29659,N_29761);
and UO_723 (O_723,N_29860,N_29629);
and UO_724 (O_724,N_29756,N_29615);
xnor UO_725 (O_725,N_29921,N_29507);
and UO_726 (O_726,N_29689,N_29922);
xnor UO_727 (O_727,N_29840,N_29982);
and UO_728 (O_728,N_29935,N_29730);
nor UO_729 (O_729,N_29812,N_29765);
xor UO_730 (O_730,N_29897,N_29777);
xnor UO_731 (O_731,N_29582,N_29521);
nand UO_732 (O_732,N_29508,N_29600);
xnor UO_733 (O_733,N_29581,N_29844);
nand UO_734 (O_734,N_29791,N_29654);
nand UO_735 (O_735,N_29791,N_29796);
and UO_736 (O_736,N_29901,N_29580);
xnor UO_737 (O_737,N_29733,N_29869);
xnor UO_738 (O_738,N_29940,N_29905);
xnor UO_739 (O_739,N_29993,N_29819);
or UO_740 (O_740,N_29867,N_29607);
xor UO_741 (O_741,N_29577,N_29750);
or UO_742 (O_742,N_29690,N_29745);
and UO_743 (O_743,N_29671,N_29717);
and UO_744 (O_744,N_29950,N_29916);
and UO_745 (O_745,N_29700,N_29586);
or UO_746 (O_746,N_29793,N_29856);
nor UO_747 (O_747,N_29774,N_29719);
or UO_748 (O_748,N_29606,N_29891);
xor UO_749 (O_749,N_29610,N_29775);
or UO_750 (O_750,N_29952,N_29594);
xnor UO_751 (O_751,N_29769,N_29855);
nand UO_752 (O_752,N_29950,N_29924);
nand UO_753 (O_753,N_29913,N_29769);
nand UO_754 (O_754,N_29602,N_29830);
and UO_755 (O_755,N_29860,N_29747);
nand UO_756 (O_756,N_29975,N_29543);
nor UO_757 (O_757,N_29612,N_29763);
or UO_758 (O_758,N_29757,N_29872);
xor UO_759 (O_759,N_29618,N_29972);
or UO_760 (O_760,N_29773,N_29537);
nor UO_761 (O_761,N_29812,N_29922);
and UO_762 (O_762,N_29682,N_29847);
or UO_763 (O_763,N_29553,N_29677);
or UO_764 (O_764,N_29950,N_29612);
and UO_765 (O_765,N_29838,N_29784);
nand UO_766 (O_766,N_29728,N_29571);
or UO_767 (O_767,N_29670,N_29593);
or UO_768 (O_768,N_29950,N_29779);
xor UO_769 (O_769,N_29537,N_29863);
nand UO_770 (O_770,N_29516,N_29830);
nand UO_771 (O_771,N_29974,N_29888);
xnor UO_772 (O_772,N_29508,N_29541);
xnor UO_773 (O_773,N_29582,N_29857);
or UO_774 (O_774,N_29819,N_29948);
xnor UO_775 (O_775,N_29663,N_29623);
or UO_776 (O_776,N_29732,N_29726);
xnor UO_777 (O_777,N_29513,N_29986);
and UO_778 (O_778,N_29560,N_29965);
nor UO_779 (O_779,N_29946,N_29574);
nor UO_780 (O_780,N_29992,N_29938);
and UO_781 (O_781,N_29886,N_29762);
nor UO_782 (O_782,N_29731,N_29914);
xor UO_783 (O_783,N_29940,N_29831);
and UO_784 (O_784,N_29644,N_29997);
nand UO_785 (O_785,N_29587,N_29713);
nand UO_786 (O_786,N_29775,N_29991);
or UO_787 (O_787,N_29920,N_29766);
xnor UO_788 (O_788,N_29638,N_29850);
or UO_789 (O_789,N_29986,N_29959);
or UO_790 (O_790,N_29509,N_29648);
or UO_791 (O_791,N_29777,N_29583);
xnor UO_792 (O_792,N_29923,N_29789);
nand UO_793 (O_793,N_29928,N_29593);
and UO_794 (O_794,N_29827,N_29744);
nand UO_795 (O_795,N_29634,N_29873);
and UO_796 (O_796,N_29754,N_29632);
nand UO_797 (O_797,N_29652,N_29719);
and UO_798 (O_798,N_29670,N_29854);
or UO_799 (O_799,N_29534,N_29638);
nand UO_800 (O_800,N_29964,N_29519);
or UO_801 (O_801,N_29565,N_29749);
nor UO_802 (O_802,N_29840,N_29709);
xnor UO_803 (O_803,N_29657,N_29605);
xor UO_804 (O_804,N_29699,N_29785);
xor UO_805 (O_805,N_29940,N_29781);
or UO_806 (O_806,N_29575,N_29557);
or UO_807 (O_807,N_29704,N_29994);
and UO_808 (O_808,N_29632,N_29625);
nand UO_809 (O_809,N_29620,N_29915);
nand UO_810 (O_810,N_29683,N_29747);
or UO_811 (O_811,N_29706,N_29641);
nor UO_812 (O_812,N_29626,N_29849);
nand UO_813 (O_813,N_29805,N_29882);
xnor UO_814 (O_814,N_29552,N_29881);
nor UO_815 (O_815,N_29833,N_29764);
and UO_816 (O_816,N_29614,N_29727);
nor UO_817 (O_817,N_29941,N_29771);
or UO_818 (O_818,N_29859,N_29738);
nand UO_819 (O_819,N_29559,N_29840);
nor UO_820 (O_820,N_29671,N_29764);
and UO_821 (O_821,N_29874,N_29565);
nand UO_822 (O_822,N_29847,N_29502);
nand UO_823 (O_823,N_29728,N_29791);
nor UO_824 (O_824,N_29823,N_29589);
and UO_825 (O_825,N_29971,N_29786);
xor UO_826 (O_826,N_29839,N_29570);
nand UO_827 (O_827,N_29852,N_29853);
and UO_828 (O_828,N_29583,N_29545);
xnor UO_829 (O_829,N_29845,N_29571);
nor UO_830 (O_830,N_29983,N_29798);
nor UO_831 (O_831,N_29769,N_29560);
nor UO_832 (O_832,N_29854,N_29919);
and UO_833 (O_833,N_29912,N_29553);
or UO_834 (O_834,N_29678,N_29501);
and UO_835 (O_835,N_29516,N_29832);
nor UO_836 (O_836,N_29746,N_29573);
nor UO_837 (O_837,N_29801,N_29637);
nand UO_838 (O_838,N_29678,N_29905);
nand UO_839 (O_839,N_29833,N_29796);
nor UO_840 (O_840,N_29873,N_29537);
and UO_841 (O_841,N_29746,N_29871);
and UO_842 (O_842,N_29820,N_29964);
or UO_843 (O_843,N_29618,N_29931);
nor UO_844 (O_844,N_29550,N_29691);
xor UO_845 (O_845,N_29968,N_29957);
nand UO_846 (O_846,N_29807,N_29629);
or UO_847 (O_847,N_29881,N_29703);
nand UO_848 (O_848,N_29915,N_29619);
and UO_849 (O_849,N_29522,N_29747);
nor UO_850 (O_850,N_29706,N_29630);
nor UO_851 (O_851,N_29554,N_29689);
or UO_852 (O_852,N_29588,N_29845);
nand UO_853 (O_853,N_29807,N_29650);
and UO_854 (O_854,N_29559,N_29904);
xnor UO_855 (O_855,N_29597,N_29749);
nor UO_856 (O_856,N_29785,N_29965);
nand UO_857 (O_857,N_29806,N_29786);
and UO_858 (O_858,N_29672,N_29923);
nor UO_859 (O_859,N_29560,N_29661);
xnor UO_860 (O_860,N_29924,N_29505);
nand UO_861 (O_861,N_29736,N_29979);
nor UO_862 (O_862,N_29945,N_29789);
and UO_863 (O_863,N_29790,N_29575);
or UO_864 (O_864,N_29617,N_29882);
or UO_865 (O_865,N_29718,N_29876);
nand UO_866 (O_866,N_29720,N_29571);
and UO_867 (O_867,N_29584,N_29768);
or UO_868 (O_868,N_29661,N_29645);
xor UO_869 (O_869,N_29972,N_29925);
and UO_870 (O_870,N_29975,N_29756);
or UO_871 (O_871,N_29570,N_29558);
and UO_872 (O_872,N_29688,N_29935);
nor UO_873 (O_873,N_29915,N_29790);
or UO_874 (O_874,N_29727,N_29630);
xor UO_875 (O_875,N_29880,N_29717);
xnor UO_876 (O_876,N_29950,N_29976);
nor UO_877 (O_877,N_29874,N_29991);
and UO_878 (O_878,N_29858,N_29629);
and UO_879 (O_879,N_29934,N_29609);
nor UO_880 (O_880,N_29529,N_29760);
nor UO_881 (O_881,N_29840,N_29831);
nor UO_882 (O_882,N_29997,N_29625);
nor UO_883 (O_883,N_29883,N_29770);
or UO_884 (O_884,N_29995,N_29517);
and UO_885 (O_885,N_29949,N_29738);
nor UO_886 (O_886,N_29851,N_29537);
nor UO_887 (O_887,N_29783,N_29966);
or UO_888 (O_888,N_29846,N_29567);
and UO_889 (O_889,N_29505,N_29953);
nand UO_890 (O_890,N_29710,N_29555);
and UO_891 (O_891,N_29595,N_29778);
nor UO_892 (O_892,N_29943,N_29754);
xnor UO_893 (O_893,N_29731,N_29880);
xor UO_894 (O_894,N_29730,N_29990);
or UO_895 (O_895,N_29866,N_29719);
nand UO_896 (O_896,N_29931,N_29531);
xor UO_897 (O_897,N_29765,N_29947);
xor UO_898 (O_898,N_29877,N_29788);
nor UO_899 (O_899,N_29935,N_29741);
nand UO_900 (O_900,N_29621,N_29971);
nor UO_901 (O_901,N_29875,N_29656);
and UO_902 (O_902,N_29552,N_29636);
or UO_903 (O_903,N_29582,N_29925);
and UO_904 (O_904,N_29719,N_29568);
xnor UO_905 (O_905,N_29954,N_29739);
xnor UO_906 (O_906,N_29796,N_29968);
xor UO_907 (O_907,N_29634,N_29881);
nand UO_908 (O_908,N_29812,N_29575);
and UO_909 (O_909,N_29864,N_29870);
nand UO_910 (O_910,N_29938,N_29659);
nand UO_911 (O_911,N_29704,N_29581);
or UO_912 (O_912,N_29940,N_29634);
and UO_913 (O_913,N_29678,N_29508);
xnor UO_914 (O_914,N_29881,N_29893);
nand UO_915 (O_915,N_29523,N_29565);
nand UO_916 (O_916,N_29604,N_29787);
nor UO_917 (O_917,N_29873,N_29679);
nand UO_918 (O_918,N_29595,N_29834);
nor UO_919 (O_919,N_29968,N_29568);
xor UO_920 (O_920,N_29879,N_29501);
xnor UO_921 (O_921,N_29803,N_29767);
nand UO_922 (O_922,N_29737,N_29514);
xor UO_923 (O_923,N_29968,N_29512);
and UO_924 (O_924,N_29505,N_29605);
and UO_925 (O_925,N_29946,N_29992);
and UO_926 (O_926,N_29583,N_29904);
and UO_927 (O_927,N_29956,N_29580);
or UO_928 (O_928,N_29540,N_29594);
xor UO_929 (O_929,N_29864,N_29862);
nor UO_930 (O_930,N_29760,N_29640);
or UO_931 (O_931,N_29568,N_29592);
xnor UO_932 (O_932,N_29718,N_29724);
or UO_933 (O_933,N_29865,N_29552);
nor UO_934 (O_934,N_29923,N_29942);
and UO_935 (O_935,N_29989,N_29675);
or UO_936 (O_936,N_29678,N_29648);
nand UO_937 (O_937,N_29936,N_29979);
and UO_938 (O_938,N_29560,N_29871);
and UO_939 (O_939,N_29653,N_29901);
and UO_940 (O_940,N_29809,N_29503);
xor UO_941 (O_941,N_29800,N_29978);
nor UO_942 (O_942,N_29850,N_29776);
and UO_943 (O_943,N_29794,N_29683);
nand UO_944 (O_944,N_29561,N_29646);
nand UO_945 (O_945,N_29921,N_29948);
nor UO_946 (O_946,N_29649,N_29525);
and UO_947 (O_947,N_29691,N_29666);
nor UO_948 (O_948,N_29656,N_29760);
nor UO_949 (O_949,N_29632,N_29782);
or UO_950 (O_950,N_29726,N_29650);
and UO_951 (O_951,N_29822,N_29929);
and UO_952 (O_952,N_29572,N_29681);
or UO_953 (O_953,N_29963,N_29686);
or UO_954 (O_954,N_29939,N_29775);
xnor UO_955 (O_955,N_29635,N_29719);
xnor UO_956 (O_956,N_29631,N_29776);
xor UO_957 (O_957,N_29762,N_29843);
and UO_958 (O_958,N_29922,N_29967);
nor UO_959 (O_959,N_29905,N_29818);
nor UO_960 (O_960,N_29569,N_29909);
xnor UO_961 (O_961,N_29513,N_29859);
xor UO_962 (O_962,N_29765,N_29764);
or UO_963 (O_963,N_29920,N_29595);
xnor UO_964 (O_964,N_29720,N_29914);
or UO_965 (O_965,N_29958,N_29840);
or UO_966 (O_966,N_29548,N_29716);
xnor UO_967 (O_967,N_29866,N_29787);
nand UO_968 (O_968,N_29692,N_29988);
or UO_969 (O_969,N_29815,N_29903);
nor UO_970 (O_970,N_29626,N_29649);
and UO_971 (O_971,N_29769,N_29503);
nor UO_972 (O_972,N_29981,N_29536);
xor UO_973 (O_973,N_29617,N_29691);
and UO_974 (O_974,N_29954,N_29883);
xnor UO_975 (O_975,N_29953,N_29840);
nor UO_976 (O_976,N_29847,N_29995);
nor UO_977 (O_977,N_29693,N_29674);
xnor UO_978 (O_978,N_29947,N_29925);
nor UO_979 (O_979,N_29622,N_29947);
or UO_980 (O_980,N_29737,N_29950);
xor UO_981 (O_981,N_29688,N_29879);
nor UO_982 (O_982,N_29795,N_29934);
or UO_983 (O_983,N_29687,N_29753);
or UO_984 (O_984,N_29797,N_29809);
nand UO_985 (O_985,N_29735,N_29527);
nor UO_986 (O_986,N_29942,N_29515);
xor UO_987 (O_987,N_29573,N_29828);
and UO_988 (O_988,N_29839,N_29971);
nor UO_989 (O_989,N_29699,N_29523);
nand UO_990 (O_990,N_29623,N_29573);
nand UO_991 (O_991,N_29794,N_29895);
xor UO_992 (O_992,N_29687,N_29910);
or UO_993 (O_993,N_29924,N_29767);
nand UO_994 (O_994,N_29994,N_29905);
nand UO_995 (O_995,N_29600,N_29520);
or UO_996 (O_996,N_29882,N_29592);
or UO_997 (O_997,N_29564,N_29684);
nor UO_998 (O_998,N_29974,N_29523);
nor UO_999 (O_999,N_29727,N_29649);
xnor UO_1000 (O_1000,N_29706,N_29734);
or UO_1001 (O_1001,N_29908,N_29568);
nand UO_1002 (O_1002,N_29761,N_29699);
or UO_1003 (O_1003,N_29939,N_29996);
and UO_1004 (O_1004,N_29521,N_29865);
nor UO_1005 (O_1005,N_29616,N_29981);
nand UO_1006 (O_1006,N_29970,N_29847);
and UO_1007 (O_1007,N_29974,N_29636);
or UO_1008 (O_1008,N_29645,N_29540);
or UO_1009 (O_1009,N_29519,N_29528);
and UO_1010 (O_1010,N_29690,N_29746);
or UO_1011 (O_1011,N_29646,N_29773);
or UO_1012 (O_1012,N_29732,N_29569);
nand UO_1013 (O_1013,N_29836,N_29613);
or UO_1014 (O_1014,N_29636,N_29706);
xor UO_1015 (O_1015,N_29993,N_29694);
xor UO_1016 (O_1016,N_29825,N_29973);
nor UO_1017 (O_1017,N_29686,N_29610);
nand UO_1018 (O_1018,N_29965,N_29706);
nor UO_1019 (O_1019,N_29910,N_29515);
xnor UO_1020 (O_1020,N_29798,N_29991);
xor UO_1021 (O_1021,N_29713,N_29683);
or UO_1022 (O_1022,N_29741,N_29688);
nand UO_1023 (O_1023,N_29900,N_29632);
nand UO_1024 (O_1024,N_29786,N_29841);
nor UO_1025 (O_1025,N_29662,N_29717);
xnor UO_1026 (O_1026,N_29841,N_29988);
nand UO_1027 (O_1027,N_29552,N_29916);
xnor UO_1028 (O_1028,N_29643,N_29976);
and UO_1029 (O_1029,N_29919,N_29860);
xor UO_1030 (O_1030,N_29660,N_29966);
nand UO_1031 (O_1031,N_29659,N_29588);
nand UO_1032 (O_1032,N_29791,N_29617);
nor UO_1033 (O_1033,N_29614,N_29580);
xor UO_1034 (O_1034,N_29940,N_29678);
and UO_1035 (O_1035,N_29718,N_29752);
or UO_1036 (O_1036,N_29792,N_29597);
xor UO_1037 (O_1037,N_29840,N_29783);
and UO_1038 (O_1038,N_29833,N_29609);
and UO_1039 (O_1039,N_29528,N_29993);
xor UO_1040 (O_1040,N_29700,N_29865);
and UO_1041 (O_1041,N_29940,N_29943);
nand UO_1042 (O_1042,N_29751,N_29863);
xor UO_1043 (O_1043,N_29760,N_29624);
and UO_1044 (O_1044,N_29897,N_29723);
and UO_1045 (O_1045,N_29988,N_29837);
xnor UO_1046 (O_1046,N_29612,N_29678);
or UO_1047 (O_1047,N_29989,N_29985);
and UO_1048 (O_1048,N_29706,N_29999);
nor UO_1049 (O_1049,N_29500,N_29679);
nor UO_1050 (O_1050,N_29702,N_29781);
and UO_1051 (O_1051,N_29977,N_29565);
or UO_1052 (O_1052,N_29883,N_29554);
and UO_1053 (O_1053,N_29736,N_29983);
nor UO_1054 (O_1054,N_29821,N_29687);
nand UO_1055 (O_1055,N_29915,N_29685);
xnor UO_1056 (O_1056,N_29652,N_29594);
nand UO_1057 (O_1057,N_29690,N_29546);
or UO_1058 (O_1058,N_29772,N_29908);
and UO_1059 (O_1059,N_29837,N_29875);
xnor UO_1060 (O_1060,N_29532,N_29774);
and UO_1061 (O_1061,N_29888,N_29771);
nand UO_1062 (O_1062,N_29715,N_29979);
or UO_1063 (O_1063,N_29526,N_29896);
and UO_1064 (O_1064,N_29753,N_29992);
xor UO_1065 (O_1065,N_29541,N_29796);
xor UO_1066 (O_1066,N_29662,N_29673);
xor UO_1067 (O_1067,N_29863,N_29950);
nand UO_1068 (O_1068,N_29763,N_29993);
nor UO_1069 (O_1069,N_29937,N_29515);
xnor UO_1070 (O_1070,N_29732,N_29584);
or UO_1071 (O_1071,N_29913,N_29619);
xor UO_1072 (O_1072,N_29595,N_29500);
nand UO_1073 (O_1073,N_29729,N_29777);
or UO_1074 (O_1074,N_29669,N_29636);
or UO_1075 (O_1075,N_29580,N_29511);
nand UO_1076 (O_1076,N_29929,N_29850);
nor UO_1077 (O_1077,N_29559,N_29683);
xor UO_1078 (O_1078,N_29679,N_29604);
nor UO_1079 (O_1079,N_29500,N_29934);
nor UO_1080 (O_1080,N_29921,N_29641);
xnor UO_1081 (O_1081,N_29958,N_29981);
and UO_1082 (O_1082,N_29833,N_29819);
nor UO_1083 (O_1083,N_29807,N_29924);
nand UO_1084 (O_1084,N_29685,N_29770);
nor UO_1085 (O_1085,N_29742,N_29853);
and UO_1086 (O_1086,N_29588,N_29746);
and UO_1087 (O_1087,N_29524,N_29867);
xnor UO_1088 (O_1088,N_29719,N_29521);
or UO_1089 (O_1089,N_29826,N_29885);
and UO_1090 (O_1090,N_29789,N_29744);
and UO_1091 (O_1091,N_29589,N_29601);
and UO_1092 (O_1092,N_29821,N_29759);
and UO_1093 (O_1093,N_29583,N_29616);
nor UO_1094 (O_1094,N_29863,N_29571);
xnor UO_1095 (O_1095,N_29588,N_29830);
and UO_1096 (O_1096,N_29852,N_29835);
nand UO_1097 (O_1097,N_29719,N_29994);
or UO_1098 (O_1098,N_29849,N_29708);
xor UO_1099 (O_1099,N_29840,N_29632);
nor UO_1100 (O_1100,N_29842,N_29949);
or UO_1101 (O_1101,N_29708,N_29636);
nand UO_1102 (O_1102,N_29659,N_29988);
xor UO_1103 (O_1103,N_29920,N_29761);
nand UO_1104 (O_1104,N_29822,N_29880);
xor UO_1105 (O_1105,N_29766,N_29883);
and UO_1106 (O_1106,N_29892,N_29887);
or UO_1107 (O_1107,N_29871,N_29824);
and UO_1108 (O_1108,N_29785,N_29781);
nor UO_1109 (O_1109,N_29995,N_29677);
and UO_1110 (O_1110,N_29693,N_29542);
or UO_1111 (O_1111,N_29770,N_29540);
and UO_1112 (O_1112,N_29513,N_29522);
or UO_1113 (O_1113,N_29546,N_29911);
nand UO_1114 (O_1114,N_29994,N_29695);
xnor UO_1115 (O_1115,N_29865,N_29977);
or UO_1116 (O_1116,N_29950,N_29722);
nand UO_1117 (O_1117,N_29824,N_29606);
or UO_1118 (O_1118,N_29704,N_29946);
nor UO_1119 (O_1119,N_29965,N_29526);
and UO_1120 (O_1120,N_29989,N_29910);
nor UO_1121 (O_1121,N_29880,N_29810);
and UO_1122 (O_1122,N_29620,N_29818);
nand UO_1123 (O_1123,N_29503,N_29639);
nand UO_1124 (O_1124,N_29617,N_29863);
or UO_1125 (O_1125,N_29641,N_29683);
nor UO_1126 (O_1126,N_29849,N_29667);
and UO_1127 (O_1127,N_29551,N_29757);
and UO_1128 (O_1128,N_29917,N_29886);
xor UO_1129 (O_1129,N_29671,N_29658);
nand UO_1130 (O_1130,N_29829,N_29534);
or UO_1131 (O_1131,N_29911,N_29992);
nor UO_1132 (O_1132,N_29523,N_29559);
xor UO_1133 (O_1133,N_29952,N_29731);
nand UO_1134 (O_1134,N_29892,N_29857);
xor UO_1135 (O_1135,N_29716,N_29755);
and UO_1136 (O_1136,N_29672,N_29946);
xor UO_1137 (O_1137,N_29875,N_29659);
nor UO_1138 (O_1138,N_29554,N_29835);
nor UO_1139 (O_1139,N_29676,N_29600);
nand UO_1140 (O_1140,N_29912,N_29877);
nand UO_1141 (O_1141,N_29683,N_29846);
or UO_1142 (O_1142,N_29509,N_29767);
nor UO_1143 (O_1143,N_29852,N_29997);
xor UO_1144 (O_1144,N_29585,N_29678);
or UO_1145 (O_1145,N_29876,N_29747);
and UO_1146 (O_1146,N_29900,N_29558);
nor UO_1147 (O_1147,N_29593,N_29739);
xnor UO_1148 (O_1148,N_29862,N_29707);
or UO_1149 (O_1149,N_29637,N_29761);
xor UO_1150 (O_1150,N_29786,N_29763);
xnor UO_1151 (O_1151,N_29900,N_29582);
or UO_1152 (O_1152,N_29669,N_29680);
or UO_1153 (O_1153,N_29608,N_29954);
nand UO_1154 (O_1154,N_29694,N_29592);
xor UO_1155 (O_1155,N_29717,N_29982);
or UO_1156 (O_1156,N_29847,N_29554);
or UO_1157 (O_1157,N_29813,N_29984);
and UO_1158 (O_1158,N_29752,N_29641);
and UO_1159 (O_1159,N_29517,N_29894);
xnor UO_1160 (O_1160,N_29721,N_29833);
nor UO_1161 (O_1161,N_29972,N_29849);
or UO_1162 (O_1162,N_29591,N_29814);
xor UO_1163 (O_1163,N_29602,N_29993);
or UO_1164 (O_1164,N_29703,N_29516);
nand UO_1165 (O_1165,N_29921,N_29587);
nor UO_1166 (O_1166,N_29539,N_29938);
and UO_1167 (O_1167,N_29658,N_29957);
or UO_1168 (O_1168,N_29610,N_29917);
nor UO_1169 (O_1169,N_29963,N_29619);
xor UO_1170 (O_1170,N_29540,N_29546);
or UO_1171 (O_1171,N_29849,N_29895);
nand UO_1172 (O_1172,N_29757,N_29858);
and UO_1173 (O_1173,N_29763,N_29832);
or UO_1174 (O_1174,N_29500,N_29893);
nor UO_1175 (O_1175,N_29939,N_29579);
or UO_1176 (O_1176,N_29924,N_29700);
nand UO_1177 (O_1177,N_29787,N_29846);
nor UO_1178 (O_1178,N_29659,N_29572);
nand UO_1179 (O_1179,N_29875,N_29529);
nor UO_1180 (O_1180,N_29998,N_29687);
xor UO_1181 (O_1181,N_29906,N_29878);
and UO_1182 (O_1182,N_29881,N_29722);
nor UO_1183 (O_1183,N_29704,N_29552);
and UO_1184 (O_1184,N_29828,N_29513);
xor UO_1185 (O_1185,N_29646,N_29707);
nand UO_1186 (O_1186,N_29732,N_29663);
and UO_1187 (O_1187,N_29988,N_29915);
nand UO_1188 (O_1188,N_29704,N_29796);
or UO_1189 (O_1189,N_29879,N_29525);
nor UO_1190 (O_1190,N_29983,N_29580);
and UO_1191 (O_1191,N_29881,N_29992);
or UO_1192 (O_1192,N_29631,N_29563);
xor UO_1193 (O_1193,N_29728,N_29784);
nor UO_1194 (O_1194,N_29999,N_29693);
nand UO_1195 (O_1195,N_29697,N_29628);
and UO_1196 (O_1196,N_29788,N_29531);
nor UO_1197 (O_1197,N_29900,N_29739);
or UO_1198 (O_1198,N_29533,N_29625);
or UO_1199 (O_1199,N_29866,N_29992);
or UO_1200 (O_1200,N_29615,N_29716);
nand UO_1201 (O_1201,N_29956,N_29514);
or UO_1202 (O_1202,N_29862,N_29797);
xnor UO_1203 (O_1203,N_29743,N_29790);
nand UO_1204 (O_1204,N_29717,N_29567);
xnor UO_1205 (O_1205,N_29856,N_29779);
or UO_1206 (O_1206,N_29923,N_29812);
and UO_1207 (O_1207,N_29726,N_29828);
xor UO_1208 (O_1208,N_29514,N_29619);
or UO_1209 (O_1209,N_29774,N_29935);
nand UO_1210 (O_1210,N_29833,N_29718);
or UO_1211 (O_1211,N_29539,N_29756);
and UO_1212 (O_1212,N_29539,N_29514);
nand UO_1213 (O_1213,N_29813,N_29735);
or UO_1214 (O_1214,N_29814,N_29804);
nand UO_1215 (O_1215,N_29963,N_29585);
xnor UO_1216 (O_1216,N_29672,N_29560);
or UO_1217 (O_1217,N_29820,N_29985);
nand UO_1218 (O_1218,N_29849,N_29510);
nor UO_1219 (O_1219,N_29802,N_29919);
nand UO_1220 (O_1220,N_29573,N_29578);
xor UO_1221 (O_1221,N_29935,N_29760);
nor UO_1222 (O_1222,N_29572,N_29940);
nor UO_1223 (O_1223,N_29694,N_29753);
or UO_1224 (O_1224,N_29616,N_29911);
xnor UO_1225 (O_1225,N_29534,N_29875);
and UO_1226 (O_1226,N_29738,N_29914);
xnor UO_1227 (O_1227,N_29927,N_29984);
or UO_1228 (O_1228,N_29556,N_29555);
nor UO_1229 (O_1229,N_29591,N_29910);
xnor UO_1230 (O_1230,N_29876,N_29792);
nor UO_1231 (O_1231,N_29969,N_29671);
nor UO_1232 (O_1232,N_29938,N_29838);
or UO_1233 (O_1233,N_29685,N_29727);
and UO_1234 (O_1234,N_29777,N_29810);
xnor UO_1235 (O_1235,N_29710,N_29914);
nor UO_1236 (O_1236,N_29704,N_29998);
or UO_1237 (O_1237,N_29693,N_29607);
nand UO_1238 (O_1238,N_29720,N_29875);
xnor UO_1239 (O_1239,N_29778,N_29981);
nand UO_1240 (O_1240,N_29777,N_29727);
or UO_1241 (O_1241,N_29560,N_29716);
and UO_1242 (O_1242,N_29523,N_29906);
nor UO_1243 (O_1243,N_29624,N_29582);
and UO_1244 (O_1244,N_29949,N_29760);
nor UO_1245 (O_1245,N_29979,N_29600);
nor UO_1246 (O_1246,N_29692,N_29570);
nand UO_1247 (O_1247,N_29730,N_29845);
nand UO_1248 (O_1248,N_29906,N_29845);
or UO_1249 (O_1249,N_29899,N_29804);
nor UO_1250 (O_1250,N_29650,N_29719);
nor UO_1251 (O_1251,N_29725,N_29799);
xnor UO_1252 (O_1252,N_29861,N_29801);
or UO_1253 (O_1253,N_29838,N_29716);
and UO_1254 (O_1254,N_29966,N_29618);
and UO_1255 (O_1255,N_29521,N_29888);
nor UO_1256 (O_1256,N_29856,N_29796);
or UO_1257 (O_1257,N_29757,N_29950);
nor UO_1258 (O_1258,N_29558,N_29678);
xor UO_1259 (O_1259,N_29720,N_29781);
and UO_1260 (O_1260,N_29756,N_29582);
nor UO_1261 (O_1261,N_29760,N_29510);
nand UO_1262 (O_1262,N_29785,N_29904);
or UO_1263 (O_1263,N_29728,N_29971);
and UO_1264 (O_1264,N_29598,N_29916);
or UO_1265 (O_1265,N_29991,N_29882);
or UO_1266 (O_1266,N_29972,N_29724);
xor UO_1267 (O_1267,N_29834,N_29663);
or UO_1268 (O_1268,N_29500,N_29604);
or UO_1269 (O_1269,N_29829,N_29728);
xor UO_1270 (O_1270,N_29963,N_29904);
xor UO_1271 (O_1271,N_29807,N_29680);
nor UO_1272 (O_1272,N_29635,N_29852);
nand UO_1273 (O_1273,N_29696,N_29704);
xnor UO_1274 (O_1274,N_29663,N_29800);
xor UO_1275 (O_1275,N_29836,N_29558);
xor UO_1276 (O_1276,N_29914,N_29612);
xor UO_1277 (O_1277,N_29618,N_29836);
nor UO_1278 (O_1278,N_29880,N_29910);
nor UO_1279 (O_1279,N_29871,N_29960);
and UO_1280 (O_1280,N_29712,N_29814);
nor UO_1281 (O_1281,N_29632,N_29811);
nor UO_1282 (O_1282,N_29989,N_29549);
xor UO_1283 (O_1283,N_29758,N_29873);
nor UO_1284 (O_1284,N_29792,N_29698);
xnor UO_1285 (O_1285,N_29501,N_29536);
and UO_1286 (O_1286,N_29897,N_29823);
and UO_1287 (O_1287,N_29604,N_29796);
xor UO_1288 (O_1288,N_29688,N_29832);
or UO_1289 (O_1289,N_29618,N_29500);
xnor UO_1290 (O_1290,N_29913,N_29783);
nand UO_1291 (O_1291,N_29569,N_29749);
or UO_1292 (O_1292,N_29898,N_29901);
xnor UO_1293 (O_1293,N_29911,N_29805);
or UO_1294 (O_1294,N_29591,N_29998);
nor UO_1295 (O_1295,N_29541,N_29634);
nand UO_1296 (O_1296,N_29657,N_29932);
xor UO_1297 (O_1297,N_29563,N_29688);
and UO_1298 (O_1298,N_29899,N_29725);
nand UO_1299 (O_1299,N_29923,N_29765);
xnor UO_1300 (O_1300,N_29538,N_29610);
or UO_1301 (O_1301,N_29858,N_29875);
nor UO_1302 (O_1302,N_29560,N_29774);
xnor UO_1303 (O_1303,N_29864,N_29701);
nand UO_1304 (O_1304,N_29669,N_29997);
nor UO_1305 (O_1305,N_29568,N_29883);
nor UO_1306 (O_1306,N_29713,N_29541);
or UO_1307 (O_1307,N_29655,N_29677);
xor UO_1308 (O_1308,N_29899,N_29760);
and UO_1309 (O_1309,N_29943,N_29657);
or UO_1310 (O_1310,N_29501,N_29975);
or UO_1311 (O_1311,N_29612,N_29587);
nand UO_1312 (O_1312,N_29797,N_29662);
xor UO_1313 (O_1313,N_29813,N_29720);
nand UO_1314 (O_1314,N_29940,N_29899);
nand UO_1315 (O_1315,N_29757,N_29556);
nor UO_1316 (O_1316,N_29543,N_29813);
or UO_1317 (O_1317,N_29936,N_29916);
xnor UO_1318 (O_1318,N_29982,N_29853);
xor UO_1319 (O_1319,N_29773,N_29745);
or UO_1320 (O_1320,N_29543,N_29598);
nor UO_1321 (O_1321,N_29853,N_29757);
nor UO_1322 (O_1322,N_29570,N_29773);
nor UO_1323 (O_1323,N_29652,N_29925);
or UO_1324 (O_1324,N_29904,N_29948);
nor UO_1325 (O_1325,N_29753,N_29787);
or UO_1326 (O_1326,N_29614,N_29891);
xnor UO_1327 (O_1327,N_29888,N_29979);
or UO_1328 (O_1328,N_29896,N_29984);
and UO_1329 (O_1329,N_29920,N_29668);
nor UO_1330 (O_1330,N_29511,N_29937);
nor UO_1331 (O_1331,N_29546,N_29952);
nand UO_1332 (O_1332,N_29556,N_29889);
or UO_1333 (O_1333,N_29794,N_29786);
nand UO_1334 (O_1334,N_29851,N_29967);
nor UO_1335 (O_1335,N_29608,N_29856);
nand UO_1336 (O_1336,N_29894,N_29516);
nand UO_1337 (O_1337,N_29913,N_29520);
nand UO_1338 (O_1338,N_29678,N_29830);
or UO_1339 (O_1339,N_29805,N_29898);
and UO_1340 (O_1340,N_29820,N_29557);
or UO_1341 (O_1341,N_29645,N_29647);
nand UO_1342 (O_1342,N_29506,N_29578);
nor UO_1343 (O_1343,N_29693,N_29893);
and UO_1344 (O_1344,N_29792,N_29731);
or UO_1345 (O_1345,N_29502,N_29830);
xnor UO_1346 (O_1346,N_29701,N_29832);
or UO_1347 (O_1347,N_29612,N_29734);
or UO_1348 (O_1348,N_29580,N_29931);
xnor UO_1349 (O_1349,N_29981,N_29866);
nand UO_1350 (O_1350,N_29667,N_29612);
or UO_1351 (O_1351,N_29605,N_29753);
nor UO_1352 (O_1352,N_29635,N_29561);
or UO_1353 (O_1353,N_29721,N_29609);
xnor UO_1354 (O_1354,N_29751,N_29664);
or UO_1355 (O_1355,N_29691,N_29894);
nand UO_1356 (O_1356,N_29710,N_29859);
nor UO_1357 (O_1357,N_29770,N_29576);
nor UO_1358 (O_1358,N_29974,N_29579);
xnor UO_1359 (O_1359,N_29759,N_29656);
and UO_1360 (O_1360,N_29697,N_29932);
nor UO_1361 (O_1361,N_29610,N_29580);
or UO_1362 (O_1362,N_29901,N_29508);
or UO_1363 (O_1363,N_29989,N_29775);
and UO_1364 (O_1364,N_29521,N_29936);
nor UO_1365 (O_1365,N_29729,N_29695);
nand UO_1366 (O_1366,N_29809,N_29720);
nor UO_1367 (O_1367,N_29614,N_29521);
nor UO_1368 (O_1368,N_29651,N_29742);
and UO_1369 (O_1369,N_29778,N_29532);
nand UO_1370 (O_1370,N_29856,N_29613);
nand UO_1371 (O_1371,N_29956,N_29613);
or UO_1372 (O_1372,N_29878,N_29804);
or UO_1373 (O_1373,N_29920,N_29916);
nor UO_1374 (O_1374,N_29657,N_29549);
nand UO_1375 (O_1375,N_29642,N_29850);
xnor UO_1376 (O_1376,N_29628,N_29510);
xor UO_1377 (O_1377,N_29553,N_29559);
nand UO_1378 (O_1378,N_29974,N_29918);
nor UO_1379 (O_1379,N_29823,N_29639);
nand UO_1380 (O_1380,N_29931,N_29664);
nand UO_1381 (O_1381,N_29554,N_29950);
xnor UO_1382 (O_1382,N_29603,N_29718);
nor UO_1383 (O_1383,N_29980,N_29593);
and UO_1384 (O_1384,N_29792,N_29996);
nand UO_1385 (O_1385,N_29571,N_29755);
nand UO_1386 (O_1386,N_29939,N_29937);
or UO_1387 (O_1387,N_29888,N_29528);
or UO_1388 (O_1388,N_29694,N_29556);
nor UO_1389 (O_1389,N_29951,N_29741);
xnor UO_1390 (O_1390,N_29584,N_29758);
or UO_1391 (O_1391,N_29906,N_29867);
or UO_1392 (O_1392,N_29866,N_29853);
and UO_1393 (O_1393,N_29998,N_29522);
nand UO_1394 (O_1394,N_29932,N_29871);
nor UO_1395 (O_1395,N_29743,N_29821);
and UO_1396 (O_1396,N_29693,N_29730);
and UO_1397 (O_1397,N_29898,N_29942);
or UO_1398 (O_1398,N_29653,N_29728);
nor UO_1399 (O_1399,N_29737,N_29604);
or UO_1400 (O_1400,N_29871,N_29849);
xor UO_1401 (O_1401,N_29938,N_29532);
and UO_1402 (O_1402,N_29601,N_29730);
xor UO_1403 (O_1403,N_29732,N_29554);
or UO_1404 (O_1404,N_29669,N_29648);
xnor UO_1405 (O_1405,N_29856,N_29931);
nand UO_1406 (O_1406,N_29615,N_29602);
or UO_1407 (O_1407,N_29804,N_29813);
and UO_1408 (O_1408,N_29533,N_29721);
or UO_1409 (O_1409,N_29665,N_29593);
or UO_1410 (O_1410,N_29895,N_29574);
and UO_1411 (O_1411,N_29663,N_29682);
nor UO_1412 (O_1412,N_29728,N_29544);
nor UO_1413 (O_1413,N_29714,N_29844);
or UO_1414 (O_1414,N_29732,N_29783);
nor UO_1415 (O_1415,N_29600,N_29700);
or UO_1416 (O_1416,N_29999,N_29936);
or UO_1417 (O_1417,N_29987,N_29525);
nand UO_1418 (O_1418,N_29957,N_29754);
nor UO_1419 (O_1419,N_29643,N_29724);
or UO_1420 (O_1420,N_29757,N_29502);
or UO_1421 (O_1421,N_29999,N_29807);
and UO_1422 (O_1422,N_29833,N_29704);
and UO_1423 (O_1423,N_29548,N_29559);
nand UO_1424 (O_1424,N_29985,N_29929);
nand UO_1425 (O_1425,N_29663,N_29863);
xnor UO_1426 (O_1426,N_29523,N_29606);
or UO_1427 (O_1427,N_29827,N_29576);
or UO_1428 (O_1428,N_29521,N_29862);
or UO_1429 (O_1429,N_29583,N_29849);
xor UO_1430 (O_1430,N_29722,N_29749);
nor UO_1431 (O_1431,N_29857,N_29695);
nand UO_1432 (O_1432,N_29922,N_29669);
nor UO_1433 (O_1433,N_29699,N_29922);
nor UO_1434 (O_1434,N_29630,N_29614);
nand UO_1435 (O_1435,N_29880,N_29696);
and UO_1436 (O_1436,N_29656,N_29986);
nand UO_1437 (O_1437,N_29687,N_29882);
nand UO_1438 (O_1438,N_29999,N_29888);
nor UO_1439 (O_1439,N_29863,N_29883);
nor UO_1440 (O_1440,N_29820,N_29552);
and UO_1441 (O_1441,N_29779,N_29519);
nand UO_1442 (O_1442,N_29529,N_29894);
or UO_1443 (O_1443,N_29774,N_29713);
or UO_1444 (O_1444,N_29910,N_29715);
or UO_1445 (O_1445,N_29587,N_29596);
xor UO_1446 (O_1446,N_29521,N_29513);
and UO_1447 (O_1447,N_29913,N_29938);
nor UO_1448 (O_1448,N_29774,N_29825);
nor UO_1449 (O_1449,N_29956,N_29511);
nand UO_1450 (O_1450,N_29744,N_29502);
xnor UO_1451 (O_1451,N_29613,N_29695);
nand UO_1452 (O_1452,N_29643,N_29801);
nand UO_1453 (O_1453,N_29780,N_29579);
nand UO_1454 (O_1454,N_29576,N_29550);
xnor UO_1455 (O_1455,N_29882,N_29585);
nor UO_1456 (O_1456,N_29981,N_29568);
xor UO_1457 (O_1457,N_29699,N_29694);
xnor UO_1458 (O_1458,N_29791,N_29565);
nor UO_1459 (O_1459,N_29761,N_29884);
nor UO_1460 (O_1460,N_29747,N_29506);
nand UO_1461 (O_1461,N_29522,N_29609);
and UO_1462 (O_1462,N_29546,N_29787);
nor UO_1463 (O_1463,N_29749,N_29635);
nand UO_1464 (O_1464,N_29500,N_29837);
xnor UO_1465 (O_1465,N_29891,N_29570);
and UO_1466 (O_1466,N_29574,N_29568);
nor UO_1467 (O_1467,N_29832,N_29938);
or UO_1468 (O_1468,N_29521,N_29525);
nand UO_1469 (O_1469,N_29930,N_29734);
nor UO_1470 (O_1470,N_29967,N_29763);
nor UO_1471 (O_1471,N_29592,N_29781);
xnor UO_1472 (O_1472,N_29568,N_29614);
nor UO_1473 (O_1473,N_29798,N_29618);
or UO_1474 (O_1474,N_29843,N_29581);
nor UO_1475 (O_1475,N_29965,N_29588);
or UO_1476 (O_1476,N_29689,N_29740);
xnor UO_1477 (O_1477,N_29753,N_29817);
or UO_1478 (O_1478,N_29879,N_29661);
or UO_1479 (O_1479,N_29793,N_29503);
or UO_1480 (O_1480,N_29906,N_29882);
or UO_1481 (O_1481,N_29648,N_29842);
nor UO_1482 (O_1482,N_29936,N_29805);
xor UO_1483 (O_1483,N_29682,N_29755);
and UO_1484 (O_1484,N_29788,N_29665);
nor UO_1485 (O_1485,N_29753,N_29941);
or UO_1486 (O_1486,N_29708,N_29665);
xor UO_1487 (O_1487,N_29969,N_29883);
xnor UO_1488 (O_1488,N_29848,N_29767);
nand UO_1489 (O_1489,N_29532,N_29678);
or UO_1490 (O_1490,N_29909,N_29972);
or UO_1491 (O_1491,N_29564,N_29862);
or UO_1492 (O_1492,N_29528,N_29940);
or UO_1493 (O_1493,N_29633,N_29761);
or UO_1494 (O_1494,N_29526,N_29999);
xnor UO_1495 (O_1495,N_29687,N_29562);
nor UO_1496 (O_1496,N_29872,N_29874);
nor UO_1497 (O_1497,N_29932,N_29746);
nand UO_1498 (O_1498,N_29822,N_29816);
nand UO_1499 (O_1499,N_29897,N_29756);
nand UO_1500 (O_1500,N_29908,N_29918);
and UO_1501 (O_1501,N_29627,N_29628);
or UO_1502 (O_1502,N_29960,N_29564);
or UO_1503 (O_1503,N_29683,N_29743);
and UO_1504 (O_1504,N_29682,N_29549);
or UO_1505 (O_1505,N_29887,N_29573);
or UO_1506 (O_1506,N_29765,N_29773);
and UO_1507 (O_1507,N_29551,N_29760);
nor UO_1508 (O_1508,N_29622,N_29765);
nand UO_1509 (O_1509,N_29696,N_29538);
and UO_1510 (O_1510,N_29535,N_29865);
and UO_1511 (O_1511,N_29638,N_29975);
nor UO_1512 (O_1512,N_29889,N_29662);
and UO_1513 (O_1513,N_29581,N_29958);
xor UO_1514 (O_1514,N_29822,N_29891);
nand UO_1515 (O_1515,N_29898,N_29864);
nor UO_1516 (O_1516,N_29619,N_29556);
and UO_1517 (O_1517,N_29640,N_29942);
nor UO_1518 (O_1518,N_29655,N_29537);
or UO_1519 (O_1519,N_29799,N_29671);
nand UO_1520 (O_1520,N_29805,N_29628);
or UO_1521 (O_1521,N_29988,N_29780);
or UO_1522 (O_1522,N_29773,N_29737);
nor UO_1523 (O_1523,N_29772,N_29781);
xnor UO_1524 (O_1524,N_29878,N_29759);
or UO_1525 (O_1525,N_29753,N_29662);
and UO_1526 (O_1526,N_29676,N_29584);
nor UO_1527 (O_1527,N_29656,N_29958);
xor UO_1528 (O_1528,N_29673,N_29962);
xor UO_1529 (O_1529,N_29831,N_29963);
nor UO_1530 (O_1530,N_29922,N_29679);
nand UO_1531 (O_1531,N_29688,N_29815);
nor UO_1532 (O_1532,N_29795,N_29792);
nand UO_1533 (O_1533,N_29942,N_29556);
and UO_1534 (O_1534,N_29869,N_29950);
nand UO_1535 (O_1535,N_29796,N_29689);
nor UO_1536 (O_1536,N_29897,N_29621);
xor UO_1537 (O_1537,N_29735,N_29502);
nand UO_1538 (O_1538,N_29651,N_29800);
and UO_1539 (O_1539,N_29539,N_29952);
or UO_1540 (O_1540,N_29755,N_29593);
nand UO_1541 (O_1541,N_29648,N_29639);
or UO_1542 (O_1542,N_29898,N_29884);
xnor UO_1543 (O_1543,N_29893,N_29825);
nand UO_1544 (O_1544,N_29895,N_29840);
xor UO_1545 (O_1545,N_29985,N_29560);
or UO_1546 (O_1546,N_29905,N_29972);
nor UO_1547 (O_1547,N_29521,N_29734);
nor UO_1548 (O_1548,N_29903,N_29654);
xor UO_1549 (O_1549,N_29618,N_29740);
nor UO_1550 (O_1550,N_29749,N_29958);
xor UO_1551 (O_1551,N_29695,N_29531);
or UO_1552 (O_1552,N_29896,N_29548);
and UO_1553 (O_1553,N_29893,N_29992);
xor UO_1554 (O_1554,N_29788,N_29688);
nor UO_1555 (O_1555,N_29724,N_29708);
or UO_1556 (O_1556,N_29945,N_29877);
or UO_1557 (O_1557,N_29535,N_29895);
nand UO_1558 (O_1558,N_29689,N_29916);
xor UO_1559 (O_1559,N_29836,N_29615);
nand UO_1560 (O_1560,N_29717,N_29645);
nor UO_1561 (O_1561,N_29816,N_29560);
nand UO_1562 (O_1562,N_29803,N_29939);
nor UO_1563 (O_1563,N_29885,N_29776);
or UO_1564 (O_1564,N_29556,N_29683);
xnor UO_1565 (O_1565,N_29653,N_29768);
nor UO_1566 (O_1566,N_29974,N_29557);
nand UO_1567 (O_1567,N_29811,N_29882);
or UO_1568 (O_1568,N_29823,N_29972);
xnor UO_1569 (O_1569,N_29713,N_29888);
or UO_1570 (O_1570,N_29820,N_29963);
nor UO_1571 (O_1571,N_29640,N_29837);
nand UO_1572 (O_1572,N_29696,N_29989);
nand UO_1573 (O_1573,N_29620,N_29860);
nor UO_1574 (O_1574,N_29815,N_29949);
xnor UO_1575 (O_1575,N_29543,N_29508);
nor UO_1576 (O_1576,N_29637,N_29632);
and UO_1577 (O_1577,N_29900,N_29716);
xnor UO_1578 (O_1578,N_29947,N_29702);
or UO_1579 (O_1579,N_29752,N_29703);
nand UO_1580 (O_1580,N_29588,N_29631);
xor UO_1581 (O_1581,N_29572,N_29989);
nor UO_1582 (O_1582,N_29512,N_29813);
nor UO_1583 (O_1583,N_29510,N_29852);
xor UO_1584 (O_1584,N_29875,N_29613);
or UO_1585 (O_1585,N_29676,N_29917);
and UO_1586 (O_1586,N_29917,N_29825);
nand UO_1587 (O_1587,N_29702,N_29751);
or UO_1588 (O_1588,N_29895,N_29999);
or UO_1589 (O_1589,N_29707,N_29666);
nand UO_1590 (O_1590,N_29614,N_29692);
nand UO_1591 (O_1591,N_29764,N_29926);
nor UO_1592 (O_1592,N_29664,N_29687);
nand UO_1593 (O_1593,N_29820,N_29790);
xnor UO_1594 (O_1594,N_29913,N_29949);
xnor UO_1595 (O_1595,N_29753,N_29520);
nand UO_1596 (O_1596,N_29673,N_29696);
nor UO_1597 (O_1597,N_29946,N_29595);
nand UO_1598 (O_1598,N_29722,N_29868);
or UO_1599 (O_1599,N_29709,N_29920);
nand UO_1600 (O_1600,N_29786,N_29860);
xor UO_1601 (O_1601,N_29744,N_29551);
xnor UO_1602 (O_1602,N_29852,N_29740);
xnor UO_1603 (O_1603,N_29692,N_29630);
nor UO_1604 (O_1604,N_29735,N_29866);
nor UO_1605 (O_1605,N_29678,N_29659);
nor UO_1606 (O_1606,N_29607,N_29770);
nor UO_1607 (O_1607,N_29787,N_29799);
xor UO_1608 (O_1608,N_29762,N_29931);
xor UO_1609 (O_1609,N_29680,N_29649);
xnor UO_1610 (O_1610,N_29752,N_29823);
or UO_1611 (O_1611,N_29804,N_29631);
nor UO_1612 (O_1612,N_29866,N_29933);
or UO_1613 (O_1613,N_29755,N_29711);
and UO_1614 (O_1614,N_29918,N_29809);
and UO_1615 (O_1615,N_29645,N_29563);
xnor UO_1616 (O_1616,N_29881,N_29757);
nand UO_1617 (O_1617,N_29620,N_29719);
and UO_1618 (O_1618,N_29604,N_29965);
and UO_1619 (O_1619,N_29820,N_29926);
or UO_1620 (O_1620,N_29835,N_29671);
nor UO_1621 (O_1621,N_29815,N_29786);
nand UO_1622 (O_1622,N_29556,N_29915);
nand UO_1623 (O_1623,N_29571,N_29869);
or UO_1624 (O_1624,N_29502,N_29531);
nor UO_1625 (O_1625,N_29929,N_29912);
nand UO_1626 (O_1626,N_29998,N_29713);
or UO_1627 (O_1627,N_29701,N_29573);
nand UO_1628 (O_1628,N_29662,N_29620);
nand UO_1629 (O_1629,N_29506,N_29877);
xor UO_1630 (O_1630,N_29744,N_29818);
xnor UO_1631 (O_1631,N_29625,N_29795);
nor UO_1632 (O_1632,N_29824,N_29878);
nor UO_1633 (O_1633,N_29831,N_29688);
and UO_1634 (O_1634,N_29666,N_29769);
nand UO_1635 (O_1635,N_29844,N_29818);
xnor UO_1636 (O_1636,N_29874,N_29681);
nor UO_1637 (O_1637,N_29638,N_29841);
nor UO_1638 (O_1638,N_29989,N_29852);
xnor UO_1639 (O_1639,N_29759,N_29929);
xor UO_1640 (O_1640,N_29952,N_29595);
nor UO_1641 (O_1641,N_29763,N_29607);
nor UO_1642 (O_1642,N_29661,N_29821);
nand UO_1643 (O_1643,N_29574,N_29588);
nor UO_1644 (O_1644,N_29941,N_29579);
xor UO_1645 (O_1645,N_29625,N_29617);
or UO_1646 (O_1646,N_29971,N_29522);
nor UO_1647 (O_1647,N_29989,N_29623);
and UO_1648 (O_1648,N_29740,N_29905);
xor UO_1649 (O_1649,N_29680,N_29523);
nand UO_1650 (O_1650,N_29985,N_29761);
nand UO_1651 (O_1651,N_29526,N_29737);
nand UO_1652 (O_1652,N_29554,N_29983);
nand UO_1653 (O_1653,N_29935,N_29953);
or UO_1654 (O_1654,N_29623,N_29895);
or UO_1655 (O_1655,N_29929,N_29875);
nand UO_1656 (O_1656,N_29658,N_29646);
and UO_1657 (O_1657,N_29741,N_29805);
or UO_1658 (O_1658,N_29806,N_29692);
nand UO_1659 (O_1659,N_29597,N_29724);
xnor UO_1660 (O_1660,N_29979,N_29835);
or UO_1661 (O_1661,N_29521,N_29793);
xnor UO_1662 (O_1662,N_29790,N_29764);
and UO_1663 (O_1663,N_29738,N_29945);
xnor UO_1664 (O_1664,N_29529,N_29735);
and UO_1665 (O_1665,N_29993,N_29902);
xor UO_1666 (O_1666,N_29814,N_29950);
and UO_1667 (O_1667,N_29765,N_29958);
or UO_1668 (O_1668,N_29728,N_29927);
xor UO_1669 (O_1669,N_29985,N_29913);
nor UO_1670 (O_1670,N_29783,N_29985);
nand UO_1671 (O_1671,N_29606,N_29785);
nand UO_1672 (O_1672,N_29567,N_29919);
or UO_1673 (O_1673,N_29680,N_29963);
or UO_1674 (O_1674,N_29734,N_29594);
or UO_1675 (O_1675,N_29590,N_29612);
xor UO_1676 (O_1676,N_29833,N_29748);
or UO_1677 (O_1677,N_29896,N_29990);
xnor UO_1678 (O_1678,N_29834,N_29901);
and UO_1679 (O_1679,N_29944,N_29612);
xor UO_1680 (O_1680,N_29562,N_29767);
xor UO_1681 (O_1681,N_29963,N_29518);
or UO_1682 (O_1682,N_29655,N_29669);
nor UO_1683 (O_1683,N_29926,N_29792);
or UO_1684 (O_1684,N_29925,N_29508);
or UO_1685 (O_1685,N_29872,N_29655);
xor UO_1686 (O_1686,N_29811,N_29981);
xnor UO_1687 (O_1687,N_29951,N_29956);
nor UO_1688 (O_1688,N_29809,N_29980);
nand UO_1689 (O_1689,N_29699,N_29816);
and UO_1690 (O_1690,N_29520,N_29716);
nor UO_1691 (O_1691,N_29884,N_29753);
or UO_1692 (O_1692,N_29700,N_29876);
nor UO_1693 (O_1693,N_29634,N_29544);
xnor UO_1694 (O_1694,N_29515,N_29928);
xor UO_1695 (O_1695,N_29699,N_29622);
nor UO_1696 (O_1696,N_29761,N_29737);
nand UO_1697 (O_1697,N_29855,N_29594);
and UO_1698 (O_1698,N_29545,N_29561);
nor UO_1699 (O_1699,N_29669,N_29943);
xnor UO_1700 (O_1700,N_29929,N_29784);
nand UO_1701 (O_1701,N_29717,N_29833);
nor UO_1702 (O_1702,N_29709,N_29703);
nand UO_1703 (O_1703,N_29636,N_29554);
or UO_1704 (O_1704,N_29971,N_29704);
and UO_1705 (O_1705,N_29943,N_29828);
nor UO_1706 (O_1706,N_29817,N_29804);
and UO_1707 (O_1707,N_29916,N_29612);
xor UO_1708 (O_1708,N_29694,N_29882);
xnor UO_1709 (O_1709,N_29757,N_29708);
xnor UO_1710 (O_1710,N_29928,N_29698);
nor UO_1711 (O_1711,N_29530,N_29787);
nor UO_1712 (O_1712,N_29517,N_29530);
nand UO_1713 (O_1713,N_29663,N_29558);
or UO_1714 (O_1714,N_29784,N_29558);
nor UO_1715 (O_1715,N_29779,N_29651);
and UO_1716 (O_1716,N_29564,N_29504);
or UO_1717 (O_1717,N_29694,N_29790);
nor UO_1718 (O_1718,N_29669,N_29749);
nand UO_1719 (O_1719,N_29846,N_29531);
or UO_1720 (O_1720,N_29886,N_29756);
nor UO_1721 (O_1721,N_29826,N_29819);
nor UO_1722 (O_1722,N_29961,N_29798);
nor UO_1723 (O_1723,N_29905,N_29893);
xor UO_1724 (O_1724,N_29865,N_29961);
nor UO_1725 (O_1725,N_29597,N_29956);
xnor UO_1726 (O_1726,N_29840,N_29940);
nand UO_1727 (O_1727,N_29710,N_29891);
nand UO_1728 (O_1728,N_29608,N_29862);
nor UO_1729 (O_1729,N_29974,N_29627);
or UO_1730 (O_1730,N_29581,N_29859);
nor UO_1731 (O_1731,N_29735,N_29977);
or UO_1732 (O_1732,N_29987,N_29780);
nor UO_1733 (O_1733,N_29560,N_29830);
or UO_1734 (O_1734,N_29880,N_29769);
or UO_1735 (O_1735,N_29836,N_29514);
nor UO_1736 (O_1736,N_29710,N_29733);
nand UO_1737 (O_1737,N_29753,N_29885);
nand UO_1738 (O_1738,N_29998,N_29927);
or UO_1739 (O_1739,N_29764,N_29640);
and UO_1740 (O_1740,N_29535,N_29989);
xnor UO_1741 (O_1741,N_29817,N_29541);
nor UO_1742 (O_1742,N_29616,N_29870);
nor UO_1743 (O_1743,N_29914,N_29856);
nand UO_1744 (O_1744,N_29584,N_29930);
or UO_1745 (O_1745,N_29588,N_29846);
nor UO_1746 (O_1746,N_29801,N_29812);
nor UO_1747 (O_1747,N_29579,N_29875);
and UO_1748 (O_1748,N_29643,N_29906);
or UO_1749 (O_1749,N_29812,N_29853);
or UO_1750 (O_1750,N_29717,N_29554);
or UO_1751 (O_1751,N_29639,N_29967);
and UO_1752 (O_1752,N_29939,N_29649);
or UO_1753 (O_1753,N_29593,N_29599);
or UO_1754 (O_1754,N_29674,N_29943);
xnor UO_1755 (O_1755,N_29501,N_29703);
nor UO_1756 (O_1756,N_29828,N_29518);
and UO_1757 (O_1757,N_29900,N_29741);
or UO_1758 (O_1758,N_29958,N_29718);
nor UO_1759 (O_1759,N_29793,N_29522);
xnor UO_1760 (O_1760,N_29625,N_29825);
and UO_1761 (O_1761,N_29527,N_29925);
nor UO_1762 (O_1762,N_29527,N_29531);
xnor UO_1763 (O_1763,N_29605,N_29742);
and UO_1764 (O_1764,N_29503,N_29975);
xor UO_1765 (O_1765,N_29935,N_29912);
or UO_1766 (O_1766,N_29793,N_29552);
xnor UO_1767 (O_1767,N_29981,N_29842);
or UO_1768 (O_1768,N_29938,N_29641);
nand UO_1769 (O_1769,N_29604,N_29983);
or UO_1770 (O_1770,N_29945,N_29540);
and UO_1771 (O_1771,N_29863,N_29985);
nand UO_1772 (O_1772,N_29686,N_29855);
and UO_1773 (O_1773,N_29751,N_29596);
nand UO_1774 (O_1774,N_29549,N_29924);
or UO_1775 (O_1775,N_29998,N_29701);
nand UO_1776 (O_1776,N_29515,N_29812);
nor UO_1777 (O_1777,N_29774,N_29660);
and UO_1778 (O_1778,N_29993,N_29747);
or UO_1779 (O_1779,N_29744,N_29629);
nand UO_1780 (O_1780,N_29905,N_29861);
or UO_1781 (O_1781,N_29965,N_29724);
and UO_1782 (O_1782,N_29705,N_29509);
or UO_1783 (O_1783,N_29553,N_29752);
nand UO_1784 (O_1784,N_29954,N_29703);
nor UO_1785 (O_1785,N_29536,N_29905);
xnor UO_1786 (O_1786,N_29622,N_29678);
nor UO_1787 (O_1787,N_29506,N_29858);
or UO_1788 (O_1788,N_29562,N_29575);
or UO_1789 (O_1789,N_29777,N_29522);
or UO_1790 (O_1790,N_29953,N_29631);
and UO_1791 (O_1791,N_29696,N_29632);
or UO_1792 (O_1792,N_29579,N_29945);
nand UO_1793 (O_1793,N_29745,N_29871);
xor UO_1794 (O_1794,N_29924,N_29706);
xnor UO_1795 (O_1795,N_29961,N_29561);
and UO_1796 (O_1796,N_29867,N_29910);
or UO_1797 (O_1797,N_29640,N_29847);
xor UO_1798 (O_1798,N_29510,N_29998);
nand UO_1799 (O_1799,N_29727,N_29617);
nor UO_1800 (O_1800,N_29761,N_29755);
nor UO_1801 (O_1801,N_29823,N_29500);
xor UO_1802 (O_1802,N_29625,N_29702);
xor UO_1803 (O_1803,N_29923,N_29550);
nor UO_1804 (O_1804,N_29884,N_29969);
xnor UO_1805 (O_1805,N_29685,N_29622);
xor UO_1806 (O_1806,N_29633,N_29648);
and UO_1807 (O_1807,N_29664,N_29577);
nand UO_1808 (O_1808,N_29734,N_29915);
nand UO_1809 (O_1809,N_29758,N_29885);
and UO_1810 (O_1810,N_29828,N_29815);
nand UO_1811 (O_1811,N_29517,N_29808);
xnor UO_1812 (O_1812,N_29635,N_29541);
and UO_1813 (O_1813,N_29877,N_29815);
nor UO_1814 (O_1814,N_29852,N_29831);
and UO_1815 (O_1815,N_29532,N_29839);
nand UO_1816 (O_1816,N_29652,N_29598);
xnor UO_1817 (O_1817,N_29588,N_29697);
nand UO_1818 (O_1818,N_29950,N_29668);
nand UO_1819 (O_1819,N_29850,N_29629);
xnor UO_1820 (O_1820,N_29813,N_29540);
or UO_1821 (O_1821,N_29855,N_29810);
and UO_1822 (O_1822,N_29652,N_29934);
nand UO_1823 (O_1823,N_29795,N_29687);
and UO_1824 (O_1824,N_29808,N_29874);
nor UO_1825 (O_1825,N_29785,N_29878);
and UO_1826 (O_1826,N_29840,N_29576);
and UO_1827 (O_1827,N_29723,N_29851);
or UO_1828 (O_1828,N_29933,N_29737);
or UO_1829 (O_1829,N_29694,N_29751);
nor UO_1830 (O_1830,N_29606,N_29694);
or UO_1831 (O_1831,N_29733,N_29927);
nor UO_1832 (O_1832,N_29855,N_29915);
xnor UO_1833 (O_1833,N_29680,N_29937);
nor UO_1834 (O_1834,N_29529,N_29574);
nand UO_1835 (O_1835,N_29808,N_29903);
nor UO_1836 (O_1836,N_29921,N_29693);
xor UO_1837 (O_1837,N_29614,N_29899);
and UO_1838 (O_1838,N_29796,N_29970);
or UO_1839 (O_1839,N_29895,N_29875);
or UO_1840 (O_1840,N_29700,N_29568);
nand UO_1841 (O_1841,N_29952,N_29761);
nor UO_1842 (O_1842,N_29918,N_29715);
xnor UO_1843 (O_1843,N_29706,N_29875);
nor UO_1844 (O_1844,N_29618,N_29715);
nand UO_1845 (O_1845,N_29707,N_29527);
xnor UO_1846 (O_1846,N_29835,N_29678);
or UO_1847 (O_1847,N_29958,N_29599);
xnor UO_1848 (O_1848,N_29521,N_29697);
nor UO_1849 (O_1849,N_29635,N_29550);
xnor UO_1850 (O_1850,N_29522,N_29958);
or UO_1851 (O_1851,N_29810,N_29804);
nand UO_1852 (O_1852,N_29534,N_29918);
nor UO_1853 (O_1853,N_29790,N_29846);
nand UO_1854 (O_1854,N_29560,N_29773);
nor UO_1855 (O_1855,N_29761,N_29565);
or UO_1856 (O_1856,N_29856,N_29523);
nand UO_1857 (O_1857,N_29503,N_29659);
nor UO_1858 (O_1858,N_29548,N_29587);
xnor UO_1859 (O_1859,N_29929,N_29697);
nand UO_1860 (O_1860,N_29604,N_29728);
nand UO_1861 (O_1861,N_29593,N_29604);
xor UO_1862 (O_1862,N_29843,N_29805);
nor UO_1863 (O_1863,N_29664,N_29843);
and UO_1864 (O_1864,N_29689,N_29820);
or UO_1865 (O_1865,N_29582,N_29716);
xor UO_1866 (O_1866,N_29597,N_29872);
nand UO_1867 (O_1867,N_29595,N_29637);
xnor UO_1868 (O_1868,N_29642,N_29848);
nand UO_1869 (O_1869,N_29830,N_29544);
xor UO_1870 (O_1870,N_29519,N_29946);
or UO_1871 (O_1871,N_29626,N_29612);
xor UO_1872 (O_1872,N_29597,N_29526);
and UO_1873 (O_1873,N_29664,N_29726);
and UO_1874 (O_1874,N_29779,N_29851);
nand UO_1875 (O_1875,N_29531,N_29743);
nand UO_1876 (O_1876,N_29892,N_29696);
or UO_1877 (O_1877,N_29983,N_29586);
xor UO_1878 (O_1878,N_29528,N_29593);
nand UO_1879 (O_1879,N_29980,N_29803);
nand UO_1880 (O_1880,N_29721,N_29588);
xnor UO_1881 (O_1881,N_29670,N_29673);
and UO_1882 (O_1882,N_29953,N_29520);
nor UO_1883 (O_1883,N_29944,N_29970);
xnor UO_1884 (O_1884,N_29858,N_29998);
nand UO_1885 (O_1885,N_29979,N_29523);
or UO_1886 (O_1886,N_29983,N_29858);
nor UO_1887 (O_1887,N_29741,N_29836);
nor UO_1888 (O_1888,N_29875,N_29532);
or UO_1889 (O_1889,N_29998,N_29800);
and UO_1890 (O_1890,N_29772,N_29593);
nor UO_1891 (O_1891,N_29770,N_29533);
nor UO_1892 (O_1892,N_29946,N_29597);
nand UO_1893 (O_1893,N_29670,N_29821);
nor UO_1894 (O_1894,N_29681,N_29976);
xnor UO_1895 (O_1895,N_29909,N_29571);
and UO_1896 (O_1896,N_29751,N_29565);
xor UO_1897 (O_1897,N_29825,N_29503);
and UO_1898 (O_1898,N_29780,N_29650);
nor UO_1899 (O_1899,N_29882,N_29781);
and UO_1900 (O_1900,N_29821,N_29735);
xnor UO_1901 (O_1901,N_29840,N_29887);
and UO_1902 (O_1902,N_29729,N_29568);
and UO_1903 (O_1903,N_29825,N_29519);
nand UO_1904 (O_1904,N_29835,N_29967);
xor UO_1905 (O_1905,N_29760,N_29694);
nor UO_1906 (O_1906,N_29533,N_29794);
nor UO_1907 (O_1907,N_29946,N_29721);
nand UO_1908 (O_1908,N_29671,N_29704);
nor UO_1909 (O_1909,N_29750,N_29565);
nand UO_1910 (O_1910,N_29778,N_29586);
nand UO_1911 (O_1911,N_29723,N_29688);
xor UO_1912 (O_1912,N_29705,N_29692);
and UO_1913 (O_1913,N_29881,N_29690);
xor UO_1914 (O_1914,N_29740,N_29983);
nand UO_1915 (O_1915,N_29968,N_29819);
or UO_1916 (O_1916,N_29872,N_29509);
or UO_1917 (O_1917,N_29510,N_29731);
nand UO_1918 (O_1918,N_29763,N_29585);
nor UO_1919 (O_1919,N_29645,N_29810);
xnor UO_1920 (O_1920,N_29613,N_29767);
and UO_1921 (O_1921,N_29977,N_29587);
xnor UO_1922 (O_1922,N_29723,N_29675);
and UO_1923 (O_1923,N_29644,N_29746);
and UO_1924 (O_1924,N_29876,N_29564);
xor UO_1925 (O_1925,N_29963,N_29687);
nand UO_1926 (O_1926,N_29896,N_29901);
nand UO_1927 (O_1927,N_29819,N_29851);
and UO_1928 (O_1928,N_29699,N_29564);
and UO_1929 (O_1929,N_29712,N_29618);
xnor UO_1930 (O_1930,N_29719,N_29536);
xnor UO_1931 (O_1931,N_29654,N_29707);
xnor UO_1932 (O_1932,N_29917,N_29747);
xor UO_1933 (O_1933,N_29950,N_29778);
xnor UO_1934 (O_1934,N_29614,N_29994);
nand UO_1935 (O_1935,N_29730,N_29894);
and UO_1936 (O_1936,N_29981,N_29992);
nand UO_1937 (O_1937,N_29531,N_29815);
or UO_1938 (O_1938,N_29677,N_29774);
and UO_1939 (O_1939,N_29977,N_29709);
or UO_1940 (O_1940,N_29908,N_29711);
xor UO_1941 (O_1941,N_29779,N_29863);
nor UO_1942 (O_1942,N_29945,N_29558);
or UO_1943 (O_1943,N_29901,N_29688);
nor UO_1944 (O_1944,N_29776,N_29675);
and UO_1945 (O_1945,N_29871,N_29857);
xor UO_1946 (O_1946,N_29651,N_29961);
xor UO_1947 (O_1947,N_29837,N_29931);
xor UO_1948 (O_1948,N_29540,N_29883);
or UO_1949 (O_1949,N_29503,N_29966);
or UO_1950 (O_1950,N_29538,N_29670);
and UO_1951 (O_1951,N_29878,N_29570);
or UO_1952 (O_1952,N_29939,N_29540);
or UO_1953 (O_1953,N_29695,N_29894);
or UO_1954 (O_1954,N_29595,N_29842);
and UO_1955 (O_1955,N_29833,N_29596);
xnor UO_1956 (O_1956,N_29592,N_29943);
or UO_1957 (O_1957,N_29927,N_29912);
nand UO_1958 (O_1958,N_29548,N_29913);
nor UO_1959 (O_1959,N_29897,N_29510);
nor UO_1960 (O_1960,N_29844,N_29893);
nand UO_1961 (O_1961,N_29768,N_29904);
xor UO_1962 (O_1962,N_29557,N_29758);
nor UO_1963 (O_1963,N_29779,N_29978);
nand UO_1964 (O_1964,N_29704,N_29834);
nor UO_1965 (O_1965,N_29689,N_29855);
xor UO_1966 (O_1966,N_29677,N_29727);
nand UO_1967 (O_1967,N_29943,N_29886);
xor UO_1968 (O_1968,N_29590,N_29967);
nor UO_1969 (O_1969,N_29757,N_29905);
nand UO_1970 (O_1970,N_29908,N_29641);
or UO_1971 (O_1971,N_29656,N_29552);
or UO_1972 (O_1972,N_29814,N_29863);
or UO_1973 (O_1973,N_29653,N_29999);
nor UO_1974 (O_1974,N_29768,N_29583);
and UO_1975 (O_1975,N_29845,N_29772);
or UO_1976 (O_1976,N_29599,N_29849);
or UO_1977 (O_1977,N_29756,N_29918);
nand UO_1978 (O_1978,N_29713,N_29764);
xor UO_1979 (O_1979,N_29848,N_29867);
nand UO_1980 (O_1980,N_29885,N_29957);
nand UO_1981 (O_1981,N_29930,N_29782);
nor UO_1982 (O_1982,N_29842,N_29733);
or UO_1983 (O_1983,N_29899,N_29852);
xor UO_1984 (O_1984,N_29678,N_29763);
xor UO_1985 (O_1985,N_29603,N_29999);
and UO_1986 (O_1986,N_29814,N_29917);
and UO_1987 (O_1987,N_29985,N_29878);
nand UO_1988 (O_1988,N_29574,N_29517);
or UO_1989 (O_1989,N_29982,N_29922);
and UO_1990 (O_1990,N_29978,N_29733);
xnor UO_1991 (O_1991,N_29708,N_29538);
xor UO_1992 (O_1992,N_29916,N_29902);
nor UO_1993 (O_1993,N_29656,N_29572);
and UO_1994 (O_1994,N_29886,N_29924);
nand UO_1995 (O_1995,N_29806,N_29511);
and UO_1996 (O_1996,N_29551,N_29886);
or UO_1997 (O_1997,N_29745,N_29867);
xor UO_1998 (O_1998,N_29579,N_29898);
nand UO_1999 (O_1999,N_29804,N_29797);
xnor UO_2000 (O_2000,N_29862,N_29990);
xnor UO_2001 (O_2001,N_29857,N_29806);
nand UO_2002 (O_2002,N_29895,N_29885);
or UO_2003 (O_2003,N_29605,N_29693);
nor UO_2004 (O_2004,N_29661,N_29838);
nor UO_2005 (O_2005,N_29953,N_29565);
and UO_2006 (O_2006,N_29850,N_29611);
and UO_2007 (O_2007,N_29996,N_29978);
or UO_2008 (O_2008,N_29993,N_29646);
nor UO_2009 (O_2009,N_29706,N_29911);
and UO_2010 (O_2010,N_29641,N_29550);
xor UO_2011 (O_2011,N_29573,N_29676);
or UO_2012 (O_2012,N_29938,N_29596);
xor UO_2013 (O_2013,N_29797,N_29805);
and UO_2014 (O_2014,N_29629,N_29927);
or UO_2015 (O_2015,N_29715,N_29811);
nor UO_2016 (O_2016,N_29717,N_29939);
nand UO_2017 (O_2017,N_29652,N_29553);
xnor UO_2018 (O_2018,N_29802,N_29749);
nand UO_2019 (O_2019,N_29776,N_29722);
nand UO_2020 (O_2020,N_29905,N_29573);
or UO_2021 (O_2021,N_29569,N_29977);
nand UO_2022 (O_2022,N_29704,N_29572);
nand UO_2023 (O_2023,N_29991,N_29595);
or UO_2024 (O_2024,N_29550,N_29723);
and UO_2025 (O_2025,N_29776,N_29863);
xor UO_2026 (O_2026,N_29683,N_29770);
nand UO_2027 (O_2027,N_29733,N_29756);
nand UO_2028 (O_2028,N_29739,N_29894);
nand UO_2029 (O_2029,N_29787,N_29557);
or UO_2030 (O_2030,N_29567,N_29569);
nand UO_2031 (O_2031,N_29862,N_29815);
nor UO_2032 (O_2032,N_29835,N_29841);
xnor UO_2033 (O_2033,N_29595,N_29522);
and UO_2034 (O_2034,N_29891,N_29882);
or UO_2035 (O_2035,N_29745,N_29849);
nand UO_2036 (O_2036,N_29747,N_29574);
xor UO_2037 (O_2037,N_29974,N_29726);
nand UO_2038 (O_2038,N_29943,N_29876);
nor UO_2039 (O_2039,N_29696,N_29732);
or UO_2040 (O_2040,N_29671,N_29944);
and UO_2041 (O_2041,N_29675,N_29783);
or UO_2042 (O_2042,N_29889,N_29522);
and UO_2043 (O_2043,N_29998,N_29863);
or UO_2044 (O_2044,N_29897,N_29953);
nor UO_2045 (O_2045,N_29979,N_29929);
and UO_2046 (O_2046,N_29771,N_29692);
nand UO_2047 (O_2047,N_29913,N_29743);
or UO_2048 (O_2048,N_29817,N_29561);
xnor UO_2049 (O_2049,N_29999,N_29644);
and UO_2050 (O_2050,N_29693,N_29938);
xor UO_2051 (O_2051,N_29700,N_29921);
nand UO_2052 (O_2052,N_29777,N_29960);
xnor UO_2053 (O_2053,N_29619,N_29523);
xnor UO_2054 (O_2054,N_29810,N_29799);
nor UO_2055 (O_2055,N_29592,N_29893);
nand UO_2056 (O_2056,N_29793,N_29908);
or UO_2057 (O_2057,N_29535,N_29658);
xor UO_2058 (O_2058,N_29825,N_29717);
nor UO_2059 (O_2059,N_29898,N_29946);
or UO_2060 (O_2060,N_29924,N_29533);
nand UO_2061 (O_2061,N_29895,N_29918);
nand UO_2062 (O_2062,N_29923,N_29786);
nor UO_2063 (O_2063,N_29867,N_29766);
and UO_2064 (O_2064,N_29508,N_29933);
nor UO_2065 (O_2065,N_29856,N_29939);
and UO_2066 (O_2066,N_29941,N_29677);
nor UO_2067 (O_2067,N_29741,N_29970);
nor UO_2068 (O_2068,N_29996,N_29843);
nand UO_2069 (O_2069,N_29601,N_29919);
nand UO_2070 (O_2070,N_29506,N_29737);
and UO_2071 (O_2071,N_29878,N_29955);
nor UO_2072 (O_2072,N_29612,N_29772);
nor UO_2073 (O_2073,N_29941,N_29738);
xnor UO_2074 (O_2074,N_29931,N_29825);
and UO_2075 (O_2075,N_29554,N_29961);
nand UO_2076 (O_2076,N_29965,N_29708);
and UO_2077 (O_2077,N_29834,N_29891);
nor UO_2078 (O_2078,N_29540,N_29835);
nor UO_2079 (O_2079,N_29678,N_29684);
xnor UO_2080 (O_2080,N_29983,N_29967);
xnor UO_2081 (O_2081,N_29541,N_29699);
nor UO_2082 (O_2082,N_29555,N_29893);
and UO_2083 (O_2083,N_29530,N_29744);
nor UO_2084 (O_2084,N_29944,N_29776);
nand UO_2085 (O_2085,N_29864,N_29754);
and UO_2086 (O_2086,N_29749,N_29792);
nand UO_2087 (O_2087,N_29563,N_29885);
or UO_2088 (O_2088,N_29514,N_29950);
nor UO_2089 (O_2089,N_29574,N_29774);
xnor UO_2090 (O_2090,N_29935,N_29957);
and UO_2091 (O_2091,N_29665,N_29925);
nand UO_2092 (O_2092,N_29520,N_29720);
xnor UO_2093 (O_2093,N_29722,N_29558);
nand UO_2094 (O_2094,N_29862,N_29941);
nor UO_2095 (O_2095,N_29585,N_29925);
and UO_2096 (O_2096,N_29511,N_29640);
nor UO_2097 (O_2097,N_29703,N_29570);
nand UO_2098 (O_2098,N_29984,N_29909);
and UO_2099 (O_2099,N_29982,N_29862);
and UO_2100 (O_2100,N_29996,N_29904);
or UO_2101 (O_2101,N_29707,N_29822);
nand UO_2102 (O_2102,N_29580,N_29640);
xor UO_2103 (O_2103,N_29600,N_29523);
nand UO_2104 (O_2104,N_29735,N_29804);
nor UO_2105 (O_2105,N_29514,N_29838);
nor UO_2106 (O_2106,N_29986,N_29980);
xnor UO_2107 (O_2107,N_29610,N_29773);
xnor UO_2108 (O_2108,N_29821,N_29785);
nor UO_2109 (O_2109,N_29834,N_29983);
and UO_2110 (O_2110,N_29514,N_29715);
nand UO_2111 (O_2111,N_29696,N_29913);
and UO_2112 (O_2112,N_29968,N_29826);
nand UO_2113 (O_2113,N_29892,N_29821);
and UO_2114 (O_2114,N_29623,N_29843);
nor UO_2115 (O_2115,N_29590,N_29631);
and UO_2116 (O_2116,N_29866,N_29794);
or UO_2117 (O_2117,N_29997,N_29878);
xnor UO_2118 (O_2118,N_29832,N_29583);
or UO_2119 (O_2119,N_29839,N_29740);
nor UO_2120 (O_2120,N_29690,N_29969);
and UO_2121 (O_2121,N_29918,N_29646);
xor UO_2122 (O_2122,N_29509,N_29540);
and UO_2123 (O_2123,N_29990,N_29624);
or UO_2124 (O_2124,N_29821,N_29504);
nand UO_2125 (O_2125,N_29715,N_29698);
xnor UO_2126 (O_2126,N_29913,N_29835);
xnor UO_2127 (O_2127,N_29727,N_29858);
and UO_2128 (O_2128,N_29910,N_29874);
and UO_2129 (O_2129,N_29673,N_29759);
and UO_2130 (O_2130,N_29715,N_29690);
and UO_2131 (O_2131,N_29972,N_29722);
or UO_2132 (O_2132,N_29596,N_29995);
and UO_2133 (O_2133,N_29532,N_29813);
nand UO_2134 (O_2134,N_29583,N_29631);
nand UO_2135 (O_2135,N_29858,N_29997);
nand UO_2136 (O_2136,N_29582,N_29608);
or UO_2137 (O_2137,N_29930,N_29558);
and UO_2138 (O_2138,N_29804,N_29703);
nor UO_2139 (O_2139,N_29976,N_29579);
nand UO_2140 (O_2140,N_29769,N_29534);
and UO_2141 (O_2141,N_29669,N_29578);
nor UO_2142 (O_2142,N_29514,N_29548);
xor UO_2143 (O_2143,N_29589,N_29727);
nor UO_2144 (O_2144,N_29813,N_29991);
nand UO_2145 (O_2145,N_29702,N_29576);
and UO_2146 (O_2146,N_29766,N_29933);
and UO_2147 (O_2147,N_29919,N_29556);
nor UO_2148 (O_2148,N_29677,N_29534);
xnor UO_2149 (O_2149,N_29503,N_29666);
xor UO_2150 (O_2150,N_29691,N_29902);
or UO_2151 (O_2151,N_29838,N_29568);
or UO_2152 (O_2152,N_29754,N_29569);
or UO_2153 (O_2153,N_29629,N_29884);
and UO_2154 (O_2154,N_29921,N_29634);
and UO_2155 (O_2155,N_29784,N_29532);
xnor UO_2156 (O_2156,N_29745,N_29853);
nand UO_2157 (O_2157,N_29931,N_29962);
or UO_2158 (O_2158,N_29667,N_29812);
nand UO_2159 (O_2159,N_29920,N_29836);
nand UO_2160 (O_2160,N_29816,N_29683);
nor UO_2161 (O_2161,N_29542,N_29705);
nand UO_2162 (O_2162,N_29535,N_29799);
or UO_2163 (O_2163,N_29576,N_29633);
xnor UO_2164 (O_2164,N_29812,N_29773);
and UO_2165 (O_2165,N_29892,N_29846);
nor UO_2166 (O_2166,N_29645,N_29758);
nand UO_2167 (O_2167,N_29874,N_29863);
and UO_2168 (O_2168,N_29617,N_29551);
and UO_2169 (O_2169,N_29840,N_29971);
nor UO_2170 (O_2170,N_29967,N_29602);
nor UO_2171 (O_2171,N_29924,N_29747);
xnor UO_2172 (O_2172,N_29586,N_29995);
and UO_2173 (O_2173,N_29940,N_29541);
and UO_2174 (O_2174,N_29803,N_29518);
and UO_2175 (O_2175,N_29724,N_29618);
and UO_2176 (O_2176,N_29868,N_29823);
xor UO_2177 (O_2177,N_29526,N_29687);
nand UO_2178 (O_2178,N_29619,N_29561);
nand UO_2179 (O_2179,N_29707,N_29501);
and UO_2180 (O_2180,N_29859,N_29845);
nand UO_2181 (O_2181,N_29601,N_29716);
and UO_2182 (O_2182,N_29868,N_29924);
xnor UO_2183 (O_2183,N_29554,N_29899);
nand UO_2184 (O_2184,N_29950,N_29798);
xor UO_2185 (O_2185,N_29833,N_29621);
and UO_2186 (O_2186,N_29676,N_29757);
or UO_2187 (O_2187,N_29976,N_29745);
nor UO_2188 (O_2188,N_29890,N_29568);
nand UO_2189 (O_2189,N_29765,N_29810);
nand UO_2190 (O_2190,N_29526,N_29704);
or UO_2191 (O_2191,N_29510,N_29970);
or UO_2192 (O_2192,N_29601,N_29659);
and UO_2193 (O_2193,N_29725,N_29509);
xnor UO_2194 (O_2194,N_29561,N_29884);
or UO_2195 (O_2195,N_29563,N_29715);
nand UO_2196 (O_2196,N_29793,N_29858);
xor UO_2197 (O_2197,N_29601,N_29986);
and UO_2198 (O_2198,N_29666,N_29837);
or UO_2199 (O_2199,N_29652,N_29570);
and UO_2200 (O_2200,N_29657,N_29865);
xor UO_2201 (O_2201,N_29872,N_29693);
and UO_2202 (O_2202,N_29992,N_29688);
and UO_2203 (O_2203,N_29645,N_29738);
nor UO_2204 (O_2204,N_29885,N_29733);
and UO_2205 (O_2205,N_29620,N_29644);
and UO_2206 (O_2206,N_29930,N_29945);
xor UO_2207 (O_2207,N_29731,N_29602);
xor UO_2208 (O_2208,N_29956,N_29590);
nor UO_2209 (O_2209,N_29731,N_29969);
nand UO_2210 (O_2210,N_29979,N_29558);
nand UO_2211 (O_2211,N_29974,N_29857);
and UO_2212 (O_2212,N_29884,N_29515);
nor UO_2213 (O_2213,N_29760,N_29580);
or UO_2214 (O_2214,N_29814,N_29682);
nand UO_2215 (O_2215,N_29918,N_29762);
nand UO_2216 (O_2216,N_29680,N_29526);
xor UO_2217 (O_2217,N_29996,N_29752);
xnor UO_2218 (O_2218,N_29797,N_29732);
xor UO_2219 (O_2219,N_29817,N_29576);
xnor UO_2220 (O_2220,N_29569,N_29607);
nand UO_2221 (O_2221,N_29518,N_29935);
nand UO_2222 (O_2222,N_29931,N_29844);
xor UO_2223 (O_2223,N_29709,N_29562);
xnor UO_2224 (O_2224,N_29818,N_29720);
xor UO_2225 (O_2225,N_29963,N_29562);
nand UO_2226 (O_2226,N_29687,N_29552);
and UO_2227 (O_2227,N_29743,N_29510);
nor UO_2228 (O_2228,N_29767,N_29990);
nor UO_2229 (O_2229,N_29909,N_29809);
or UO_2230 (O_2230,N_29915,N_29962);
nand UO_2231 (O_2231,N_29660,N_29506);
nor UO_2232 (O_2232,N_29522,N_29664);
nand UO_2233 (O_2233,N_29757,N_29553);
nor UO_2234 (O_2234,N_29516,N_29866);
or UO_2235 (O_2235,N_29918,N_29884);
xor UO_2236 (O_2236,N_29809,N_29970);
nor UO_2237 (O_2237,N_29818,N_29908);
xor UO_2238 (O_2238,N_29557,N_29824);
xor UO_2239 (O_2239,N_29777,N_29563);
nor UO_2240 (O_2240,N_29560,N_29764);
or UO_2241 (O_2241,N_29694,N_29535);
and UO_2242 (O_2242,N_29613,N_29928);
nor UO_2243 (O_2243,N_29910,N_29651);
and UO_2244 (O_2244,N_29544,N_29723);
and UO_2245 (O_2245,N_29979,N_29571);
and UO_2246 (O_2246,N_29802,N_29613);
nor UO_2247 (O_2247,N_29884,N_29900);
and UO_2248 (O_2248,N_29838,N_29924);
xnor UO_2249 (O_2249,N_29997,N_29693);
and UO_2250 (O_2250,N_29747,N_29505);
nand UO_2251 (O_2251,N_29711,N_29856);
nand UO_2252 (O_2252,N_29922,N_29856);
xnor UO_2253 (O_2253,N_29896,N_29710);
or UO_2254 (O_2254,N_29699,N_29725);
xor UO_2255 (O_2255,N_29681,N_29716);
or UO_2256 (O_2256,N_29763,N_29737);
xor UO_2257 (O_2257,N_29764,N_29878);
or UO_2258 (O_2258,N_29693,N_29788);
and UO_2259 (O_2259,N_29670,N_29632);
xnor UO_2260 (O_2260,N_29817,N_29735);
and UO_2261 (O_2261,N_29892,N_29648);
or UO_2262 (O_2262,N_29875,N_29628);
and UO_2263 (O_2263,N_29602,N_29559);
or UO_2264 (O_2264,N_29626,N_29706);
nand UO_2265 (O_2265,N_29673,N_29886);
nor UO_2266 (O_2266,N_29763,N_29728);
or UO_2267 (O_2267,N_29746,N_29737);
nand UO_2268 (O_2268,N_29801,N_29738);
nor UO_2269 (O_2269,N_29776,N_29818);
or UO_2270 (O_2270,N_29560,N_29843);
nor UO_2271 (O_2271,N_29827,N_29908);
and UO_2272 (O_2272,N_29652,N_29676);
or UO_2273 (O_2273,N_29775,N_29719);
and UO_2274 (O_2274,N_29878,N_29987);
or UO_2275 (O_2275,N_29706,N_29688);
xnor UO_2276 (O_2276,N_29998,N_29793);
or UO_2277 (O_2277,N_29703,N_29775);
nand UO_2278 (O_2278,N_29688,N_29993);
xnor UO_2279 (O_2279,N_29687,N_29939);
or UO_2280 (O_2280,N_29577,N_29712);
nor UO_2281 (O_2281,N_29852,N_29914);
and UO_2282 (O_2282,N_29897,N_29892);
or UO_2283 (O_2283,N_29553,N_29666);
or UO_2284 (O_2284,N_29761,N_29601);
nand UO_2285 (O_2285,N_29769,N_29625);
nor UO_2286 (O_2286,N_29784,N_29525);
nor UO_2287 (O_2287,N_29721,N_29889);
nor UO_2288 (O_2288,N_29554,N_29515);
nand UO_2289 (O_2289,N_29955,N_29742);
and UO_2290 (O_2290,N_29647,N_29768);
or UO_2291 (O_2291,N_29681,N_29845);
nand UO_2292 (O_2292,N_29646,N_29780);
or UO_2293 (O_2293,N_29954,N_29826);
nor UO_2294 (O_2294,N_29560,N_29949);
or UO_2295 (O_2295,N_29919,N_29796);
and UO_2296 (O_2296,N_29968,N_29825);
nor UO_2297 (O_2297,N_29853,N_29903);
nand UO_2298 (O_2298,N_29984,N_29894);
and UO_2299 (O_2299,N_29558,N_29767);
nand UO_2300 (O_2300,N_29877,N_29919);
nand UO_2301 (O_2301,N_29646,N_29655);
or UO_2302 (O_2302,N_29694,N_29886);
or UO_2303 (O_2303,N_29957,N_29771);
nor UO_2304 (O_2304,N_29959,N_29726);
nor UO_2305 (O_2305,N_29749,N_29937);
xor UO_2306 (O_2306,N_29856,N_29616);
xor UO_2307 (O_2307,N_29585,N_29511);
nor UO_2308 (O_2308,N_29666,N_29908);
and UO_2309 (O_2309,N_29914,N_29747);
xnor UO_2310 (O_2310,N_29884,N_29887);
and UO_2311 (O_2311,N_29745,N_29870);
and UO_2312 (O_2312,N_29956,N_29561);
nor UO_2313 (O_2313,N_29577,N_29551);
and UO_2314 (O_2314,N_29654,N_29764);
nor UO_2315 (O_2315,N_29742,N_29843);
xnor UO_2316 (O_2316,N_29683,N_29665);
nand UO_2317 (O_2317,N_29800,N_29591);
and UO_2318 (O_2318,N_29661,N_29672);
nor UO_2319 (O_2319,N_29698,N_29545);
nor UO_2320 (O_2320,N_29585,N_29659);
nor UO_2321 (O_2321,N_29997,N_29874);
nand UO_2322 (O_2322,N_29652,N_29879);
and UO_2323 (O_2323,N_29983,N_29553);
or UO_2324 (O_2324,N_29645,N_29528);
and UO_2325 (O_2325,N_29755,N_29725);
nand UO_2326 (O_2326,N_29940,N_29950);
or UO_2327 (O_2327,N_29971,N_29675);
or UO_2328 (O_2328,N_29777,N_29833);
nand UO_2329 (O_2329,N_29871,N_29943);
and UO_2330 (O_2330,N_29954,N_29818);
nand UO_2331 (O_2331,N_29787,N_29969);
and UO_2332 (O_2332,N_29872,N_29691);
or UO_2333 (O_2333,N_29821,N_29755);
nor UO_2334 (O_2334,N_29829,N_29863);
or UO_2335 (O_2335,N_29978,N_29787);
or UO_2336 (O_2336,N_29616,N_29812);
nand UO_2337 (O_2337,N_29624,N_29542);
nand UO_2338 (O_2338,N_29562,N_29715);
or UO_2339 (O_2339,N_29907,N_29576);
and UO_2340 (O_2340,N_29949,N_29626);
xnor UO_2341 (O_2341,N_29670,N_29928);
and UO_2342 (O_2342,N_29987,N_29508);
xnor UO_2343 (O_2343,N_29754,N_29517);
xor UO_2344 (O_2344,N_29723,N_29726);
nand UO_2345 (O_2345,N_29879,N_29955);
nand UO_2346 (O_2346,N_29587,N_29644);
xor UO_2347 (O_2347,N_29580,N_29712);
or UO_2348 (O_2348,N_29675,N_29604);
nor UO_2349 (O_2349,N_29685,N_29937);
xnor UO_2350 (O_2350,N_29992,N_29862);
nand UO_2351 (O_2351,N_29741,N_29977);
or UO_2352 (O_2352,N_29942,N_29787);
xnor UO_2353 (O_2353,N_29590,N_29522);
nand UO_2354 (O_2354,N_29562,N_29794);
nor UO_2355 (O_2355,N_29870,N_29535);
nand UO_2356 (O_2356,N_29684,N_29993);
nor UO_2357 (O_2357,N_29549,N_29981);
nor UO_2358 (O_2358,N_29907,N_29664);
nor UO_2359 (O_2359,N_29726,N_29509);
xnor UO_2360 (O_2360,N_29814,N_29878);
nand UO_2361 (O_2361,N_29599,N_29776);
nor UO_2362 (O_2362,N_29710,N_29964);
and UO_2363 (O_2363,N_29783,N_29961);
or UO_2364 (O_2364,N_29764,N_29646);
xnor UO_2365 (O_2365,N_29821,N_29803);
and UO_2366 (O_2366,N_29861,N_29529);
xor UO_2367 (O_2367,N_29630,N_29681);
and UO_2368 (O_2368,N_29754,N_29583);
xor UO_2369 (O_2369,N_29738,N_29993);
nor UO_2370 (O_2370,N_29841,N_29676);
and UO_2371 (O_2371,N_29556,N_29642);
or UO_2372 (O_2372,N_29684,N_29970);
nand UO_2373 (O_2373,N_29560,N_29969);
nand UO_2374 (O_2374,N_29543,N_29867);
nand UO_2375 (O_2375,N_29998,N_29563);
nor UO_2376 (O_2376,N_29753,N_29927);
and UO_2377 (O_2377,N_29598,N_29897);
nor UO_2378 (O_2378,N_29959,N_29606);
or UO_2379 (O_2379,N_29887,N_29806);
or UO_2380 (O_2380,N_29951,N_29678);
or UO_2381 (O_2381,N_29688,N_29556);
and UO_2382 (O_2382,N_29797,N_29825);
and UO_2383 (O_2383,N_29945,N_29653);
or UO_2384 (O_2384,N_29648,N_29580);
or UO_2385 (O_2385,N_29604,N_29630);
and UO_2386 (O_2386,N_29888,N_29997);
nand UO_2387 (O_2387,N_29577,N_29964);
and UO_2388 (O_2388,N_29714,N_29523);
nand UO_2389 (O_2389,N_29956,N_29815);
nor UO_2390 (O_2390,N_29820,N_29623);
or UO_2391 (O_2391,N_29716,N_29524);
nor UO_2392 (O_2392,N_29908,N_29951);
or UO_2393 (O_2393,N_29982,N_29689);
nand UO_2394 (O_2394,N_29846,N_29553);
nand UO_2395 (O_2395,N_29669,N_29626);
nor UO_2396 (O_2396,N_29923,N_29844);
nand UO_2397 (O_2397,N_29843,N_29642);
and UO_2398 (O_2398,N_29773,N_29912);
nand UO_2399 (O_2399,N_29904,N_29592);
or UO_2400 (O_2400,N_29790,N_29574);
xor UO_2401 (O_2401,N_29971,N_29631);
or UO_2402 (O_2402,N_29676,N_29814);
or UO_2403 (O_2403,N_29762,N_29648);
and UO_2404 (O_2404,N_29551,N_29985);
nor UO_2405 (O_2405,N_29968,N_29597);
or UO_2406 (O_2406,N_29650,N_29966);
xnor UO_2407 (O_2407,N_29627,N_29849);
nand UO_2408 (O_2408,N_29643,N_29992);
nand UO_2409 (O_2409,N_29819,N_29589);
xnor UO_2410 (O_2410,N_29869,N_29568);
and UO_2411 (O_2411,N_29707,N_29540);
and UO_2412 (O_2412,N_29803,N_29741);
nand UO_2413 (O_2413,N_29888,N_29563);
nor UO_2414 (O_2414,N_29594,N_29633);
nand UO_2415 (O_2415,N_29887,N_29870);
nand UO_2416 (O_2416,N_29855,N_29562);
nor UO_2417 (O_2417,N_29656,N_29777);
nor UO_2418 (O_2418,N_29951,N_29538);
xnor UO_2419 (O_2419,N_29630,N_29856);
nand UO_2420 (O_2420,N_29791,N_29842);
or UO_2421 (O_2421,N_29891,N_29697);
or UO_2422 (O_2422,N_29914,N_29756);
and UO_2423 (O_2423,N_29845,N_29888);
nand UO_2424 (O_2424,N_29980,N_29903);
nand UO_2425 (O_2425,N_29783,N_29611);
nor UO_2426 (O_2426,N_29949,N_29989);
and UO_2427 (O_2427,N_29956,N_29706);
and UO_2428 (O_2428,N_29616,N_29539);
nor UO_2429 (O_2429,N_29854,N_29923);
nand UO_2430 (O_2430,N_29601,N_29782);
or UO_2431 (O_2431,N_29844,N_29660);
xnor UO_2432 (O_2432,N_29607,N_29978);
nand UO_2433 (O_2433,N_29822,N_29807);
or UO_2434 (O_2434,N_29686,N_29708);
nor UO_2435 (O_2435,N_29987,N_29865);
and UO_2436 (O_2436,N_29554,N_29604);
or UO_2437 (O_2437,N_29542,N_29999);
xor UO_2438 (O_2438,N_29991,N_29784);
xor UO_2439 (O_2439,N_29832,N_29572);
nand UO_2440 (O_2440,N_29866,N_29777);
and UO_2441 (O_2441,N_29751,N_29697);
nor UO_2442 (O_2442,N_29529,N_29626);
and UO_2443 (O_2443,N_29793,N_29519);
or UO_2444 (O_2444,N_29581,N_29842);
nor UO_2445 (O_2445,N_29894,N_29557);
and UO_2446 (O_2446,N_29684,N_29738);
and UO_2447 (O_2447,N_29543,N_29546);
or UO_2448 (O_2448,N_29632,N_29541);
and UO_2449 (O_2449,N_29977,N_29547);
nor UO_2450 (O_2450,N_29772,N_29611);
and UO_2451 (O_2451,N_29578,N_29819);
xnor UO_2452 (O_2452,N_29666,N_29813);
or UO_2453 (O_2453,N_29810,N_29643);
nand UO_2454 (O_2454,N_29607,N_29741);
or UO_2455 (O_2455,N_29693,N_29610);
or UO_2456 (O_2456,N_29705,N_29970);
or UO_2457 (O_2457,N_29612,N_29931);
xor UO_2458 (O_2458,N_29980,N_29699);
xor UO_2459 (O_2459,N_29838,N_29506);
xor UO_2460 (O_2460,N_29900,N_29675);
nand UO_2461 (O_2461,N_29524,N_29955);
nor UO_2462 (O_2462,N_29559,N_29946);
and UO_2463 (O_2463,N_29647,N_29508);
and UO_2464 (O_2464,N_29986,N_29996);
and UO_2465 (O_2465,N_29885,N_29672);
nor UO_2466 (O_2466,N_29766,N_29978);
nand UO_2467 (O_2467,N_29603,N_29954);
or UO_2468 (O_2468,N_29609,N_29698);
or UO_2469 (O_2469,N_29637,N_29514);
nor UO_2470 (O_2470,N_29976,N_29890);
or UO_2471 (O_2471,N_29814,N_29699);
xor UO_2472 (O_2472,N_29658,N_29606);
nor UO_2473 (O_2473,N_29517,N_29643);
xor UO_2474 (O_2474,N_29990,N_29946);
xnor UO_2475 (O_2475,N_29757,N_29574);
or UO_2476 (O_2476,N_29618,N_29510);
nand UO_2477 (O_2477,N_29696,N_29834);
and UO_2478 (O_2478,N_29854,N_29555);
and UO_2479 (O_2479,N_29730,N_29719);
or UO_2480 (O_2480,N_29908,N_29661);
or UO_2481 (O_2481,N_29985,N_29904);
or UO_2482 (O_2482,N_29727,N_29650);
nor UO_2483 (O_2483,N_29979,N_29762);
nor UO_2484 (O_2484,N_29502,N_29872);
nand UO_2485 (O_2485,N_29759,N_29576);
nand UO_2486 (O_2486,N_29897,N_29877);
nand UO_2487 (O_2487,N_29690,N_29643);
nor UO_2488 (O_2488,N_29878,N_29915);
or UO_2489 (O_2489,N_29620,N_29612);
xnor UO_2490 (O_2490,N_29562,N_29780);
nand UO_2491 (O_2491,N_29958,N_29961);
nor UO_2492 (O_2492,N_29531,N_29996);
nor UO_2493 (O_2493,N_29682,N_29554);
xnor UO_2494 (O_2494,N_29694,N_29832);
xor UO_2495 (O_2495,N_29855,N_29647);
xnor UO_2496 (O_2496,N_29539,N_29745);
nor UO_2497 (O_2497,N_29789,N_29682);
nand UO_2498 (O_2498,N_29696,N_29891);
nor UO_2499 (O_2499,N_29835,N_29718);
nand UO_2500 (O_2500,N_29648,N_29586);
or UO_2501 (O_2501,N_29786,N_29640);
or UO_2502 (O_2502,N_29836,N_29686);
and UO_2503 (O_2503,N_29636,N_29665);
xnor UO_2504 (O_2504,N_29572,N_29570);
or UO_2505 (O_2505,N_29873,N_29987);
or UO_2506 (O_2506,N_29762,N_29813);
and UO_2507 (O_2507,N_29859,N_29557);
or UO_2508 (O_2508,N_29806,N_29747);
nand UO_2509 (O_2509,N_29882,N_29905);
nand UO_2510 (O_2510,N_29845,N_29800);
nor UO_2511 (O_2511,N_29845,N_29649);
and UO_2512 (O_2512,N_29577,N_29779);
and UO_2513 (O_2513,N_29581,N_29791);
xor UO_2514 (O_2514,N_29540,N_29642);
xnor UO_2515 (O_2515,N_29825,N_29942);
or UO_2516 (O_2516,N_29811,N_29707);
or UO_2517 (O_2517,N_29976,N_29906);
nor UO_2518 (O_2518,N_29970,N_29631);
nor UO_2519 (O_2519,N_29723,N_29745);
xnor UO_2520 (O_2520,N_29642,N_29978);
nor UO_2521 (O_2521,N_29973,N_29879);
xor UO_2522 (O_2522,N_29851,N_29538);
xnor UO_2523 (O_2523,N_29700,N_29627);
xor UO_2524 (O_2524,N_29661,N_29655);
nand UO_2525 (O_2525,N_29669,N_29651);
nor UO_2526 (O_2526,N_29520,N_29768);
nor UO_2527 (O_2527,N_29745,N_29799);
nor UO_2528 (O_2528,N_29577,N_29525);
and UO_2529 (O_2529,N_29540,N_29787);
and UO_2530 (O_2530,N_29847,N_29954);
or UO_2531 (O_2531,N_29843,N_29919);
nand UO_2532 (O_2532,N_29922,N_29985);
xor UO_2533 (O_2533,N_29744,N_29655);
or UO_2534 (O_2534,N_29696,N_29772);
or UO_2535 (O_2535,N_29669,N_29714);
and UO_2536 (O_2536,N_29933,N_29756);
nand UO_2537 (O_2537,N_29726,N_29556);
nand UO_2538 (O_2538,N_29735,N_29710);
and UO_2539 (O_2539,N_29949,N_29620);
nor UO_2540 (O_2540,N_29888,N_29791);
xnor UO_2541 (O_2541,N_29649,N_29631);
nor UO_2542 (O_2542,N_29513,N_29972);
and UO_2543 (O_2543,N_29544,N_29721);
and UO_2544 (O_2544,N_29948,N_29784);
and UO_2545 (O_2545,N_29669,N_29570);
or UO_2546 (O_2546,N_29744,N_29847);
and UO_2547 (O_2547,N_29662,N_29557);
nor UO_2548 (O_2548,N_29999,N_29651);
xor UO_2549 (O_2549,N_29924,N_29618);
and UO_2550 (O_2550,N_29625,N_29902);
nor UO_2551 (O_2551,N_29635,N_29687);
nand UO_2552 (O_2552,N_29546,N_29600);
and UO_2553 (O_2553,N_29514,N_29570);
nand UO_2554 (O_2554,N_29866,N_29699);
and UO_2555 (O_2555,N_29614,N_29518);
nor UO_2556 (O_2556,N_29921,N_29721);
nand UO_2557 (O_2557,N_29779,N_29714);
or UO_2558 (O_2558,N_29692,N_29671);
nand UO_2559 (O_2559,N_29962,N_29940);
or UO_2560 (O_2560,N_29588,N_29767);
and UO_2561 (O_2561,N_29941,N_29885);
nor UO_2562 (O_2562,N_29803,N_29950);
or UO_2563 (O_2563,N_29865,N_29570);
or UO_2564 (O_2564,N_29954,N_29508);
and UO_2565 (O_2565,N_29672,N_29714);
nor UO_2566 (O_2566,N_29895,N_29558);
xnor UO_2567 (O_2567,N_29954,N_29511);
and UO_2568 (O_2568,N_29767,N_29879);
nand UO_2569 (O_2569,N_29580,N_29847);
nand UO_2570 (O_2570,N_29963,N_29735);
and UO_2571 (O_2571,N_29668,N_29585);
nand UO_2572 (O_2572,N_29613,N_29905);
and UO_2573 (O_2573,N_29866,N_29911);
nor UO_2574 (O_2574,N_29666,N_29686);
nor UO_2575 (O_2575,N_29903,N_29718);
nand UO_2576 (O_2576,N_29794,N_29841);
or UO_2577 (O_2577,N_29913,N_29989);
or UO_2578 (O_2578,N_29554,N_29829);
xor UO_2579 (O_2579,N_29818,N_29732);
and UO_2580 (O_2580,N_29608,N_29941);
nor UO_2581 (O_2581,N_29878,N_29760);
xnor UO_2582 (O_2582,N_29750,N_29633);
xor UO_2583 (O_2583,N_29508,N_29536);
nand UO_2584 (O_2584,N_29817,N_29829);
nor UO_2585 (O_2585,N_29508,N_29816);
and UO_2586 (O_2586,N_29610,N_29620);
or UO_2587 (O_2587,N_29584,N_29885);
nand UO_2588 (O_2588,N_29899,N_29777);
and UO_2589 (O_2589,N_29590,N_29589);
nand UO_2590 (O_2590,N_29664,N_29936);
xor UO_2591 (O_2591,N_29660,N_29866);
nor UO_2592 (O_2592,N_29729,N_29558);
or UO_2593 (O_2593,N_29721,N_29550);
nor UO_2594 (O_2594,N_29645,N_29511);
and UO_2595 (O_2595,N_29978,N_29598);
nand UO_2596 (O_2596,N_29734,N_29605);
or UO_2597 (O_2597,N_29896,N_29583);
and UO_2598 (O_2598,N_29506,N_29979);
or UO_2599 (O_2599,N_29927,N_29668);
nand UO_2600 (O_2600,N_29628,N_29730);
and UO_2601 (O_2601,N_29615,N_29984);
nand UO_2602 (O_2602,N_29964,N_29793);
and UO_2603 (O_2603,N_29693,N_29584);
or UO_2604 (O_2604,N_29593,N_29821);
xnor UO_2605 (O_2605,N_29568,N_29593);
xnor UO_2606 (O_2606,N_29615,N_29808);
nand UO_2607 (O_2607,N_29621,N_29735);
or UO_2608 (O_2608,N_29947,N_29726);
and UO_2609 (O_2609,N_29581,N_29677);
nand UO_2610 (O_2610,N_29511,N_29700);
or UO_2611 (O_2611,N_29592,N_29992);
and UO_2612 (O_2612,N_29810,N_29714);
and UO_2613 (O_2613,N_29740,N_29972);
nand UO_2614 (O_2614,N_29588,N_29512);
and UO_2615 (O_2615,N_29717,N_29507);
nor UO_2616 (O_2616,N_29766,N_29548);
or UO_2617 (O_2617,N_29727,N_29837);
nor UO_2618 (O_2618,N_29503,N_29506);
nand UO_2619 (O_2619,N_29803,N_29761);
or UO_2620 (O_2620,N_29655,N_29936);
nand UO_2621 (O_2621,N_29687,N_29554);
xor UO_2622 (O_2622,N_29917,N_29560);
or UO_2623 (O_2623,N_29555,N_29868);
xor UO_2624 (O_2624,N_29698,N_29616);
nor UO_2625 (O_2625,N_29583,N_29681);
xor UO_2626 (O_2626,N_29688,N_29707);
nor UO_2627 (O_2627,N_29766,N_29946);
nand UO_2628 (O_2628,N_29760,N_29693);
nor UO_2629 (O_2629,N_29532,N_29502);
nor UO_2630 (O_2630,N_29600,N_29966);
and UO_2631 (O_2631,N_29503,N_29721);
nor UO_2632 (O_2632,N_29650,N_29619);
nor UO_2633 (O_2633,N_29916,N_29824);
nand UO_2634 (O_2634,N_29665,N_29830);
and UO_2635 (O_2635,N_29750,N_29652);
or UO_2636 (O_2636,N_29604,N_29528);
or UO_2637 (O_2637,N_29591,N_29933);
nor UO_2638 (O_2638,N_29512,N_29815);
and UO_2639 (O_2639,N_29891,N_29569);
nand UO_2640 (O_2640,N_29533,N_29608);
xnor UO_2641 (O_2641,N_29735,N_29818);
xnor UO_2642 (O_2642,N_29700,N_29721);
nand UO_2643 (O_2643,N_29936,N_29541);
or UO_2644 (O_2644,N_29684,N_29579);
xnor UO_2645 (O_2645,N_29654,N_29915);
nor UO_2646 (O_2646,N_29957,N_29723);
and UO_2647 (O_2647,N_29874,N_29914);
nor UO_2648 (O_2648,N_29929,N_29646);
and UO_2649 (O_2649,N_29658,N_29862);
xnor UO_2650 (O_2650,N_29956,N_29556);
or UO_2651 (O_2651,N_29952,N_29861);
xnor UO_2652 (O_2652,N_29599,N_29953);
nand UO_2653 (O_2653,N_29725,N_29595);
nand UO_2654 (O_2654,N_29965,N_29891);
nor UO_2655 (O_2655,N_29947,N_29861);
nand UO_2656 (O_2656,N_29542,N_29558);
and UO_2657 (O_2657,N_29981,N_29533);
or UO_2658 (O_2658,N_29928,N_29805);
xor UO_2659 (O_2659,N_29743,N_29734);
nor UO_2660 (O_2660,N_29642,N_29817);
and UO_2661 (O_2661,N_29500,N_29846);
and UO_2662 (O_2662,N_29717,N_29872);
and UO_2663 (O_2663,N_29838,N_29939);
nand UO_2664 (O_2664,N_29781,N_29564);
and UO_2665 (O_2665,N_29625,N_29980);
xnor UO_2666 (O_2666,N_29937,N_29717);
nor UO_2667 (O_2667,N_29705,N_29798);
nand UO_2668 (O_2668,N_29879,N_29507);
nor UO_2669 (O_2669,N_29843,N_29854);
nor UO_2670 (O_2670,N_29773,N_29861);
or UO_2671 (O_2671,N_29993,N_29938);
or UO_2672 (O_2672,N_29705,N_29589);
or UO_2673 (O_2673,N_29819,N_29849);
nand UO_2674 (O_2674,N_29622,N_29693);
and UO_2675 (O_2675,N_29650,N_29795);
xor UO_2676 (O_2676,N_29833,N_29720);
or UO_2677 (O_2677,N_29771,N_29566);
xor UO_2678 (O_2678,N_29567,N_29962);
xnor UO_2679 (O_2679,N_29688,N_29522);
nor UO_2680 (O_2680,N_29827,N_29716);
and UO_2681 (O_2681,N_29763,N_29716);
and UO_2682 (O_2682,N_29833,N_29723);
nor UO_2683 (O_2683,N_29867,N_29925);
and UO_2684 (O_2684,N_29552,N_29640);
nor UO_2685 (O_2685,N_29838,N_29778);
or UO_2686 (O_2686,N_29947,N_29867);
and UO_2687 (O_2687,N_29774,N_29945);
xor UO_2688 (O_2688,N_29827,N_29621);
nor UO_2689 (O_2689,N_29656,N_29588);
nand UO_2690 (O_2690,N_29597,N_29573);
nand UO_2691 (O_2691,N_29943,N_29829);
xnor UO_2692 (O_2692,N_29655,N_29852);
xor UO_2693 (O_2693,N_29671,N_29705);
nor UO_2694 (O_2694,N_29692,N_29821);
and UO_2695 (O_2695,N_29781,N_29933);
nand UO_2696 (O_2696,N_29511,N_29939);
or UO_2697 (O_2697,N_29605,N_29853);
nor UO_2698 (O_2698,N_29532,N_29829);
xnor UO_2699 (O_2699,N_29960,N_29950);
and UO_2700 (O_2700,N_29966,N_29911);
and UO_2701 (O_2701,N_29668,N_29675);
nor UO_2702 (O_2702,N_29721,N_29959);
xnor UO_2703 (O_2703,N_29940,N_29729);
nor UO_2704 (O_2704,N_29554,N_29608);
nor UO_2705 (O_2705,N_29907,N_29610);
xnor UO_2706 (O_2706,N_29506,N_29848);
or UO_2707 (O_2707,N_29600,N_29800);
nor UO_2708 (O_2708,N_29994,N_29523);
nand UO_2709 (O_2709,N_29577,N_29583);
and UO_2710 (O_2710,N_29905,N_29783);
or UO_2711 (O_2711,N_29590,N_29687);
nor UO_2712 (O_2712,N_29884,N_29874);
nor UO_2713 (O_2713,N_29702,N_29731);
xor UO_2714 (O_2714,N_29576,N_29762);
and UO_2715 (O_2715,N_29776,N_29736);
xor UO_2716 (O_2716,N_29918,N_29787);
nor UO_2717 (O_2717,N_29768,N_29750);
nor UO_2718 (O_2718,N_29913,N_29670);
xnor UO_2719 (O_2719,N_29577,N_29815);
nor UO_2720 (O_2720,N_29731,N_29538);
nor UO_2721 (O_2721,N_29735,N_29980);
or UO_2722 (O_2722,N_29740,N_29791);
and UO_2723 (O_2723,N_29547,N_29734);
and UO_2724 (O_2724,N_29882,N_29856);
or UO_2725 (O_2725,N_29637,N_29581);
nor UO_2726 (O_2726,N_29801,N_29570);
xor UO_2727 (O_2727,N_29570,N_29737);
or UO_2728 (O_2728,N_29754,N_29658);
nand UO_2729 (O_2729,N_29754,N_29510);
nand UO_2730 (O_2730,N_29799,N_29539);
nor UO_2731 (O_2731,N_29763,N_29989);
or UO_2732 (O_2732,N_29613,N_29965);
or UO_2733 (O_2733,N_29560,N_29936);
xor UO_2734 (O_2734,N_29911,N_29606);
xnor UO_2735 (O_2735,N_29639,N_29822);
nor UO_2736 (O_2736,N_29633,N_29940);
nor UO_2737 (O_2737,N_29754,N_29732);
xor UO_2738 (O_2738,N_29547,N_29649);
nor UO_2739 (O_2739,N_29912,N_29606);
or UO_2740 (O_2740,N_29562,N_29787);
and UO_2741 (O_2741,N_29524,N_29850);
nor UO_2742 (O_2742,N_29521,N_29516);
and UO_2743 (O_2743,N_29866,N_29874);
or UO_2744 (O_2744,N_29505,N_29897);
nor UO_2745 (O_2745,N_29869,N_29545);
nand UO_2746 (O_2746,N_29649,N_29898);
or UO_2747 (O_2747,N_29520,N_29683);
or UO_2748 (O_2748,N_29675,N_29968);
xor UO_2749 (O_2749,N_29940,N_29548);
nor UO_2750 (O_2750,N_29527,N_29663);
or UO_2751 (O_2751,N_29990,N_29995);
xor UO_2752 (O_2752,N_29931,N_29552);
nor UO_2753 (O_2753,N_29670,N_29865);
and UO_2754 (O_2754,N_29784,N_29758);
xnor UO_2755 (O_2755,N_29816,N_29543);
nor UO_2756 (O_2756,N_29765,N_29870);
xnor UO_2757 (O_2757,N_29674,N_29684);
and UO_2758 (O_2758,N_29605,N_29988);
nor UO_2759 (O_2759,N_29729,N_29820);
nand UO_2760 (O_2760,N_29661,N_29941);
nand UO_2761 (O_2761,N_29888,N_29884);
xor UO_2762 (O_2762,N_29966,N_29560);
nand UO_2763 (O_2763,N_29740,N_29739);
nor UO_2764 (O_2764,N_29686,N_29687);
or UO_2765 (O_2765,N_29992,N_29844);
nor UO_2766 (O_2766,N_29912,N_29816);
xnor UO_2767 (O_2767,N_29535,N_29786);
and UO_2768 (O_2768,N_29537,N_29960);
and UO_2769 (O_2769,N_29969,N_29828);
nand UO_2770 (O_2770,N_29652,N_29505);
or UO_2771 (O_2771,N_29998,N_29589);
nor UO_2772 (O_2772,N_29659,N_29788);
nor UO_2773 (O_2773,N_29699,N_29537);
or UO_2774 (O_2774,N_29568,N_29668);
or UO_2775 (O_2775,N_29970,N_29721);
and UO_2776 (O_2776,N_29943,N_29834);
nor UO_2777 (O_2777,N_29632,N_29565);
nand UO_2778 (O_2778,N_29926,N_29754);
and UO_2779 (O_2779,N_29802,N_29690);
xnor UO_2780 (O_2780,N_29716,N_29697);
or UO_2781 (O_2781,N_29578,N_29728);
or UO_2782 (O_2782,N_29857,N_29578);
xnor UO_2783 (O_2783,N_29863,N_29908);
and UO_2784 (O_2784,N_29925,N_29507);
xnor UO_2785 (O_2785,N_29577,N_29980);
xnor UO_2786 (O_2786,N_29682,N_29863);
xnor UO_2787 (O_2787,N_29712,N_29785);
or UO_2788 (O_2788,N_29611,N_29543);
and UO_2789 (O_2789,N_29655,N_29934);
nand UO_2790 (O_2790,N_29642,N_29677);
and UO_2791 (O_2791,N_29509,N_29672);
nor UO_2792 (O_2792,N_29701,N_29697);
nand UO_2793 (O_2793,N_29787,N_29640);
xnor UO_2794 (O_2794,N_29885,N_29750);
nor UO_2795 (O_2795,N_29664,N_29981);
and UO_2796 (O_2796,N_29840,N_29731);
nand UO_2797 (O_2797,N_29953,N_29604);
nand UO_2798 (O_2798,N_29613,N_29699);
or UO_2799 (O_2799,N_29672,N_29872);
and UO_2800 (O_2800,N_29667,N_29935);
nor UO_2801 (O_2801,N_29551,N_29980);
and UO_2802 (O_2802,N_29572,N_29502);
xnor UO_2803 (O_2803,N_29829,N_29979);
nor UO_2804 (O_2804,N_29519,N_29773);
and UO_2805 (O_2805,N_29805,N_29505);
xor UO_2806 (O_2806,N_29841,N_29728);
nand UO_2807 (O_2807,N_29691,N_29586);
nor UO_2808 (O_2808,N_29693,N_29865);
xor UO_2809 (O_2809,N_29871,N_29664);
xnor UO_2810 (O_2810,N_29723,N_29604);
and UO_2811 (O_2811,N_29514,N_29876);
and UO_2812 (O_2812,N_29719,N_29716);
xor UO_2813 (O_2813,N_29882,N_29755);
and UO_2814 (O_2814,N_29877,N_29500);
and UO_2815 (O_2815,N_29918,N_29907);
and UO_2816 (O_2816,N_29527,N_29526);
or UO_2817 (O_2817,N_29990,N_29621);
or UO_2818 (O_2818,N_29586,N_29713);
nor UO_2819 (O_2819,N_29677,N_29851);
and UO_2820 (O_2820,N_29555,N_29891);
nand UO_2821 (O_2821,N_29691,N_29613);
or UO_2822 (O_2822,N_29544,N_29825);
nand UO_2823 (O_2823,N_29643,N_29904);
or UO_2824 (O_2824,N_29762,N_29735);
nand UO_2825 (O_2825,N_29590,N_29926);
or UO_2826 (O_2826,N_29808,N_29717);
and UO_2827 (O_2827,N_29986,N_29853);
nor UO_2828 (O_2828,N_29963,N_29616);
nand UO_2829 (O_2829,N_29669,N_29520);
nand UO_2830 (O_2830,N_29713,N_29552);
nor UO_2831 (O_2831,N_29554,N_29971);
or UO_2832 (O_2832,N_29803,N_29532);
and UO_2833 (O_2833,N_29502,N_29953);
and UO_2834 (O_2834,N_29893,N_29884);
and UO_2835 (O_2835,N_29856,N_29776);
or UO_2836 (O_2836,N_29584,N_29614);
nand UO_2837 (O_2837,N_29731,N_29768);
nor UO_2838 (O_2838,N_29802,N_29680);
and UO_2839 (O_2839,N_29863,N_29593);
nand UO_2840 (O_2840,N_29533,N_29613);
xor UO_2841 (O_2841,N_29537,N_29503);
or UO_2842 (O_2842,N_29655,N_29720);
nand UO_2843 (O_2843,N_29796,N_29902);
nor UO_2844 (O_2844,N_29752,N_29578);
xor UO_2845 (O_2845,N_29953,N_29718);
and UO_2846 (O_2846,N_29831,N_29685);
nor UO_2847 (O_2847,N_29730,N_29735);
xor UO_2848 (O_2848,N_29638,N_29958);
xor UO_2849 (O_2849,N_29574,N_29823);
nand UO_2850 (O_2850,N_29813,N_29564);
or UO_2851 (O_2851,N_29632,N_29697);
nor UO_2852 (O_2852,N_29570,N_29870);
nor UO_2853 (O_2853,N_29804,N_29509);
and UO_2854 (O_2854,N_29683,N_29921);
or UO_2855 (O_2855,N_29552,N_29596);
xnor UO_2856 (O_2856,N_29850,N_29900);
xor UO_2857 (O_2857,N_29755,N_29865);
xor UO_2858 (O_2858,N_29965,N_29742);
xor UO_2859 (O_2859,N_29625,N_29759);
or UO_2860 (O_2860,N_29963,N_29898);
nor UO_2861 (O_2861,N_29905,N_29863);
and UO_2862 (O_2862,N_29691,N_29856);
xnor UO_2863 (O_2863,N_29663,N_29997);
and UO_2864 (O_2864,N_29932,N_29525);
and UO_2865 (O_2865,N_29613,N_29844);
or UO_2866 (O_2866,N_29818,N_29810);
or UO_2867 (O_2867,N_29721,N_29916);
xnor UO_2868 (O_2868,N_29806,N_29937);
nand UO_2869 (O_2869,N_29588,N_29971);
and UO_2870 (O_2870,N_29847,N_29824);
and UO_2871 (O_2871,N_29875,N_29918);
nand UO_2872 (O_2872,N_29804,N_29788);
nand UO_2873 (O_2873,N_29783,N_29652);
xor UO_2874 (O_2874,N_29724,N_29511);
nand UO_2875 (O_2875,N_29846,N_29587);
nand UO_2876 (O_2876,N_29885,N_29570);
nand UO_2877 (O_2877,N_29641,N_29544);
nand UO_2878 (O_2878,N_29707,N_29755);
and UO_2879 (O_2879,N_29755,N_29900);
or UO_2880 (O_2880,N_29900,N_29616);
or UO_2881 (O_2881,N_29615,N_29920);
nor UO_2882 (O_2882,N_29822,N_29722);
or UO_2883 (O_2883,N_29821,N_29819);
nor UO_2884 (O_2884,N_29848,N_29959);
xnor UO_2885 (O_2885,N_29805,N_29749);
xnor UO_2886 (O_2886,N_29573,N_29552);
and UO_2887 (O_2887,N_29686,N_29619);
xor UO_2888 (O_2888,N_29860,N_29723);
or UO_2889 (O_2889,N_29540,N_29669);
nand UO_2890 (O_2890,N_29717,N_29523);
or UO_2891 (O_2891,N_29637,N_29972);
nand UO_2892 (O_2892,N_29660,N_29703);
nand UO_2893 (O_2893,N_29690,N_29705);
nor UO_2894 (O_2894,N_29902,N_29823);
or UO_2895 (O_2895,N_29840,N_29631);
nand UO_2896 (O_2896,N_29799,N_29557);
and UO_2897 (O_2897,N_29585,N_29947);
or UO_2898 (O_2898,N_29599,N_29845);
nor UO_2899 (O_2899,N_29662,N_29636);
or UO_2900 (O_2900,N_29736,N_29730);
and UO_2901 (O_2901,N_29783,N_29969);
and UO_2902 (O_2902,N_29662,N_29514);
nand UO_2903 (O_2903,N_29941,N_29851);
xor UO_2904 (O_2904,N_29566,N_29901);
nand UO_2905 (O_2905,N_29857,N_29922);
nor UO_2906 (O_2906,N_29976,N_29904);
xnor UO_2907 (O_2907,N_29729,N_29589);
nand UO_2908 (O_2908,N_29556,N_29742);
xor UO_2909 (O_2909,N_29751,N_29901);
nand UO_2910 (O_2910,N_29982,N_29590);
nand UO_2911 (O_2911,N_29532,N_29901);
xor UO_2912 (O_2912,N_29904,N_29950);
and UO_2913 (O_2913,N_29977,N_29581);
xnor UO_2914 (O_2914,N_29533,N_29995);
xor UO_2915 (O_2915,N_29821,N_29823);
nand UO_2916 (O_2916,N_29831,N_29725);
or UO_2917 (O_2917,N_29508,N_29702);
nor UO_2918 (O_2918,N_29676,N_29822);
and UO_2919 (O_2919,N_29901,N_29930);
xor UO_2920 (O_2920,N_29925,N_29629);
or UO_2921 (O_2921,N_29927,N_29544);
nor UO_2922 (O_2922,N_29509,N_29641);
xor UO_2923 (O_2923,N_29945,N_29846);
or UO_2924 (O_2924,N_29713,N_29990);
and UO_2925 (O_2925,N_29733,N_29617);
and UO_2926 (O_2926,N_29859,N_29965);
or UO_2927 (O_2927,N_29898,N_29679);
nor UO_2928 (O_2928,N_29606,N_29975);
nor UO_2929 (O_2929,N_29508,N_29540);
nand UO_2930 (O_2930,N_29790,N_29563);
nand UO_2931 (O_2931,N_29705,N_29723);
nor UO_2932 (O_2932,N_29645,N_29736);
or UO_2933 (O_2933,N_29827,N_29628);
xor UO_2934 (O_2934,N_29649,N_29558);
nand UO_2935 (O_2935,N_29570,N_29889);
nor UO_2936 (O_2936,N_29830,N_29629);
and UO_2937 (O_2937,N_29939,N_29743);
xor UO_2938 (O_2938,N_29627,N_29541);
nor UO_2939 (O_2939,N_29858,N_29537);
and UO_2940 (O_2940,N_29589,N_29535);
or UO_2941 (O_2941,N_29805,N_29712);
nor UO_2942 (O_2942,N_29775,N_29903);
nor UO_2943 (O_2943,N_29636,N_29587);
and UO_2944 (O_2944,N_29678,N_29591);
nand UO_2945 (O_2945,N_29627,N_29622);
nor UO_2946 (O_2946,N_29578,N_29949);
and UO_2947 (O_2947,N_29706,N_29894);
or UO_2948 (O_2948,N_29613,N_29764);
and UO_2949 (O_2949,N_29544,N_29669);
or UO_2950 (O_2950,N_29641,N_29711);
nand UO_2951 (O_2951,N_29959,N_29597);
nor UO_2952 (O_2952,N_29539,N_29800);
xnor UO_2953 (O_2953,N_29608,N_29830);
nor UO_2954 (O_2954,N_29669,N_29942);
nor UO_2955 (O_2955,N_29806,N_29526);
or UO_2956 (O_2956,N_29853,N_29788);
and UO_2957 (O_2957,N_29576,N_29924);
xnor UO_2958 (O_2958,N_29932,N_29801);
nand UO_2959 (O_2959,N_29842,N_29616);
nor UO_2960 (O_2960,N_29867,N_29780);
xnor UO_2961 (O_2961,N_29679,N_29627);
nand UO_2962 (O_2962,N_29795,N_29601);
xor UO_2963 (O_2963,N_29803,N_29554);
nand UO_2964 (O_2964,N_29631,N_29551);
or UO_2965 (O_2965,N_29734,N_29520);
nor UO_2966 (O_2966,N_29906,N_29691);
nand UO_2967 (O_2967,N_29638,N_29930);
or UO_2968 (O_2968,N_29720,N_29565);
or UO_2969 (O_2969,N_29945,N_29982);
nor UO_2970 (O_2970,N_29782,N_29579);
nor UO_2971 (O_2971,N_29643,N_29933);
or UO_2972 (O_2972,N_29556,N_29655);
or UO_2973 (O_2973,N_29990,N_29627);
xor UO_2974 (O_2974,N_29594,N_29718);
xor UO_2975 (O_2975,N_29663,N_29958);
and UO_2976 (O_2976,N_29801,N_29659);
or UO_2977 (O_2977,N_29888,N_29680);
nand UO_2978 (O_2978,N_29649,N_29982);
nor UO_2979 (O_2979,N_29758,N_29622);
nand UO_2980 (O_2980,N_29531,N_29924);
nor UO_2981 (O_2981,N_29793,N_29515);
or UO_2982 (O_2982,N_29866,N_29585);
xor UO_2983 (O_2983,N_29604,N_29620);
xnor UO_2984 (O_2984,N_29758,N_29790);
nor UO_2985 (O_2985,N_29750,N_29797);
nor UO_2986 (O_2986,N_29672,N_29995);
nor UO_2987 (O_2987,N_29697,N_29944);
and UO_2988 (O_2988,N_29885,N_29855);
nand UO_2989 (O_2989,N_29537,N_29528);
and UO_2990 (O_2990,N_29880,N_29502);
or UO_2991 (O_2991,N_29563,N_29921);
or UO_2992 (O_2992,N_29602,N_29789);
or UO_2993 (O_2993,N_29756,N_29766);
and UO_2994 (O_2994,N_29512,N_29890);
xnor UO_2995 (O_2995,N_29598,N_29821);
xor UO_2996 (O_2996,N_29720,N_29974);
nand UO_2997 (O_2997,N_29890,N_29692);
xnor UO_2998 (O_2998,N_29819,N_29697);
and UO_2999 (O_2999,N_29732,N_29937);
nand UO_3000 (O_3000,N_29562,N_29674);
nor UO_3001 (O_3001,N_29973,N_29693);
nand UO_3002 (O_3002,N_29909,N_29902);
xor UO_3003 (O_3003,N_29768,N_29597);
xor UO_3004 (O_3004,N_29543,N_29997);
nand UO_3005 (O_3005,N_29734,N_29807);
xnor UO_3006 (O_3006,N_29792,N_29673);
or UO_3007 (O_3007,N_29703,N_29963);
and UO_3008 (O_3008,N_29573,N_29654);
xnor UO_3009 (O_3009,N_29565,N_29866);
or UO_3010 (O_3010,N_29720,N_29669);
or UO_3011 (O_3011,N_29836,N_29990);
xnor UO_3012 (O_3012,N_29507,N_29941);
or UO_3013 (O_3013,N_29867,N_29959);
nor UO_3014 (O_3014,N_29574,N_29719);
nand UO_3015 (O_3015,N_29648,N_29622);
nand UO_3016 (O_3016,N_29732,N_29999);
xnor UO_3017 (O_3017,N_29785,N_29903);
xor UO_3018 (O_3018,N_29808,N_29999);
and UO_3019 (O_3019,N_29621,N_29937);
nor UO_3020 (O_3020,N_29503,N_29730);
xor UO_3021 (O_3021,N_29938,N_29729);
nor UO_3022 (O_3022,N_29867,N_29751);
and UO_3023 (O_3023,N_29789,N_29713);
and UO_3024 (O_3024,N_29819,N_29529);
xnor UO_3025 (O_3025,N_29935,N_29864);
and UO_3026 (O_3026,N_29558,N_29584);
or UO_3027 (O_3027,N_29854,N_29502);
or UO_3028 (O_3028,N_29662,N_29525);
xnor UO_3029 (O_3029,N_29864,N_29735);
nor UO_3030 (O_3030,N_29610,N_29829);
nand UO_3031 (O_3031,N_29727,N_29972);
and UO_3032 (O_3032,N_29945,N_29593);
nand UO_3033 (O_3033,N_29878,N_29645);
nand UO_3034 (O_3034,N_29626,N_29791);
nand UO_3035 (O_3035,N_29767,N_29953);
nand UO_3036 (O_3036,N_29892,N_29983);
or UO_3037 (O_3037,N_29714,N_29871);
nor UO_3038 (O_3038,N_29527,N_29533);
nand UO_3039 (O_3039,N_29555,N_29831);
xnor UO_3040 (O_3040,N_29585,N_29908);
or UO_3041 (O_3041,N_29735,N_29668);
nor UO_3042 (O_3042,N_29873,N_29999);
nand UO_3043 (O_3043,N_29924,N_29565);
nor UO_3044 (O_3044,N_29612,N_29974);
or UO_3045 (O_3045,N_29506,N_29686);
nor UO_3046 (O_3046,N_29910,N_29762);
and UO_3047 (O_3047,N_29661,N_29798);
nand UO_3048 (O_3048,N_29976,N_29645);
nor UO_3049 (O_3049,N_29819,N_29705);
and UO_3050 (O_3050,N_29915,N_29732);
and UO_3051 (O_3051,N_29555,N_29687);
and UO_3052 (O_3052,N_29984,N_29999);
nand UO_3053 (O_3053,N_29854,N_29983);
or UO_3054 (O_3054,N_29810,N_29745);
and UO_3055 (O_3055,N_29821,N_29734);
nor UO_3056 (O_3056,N_29916,N_29988);
and UO_3057 (O_3057,N_29898,N_29977);
or UO_3058 (O_3058,N_29677,N_29559);
xnor UO_3059 (O_3059,N_29965,N_29559);
nand UO_3060 (O_3060,N_29740,N_29681);
nor UO_3061 (O_3061,N_29628,N_29868);
xor UO_3062 (O_3062,N_29896,N_29643);
or UO_3063 (O_3063,N_29556,N_29740);
or UO_3064 (O_3064,N_29840,N_29570);
xor UO_3065 (O_3065,N_29967,N_29653);
or UO_3066 (O_3066,N_29616,N_29831);
nand UO_3067 (O_3067,N_29669,N_29927);
and UO_3068 (O_3068,N_29713,N_29955);
nand UO_3069 (O_3069,N_29996,N_29566);
nor UO_3070 (O_3070,N_29550,N_29617);
and UO_3071 (O_3071,N_29918,N_29523);
or UO_3072 (O_3072,N_29879,N_29646);
or UO_3073 (O_3073,N_29587,N_29856);
nand UO_3074 (O_3074,N_29526,N_29915);
and UO_3075 (O_3075,N_29687,N_29689);
or UO_3076 (O_3076,N_29865,N_29849);
and UO_3077 (O_3077,N_29738,N_29778);
nand UO_3078 (O_3078,N_29921,N_29952);
xnor UO_3079 (O_3079,N_29737,N_29724);
xor UO_3080 (O_3080,N_29623,N_29539);
xor UO_3081 (O_3081,N_29562,N_29519);
xnor UO_3082 (O_3082,N_29893,N_29610);
or UO_3083 (O_3083,N_29918,N_29755);
and UO_3084 (O_3084,N_29831,N_29839);
and UO_3085 (O_3085,N_29930,N_29639);
nand UO_3086 (O_3086,N_29611,N_29681);
xor UO_3087 (O_3087,N_29959,N_29769);
or UO_3088 (O_3088,N_29538,N_29511);
nand UO_3089 (O_3089,N_29943,N_29564);
or UO_3090 (O_3090,N_29768,N_29623);
nand UO_3091 (O_3091,N_29761,N_29672);
nor UO_3092 (O_3092,N_29837,N_29687);
and UO_3093 (O_3093,N_29889,N_29733);
nand UO_3094 (O_3094,N_29826,N_29803);
nand UO_3095 (O_3095,N_29970,N_29746);
or UO_3096 (O_3096,N_29610,N_29868);
xor UO_3097 (O_3097,N_29580,N_29986);
or UO_3098 (O_3098,N_29839,N_29790);
and UO_3099 (O_3099,N_29509,N_29803);
nand UO_3100 (O_3100,N_29605,N_29875);
nor UO_3101 (O_3101,N_29795,N_29699);
nand UO_3102 (O_3102,N_29892,N_29681);
nand UO_3103 (O_3103,N_29745,N_29623);
xnor UO_3104 (O_3104,N_29857,N_29671);
nand UO_3105 (O_3105,N_29538,N_29501);
nand UO_3106 (O_3106,N_29867,N_29978);
nor UO_3107 (O_3107,N_29739,N_29816);
nor UO_3108 (O_3108,N_29518,N_29609);
nor UO_3109 (O_3109,N_29809,N_29804);
and UO_3110 (O_3110,N_29712,N_29877);
or UO_3111 (O_3111,N_29859,N_29879);
nor UO_3112 (O_3112,N_29805,N_29600);
or UO_3113 (O_3113,N_29819,N_29870);
nor UO_3114 (O_3114,N_29738,N_29553);
nor UO_3115 (O_3115,N_29600,N_29505);
xnor UO_3116 (O_3116,N_29767,N_29995);
nand UO_3117 (O_3117,N_29916,N_29814);
xnor UO_3118 (O_3118,N_29895,N_29812);
or UO_3119 (O_3119,N_29989,N_29893);
nand UO_3120 (O_3120,N_29750,N_29794);
or UO_3121 (O_3121,N_29822,N_29766);
or UO_3122 (O_3122,N_29593,N_29861);
and UO_3123 (O_3123,N_29964,N_29988);
nor UO_3124 (O_3124,N_29888,N_29692);
nor UO_3125 (O_3125,N_29874,N_29698);
or UO_3126 (O_3126,N_29798,N_29851);
and UO_3127 (O_3127,N_29522,N_29922);
and UO_3128 (O_3128,N_29583,N_29892);
and UO_3129 (O_3129,N_29687,N_29752);
or UO_3130 (O_3130,N_29525,N_29786);
or UO_3131 (O_3131,N_29866,N_29659);
and UO_3132 (O_3132,N_29842,N_29883);
nor UO_3133 (O_3133,N_29911,N_29737);
nor UO_3134 (O_3134,N_29788,N_29667);
xnor UO_3135 (O_3135,N_29679,N_29802);
nor UO_3136 (O_3136,N_29988,N_29939);
xnor UO_3137 (O_3137,N_29595,N_29944);
or UO_3138 (O_3138,N_29550,N_29777);
xor UO_3139 (O_3139,N_29994,N_29554);
or UO_3140 (O_3140,N_29905,N_29851);
and UO_3141 (O_3141,N_29550,N_29701);
or UO_3142 (O_3142,N_29762,N_29658);
and UO_3143 (O_3143,N_29724,N_29588);
xnor UO_3144 (O_3144,N_29926,N_29812);
nor UO_3145 (O_3145,N_29714,N_29725);
nand UO_3146 (O_3146,N_29670,N_29581);
or UO_3147 (O_3147,N_29599,N_29826);
nand UO_3148 (O_3148,N_29613,N_29850);
xnor UO_3149 (O_3149,N_29615,N_29911);
or UO_3150 (O_3150,N_29594,N_29888);
xnor UO_3151 (O_3151,N_29755,N_29500);
or UO_3152 (O_3152,N_29595,N_29677);
xor UO_3153 (O_3153,N_29648,N_29504);
or UO_3154 (O_3154,N_29670,N_29880);
and UO_3155 (O_3155,N_29772,N_29918);
nor UO_3156 (O_3156,N_29903,N_29568);
and UO_3157 (O_3157,N_29890,N_29760);
nand UO_3158 (O_3158,N_29903,N_29534);
and UO_3159 (O_3159,N_29518,N_29992);
xnor UO_3160 (O_3160,N_29855,N_29659);
nand UO_3161 (O_3161,N_29566,N_29524);
nand UO_3162 (O_3162,N_29767,N_29540);
or UO_3163 (O_3163,N_29997,N_29760);
nor UO_3164 (O_3164,N_29892,N_29646);
nand UO_3165 (O_3165,N_29777,N_29763);
nor UO_3166 (O_3166,N_29943,N_29693);
or UO_3167 (O_3167,N_29602,N_29633);
nand UO_3168 (O_3168,N_29790,N_29824);
or UO_3169 (O_3169,N_29538,N_29553);
and UO_3170 (O_3170,N_29595,N_29682);
nor UO_3171 (O_3171,N_29759,N_29767);
nand UO_3172 (O_3172,N_29939,N_29868);
nor UO_3173 (O_3173,N_29708,N_29567);
and UO_3174 (O_3174,N_29997,N_29779);
nand UO_3175 (O_3175,N_29711,N_29970);
and UO_3176 (O_3176,N_29779,N_29527);
xnor UO_3177 (O_3177,N_29608,N_29745);
nor UO_3178 (O_3178,N_29555,N_29728);
or UO_3179 (O_3179,N_29764,N_29839);
nor UO_3180 (O_3180,N_29942,N_29715);
xor UO_3181 (O_3181,N_29728,N_29621);
and UO_3182 (O_3182,N_29927,N_29786);
nor UO_3183 (O_3183,N_29545,N_29731);
nand UO_3184 (O_3184,N_29672,N_29870);
xor UO_3185 (O_3185,N_29949,N_29972);
nor UO_3186 (O_3186,N_29951,N_29791);
or UO_3187 (O_3187,N_29810,N_29696);
nor UO_3188 (O_3188,N_29624,N_29547);
and UO_3189 (O_3189,N_29750,N_29728);
nor UO_3190 (O_3190,N_29687,N_29952);
nand UO_3191 (O_3191,N_29968,N_29916);
and UO_3192 (O_3192,N_29659,N_29531);
nor UO_3193 (O_3193,N_29640,N_29719);
or UO_3194 (O_3194,N_29702,N_29816);
and UO_3195 (O_3195,N_29839,N_29686);
nor UO_3196 (O_3196,N_29937,N_29767);
nor UO_3197 (O_3197,N_29659,N_29824);
nor UO_3198 (O_3198,N_29782,N_29821);
or UO_3199 (O_3199,N_29739,N_29846);
and UO_3200 (O_3200,N_29777,N_29537);
xor UO_3201 (O_3201,N_29720,N_29748);
xor UO_3202 (O_3202,N_29739,N_29689);
nand UO_3203 (O_3203,N_29643,N_29627);
nor UO_3204 (O_3204,N_29594,N_29921);
and UO_3205 (O_3205,N_29958,N_29951);
xor UO_3206 (O_3206,N_29587,N_29997);
or UO_3207 (O_3207,N_29880,N_29581);
xor UO_3208 (O_3208,N_29645,N_29885);
or UO_3209 (O_3209,N_29612,N_29827);
nand UO_3210 (O_3210,N_29717,N_29648);
xor UO_3211 (O_3211,N_29930,N_29875);
nor UO_3212 (O_3212,N_29726,N_29789);
and UO_3213 (O_3213,N_29648,N_29883);
or UO_3214 (O_3214,N_29541,N_29986);
nor UO_3215 (O_3215,N_29613,N_29734);
or UO_3216 (O_3216,N_29693,N_29738);
xnor UO_3217 (O_3217,N_29715,N_29592);
nand UO_3218 (O_3218,N_29860,N_29866);
xor UO_3219 (O_3219,N_29892,N_29513);
or UO_3220 (O_3220,N_29982,N_29783);
nor UO_3221 (O_3221,N_29702,N_29569);
and UO_3222 (O_3222,N_29572,N_29747);
xor UO_3223 (O_3223,N_29757,N_29877);
and UO_3224 (O_3224,N_29962,N_29700);
nand UO_3225 (O_3225,N_29616,N_29565);
nor UO_3226 (O_3226,N_29919,N_29855);
xor UO_3227 (O_3227,N_29544,N_29762);
and UO_3228 (O_3228,N_29825,N_29672);
xnor UO_3229 (O_3229,N_29636,N_29664);
nor UO_3230 (O_3230,N_29921,N_29742);
and UO_3231 (O_3231,N_29637,N_29843);
nor UO_3232 (O_3232,N_29589,N_29712);
and UO_3233 (O_3233,N_29819,N_29692);
nor UO_3234 (O_3234,N_29881,N_29878);
nand UO_3235 (O_3235,N_29709,N_29684);
or UO_3236 (O_3236,N_29604,N_29831);
xor UO_3237 (O_3237,N_29515,N_29917);
or UO_3238 (O_3238,N_29748,N_29918);
xor UO_3239 (O_3239,N_29716,N_29790);
xor UO_3240 (O_3240,N_29571,N_29844);
nand UO_3241 (O_3241,N_29759,N_29726);
and UO_3242 (O_3242,N_29594,N_29885);
nand UO_3243 (O_3243,N_29728,N_29688);
and UO_3244 (O_3244,N_29974,N_29995);
nand UO_3245 (O_3245,N_29674,N_29960);
nor UO_3246 (O_3246,N_29590,N_29871);
xnor UO_3247 (O_3247,N_29775,N_29978);
xnor UO_3248 (O_3248,N_29517,N_29575);
nand UO_3249 (O_3249,N_29781,N_29948);
and UO_3250 (O_3250,N_29940,N_29757);
or UO_3251 (O_3251,N_29596,N_29538);
or UO_3252 (O_3252,N_29978,N_29963);
nand UO_3253 (O_3253,N_29989,N_29952);
nand UO_3254 (O_3254,N_29895,N_29556);
and UO_3255 (O_3255,N_29877,N_29672);
and UO_3256 (O_3256,N_29532,N_29501);
or UO_3257 (O_3257,N_29685,N_29934);
nand UO_3258 (O_3258,N_29645,N_29915);
nand UO_3259 (O_3259,N_29730,N_29822);
nor UO_3260 (O_3260,N_29774,N_29850);
nand UO_3261 (O_3261,N_29806,N_29573);
nand UO_3262 (O_3262,N_29936,N_29792);
xor UO_3263 (O_3263,N_29684,N_29549);
nand UO_3264 (O_3264,N_29895,N_29925);
nand UO_3265 (O_3265,N_29763,N_29720);
and UO_3266 (O_3266,N_29619,N_29928);
nand UO_3267 (O_3267,N_29666,N_29652);
xnor UO_3268 (O_3268,N_29977,N_29924);
or UO_3269 (O_3269,N_29631,N_29712);
and UO_3270 (O_3270,N_29543,N_29746);
nand UO_3271 (O_3271,N_29780,N_29580);
nand UO_3272 (O_3272,N_29702,N_29647);
and UO_3273 (O_3273,N_29827,N_29558);
xnor UO_3274 (O_3274,N_29633,N_29510);
nand UO_3275 (O_3275,N_29692,N_29783);
and UO_3276 (O_3276,N_29875,N_29637);
nor UO_3277 (O_3277,N_29812,N_29962);
and UO_3278 (O_3278,N_29864,N_29945);
nor UO_3279 (O_3279,N_29973,N_29759);
or UO_3280 (O_3280,N_29710,N_29584);
xor UO_3281 (O_3281,N_29615,N_29773);
nor UO_3282 (O_3282,N_29529,N_29837);
xor UO_3283 (O_3283,N_29618,N_29580);
and UO_3284 (O_3284,N_29558,N_29704);
and UO_3285 (O_3285,N_29995,N_29644);
or UO_3286 (O_3286,N_29524,N_29589);
and UO_3287 (O_3287,N_29656,N_29780);
nand UO_3288 (O_3288,N_29913,N_29643);
nor UO_3289 (O_3289,N_29978,N_29823);
or UO_3290 (O_3290,N_29663,N_29908);
and UO_3291 (O_3291,N_29803,N_29791);
or UO_3292 (O_3292,N_29780,N_29752);
nor UO_3293 (O_3293,N_29960,N_29928);
xor UO_3294 (O_3294,N_29989,N_29548);
xor UO_3295 (O_3295,N_29964,N_29581);
nor UO_3296 (O_3296,N_29535,N_29977);
xnor UO_3297 (O_3297,N_29599,N_29854);
xor UO_3298 (O_3298,N_29580,N_29782);
nor UO_3299 (O_3299,N_29866,N_29808);
nor UO_3300 (O_3300,N_29767,N_29764);
nor UO_3301 (O_3301,N_29604,N_29727);
or UO_3302 (O_3302,N_29581,N_29917);
or UO_3303 (O_3303,N_29635,N_29778);
xnor UO_3304 (O_3304,N_29921,N_29962);
nand UO_3305 (O_3305,N_29634,N_29615);
or UO_3306 (O_3306,N_29703,N_29781);
nand UO_3307 (O_3307,N_29811,N_29907);
nand UO_3308 (O_3308,N_29981,N_29955);
nand UO_3309 (O_3309,N_29629,N_29670);
xnor UO_3310 (O_3310,N_29720,N_29829);
xnor UO_3311 (O_3311,N_29782,N_29504);
nand UO_3312 (O_3312,N_29606,N_29854);
xnor UO_3313 (O_3313,N_29915,N_29798);
nand UO_3314 (O_3314,N_29811,N_29822);
and UO_3315 (O_3315,N_29500,N_29784);
or UO_3316 (O_3316,N_29529,N_29528);
or UO_3317 (O_3317,N_29861,N_29965);
or UO_3318 (O_3318,N_29959,N_29611);
nor UO_3319 (O_3319,N_29753,N_29856);
xor UO_3320 (O_3320,N_29685,N_29905);
or UO_3321 (O_3321,N_29818,N_29711);
xnor UO_3322 (O_3322,N_29978,N_29781);
nor UO_3323 (O_3323,N_29880,N_29518);
xor UO_3324 (O_3324,N_29710,N_29665);
nand UO_3325 (O_3325,N_29682,N_29956);
nor UO_3326 (O_3326,N_29775,N_29627);
or UO_3327 (O_3327,N_29835,N_29694);
nand UO_3328 (O_3328,N_29829,N_29736);
and UO_3329 (O_3329,N_29861,N_29699);
and UO_3330 (O_3330,N_29547,N_29918);
xor UO_3331 (O_3331,N_29745,N_29616);
or UO_3332 (O_3332,N_29805,N_29516);
xor UO_3333 (O_3333,N_29766,N_29539);
and UO_3334 (O_3334,N_29819,N_29858);
nand UO_3335 (O_3335,N_29511,N_29543);
xor UO_3336 (O_3336,N_29572,N_29622);
and UO_3337 (O_3337,N_29575,N_29910);
nor UO_3338 (O_3338,N_29963,N_29832);
and UO_3339 (O_3339,N_29974,N_29567);
nor UO_3340 (O_3340,N_29715,N_29834);
nor UO_3341 (O_3341,N_29750,N_29528);
xnor UO_3342 (O_3342,N_29605,N_29917);
xnor UO_3343 (O_3343,N_29987,N_29706);
nor UO_3344 (O_3344,N_29888,N_29775);
nor UO_3345 (O_3345,N_29750,N_29520);
and UO_3346 (O_3346,N_29676,N_29912);
and UO_3347 (O_3347,N_29756,N_29738);
or UO_3348 (O_3348,N_29893,N_29659);
xor UO_3349 (O_3349,N_29893,N_29831);
xnor UO_3350 (O_3350,N_29553,N_29980);
xnor UO_3351 (O_3351,N_29579,N_29778);
and UO_3352 (O_3352,N_29985,N_29698);
and UO_3353 (O_3353,N_29631,N_29871);
xnor UO_3354 (O_3354,N_29844,N_29627);
xnor UO_3355 (O_3355,N_29511,N_29814);
nor UO_3356 (O_3356,N_29735,N_29796);
and UO_3357 (O_3357,N_29853,N_29983);
xor UO_3358 (O_3358,N_29684,N_29758);
nor UO_3359 (O_3359,N_29882,N_29919);
xor UO_3360 (O_3360,N_29931,N_29749);
nand UO_3361 (O_3361,N_29585,N_29563);
and UO_3362 (O_3362,N_29970,N_29686);
nor UO_3363 (O_3363,N_29930,N_29726);
xor UO_3364 (O_3364,N_29880,N_29964);
or UO_3365 (O_3365,N_29556,N_29855);
xor UO_3366 (O_3366,N_29924,N_29828);
and UO_3367 (O_3367,N_29544,N_29991);
nand UO_3368 (O_3368,N_29584,N_29817);
or UO_3369 (O_3369,N_29840,N_29716);
and UO_3370 (O_3370,N_29665,N_29854);
nand UO_3371 (O_3371,N_29807,N_29922);
nor UO_3372 (O_3372,N_29809,N_29595);
or UO_3373 (O_3373,N_29809,N_29859);
nor UO_3374 (O_3374,N_29895,N_29526);
nand UO_3375 (O_3375,N_29601,N_29548);
nand UO_3376 (O_3376,N_29880,N_29613);
or UO_3377 (O_3377,N_29639,N_29684);
or UO_3378 (O_3378,N_29867,N_29851);
nor UO_3379 (O_3379,N_29757,N_29661);
xor UO_3380 (O_3380,N_29843,N_29782);
xnor UO_3381 (O_3381,N_29878,N_29833);
nor UO_3382 (O_3382,N_29767,N_29792);
or UO_3383 (O_3383,N_29505,N_29542);
or UO_3384 (O_3384,N_29668,N_29687);
xnor UO_3385 (O_3385,N_29670,N_29998);
nor UO_3386 (O_3386,N_29575,N_29825);
or UO_3387 (O_3387,N_29719,N_29557);
nor UO_3388 (O_3388,N_29670,N_29933);
nand UO_3389 (O_3389,N_29943,N_29619);
nand UO_3390 (O_3390,N_29982,N_29901);
xnor UO_3391 (O_3391,N_29986,N_29760);
nand UO_3392 (O_3392,N_29978,N_29643);
xor UO_3393 (O_3393,N_29665,N_29538);
nor UO_3394 (O_3394,N_29659,N_29609);
or UO_3395 (O_3395,N_29990,N_29514);
nor UO_3396 (O_3396,N_29950,N_29817);
nand UO_3397 (O_3397,N_29584,N_29677);
nor UO_3398 (O_3398,N_29821,N_29937);
nand UO_3399 (O_3399,N_29687,N_29579);
xnor UO_3400 (O_3400,N_29609,N_29790);
or UO_3401 (O_3401,N_29812,N_29653);
nor UO_3402 (O_3402,N_29684,N_29948);
xor UO_3403 (O_3403,N_29834,N_29612);
and UO_3404 (O_3404,N_29691,N_29983);
and UO_3405 (O_3405,N_29887,N_29985);
nor UO_3406 (O_3406,N_29534,N_29739);
nand UO_3407 (O_3407,N_29835,N_29705);
xor UO_3408 (O_3408,N_29563,N_29889);
and UO_3409 (O_3409,N_29600,N_29549);
nand UO_3410 (O_3410,N_29563,N_29797);
nand UO_3411 (O_3411,N_29640,N_29730);
and UO_3412 (O_3412,N_29949,N_29812);
nor UO_3413 (O_3413,N_29947,N_29742);
nand UO_3414 (O_3414,N_29577,N_29714);
nor UO_3415 (O_3415,N_29827,N_29749);
xor UO_3416 (O_3416,N_29768,N_29625);
and UO_3417 (O_3417,N_29747,N_29577);
nand UO_3418 (O_3418,N_29535,N_29759);
or UO_3419 (O_3419,N_29905,N_29915);
nor UO_3420 (O_3420,N_29627,N_29507);
nand UO_3421 (O_3421,N_29893,N_29904);
nand UO_3422 (O_3422,N_29742,N_29693);
nor UO_3423 (O_3423,N_29993,N_29825);
or UO_3424 (O_3424,N_29626,N_29609);
nand UO_3425 (O_3425,N_29650,N_29773);
nand UO_3426 (O_3426,N_29682,N_29540);
xor UO_3427 (O_3427,N_29965,N_29873);
nor UO_3428 (O_3428,N_29564,N_29978);
nor UO_3429 (O_3429,N_29959,N_29624);
xor UO_3430 (O_3430,N_29694,N_29879);
nand UO_3431 (O_3431,N_29944,N_29704);
and UO_3432 (O_3432,N_29742,N_29746);
nand UO_3433 (O_3433,N_29613,N_29882);
nand UO_3434 (O_3434,N_29643,N_29831);
nand UO_3435 (O_3435,N_29558,N_29926);
nand UO_3436 (O_3436,N_29551,N_29607);
and UO_3437 (O_3437,N_29813,N_29952);
or UO_3438 (O_3438,N_29618,N_29747);
xnor UO_3439 (O_3439,N_29801,N_29844);
and UO_3440 (O_3440,N_29671,N_29783);
nor UO_3441 (O_3441,N_29631,N_29901);
or UO_3442 (O_3442,N_29997,N_29780);
nand UO_3443 (O_3443,N_29853,N_29820);
or UO_3444 (O_3444,N_29506,N_29825);
or UO_3445 (O_3445,N_29871,N_29945);
nor UO_3446 (O_3446,N_29636,N_29840);
or UO_3447 (O_3447,N_29526,N_29521);
or UO_3448 (O_3448,N_29824,N_29508);
and UO_3449 (O_3449,N_29503,N_29810);
nand UO_3450 (O_3450,N_29945,N_29618);
or UO_3451 (O_3451,N_29631,N_29767);
and UO_3452 (O_3452,N_29830,N_29512);
or UO_3453 (O_3453,N_29703,N_29589);
or UO_3454 (O_3454,N_29646,N_29663);
and UO_3455 (O_3455,N_29670,N_29598);
xnor UO_3456 (O_3456,N_29701,N_29984);
nand UO_3457 (O_3457,N_29859,N_29974);
nor UO_3458 (O_3458,N_29969,N_29712);
and UO_3459 (O_3459,N_29594,N_29909);
and UO_3460 (O_3460,N_29508,N_29865);
nor UO_3461 (O_3461,N_29784,N_29501);
and UO_3462 (O_3462,N_29567,N_29553);
or UO_3463 (O_3463,N_29998,N_29945);
nor UO_3464 (O_3464,N_29802,N_29615);
or UO_3465 (O_3465,N_29569,N_29807);
nand UO_3466 (O_3466,N_29881,N_29704);
nor UO_3467 (O_3467,N_29568,N_29575);
or UO_3468 (O_3468,N_29706,N_29805);
nor UO_3469 (O_3469,N_29665,N_29760);
and UO_3470 (O_3470,N_29685,N_29942);
nor UO_3471 (O_3471,N_29718,N_29539);
nor UO_3472 (O_3472,N_29558,N_29889);
nand UO_3473 (O_3473,N_29917,N_29874);
xor UO_3474 (O_3474,N_29723,N_29654);
xnor UO_3475 (O_3475,N_29786,N_29563);
or UO_3476 (O_3476,N_29680,N_29627);
xnor UO_3477 (O_3477,N_29637,N_29824);
xor UO_3478 (O_3478,N_29978,N_29797);
and UO_3479 (O_3479,N_29980,N_29794);
nor UO_3480 (O_3480,N_29705,N_29996);
and UO_3481 (O_3481,N_29990,N_29939);
or UO_3482 (O_3482,N_29591,N_29750);
xor UO_3483 (O_3483,N_29696,N_29661);
and UO_3484 (O_3484,N_29744,N_29723);
and UO_3485 (O_3485,N_29782,N_29572);
or UO_3486 (O_3486,N_29870,N_29998);
xnor UO_3487 (O_3487,N_29572,N_29924);
and UO_3488 (O_3488,N_29504,N_29526);
nand UO_3489 (O_3489,N_29652,N_29870);
nor UO_3490 (O_3490,N_29619,N_29609);
nor UO_3491 (O_3491,N_29637,N_29952);
or UO_3492 (O_3492,N_29807,N_29797);
or UO_3493 (O_3493,N_29773,N_29543);
and UO_3494 (O_3494,N_29648,N_29944);
and UO_3495 (O_3495,N_29874,N_29897);
nand UO_3496 (O_3496,N_29967,N_29898);
and UO_3497 (O_3497,N_29895,N_29854);
xnor UO_3498 (O_3498,N_29811,N_29713);
nand UO_3499 (O_3499,N_29571,N_29667);
endmodule