module basic_2000_20000_2500_50_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_96,In_773);
or U1 (N_1,In_1812,In_984);
and U2 (N_2,In_920,In_551);
xor U3 (N_3,In_1443,In_194);
and U4 (N_4,In_1749,In_44);
xnor U5 (N_5,In_614,In_161);
and U6 (N_6,In_1767,In_1714);
nand U7 (N_7,In_1103,In_777);
or U8 (N_8,In_723,In_808);
nor U9 (N_9,In_1913,In_438);
nor U10 (N_10,In_343,In_959);
or U11 (N_11,In_1455,In_380);
and U12 (N_12,In_1817,In_856);
nor U13 (N_13,In_1199,In_1206);
nor U14 (N_14,In_368,In_311);
or U15 (N_15,In_1622,In_1065);
nand U16 (N_16,In_1953,In_539);
or U17 (N_17,In_1368,In_1915);
or U18 (N_18,In_1766,In_210);
or U19 (N_19,In_1142,In_475);
nor U20 (N_20,In_560,In_1225);
nand U21 (N_21,In_819,In_993);
and U22 (N_22,In_576,In_1193);
nand U23 (N_23,In_1783,In_133);
nand U24 (N_24,In_1623,In_1456);
xor U25 (N_25,In_989,In_1008);
nand U26 (N_26,In_1824,In_153);
xnor U27 (N_27,In_1938,In_1706);
or U28 (N_28,In_1727,In_574);
xor U29 (N_29,In_277,In_1656);
nor U30 (N_30,In_1614,In_945);
or U31 (N_31,In_1995,In_1703);
and U32 (N_32,In_1069,In_1360);
nand U33 (N_33,In_591,In_1599);
or U34 (N_34,In_1990,In_1412);
xnor U35 (N_35,In_493,In_1461);
and U36 (N_36,In_215,In_689);
xnor U37 (N_37,In_359,In_981);
nand U38 (N_38,In_809,In_676);
nor U39 (N_39,In_1753,In_712);
xor U40 (N_40,In_1234,In_1722);
nand U41 (N_41,In_80,In_1440);
nand U42 (N_42,In_352,In_845);
nand U43 (N_43,In_1123,In_526);
or U44 (N_44,In_1037,In_1537);
xnor U45 (N_45,In_1354,In_1305);
xnor U46 (N_46,In_1728,In_1802);
xor U47 (N_47,In_188,In_319);
or U48 (N_48,In_1473,In_527);
xnor U49 (N_49,In_1469,In_241);
xor U50 (N_50,In_675,In_1764);
nand U51 (N_51,In_1215,In_668);
and U52 (N_52,In_838,In_916);
nand U53 (N_53,In_1272,In_1536);
nor U54 (N_54,In_59,In_66);
xor U55 (N_55,In_1523,In_944);
nor U56 (N_56,In_738,In_1459);
nor U57 (N_57,In_1933,In_740);
or U58 (N_58,In_203,In_181);
nand U59 (N_59,In_1160,In_63);
or U60 (N_60,In_1422,In_837);
nand U61 (N_61,In_14,In_1058);
or U62 (N_62,In_653,In_1270);
nor U63 (N_63,In_1046,In_165);
xor U64 (N_64,In_1260,In_1229);
xor U65 (N_65,In_100,In_1314);
and U66 (N_66,In_234,In_73);
or U67 (N_67,In_1488,In_1197);
or U68 (N_68,In_1947,In_111);
nor U69 (N_69,In_1319,In_1431);
nor U70 (N_70,In_1268,In_163);
and U71 (N_71,In_851,In_720);
or U72 (N_72,In_197,In_204);
nand U73 (N_73,In_439,In_731);
nand U74 (N_74,In_106,In_980);
nor U75 (N_75,In_403,In_283);
nand U76 (N_76,In_1711,In_1717);
and U77 (N_77,In_324,In_47);
nor U78 (N_78,In_169,In_1654);
and U79 (N_79,In_1541,In_1552);
and U80 (N_80,In_546,In_681);
nor U81 (N_81,In_1345,In_1575);
nor U82 (N_82,In_1060,In_780);
nor U83 (N_83,In_1895,In_1211);
or U84 (N_84,In_971,In_791);
nor U85 (N_85,In_365,In_1719);
nor U86 (N_86,In_1021,In_101);
nor U87 (N_87,In_1985,In_1191);
and U88 (N_88,In_1054,In_485);
or U89 (N_89,In_933,In_1245);
nor U90 (N_90,In_1850,In_1332);
and U91 (N_91,In_545,In_1872);
nand U92 (N_92,In_1988,In_156);
and U93 (N_93,In_1881,In_1587);
xnor U94 (N_94,In_1289,In_119);
or U95 (N_95,In_1873,In_596);
nor U96 (N_96,In_1896,In_1048);
and U97 (N_97,In_1864,In_1438);
xor U98 (N_98,In_470,In_262);
nand U99 (N_99,In_1586,In_1646);
nor U100 (N_100,In_744,In_1484);
xor U101 (N_101,In_224,In_99);
nor U102 (N_102,In_1047,In_1430);
xnor U103 (N_103,In_1176,In_1448);
and U104 (N_104,In_406,In_444);
or U105 (N_105,In_999,In_1464);
nand U106 (N_106,In_1445,In_1326);
nand U107 (N_107,In_673,In_714);
xnor U108 (N_108,In_1704,In_1528);
or U109 (N_109,In_986,In_226);
xor U110 (N_110,In_1814,In_1909);
or U111 (N_111,In_1013,In_214);
and U112 (N_112,In_1477,In_647);
or U113 (N_113,In_1689,In_634);
nor U114 (N_114,In_537,In_310);
xor U115 (N_115,In_1041,In_1874);
xnor U116 (N_116,In_510,In_1554);
xor U117 (N_117,In_503,In_1153);
nor U118 (N_118,In_1118,In_458);
nor U119 (N_119,In_1468,In_1325);
xnor U120 (N_120,In_1967,In_185);
and U121 (N_121,In_568,In_1378);
and U122 (N_122,In_1070,In_886);
xnor U123 (N_123,In_1009,In_1939);
or U124 (N_124,In_1267,In_1243);
or U125 (N_125,In_1594,In_1089);
or U126 (N_126,In_222,In_255);
xor U127 (N_127,In_4,In_405);
and U128 (N_128,In_1501,In_1603);
or U129 (N_129,In_82,In_221);
nand U130 (N_130,In_23,In_1441);
nor U131 (N_131,In_1663,In_33);
or U132 (N_132,In_1961,In_40);
nor U133 (N_133,In_1044,In_937);
or U134 (N_134,In_1017,In_1127);
nor U135 (N_135,In_1334,In_1572);
nand U136 (N_136,In_963,In_321);
nand U137 (N_137,In_1163,In_1258);
and U138 (N_138,In_825,In_20);
nor U139 (N_139,In_563,In_1558);
or U140 (N_140,In_1490,In_567);
nand U141 (N_141,In_90,In_913);
or U142 (N_142,In_788,In_1034);
nand U143 (N_143,In_1213,In_1216);
nor U144 (N_144,In_822,In_132);
xnor U145 (N_145,In_1097,In_1524);
nor U146 (N_146,In_431,In_1989);
xor U147 (N_147,In_620,In_330);
and U148 (N_148,In_954,In_1836);
nand U149 (N_149,In_1450,In_1503);
xor U150 (N_150,In_1716,In_1724);
xnor U151 (N_151,In_915,In_656);
nand U152 (N_152,In_570,In_1534);
nor U153 (N_153,In_1124,In_1715);
or U154 (N_154,In_461,In_1307);
nand U155 (N_155,In_347,In_480);
and U156 (N_156,In_1186,In_1679);
or U157 (N_157,In_985,In_171);
nor U158 (N_158,In_337,In_1994);
or U159 (N_159,In_1694,In_1849);
nor U160 (N_160,In_473,In_1533);
or U161 (N_161,In_768,In_1472);
and U162 (N_162,In_1776,In_870);
or U163 (N_163,In_756,In_521);
xor U164 (N_164,In_1875,In_238);
xnor U165 (N_165,In_1797,In_1929);
or U166 (N_166,In_680,In_1347);
nand U167 (N_167,In_1863,In_1302);
or U168 (N_168,In_27,In_97);
or U169 (N_169,In_734,In_1079);
nor U170 (N_170,In_1684,In_659);
or U171 (N_171,In_1545,In_1948);
or U172 (N_172,In_1734,In_706);
nor U173 (N_173,In_1512,In_960);
and U174 (N_174,In_623,In_1607);
xor U175 (N_175,In_1886,In_1498);
nor U176 (N_176,In_144,In_1943);
and U177 (N_177,In_1815,In_1866);
and U178 (N_178,In_1106,In_422);
nor U179 (N_179,In_412,In_1742);
xnor U180 (N_180,In_605,In_1283);
and U181 (N_181,In_1978,In_74);
or U182 (N_182,In_663,In_1601);
or U183 (N_183,In_1642,In_864);
or U184 (N_184,In_1649,In_1736);
or U185 (N_185,In_15,In_1958);
xnor U186 (N_186,In_1322,In_54);
or U187 (N_187,In_1239,In_1867);
and U188 (N_188,In_1798,In_1219);
or U189 (N_189,In_432,In_417);
nor U190 (N_190,In_1491,In_292);
xnor U191 (N_191,In_1129,In_832);
and U192 (N_192,In_1592,In_435);
nand U193 (N_193,In_278,In_1000);
nand U194 (N_194,In_1936,In_145);
xnor U195 (N_195,In_416,In_492);
or U196 (N_196,In_1265,In_1999);
xor U197 (N_197,In_1262,In_1261);
or U198 (N_198,In_861,In_1497);
or U199 (N_199,In_968,In_1204);
xnor U200 (N_200,In_1128,In_1963);
nand U201 (N_201,In_328,In_1381);
nand U202 (N_202,In_718,In_445);
or U203 (N_203,In_388,In_637);
xor U204 (N_204,In_24,In_1417);
nand U205 (N_205,In_1135,In_1604);
nand U206 (N_206,In_386,In_1022);
xor U207 (N_207,In_442,In_1861);
nor U208 (N_208,In_217,In_1033);
and U209 (N_209,In_50,In_1208);
or U210 (N_210,In_1007,In_424);
or U211 (N_211,In_409,In_1937);
xnor U212 (N_212,In_1500,In_402);
xor U213 (N_213,In_29,In_1284);
and U214 (N_214,In_31,In_1650);
nor U215 (N_215,In_401,In_291);
nor U216 (N_216,In_695,In_1035);
and U217 (N_217,In_1231,In_1910);
nand U218 (N_218,In_522,In_1379);
nand U219 (N_219,In_1226,In_1294);
nand U220 (N_220,In_1580,In_7);
xnor U221 (N_221,In_275,In_309);
and U222 (N_222,In_441,In_8);
or U223 (N_223,In_1494,In_1955);
nand U224 (N_224,In_108,In_253);
xor U225 (N_225,In_1308,In_1709);
and U226 (N_226,In_376,In_1303);
and U227 (N_227,In_396,In_1840);
or U228 (N_228,In_1670,In_1757);
or U229 (N_229,In_1432,In_116);
or U230 (N_230,In_1457,In_1300);
nand U231 (N_231,In_1241,In_176);
or U232 (N_232,In_11,In_557);
or U233 (N_233,In_327,In_455);
nor U234 (N_234,In_237,In_1969);
nor U235 (N_235,In_554,In_407);
and U236 (N_236,In_64,In_1718);
nor U237 (N_237,In_6,In_918);
nand U238 (N_238,In_143,In_1353);
nor U239 (N_239,In_1145,In_60);
xor U240 (N_240,In_1098,In_1419);
nor U241 (N_241,In_1957,In_797);
or U242 (N_242,In_582,In_1610);
xnor U243 (N_243,In_812,In_28);
or U244 (N_244,In_1600,In_682);
and U245 (N_245,In_1737,In_610);
and U246 (N_246,In_55,In_393);
nor U247 (N_247,In_49,In_899);
nor U248 (N_248,In_489,In_426);
xnor U249 (N_249,In_69,In_816);
nand U250 (N_250,In_789,In_1073);
and U251 (N_251,In_1565,In_1371);
nand U252 (N_252,In_1346,In_1359);
and U253 (N_253,In_894,In_182);
xor U254 (N_254,In_1898,In_589);
nand U255 (N_255,In_774,In_361);
or U256 (N_256,In_326,In_79);
nor U257 (N_257,In_664,In_314);
nand U258 (N_258,In_826,In_331);
nor U259 (N_259,In_708,In_1810);
and U260 (N_260,In_1299,In_2);
and U261 (N_261,In_855,In_1885);
or U262 (N_262,In_779,In_906);
xnor U263 (N_263,In_123,In_1608);
xor U264 (N_264,In_1252,In_935);
and U265 (N_265,In_1190,In_824);
and U266 (N_266,In_471,In_518);
nand U267 (N_267,In_1993,In_295);
nor U268 (N_268,In_1185,In_1436);
xnor U269 (N_269,In_1315,In_757);
and U270 (N_270,In_1792,In_921);
nand U271 (N_271,In_1442,In_198);
or U272 (N_272,In_1400,In_1446);
xnor U273 (N_273,In_1838,In_1925);
and U274 (N_274,In_770,In_1621);
nand U275 (N_275,In_1212,In_674);
xor U276 (N_276,In_1667,In_476);
and U277 (N_277,In_1550,In_1004);
and U278 (N_278,In_644,In_1331);
nand U279 (N_279,In_1201,In_120);
or U280 (N_280,In_76,In_93);
nor U281 (N_281,In_1996,In_823);
nand U282 (N_282,In_1149,In_1529);
or U283 (N_283,In_1750,In_1071);
or U284 (N_284,In_948,In_752);
nor U285 (N_285,In_1235,In_932);
nor U286 (N_286,In_763,In_1602);
xnor U287 (N_287,In_754,In_1221);
nor U288 (N_288,In_1923,In_1641);
xnor U289 (N_289,In_244,In_354);
and U290 (N_290,In_394,In_1084);
nand U291 (N_291,In_1083,In_246);
nor U292 (N_292,In_942,In_1248);
nor U293 (N_293,In_1174,In_1854);
nor U294 (N_294,In_715,In_1743);
and U295 (N_295,In_1390,In_566);
xor U296 (N_296,In_1609,In_201);
xor U297 (N_297,In_317,In_1433);
and U298 (N_298,In_1721,In_1944);
xnor U299 (N_299,In_1591,In_1504);
nor U300 (N_300,In_1730,In_1851);
and U301 (N_301,In_827,In_1370);
nand U302 (N_302,In_1829,In_1232);
nor U303 (N_303,In_177,In_1538);
and U304 (N_304,In_423,In_1489);
nand U305 (N_305,In_645,In_626);
xor U306 (N_306,In_949,In_1356);
xor U307 (N_307,In_1522,In_709);
or U308 (N_308,In_1903,In_155);
xnor U309 (N_309,In_1362,In_820);
or U310 (N_310,In_1647,In_440);
and U311 (N_311,In_301,In_287);
nor U312 (N_312,In_71,In_1920);
nor U313 (N_313,In_872,In_549);
nand U314 (N_314,In_1942,In_225);
nand U315 (N_315,In_1198,In_924);
xnor U316 (N_316,In_136,In_1902);
nor U317 (N_317,In_1297,In_1796);
xor U318 (N_318,In_1793,In_1935);
xor U319 (N_319,In_869,In_446);
nor U320 (N_320,In_271,In_1570);
or U321 (N_321,In_686,In_1148);
or U322 (N_322,In_379,In_1639);
and U323 (N_323,In_951,In_158);
nand U324 (N_324,In_1625,In_931);
nor U325 (N_325,In_1482,In_1805);
and U326 (N_326,In_276,In_1751);
or U327 (N_327,In_477,In_964);
xnor U328 (N_328,In_364,In_1077);
nand U329 (N_329,In_1237,In_1962);
nor U330 (N_330,In_342,In_594);
xor U331 (N_331,In_1959,In_509);
nand U332 (N_332,In_1606,In_146);
and U333 (N_333,In_642,In_178);
nor U334 (N_334,In_1223,In_1343);
or U335 (N_335,In_360,In_600);
nand U336 (N_336,In_129,In_1399);
and U337 (N_337,In_1428,In_124);
nand U338 (N_338,In_86,In_632);
and U339 (N_339,In_1723,In_1982);
or U340 (N_340,In_1871,In_1351);
nor U341 (N_341,In_304,In_131);
xnor U342 (N_342,In_604,In_633);
xnor U343 (N_343,In_1568,In_781);
nor U344 (N_344,In_577,In_1027);
or U345 (N_345,In_1099,In_1141);
nor U346 (N_346,In_1402,In_1414);
and U347 (N_347,In_507,In_308);
and U348 (N_348,In_1555,In_420);
and U349 (N_349,In_172,In_1023);
nor U350 (N_350,In_1110,In_1847);
nor U351 (N_351,In_990,In_1107);
and U352 (N_352,In_1429,In_1596);
or U353 (N_353,In_996,In_843);
xnor U354 (N_354,In_1288,In_1540);
nor U355 (N_355,In_1405,In_553);
nand U356 (N_356,In_1760,In_1638);
nand U357 (N_357,In_1870,In_854);
xor U358 (N_358,In_1478,In_707);
nand U359 (N_359,In_1180,In_385);
and U360 (N_360,In_1165,In_1031);
nor U361 (N_361,In_749,In_57);
or U362 (N_362,In_413,In_922);
or U363 (N_363,In_112,In_547);
nor U364 (N_364,In_1499,In_247);
or U365 (N_365,In_1761,In_252);
nor U366 (N_366,In_1408,In_810);
nor U367 (N_367,In_598,In_1401);
and U368 (N_368,In_1777,In_1310);
nor U369 (N_369,In_1756,In_53);
or U370 (N_370,In_655,In_884);
nand U371 (N_371,In_641,In_1597);
nor U372 (N_372,In_332,In_355);
and U373 (N_373,In_481,In_1518);
nor U374 (N_374,In_46,In_375);
nor U375 (N_375,In_1574,In_1111);
nor U376 (N_376,In_573,In_1474);
or U377 (N_377,In_1074,In_885);
xnor U378 (N_378,In_1067,In_1183);
xnor U379 (N_379,In_282,In_256);
or U380 (N_380,In_1264,In_1746);
xnor U381 (N_381,In_85,In_266);
xnor U382 (N_382,In_279,In_1157);
nand U383 (N_383,In_5,In_87);
or U384 (N_384,In_1908,In_575);
xor U385 (N_385,In_929,In_1344);
or U386 (N_386,In_1336,In_335);
or U387 (N_387,In_1094,In_1683);
nand U388 (N_388,In_1513,In_802);
and U389 (N_389,In_1553,In_662);
xor U390 (N_390,In_91,In_588);
or U391 (N_391,In_251,In_1626);
and U392 (N_392,In_333,In_1105);
or U393 (N_393,In_366,In_1122);
xor U394 (N_394,In_806,In_535);
nor U395 (N_395,In_1517,In_1678);
or U396 (N_396,In_1062,In_1480);
nor U397 (N_397,In_508,In_722);
and U398 (N_398,In_427,In_1636);
xor U399 (N_399,In_1551,In_1154);
or U400 (N_400,N_292,In_1010);
and U401 (N_401,In_687,In_1876);
nand U402 (N_402,In_1209,In_1133);
nand U403 (N_403,In_149,In_164);
and U404 (N_404,N_259,In_743);
or U405 (N_405,In_367,In_1335);
xor U406 (N_406,In_698,In_1170);
and U407 (N_407,In_286,N_372);
xor U408 (N_408,In_1196,In_1583);
nand U409 (N_409,In_260,In_1279);
nand U410 (N_410,In_1341,In_351);
nand U411 (N_411,In_336,In_1960);
xor U412 (N_412,In_1271,N_71);
and U413 (N_413,In_1577,In_1858);
or U414 (N_414,N_7,In_1389);
and U415 (N_415,In_459,In_18);
nor U416 (N_416,N_377,N_366);
nand U417 (N_417,In_1807,In_199);
nand U418 (N_418,In_1470,N_23);
or U419 (N_419,In_1693,N_315);
nor U420 (N_420,N_176,In_519);
nand U421 (N_421,In_72,In_1934);
or U422 (N_422,In_1406,In_1624);
nand U423 (N_423,In_1690,In_1945);
nor U424 (N_424,In_1664,In_150);
xor U425 (N_425,In_506,In_1924);
or U426 (N_426,In_771,In_1671);
nand U427 (N_427,In_273,In_1894);
nor U428 (N_428,In_41,In_939);
xor U429 (N_429,In_1806,In_1560);
nand U430 (N_430,In_688,In_486);
and U431 (N_431,In_142,N_110);
xnor U432 (N_432,In_995,N_278);
or U433 (N_433,In_1525,In_390);
and U434 (N_434,N_209,N_145);
nor U435 (N_435,N_165,N_252);
xor U436 (N_436,N_150,In_1296);
nor U437 (N_437,In_305,In_1901);
or U438 (N_438,N_310,In_1788);
and U439 (N_439,In_1434,In_733);
and U440 (N_440,In_910,N_194);
and U441 (N_441,In_631,N_362);
and U442 (N_442,In_1747,In_988);
xnor U443 (N_443,N_63,In_1868);
or U444 (N_444,In_1927,In_382);
nor U445 (N_445,In_115,In_905);
nand U446 (N_446,In_776,In_807);
nor U447 (N_447,In_958,In_1246);
xnor U448 (N_448,In_672,In_1882);
and U449 (N_449,In_801,In_1045);
nor U450 (N_450,In_1712,In_1147);
nand U451 (N_451,In_257,N_198);
xnor U452 (N_452,N_171,In_428);
and U453 (N_453,In_1210,In_817);
xor U454 (N_454,In_829,In_755);
xnor U455 (N_455,In_624,In_1029);
nor U456 (N_456,In_448,In_1161);
nor U457 (N_457,N_149,In_1979);
or U458 (N_458,In_315,In_1877);
or U459 (N_459,In_127,In_490);
and U460 (N_460,N_395,In_1404);
xnor U461 (N_461,In_1765,In_1324);
nand U462 (N_462,In_1818,N_268);
nor U463 (N_463,In_358,In_1295);
and U464 (N_464,In_88,In_1804);
nand U465 (N_465,In_1543,In_1784);
xnor U466 (N_466,In_1926,In_1505);
and U467 (N_467,In_1358,In_881);
xor U468 (N_468,In_1508,In_1130);
xor U469 (N_469,In_469,In_289);
nand U470 (N_470,In_1892,N_258);
nor U471 (N_471,In_1635,In_205);
nand U472 (N_472,In_1830,N_294);
nand U473 (N_473,In_1841,N_137);
nor U474 (N_474,In_494,In_1782);
or U475 (N_475,N_375,In_792);
nand U476 (N_476,In_593,In_1502);
and U477 (N_477,In_103,In_1862);
nor U478 (N_478,N_173,In_1274);
or U479 (N_479,In_193,In_1420);
xor U480 (N_480,N_73,In_65);
or U481 (N_481,In_540,N_223);
or U482 (N_482,In_1666,In_1855);
xnor U483 (N_483,In_258,N_179);
or U484 (N_484,In_622,In_34);
or U485 (N_485,In_717,In_70);
and U486 (N_486,N_161,In_638);
and U487 (N_487,In_1391,In_901);
nor U488 (N_488,In_1152,In_943);
and U489 (N_489,In_1171,In_1159);
or U490 (N_490,N_323,In_498);
and U491 (N_491,In_798,In_1768);
and U492 (N_492,In_186,In_1321);
or U493 (N_493,N_199,N_111);
xnor U494 (N_494,In_1453,In_1922);
and U495 (N_495,In_19,In_1844);
xor U496 (N_496,In_1364,In_1072);
xnor U497 (N_497,In_579,In_1816);
or U498 (N_498,In_846,In_1019);
or U499 (N_499,N_228,In_767);
or U500 (N_500,N_351,N_300);
nor U501 (N_501,In_1547,In_660);
and U502 (N_502,In_1476,In_1964);
and U503 (N_503,In_1424,In_1257);
or U504 (N_504,In_1549,In_1195);
and U505 (N_505,N_144,In_1318);
and U506 (N_506,In_1151,In_290);
xor U507 (N_507,In_313,N_112);
xor U508 (N_508,N_273,In_1674);
nor U509 (N_509,In_147,In_130);
nor U510 (N_510,In_1631,In_1794);
xor U511 (N_511,In_43,In_857);
and U512 (N_512,In_318,In_840);
nor U513 (N_513,In_138,In_1306);
xor U514 (N_514,In_1511,N_162);
xnor U515 (N_515,In_216,In_1410);
nor U516 (N_516,In_1179,In_491);
nand U517 (N_517,N_70,In_1355);
xor U518 (N_518,N_382,N_324);
xnor U519 (N_519,In_395,In_160);
xor U520 (N_520,N_134,In_994);
nor U521 (N_521,In_764,In_772);
xor U522 (N_522,In_976,In_1984);
nor U523 (N_523,In_1061,In_1976);
nor U524 (N_524,N_299,In_1705);
nand U525 (N_525,In_1630,In_1397);
and U526 (N_526,In_1931,In_880);
nand U527 (N_527,In_1648,In_472);
and U528 (N_528,N_232,In_1175);
and U529 (N_529,In_220,In_209);
nand U530 (N_530,In_1042,N_373);
nand U531 (N_531,N_135,In_1755);
nand U532 (N_532,In_616,In_152);
or U533 (N_533,In_3,N_379);
and U534 (N_534,In_515,In_1563);
nor U535 (N_535,N_226,In_323);
nor U536 (N_536,N_383,In_1643);
xor U537 (N_537,In_1891,In_1119);
and U538 (N_538,In_1842,N_82);
and U539 (N_539,In_1427,In_1658);
xor U540 (N_540,In_800,N_260);
and U541 (N_541,N_50,In_955);
and U542 (N_542,N_66,In_1465);
xnor U543 (N_543,In_552,In_1754);
nand U544 (N_544,N_237,N_92);
and U545 (N_545,N_381,In_1506);
nor U546 (N_546,In_272,In_735);
or U547 (N_547,In_934,In_1822);
and U548 (N_548,In_926,N_35);
and U549 (N_549,In_179,N_106);
xnor U550 (N_550,N_116,In_303);
nand U551 (N_551,In_1825,In_587);
xnor U552 (N_552,In_1169,In_229);
nor U553 (N_553,In_418,In_1291);
nor U554 (N_554,In_1620,In_1696);
and U555 (N_555,In_1282,In_81);
and U556 (N_556,N_319,N_276);
and U557 (N_557,In_578,In_543);
or U558 (N_558,N_157,In_874);
nor U559 (N_559,In_464,N_271);
nand U560 (N_560,In_833,In_1143);
and U561 (N_561,In_1230,In_77);
nand U562 (N_562,In_1038,N_96);
or U563 (N_563,In_1556,N_141);
and U564 (N_564,In_1222,In_1809);
nand U565 (N_565,N_166,In_383);
and U566 (N_566,In_848,N_20);
nand U567 (N_567,N_288,N_220);
nand U568 (N_568,In_1328,N_341);
nand U569 (N_569,In_1114,In_1348);
and U570 (N_570,In_1286,In_1189);
or U571 (N_571,In_1251,In_1653);
and U572 (N_572,N_224,In_860);
or U573 (N_573,In_1585,In_762);
or U574 (N_574,In_790,In_1376);
nand U575 (N_575,N_396,In_1372);
nor U576 (N_576,N_127,In_1155);
xor U577 (N_577,In_297,N_3);
and U578 (N_578,In_148,N_87);
nand U579 (N_579,In_648,N_67);
or U580 (N_580,In_1731,In_759);
or U581 (N_581,In_1691,In_1116);
xnor U582 (N_582,In_316,In_684);
nand U583 (N_583,In_1373,In_1845);
and U584 (N_584,In_1645,N_321);
xor U585 (N_585,In_862,In_9);
nor U586 (N_586,In_189,In_92);
nor U587 (N_587,N_143,In_670);
nor U588 (N_588,In_1131,N_120);
nand U589 (N_589,In_1573,N_74);
or U590 (N_590,In_1380,In_1005);
xor U591 (N_591,In_1285,In_636);
nor U592 (N_592,In_329,In_269);
or U593 (N_593,In_1396,In_357);
xor U594 (N_594,In_168,N_213);
nand U595 (N_595,In_1733,N_10);
nor U596 (N_596,In_739,In_61);
nor U597 (N_597,In_555,In_398);
xnor U598 (N_598,In_1584,In_821);
nand U599 (N_599,In_202,In_1790);
nand U600 (N_600,N_225,In_583);
and U601 (N_601,In_1971,In_962);
nor U602 (N_602,In_1839,N_76);
and U603 (N_603,In_363,In_1542);
or U604 (N_604,In_1848,N_79);
and U605 (N_605,In_325,In_1014);
nand U606 (N_606,In_1972,In_1177);
xnor U607 (N_607,In_1120,In_803);
or U608 (N_608,In_903,In_1853);
or U609 (N_609,In_621,In_454);
or U610 (N_610,In_952,N_138);
or U611 (N_611,N_325,In_1637);
nand U612 (N_612,N_371,In_879);
or U613 (N_613,N_42,In_1087);
or U614 (N_614,In_1852,In_261);
xor U615 (N_615,In_499,In_462);
nand U616 (N_616,In_1278,In_1057);
nand U617 (N_617,N_307,N_397);
and U618 (N_618,N_392,In_411);
or U619 (N_619,N_245,In_1333);
or U620 (N_620,In_1827,In_369);
nand U621 (N_621,In_374,In_1582);
and U622 (N_622,N_31,In_1415);
xnor U623 (N_623,In_895,In_1800);
xor U624 (N_624,In_190,N_230);
nand U625 (N_625,In_1056,In_128);
nor U626 (N_626,In_669,N_277);
nand U627 (N_627,In_930,In_1987);
nor U628 (N_628,In_1832,In_1578);
nor U629 (N_629,In_1786,In_102);
and U630 (N_630,In_1247,In_1374);
nor U631 (N_631,In_1998,N_86);
nand U632 (N_632,In_737,In_1095);
and U633 (N_633,N_88,In_1275);
and U634 (N_634,In_883,In_1672);
xnor U635 (N_635,In_362,N_304);
nand U636 (N_636,In_1566,In_1188);
xnor U637 (N_637,In_1144,N_27);
and U638 (N_638,In_599,N_202);
xnor U639 (N_639,In_430,In_978);
and U640 (N_640,In_852,In_1616);
nor U641 (N_641,In_1820,In_908);
or U642 (N_642,In_1659,In_1527);
or U643 (N_643,In_983,In_818);
and U644 (N_644,N_151,In_1617);
and U645 (N_645,N_37,In_1644);
nor U646 (N_646,In_1521,In_338);
nand U647 (N_647,In_564,N_78);
or U648 (N_648,In_1053,In_1949);
xor U649 (N_649,In_612,In_1605);
or U650 (N_650,In_799,In_736);
nand U651 (N_651,In_1228,In_1425);
nor U652 (N_652,In_1100,In_371);
nand U653 (N_653,In_353,In_1865);
and U654 (N_654,In_419,In_666);
or U655 (N_655,N_338,N_337);
xnor U656 (N_656,In_1317,In_425);
nor U657 (N_657,In_1661,N_72);
nand U658 (N_658,N_285,N_38);
xor U659 (N_659,In_151,In_1117);
and U660 (N_660,In_141,N_242);
or U661 (N_661,In_1011,N_255);
nand U662 (N_662,N_125,N_249);
nand U663 (N_663,In_1769,In_769);
or U664 (N_664,N_222,N_196);
nand U665 (N_665,In_1090,In_565);
and U666 (N_666,In_1173,In_1249);
xor U667 (N_667,In_12,N_227);
and U668 (N_668,In_732,In_447);
xnor U669 (N_669,N_130,N_142);
xor U670 (N_670,In_842,In_307);
or U671 (N_671,In_48,N_295);
or U672 (N_672,N_190,In_1259);
nand U673 (N_673,N_197,N_182);
nand U674 (N_674,In_595,In_265);
nor U675 (N_675,In_1946,N_283);
nor U676 (N_676,In_1860,N_336);
and U677 (N_677,In_1564,In_306);
and U678 (N_678,In_1150,N_286);
or U679 (N_679,N_4,In_1991);
nor U680 (N_680,In_581,In_1435);
xor U681 (N_681,In_1956,In_83);
xnor U682 (N_682,In_630,In_1466);
nand U683 (N_683,In_1514,N_298);
nor U684 (N_684,In_200,N_129);
xor U685 (N_685,N_104,In_654);
nand U686 (N_686,In_909,N_164);
nand U687 (N_687,In_1657,In_987);
xor U688 (N_688,In_339,In_1611);
nand U689 (N_689,In_1387,In_961);
xnor U690 (N_690,In_243,N_345);
xnor U691 (N_691,N_342,In_1739);
nand U692 (N_692,In_538,N_49);
or U693 (N_693,In_890,In_523);
nor U694 (N_694,N_133,In_1952);
nand U695 (N_695,In_746,In_725);
or U696 (N_696,In_1421,In_724);
nand U697 (N_697,In_1811,N_339);
nand U698 (N_698,In_1184,In_1682);
xor U699 (N_699,In_1463,In_1426);
and U700 (N_700,In_1411,In_293);
or U701 (N_701,N_257,In_646);
xnor U702 (N_702,N_58,In_1088);
and U703 (N_703,In_1673,In_1544);
or U704 (N_704,In_1316,In_1330);
xnor U705 (N_705,In_804,In_1140);
nand U706 (N_706,In_414,In_831);
or U707 (N_707,In_1803,In_1006);
nand U708 (N_708,In_1495,In_465);
xor U709 (N_709,N_183,N_378);
and U710 (N_710,In_312,In_531);
nor U711 (N_711,N_250,In_1365);
and U712 (N_712,In_956,In_1539);
xnor U713 (N_713,N_254,In_550);
nand U714 (N_714,In_1451,N_184);
xor U715 (N_715,In_690,In_1595);
xor U716 (N_716,In_242,In_195);
and U717 (N_717,In_683,In_1329);
and U718 (N_718,In_1108,In_1063);
nand U719 (N_719,N_376,In_1752);
xor U720 (N_720,In_1808,In_211);
and U721 (N_721,N_363,In_104);
nand U722 (N_722,In_558,N_45);
nand U723 (N_723,In_1859,In_1439);
xor U724 (N_724,In_1899,In_1162);
or U725 (N_725,In_504,In_517);
nand U726 (N_726,In_957,In_1593);
and U727 (N_727,N_174,In_453);
and U728 (N_728,In_1688,N_368);
and U729 (N_729,In_979,N_287);
nor U730 (N_730,N_279,N_75);
nor U731 (N_731,In_1242,In_1762);
and U732 (N_732,In_677,In_1172);
xnor U733 (N_733,In_1398,In_245);
nand U734 (N_734,In_601,In_1676);
xnor U735 (N_735,N_360,N_326);
xnor U736 (N_736,In_745,In_778);
or U737 (N_737,In_693,N_263);
xor U738 (N_738,In_761,In_1486);
xnor U739 (N_739,In_1707,In_1613);
or U740 (N_740,In_1394,In_387);
or U741 (N_741,In_859,In_516);
nor U742 (N_742,In_580,In_1051);
xnor U743 (N_743,In_68,In_457);
nor U744 (N_744,In_1313,N_394);
nand U745 (N_745,In_1064,In_373);
xnor U746 (N_746,In_1413,In_835);
and U747 (N_747,In_927,In_1187);
and U748 (N_748,In_699,In_657);
nor U749 (N_749,In_139,In_372);
and U750 (N_750,N_346,In_1557);
xor U751 (N_751,In_268,N_126);
or U752 (N_752,In_1139,In_1970);
nor U753 (N_753,In_415,N_114);
nor U754 (N_754,In_1932,In_502);
nor U755 (N_755,N_251,In_1628);
and U756 (N_756,In_844,In_705);
and U757 (N_757,In_805,In_408);
nand U758 (N_758,In_496,In_1519);
or U759 (N_759,In_240,N_231);
nor U760 (N_760,In_184,N_332);
nand U761 (N_761,N_301,In_105);
and U762 (N_762,In_1409,In_1738);
nor U763 (N_763,In_1774,In_1026);
nor U764 (N_764,In_1214,In_1968);
and U765 (N_765,In_1085,In_1917);
or U766 (N_766,N_253,In_1813);
nor U767 (N_767,In_928,In_298);
and U768 (N_768,In_665,In_559);
xnor U769 (N_769,In_479,N_239);
nor U770 (N_770,In_227,In_299);
nand U771 (N_771,N_28,In_1975);
and U772 (N_772,In_391,In_1581);
xor U773 (N_773,In_1904,In_89);
nand U774 (N_774,In_898,In_1652);
xnor U775 (N_775,N_91,In_1590);
xnor U776 (N_776,In_36,N_270);
xnor U777 (N_777,N_272,In_1612);
and U778 (N_778,N_216,In_487);
and U779 (N_779,In_1973,In_230);
nor U780 (N_780,In_1254,In_571);
or U781 (N_781,In_1758,In_618);
xor U782 (N_782,In_1385,In_250);
or U783 (N_783,In_1835,In_22);
nand U784 (N_784,N_172,In_1377);
nor U785 (N_785,In_285,N_269);
xor U786 (N_786,N_354,In_1255);
xnor U787 (N_787,In_729,N_241);
nand U788 (N_788,In_1481,N_41);
nand U789 (N_789,In_888,In_667);
nor U790 (N_790,In_1843,In_1068);
nand U791 (N_791,In_513,In_544);
and U792 (N_792,In_1725,In_1178);
xnor U793 (N_793,In_1146,In_1589);
nand U794 (N_794,In_1531,In_902);
nor U795 (N_795,N_121,In_267);
or U796 (N_796,In_1986,In_1327);
xnor U797 (N_797,In_219,N_68);
nand U798 (N_798,In_56,In_524);
and U799 (N_799,N_93,In_783);
or U800 (N_800,N_798,In_1668);
and U801 (N_801,In_530,In_1831);
xnor U802 (N_802,In_1997,In_1535);
and U803 (N_803,N_479,N_316);
nand U804 (N_804,In_1681,In_828);
nand U805 (N_805,In_284,N_17);
or U806 (N_806,In_786,N_632);
or U807 (N_807,N_462,In_858);
and U808 (N_808,N_105,In_162);
and U809 (N_809,In_501,In_766);
nand U810 (N_810,N_573,In_1449);
and U811 (N_811,N_189,In_1393);
xnor U812 (N_812,N_779,N_428);
nor U813 (N_813,In_1744,N_13);
or U814 (N_814,N_390,N_597);
nor U815 (N_815,In_263,In_536);
and U816 (N_816,N_5,N_499);
nor U817 (N_817,In_607,In_1269);
and U818 (N_818,N_580,N_435);
xnor U819 (N_819,N_689,In_893);
nor U820 (N_820,In_348,N_303);
nand U821 (N_821,N_80,In_1791);
and U822 (N_822,In_1167,N_668);
and U823 (N_823,N_730,N_669);
xnor U824 (N_824,In_340,In_572);
and U825 (N_825,N_706,N_90);
xor U826 (N_826,In_434,In_1015);
or U827 (N_827,In_1253,N_99);
xor U828 (N_828,N_247,N_623);
and U829 (N_829,N_476,N_607);
or U830 (N_830,In_974,In_1338);
or U831 (N_831,In_940,In_1028);
xnor U832 (N_832,In_529,N_795);
xnor U833 (N_833,In_58,N_529);
or U834 (N_834,N_671,N_485);
and U835 (N_835,In_1735,N_438);
nand U836 (N_836,In_1382,In_896);
xnor U837 (N_837,In_17,N_94);
xnor U838 (N_838,N_691,In_1080);
or U839 (N_839,N_101,N_444);
nand U840 (N_840,N_217,In_1104);
xor U841 (N_841,N_477,In_873);
nor U842 (N_842,In_280,N_692);
xor U843 (N_843,In_1016,In_39);
xor U844 (N_844,N_638,N_480);
nand U845 (N_845,In_938,N_451);
xnor U846 (N_846,N_686,In_1138);
or U847 (N_847,In_1710,In_671);
xnor U848 (N_848,N_519,N_556);
nand U849 (N_849,In_1833,N_570);
nand U850 (N_850,In_1323,In_1977);
xnor U851 (N_851,N_553,N_786);
nor U852 (N_852,N_108,N_11);
xnor U853 (N_853,In_1516,In_514);
and U854 (N_854,In_953,N_550);
or U855 (N_855,In_649,In_159);
and U856 (N_856,N_587,In_585);
nand U857 (N_857,N_512,N_541);
or U858 (N_858,N_448,In_1965);
or U859 (N_859,N_455,N_432);
nand U860 (N_860,In_1520,N_293);
nand U861 (N_861,In_231,In_972);
or U862 (N_862,N_404,N_723);
nor U863 (N_863,N_643,In_377);
or U864 (N_864,N_624,In_350);
and U865 (N_865,In_794,In_1884);
and U866 (N_866,N_744,N_520);
or U867 (N_867,In_1066,N_522);
nor U868 (N_868,N_571,N_313);
and U869 (N_869,In_849,In_1759);
nor U870 (N_870,N_728,N_646);
xor U871 (N_871,N_421,N_210);
nor U872 (N_872,In_1340,In_1883);
and U873 (N_873,N_318,In_640);
or U874 (N_874,In_556,In_1479);
nand U875 (N_875,N_200,N_586);
and U876 (N_876,N_704,In_166);
and U877 (N_877,In_703,N_653);
nand U878 (N_878,In_534,N_393);
xnor U879 (N_879,In_228,In_753);
nand U880 (N_880,In_967,In_235);
and U881 (N_881,N_14,N_690);
xnor U882 (N_882,In_1076,In_658);
and U883 (N_883,N_402,In_1632);
xnor U884 (N_884,N_746,In_1559);
nor U885 (N_885,N_611,N_411);
nand U886 (N_886,N_353,N_465);
or U887 (N_887,In_484,In_1515);
and U888 (N_888,N_290,In_21);
nand U889 (N_889,N_559,In_456);
xnor U890 (N_890,N_718,In_697);
and U891 (N_891,N_352,N_170);
or U892 (N_892,N_794,In_51);
or U893 (N_893,In_1025,In_635);
nor U894 (N_894,In_1576,In_904);
nor U895 (N_895,N_538,In_702);
xnor U896 (N_896,In_1050,N_507);
and U897 (N_897,N_628,N_478);
or U898 (N_898,N_439,In_1121);
xnor U899 (N_899,N_688,N_540);
nand U900 (N_900,In_679,N_561);
xnor U901 (N_901,N_585,In_302);
nand U902 (N_902,In_887,N_431);
xor U903 (N_903,In_977,In_1579);
xnor U904 (N_904,In_505,In_1369);
or U905 (N_905,In_463,In_973);
or U906 (N_906,In_1510,N_747);
nor U907 (N_907,N_756,In_137);
nand U908 (N_908,In_1036,In_1496);
and U909 (N_909,N_772,N_552);
and U910 (N_910,In_1921,In_907);
and U911 (N_911,In_1916,In_274);
nand U912 (N_912,In_615,In_135);
nand U913 (N_913,In_1801,In_721);
or U914 (N_914,N_349,In_95);
xor U915 (N_915,N_244,In_1375);
or U916 (N_916,N_54,In_125);
xnor U917 (N_917,In_1293,In_911);
xnor U918 (N_918,N_769,N_22);
and U919 (N_919,N_443,In_1819);
or U920 (N_920,In_1532,In_1049);
or U921 (N_921,N_777,N_344);
or U922 (N_922,N_634,In_853);
nand U923 (N_923,In_584,In_1770);
and U924 (N_924,N_365,N_51);
or U925 (N_925,In_1546,In_1487);
nand U926 (N_926,In_474,In_404);
or U927 (N_927,In_1483,N_655);
nor U928 (N_928,N_618,N_136);
or U929 (N_929,N_694,N_763);
xnor U930 (N_930,In_1220,N_535);
and U931 (N_931,In_1828,N_679);
xor U932 (N_932,In_1352,In_1732);
nand U933 (N_933,In_751,N_602);
nor U934 (N_934,N_471,In_1);
nor U935 (N_935,N_474,N_401);
nor U936 (N_936,N_98,N_713);
or U937 (N_937,In_512,In_1548);
nor U938 (N_938,In_878,N_83);
and U939 (N_939,N_588,N_739);
nand U940 (N_940,In_813,In_1454);
nor U941 (N_941,In_815,In_1075);
and U942 (N_942,In_650,In_0);
nor U943 (N_943,N_729,N_238);
nand U944 (N_944,In_400,N_487);
or U945 (N_945,N_648,In_1350);
xor U946 (N_946,N_639,N_500);
nand U947 (N_947,N_714,N_766);
or U948 (N_948,In_1287,N_215);
nand U949 (N_949,N_350,In_871);
nand U950 (N_950,In_236,N_755);
nor U951 (N_951,In_35,N_115);
nand U952 (N_952,N_163,In_866);
nor U953 (N_953,In_1366,N_155);
nand U954 (N_954,N_427,N_409);
or U955 (N_955,N_612,N_486);
nor U956 (N_956,In_975,In_1748);
and U957 (N_957,N_422,N_617);
and U958 (N_958,N_651,In_1202);
and U959 (N_959,In_1203,In_1588);
nor U960 (N_960,N_636,N_659);
and U961 (N_961,N_656,N_436);
nor U962 (N_962,In_1928,In_520);
nand U963 (N_963,In_495,In_37);
nor U964 (N_964,N_470,In_1475);
or U965 (N_965,In_1562,N_491);
xnor U966 (N_966,N_329,In_1001);
or U967 (N_967,N_518,In_1290);
and U968 (N_968,In_1194,In_726);
or U969 (N_969,In_836,N_582);
nand U970 (N_970,N_621,N_457);
or U971 (N_971,In_1697,In_1912);
nand U972 (N_972,In_10,N_128);
xnor U973 (N_973,In_811,In_1273);
or U974 (N_974,In_628,N_400);
nand U975 (N_975,N_726,N_554);
or U976 (N_976,N_367,In_114);
nor U977 (N_977,In_218,In_1911);
or U978 (N_978,In_1780,In_966);
nor U979 (N_979,N_716,N_356);
and U980 (N_980,In_1311,N_389);
or U981 (N_981,N_685,In_1277);
or U982 (N_982,N_654,N_454);
xor U983 (N_983,N_97,In_288);
nand U984 (N_984,N_464,N_591);
or U985 (N_985,In_892,In_239);
nand U986 (N_986,N_568,N_717);
nor U987 (N_987,In_1281,N_410);
xnor U988 (N_988,N_776,In_296);
nand U989 (N_989,N_715,N_168);
nand U990 (N_990,N_564,In_1698);
or U991 (N_991,N_358,N_243);
nand U992 (N_992,In_196,In_1301);
xor U993 (N_993,N_560,In_1256);
xor U994 (N_994,In_191,N_9);
nand U995 (N_995,In_548,In_25);
or U996 (N_996,In_208,In_1137);
or U997 (N_997,N_677,In_1775);
nor U998 (N_998,N_2,In_1055);
nand U999 (N_999,In_16,N_322);
xor U1000 (N_1000,In_696,N_331);
nor U1001 (N_1001,In_1437,In_1685);
nand U1002 (N_1002,In_1720,In_1787);
nor U1003 (N_1003,In_912,N_398);
or U1004 (N_1004,N_460,N_665);
nand U1005 (N_1005,In_692,N_355);
and U1006 (N_1006,In_78,N_473);
and U1007 (N_1007,N_737,N_767);
nor U1008 (N_1008,In_206,In_917);
nor U1009 (N_1009,N_630,N_32);
and U1010 (N_1010,In_1032,In_1462);
xnor U1011 (N_1011,N_749,N_467);
nand U1012 (N_1012,N_445,N_296);
nor U1013 (N_1013,N_525,In_436);
nand U1014 (N_1014,N_534,N_645);
or U1015 (N_1015,N_36,N_562);
and U1016 (N_1016,N_509,N_340);
and U1017 (N_1017,In_889,In_1686);
or U1018 (N_1018,N_413,In_713);
nand U1019 (N_1019,In_561,N_557);
nor U1020 (N_1020,In_1633,In_1298);
or U1021 (N_1021,In_1890,N_530);
xnor U1022 (N_1022,In_320,In_1156);
nor U1023 (N_1023,In_300,In_1217);
nand U1024 (N_1024,N_725,In_1236);
and U1025 (N_1025,In_450,In_223);
nand U1026 (N_1026,N_733,In_1888);
and U1027 (N_1027,N_765,N_330);
or U1028 (N_1028,N_569,In_1918);
and U1029 (N_1029,N_388,N_440);
nor U1030 (N_1030,N_600,N_792);
xor U1031 (N_1031,In_1349,In_1950);
xnor U1032 (N_1032,In_1101,N_204);
xnor U1033 (N_1033,N_770,N_19);
xnor U1034 (N_1034,In_1312,In_121);
or U1035 (N_1035,N_328,In_1837);
and U1036 (N_1036,N_34,In_107);
nand U1037 (N_1037,In_30,In_617);
xor U1038 (N_1038,In_1091,N_761);
and U1039 (N_1039,In_704,In_1966);
nand U1040 (N_1040,In_1680,N_117);
xnor U1041 (N_1041,N_731,N_48);
or U1042 (N_1042,In_613,In_830);
or U1043 (N_1043,N_218,N_768);
nand U1044 (N_1044,N_791,N_282);
nand U1045 (N_1045,N_456,In_1407);
and U1046 (N_1046,N_160,N_419);
or U1047 (N_1047,In_270,N_546);
nand U1048 (N_1048,N_275,In_727);
or U1049 (N_1049,In_1458,N_595);
and U1050 (N_1050,N_528,N_584);
nor U1051 (N_1051,In_991,In_1857);
nand U1052 (N_1052,In_322,In_1880);
nor U1053 (N_1053,In_482,In_281);
and U1054 (N_1054,N_610,N_306);
or U1055 (N_1055,N_357,In_187);
xor U1056 (N_1056,N_762,In_1164);
or U1057 (N_1057,In_1388,In_1113);
nand U1058 (N_1058,N_132,In_397);
nand U1059 (N_1059,In_1651,In_950);
nor U1060 (N_1060,In_75,In_249);
nor U1061 (N_1061,In_597,In_1598);
xor U1062 (N_1062,In_421,In_1907);
xor U1063 (N_1063,N_466,N_506);
or U1064 (N_1064,In_26,N_16);
and U1065 (N_1065,N_721,N_743);
nand U1066 (N_1066,In_1395,N_724);
nand U1067 (N_1067,In_497,In_1416);
nand U1068 (N_1068,In_730,N_505);
xor U1069 (N_1069,N_408,In_294);
or U1070 (N_1070,N_264,In_1773);
nand U1071 (N_1071,N_384,N_619);
nand U1072 (N_1072,N_631,In_429);
nand U1073 (N_1073,In_1392,In_449);
xnor U1074 (N_1074,In_1763,In_467);
xor U1075 (N_1075,N_748,In_710);
nand U1076 (N_1076,In_1003,N_493);
nor U1077 (N_1077,In_795,N_463);
nand U1078 (N_1078,N_510,In_1418);
nand U1079 (N_1079,N_449,In_1713);
or U1080 (N_1080,In_1526,N_370);
or U1081 (N_1081,In_1304,N_543);
nand U1082 (N_1082,N_280,In_1078);
and U1083 (N_1083,N_208,N_343);
xnor U1084 (N_1084,In_1227,N_52);
and U1085 (N_1085,N_195,In_356);
xnor U1086 (N_1086,In_334,In_750);
or U1087 (N_1087,N_236,N_537);
xor U1088 (N_1088,In_212,In_542);
and U1089 (N_1089,N_698,In_466);
or U1090 (N_1090,In_207,In_1692);
xnor U1091 (N_1091,In_1699,In_1224);
nor U1092 (N_1092,In_651,N_361);
nor U1093 (N_1093,In_433,In_1115);
nand U1094 (N_1094,N_185,N_77);
nand U1095 (N_1095,In_608,In_925);
and U1096 (N_1096,N_309,In_1081);
and U1097 (N_1097,In_839,N_274);
nor U1098 (N_1098,N_446,N_177);
or U1099 (N_1099,N_709,N_423);
nand U1100 (N_1100,In_232,N_489);
and U1101 (N_1101,In_1040,N_757);
and U1102 (N_1102,In_264,In_1729);
nand U1103 (N_1103,N_61,N_212);
nand U1104 (N_1104,N_676,N_148);
or U1105 (N_1105,N_539,In_643);
or U1106 (N_1106,N_567,In_1781);
nor U1107 (N_1107,N_407,N_308);
and U1108 (N_1108,N_710,N_785);
nor U1109 (N_1109,In_117,N_650);
xnor U1110 (N_1110,In_639,In_1126);
nand U1111 (N_1111,N_695,N_751);
or U1112 (N_1112,N_707,N_156);
and U1113 (N_1113,In_1043,In_154);
nand U1114 (N_1114,N_314,N_614);
xnor U1115 (N_1115,In_1363,N_483);
and U1116 (N_1116,N_385,In_1530);
nand U1117 (N_1117,N_459,In_678);
xnor U1118 (N_1118,N_1,N_380);
nor U1119 (N_1119,N_592,N_745);
and U1120 (N_1120,N_593,N_442);
xor U1121 (N_1121,N_784,In_627);
xor U1122 (N_1122,N_302,N_548);
and U1123 (N_1123,N_107,N_233);
xnor U1124 (N_1124,In_876,In_1020);
xnor U1125 (N_1125,In_1134,N_754);
xor U1126 (N_1126,In_691,In_1618);
nor U1127 (N_1127,In_1082,N_312);
nor U1128 (N_1128,N_598,In_796);
and U1129 (N_1129,N_517,N_441);
nor U1130 (N_1130,In_94,N_100);
or U1131 (N_1131,N_180,In_1930);
xor U1132 (N_1132,In_122,N_8);
nor U1133 (N_1133,In_468,In_98);
nor U1134 (N_1134,N_793,N_496);
nor U1135 (N_1135,N_248,In_32);
or U1136 (N_1136,N_191,N_601);
nand U1137 (N_1137,In_897,N_536);
or U1138 (N_1138,N_753,N_418);
and U1139 (N_1139,N_187,N_760);
xnor U1140 (N_1140,N_702,N_705);
or U1141 (N_1141,N_750,N_39);
and U1142 (N_1142,In_1700,In_174);
and U1143 (N_1143,In_562,N_708);
nor U1144 (N_1144,N_640,In_1919);
or U1145 (N_1145,N_513,N_414);
nor U1146 (N_1146,N_240,In_863);
or U1147 (N_1147,In_865,In_1695);
or U1148 (N_1148,N_663,N_417);
nand U1149 (N_1149,In_787,N_57);
nor U1150 (N_1150,In_1112,N_635);
xor U1151 (N_1151,In_1096,N_508);
or U1152 (N_1152,In_1701,N_759);
xnor U1153 (N_1153,N_682,N_796);
or U1154 (N_1154,In_946,In_1640);
nand U1155 (N_1155,N_615,In_784);
nand U1156 (N_1156,In_742,In_511);
and U1157 (N_1157,N_625,N_524);
and U1158 (N_1158,N_26,N_494);
or U1159 (N_1159,In_170,In_346);
xor U1160 (N_1160,N_565,In_941);
or U1161 (N_1161,In_392,N_735);
or U1162 (N_1162,In_1263,In_719);
xnor U1163 (N_1163,In_1834,N_616);
nand U1164 (N_1164,N_790,N_12);
and U1165 (N_1165,In_1677,N_426);
and U1166 (N_1166,In_399,N_566);
and U1167 (N_1167,In_451,N_697);
xor U1168 (N_1168,N_629,In_1292);
nand U1169 (N_1169,In_1785,N_289);
xor U1170 (N_1170,In_1887,N_123);
or U1171 (N_1171,N_599,In_1846);
and U1172 (N_1172,In_1879,N_633);
nor U1173 (N_1173,In_1109,In_1708);
and U1174 (N_1174,In_1779,In_13);
xnor U1175 (N_1175,In_716,In_758);
xnor U1176 (N_1176,N_780,In_192);
or U1177 (N_1177,In_1951,N_771);
and U1178 (N_1178,N_192,In_661);
nand U1179 (N_1179,N_604,In_1615);
nand U1180 (N_1180,In_814,In_760);
nor U1181 (N_1181,N_775,N_532);
xnor U1182 (N_1182,N_469,N_558);
and U1183 (N_1183,In_1132,N_262);
and U1184 (N_1184,N_450,N_152);
and U1185 (N_1185,N_683,In_1662);
nand U1186 (N_1186,N_742,N_551);
xor U1187 (N_1187,In_970,N_154);
nand U1188 (N_1188,N_201,N_335);
xnor U1189 (N_1189,N_475,N_603);
and U1190 (N_1190,N_533,N_589);
nor U1191 (N_1191,N_317,N_658);
nor U1192 (N_1192,N_576,N_797);
nor U1193 (N_1193,In_1361,N_672);
nor U1194 (N_1194,N_720,N_641);
xor U1195 (N_1195,N_608,N_497);
xnor U1196 (N_1196,In_1629,In_1569);
xor U1197 (N_1197,N_85,In_1823);
nor U1198 (N_1198,N_44,N_403);
nor U1199 (N_1199,In_1309,N_320);
nand U1200 (N_1200,N_613,N_657);
and U1201 (N_1201,N_140,In_254);
nand U1202 (N_1202,N_924,In_134);
xnor U1203 (N_1203,N_458,N_158);
nand U1204 (N_1204,N_1181,In_1940);
nor U1205 (N_1205,In_1771,N_825);
nand U1206 (N_1206,N_804,N_1091);
xnor U1207 (N_1207,N_1100,In_183);
and U1208 (N_1208,In_603,In_1386);
xnor U1209 (N_1209,N_1187,N_889);
and U1210 (N_1210,N_1017,N_836);
and U1211 (N_1211,N_978,In_1136);
xor U1212 (N_1212,N_1182,N_970);
or U1213 (N_1213,N_788,N_1174);
nand U1214 (N_1214,N_987,N_962);
nor U1215 (N_1215,In_1030,N_963);
nor U1216 (N_1216,In_109,N_661);
nor U1217 (N_1217,N_899,N_622);
nand U1218 (N_1218,N_504,N_1160);
or U1219 (N_1219,In_1093,N_575);
nand U1220 (N_1220,N_495,N_1132);
and U1221 (N_1221,N_860,N_25);
and U1222 (N_1222,N_935,N_859);
xor U1223 (N_1223,N_673,N_461);
nand U1224 (N_1224,In_834,N_817);
nand U1225 (N_1225,N_896,N_781);
nor U1226 (N_1226,N_1113,N_711);
nor U1227 (N_1227,N_297,N_865);
xor U1228 (N_1228,N_972,N_542);
or U1229 (N_1229,N_903,N_327);
nor U1230 (N_1230,N_503,N_590);
nand U1231 (N_1231,N_1128,N_1010);
nand U1232 (N_1232,N_960,In_868);
nor U1233 (N_1233,N_1120,N_1111);
xnor U1234 (N_1234,N_722,N_1038);
nor U1235 (N_1235,N_1008,N_6);
and U1236 (N_1236,N_916,N_928);
xor U1237 (N_1237,N_424,In_1052);
and U1238 (N_1238,In_113,In_619);
nor U1239 (N_1239,N_547,N_387);
xor U1240 (N_1240,N_305,N_447);
xnor U1241 (N_1241,In_45,N_773);
xor U1242 (N_1242,N_835,N_696);
nor U1243 (N_1243,N_1068,In_1039);
nand U1244 (N_1244,In_1485,N_1095);
nor U1245 (N_1245,N_902,N_1050);
nor U1246 (N_1246,N_894,N_1196);
nor U1247 (N_1247,N_814,N_1150);
and U1248 (N_1248,In_84,N_1199);
nor U1249 (N_1249,N_674,N_898);
and U1250 (N_1250,N_843,In_410);
or U1251 (N_1251,In_259,N_1109);
nand U1252 (N_1252,In_452,N_53);
nor U1253 (N_1253,In_609,In_180);
nand U1254 (N_1254,N_81,N_989);
nand U1255 (N_1255,In_38,N_869);
xor U1256 (N_1256,N_823,N_855);
xnor U1257 (N_1257,In_590,In_1276);
xnor U1258 (N_1258,N_235,N_1134);
nand U1259 (N_1259,N_936,N_103);
nor U1260 (N_1260,N_1048,In_233);
nand U1261 (N_1261,In_694,N_652);
xnor U1262 (N_1262,N_862,In_1869);
or U1263 (N_1263,N_1164,N_1157);
nand U1264 (N_1264,In_1983,N_1082);
or U1265 (N_1265,N_809,N_62);
or U1266 (N_1266,In_891,In_629);
xor U1267 (N_1267,N_853,In_900);
xnor U1268 (N_1268,In_478,N_841);
nand U1269 (N_1269,N_895,N_911);
nand U1270 (N_1270,N_555,N_1012);
and U1271 (N_1271,N_941,In_782);
and U1272 (N_1272,N_1186,N_1125);
or U1273 (N_1273,N_1135,In_700);
nand U1274 (N_1274,N_1178,N_662);
nand U1275 (N_1275,N_1032,N_909);
nor U1276 (N_1276,N_912,N_1141);
nor U1277 (N_1277,N_995,N_95);
or U1278 (N_1278,N_799,N_1108);
and U1279 (N_1279,N_866,N_490);
xnor U1280 (N_1280,N_983,In_569);
nor U1281 (N_1281,N_1074,N_701);
and U1282 (N_1282,N_1153,In_1900);
nand U1283 (N_1283,In_1906,N_1115);
nand U1284 (N_1284,N_783,N_990);
xnor U1285 (N_1285,N_545,N_1004);
and U1286 (N_1286,N_15,In_1941);
or U1287 (N_1287,N_881,N_1000);
nor U1288 (N_1288,N_920,N_572);
nor U1289 (N_1289,N_808,In_381);
xnor U1290 (N_1290,N_727,In_370);
nor U1291 (N_1291,N_1170,N_849);
nor U1292 (N_1292,N_1051,In_42);
and U1293 (N_1293,N_1148,N_666);
nand U1294 (N_1294,N_169,N_429);
nand U1295 (N_1295,N_877,N_815);
or U1296 (N_1296,N_922,N_985);
or U1297 (N_1297,N_1195,In_173);
nand U1298 (N_1298,N_945,N_40);
and U1299 (N_1299,In_1567,N_1173);
nor U1300 (N_1300,In_1687,In_914);
or U1301 (N_1301,N_1177,N_1029);
and U1302 (N_1302,N_1027,N_359);
nand U1303 (N_1303,N_734,In_1669);
nor U1304 (N_1304,N_1042,N_845);
or U1305 (N_1305,N_829,In_1125);
nor U1306 (N_1306,N_234,N_863);
xnor U1307 (N_1307,N_947,N_940);
nor U1308 (N_1308,N_47,N_789);
xor U1309 (N_1309,N_1156,N_594);
xnor U1310 (N_1310,N_1147,N_967);
nor U1311 (N_1311,N_637,N_481);
and U1312 (N_1312,In_1675,In_775);
and U1313 (N_1313,N_937,In_378);
or U1314 (N_1314,N_930,In_701);
nor U1315 (N_1315,In_525,In_1509);
nand U1316 (N_1316,N_1175,In_345);
or U1317 (N_1317,N_1163,N_131);
and U1318 (N_1318,N_291,In_1238);
and U1319 (N_1319,N_1101,N_1024);
xnor U1320 (N_1320,N_1072,N_848);
or U1321 (N_1321,N_205,In_1012);
or U1322 (N_1322,N_1116,N_918);
nand U1323 (N_1323,N_1180,N_482);
nand U1324 (N_1324,In_1471,N_1040);
or U1325 (N_1325,In_1561,N_880);
nand U1326 (N_1326,N_1098,N_805);
xor U1327 (N_1327,N_207,In_118);
and U1328 (N_1328,In_488,N_738);
xor U1329 (N_1329,N_965,N_55);
xnor U1330 (N_1330,N_84,N_732);
xor U1331 (N_1331,In_1460,N_113);
or U1332 (N_1332,N_931,N_906);
and U1333 (N_1333,In_748,In_1452);
or U1334 (N_1334,N_498,In_1740);
nor U1335 (N_1335,N_961,N_374);
xor U1336 (N_1336,N_801,In_1018);
nand U1337 (N_1337,N_265,N_284);
and U1338 (N_1338,In_875,N_256);
nor U1339 (N_1339,N_758,N_907);
nand U1340 (N_1340,N_951,N_812);
and U1341 (N_1341,N_981,In_1337);
xnor U1342 (N_1342,N_973,N_577);
nand U1343 (N_1343,N_1064,In_1205);
nor U1344 (N_1344,In_850,N_1022);
or U1345 (N_1345,In_1244,N_531);
or U1346 (N_1346,N_1028,N_800);
nor U1347 (N_1347,N_678,N_974);
or U1348 (N_1348,In_685,In_936);
xor U1349 (N_1349,N_703,N_667);
xor U1350 (N_1350,In_793,N_670);
or U1351 (N_1351,N_774,In_1059);
and U1352 (N_1352,In_1339,N_221);
nand U1353 (N_1353,N_647,N_523);
nand U1354 (N_1354,In_500,N_926);
xnor U1355 (N_1355,N_917,N_229);
nand U1356 (N_1356,In_483,In_248);
xnor U1357 (N_1357,In_1795,N_660);
and U1358 (N_1358,N_878,N_1105);
or U1359 (N_1359,N_802,N_992);
nor U1360 (N_1360,N_1142,In_1403);
or U1361 (N_1361,In_1467,In_611);
and U1362 (N_1362,N_472,N_1037);
or U1363 (N_1363,N_1081,N_311);
or U1364 (N_1364,In_140,N_991);
nor U1365 (N_1365,N_986,N_871);
and U1366 (N_1366,N_684,N_856);
nor U1367 (N_1367,N_348,N_1118);
and U1368 (N_1368,N_122,In_741);
xor U1369 (N_1369,N_1071,In_1789);
nand U1370 (N_1370,N_816,N_741);
and U1371 (N_1371,N_958,In_1092);
nand U1372 (N_1372,N_910,N_1192);
or U1373 (N_1373,N_1015,N_1014);
or U1374 (N_1374,N_919,N_1198);
xnor U1375 (N_1375,N_64,N_488);
xor U1376 (N_1376,N_813,N_1171);
nand U1377 (N_1377,In_1342,In_877);
nand U1378 (N_1378,In_1200,N_596);
xor U1379 (N_1379,N_1126,In_349);
xor U1380 (N_1380,In_919,In_785);
xor U1381 (N_1381,N_1070,N_1011);
xnor U1382 (N_1382,N_124,N_1059);
or U1383 (N_1383,N_1054,N_579);
or U1384 (N_1384,N_925,In_384);
nor U1385 (N_1385,In_998,In_110);
nand U1386 (N_1386,N_832,N_834);
nor U1387 (N_1387,In_1182,N_1033);
nand U1388 (N_1388,N_1197,N_159);
and U1389 (N_1389,N_994,N_153);
nor U1390 (N_1390,N_975,N_1007);
or U1391 (N_1391,N_56,N_933);
nand U1392 (N_1392,N_399,N_1103);
nor U1393 (N_1393,N_851,N_891);
xnor U1394 (N_1394,N_782,In_126);
and U1395 (N_1395,In_1799,N_1021);
nor U1396 (N_1396,N_1046,N_885);
nand U1397 (N_1397,N_644,N_1045);
or U1398 (N_1398,N_1121,N_977);
and U1399 (N_1399,N_1035,N_1047);
or U1400 (N_1400,In_1655,N_430);
xnor U1401 (N_1401,In_62,N_1030);
nor U1402 (N_1402,N_839,N_642);
or U1403 (N_1403,N_415,N_1026);
nand U1404 (N_1404,N_433,In_1745);
xor U1405 (N_1405,N_347,N_831);
or U1406 (N_1406,N_627,In_1889);
nand U1407 (N_1407,N_950,N_886);
nand U1408 (N_1408,N_1152,In_1233);
nor U1409 (N_1409,In_1778,N_955);
xnor U1410 (N_1410,In_982,N_675);
and U1411 (N_1411,N_1090,N_664);
or U1412 (N_1412,N_1119,N_687);
xor U1413 (N_1413,N_24,N_897);
and U1414 (N_1414,N_605,N_1191);
nor U1415 (N_1415,In_1974,N_406);
xor U1416 (N_1416,N_1190,In_1166);
nand U1417 (N_1417,N_219,N_281);
or U1418 (N_1418,N_516,N_1075);
nand U1419 (N_1419,N_1025,N_1086);
and U1420 (N_1420,N_1139,N_904);
or U1421 (N_1421,N_953,N_943);
or U1422 (N_1422,N_861,In_1492);
xor U1423 (N_1423,N_700,N_984);
nand U1424 (N_1424,N_997,N_929);
and U1425 (N_1425,N_699,In_437);
nor U1426 (N_1426,In_1367,N_858);
xnor U1427 (N_1427,N_1001,N_1066);
xnor U1428 (N_1428,N_333,In_1423);
nand U1429 (N_1429,N_712,N_870);
nand U1430 (N_1430,In_765,N_1020);
or U1431 (N_1431,N_1052,N_887);
and U1432 (N_1432,N_719,N_118);
and U1433 (N_1433,N_1154,N_980);
xor U1434 (N_1434,N_1080,In_969);
xnor U1435 (N_1435,N_828,N_30);
nand U1436 (N_1436,N_43,In_841);
and U1437 (N_1437,In_1181,N_193);
nor U1438 (N_1438,N_1131,N_913);
or U1439 (N_1439,N_1151,N_1041);
and U1440 (N_1440,N_266,N_549);
and U1441 (N_1441,N_511,N_693);
and U1442 (N_1442,In_1821,N_908);
or U1443 (N_1443,In_602,N_948);
or U1444 (N_1444,In_157,N_956);
or U1445 (N_1445,N_764,N_944);
or U1446 (N_1446,In_533,N_1060);
nand U1447 (N_1447,N_581,N_1194);
or U1448 (N_1448,N_33,N_1102);
nand U1449 (N_1449,N_1165,In_997);
or U1450 (N_1450,N_521,N_1137);
xor U1451 (N_1451,N_957,N_412);
xnor U1452 (N_1452,N_186,In_1507);
xor U1453 (N_1453,N_778,N_1044);
nand U1454 (N_1454,N_923,In_213);
or U1455 (N_1455,N_1133,N_1055);
and U1456 (N_1456,N_391,N_59);
xor U1457 (N_1457,N_979,N_1129);
and U1458 (N_1458,In_1627,N_1073);
or U1459 (N_1459,In_1383,N_1078);
xor U1460 (N_1460,N_1062,N_526);
nand U1461 (N_1461,N_211,In_1571);
nor U1462 (N_1462,N_181,N_681);
or U1463 (N_1463,In_1357,N_736);
nor U1464 (N_1464,N_405,N_1009);
nand U1465 (N_1465,In_882,N_842);
or U1466 (N_1466,N_468,N_752);
xnor U1467 (N_1467,N_921,N_649);
nand U1468 (N_1468,N_982,N_819);
and U1469 (N_1469,N_1063,N_267);
and U1470 (N_1470,N_502,N_939);
xor U1471 (N_1471,N_1172,N_1031);
and U1472 (N_1472,N_1013,N_1099);
nor U1473 (N_1473,N_1053,In_1384);
nand U1474 (N_1474,In_1893,In_1741);
xor U1475 (N_1475,N_1005,In_1954);
and U1476 (N_1476,In_1250,N_1112);
nand U1477 (N_1477,N_1034,In_728);
or U1478 (N_1478,N_833,N_821);
or U1479 (N_1479,N_109,N_1110);
xor U1480 (N_1480,N_803,In_1992);
nor U1481 (N_1481,N_514,N_946);
nor U1482 (N_1482,N_1092,N_386);
or U1483 (N_1483,N_21,In_443);
and U1484 (N_1484,In_1772,N_1167);
nand U1485 (N_1485,N_914,In_923);
or U1486 (N_1486,In_52,N_1104);
xor U1487 (N_1487,N_1188,N_954);
xor U1488 (N_1488,N_1184,N_949);
and U1489 (N_1489,N_806,N_905);
nor U1490 (N_1490,N_1093,N_838);
nor U1491 (N_1491,N_1168,N_876);
nand U1492 (N_1492,N_102,N_847);
nor U1493 (N_1493,In_1878,N_1144);
nand U1494 (N_1494,N_334,N_1124);
nor U1495 (N_1495,N_1162,N_822);
nand U1496 (N_1496,In_1660,In_1980);
xnor U1497 (N_1497,In_1024,N_65);
or U1498 (N_1498,In_992,N_178);
nor U1499 (N_1499,N_840,In_1905);
nor U1500 (N_1500,N_1145,N_515);
nand U1501 (N_1501,N_261,N_850);
nand U1502 (N_1502,N_453,N_999);
xnor U1503 (N_1503,In_175,N_874);
and U1504 (N_1504,In_1444,N_484);
or U1505 (N_1505,N_857,In_528);
nor U1506 (N_1506,N_1161,In_1240);
xnor U1507 (N_1507,N_1127,N_1069);
xnor U1508 (N_1508,N_1003,N_18);
and U1509 (N_1509,In_1207,N_971);
nand U1510 (N_1510,In_167,N_139);
xor U1511 (N_1511,N_1067,N_1107);
nor U1512 (N_1512,In_1102,N_1136);
xor U1513 (N_1513,N_1087,In_1493);
xor U1514 (N_1514,N_811,N_942);
nand U1515 (N_1515,N_988,In_1447);
nor U1516 (N_1516,N_852,In_344);
nor U1517 (N_1517,N_900,N_867);
or U1518 (N_1518,N_206,In_592);
or U1519 (N_1519,N_437,N_1149);
nor U1520 (N_1520,N_606,N_1096);
nor U1521 (N_1521,N_810,N_915);
nor U1522 (N_1522,In_1702,N_1056);
or U1523 (N_1523,N_527,N_844);
nand U1524 (N_1524,N_1179,N_1083);
or U1525 (N_1525,N_1143,N_820);
or U1526 (N_1526,N_1088,In_1002);
or U1527 (N_1527,N_934,In_1897);
or U1528 (N_1528,In_1914,N_175);
nand U1529 (N_1529,N_1076,N_583);
nor U1530 (N_1530,N_609,N_1097);
or U1531 (N_1531,N_420,In_389);
and U1532 (N_1532,In_1158,In_1280);
xor U1533 (N_1533,N_787,In_1266);
or U1534 (N_1534,N_959,In_1981);
nor U1535 (N_1535,N_1016,In_1320);
and U1536 (N_1536,N_89,N_868);
nand U1537 (N_1537,N_1077,N_492);
nor U1538 (N_1538,N_818,N_966);
nor U1539 (N_1539,N_1043,N_578);
nor U1540 (N_1540,N_1094,In_867);
nor U1541 (N_1541,N_890,N_46);
xnor U1542 (N_1542,N_501,N_893);
nand U1543 (N_1543,N_452,N_1023);
xor U1544 (N_1544,N_892,N_1019);
and U1545 (N_1545,N_837,N_1130);
and U1546 (N_1546,N_1140,In_965);
and U1547 (N_1547,N_1089,N_883);
nand U1548 (N_1548,N_0,N_938);
or U1549 (N_1549,N_1036,N_1079);
xor U1550 (N_1550,N_827,N_1189);
xor U1551 (N_1551,N_147,N_873);
nand U1552 (N_1552,N_964,In_341);
nor U1553 (N_1553,In_67,In_652);
and U1554 (N_1554,N_996,N_1185);
or U1555 (N_1555,In_541,N_1146);
or U1556 (N_1556,N_167,N_425);
and U1557 (N_1557,N_952,In_1192);
or U1558 (N_1558,In_1086,N_246);
and U1559 (N_1559,N_968,N_1061);
xor U1560 (N_1560,N_824,N_369);
and U1561 (N_1561,N_620,N_830);
nor U1562 (N_1562,N_1138,In_586);
and U1563 (N_1563,N_969,N_680);
xor U1564 (N_1564,N_888,N_1039);
and U1565 (N_1565,N_1057,N_1166);
nand U1566 (N_1566,N_1122,N_1018);
and U1567 (N_1567,N_1085,In_947);
nor U1568 (N_1568,N_976,N_416);
or U1569 (N_1569,N_884,N_364);
or U1570 (N_1570,N_872,N_1193);
nor U1571 (N_1571,N_1106,N_119);
xnor U1572 (N_1572,N_1117,N_1114);
nor U1573 (N_1573,N_1169,In_532);
and U1574 (N_1574,In_1726,N_879);
nor U1575 (N_1575,N_875,In_1665);
or U1576 (N_1576,In_1168,N_1084);
nand U1577 (N_1577,In_747,N_882);
nor U1578 (N_1578,N_826,N_214);
or U1579 (N_1579,N_60,N_864);
nor U1580 (N_1580,N_927,N_1158);
nor U1581 (N_1581,N_1183,In_606);
or U1582 (N_1582,N_1155,In_460);
or U1583 (N_1583,N_29,N_998);
nand U1584 (N_1584,N_1123,N_146);
nand U1585 (N_1585,In_1218,N_1049);
nor U1586 (N_1586,In_847,N_1006);
xor U1587 (N_1587,N_69,N_993);
and U1588 (N_1588,In_1826,N_901);
nor U1589 (N_1589,N_1058,N_1002);
or U1590 (N_1590,N_626,N_188);
xor U1591 (N_1591,In_625,N_846);
or U1592 (N_1592,N_434,In_1856);
nor U1593 (N_1593,N_1065,N_1159);
xnor U1594 (N_1594,N_740,In_1634);
xor U1595 (N_1595,N_203,N_544);
nand U1596 (N_1596,N_854,In_711);
nor U1597 (N_1597,N_563,N_932);
xnor U1598 (N_1598,N_1176,N_807);
and U1599 (N_1599,N_574,In_1619);
or U1600 (N_1600,N_1296,N_1377);
and U1601 (N_1601,N_1262,N_1385);
and U1602 (N_1602,N_1384,N_1362);
or U1603 (N_1603,N_1520,N_1367);
nor U1604 (N_1604,N_1595,N_1457);
nand U1605 (N_1605,N_1229,N_1586);
or U1606 (N_1606,N_1577,N_1331);
nand U1607 (N_1607,N_1318,N_1383);
nor U1608 (N_1608,N_1584,N_1509);
nand U1609 (N_1609,N_1363,N_1414);
and U1610 (N_1610,N_1329,N_1497);
nor U1611 (N_1611,N_1312,N_1568);
nand U1612 (N_1612,N_1453,N_1592);
nand U1613 (N_1613,N_1437,N_1463);
nor U1614 (N_1614,N_1458,N_1292);
xnor U1615 (N_1615,N_1464,N_1371);
nand U1616 (N_1616,N_1373,N_1476);
nand U1617 (N_1617,N_1554,N_1369);
xnor U1618 (N_1618,N_1451,N_1534);
and U1619 (N_1619,N_1308,N_1269);
nor U1620 (N_1620,N_1200,N_1250);
or U1621 (N_1621,N_1465,N_1215);
xor U1622 (N_1622,N_1406,N_1306);
or U1623 (N_1623,N_1533,N_1264);
or U1624 (N_1624,N_1452,N_1526);
xnor U1625 (N_1625,N_1543,N_1222);
xnor U1626 (N_1626,N_1338,N_1203);
nand U1627 (N_1627,N_1237,N_1540);
and U1628 (N_1628,N_1395,N_1346);
xor U1629 (N_1629,N_1583,N_1320);
or U1630 (N_1630,N_1443,N_1211);
nand U1631 (N_1631,N_1496,N_1353);
and U1632 (N_1632,N_1302,N_1455);
nand U1633 (N_1633,N_1501,N_1223);
or U1634 (N_1634,N_1295,N_1566);
xor U1635 (N_1635,N_1252,N_1322);
xnor U1636 (N_1636,N_1500,N_1396);
or U1637 (N_1637,N_1364,N_1472);
nor U1638 (N_1638,N_1488,N_1251);
nand U1639 (N_1639,N_1404,N_1527);
and U1640 (N_1640,N_1254,N_1206);
nand U1641 (N_1641,N_1432,N_1265);
nor U1642 (N_1642,N_1522,N_1301);
or U1643 (N_1643,N_1557,N_1505);
and U1644 (N_1644,N_1475,N_1585);
nor U1645 (N_1645,N_1281,N_1575);
nand U1646 (N_1646,N_1562,N_1234);
xnor U1647 (N_1647,N_1518,N_1340);
nor U1648 (N_1648,N_1286,N_1225);
nor U1649 (N_1649,N_1298,N_1521);
nor U1650 (N_1650,N_1293,N_1567);
and U1651 (N_1651,N_1227,N_1220);
nor U1652 (N_1652,N_1244,N_1544);
or U1653 (N_1653,N_1291,N_1563);
or U1654 (N_1654,N_1548,N_1224);
xor U1655 (N_1655,N_1310,N_1282);
nor U1656 (N_1656,N_1305,N_1307);
xor U1657 (N_1657,N_1528,N_1564);
and U1658 (N_1658,N_1415,N_1366);
nand U1659 (N_1659,N_1515,N_1311);
nor U1660 (N_1660,N_1536,N_1235);
xnor U1661 (N_1661,N_1506,N_1428);
nor U1662 (N_1662,N_1560,N_1429);
or U1663 (N_1663,N_1398,N_1394);
xnor U1664 (N_1664,N_1407,N_1402);
and U1665 (N_1665,N_1449,N_1438);
and U1666 (N_1666,N_1423,N_1596);
or U1667 (N_1667,N_1579,N_1593);
nor U1668 (N_1668,N_1448,N_1261);
xor U1669 (N_1669,N_1558,N_1571);
xnor U1670 (N_1670,N_1489,N_1258);
nand U1671 (N_1671,N_1469,N_1487);
nor U1672 (N_1672,N_1454,N_1350);
and U1673 (N_1673,N_1594,N_1445);
or U1674 (N_1674,N_1442,N_1565);
and U1675 (N_1675,N_1321,N_1470);
xor U1676 (N_1676,N_1493,N_1559);
nand U1677 (N_1677,N_1208,N_1349);
or U1678 (N_1678,N_1341,N_1555);
or U1679 (N_1679,N_1513,N_1283);
and U1680 (N_1680,N_1332,N_1273);
xnor U1681 (N_1681,N_1374,N_1326);
nor U1682 (N_1682,N_1249,N_1551);
xnor U1683 (N_1683,N_1379,N_1263);
and U1684 (N_1684,N_1217,N_1473);
or U1685 (N_1685,N_1532,N_1257);
nand U1686 (N_1686,N_1380,N_1529);
nor U1687 (N_1687,N_1337,N_1356);
nor U1688 (N_1688,N_1360,N_1289);
nor U1689 (N_1689,N_1446,N_1433);
nand U1690 (N_1690,N_1477,N_1492);
and U1691 (N_1691,N_1504,N_1545);
and U1692 (N_1692,N_1430,N_1248);
xor U1693 (N_1693,N_1403,N_1230);
nand U1694 (N_1694,N_1315,N_1507);
nor U1695 (N_1695,N_1347,N_1351);
and U1696 (N_1696,N_1270,N_1569);
nor U1697 (N_1697,N_1212,N_1421);
xnor U1698 (N_1698,N_1354,N_1556);
or U1699 (N_1699,N_1440,N_1549);
or U1700 (N_1700,N_1239,N_1255);
or U1701 (N_1701,N_1519,N_1578);
or U1702 (N_1702,N_1355,N_1561);
or U1703 (N_1703,N_1238,N_1400);
xor U1704 (N_1704,N_1344,N_1274);
and U1705 (N_1705,N_1570,N_1219);
nand U1706 (N_1706,N_1241,N_1267);
nor U1707 (N_1707,N_1462,N_1524);
nand U1708 (N_1708,N_1378,N_1266);
nor U1709 (N_1709,N_1553,N_1348);
or U1710 (N_1710,N_1277,N_1461);
nand U1711 (N_1711,N_1427,N_1372);
xor U1712 (N_1712,N_1375,N_1231);
nand U1713 (N_1713,N_1580,N_1323);
nand U1714 (N_1714,N_1581,N_1368);
xnor U1715 (N_1715,N_1299,N_1479);
or U1716 (N_1716,N_1358,N_1508);
xnor U1717 (N_1717,N_1253,N_1468);
and U1718 (N_1718,N_1303,N_1214);
and U1719 (N_1719,N_1202,N_1478);
xor U1720 (N_1720,N_1588,N_1444);
or U1721 (N_1721,N_1459,N_1491);
nand U1722 (N_1722,N_1242,N_1447);
and U1723 (N_1723,N_1345,N_1539);
xnor U1724 (N_1724,N_1409,N_1330);
xor U1725 (N_1725,N_1480,N_1236);
nor U1726 (N_1726,N_1300,N_1376);
and U1727 (N_1727,N_1268,N_1550);
xnor U1728 (N_1728,N_1436,N_1247);
xnor U1729 (N_1729,N_1297,N_1399);
and U1730 (N_1730,N_1413,N_1598);
and U1731 (N_1731,N_1483,N_1397);
nand U1732 (N_1732,N_1393,N_1359);
nor U1733 (N_1733,N_1205,N_1523);
nor U1734 (N_1734,N_1386,N_1481);
or U1735 (N_1735,N_1466,N_1294);
nor U1736 (N_1736,N_1499,N_1391);
nor U1737 (N_1737,N_1390,N_1304);
xor U1738 (N_1738,N_1228,N_1343);
xnor U1739 (N_1739,N_1514,N_1490);
and U1740 (N_1740,N_1256,N_1284);
nand U1741 (N_1741,N_1275,N_1599);
nor U1742 (N_1742,N_1552,N_1495);
nor U1743 (N_1743,N_1582,N_1342);
nand U1744 (N_1744,N_1510,N_1309);
and U1745 (N_1745,N_1426,N_1213);
and U1746 (N_1746,N_1285,N_1313);
or U1747 (N_1747,N_1334,N_1482);
or U1748 (N_1748,N_1417,N_1485);
or U1749 (N_1749,N_1381,N_1226);
xor U1750 (N_1750,N_1216,N_1232);
or U1751 (N_1751,N_1387,N_1240);
nor U1752 (N_1752,N_1271,N_1339);
or U1753 (N_1753,N_1530,N_1410);
nand U1754 (N_1754,N_1319,N_1576);
nor U1755 (N_1755,N_1498,N_1572);
or U1756 (N_1756,N_1486,N_1537);
xnor U1757 (N_1757,N_1218,N_1209);
and U1758 (N_1758,N_1280,N_1370);
or U1759 (N_1759,N_1535,N_1434);
nand U1760 (N_1760,N_1547,N_1516);
or U1761 (N_1761,N_1365,N_1233);
and U1762 (N_1762,N_1474,N_1531);
or U1763 (N_1763,N_1333,N_1260);
and U1764 (N_1764,N_1538,N_1401);
nand U1765 (N_1765,N_1431,N_1589);
xor U1766 (N_1766,N_1591,N_1336);
nand U1767 (N_1767,N_1456,N_1288);
or U1768 (N_1768,N_1494,N_1422);
xor U1769 (N_1769,N_1411,N_1278);
or U1770 (N_1770,N_1512,N_1388);
and U1771 (N_1771,N_1335,N_1587);
nand U1772 (N_1772,N_1467,N_1574);
or U1773 (N_1773,N_1361,N_1525);
xor U1774 (N_1774,N_1420,N_1352);
nand U1775 (N_1775,N_1542,N_1357);
and U1776 (N_1776,N_1408,N_1419);
xor U1777 (N_1777,N_1597,N_1450);
nand U1778 (N_1778,N_1327,N_1221);
or U1779 (N_1779,N_1317,N_1287);
or U1780 (N_1780,N_1245,N_1416);
nand U1781 (N_1781,N_1511,N_1314);
xor U1782 (N_1782,N_1418,N_1590);
or U1783 (N_1783,N_1435,N_1503);
and U1784 (N_1784,N_1541,N_1201);
nor U1785 (N_1785,N_1259,N_1441);
nand U1786 (N_1786,N_1246,N_1424);
or U1787 (N_1787,N_1382,N_1412);
and U1788 (N_1788,N_1405,N_1204);
or U1789 (N_1789,N_1272,N_1392);
nand U1790 (N_1790,N_1276,N_1279);
or U1791 (N_1791,N_1324,N_1325);
or U1792 (N_1792,N_1207,N_1471);
nor U1793 (N_1793,N_1502,N_1210);
nor U1794 (N_1794,N_1425,N_1484);
nor U1795 (N_1795,N_1328,N_1316);
or U1796 (N_1796,N_1290,N_1460);
nand U1797 (N_1797,N_1573,N_1517);
or U1798 (N_1798,N_1546,N_1439);
nand U1799 (N_1799,N_1389,N_1243);
nand U1800 (N_1800,N_1364,N_1378);
and U1801 (N_1801,N_1276,N_1222);
xor U1802 (N_1802,N_1441,N_1551);
nand U1803 (N_1803,N_1479,N_1257);
nand U1804 (N_1804,N_1572,N_1237);
or U1805 (N_1805,N_1207,N_1594);
nand U1806 (N_1806,N_1466,N_1276);
nand U1807 (N_1807,N_1533,N_1325);
nor U1808 (N_1808,N_1305,N_1274);
and U1809 (N_1809,N_1412,N_1564);
or U1810 (N_1810,N_1437,N_1364);
xor U1811 (N_1811,N_1255,N_1236);
and U1812 (N_1812,N_1401,N_1434);
xor U1813 (N_1813,N_1379,N_1393);
nand U1814 (N_1814,N_1409,N_1486);
nand U1815 (N_1815,N_1435,N_1313);
nor U1816 (N_1816,N_1320,N_1294);
or U1817 (N_1817,N_1472,N_1569);
nand U1818 (N_1818,N_1583,N_1409);
or U1819 (N_1819,N_1209,N_1488);
or U1820 (N_1820,N_1421,N_1342);
xnor U1821 (N_1821,N_1402,N_1464);
and U1822 (N_1822,N_1318,N_1582);
and U1823 (N_1823,N_1348,N_1420);
and U1824 (N_1824,N_1323,N_1499);
nor U1825 (N_1825,N_1300,N_1279);
or U1826 (N_1826,N_1331,N_1252);
or U1827 (N_1827,N_1386,N_1363);
or U1828 (N_1828,N_1329,N_1400);
or U1829 (N_1829,N_1410,N_1228);
and U1830 (N_1830,N_1221,N_1507);
and U1831 (N_1831,N_1505,N_1590);
and U1832 (N_1832,N_1250,N_1370);
or U1833 (N_1833,N_1596,N_1294);
nand U1834 (N_1834,N_1482,N_1485);
or U1835 (N_1835,N_1270,N_1255);
or U1836 (N_1836,N_1455,N_1317);
nor U1837 (N_1837,N_1419,N_1389);
and U1838 (N_1838,N_1314,N_1244);
nor U1839 (N_1839,N_1529,N_1389);
nand U1840 (N_1840,N_1531,N_1264);
and U1841 (N_1841,N_1549,N_1484);
xnor U1842 (N_1842,N_1453,N_1226);
or U1843 (N_1843,N_1535,N_1226);
or U1844 (N_1844,N_1529,N_1209);
nor U1845 (N_1845,N_1528,N_1378);
xor U1846 (N_1846,N_1344,N_1261);
nor U1847 (N_1847,N_1217,N_1554);
and U1848 (N_1848,N_1569,N_1480);
and U1849 (N_1849,N_1415,N_1582);
or U1850 (N_1850,N_1209,N_1223);
nor U1851 (N_1851,N_1556,N_1562);
nor U1852 (N_1852,N_1313,N_1261);
or U1853 (N_1853,N_1273,N_1442);
nand U1854 (N_1854,N_1457,N_1523);
or U1855 (N_1855,N_1430,N_1573);
and U1856 (N_1856,N_1506,N_1408);
and U1857 (N_1857,N_1200,N_1234);
or U1858 (N_1858,N_1538,N_1301);
nand U1859 (N_1859,N_1404,N_1309);
xnor U1860 (N_1860,N_1566,N_1431);
and U1861 (N_1861,N_1436,N_1283);
xnor U1862 (N_1862,N_1398,N_1222);
nand U1863 (N_1863,N_1511,N_1518);
or U1864 (N_1864,N_1314,N_1493);
xnor U1865 (N_1865,N_1468,N_1396);
and U1866 (N_1866,N_1289,N_1469);
xor U1867 (N_1867,N_1432,N_1375);
and U1868 (N_1868,N_1201,N_1387);
nor U1869 (N_1869,N_1466,N_1420);
nor U1870 (N_1870,N_1222,N_1403);
nand U1871 (N_1871,N_1225,N_1422);
and U1872 (N_1872,N_1385,N_1300);
nand U1873 (N_1873,N_1289,N_1490);
xnor U1874 (N_1874,N_1381,N_1481);
nand U1875 (N_1875,N_1512,N_1400);
nand U1876 (N_1876,N_1466,N_1342);
and U1877 (N_1877,N_1209,N_1410);
nand U1878 (N_1878,N_1359,N_1365);
and U1879 (N_1879,N_1541,N_1431);
xor U1880 (N_1880,N_1315,N_1283);
nor U1881 (N_1881,N_1586,N_1588);
nor U1882 (N_1882,N_1599,N_1587);
or U1883 (N_1883,N_1357,N_1221);
and U1884 (N_1884,N_1217,N_1293);
or U1885 (N_1885,N_1453,N_1216);
or U1886 (N_1886,N_1595,N_1265);
or U1887 (N_1887,N_1398,N_1462);
and U1888 (N_1888,N_1364,N_1225);
nand U1889 (N_1889,N_1228,N_1452);
and U1890 (N_1890,N_1518,N_1381);
nor U1891 (N_1891,N_1206,N_1584);
xor U1892 (N_1892,N_1295,N_1293);
nand U1893 (N_1893,N_1578,N_1463);
and U1894 (N_1894,N_1396,N_1597);
nor U1895 (N_1895,N_1482,N_1573);
and U1896 (N_1896,N_1318,N_1204);
xnor U1897 (N_1897,N_1234,N_1228);
nand U1898 (N_1898,N_1227,N_1329);
nand U1899 (N_1899,N_1369,N_1348);
and U1900 (N_1900,N_1325,N_1215);
and U1901 (N_1901,N_1369,N_1450);
and U1902 (N_1902,N_1542,N_1437);
nand U1903 (N_1903,N_1350,N_1295);
or U1904 (N_1904,N_1398,N_1592);
or U1905 (N_1905,N_1552,N_1216);
or U1906 (N_1906,N_1441,N_1205);
nand U1907 (N_1907,N_1285,N_1471);
or U1908 (N_1908,N_1296,N_1258);
nand U1909 (N_1909,N_1342,N_1577);
and U1910 (N_1910,N_1362,N_1548);
or U1911 (N_1911,N_1515,N_1482);
or U1912 (N_1912,N_1252,N_1483);
and U1913 (N_1913,N_1381,N_1391);
nor U1914 (N_1914,N_1245,N_1251);
and U1915 (N_1915,N_1433,N_1333);
nand U1916 (N_1916,N_1316,N_1229);
and U1917 (N_1917,N_1397,N_1598);
and U1918 (N_1918,N_1380,N_1528);
or U1919 (N_1919,N_1275,N_1221);
xor U1920 (N_1920,N_1437,N_1303);
nand U1921 (N_1921,N_1290,N_1345);
and U1922 (N_1922,N_1341,N_1258);
nand U1923 (N_1923,N_1442,N_1489);
and U1924 (N_1924,N_1514,N_1569);
or U1925 (N_1925,N_1345,N_1439);
and U1926 (N_1926,N_1514,N_1449);
xnor U1927 (N_1927,N_1234,N_1311);
or U1928 (N_1928,N_1508,N_1284);
or U1929 (N_1929,N_1344,N_1405);
and U1930 (N_1930,N_1406,N_1505);
nand U1931 (N_1931,N_1330,N_1253);
nor U1932 (N_1932,N_1293,N_1406);
and U1933 (N_1933,N_1454,N_1493);
nor U1934 (N_1934,N_1278,N_1276);
and U1935 (N_1935,N_1455,N_1321);
or U1936 (N_1936,N_1598,N_1388);
or U1937 (N_1937,N_1538,N_1380);
and U1938 (N_1938,N_1362,N_1373);
nand U1939 (N_1939,N_1391,N_1378);
nand U1940 (N_1940,N_1505,N_1434);
nor U1941 (N_1941,N_1471,N_1286);
nor U1942 (N_1942,N_1466,N_1569);
and U1943 (N_1943,N_1495,N_1524);
or U1944 (N_1944,N_1221,N_1323);
xor U1945 (N_1945,N_1268,N_1514);
nand U1946 (N_1946,N_1571,N_1577);
and U1947 (N_1947,N_1302,N_1255);
nor U1948 (N_1948,N_1486,N_1234);
nand U1949 (N_1949,N_1487,N_1380);
nand U1950 (N_1950,N_1526,N_1475);
xnor U1951 (N_1951,N_1526,N_1506);
nand U1952 (N_1952,N_1501,N_1246);
nand U1953 (N_1953,N_1200,N_1403);
nor U1954 (N_1954,N_1297,N_1495);
nor U1955 (N_1955,N_1437,N_1363);
or U1956 (N_1956,N_1362,N_1411);
nand U1957 (N_1957,N_1506,N_1383);
and U1958 (N_1958,N_1300,N_1222);
nor U1959 (N_1959,N_1297,N_1368);
or U1960 (N_1960,N_1388,N_1212);
or U1961 (N_1961,N_1475,N_1319);
and U1962 (N_1962,N_1350,N_1294);
xnor U1963 (N_1963,N_1568,N_1451);
xor U1964 (N_1964,N_1276,N_1415);
and U1965 (N_1965,N_1370,N_1554);
or U1966 (N_1966,N_1360,N_1201);
nor U1967 (N_1967,N_1537,N_1259);
xor U1968 (N_1968,N_1241,N_1237);
and U1969 (N_1969,N_1588,N_1324);
nor U1970 (N_1970,N_1224,N_1252);
and U1971 (N_1971,N_1206,N_1202);
and U1972 (N_1972,N_1273,N_1481);
nor U1973 (N_1973,N_1215,N_1274);
nor U1974 (N_1974,N_1477,N_1292);
nor U1975 (N_1975,N_1470,N_1220);
nor U1976 (N_1976,N_1430,N_1309);
or U1977 (N_1977,N_1492,N_1527);
and U1978 (N_1978,N_1547,N_1328);
nor U1979 (N_1979,N_1573,N_1463);
or U1980 (N_1980,N_1593,N_1200);
xnor U1981 (N_1981,N_1520,N_1276);
nor U1982 (N_1982,N_1379,N_1492);
or U1983 (N_1983,N_1533,N_1413);
xnor U1984 (N_1984,N_1412,N_1470);
or U1985 (N_1985,N_1341,N_1290);
xor U1986 (N_1986,N_1599,N_1211);
nand U1987 (N_1987,N_1291,N_1337);
or U1988 (N_1988,N_1281,N_1556);
nand U1989 (N_1989,N_1274,N_1286);
and U1990 (N_1990,N_1545,N_1291);
or U1991 (N_1991,N_1227,N_1590);
xor U1992 (N_1992,N_1392,N_1263);
xor U1993 (N_1993,N_1279,N_1463);
xor U1994 (N_1994,N_1515,N_1303);
nor U1995 (N_1995,N_1323,N_1509);
nor U1996 (N_1996,N_1302,N_1303);
xor U1997 (N_1997,N_1491,N_1315);
or U1998 (N_1998,N_1409,N_1324);
and U1999 (N_1999,N_1434,N_1221);
nand U2000 (N_2000,N_1900,N_1918);
nor U2001 (N_2001,N_1788,N_1831);
or U2002 (N_2002,N_1655,N_1733);
xnor U2003 (N_2003,N_1698,N_1896);
or U2004 (N_2004,N_1968,N_1928);
nor U2005 (N_2005,N_1726,N_1889);
nand U2006 (N_2006,N_1837,N_1632);
xnor U2007 (N_2007,N_1700,N_1704);
and U2008 (N_2008,N_1670,N_1775);
nand U2009 (N_2009,N_1600,N_1662);
and U2010 (N_2010,N_1610,N_1876);
nand U2011 (N_2011,N_1980,N_1944);
xnor U2012 (N_2012,N_1695,N_1903);
nor U2013 (N_2013,N_1699,N_1617);
or U2014 (N_2014,N_1664,N_1798);
nor U2015 (N_2015,N_1741,N_1866);
and U2016 (N_2016,N_1636,N_1743);
xnor U2017 (N_2017,N_1826,N_1608);
xnor U2018 (N_2018,N_1772,N_1683);
nor U2019 (N_2019,N_1795,N_1823);
and U2020 (N_2020,N_1891,N_1828);
xor U2021 (N_2021,N_1941,N_1945);
xnor U2022 (N_2022,N_1899,N_1997);
nor U2023 (N_2023,N_1692,N_1785);
and U2024 (N_2024,N_1760,N_1719);
nand U2025 (N_2025,N_1784,N_1971);
and U2026 (N_2026,N_1649,N_1761);
xnor U2027 (N_2027,N_1663,N_1897);
xor U2028 (N_2028,N_1961,N_1815);
nor U2029 (N_2029,N_1863,N_1865);
and U2030 (N_2030,N_1697,N_1856);
nor U2031 (N_2031,N_1979,N_1782);
xnor U2032 (N_2032,N_1757,N_1773);
nor U2033 (N_2033,N_1985,N_1710);
xnor U2034 (N_2034,N_1882,N_1931);
or U2035 (N_2035,N_1749,N_1770);
xor U2036 (N_2036,N_1615,N_1998);
nand U2037 (N_2037,N_1845,N_1652);
or U2038 (N_2038,N_1807,N_1768);
or U2039 (N_2039,N_1675,N_1701);
nand U2040 (N_2040,N_1707,N_1929);
and U2041 (N_2041,N_1799,N_1680);
xnor U2042 (N_2042,N_1694,N_1739);
nand U2043 (N_2043,N_1748,N_1960);
nand U2044 (N_2044,N_1672,N_1629);
xor U2045 (N_2045,N_1814,N_1917);
nor U2046 (N_2046,N_1752,N_1919);
xor U2047 (N_2047,N_1852,N_1989);
nand U2048 (N_2048,N_1651,N_1999);
xor U2049 (N_2049,N_1661,N_1860);
or U2050 (N_2050,N_1958,N_1601);
nand U2051 (N_2051,N_1786,N_1671);
and U2052 (N_2052,N_1921,N_1902);
nand U2053 (N_2053,N_1875,N_1774);
and U2054 (N_2054,N_1614,N_1650);
and U2055 (N_2055,N_1794,N_1718);
nand U2056 (N_2056,N_1816,N_1677);
or U2057 (N_2057,N_1853,N_1943);
or U2058 (N_2058,N_1656,N_1744);
and U2059 (N_2059,N_1708,N_1643);
and U2060 (N_2060,N_1705,N_1981);
nor U2061 (N_2061,N_1877,N_1764);
or U2062 (N_2062,N_1604,N_1809);
and U2063 (N_2063,N_1793,N_1893);
or U2064 (N_2064,N_1910,N_1642);
and U2065 (N_2065,N_1612,N_1874);
or U2066 (N_2066,N_1754,N_1800);
xor U2067 (N_2067,N_1727,N_1712);
xnor U2068 (N_2068,N_1844,N_1940);
nand U2069 (N_2069,N_1690,N_1916);
or U2070 (N_2070,N_1962,N_1953);
nand U2071 (N_2071,N_1992,N_1647);
or U2072 (N_2072,N_1638,N_1869);
or U2073 (N_2073,N_1603,N_1635);
or U2074 (N_2074,N_1821,N_1850);
xor U2075 (N_2075,N_1818,N_1973);
xor U2076 (N_2076,N_1802,N_1616);
or U2077 (N_2077,N_1849,N_1624);
xor U2078 (N_2078,N_1644,N_1938);
or U2079 (N_2079,N_1970,N_1817);
or U2080 (N_2080,N_1666,N_1711);
nor U2081 (N_2081,N_1868,N_1822);
nand U2082 (N_2082,N_1731,N_1829);
or U2083 (N_2083,N_1637,N_1976);
nor U2084 (N_2084,N_1605,N_1892);
and U2085 (N_2085,N_1618,N_1932);
nor U2086 (N_2086,N_1621,N_1687);
xnor U2087 (N_2087,N_1625,N_1842);
xnor U2088 (N_2088,N_1676,N_1854);
and U2089 (N_2089,N_1791,N_1833);
or U2090 (N_2090,N_1847,N_1789);
nor U2091 (N_2091,N_1862,N_1703);
nand U2092 (N_2092,N_1622,N_1740);
xor U2093 (N_2093,N_1763,N_1846);
nor U2094 (N_2094,N_1606,N_1836);
or U2095 (N_2095,N_1732,N_1950);
and U2096 (N_2096,N_1735,N_1648);
or U2097 (N_2097,N_1839,N_1769);
nor U2098 (N_2098,N_1668,N_1657);
nor U2099 (N_2099,N_1631,N_1885);
or U2100 (N_2100,N_1665,N_1646);
nand U2101 (N_2101,N_1915,N_1872);
and U2102 (N_2102,N_1939,N_1923);
and U2103 (N_2103,N_1859,N_1991);
nand U2104 (N_2104,N_1830,N_1767);
xor U2105 (N_2105,N_1654,N_1925);
and U2106 (N_2106,N_1906,N_1963);
nor U2107 (N_2107,N_1688,N_1952);
nor U2108 (N_2108,N_1641,N_1790);
or U2109 (N_2109,N_1954,N_1972);
or U2110 (N_2110,N_1681,N_1895);
nand U2111 (N_2111,N_1905,N_1684);
xor U2112 (N_2112,N_1888,N_1721);
nor U2113 (N_2113,N_1607,N_1913);
nor U2114 (N_2114,N_1645,N_1619);
or U2115 (N_2115,N_1682,N_1955);
or U2116 (N_2116,N_1620,N_1977);
and U2117 (N_2117,N_1717,N_1949);
nor U2118 (N_2118,N_1870,N_1734);
xor U2119 (N_2119,N_1861,N_1667);
and U2120 (N_2120,N_1602,N_1990);
nand U2121 (N_2121,N_1777,N_1627);
and U2122 (N_2122,N_1723,N_1937);
and U2123 (N_2123,N_1765,N_1674);
and U2124 (N_2124,N_1766,N_1956);
nand U2125 (N_2125,N_1908,N_1779);
xor U2126 (N_2126,N_1696,N_1959);
nand U2127 (N_2127,N_1867,N_1927);
nand U2128 (N_2128,N_1611,N_1737);
and U2129 (N_2129,N_1805,N_1801);
and U2130 (N_2130,N_1673,N_1806);
nor U2131 (N_2131,N_1901,N_1843);
nand U2132 (N_2132,N_1912,N_1738);
and U2133 (N_2133,N_1781,N_1640);
nor U2134 (N_2134,N_1907,N_1909);
nor U2135 (N_2135,N_1841,N_1827);
nand U2136 (N_2136,N_1848,N_1883);
xnor U2137 (N_2137,N_1878,N_1988);
or U2138 (N_2138,N_1825,N_1948);
and U2139 (N_2139,N_1851,N_1678);
or U2140 (N_2140,N_1904,N_1762);
or U2141 (N_2141,N_1759,N_1804);
and U2142 (N_2142,N_1924,N_1969);
nand U2143 (N_2143,N_1886,N_1630);
nand U2144 (N_2144,N_1634,N_1623);
and U2145 (N_2145,N_1855,N_1780);
and U2146 (N_2146,N_1982,N_1736);
xor U2147 (N_2147,N_1691,N_1722);
xor U2148 (N_2148,N_1942,N_1838);
nor U2149 (N_2149,N_1808,N_1986);
xor U2150 (N_2150,N_1810,N_1713);
and U2151 (N_2151,N_1898,N_1751);
xor U2152 (N_2152,N_1946,N_1796);
xor U2153 (N_2153,N_1922,N_1813);
and U2154 (N_2154,N_1840,N_1613);
nand U2155 (N_2155,N_1720,N_1714);
nor U2156 (N_2156,N_1884,N_1819);
and U2157 (N_2157,N_1964,N_1935);
or U2158 (N_2158,N_1725,N_1715);
and U2159 (N_2159,N_1706,N_1887);
xnor U2160 (N_2160,N_1993,N_1832);
and U2161 (N_2161,N_1994,N_1873);
nor U2162 (N_2162,N_1864,N_1936);
or U2163 (N_2163,N_1753,N_1659);
nand U2164 (N_2164,N_1881,N_1716);
nor U2165 (N_2165,N_1746,N_1756);
or U2166 (N_2166,N_1724,N_1783);
nor U2167 (N_2167,N_1965,N_1686);
xor U2168 (N_2168,N_1778,N_1633);
nand U2169 (N_2169,N_1658,N_1983);
xor U2170 (N_2170,N_1811,N_1995);
nor U2171 (N_2171,N_1880,N_1975);
nand U2172 (N_2172,N_1934,N_1679);
and U2173 (N_2173,N_1812,N_1626);
xor U2174 (N_2174,N_1660,N_1920);
and U2175 (N_2175,N_1787,N_1628);
and U2176 (N_2176,N_1951,N_1835);
nor U2177 (N_2177,N_1967,N_1792);
nor U2178 (N_2178,N_1978,N_1930);
nor U2179 (N_2179,N_1747,N_1974);
or U2180 (N_2180,N_1776,N_1797);
or U2181 (N_2181,N_1984,N_1996);
and U2182 (N_2182,N_1669,N_1689);
xnor U2183 (N_2183,N_1987,N_1685);
and U2184 (N_2184,N_1894,N_1858);
nor U2185 (N_2185,N_1824,N_1933);
or U2186 (N_2186,N_1745,N_1914);
and U2187 (N_2187,N_1890,N_1803);
and U2188 (N_2188,N_1834,N_1639);
xnor U2189 (N_2189,N_1730,N_1755);
or U2190 (N_2190,N_1728,N_1966);
and U2191 (N_2191,N_1693,N_1709);
xor U2192 (N_2192,N_1729,N_1871);
and U2193 (N_2193,N_1702,N_1857);
or U2194 (N_2194,N_1653,N_1742);
nor U2195 (N_2195,N_1609,N_1771);
xnor U2196 (N_2196,N_1957,N_1926);
nand U2197 (N_2197,N_1820,N_1879);
nand U2198 (N_2198,N_1947,N_1758);
xor U2199 (N_2199,N_1911,N_1750);
and U2200 (N_2200,N_1792,N_1776);
nor U2201 (N_2201,N_1892,N_1756);
nand U2202 (N_2202,N_1993,N_1715);
nand U2203 (N_2203,N_1741,N_1835);
nor U2204 (N_2204,N_1749,N_1634);
nand U2205 (N_2205,N_1671,N_1987);
xnor U2206 (N_2206,N_1677,N_1624);
nand U2207 (N_2207,N_1985,N_1845);
or U2208 (N_2208,N_1719,N_1952);
nor U2209 (N_2209,N_1827,N_1749);
or U2210 (N_2210,N_1687,N_1960);
or U2211 (N_2211,N_1794,N_1642);
and U2212 (N_2212,N_1981,N_1940);
xor U2213 (N_2213,N_1617,N_1745);
and U2214 (N_2214,N_1714,N_1918);
nand U2215 (N_2215,N_1727,N_1817);
xor U2216 (N_2216,N_1856,N_1706);
xor U2217 (N_2217,N_1863,N_1682);
and U2218 (N_2218,N_1703,N_1606);
or U2219 (N_2219,N_1753,N_1979);
nand U2220 (N_2220,N_1634,N_1900);
xnor U2221 (N_2221,N_1719,N_1917);
or U2222 (N_2222,N_1878,N_1919);
nor U2223 (N_2223,N_1961,N_1709);
and U2224 (N_2224,N_1676,N_1936);
xnor U2225 (N_2225,N_1764,N_1754);
nor U2226 (N_2226,N_1671,N_1779);
xnor U2227 (N_2227,N_1796,N_1944);
nor U2228 (N_2228,N_1735,N_1687);
or U2229 (N_2229,N_1858,N_1978);
nand U2230 (N_2230,N_1726,N_1850);
nand U2231 (N_2231,N_1649,N_1646);
xnor U2232 (N_2232,N_1634,N_1602);
nand U2233 (N_2233,N_1823,N_1831);
nand U2234 (N_2234,N_1733,N_1783);
nand U2235 (N_2235,N_1799,N_1705);
xor U2236 (N_2236,N_1625,N_1996);
xor U2237 (N_2237,N_1738,N_1866);
and U2238 (N_2238,N_1700,N_1796);
xor U2239 (N_2239,N_1766,N_1686);
xnor U2240 (N_2240,N_1994,N_1978);
and U2241 (N_2241,N_1993,N_1655);
xor U2242 (N_2242,N_1708,N_1681);
or U2243 (N_2243,N_1843,N_1873);
or U2244 (N_2244,N_1777,N_1973);
nor U2245 (N_2245,N_1692,N_1914);
or U2246 (N_2246,N_1636,N_1759);
or U2247 (N_2247,N_1746,N_1892);
or U2248 (N_2248,N_1790,N_1748);
or U2249 (N_2249,N_1615,N_1693);
nand U2250 (N_2250,N_1829,N_1724);
nand U2251 (N_2251,N_1619,N_1940);
nand U2252 (N_2252,N_1647,N_1613);
xnor U2253 (N_2253,N_1986,N_1870);
or U2254 (N_2254,N_1703,N_1861);
nor U2255 (N_2255,N_1823,N_1833);
or U2256 (N_2256,N_1665,N_1752);
xor U2257 (N_2257,N_1660,N_1767);
nor U2258 (N_2258,N_1638,N_1677);
nor U2259 (N_2259,N_1677,N_1956);
or U2260 (N_2260,N_1707,N_1979);
xor U2261 (N_2261,N_1692,N_1836);
or U2262 (N_2262,N_1657,N_1865);
nand U2263 (N_2263,N_1982,N_1987);
nand U2264 (N_2264,N_1897,N_1972);
nand U2265 (N_2265,N_1826,N_1668);
or U2266 (N_2266,N_1944,N_1627);
or U2267 (N_2267,N_1815,N_1628);
or U2268 (N_2268,N_1691,N_1686);
xnor U2269 (N_2269,N_1831,N_1944);
nor U2270 (N_2270,N_1676,N_1701);
and U2271 (N_2271,N_1927,N_1880);
and U2272 (N_2272,N_1607,N_1793);
nor U2273 (N_2273,N_1794,N_1915);
or U2274 (N_2274,N_1960,N_1840);
nor U2275 (N_2275,N_1750,N_1678);
and U2276 (N_2276,N_1947,N_1787);
or U2277 (N_2277,N_1744,N_1719);
and U2278 (N_2278,N_1841,N_1723);
nand U2279 (N_2279,N_1617,N_1899);
or U2280 (N_2280,N_1700,N_1894);
xor U2281 (N_2281,N_1795,N_1620);
nand U2282 (N_2282,N_1821,N_1643);
xnor U2283 (N_2283,N_1636,N_1706);
and U2284 (N_2284,N_1992,N_1782);
nand U2285 (N_2285,N_1770,N_1842);
nor U2286 (N_2286,N_1817,N_1785);
nand U2287 (N_2287,N_1858,N_1708);
or U2288 (N_2288,N_1721,N_1666);
or U2289 (N_2289,N_1946,N_1888);
nor U2290 (N_2290,N_1957,N_1726);
and U2291 (N_2291,N_1823,N_1976);
or U2292 (N_2292,N_1954,N_1673);
xor U2293 (N_2293,N_1905,N_1823);
and U2294 (N_2294,N_1617,N_1784);
xnor U2295 (N_2295,N_1967,N_1769);
nor U2296 (N_2296,N_1753,N_1631);
xnor U2297 (N_2297,N_1720,N_1775);
nand U2298 (N_2298,N_1742,N_1778);
xnor U2299 (N_2299,N_1647,N_1786);
or U2300 (N_2300,N_1760,N_1941);
nand U2301 (N_2301,N_1605,N_1843);
or U2302 (N_2302,N_1616,N_1976);
and U2303 (N_2303,N_1639,N_1867);
nor U2304 (N_2304,N_1697,N_1627);
or U2305 (N_2305,N_1989,N_1620);
or U2306 (N_2306,N_1875,N_1855);
and U2307 (N_2307,N_1682,N_1606);
or U2308 (N_2308,N_1968,N_1890);
and U2309 (N_2309,N_1709,N_1881);
and U2310 (N_2310,N_1934,N_1962);
nand U2311 (N_2311,N_1671,N_1711);
nor U2312 (N_2312,N_1816,N_1872);
nor U2313 (N_2313,N_1960,N_1957);
xor U2314 (N_2314,N_1745,N_1835);
nor U2315 (N_2315,N_1617,N_1607);
xor U2316 (N_2316,N_1615,N_1903);
xnor U2317 (N_2317,N_1972,N_1931);
and U2318 (N_2318,N_1963,N_1866);
nand U2319 (N_2319,N_1933,N_1714);
nand U2320 (N_2320,N_1737,N_1968);
nor U2321 (N_2321,N_1926,N_1801);
and U2322 (N_2322,N_1801,N_1997);
nor U2323 (N_2323,N_1979,N_1909);
nand U2324 (N_2324,N_1881,N_1677);
or U2325 (N_2325,N_1916,N_1748);
and U2326 (N_2326,N_1628,N_1667);
nor U2327 (N_2327,N_1601,N_1803);
xnor U2328 (N_2328,N_1975,N_1973);
xor U2329 (N_2329,N_1817,N_1923);
and U2330 (N_2330,N_1826,N_1946);
nand U2331 (N_2331,N_1915,N_1783);
or U2332 (N_2332,N_1729,N_1703);
and U2333 (N_2333,N_1904,N_1853);
nor U2334 (N_2334,N_1883,N_1773);
xor U2335 (N_2335,N_1975,N_1845);
nand U2336 (N_2336,N_1696,N_1838);
and U2337 (N_2337,N_1953,N_1820);
and U2338 (N_2338,N_1958,N_1603);
nor U2339 (N_2339,N_1704,N_1874);
xor U2340 (N_2340,N_1840,N_1796);
and U2341 (N_2341,N_1966,N_1862);
xor U2342 (N_2342,N_1826,N_1733);
xnor U2343 (N_2343,N_1747,N_1965);
nand U2344 (N_2344,N_1655,N_1709);
nand U2345 (N_2345,N_1651,N_1798);
nor U2346 (N_2346,N_1962,N_1909);
nor U2347 (N_2347,N_1774,N_1964);
or U2348 (N_2348,N_1630,N_1640);
and U2349 (N_2349,N_1703,N_1833);
and U2350 (N_2350,N_1809,N_1926);
nor U2351 (N_2351,N_1729,N_1726);
nor U2352 (N_2352,N_1836,N_1653);
and U2353 (N_2353,N_1729,N_1995);
nand U2354 (N_2354,N_1709,N_1818);
nand U2355 (N_2355,N_1686,N_1928);
nor U2356 (N_2356,N_1856,N_1728);
nand U2357 (N_2357,N_1959,N_1977);
nand U2358 (N_2358,N_1786,N_1971);
or U2359 (N_2359,N_1767,N_1945);
nor U2360 (N_2360,N_1653,N_1773);
xor U2361 (N_2361,N_1879,N_1749);
xnor U2362 (N_2362,N_1855,N_1664);
or U2363 (N_2363,N_1771,N_1696);
or U2364 (N_2364,N_1727,N_1606);
or U2365 (N_2365,N_1748,N_1803);
nor U2366 (N_2366,N_1849,N_1916);
xor U2367 (N_2367,N_1786,N_1698);
and U2368 (N_2368,N_1609,N_1770);
nand U2369 (N_2369,N_1625,N_1712);
nor U2370 (N_2370,N_1851,N_1761);
nand U2371 (N_2371,N_1645,N_1628);
nor U2372 (N_2372,N_1875,N_1843);
and U2373 (N_2373,N_1748,N_1853);
and U2374 (N_2374,N_1804,N_1737);
or U2375 (N_2375,N_1755,N_1702);
and U2376 (N_2376,N_1974,N_1911);
nand U2377 (N_2377,N_1898,N_1780);
nand U2378 (N_2378,N_1853,N_1966);
nor U2379 (N_2379,N_1944,N_1802);
and U2380 (N_2380,N_1694,N_1742);
and U2381 (N_2381,N_1643,N_1685);
and U2382 (N_2382,N_1788,N_1846);
or U2383 (N_2383,N_1769,N_1957);
nand U2384 (N_2384,N_1890,N_1957);
xnor U2385 (N_2385,N_1872,N_1732);
xnor U2386 (N_2386,N_1703,N_1832);
xnor U2387 (N_2387,N_1830,N_1661);
nor U2388 (N_2388,N_1756,N_1783);
or U2389 (N_2389,N_1746,N_1814);
nor U2390 (N_2390,N_1662,N_1800);
xor U2391 (N_2391,N_1986,N_1695);
xnor U2392 (N_2392,N_1870,N_1980);
or U2393 (N_2393,N_1668,N_1710);
nor U2394 (N_2394,N_1922,N_1717);
xor U2395 (N_2395,N_1638,N_1620);
nor U2396 (N_2396,N_1958,N_1716);
nor U2397 (N_2397,N_1705,N_1810);
xor U2398 (N_2398,N_1956,N_1792);
nand U2399 (N_2399,N_1624,N_1658);
nor U2400 (N_2400,N_2126,N_2071);
xor U2401 (N_2401,N_2103,N_2381);
nor U2402 (N_2402,N_2356,N_2233);
and U2403 (N_2403,N_2241,N_2360);
nand U2404 (N_2404,N_2127,N_2211);
xor U2405 (N_2405,N_2017,N_2387);
or U2406 (N_2406,N_2033,N_2083);
nand U2407 (N_2407,N_2161,N_2191);
and U2408 (N_2408,N_2332,N_2020);
nand U2409 (N_2409,N_2198,N_2039);
and U2410 (N_2410,N_2263,N_2031);
or U2411 (N_2411,N_2340,N_2245);
nor U2412 (N_2412,N_2056,N_2388);
nand U2413 (N_2413,N_2058,N_2094);
nand U2414 (N_2414,N_2212,N_2029);
nand U2415 (N_2415,N_2073,N_2293);
and U2416 (N_2416,N_2288,N_2396);
and U2417 (N_2417,N_2311,N_2266);
nand U2418 (N_2418,N_2345,N_2243);
nor U2419 (N_2419,N_2256,N_2213);
and U2420 (N_2420,N_2069,N_2346);
and U2421 (N_2421,N_2242,N_2115);
or U2422 (N_2422,N_2010,N_2085);
nor U2423 (N_2423,N_2199,N_2268);
and U2424 (N_2424,N_2232,N_2244);
nor U2425 (N_2425,N_2361,N_2038);
and U2426 (N_2426,N_2362,N_2118);
xor U2427 (N_2427,N_2062,N_2076);
nand U2428 (N_2428,N_2261,N_2027);
nor U2429 (N_2429,N_2229,N_2008);
and U2430 (N_2430,N_2303,N_2307);
xnor U2431 (N_2431,N_2373,N_2299);
xor U2432 (N_2432,N_2300,N_2078);
nand U2433 (N_2433,N_2391,N_2182);
xor U2434 (N_2434,N_2220,N_2023);
xor U2435 (N_2435,N_2044,N_2190);
nand U2436 (N_2436,N_2389,N_2231);
or U2437 (N_2437,N_2317,N_2137);
nor U2438 (N_2438,N_2016,N_2223);
or U2439 (N_2439,N_2368,N_2336);
nand U2440 (N_2440,N_2239,N_2065);
or U2441 (N_2441,N_2128,N_2301);
nor U2442 (N_2442,N_2072,N_2376);
nor U2443 (N_2443,N_2117,N_2070);
and U2444 (N_2444,N_2207,N_2259);
nand U2445 (N_2445,N_2315,N_2159);
and U2446 (N_2446,N_2377,N_2155);
nand U2447 (N_2447,N_2393,N_2250);
nor U2448 (N_2448,N_2153,N_2310);
or U2449 (N_2449,N_2102,N_2348);
nor U2450 (N_2450,N_2059,N_2166);
nor U2451 (N_2451,N_2347,N_2181);
or U2452 (N_2452,N_2079,N_2095);
xnor U2453 (N_2453,N_2113,N_2122);
nand U2454 (N_2454,N_2157,N_2134);
nor U2455 (N_2455,N_2353,N_2382);
nor U2456 (N_2456,N_2035,N_2004);
xor U2457 (N_2457,N_2052,N_2331);
xor U2458 (N_2458,N_2110,N_2168);
and U2459 (N_2459,N_2338,N_2247);
xor U2460 (N_2460,N_2025,N_2274);
and U2461 (N_2461,N_2218,N_2097);
xnor U2462 (N_2462,N_2143,N_2375);
nor U2463 (N_2463,N_2148,N_2398);
xnor U2464 (N_2464,N_2173,N_2125);
or U2465 (N_2465,N_2142,N_2321);
or U2466 (N_2466,N_2172,N_2390);
nor U2467 (N_2467,N_2319,N_2325);
nand U2468 (N_2468,N_2219,N_2013);
nand U2469 (N_2469,N_2209,N_2099);
xor U2470 (N_2470,N_2129,N_2253);
nand U2471 (N_2471,N_2341,N_2032);
and U2472 (N_2472,N_2189,N_2342);
nand U2473 (N_2473,N_2357,N_2162);
nand U2474 (N_2474,N_2320,N_2399);
nor U2475 (N_2475,N_2318,N_2369);
nand U2476 (N_2476,N_2251,N_2109);
or U2477 (N_2477,N_2187,N_2074);
xnor U2478 (N_2478,N_2176,N_2184);
and U2479 (N_2479,N_2350,N_2053);
nand U2480 (N_2480,N_2291,N_2230);
and U2481 (N_2481,N_2177,N_2269);
and U2482 (N_2482,N_2111,N_2091);
and U2483 (N_2483,N_2383,N_2283);
xor U2484 (N_2484,N_2343,N_2135);
nand U2485 (N_2485,N_2281,N_2297);
and U2486 (N_2486,N_2011,N_2280);
and U2487 (N_2487,N_2121,N_2260);
and U2488 (N_2488,N_2395,N_2224);
or U2489 (N_2489,N_2156,N_2370);
nor U2490 (N_2490,N_2141,N_2374);
and U2491 (N_2491,N_2067,N_2202);
or U2492 (N_2492,N_2064,N_2276);
nand U2493 (N_2493,N_2208,N_2354);
xnor U2494 (N_2494,N_2167,N_2150);
or U2495 (N_2495,N_2270,N_2175);
nand U2496 (N_2496,N_2132,N_2235);
nand U2497 (N_2497,N_2015,N_2312);
xor U2498 (N_2498,N_2019,N_2334);
xnor U2499 (N_2499,N_2145,N_2386);
nand U2500 (N_2500,N_2131,N_2041);
or U2501 (N_2501,N_2306,N_2363);
or U2502 (N_2502,N_2042,N_2192);
nor U2503 (N_2503,N_2367,N_2246);
or U2504 (N_2504,N_2215,N_2164);
nor U2505 (N_2505,N_2170,N_2080);
nand U2506 (N_2506,N_2014,N_2339);
or U2507 (N_2507,N_2214,N_2180);
and U2508 (N_2508,N_2105,N_2359);
or U2509 (N_2509,N_2206,N_2018);
nor U2510 (N_2510,N_2292,N_2249);
and U2511 (N_2511,N_2258,N_2050);
nor U2512 (N_2512,N_2328,N_2380);
nor U2513 (N_2513,N_2036,N_2098);
or U2514 (N_2514,N_2136,N_2275);
nor U2515 (N_2515,N_2308,N_2290);
nand U2516 (N_2516,N_2333,N_2397);
and U2517 (N_2517,N_2324,N_2257);
or U2518 (N_2518,N_2364,N_2335);
nor U2519 (N_2519,N_2101,N_2195);
xor U2520 (N_2520,N_2355,N_2327);
and U2521 (N_2521,N_2267,N_2197);
xnor U2522 (N_2522,N_2394,N_2048);
nor U2523 (N_2523,N_2221,N_2055);
nor U2524 (N_2524,N_2273,N_2084);
nor U2525 (N_2525,N_2179,N_2282);
xor U2526 (N_2526,N_2082,N_2133);
and U2527 (N_2527,N_2045,N_2194);
and U2528 (N_2528,N_2089,N_2130);
or U2529 (N_2529,N_2146,N_2112);
and U2530 (N_2530,N_2200,N_2144);
nor U2531 (N_2531,N_2061,N_2123);
or U2532 (N_2532,N_2185,N_2271);
or U2533 (N_2533,N_2330,N_2088);
xnor U2534 (N_2534,N_2349,N_2304);
and U2535 (N_2535,N_2188,N_2205);
or U2536 (N_2536,N_2222,N_2240);
xnor U2537 (N_2537,N_2314,N_2138);
nand U2538 (N_2538,N_2277,N_2124);
xor U2539 (N_2539,N_2051,N_2272);
and U2540 (N_2540,N_2228,N_2178);
nor U2541 (N_2541,N_2237,N_2116);
xnor U2542 (N_2542,N_2385,N_2068);
and U2543 (N_2543,N_2003,N_2234);
or U2544 (N_2544,N_2337,N_2057);
nand U2545 (N_2545,N_2286,N_2236);
and U2546 (N_2546,N_2047,N_2030);
nor U2547 (N_2547,N_2040,N_2028);
nand U2548 (N_2548,N_2002,N_2392);
and U2549 (N_2549,N_2075,N_2278);
or U2550 (N_2550,N_2007,N_2226);
and U2551 (N_2551,N_2108,N_2217);
nor U2552 (N_2552,N_2298,N_2165);
nand U2553 (N_2553,N_2227,N_2024);
or U2554 (N_2554,N_2092,N_2366);
and U2555 (N_2555,N_2284,N_2066);
nor U2556 (N_2556,N_2140,N_2210);
and U2557 (N_2557,N_2037,N_2305);
nor U2558 (N_2558,N_2279,N_2021);
xnor U2559 (N_2559,N_2201,N_2351);
nand U2560 (N_2560,N_2326,N_2034);
nor U2561 (N_2561,N_2225,N_2255);
xor U2562 (N_2562,N_2171,N_2186);
nand U2563 (N_2563,N_2009,N_2285);
or U2564 (N_2564,N_2077,N_2158);
or U2565 (N_2565,N_2294,N_2196);
xnor U2566 (N_2566,N_2005,N_2254);
nand U2567 (N_2567,N_2203,N_2262);
or U2568 (N_2568,N_2365,N_2006);
xor U2569 (N_2569,N_2372,N_2302);
xor U2570 (N_2570,N_2169,N_2152);
or U2571 (N_2571,N_2090,N_2096);
and U2572 (N_2572,N_2163,N_2043);
xor U2573 (N_2573,N_2344,N_2026);
or U2574 (N_2574,N_2193,N_2087);
nand U2575 (N_2575,N_2114,N_2296);
xor U2576 (N_2576,N_2379,N_2160);
and U2577 (N_2577,N_2216,N_2384);
nor U2578 (N_2578,N_2049,N_2120);
or U2579 (N_2579,N_2264,N_2093);
nor U2580 (N_2580,N_2238,N_2139);
nor U2581 (N_2581,N_2289,N_2378);
and U2582 (N_2582,N_2104,N_2358);
nand U2583 (N_2583,N_2316,N_2371);
and U2584 (N_2584,N_2119,N_2046);
nand U2585 (N_2585,N_2323,N_2309);
xnor U2586 (N_2586,N_2174,N_2265);
or U2587 (N_2587,N_2149,N_2000);
xor U2588 (N_2588,N_2322,N_2204);
xnor U2589 (N_2589,N_2151,N_2107);
nand U2590 (N_2590,N_2012,N_2313);
xor U2591 (N_2591,N_2154,N_2063);
and U2592 (N_2592,N_2081,N_2106);
nand U2593 (N_2593,N_2329,N_2054);
xor U2594 (N_2594,N_2001,N_2183);
nand U2595 (N_2595,N_2060,N_2252);
nor U2596 (N_2596,N_2248,N_2086);
nor U2597 (N_2597,N_2295,N_2100);
and U2598 (N_2598,N_2287,N_2147);
or U2599 (N_2599,N_2352,N_2022);
and U2600 (N_2600,N_2342,N_2326);
nand U2601 (N_2601,N_2223,N_2140);
nand U2602 (N_2602,N_2081,N_2273);
nor U2603 (N_2603,N_2328,N_2381);
nor U2604 (N_2604,N_2012,N_2106);
and U2605 (N_2605,N_2176,N_2360);
nand U2606 (N_2606,N_2073,N_2275);
nand U2607 (N_2607,N_2029,N_2085);
or U2608 (N_2608,N_2388,N_2157);
and U2609 (N_2609,N_2023,N_2376);
and U2610 (N_2610,N_2110,N_2090);
xor U2611 (N_2611,N_2174,N_2003);
nand U2612 (N_2612,N_2025,N_2248);
nor U2613 (N_2613,N_2068,N_2354);
xor U2614 (N_2614,N_2208,N_2221);
xnor U2615 (N_2615,N_2022,N_2382);
nor U2616 (N_2616,N_2133,N_2038);
nor U2617 (N_2617,N_2273,N_2293);
nand U2618 (N_2618,N_2246,N_2034);
nor U2619 (N_2619,N_2142,N_2197);
nor U2620 (N_2620,N_2259,N_2215);
nor U2621 (N_2621,N_2274,N_2277);
and U2622 (N_2622,N_2211,N_2246);
or U2623 (N_2623,N_2357,N_2101);
nor U2624 (N_2624,N_2080,N_2112);
and U2625 (N_2625,N_2382,N_2385);
nor U2626 (N_2626,N_2075,N_2357);
or U2627 (N_2627,N_2202,N_2062);
xor U2628 (N_2628,N_2299,N_2086);
xor U2629 (N_2629,N_2271,N_2273);
xor U2630 (N_2630,N_2221,N_2215);
nor U2631 (N_2631,N_2102,N_2078);
nor U2632 (N_2632,N_2319,N_2276);
nor U2633 (N_2633,N_2022,N_2181);
and U2634 (N_2634,N_2154,N_2367);
xnor U2635 (N_2635,N_2040,N_2065);
xor U2636 (N_2636,N_2050,N_2343);
and U2637 (N_2637,N_2362,N_2165);
or U2638 (N_2638,N_2095,N_2307);
and U2639 (N_2639,N_2318,N_2121);
nor U2640 (N_2640,N_2364,N_2161);
or U2641 (N_2641,N_2060,N_2251);
and U2642 (N_2642,N_2067,N_2076);
nand U2643 (N_2643,N_2227,N_2297);
or U2644 (N_2644,N_2092,N_2026);
nor U2645 (N_2645,N_2392,N_2094);
nand U2646 (N_2646,N_2323,N_2322);
or U2647 (N_2647,N_2238,N_2090);
nor U2648 (N_2648,N_2106,N_2296);
or U2649 (N_2649,N_2388,N_2294);
nand U2650 (N_2650,N_2305,N_2134);
xnor U2651 (N_2651,N_2221,N_2282);
or U2652 (N_2652,N_2373,N_2347);
nand U2653 (N_2653,N_2103,N_2327);
nor U2654 (N_2654,N_2393,N_2239);
nor U2655 (N_2655,N_2220,N_2115);
xnor U2656 (N_2656,N_2287,N_2279);
nor U2657 (N_2657,N_2213,N_2278);
and U2658 (N_2658,N_2271,N_2028);
nand U2659 (N_2659,N_2288,N_2046);
xor U2660 (N_2660,N_2020,N_2310);
xor U2661 (N_2661,N_2363,N_2289);
or U2662 (N_2662,N_2209,N_2108);
or U2663 (N_2663,N_2269,N_2283);
xor U2664 (N_2664,N_2353,N_2338);
or U2665 (N_2665,N_2027,N_2011);
nor U2666 (N_2666,N_2036,N_2242);
nand U2667 (N_2667,N_2215,N_2055);
xnor U2668 (N_2668,N_2300,N_2297);
nor U2669 (N_2669,N_2262,N_2301);
or U2670 (N_2670,N_2248,N_2301);
nor U2671 (N_2671,N_2117,N_2103);
xnor U2672 (N_2672,N_2230,N_2319);
or U2673 (N_2673,N_2303,N_2224);
nor U2674 (N_2674,N_2377,N_2140);
xor U2675 (N_2675,N_2329,N_2137);
or U2676 (N_2676,N_2120,N_2057);
or U2677 (N_2677,N_2107,N_2179);
or U2678 (N_2678,N_2251,N_2317);
nand U2679 (N_2679,N_2112,N_2120);
nor U2680 (N_2680,N_2339,N_2100);
or U2681 (N_2681,N_2310,N_2334);
and U2682 (N_2682,N_2189,N_2374);
xnor U2683 (N_2683,N_2258,N_2354);
nand U2684 (N_2684,N_2027,N_2062);
nand U2685 (N_2685,N_2275,N_2040);
xnor U2686 (N_2686,N_2263,N_2192);
xor U2687 (N_2687,N_2375,N_2192);
or U2688 (N_2688,N_2393,N_2146);
or U2689 (N_2689,N_2285,N_2139);
and U2690 (N_2690,N_2047,N_2243);
nor U2691 (N_2691,N_2259,N_2327);
or U2692 (N_2692,N_2276,N_2359);
xor U2693 (N_2693,N_2205,N_2244);
xnor U2694 (N_2694,N_2017,N_2164);
nor U2695 (N_2695,N_2162,N_2298);
and U2696 (N_2696,N_2326,N_2306);
nand U2697 (N_2697,N_2198,N_2370);
or U2698 (N_2698,N_2104,N_2391);
and U2699 (N_2699,N_2391,N_2087);
nor U2700 (N_2700,N_2335,N_2349);
nand U2701 (N_2701,N_2360,N_2181);
and U2702 (N_2702,N_2312,N_2329);
or U2703 (N_2703,N_2273,N_2355);
xor U2704 (N_2704,N_2259,N_2123);
xnor U2705 (N_2705,N_2343,N_2038);
nand U2706 (N_2706,N_2050,N_2095);
nand U2707 (N_2707,N_2075,N_2218);
and U2708 (N_2708,N_2043,N_2364);
or U2709 (N_2709,N_2284,N_2322);
nor U2710 (N_2710,N_2149,N_2011);
or U2711 (N_2711,N_2297,N_2067);
and U2712 (N_2712,N_2276,N_2348);
nand U2713 (N_2713,N_2212,N_2031);
nor U2714 (N_2714,N_2312,N_2053);
or U2715 (N_2715,N_2101,N_2302);
xor U2716 (N_2716,N_2051,N_2035);
nand U2717 (N_2717,N_2064,N_2199);
nand U2718 (N_2718,N_2246,N_2212);
xor U2719 (N_2719,N_2121,N_2143);
and U2720 (N_2720,N_2243,N_2003);
xor U2721 (N_2721,N_2310,N_2349);
or U2722 (N_2722,N_2335,N_2111);
nor U2723 (N_2723,N_2263,N_2296);
nand U2724 (N_2724,N_2308,N_2181);
or U2725 (N_2725,N_2303,N_2286);
nand U2726 (N_2726,N_2072,N_2332);
and U2727 (N_2727,N_2296,N_2346);
and U2728 (N_2728,N_2209,N_2307);
xor U2729 (N_2729,N_2220,N_2032);
nand U2730 (N_2730,N_2185,N_2288);
nand U2731 (N_2731,N_2093,N_2242);
and U2732 (N_2732,N_2344,N_2287);
nor U2733 (N_2733,N_2355,N_2342);
xor U2734 (N_2734,N_2028,N_2275);
nor U2735 (N_2735,N_2024,N_2205);
and U2736 (N_2736,N_2117,N_2050);
nor U2737 (N_2737,N_2389,N_2248);
or U2738 (N_2738,N_2021,N_2367);
nand U2739 (N_2739,N_2244,N_2030);
or U2740 (N_2740,N_2385,N_2060);
xor U2741 (N_2741,N_2202,N_2397);
nand U2742 (N_2742,N_2119,N_2075);
or U2743 (N_2743,N_2045,N_2212);
nand U2744 (N_2744,N_2156,N_2266);
and U2745 (N_2745,N_2138,N_2172);
and U2746 (N_2746,N_2209,N_2228);
nor U2747 (N_2747,N_2391,N_2134);
or U2748 (N_2748,N_2158,N_2361);
xor U2749 (N_2749,N_2122,N_2042);
or U2750 (N_2750,N_2168,N_2343);
and U2751 (N_2751,N_2328,N_2371);
xor U2752 (N_2752,N_2297,N_2352);
or U2753 (N_2753,N_2053,N_2153);
xor U2754 (N_2754,N_2199,N_2313);
nor U2755 (N_2755,N_2159,N_2177);
or U2756 (N_2756,N_2159,N_2201);
and U2757 (N_2757,N_2161,N_2266);
nand U2758 (N_2758,N_2233,N_2176);
nor U2759 (N_2759,N_2102,N_2366);
or U2760 (N_2760,N_2042,N_2317);
xor U2761 (N_2761,N_2311,N_2038);
nor U2762 (N_2762,N_2009,N_2093);
and U2763 (N_2763,N_2194,N_2078);
and U2764 (N_2764,N_2334,N_2353);
nand U2765 (N_2765,N_2342,N_2041);
nor U2766 (N_2766,N_2349,N_2327);
and U2767 (N_2767,N_2184,N_2376);
nand U2768 (N_2768,N_2117,N_2206);
nand U2769 (N_2769,N_2219,N_2225);
nor U2770 (N_2770,N_2069,N_2158);
or U2771 (N_2771,N_2126,N_2159);
and U2772 (N_2772,N_2248,N_2208);
xor U2773 (N_2773,N_2008,N_2292);
nor U2774 (N_2774,N_2089,N_2277);
or U2775 (N_2775,N_2093,N_2359);
and U2776 (N_2776,N_2106,N_2295);
and U2777 (N_2777,N_2129,N_2309);
xnor U2778 (N_2778,N_2131,N_2202);
and U2779 (N_2779,N_2334,N_2272);
nor U2780 (N_2780,N_2383,N_2102);
xor U2781 (N_2781,N_2391,N_2175);
xnor U2782 (N_2782,N_2155,N_2076);
and U2783 (N_2783,N_2331,N_2303);
xor U2784 (N_2784,N_2204,N_2276);
and U2785 (N_2785,N_2000,N_2020);
and U2786 (N_2786,N_2224,N_2108);
nand U2787 (N_2787,N_2251,N_2151);
nand U2788 (N_2788,N_2218,N_2120);
or U2789 (N_2789,N_2216,N_2118);
nor U2790 (N_2790,N_2032,N_2188);
xnor U2791 (N_2791,N_2103,N_2378);
nor U2792 (N_2792,N_2238,N_2078);
nor U2793 (N_2793,N_2138,N_2281);
and U2794 (N_2794,N_2387,N_2373);
and U2795 (N_2795,N_2106,N_2234);
nand U2796 (N_2796,N_2269,N_2320);
nand U2797 (N_2797,N_2244,N_2349);
or U2798 (N_2798,N_2005,N_2397);
or U2799 (N_2799,N_2163,N_2155);
or U2800 (N_2800,N_2617,N_2795);
xnor U2801 (N_2801,N_2476,N_2533);
and U2802 (N_2802,N_2701,N_2454);
xor U2803 (N_2803,N_2598,N_2740);
and U2804 (N_2804,N_2716,N_2408);
xnor U2805 (N_2805,N_2775,N_2767);
or U2806 (N_2806,N_2436,N_2559);
xor U2807 (N_2807,N_2681,N_2410);
xnor U2808 (N_2808,N_2616,N_2553);
nor U2809 (N_2809,N_2554,N_2450);
nor U2810 (N_2810,N_2464,N_2516);
and U2811 (N_2811,N_2578,N_2614);
nor U2812 (N_2812,N_2482,N_2550);
or U2813 (N_2813,N_2503,N_2609);
xor U2814 (N_2814,N_2677,N_2526);
xor U2815 (N_2815,N_2600,N_2509);
or U2816 (N_2816,N_2741,N_2678);
xnor U2817 (N_2817,N_2437,N_2539);
xnor U2818 (N_2818,N_2796,N_2702);
and U2819 (N_2819,N_2655,N_2529);
xor U2820 (N_2820,N_2523,N_2628);
or U2821 (N_2821,N_2571,N_2440);
nand U2822 (N_2822,N_2470,N_2764);
xnor U2823 (N_2823,N_2403,N_2487);
and U2824 (N_2824,N_2786,N_2490);
nand U2825 (N_2825,N_2545,N_2738);
or U2826 (N_2826,N_2783,N_2669);
or U2827 (N_2827,N_2698,N_2718);
nor U2828 (N_2828,N_2438,N_2719);
nor U2829 (N_2829,N_2590,N_2615);
nor U2830 (N_2830,N_2761,N_2508);
nand U2831 (N_2831,N_2602,N_2491);
and U2832 (N_2832,N_2452,N_2652);
and U2833 (N_2833,N_2630,N_2460);
or U2834 (N_2834,N_2595,N_2624);
xor U2835 (N_2835,N_2426,N_2721);
and U2836 (N_2836,N_2720,N_2710);
or U2837 (N_2837,N_2463,N_2484);
or U2838 (N_2838,N_2787,N_2404);
xor U2839 (N_2839,N_2688,N_2512);
xor U2840 (N_2840,N_2453,N_2423);
xnor U2841 (N_2841,N_2755,N_2501);
nor U2842 (N_2842,N_2723,N_2548);
or U2843 (N_2843,N_2734,N_2537);
nor U2844 (N_2844,N_2599,N_2750);
nand U2845 (N_2845,N_2444,N_2733);
and U2846 (N_2846,N_2686,N_2531);
nor U2847 (N_2847,N_2447,N_2699);
nand U2848 (N_2848,N_2471,N_2564);
xnor U2849 (N_2849,N_2419,N_2735);
and U2850 (N_2850,N_2416,N_2695);
xor U2851 (N_2851,N_2782,N_2746);
nand U2852 (N_2852,N_2791,N_2751);
nor U2853 (N_2853,N_2629,N_2499);
xor U2854 (N_2854,N_2752,N_2502);
and U2855 (N_2855,N_2400,N_2632);
or U2856 (N_2856,N_2789,N_2724);
or U2857 (N_2857,N_2430,N_2558);
and U2858 (N_2858,N_2648,N_2418);
or U2859 (N_2859,N_2625,N_2428);
nor U2860 (N_2860,N_2663,N_2610);
and U2861 (N_2861,N_2572,N_2641);
or U2862 (N_2862,N_2448,N_2676);
nand U2863 (N_2863,N_2519,N_2459);
and U2864 (N_2864,N_2794,N_2635);
or U2865 (N_2865,N_2504,N_2722);
or U2866 (N_2866,N_2776,N_2777);
xor U2867 (N_2867,N_2665,N_2462);
nand U2868 (N_2868,N_2511,N_2666);
nor U2869 (N_2869,N_2644,N_2481);
xnor U2870 (N_2870,N_2736,N_2797);
nand U2871 (N_2871,N_2506,N_2611);
nand U2872 (N_2872,N_2588,N_2479);
nor U2873 (N_2873,N_2542,N_2662);
nor U2874 (N_2874,N_2445,N_2778);
or U2875 (N_2875,N_2689,N_2427);
or U2876 (N_2876,N_2573,N_2670);
or U2877 (N_2877,N_2601,N_2441);
nand U2878 (N_2878,N_2674,N_2744);
and U2879 (N_2879,N_2684,N_2647);
nand U2880 (N_2880,N_2696,N_2737);
xnor U2881 (N_2881,N_2488,N_2420);
nor U2882 (N_2882,N_2685,N_2730);
or U2883 (N_2883,N_2556,N_2623);
nor U2884 (N_2884,N_2486,N_2691);
nand U2885 (N_2885,N_2792,N_2725);
or U2886 (N_2886,N_2757,N_2726);
xnor U2887 (N_2887,N_2413,N_2434);
or U2888 (N_2888,N_2535,N_2612);
or U2889 (N_2889,N_2580,N_2745);
and U2890 (N_2890,N_2765,N_2525);
and U2891 (N_2891,N_2515,N_2587);
nand U2892 (N_2892,N_2653,N_2498);
and U2893 (N_2893,N_2522,N_2579);
xor U2894 (N_2894,N_2766,N_2443);
nor U2895 (N_2895,N_2524,N_2634);
or U2896 (N_2896,N_2622,N_2705);
xor U2897 (N_2897,N_2402,N_2456);
and U2898 (N_2898,N_2687,N_2620);
xnor U2899 (N_2899,N_2566,N_2603);
or U2900 (N_2900,N_2656,N_2500);
and U2901 (N_2901,N_2706,N_2704);
xor U2902 (N_2902,N_2754,N_2461);
and U2903 (N_2903,N_2497,N_2478);
nand U2904 (N_2904,N_2439,N_2798);
or U2905 (N_2905,N_2412,N_2520);
or U2906 (N_2906,N_2651,N_2582);
nor U2907 (N_2907,N_2492,N_2465);
or U2908 (N_2908,N_2435,N_2643);
nand U2909 (N_2909,N_2591,N_2790);
nand U2910 (N_2910,N_2679,N_2496);
or U2911 (N_2911,N_2561,N_2536);
and U2912 (N_2912,N_2528,N_2668);
nand U2913 (N_2913,N_2407,N_2417);
xnor U2914 (N_2914,N_2715,N_2514);
and U2915 (N_2915,N_2494,N_2594);
nand U2916 (N_2916,N_2631,N_2619);
nand U2917 (N_2917,N_2527,N_2431);
and U2918 (N_2918,N_2432,N_2645);
xnor U2919 (N_2919,N_2758,N_2727);
or U2920 (N_2920,N_2469,N_2749);
nor U2921 (N_2921,N_2414,N_2664);
nor U2922 (N_2922,N_2411,N_2541);
and U2923 (N_2923,N_2785,N_2521);
and U2924 (N_2924,N_2485,N_2592);
nor U2925 (N_2925,N_2781,N_2732);
nand U2926 (N_2926,N_2661,N_2711);
and U2927 (N_2927,N_2583,N_2731);
or U2928 (N_2928,N_2690,N_2707);
nor U2929 (N_2929,N_2557,N_2532);
xnor U2930 (N_2930,N_2607,N_2473);
nor U2931 (N_2931,N_2646,N_2513);
nor U2932 (N_2932,N_2567,N_2683);
or U2933 (N_2933,N_2467,N_2475);
or U2934 (N_2934,N_2618,N_2709);
xnor U2935 (N_2935,N_2784,N_2534);
nor U2936 (N_2936,N_2405,N_2458);
or U2937 (N_2937,N_2593,N_2507);
nand U2938 (N_2938,N_2597,N_2799);
xnor U2939 (N_2939,N_2409,N_2585);
nand U2940 (N_2940,N_2574,N_2606);
nand U2941 (N_2941,N_2640,N_2763);
or U2942 (N_2942,N_2480,N_2449);
or U2943 (N_2943,N_2472,N_2576);
or U2944 (N_2944,N_2633,N_2667);
nand U2945 (N_2945,N_2466,N_2760);
nor U2946 (N_2946,N_2682,N_2510);
xor U2947 (N_2947,N_2788,N_2406);
and U2948 (N_2948,N_2742,N_2717);
xnor U2949 (N_2949,N_2756,N_2672);
or U2950 (N_2950,N_2729,N_2659);
or U2951 (N_2951,N_2739,N_2547);
nor U2952 (N_2952,N_2642,N_2446);
or U2953 (N_2953,N_2621,N_2650);
or U2954 (N_2954,N_2489,N_2604);
and U2955 (N_2955,N_2581,N_2455);
and U2956 (N_2956,N_2433,N_2584);
and U2957 (N_2957,N_2565,N_2560);
nand U2958 (N_2958,N_2425,N_2713);
and U2959 (N_2959,N_2401,N_2636);
and U2960 (N_2960,N_2546,N_2575);
nor U2961 (N_2961,N_2549,N_2654);
nor U2962 (N_2962,N_2468,N_2517);
xor U2963 (N_2963,N_2712,N_2700);
nor U2964 (N_2964,N_2743,N_2657);
and U2965 (N_2965,N_2769,N_2770);
and U2966 (N_2966,N_2552,N_2639);
nor U2967 (N_2967,N_2596,N_2483);
nand U2968 (N_2968,N_2540,N_2728);
nor U2969 (N_2969,N_2569,N_2538);
and U2970 (N_2970,N_2518,N_2673);
and U2971 (N_2971,N_2694,N_2772);
xor U2972 (N_2972,N_2793,N_2671);
or U2973 (N_2973,N_2530,N_2442);
or U2974 (N_2974,N_2780,N_2543);
and U2975 (N_2975,N_2568,N_2779);
or U2976 (N_2976,N_2577,N_2774);
nand U2977 (N_2977,N_2626,N_2697);
nand U2978 (N_2978,N_2605,N_2457);
nor U2979 (N_2979,N_2675,N_2768);
nand U2980 (N_2980,N_2773,N_2747);
xor U2981 (N_2981,N_2563,N_2692);
or U2982 (N_2982,N_2680,N_2429);
and U2983 (N_2983,N_2703,N_2748);
xnor U2984 (N_2984,N_2493,N_2608);
and U2985 (N_2985,N_2555,N_2708);
and U2986 (N_2986,N_2714,N_2762);
nor U2987 (N_2987,N_2570,N_2562);
or U2988 (N_2988,N_2753,N_2759);
nor U2989 (N_2989,N_2627,N_2638);
and U2990 (N_2990,N_2415,N_2505);
nor U2991 (N_2991,N_2771,N_2474);
nand U2992 (N_2992,N_2451,N_2637);
nor U2993 (N_2993,N_2477,N_2422);
xnor U2994 (N_2994,N_2660,N_2495);
xnor U2995 (N_2995,N_2693,N_2544);
or U2996 (N_2996,N_2424,N_2649);
nand U2997 (N_2997,N_2586,N_2551);
xor U2998 (N_2998,N_2613,N_2658);
nor U2999 (N_2999,N_2421,N_2589);
nor U3000 (N_3000,N_2642,N_2402);
nand U3001 (N_3001,N_2787,N_2770);
or U3002 (N_3002,N_2463,N_2776);
nor U3003 (N_3003,N_2631,N_2479);
nand U3004 (N_3004,N_2777,N_2488);
xor U3005 (N_3005,N_2727,N_2726);
xnor U3006 (N_3006,N_2435,N_2420);
nand U3007 (N_3007,N_2499,N_2756);
nor U3008 (N_3008,N_2658,N_2536);
or U3009 (N_3009,N_2476,N_2464);
nand U3010 (N_3010,N_2627,N_2731);
xor U3011 (N_3011,N_2699,N_2764);
xor U3012 (N_3012,N_2659,N_2767);
or U3013 (N_3013,N_2463,N_2671);
and U3014 (N_3014,N_2777,N_2746);
nand U3015 (N_3015,N_2478,N_2703);
xor U3016 (N_3016,N_2630,N_2685);
and U3017 (N_3017,N_2531,N_2774);
nor U3018 (N_3018,N_2506,N_2551);
or U3019 (N_3019,N_2404,N_2620);
xnor U3020 (N_3020,N_2690,N_2532);
and U3021 (N_3021,N_2632,N_2456);
nor U3022 (N_3022,N_2649,N_2407);
nand U3023 (N_3023,N_2576,N_2450);
or U3024 (N_3024,N_2719,N_2767);
or U3025 (N_3025,N_2767,N_2578);
nor U3026 (N_3026,N_2469,N_2408);
xor U3027 (N_3027,N_2592,N_2506);
nand U3028 (N_3028,N_2798,N_2548);
or U3029 (N_3029,N_2614,N_2684);
nand U3030 (N_3030,N_2620,N_2666);
xnor U3031 (N_3031,N_2517,N_2606);
or U3032 (N_3032,N_2527,N_2745);
nor U3033 (N_3033,N_2549,N_2562);
nor U3034 (N_3034,N_2477,N_2629);
and U3035 (N_3035,N_2405,N_2723);
nor U3036 (N_3036,N_2473,N_2664);
and U3037 (N_3037,N_2552,N_2643);
or U3038 (N_3038,N_2554,N_2429);
nand U3039 (N_3039,N_2754,N_2645);
nand U3040 (N_3040,N_2425,N_2484);
xor U3041 (N_3041,N_2658,N_2703);
and U3042 (N_3042,N_2497,N_2736);
and U3043 (N_3043,N_2487,N_2576);
nor U3044 (N_3044,N_2579,N_2689);
and U3045 (N_3045,N_2596,N_2768);
nor U3046 (N_3046,N_2584,N_2446);
and U3047 (N_3047,N_2796,N_2622);
nor U3048 (N_3048,N_2430,N_2530);
nand U3049 (N_3049,N_2546,N_2442);
nor U3050 (N_3050,N_2779,N_2644);
nor U3051 (N_3051,N_2516,N_2424);
nand U3052 (N_3052,N_2759,N_2537);
nand U3053 (N_3053,N_2700,N_2467);
and U3054 (N_3054,N_2622,N_2699);
or U3055 (N_3055,N_2544,N_2526);
xnor U3056 (N_3056,N_2731,N_2452);
or U3057 (N_3057,N_2441,N_2532);
and U3058 (N_3058,N_2498,N_2441);
and U3059 (N_3059,N_2645,N_2623);
nor U3060 (N_3060,N_2539,N_2411);
or U3061 (N_3061,N_2701,N_2767);
xnor U3062 (N_3062,N_2690,N_2452);
nor U3063 (N_3063,N_2688,N_2670);
or U3064 (N_3064,N_2618,N_2426);
nand U3065 (N_3065,N_2451,N_2553);
xnor U3066 (N_3066,N_2538,N_2589);
or U3067 (N_3067,N_2591,N_2561);
or U3068 (N_3068,N_2506,N_2748);
and U3069 (N_3069,N_2685,N_2505);
and U3070 (N_3070,N_2446,N_2497);
or U3071 (N_3071,N_2475,N_2743);
nand U3072 (N_3072,N_2478,N_2513);
nand U3073 (N_3073,N_2659,N_2462);
nor U3074 (N_3074,N_2790,N_2428);
or U3075 (N_3075,N_2741,N_2544);
nand U3076 (N_3076,N_2699,N_2565);
xor U3077 (N_3077,N_2515,N_2606);
xnor U3078 (N_3078,N_2764,N_2672);
and U3079 (N_3079,N_2513,N_2451);
and U3080 (N_3080,N_2465,N_2613);
and U3081 (N_3081,N_2777,N_2587);
xnor U3082 (N_3082,N_2723,N_2749);
nand U3083 (N_3083,N_2582,N_2568);
nor U3084 (N_3084,N_2485,N_2672);
or U3085 (N_3085,N_2410,N_2640);
or U3086 (N_3086,N_2660,N_2609);
and U3087 (N_3087,N_2649,N_2664);
xnor U3088 (N_3088,N_2503,N_2716);
nor U3089 (N_3089,N_2641,N_2630);
and U3090 (N_3090,N_2492,N_2772);
and U3091 (N_3091,N_2663,N_2720);
xor U3092 (N_3092,N_2777,N_2453);
nand U3093 (N_3093,N_2428,N_2678);
nor U3094 (N_3094,N_2622,N_2546);
and U3095 (N_3095,N_2663,N_2606);
xnor U3096 (N_3096,N_2511,N_2573);
nand U3097 (N_3097,N_2784,N_2602);
xnor U3098 (N_3098,N_2781,N_2774);
and U3099 (N_3099,N_2742,N_2796);
xor U3100 (N_3100,N_2603,N_2597);
xnor U3101 (N_3101,N_2588,N_2650);
xnor U3102 (N_3102,N_2706,N_2510);
nand U3103 (N_3103,N_2512,N_2687);
nand U3104 (N_3104,N_2793,N_2425);
xor U3105 (N_3105,N_2490,N_2778);
xnor U3106 (N_3106,N_2483,N_2612);
nand U3107 (N_3107,N_2637,N_2770);
and U3108 (N_3108,N_2490,N_2738);
nor U3109 (N_3109,N_2457,N_2703);
nand U3110 (N_3110,N_2408,N_2479);
or U3111 (N_3111,N_2597,N_2515);
xnor U3112 (N_3112,N_2622,N_2497);
xnor U3113 (N_3113,N_2706,N_2619);
nand U3114 (N_3114,N_2658,N_2540);
and U3115 (N_3115,N_2778,N_2524);
xnor U3116 (N_3116,N_2508,N_2491);
nor U3117 (N_3117,N_2473,N_2763);
xor U3118 (N_3118,N_2583,N_2506);
nand U3119 (N_3119,N_2457,N_2639);
or U3120 (N_3120,N_2492,N_2447);
or U3121 (N_3121,N_2540,N_2428);
nor U3122 (N_3122,N_2580,N_2528);
or U3123 (N_3123,N_2495,N_2684);
and U3124 (N_3124,N_2469,N_2624);
nor U3125 (N_3125,N_2475,N_2450);
nand U3126 (N_3126,N_2552,N_2785);
xor U3127 (N_3127,N_2536,N_2428);
or U3128 (N_3128,N_2513,N_2536);
or U3129 (N_3129,N_2424,N_2735);
and U3130 (N_3130,N_2712,N_2611);
nand U3131 (N_3131,N_2434,N_2545);
nand U3132 (N_3132,N_2655,N_2698);
nor U3133 (N_3133,N_2711,N_2797);
xor U3134 (N_3134,N_2495,N_2469);
and U3135 (N_3135,N_2627,N_2568);
nand U3136 (N_3136,N_2786,N_2781);
xnor U3137 (N_3137,N_2658,N_2701);
xnor U3138 (N_3138,N_2642,N_2694);
xor U3139 (N_3139,N_2519,N_2495);
xnor U3140 (N_3140,N_2422,N_2591);
or U3141 (N_3141,N_2791,N_2754);
xnor U3142 (N_3142,N_2611,N_2488);
or U3143 (N_3143,N_2793,N_2443);
or U3144 (N_3144,N_2699,N_2525);
nand U3145 (N_3145,N_2512,N_2785);
or U3146 (N_3146,N_2574,N_2422);
and U3147 (N_3147,N_2516,N_2445);
nand U3148 (N_3148,N_2726,N_2423);
nand U3149 (N_3149,N_2675,N_2488);
nand U3150 (N_3150,N_2622,N_2634);
and U3151 (N_3151,N_2618,N_2487);
xnor U3152 (N_3152,N_2421,N_2726);
xor U3153 (N_3153,N_2745,N_2758);
nor U3154 (N_3154,N_2776,N_2575);
nand U3155 (N_3155,N_2444,N_2430);
nor U3156 (N_3156,N_2603,N_2568);
nand U3157 (N_3157,N_2676,N_2721);
and U3158 (N_3158,N_2753,N_2587);
or U3159 (N_3159,N_2731,N_2521);
nand U3160 (N_3160,N_2629,N_2405);
xnor U3161 (N_3161,N_2685,N_2788);
nor U3162 (N_3162,N_2466,N_2519);
nand U3163 (N_3163,N_2685,N_2634);
xnor U3164 (N_3164,N_2564,N_2615);
xnor U3165 (N_3165,N_2700,N_2592);
nand U3166 (N_3166,N_2660,N_2741);
and U3167 (N_3167,N_2720,N_2587);
xor U3168 (N_3168,N_2518,N_2563);
xor U3169 (N_3169,N_2569,N_2773);
or U3170 (N_3170,N_2738,N_2429);
xor U3171 (N_3171,N_2716,N_2645);
and U3172 (N_3172,N_2542,N_2421);
and U3173 (N_3173,N_2661,N_2655);
xor U3174 (N_3174,N_2767,N_2588);
xor U3175 (N_3175,N_2415,N_2730);
xnor U3176 (N_3176,N_2456,N_2451);
nor U3177 (N_3177,N_2487,N_2474);
and U3178 (N_3178,N_2708,N_2596);
nand U3179 (N_3179,N_2481,N_2600);
or U3180 (N_3180,N_2595,N_2452);
xor U3181 (N_3181,N_2775,N_2665);
xnor U3182 (N_3182,N_2747,N_2683);
or U3183 (N_3183,N_2547,N_2478);
nor U3184 (N_3184,N_2466,N_2623);
xnor U3185 (N_3185,N_2754,N_2710);
and U3186 (N_3186,N_2756,N_2767);
xnor U3187 (N_3187,N_2652,N_2680);
nand U3188 (N_3188,N_2585,N_2782);
nand U3189 (N_3189,N_2497,N_2419);
and U3190 (N_3190,N_2609,N_2681);
and U3191 (N_3191,N_2455,N_2740);
nor U3192 (N_3192,N_2784,N_2601);
nand U3193 (N_3193,N_2722,N_2602);
nand U3194 (N_3194,N_2796,N_2736);
nand U3195 (N_3195,N_2753,N_2603);
nand U3196 (N_3196,N_2476,N_2635);
nor U3197 (N_3197,N_2674,N_2644);
nor U3198 (N_3198,N_2671,N_2752);
xnor U3199 (N_3199,N_2478,N_2483);
nand U3200 (N_3200,N_3174,N_3087);
nor U3201 (N_3201,N_2997,N_2980);
or U3202 (N_3202,N_2954,N_2832);
nor U3203 (N_3203,N_2895,N_2900);
nor U3204 (N_3204,N_2800,N_2872);
and U3205 (N_3205,N_3197,N_2886);
xnor U3206 (N_3206,N_3120,N_3117);
nor U3207 (N_3207,N_2890,N_3078);
nand U3208 (N_3208,N_2998,N_2920);
or U3209 (N_3209,N_2961,N_3046);
nand U3210 (N_3210,N_3155,N_2993);
xor U3211 (N_3211,N_3157,N_2973);
nor U3212 (N_3212,N_3070,N_2976);
or U3213 (N_3213,N_2873,N_3053);
nand U3214 (N_3214,N_3129,N_2851);
nand U3215 (N_3215,N_3131,N_3082);
nand U3216 (N_3216,N_3011,N_2987);
nor U3217 (N_3217,N_2990,N_3090);
and U3218 (N_3218,N_2807,N_3041);
nand U3219 (N_3219,N_2950,N_3072);
and U3220 (N_3220,N_3153,N_2805);
nand U3221 (N_3221,N_2971,N_3170);
xnor U3222 (N_3222,N_3056,N_3002);
and U3223 (N_3223,N_2836,N_2910);
and U3224 (N_3224,N_2866,N_3022);
and U3225 (N_3225,N_2929,N_3043);
and U3226 (N_3226,N_3029,N_2962);
nor U3227 (N_3227,N_2880,N_3137);
xor U3228 (N_3228,N_3091,N_2983);
and U3229 (N_3229,N_3037,N_3190);
and U3230 (N_3230,N_2869,N_3062);
xor U3231 (N_3231,N_3024,N_2948);
nor U3232 (N_3232,N_3001,N_2808);
xor U3233 (N_3233,N_2943,N_3086);
and U3234 (N_3234,N_3150,N_2887);
nand U3235 (N_3235,N_3135,N_2958);
or U3236 (N_3236,N_2906,N_3069);
and U3237 (N_3237,N_3165,N_3143);
nand U3238 (N_3238,N_2904,N_2848);
nor U3239 (N_3239,N_3154,N_3030);
or U3240 (N_3240,N_2926,N_3144);
nand U3241 (N_3241,N_3164,N_2953);
xor U3242 (N_3242,N_3012,N_2828);
and U3243 (N_3243,N_2879,N_2989);
and U3244 (N_3244,N_2889,N_2806);
and U3245 (N_3245,N_2944,N_2902);
or U3246 (N_3246,N_2975,N_3077);
nand U3247 (N_3247,N_2901,N_3175);
xnor U3248 (N_3248,N_2974,N_2838);
or U3249 (N_3249,N_2982,N_2959);
and U3250 (N_3250,N_2915,N_3100);
nand U3251 (N_3251,N_2858,N_2937);
xnor U3252 (N_3252,N_3179,N_3139);
nor U3253 (N_3253,N_3092,N_3027);
nand U3254 (N_3254,N_2995,N_3187);
xnor U3255 (N_3255,N_2899,N_2924);
xor U3256 (N_3256,N_2933,N_3186);
nand U3257 (N_3257,N_2951,N_2865);
xnor U3258 (N_3258,N_3066,N_2883);
nand U3259 (N_3259,N_3020,N_2857);
and U3260 (N_3260,N_3196,N_3096);
and U3261 (N_3261,N_2907,N_2863);
nand U3262 (N_3262,N_2957,N_2918);
xnor U3263 (N_3263,N_3185,N_2817);
or U3264 (N_3264,N_3004,N_2970);
nor U3265 (N_3265,N_3057,N_2809);
or U3266 (N_3266,N_3158,N_3166);
or U3267 (N_3267,N_2853,N_3149);
xnor U3268 (N_3268,N_3048,N_2979);
and U3269 (N_3269,N_2823,N_3050);
nor U3270 (N_3270,N_3036,N_3095);
or U3271 (N_3271,N_3097,N_3010);
and U3272 (N_3272,N_2803,N_3108);
and U3273 (N_3273,N_3146,N_3047);
and U3274 (N_3274,N_3122,N_2927);
nor U3275 (N_3275,N_2855,N_3008);
nand U3276 (N_3276,N_3184,N_3017);
and U3277 (N_3277,N_3136,N_3189);
nand U3278 (N_3278,N_3064,N_3128);
nand U3279 (N_3279,N_3198,N_2934);
nand U3280 (N_3280,N_2938,N_2964);
and U3281 (N_3281,N_3034,N_2871);
or U3282 (N_3282,N_2942,N_2860);
or U3283 (N_3283,N_2963,N_2984);
or U3284 (N_3284,N_2816,N_3065);
nand U3285 (N_3285,N_3089,N_3079);
nand U3286 (N_3286,N_2829,N_3102);
nand U3287 (N_3287,N_3044,N_3052);
xnor U3288 (N_3288,N_2815,N_2847);
and U3289 (N_3289,N_2876,N_2814);
and U3290 (N_3290,N_3073,N_2822);
or U3291 (N_3291,N_3031,N_2881);
nand U3292 (N_3292,N_3173,N_3023);
xor U3293 (N_3293,N_3183,N_2986);
xor U3294 (N_3294,N_3105,N_3101);
nand U3295 (N_3295,N_3076,N_2968);
nand U3296 (N_3296,N_3114,N_2852);
nand U3297 (N_3297,N_2845,N_3060);
nand U3298 (N_3298,N_3177,N_3025);
or U3299 (N_3299,N_2992,N_3113);
or U3300 (N_3300,N_3075,N_2875);
nor U3301 (N_3301,N_2884,N_2894);
xor U3302 (N_3302,N_3099,N_2801);
xnor U3303 (N_3303,N_3007,N_3033);
nor U3304 (N_3304,N_2932,N_2820);
xnor U3305 (N_3305,N_2867,N_3140);
and U3306 (N_3306,N_2916,N_2825);
nor U3307 (N_3307,N_3009,N_2818);
xor U3308 (N_3308,N_2912,N_2956);
nor U3309 (N_3309,N_3182,N_3018);
nand U3310 (N_3310,N_3055,N_3093);
and U3311 (N_3311,N_3045,N_2905);
nor U3312 (N_3312,N_3195,N_2988);
nand U3313 (N_3313,N_2911,N_3125);
or U3314 (N_3314,N_3172,N_2922);
and U3315 (N_3315,N_3094,N_3199);
and U3316 (N_3316,N_3112,N_2877);
nor U3317 (N_3317,N_3019,N_3147);
or U3318 (N_3318,N_2966,N_2892);
nand U3319 (N_3319,N_3000,N_2999);
nor U3320 (N_3320,N_3088,N_2947);
nand U3321 (N_3321,N_2952,N_2827);
nand U3322 (N_3322,N_3071,N_3104);
or U3323 (N_3323,N_3014,N_2914);
or U3324 (N_3324,N_3039,N_3051);
nor U3325 (N_3325,N_2885,N_3188);
nand U3326 (N_3326,N_3171,N_2903);
nand U3327 (N_3327,N_3123,N_3110);
nor U3328 (N_3328,N_3168,N_2967);
nand U3329 (N_3329,N_3119,N_3180);
nor U3330 (N_3330,N_2991,N_2931);
nand U3331 (N_3331,N_2965,N_3169);
xor U3332 (N_3332,N_2891,N_3016);
nor U3333 (N_3333,N_2882,N_3124);
xor U3334 (N_3334,N_3005,N_3006);
xor U3335 (N_3335,N_3059,N_3049);
xnor U3336 (N_3336,N_3159,N_3152);
nand U3337 (N_3337,N_2996,N_2945);
xnor U3338 (N_3338,N_3163,N_3015);
nor U3339 (N_3339,N_3126,N_2859);
nor U3340 (N_3340,N_3103,N_3080);
and U3341 (N_3341,N_2981,N_3028);
or U3342 (N_3342,N_2844,N_2834);
or U3343 (N_3343,N_2960,N_3121);
and U3344 (N_3344,N_2969,N_2977);
xor U3345 (N_3345,N_3148,N_3074);
xor U3346 (N_3346,N_3040,N_3111);
or U3347 (N_3347,N_2955,N_3176);
nor U3348 (N_3348,N_3138,N_3161);
or U3349 (N_3349,N_2917,N_3181);
nor U3350 (N_3350,N_3107,N_2862);
or U3351 (N_3351,N_3061,N_2821);
xor U3352 (N_3352,N_2925,N_3116);
or U3353 (N_3353,N_2921,N_2843);
nor U3354 (N_3354,N_2939,N_2861);
and U3355 (N_3355,N_3191,N_2802);
and U3356 (N_3356,N_2854,N_2849);
or U3357 (N_3357,N_2833,N_2878);
and U3358 (N_3358,N_3142,N_3141);
xnor U3359 (N_3359,N_3083,N_2830);
nor U3360 (N_3360,N_3162,N_3167);
nand U3361 (N_3361,N_3021,N_3085);
and U3362 (N_3362,N_3134,N_3194);
nand U3363 (N_3363,N_3035,N_2874);
or U3364 (N_3364,N_2864,N_2897);
nor U3365 (N_3365,N_3151,N_2811);
nand U3366 (N_3366,N_3003,N_2919);
xnor U3367 (N_3367,N_2946,N_3058);
nand U3368 (N_3368,N_3063,N_3133);
xnor U3369 (N_3369,N_2985,N_2826);
xnor U3370 (N_3370,N_2935,N_2941);
xor U3371 (N_3371,N_3192,N_2936);
and U3372 (N_3372,N_2923,N_3081);
nand U3373 (N_3373,N_3067,N_2837);
and U3374 (N_3374,N_2850,N_2846);
nand U3375 (N_3375,N_3145,N_3068);
xor U3376 (N_3376,N_3130,N_3098);
and U3377 (N_3377,N_2870,N_3013);
nand U3378 (N_3378,N_2930,N_3156);
xnor U3379 (N_3379,N_2978,N_2908);
and U3380 (N_3380,N_2813,N_2893);
nor U3381 (N_3381,N_3118,N_3038);
or U3382 (N_3382,N_2831,N_2824);
xor U3383 (N_3383,N_3032,N_3193);
and U3384 (N_3384,N_2909,N_2949);
xnor U3385 (N_3385,N_3132,N_2898);
nor U3386 (N_3386,N_2804,N_2842);
or U3387 (N_3387,N_3127,N_2913);
and U3388 (N_3388,N_2928,N_2839);
nand U3389 (N_3389,N_2994,N_3115);
nand U3390 (N_3390,N_2888,N_2940);
and U3391 (N_3391,N_3084,N_2812);
nor U3392 (N_3392,N_3042,N_2841);
or U3393 (N_3393,N_3178,N_3160);
nor U3394 (N_3394,N_2810,N_3054);
nor U3395 (N_3395,N_3106,N_3026);
and U3396 (N_3396,N_2819,N_2972);
xor U3397 (N_3397,N_3109,N_2896);
or U3398 (N_3398,N_2868,N_2835);
nand U3399 (N_3399,N_2840,N_2856);
or U3400 (N_3400,N_3174,N_3044);
nor U3401 (N_3401,N_3065,N_2966);
or U3402 (N_3402,N_3167,N_3094);
nor U3403 (N_3403,N_2952,N_3044);
or U3404 (N_3404,N_2864,N_2978);
nand U3405 (N_3405,N_2901,N_2868);
xor U3406 (N_3406,N_2963,N_3112);
xor U3407 (N_3407,N_3121,N_3039);
nand U3408 (N_3408,N_2803,N_2919);
or U3409 (N_3409,N_3198,N_2809);
and U3410 (N_3410,N_2947,N_2991);
nand U3411 (N_3411,N_3160,N_2813);
nand U3412 (N_3412,N_2838,N_3019);
or U3413 (N_3413,N_3043,N_2916);
or U3414 (N_3414,N_2828,N_2944);
nand U3415 (N_3415,N_2889,N_2910);
and U3416 (N_3416,N_3057,N_2864);
xor U3417 (N_3417,N_3190,N_3088);
and U3418 (N_3418,N_2852,N_2903);
nand U3419 (N_3419,N_2928,N_2810);
or U3420 (N_3420,N_2947,N_3026);
and U3421 (N_3421,N_2818,N_3090);
xor U3422 (N_3422,N_3111,N_2801);
and U3423 (N_3423,N_2861,N_3006);
or U3424 (N_3424,N_3053,N_2871);
or U3425 (N_3425,N_3170,N_3040);
xnor U3426 (N_3426,N_3047,N_3111);
xnor U3427 (N_3427,N_2900,N_2905);
or U3428 (N_3428,N_2832,N_3078);
nand U3429 (N_3429,N_2875,N_2920);
and U3430 (N_3430,N_2892,N_3098);
nor U3431 (N_3431,N_2861,N_2890);
xnor U3432 (N_3432,N_3124,N_3188);
nand U3433 (N_3433,N_2923,N_2867);
or U3434 (N_3434,N_3178,N_3122);
xor U3435 (N_3435,N_3135,N_3188);
or U3436 (N_3436,N_2905,N_3105);
xor U3437 (N_3437,N_2858,N_3099);
and U3438 (N_3438,N_3161,N_3074);
xor U3439 (N_3439,N_2813,N_2864);
or U3440 (N_3440,N_2887,N_2961);
or U3441 (N_3441,N_2844,N_2812);
nor U3442 (N_3442,N_2805,N_2873);
xor U3443 (N_3443,N_2937,N_3011);
nor U3444 (N_3444,N_2967,N_2887);
and U3445 (N_3445,N_3197,N_3015);
nor U3446 (N_3446,N_2944,N_3002);
xor U3447 (N_3447,N_2825,N_2939);
nor U3448 (N_3448,N_2989,N_3067);
nand U3449 (N_3449,N_2853,N_3193);
xnor U3450 (N_3450,N_2852,N_3044);
or U3451 (N_3451,N_3045,N_3117);
or U3452 (N_3452,N_3154,N_3182);
xor U3453 (N_3453,N_2913,N_2918);
nand U3454 (N_3454,N_3128,N_3119);
nor U3455 (N_3455,N_2886,N_2922);
nor U3456 (N_3456,N_3066,N_2897);
and U3457 (N_3457,N_2890,N_2935);
nor U3458 (N_3458,N_2839,N_2982);
xor U3459 (N_3459,N_2845,N_2993);
and U3460 (N_3460,N_2855,N_2853);
xnor U3461 (N_3461,N_2982,N_2967);
nor U3462 (N_3462,N_2825,N_3160);
nor U3463 (N_3463,N_2916,N_3137);
xnor U3464 (N_3464,N_3050,N_3195);
nand U3465 (N_3465,N_3082,N_3087);
nor U3466 (N_3466,N_3148,N_3008);
nand U3467 (N_3467,N_2826,N_2955);
or U3468 (N_3468,N_2803,N_2866);
or U3469 (N_3469,N_2905,N_3124);
nand U3470 (N_3470,N_3114,N_2815);
and U3471 (N_3471,N_2935,N_3063);
and U3472 (N_3472,N_2989,N_3028);
nand U3473 (N_3473,N_2971,N_2927);
xnor U3474 (N_3474,N_2941,N_3078);
nand U3475 (N_3475,N_2896,N_3151);
xnor U3476 (N_3476,N_2842,N_2923);
xnor U3477 (N_3477,N_2875,N_3063);
nand U3478 (N_3478,N_2868,N_3164);
or U3479 (N_3479,N_3190,N_3014);
xnor U3480 (N_3480,N_3060,N_2816);
nand U3481 (N_3481,N_3152,N_2828);
nand U3482 (N_3482,N_2877,N_3098);
nand U3483 (N_3483,N_3104,N_2959);
nand U3484 (N_3484,N_3081,N_3168);
nor U3485 (N_3485,N_3070,N_2921);
xnor U3486 (N_3486,N_3101,N_3047);
xor U3487 (N_3487,N_3156,N_2859);
xnor U3488 (N_3488,N_3143,N_3159);
and U3489 (N_3489,N_2831,N_3064);
xor U3490 (N_3490,N_2922,N_3136);
xnor U3491 (N_3491,N_2962,N_3080);
and U3492 (N_3492,N_2847,N_3085);
and U3493 (N_3493,N_2878,N_3055);
nand U3494 (N_3494,N_3036,N_2981);
or U3495 (N_3495,N_3032,N_2897);
nand U3496 (N_3496,N_2946,N_2954);
nand U3497 (N_3497,N_3195,N_2996);
nand U3498 (N_3498,N_2998,N_2901);
xnor U3499 (N_3499,N_2855,N_2978);
nand U3500 (N_3500,N_3146,N_3193);
xnor U3501 (N_3501,N_3055,N_2909);
and U3502 (N_3502,N_2879,N_2977);
nor U3503 (N_3503,N_2873,N_2908);
nor U3504 (N_3504,N_2929,N_2850);
or U3505 (N_3505,N_2821,N_2838);
nor U3506 (N_3506,N_2926,N_2816);
xor U3507 (N_3507,N_2801,N_2887);
xnor U3508 (N_3508,N_3093,N_2832);
nor U3509 (N_3509,N_3130,N_3180);
xnor U3510 (N_3510,N_3166,N_2918);
or U3511 (N_3511,N_2829,N_3116);
nand U3512 (N_3512,N_2902,N_2928);
and U3513 (N_3513,N_3138,N_3046);
nand U3514 (N_3514,N_3050,N_2907);
or U3515 (N_3515,N_3101,N_3069);
nand U3516 (N_3516,N_2839,N_2804);
nand U3517 (N_3517,N_3143,N_3073);
or U3518 (N_3518,N_2946,N_3082);
xnor U3519 (N_3519,N_2979,N_2997);
nor U3520 (N_3520,N_2801,N_3172);
or U3521 (N_3521,N_2829,N_3049);
or U3522 (N_3522,N_2934,N_3159);
and U3523 (N_3523,N_2937,N_3158);
nand U3524 (N_3524,N_2846,N_2933);
or U3525 (N_3525,N_3083,N_3105);
xor U3526 (N_3526,N_2938,N_3052);
nand U3527 (N_3527,N_2926,N_3141);
nand U3528 (N_3528,N_3004,N_3133);
and U3529 (N_3529,N_2837,N_2996);
nand U3530 (N_3530,N_2856,N_2972);
and U3531 (N_3531,N_3119,N_3089);
nand U3532 (N_3532,N_2887,N_3044);
nor U3533 (N_3533,N_2984,N_2824);
nand U3534 (N_3534,N_3000,N_3041);
or U3535 (N_3535,N_3125,N_2914);
or U3536 (N_3536,N_2848,N_2993);
and U3537 (N_3537,N_2896,N_3113);
or U3538 (N_3538,N_2908,N_3178);
nand U3539 (N_3539,N_2917,N_3023);
and U3540 (N_3540,N_2915,N_3107);
nor U3541 (N_3541,N_2853,N_3054);
or U3542 (N_3542,N_2824,N_3027);
xor U3543 (N_3543,N_2924,N_2908);
xor U3544 (N_3544,N_2854,N_2907);
xnor U3545 (N_3545,N_3052,N_3194);
nor U3546 (N_3546,N_2974,N_3040);
and U3547 (N_3547,N_3056,N_3137);
xor U3548 (N_3548,N_3039,N_3079);
or U3549 (N_3549,N_2825,N_3086);
xnor U3550 (N_3550,N_3117,N_3063);
nor U3551 (N_3551,N_2896,N_2997);
and U3552 (N_3552,N_3126,N_3029);
xor U3553 (N_3553,N_2928,N_3058);
or U3554 (N_3554,N_3098,N_2994);
xor U3555 (N_3555,N_2896,N_2943);
or U3556 (N_3556,N_2828,N_2876);
nor U3557 (N_3557,N_2822,N_2971);
xnor U3558 (N_3558,N_3020,N_2807);
or U3559 (N_3559,N_3139,N_3107);
nand U3560 (N_3560,N_2958,N_3165);
and U3561 (N_3561,N_2950,N_3153);
nor U3562 (N_3562,N_3082,N_2960);
or U3563 (N_3563,N_3185,N_2994);
nor U3564 (N_3564,N_3120,N_2880);
nor U3565 (N_3565,N_2811,N_2800);
and U3566 (N_3566,N_3182,N_3176);
and U3567 (N_3567,N_3092,N_2920);
xor U3568 (N_3568,N_2853,N_2965);
nand U3569 (N_3569,N_2872,N_3145);
or U3570 (N_3570,N_2820,N_3014);
nor U3571 (N_3571,N_3135,N_3102);
nor U3572 (N_3572,N_3128,N_3138);
nand U3573 (N_3573,N_3050,N_3198);
nor U3574 (N_3574,N_3022,N_2891);
and U3575 (N_3575,N_2879,N_2914);
or U3576 (N_3576,N_3099,N_2957);
nand U3577 (N_3577,N_3018,N_2812);
nand U3578 (N_3578,N_3116,N_3168);
or U3579 (N_3579,N_3117,N_2833);
xnor U3580 (N_3580,N_3122,N_2954);
nand U3581 (N_3581,N_3097,N_3135);
or U3582 (N_3582,N_2942,N_2941);
and U3583 (N_3583,N_2977,N_2862);
nand U3584 (N_3584,N_3085,N_2912);
xnor U3585 (N_3585,N_2993,N_3117);
xor U3586 (N_3586,N_2816,N_2895);
nor U3587 (N_3587,N_2913,N_2874);
and U3588 (N_3588,N_2964,N_2930);
nand U3589 (N_3589,N_3157,N_2887);
or U3590 (N_3590,N_2820,N_3020);
or U3591 (N_3591,N_2928,N_3124);
nand U3592 (N_3592,N_2893,N_2938);
nand U3593 (N_3593,N_3142,N_2993);
xor U3594 (N_3594,N_2853,N_2966);
nor U3595 (N_3595,N_2968,N_3089);
or U3596 (N_3596,N_3060,N_2856);
and U3597 (N_3597,N_3071,N_2813);
nand U3598 (N_3598,N_2852,N_3018);
xor U3599 (N_3599,N_2893,N_2923);
or U3600 (N_3600,N_3339,N_3320);
xnor U3601 (N_3601,N_3562,N_3228);
nand U3602 (N_3602,N_3356,N_3210);
or U3603 (N_3603,N_3520,N_3256);
or U3604 (N_3604,N_3472,N_3371);
nand U3605 (N_3605,N_3357,N_3461);
and U3606 (N_3606,N_3515,N_3566);
nor U3607 (N_3607,N_3572,N_3418);
nand U3608 (N_3608,N_3502,N_3442);
nand U3609 (N_3609,N_3259,N_3488);
nor U3610 (N_3610,N_3550,N_3582);
and U3611 (N_3611,N_3401,N_3290);
xnor U3612 (N_3612,N_3263,N_3523);
or U3613 (N_3613,N_3402,N_3473);
or U3614 (N_3614,N_3456,N_3241);
nor U3615 (N_3615,N_3432,N_3574);
nor U3616 (N_3616,N_3245,N_3340);
or U3617 (N_3617,N_3318,N_3467);
and U3618 (N_3618,N_3492,N_3338);
nand U3619 (N_3619,N_3355,N_3407);
nand U3620 (N_3620,N_3301,N_3203);
nor U3621 (N_3621,N_3552,N_3380);
xnor U3622 (N_3622,N_3466,N_3229);
and U3623 (N_3623,N_3501,N_3490);
or U3624 (N_3624,N_3565,N_3253);
nand U3625 (N_3625,N_3348,N_3496);
and U3626 (N_3626,N_3494,N_3400);
nor U3627 (N_3627,N_3462,N_3249);
nand U3628 (N_3628,N_3555,N_3266);
xnor U3629 (N_3629,N_3262,N_3570);
xnor U3630 (N_3630,N_3531,N_3248);
and U3631 (N_3631,N_3378,N_3399);
or U3632 (N_3632,N_3469,N_3295);
xor U3633 (N_3633,N_3573,N_3584);
nand U3634 (N_3634,N_3351,N_3436);
nand U3635 (N_3635,N_3302,N_3423);
nor U3636 (N_3636,N_3445,N_3200);
nand U3637 (N_3637,N_3592,N_3597);
and U3638 (N_3638,N_3571,N_3403);
xor U3639 (N_3639,N_3451,N_3580);
nor U3640 (N_3640,N_3453,N_3590);
nand U3641 (N_3641,N_3267,N_3386);
xnor U3642 (N_3642,N_3519,N_3420);
and U3643 (N_3643,N_3535,N_3376);
nor U3644 (N_3644,N_3435,N_3285);
nand U3645 (N_3645,N_3437,N_3575);
nor U3646 (N_3646,N_3491,N_3391);
xnor U3647 (N_3647,N_3223,N_3438);
nand U3648 (N_3648,N_3413,N_3329);
nand U3649 (N_3649,N_3294,N_3583);
nand U3650 (N_3650,N_3258,N_3291);
or U3651 (N_3651,N_3220,N_3206);
and U3652 (N_3652,N_3465,N_3533);
xnor U3653 (N_3653,N_3595,N_3553);
or U3654 (N_3654,N_3486,N_3449);
and U3655 (N_3655,N_3510,N_3459);
or U3656 (N_3656,N_3484,N_3460);
or U3657 (N_3657,N_3498,N_3385);
nor U3658 (N_3658,N_3325,N_3579);
nand U3659 (N_3659,N_3271,N_3541);
and U3660 (N_3660,N_3563,N_3347);
and U3661 (N_3661,N_3482,N_3361);
or U3662 (N_3662,N_3441,N_3373);
and U3663 (N_3663,N_3322,N_3489);
nand U3664 (N_3664,N_3365,N_3448);
nand U3665 (N_3665,N_3350,N_3521);
nor U3666 (N_3666,N_3543,N_3447);
nor U3667 (N_3667,N_3292,N_3260);
xor U3668 (N_3668,N_3527,N_3299);
or U3669 (N_3669,N_3327,N_3217);
xnor U3670 (N_3670,N_3560,N_3564);
or U3671 (N_3671,N_3377,N_3323);
nand U3672 (N_3672,N_3280,N_3443);
or U3673 (N_3673,N_3479,N_3336);
or U3674 (N_3674,N_3485,N_3227);
and U3675 (N_3675,N_3440,N_3216);
xnor U3676 (N_3676,N_3374,N_3547);
or U3677 (N_3677,N_3429,N_3213);
or U3678 (N_3678,N_3317,N_3414);
xnor U3679 (N_3679,N_3507,N_3589);
nand U3680 (N_3680,N_3246,N_3304);
nor U3681 (N_3681,N_3360,N_3239);
nor U3682 (N_3682,N_3556,N_3261);
or U3683 (N_3683,N_3214,N_3395);
and U3684 (N_3684,N_3549,N_3251);
nand U3685 (N_3685,N_3506,N_3289);
nor U3686 (N_3686,N_3212,N_3303);
nand U3687 (N_3687,N_3559,N_3567);
nand U3688 (N_3688,N_3421,N_3530);
nand U3689 (N_3689,N_3536,N_3593);
xor U3690 (N_3690,N_3288,N_3487);
nor U3691 (N_3691,N_3284,N_3231);
and U3692 (N_3692,N_3334,N_3450);
xnor U3693 (N_3693,N_3232,N_3305);
nor U3694 (N_3694,N_3422,N_3281);
xnor U3695 (N_3695,N_3242,N_3477);
nor U3696 (N_3696,N_3311,N_3319);
nand U3697 (N_3697,N_3298,N_3393);
or U3698 (N_3698,N_3381,N_3481);
nor U3699 (N_3699,N_3455,N_3343);
nand U3700 (N_3700,N_3276,N_3211);
xor U3701 (N_3701,N_3250,N_3369);
xor U3702 (N_3702,N_3277,N_3554);
xor U3703 (N_3703,N_3341,N_3430);
and U3704 (N_3704,N_3201,N_3204);
xnor U3705 (N_3705,N_3410,N_3500);
xor U3706 (N_3706,N_3247,N_3363);
and U3707 (N_3707,N_3537,N_3508);
xnor U3708 (N_3708,N_3480,N_3427);
nand U3709 (N_3709,N_3324,N_3254);
and U3710 (N_3710,N_3306,N_3202);
and U3711 (N_3711,N_3240,N_3208);
nor U3712 (N_3712,N_3222,N_3561);
or U3713 (N_3713,N_3342,N_3557);
and U3714 (N_3714,N_3207,N_3372);
nor U3715 (N_3715,N_3265,N_3394);
nand U3716 (N_3716,N_3300,N_3568);
or U3717 (N_3717,N_3274,N_3470);
and U3718 (N_3718,N_3383,N_3236);
and U3719 (N_3719,N_3569,N_3346);
nand U3720 (N_3720,N_3352,N_3596);
nand U3721 (N_3721,N_3364,N_3475);
xnor U3722 (N_3722,N_3517,N_3358);
or U3723 (N_3723,N_3476,N_3431);
xnor U3724 (N_3724,N_3359,N_3512);
or U3725 (N_3725,N_3599,N_3332);
nor U3726 (N_3726,N_3273,N_3296);
nor U3727 (N_3727,N_3411,N_3215);
and U3728 (N_3728,N_3349,N_3233);
or U3729 (N_3729,N_3270,N_3406);
nand U3730 (N_3730,N_3225,N_3551);
nor U3731 (N_3731,N_3457,N_3424);
and U3732 (N_3732,N_3268,N_3483);
and U3733 (N_3733,N_3416,N_3545);
and U3734 (N_3734,N_3439,N_3591);
xor U3735 (N_3735,N_3283,N_3375);
xor U3736 (N_3736,N_3243,N_3528);
nor U3737 (N_3737,N_3235,N_3272);
or U3738 (N_3738,N_3282,N_3581);
or U3739 (N_3739,N_3474,N_3587);
nand U3740 (N_3740,N_3224,N_3513);
xnor U3741 (N_3741,N_3367,N_3219);
nor U3742 (N_3742,N_3576,N_3594);
nand U3743 (N_3743,N_3514,N_3337);
nor U3744 (N_3744,N_3518,N_3412);
nand U3745 (N_3745,N_3452,N_3434);
nor U3746 (N_3746,N_3275,N_3495);
nand U3747 (N_3747,N_3390,N_3379);
xnor U3748 (N_3748,N_3586,N_3546);
xor U3749 (N_3749,N_3522,N_3396);
nand U3750 (N_3750,N_3493,N_3345);
nor U3751 (N_3751,N_3230,N_3542);
nand U3752 (N_3752,N_3331,N_3409);
nor U3753 (N_3753,N_3578,N_3511);
nand U3754 (N_3754,N_3417,N_3330);
or U3755 (N_3755,N_3588,N_3382);
nor U3756 (N_3756,N_3468,N_3252);
or U3757 (N_3757,N_3209,N_3314);
or U3758 (N_3758,N_3525,N_3279);
and U3759 (N_3759,N_3539,N_3398);
nand U3760 (N_3760,N_3454,N_3315);
nand U3761 (N_3761,N_3366,N_3505);
xor U3762 (N_3762,N_3316,N_3205);
or U3763 (N_3763,N_3548,N_3226);
or U3764 (N_3764,N_3478,N_3384);
xor U3765 (N_3765,N_3238,N_3293);
nor U3766 (N_3766,N_3297,N_3426);
xor U3767 (N_3767,N_3362,N_3464);
nand U3768 (N_3768,N_3538,N_3446);
nand U3769 (N_3769,N_3237,N_3387);
nor U3770 (N_3770,N_3264,N_3503);
and U3771 (N_3771,N_3218,N_3499);
or U3772 (N_3772,N_3344,N_3221);
xnor U3773 (N_3773,N_3368,N_3310);
xor U3774 (N_3774,N_3544,N_3370);
nand U3775 (N_3775,N_3269,N_3255);
or U3776 (N_3776,N_3458,N_3405);
nand U3777 (N_3777,N_3326,N_3333);
and U3778 (N_3778,N_3509,N_3444);
or U3779 (N_3779,N_3524,N_3287);
xor U3780 (N_3780,N_3516,N_3234);
nand U3781 (N_3781,N_3497,N_3471);
or U3782 (N_3782,N_3353,N_3415);
or U3783 (N_3783,N_3312,N_3328);
or U3784 (N_3784,N_3526,N_3397);
and U3785 (N_3785,N_3308,N_3532);
nand U3786 (N_3786,N_3354,N_3585);
nand U3787 (N_3787,N_3504,N_3335);
or U3788 (N_3788,N_3534,N_3425);
nand U3789 (N_3789,N_3529,N_3463);
nor U3790 (N_3790,N_3389,N_3278);
nand U3791 (N_3791,N_3577,N_3313);
nor U3792 (N_3792,N_3388,N_3419);
and U3793 (N_3793,N_3286,N_3598);
and U3794 (N_3794,N_3244,N_3257);
and U3795 (N_3795,N_3392,N_3540);
nor U3796 (N_3796,N_3433,N_3404);
xnor U3797 (N_3797,N_3558,N_3309);
nand U3798 (N_3798,N_3321,N_3408);
or U3799 (N_3799,N_3428,N_3307);
and U3800 (N_3800,N_3288,N_3304);
xnor U3801 (N_3801,N_3582,N_3354);
and U3802 (N_3802,N_3320,N_3311);
or U3803 (N_3803,N_3396,N_3592);
nor U3804 (N_3804,N_3318,N_3217);
xor U3805 (N_3805,N_3476,N_3549);
xor U3806 (N_3806,N_3237,N_3406);
nor U3807 (N_3807,N_3471,N_3590);
nor U3808 (N_3808,N_3455,N_3435);
or U3809 (N_3809,N_3413,N_3383);
nand U3810 (N_3810,N_3424,N_3221);
or U3811 (N_3811,N_3453,N_3268);
or U3812 (N_3812,N_3265,N_3309);
xor U3813 (N_3813,N_3421,N_3236);
nand U3814 (N_3814,N_3502,N_3293);
or U3815 (N_3815,N_3581,N_3445);
nor U3816 (N_3816,N_3555,N_3293);
or U3817 (N_3817,N_3231,N_3222);
nor U3818 (N_3818,N_3232,N_3280);
xnor U3819 (N_3819,N_3582,N_3504);
or U3820 (N_3820,N_3527,N_3265);
and U3821 (N_3821,N_3421,N_3560);
nor U3822 (N_3822,N_3473,N_3529);
xor U3823 (N_3823,N_3537,N_3469);
xor U3824 (N_3824,N_3492,N_3226);
nor U3825 (N_3825,N_3406,N_3385);
and U3826 (N_3826,N_3410,N_3300);
or U3827 (N_3827,N_3547,N_3372);
nor U3828 (N_3828,N_3331,N_3428);
and U3829 (N_3829,N_3478,N_3503);
xnor U3830 (N_3830,N_3425,N_3271);
nor U3831 (N_3831,N_3294,N_3422);
nor U3832 (N_3832,N_3242,N_3354);
nor U3833 (N_3833,N_3268,N_3539);
nand U3834 (N_3834,N_3583,N_3335);
nand U3835 (N_3835,N_3321,N_3546);
nor U3836 (N_3836,N_3309,N_3591);
or U3837 (N_3837,N_3329,N_3443);
xnor U3838 (N_3838,N_3366,N_3428);
xnor U3839 (N_3839,N_3562,N_3232);
nor U3840 (N_3840,N_3308,N_3232);
nor U3841 (N_3841,N_3590,N_3413);
nor U3842 (N_3842,N_3479,N_3343);
or U3843 (N_3843,N_3420,N_3480);
xnor U3844 (N_3844,N_3214,N_3488);
nand U3845 (N_3845,N_3474,N_3211);
or U3846 (N_3846,N_3296,N_3319);
and U3847 (N_3847,N_3231,N_3558);
or U3848 (N_3848,N_3309,N_3256);
and U3849 (N_3849,N_3236,N_3538);
nor U3850 (N_3850,N_3438,N_3429);
nor U3851 (N_3851,N_3219,N_3305);
or U3852 (N_3852,N_3219,N_3362);
and U3853 (N_3853,N_3216,N_3514);
and U3854 (N_3854,N_3303,N_3267);
nor U3855 (N_3855,N_3498,N_3340);
nand U3856 (N_3856,N_3345,N_3289);
or U3857 (N_3857,N_3361,N_3348);
and U3858 (N_3858,N_3562,N_3515);
or U3859 (N_3859,N_3593,N_3364);
xor U3860 (N_3860,N_3440,N_3394);
or U3861 (N_3861,N_3411,N_3409);
xor U3862 (N_3862,N_3304,N_3368);
xor U3863 (N_3863,N_3568,N_3383);
and U3864 (N_3864,N_3493,N_3420);
nor U3865 (N_3865,N_3351,N_3337);
nor U3866 (N_3866,N_3494,N_3574);
xor U3867 (N_3867,N_3372,N_3488);
or U3868 (N_3868,N_3285,N_3319);
or U3869 (N_3869,N_3457,N_3326);
xnor U3870 (N_3870,N_3415,N_3213);
or U3871 (N_3871,N_3436,N_3238);
or U3872 (N_3872,N_3506,N_3262);
nand U3873 (N_3873,N_3417,N_3490);
xnor U3874 (N_3874,N_3575,N_3580);
xnor U3875 (N_3875,N_3507,N_3519);
xnor U3876 (N_3876,N_3399,N_3421);
nand U3877 (N_3877,N_3209,N_3288);
nand U3878 (N_3878,N_3466,N_3388);
and U3879 (N_3879,N_3526,N_3472);
nor U3880 (N_3880,N_3544,N_3452);
nor U3881 (N_3881,N_3350,N_3246);
and U3882 (N_3882,N_3554,N_3432);
xor U3883 (N_3883,N_3534,N_3200);
nand U3884 (N_3884,N_3524,N_3378);
xnor U3885 (N_3885,N_3427,N_3341);
nor U3886 (N_3886,N_3439,N_3232);
or U3887 (N_3887,N_3464,N_3402);
or U3888 (N_3888,N_3543,N_3277);
nor U3889 (N_3889,N_3270,N_3548);
nand U3890 (N_3890,N_3419,N_3559);
and U3891 (N_3891,N_3280,N_3460);
xnor U3892 (N_3892,N_3353,N_3308);
xnor U3893 (N_3893,N_3351,N_3327);
nor U3894 (N_3894,N_3269,N_3594);
nor U3895 (N_3895,N_3465,N_3322);
nor U3896 (N_3896,N_3491,N_3445);
xnor U3897 (N_3897,N_3585,N_3331);
nand U3898 (N_3898,N_3474,N_3305);
or U3899 (N_3899,N_3390,N_3402);
and U3900 (N_3900,N_3570,N_3340);
or U3901 (N_3901,N_3278,N_3416);
nor U3902 (N_3902,N_3582,N_3574);
and U3903 (N_3903,N_3305,N_3274);
nor U3904 (N_3904,N_3492,N_3408);
xnor U3905 (N_3905,N_3398,N_3272);
xor U3906 (N_3906,N_3513,N_3551);
and U3907 (N_3907,N_3451,N_3373);
nand U3908 (N_3908,N_3380,N_3549);
nand U3909 (N_3909,N_3534,N_3521);
nand U3910 (N_3910,N_3430,N_3230);
and U3911 (N_3911,N_3429,N_3354);
or U3912 (N_3912,N_3480,N_3327);
and U3913 (N_3913,N_3502,N_3495);
xor U3914 (N_3914,N_3579,N_3284);
nor U3915 (N_3915,N_3209,N_3279);
nand U3916 (N_3916,N_3507,N_3300);
or U3917 (N_3917,N_3386,N_3369);
nand U3918 (N_3918,N_3454,N_3250);
or U3919 (N_3919,N_3460,N_3492);
xnor U3920 (N_3920,N_3497,N_3485);
nor U3921 (N_3921,N_3272,N_3391);
or U3922 (N_3922,N_3218,N_3424);
xor U3923 (N_3923,N_3594,N_3332);
or U3924 (N_3924,N_3275,N_3440);
nor U3925 (N_3925,N_3268,N_3491);
or U3926 (N_3926,N_3424,N_3280);
xor U3927 (N_3927,N_3436,N_3489);
nor U3928 (N_3928,N_3439,N_3578);
nand U3929 (N_3929,N_3465,N_3571);
or U3930 (N_3930,N_3334,N_3506);
or U3931 (N_3931,N_3422,N_3383);
xor U3932 (N_3932,N_3439,N_3300);
xor U3933 (N_3933,N_3312,N_3516);
or U3934 (N_3934,N_3387,N_3223);
xor U3935 (N_3935,N_3306,N_3506);
xnor U3936 (N_3936,N_3427,N_3273);
and U3937 (N_3937,N_3351,N_3547);
nand U3938 (N_3938,N_3348,N_3436);
nor U3939 (N_3939,N_3578,N_3483);
and U3940 (N_3940,N_3523,N_3500);
and U3941 (N_3941,N_3323,N_3389);
xnor U3942 (N_3942,N_3347,N_3495);
nand U3943 (N_3943,N_3540,N_3526);
or U3944 (N_3944,N_3514,N_3369);
nor U3945 (N_3945,N_3291,N_3367);
nand U3946 (N_3946,N_3340,N_3545);
nand U3947 (N_3947,N_3591,N_3246);
and U3948 (N_3948,N_3595,N_3473);
nor U3949 (N_3949,N_3373,N_3426);
nand U3950 (N_3950,N_3327,N_3336);
nand U3951 (N_3951,N_3274,N_3583);
xnor U3952 (N_3952,N_3264,N_3371);
nor U3953 (N_3953,N_3540,N_3447);
and U3954 (N_3954,N_3558,N_3403);
and U3955 (N_3955,N_3327,N_3532);
xnor U3956 (N_3956,N_3508,N_3246);
xnor U3957 (N_3957,N_3403,N_3436);
nor U3958 (N_3958,N_3450,N_3575);
nand U3959 (N_3959,N_3580,N_3545);
nor U3960 (N_3960,N_3502,N_3335);
and U3961 (N_3961,N_3296,N_3370);
nand U3962 (N_3962,N_3455,N_3591);
nand U3963 (N_3963,N_3215,N_3201);
or U3964 (N_3964,N_3434,N_3466);
nand U3965 (N_3965,N_3566,N_3555);
nand U3966 (N_3966,N_3370,N_3463);
nand U3967 (N_3967,N_3231,N_3253);
and U3968 (N_3968,N_3303,N_3432);
or U3969 (N_3969,N_3440,N_3376);
and U3970 (N_3970,N_3514,N_3352);
or U3971 (N_3971,N_3540,N_3559);
xnor U3972 (N_3972,N_3504,N_3420);
or U3973 (N_3973,N_3544,N_3398);
nor U3974 (N_3974,N_3505,N_3549);
or U3975 (N_3975,N_3584,N_3578);
nor U3976 (N_3976,N_3350,N_3423);
nand U3977 (N_3977,N_3448,N_3337);
nand U3978 (N_3978,N_3534,N_3311);
and U3979 (N_3979,N_3209,N_3353);
xor U3980 (N_3980,N_3518,N_3238);
nand U3981 (N_3981,N_3260,N_3211);
nand U3982 (N_3982,N_3593,N_3567);
nand U3983 (N_3983,N_3236,N_3439);
nand U3984 (N_3984,N_3338,N_3247);
nor U3985 (N_3985,N_3309,N_3359);
or U3986 (N_3986,N_3206,N_3599);
and U3987 (N_3987,N_3586,N_3508);
and U3988 (N_3988,N_3362,N_3228);
nand U3989 (N_3989,N_3289,N_3510);
nand U3990 (N_3990,N_3565,N_3418);
nand U3991 (N_3991,N_3532,N_3384);
and U3992 (N_3992,N_3493,N_3408);
nor U3993 (N_3993,N_3482,N_3472);
nor U3994 (N_3994,N_3266,N_3575);
or U3995 (N_3995,N_3510,N_3444);
nand U3996 (N_3996,N_3546,N_3487);
nor U3997 (N_3997,N_3516,N_3381);
xor U3998 (N_3998,N_3559,N_3355);
nor U3999 (N_3999,N_3531,N_3332);
xnor U4000 (N_4000,N_3659,N_3705);
xor U4001 (N_4001,N_3862,N_3614);
and U4002 (N_4002,N_3927,N_3835);
xor U4003 (N_4003,N_3724,N_3609);
nand U4004 (N_4004,N_3980,N_3848);
xnor U4005 (N_4005,N_3839,N_3982);
and U4006 (N_4006,N_3718,N_3865);
nor U4007 (N_4007,N_3843,N_3920);
xnor U4008 (N_4008,N_3624,N_3880);
xor U4009 (N_4009,N_3756,N_3825);
nand U4010 (N_4010,N_3611,N_3665);
and U4011 (N_4011,N_3969,N_3988);
or U4012 (N_4012,N_3677,N_3966);
xor U4013 (N_4013,N_3890,N_3671);
and U4014 (N_4014,N_3815,N_3783);
xnor U4015 (N_4015,N_3853,N_3902);
nor U4016 (N_4016,N_3951,N_3745);
nand U4017 (N_4017,N_3735,N_3943);
xor U4018 (N_4018,N_3607,N_3773);
xor U4019 (N_4019,N_3897,N_3791);
and U4020 (N_4020,N_3631,N_3806);
or U4021 (N_4021,N_3714,N_3940);
xnor U4022 (N_4022,N_3838,N_3716);
or U4023 (N_4023,N_3958,N_3643);
or U4024 (N_4024,N_3952,N_3680);
nor U4025 (N_4025,N_3874,N_3893);
xor U4026 (N_4026,N_3993,N_3936);
or U4027 (N_4027,N_3805,N_3775);
and U4028 (N_4028,N_3871,N_3780);
and U4029 (N_4029,N_3821,N_3983);
or U4030 (N_4030,N_3828,N_3715);
nand U4031 (N_4031,N_3733,N_3883);
xnor U4032 (N_4032,N_3987,N_3759);
xnor U4033 (N_4033,N_3700,N_3930);
nor U4034 (N_4034,N_3693,N_3931);
xor U4035 (N_4035,N_3955,N_3661);
nor U4036 (N_4036,N_3933,N_3709);
xnor U4037 (N_4037,N_3888,N_3856);
or U4038 (N_4038,N_3637,N_3689);
nand U4039 (N_4039,N_3896,N_3879);
nor U4040 (N_4040,N_3986,N_3816);
or U4041 (N_4041,N_3914,N_3663);
and U4042 (N_4042,N_3906,N_3777);
nor U4043 (N_4043,N_3687,N_3617);
xor U4044 (N_4044,N_3976,N_3907);
or U4045 (N_4045,N_3905,N_3669);
and U4046 (N_4046,N_3984,N_3970);
nand U4047 (N_4047,N_3956,N_3625);
nand U4048 (N_4048,N_3675,N_3836);
xnor U4049 (N_4049,N_3834,N_3639);
or U4050 (N_4050,N_3647,N_3918);
xnor U4051 (N_4051,N_3847,N_3863);
nand U4052 (N_4052,N_3696,N_3868);
xor U4053 (N_4053,N_3662,N_3641);
or U4054 (N_4054,N_3630,N_3842);
nand U4055 (N_4055,N_3889,N_3823);
nor U4056 (N_4056,N_3990,N_3748);
and U4057 (N_4057,N_3610,N_3939);
and U4058 (N_4058,N_3787,N_3749);
nor U4059 (N_4059,N_3997,N_3707);
xor U4060 (N_4060,N_3965,N_3796);
xnor U4061 (N_4061,N_3720,N_3899);
and U4062 (N_4062,N_3964,N_3959);
nand U4063 (N_4063,N_3795,N_3615);
nand U4064 (N_4064,N_3695,N_3672);
xor U4065 (N_4065,N_3750,N_3919);
and U4066 (N_4066,N_3845,N_3711);
nor U4067 (N_4067,N_3618,N_3992);
nor U4068 (N_4068,N_3928,N_3649);
or U4069 (N_4069,N_3870,N_3938);
and U4070 (N_4070,N_3786,N_3627);
or U4071 (N_4071,N_3797,N_3784);
and U4072 (N_4072,N_3668,N_3739);
and U4073 (N_4073,N_3638,N_3832);
nor U4074 (N_4074,N_3656,N_3894);
nand U4075 (N_4075,N_3855,N_3814);
nand U4076 (N_4076,N_3683,N_3804);
and U4077 (N_4077,N_3803,N_3728);
and U4078 (N_4078,N_3681,N_3660);
and U4079 (N_4079,N_3979,N_3690);
or U4080 (N_4080,N_3860,N_3732);
and U4081 (N_4081,N_3974,N_3658);
and U4082 (N_4082,N_3881,N_3875);
xor U4083 (N_4083,N_3721,N_3751);
or U4084 (N_4084,N_3770,N_3697);
and U4085 (N_4085,N_3717,N_3950);
nand U4086 (N_4086,N_3760,N_3606);
nor U4087 (N_4087,N_3948,N_3774);
nor U4088 (N_4088,N_3971,N_3788);
or U4089 (N_4089,N_3794,N_3736);
nand U4090 (N_4090,N_3792,N_3785);
or U4091 (N_4091,N_3674,N_3954);
nand U4092 (N_4092,N_3935,N_3692);
and U4093 (N_4093,N_3782,N_3876);
and U4094 (N_4094,N_3670,N_3781);
and U4095 (N_4095,N_3629,N_3947);
or U4096 (N_4096,N_3762,N_3912);
nor U4097 (N_4097,N_3702,N_3691);
nor U4098 (N_4098,N_3961,N_3703);
nand U4099 (N_4099,N_3813,N_3685);
xnor U4100 (N_4100,N_3613,N_3994);
nor U4101 (N_4101,N_3995,N_3667);
or U4102 (N_4102,N_3633,N_3701);
nand U4103 (N_4103,N_3651,N_3887);
and U4104 (N_4104,N_3829,N_3898);
and U4105 (N_4105,N_3758,N_3727);
nand U4106 (N_4106,N_3934,N_3867);
nand U4107 (N_4107,N_3892,N_3761);
nand U4108 (N_4108,N_3837,N_3741);
nand U4109 (N_4109,N_3650,N_3740);
nand U4110 (N_4110,N_3967,N_3981);
xor U4111 (N_4111,N_3913,N_3730);
xnor U4112 (N_4112,N_3908,N_3901);
nand U4113 (N_4113,N_3852,N_3746);
xnor U4114 (N_4114,N_3826,N_3694);
xnor U4115 (N_4115,N_3801,N_3726);
nor U4116 (N_4116,N_3957,N_3772);
and U4117 (N_4117,N_3989,N_3942);
nor U4118 (N_4118,N_3802,N_3960);
xor U4119 (N_4119,N_3771,N_3653);
and U4120 (N_4120,N_3818,N_3962);
nor U4121 (N_4121,N_3686,N_3991);
nor U4122 (N_4122,N_3657,N_3910);
and U4123 (N_4123,N_3640,N_3877);
xor U4124 (N_4124,N_3808,N_3635);
nand U4125 (N_4125,N_3642,N_3858);
and U4126 (N_4126,N_3811,N_3975);
nor U4127 (N_4127,N_3648,N_3926);
nor U4128 (N_4128,N_3623,N_3944);
or U4129 (N_4129,N_3622,N_3602);
and U4130 (N_4130,N_3820,N_3723);
xnor U4131 (N_4131,N_3904,N_3654);
nand U4132 (N_4132,N_3827,N_3619);
xor U4133 (N_4133,N_3882,N_3793);
and U4134 (N_4134,N_3753,N_3999);
and U4135 (N_4135,N_3911,N_3612);
nor U4136 (N_4136,N_3719,N_3937);
or U4137 (N_4137,N_3866,N_3699);
or U4138 (N_4138,N_3946,N_3812);
xnor U4139 (N_4139,N_3755,N_3850);
or U4140 (N_4140,N_3909,N_3810);
xor U4141 (N_4141,N_3932,N_3688);
nor U4142 (N_4142,N_3645,N_3600);
and U4143 (N_4143,N_3886,N_3953);
or U4144 (N_4144,N_3722,N_3923);
nand U4145 (N_4145,N_3620,N_3800);
nand U4146 (N_4146,N_3757,N_3632);
nor U4147 (N_4147,N_3900,N_3601);
nor U4148 (N_4148,N_3963,N_3895);
nand U4149 (N_4149,N_3830,N_3676);
xnor U4150 (N_4150,N_3731,N_3846);
nor U4151 (N_4151,N_3949,N_3608);
or U4152 (N_4152,N_3844,N_3776);
nor U4153 (N_4153,N_3752,N_3704);
or U4154 (N_4154,N_3767,N_3929);
nor U4155 (N_4155,N_3873,N_3725);
nand U4156 (N_4156,N_3744,N_3973);
nand U4157 (N_4157,N_3754,N_3605);
and U4158 (N_4158,N_3706,N_3972);
or U4159 (N_4159,N_3708,N_3790);
nand U4160 (N_4160,N_3941,N_3840);
nand U4161 (N_4161,N_3903,N_3710);
nand U4162 (N_4162,N_3678,N_3985);
nand U4163 (N_4163,N_3684,N_3636);
and U4164 (N_4164,N_3621,N_3764);
and U4165 (N_4165,N_3807,N_3859);
and U4166 (N_4166,N_3673,N_3628);
nor U4167 (N_4167,N_3778,N_3789);
nand U4168 (N_4168,N_3916,N_3779);
nor U4169 (N_4169,N_3864,N_3616);
or U4170 (N_4170,N_3833,N_3924);
and U4171 (N_4171,N_3769,N_3884);
nand U4172 (N_4172,N_3854,N_3885);
xor U4173 (N_4173,N_3646,N_3604);
xor U4174 (N_4174,N_3819,N_3798);
or U4175 (N_4175,N_3652,N_3872);
xnor U4176 (N_4176,N_3766,N_3841);
nor U4177 (N_4177,N_3738,N_3878);
nand U4178 (N_4178,N_3978,N_3664);
nor U4179 (N_4179,N_3679,N_3713);
xor U4180 (N_4180,N_3765,N_3729);
xor U4181 (N_4181,N_3666,N_3626);
nand U4182 (N_4182,N_3824,N_3998);
nand U4183 (N_4183,N_3945,N_3891);
nand U4184 (N_4184,N_3655,N_3977);
nand U4185 (N_4185,N_3768,N_3634);
nor U4186 (N_4186,N_3737,N_3809);
and U4187 (N_4187,N_3922,N_3698);
or U4188 (N_4188,N_3861,N_3869);
and U4189 (N_4189,N_3857,N_3849);
xnor U4190 (N_4190,N_3817,N_3921);
or U4191 (N_4191,N_3742,N_3822);
nor U4192 (N_4192,N_3747,N_3644);
nand U4193 (N_4193,N_3917,N_3743);
xor U4194 (N_4194,N_3763,N_3915);
nor U4195 (N_4195,N_3851,N_3831);
and U4196 (N_4196,N_3682,N_3799);
or U4197 (N_4197,N_3925,N_3734);
nor U4198 (N_4198,N_3603,N_3712);
or U4199 (N_4199,N_3996,N_3968);
nor U4200 (N_4200,N_3915,N_3779);
nand U4201 (N_4201,N_3705,N_3600);
or U4202 (N_4202,N_3696,N_3623);
or U4203 (N_4203,N_3946,N_3958);
and U4204 (N_4204,N_3943,N_3627);
and U4205 (N_4205,N_3639,N_3736);
xor U4206 (N_4206,N_3747,N_3698);
nand U4207 (N_4207,N_3857,N_3749);
nand U4208 (N_4208,N_3917,N_3763);
and U4209 (N_4209,N_3958,N_3719);
xor U4210 (N_4210,N_3601,N_3605);
or U4211 (N_4211,N_3666,N_3945);
or U4212 (N_4212,N_3882,N_3903);
or U4213 (N_4213,N_3649,N_3642);
nor U4214 (N_4214,N_3809,N_3794);
or U4215 (N_4215,N_3894,N_3920);
nor U4216 (N_4216,N_3655,N_3676);
and U4217 (N_4217,N_3957,N_3827);
and U4218 (N_4218,N_3622,N_3819);
nand U4219 (N_4219,N_3800,N_3674);
xor U4220 (N_4220,N_3686,N_3918);
and U4221 (N_4221,N_3724,N_3785);
xnor U4222 (N_4222,N_3707,N_3975);
or U4223 (N_4223,N_3925,N_3650);
nand U4224 (N_4224,N_3674,N_3952);
or U4225 (N_4225,N_3662,N_3844);
or U4226 (N_4226,N_3783,N_3875);
nor U4227 (N_4227,N_3941,N_3718);
nand U4228 (N_4228,N_3953,N_3851);
nor U4229 (N_4229,N_3639,N_3689);
nand U4230 (N_4230,N_3935,N_3695);
or U4231 (N_4231,N_3912,N_3892);
or U4232 (N_4232,N_3707,N_3723);
nor U4233 (N_4233,N_3774,N_3923);
nor U4234 (N_4234,N_3723,N_3708);
nor U4235 (N_4235,N_3959,N_3986);
or U4236 (N_4236,N_3609,N_3782);
xor U4237 (N_4237,N_3793,N_3996);
and U4238 (N_4238,N_3874,N_3907);
xnor U4239 (N_4239,N_3679,N_3653);
nand U4240 (N_4240,N_3767,N_3701);
and U4241 (N_4241,N_3622,N_3826);
or U4242 (N_4242,N_3686,N_3970);
nor U4243 (N_4243,N_3812,N_3623);
xnor U4244 (N_4244,N_3706,N_3757);
nand U4245 (N_4245,N_3687,N_3942);
or U4246 (N_4246,N_3667,N_3713);
xnor U4247 (N_4247,N_3891,N_3900);
and U4248 (N_4248,N_3982,N_3891);
and U4249 (N_4249,N_3759,N_3899);
nand U4250 (N_4250,N_3634,N_3874);
nor U4251 (N_4251,N_3613,N_3914);
xnor U4252 (N_4252,N_3976,N_3713);
nand U4253 (N_4253,N_3798,N_3606);
or U4254 (N_4254,N_3853,N_3614);
and U4255 (N_4255,N_3822,N_3909);
or U4256 (N_4256,N_3904,N_3709);
xor U4257 (N_4257,N_3716,N_3614);
and U4258 (N_4258,N_3808,N_3976);
and U4259 (N_4259,N_3994,N_3908);
xor U4260 (N_4260,N_3916,N_3664);
nand U4261 (N_4261,N_3773,N_3614);
nand U4262 (N_4262,N_3861,N_3933);
nor U4263 (N_4263,N_3650,N_3931);
xnor U4264 (N_4264,N_3931,N_3661);
nor U4265 (N_4265,N_3928,N_3869);
nand U4266 (N_4266,N_3934,N_3917);
xnor U4267 (N_4267,N_3886,N_3857);
and U4268 (N_4268,N_3762,N_3654);
or U4269 (N_4269,N_3735,N_3611);
xnor U4270 (N_4270,N_3842,N_3916);
or U4271 (N_4271,N_3908,N_3947);
nor U4272 (N_4272,N_3864,N_3788);
and U4273 (N_4273,N_3638,N_3883);
xor U4274 (N_4274,N_3696,N_3603);
or U4275 (N_4275,N_3702,N_3803);
xnor U4276 (N_4276,N_3663,N_3815);
nor U4277 (N_4277,N_3889,N_3868);
or U4278 (N_4278,N_3805,N_3939);
or U4279 (N_4279,N_3619,N_3665);
nand U4280 (N_4280,N_3715,N_3646);
xnor U4281 (N_4281,N_3755,N_3946);
xor U4282 (N_4282,N_3774,N_3927);
nand U4283 (N_4283,N_3778,N_3728);
xnor U4284 (N_4284,N_3967,N_3901);
nor U4285 (N_4285,N_3650,N_3998);
nor U4286 (N_4286,N_3791,N_3778);
xnor U4287 (N_4287,N_3832,N_3614);
xnor U4288 (N_4288,N_3945,N_3625);
and U4289 (N_4289,N_3901,N_3793);
nor U4290 (N_4290,N_3937,N_3863);
nand U4291 (N_4291,N_3697,N_3704);
xor U4292 (N_4292,N_3893,N_3865);
nor U4293 (N_4293,N_3632,N_3899);
nand U4294 (N_4294,N_3826,N_3714);
nor U4295 (N_4295,N_3771,N_3939);
or U4296 (N_4296,N_3659,N_3627);
nor U4297 (N_4297,N_3660,N_3723);
nand U4298 (N_4298,N_3758,N_3707);
nor U4299 (N_4299,N_3793,N_3778);
and U4300 (N_4300,N_3908,N_3913);
nor U4301 (N_4301,N_3744,N_3747);
or U4302 (N_4302,N_3635,N_3875);
nor U4303 (N_4303,N_3959,N_3842);
xor U4304 (N_4304,N_3793,N_3877);
or U4305 (N_4305,N_3606,N_3603);
nor U4306 (N_4306,N_3808,N_3684);
nor U4307 (N_4307,N_3918,N_3760);
nand U4308 (N_4308,N_3901,N_3688);
xor U4309 (N_4309,N_3807,N_3697);
xnor U4310 (N_4310,N_3649,N_3901);
nand U4311 (N_4311,N_3666,N_3749);
xor U4312 (N_4312,N_3712,N_3727);
nor U4313 (N_4313,N_3939,N_3908);
xor U4314 (N_4314,N_3923,N_3909);
and U4315 (N_4315,N_3993,N_3974);
xnor U4316 (N_4316,N_3621,N_3712);
nand U4317 (N_4317,N_3815,N_3686);
nor U4318 (N_4318,N_3813,N_3738);
nand U4319 (N_4319,N_3829,N_3776);
nand U4320 (N_4320,N_3755,N_3629);
and U4321 (N_4321,N_3896,N_3763);
nand U4322 (N_4322,N_3899,N_3663);
nor U4323 (N_4323,N_3873,N_3826);
nor U4324 (N_4324,N_3647,N_3723);
xnor U4325 (N_4325,N_3922,N_3928);
nand U4326 (N_4326,N_3745,N_3976);
or U4327 (N_4327,N_3739,N_3968);
and U4328 (N_4328,N_3643,N_3868);
nand U4329 (N_4329,N_3715,N_3805);
nor U4330 (N_4330,N_3939,N_3903);
or U4331 (N_4331,N_3834,N_3752);
xnor U4332 (N_4332,N_3669,N_3640);
and U4333 (N_4333,N_3898,N_3862);
nand U4334 (N_4334,N_3886,N_3950);
nand U4335 (N_4335,N_3717,N_3961);
xor U4336 (N_4336,N_3727,N_3655);
nand U4337 (N_4337,N_3844,N_3735);
or U4338 (N_4338,N_3951,N_3735);
xnor U4339 (N_4339,N_3608,N_3841);
xnor U4340 (N_4340,N_3740,N_3879);
xor U4341 (N_4341,N_3812,N_3874);
or U4342 (N_4342,N_3839,N_3887);
and U4343 (N_4343,N_3602,N_3607);
or U4344 (N_4344,N_3950,N_3913);
nor U4345 (N_4345,N_3608,N_3872);
nand U4346 (N_4346,N_3667,N_3775);
nor U4347 (N_4347,N_3881,N_3972);
or U4348 (N_4348,N_3979,N_3953);
nand U4349 (N_4349,N_3709,N_3624);
nor U4350 (N_4350,N_3800,N_3884);
xor U4351 (N_4351,N_3974,N_3726);
xor U4352 (N_4352,N_3918,N_3644);
nand U4353 (N_4353,N_3714,N_3720);
nand U4354 (N_4354,N_3669,N_3699);
or U4355 (N_4355,N_3780,N_3656);
nand U4356 (N_4356,N_3730,N_3688);
and U4357 (N_4357,N_3804,N_3914);
or U4358 (N_4358,N_3910,N_3902);
nor U4359 (N_4359,N_3797,N_3832);
nand U4360 (N_4360,N_3655,N_3662);
or U4361 (N_4361,N_3955,N_3916);
nor U4362 (N_4362,N_3937,N_3792);
and U4363 (N_4363,N_3933,N_3802);
or U4364 (N_4364,N_3715,N_3721);
nand U4365 (N_4365,N_3977,N_3986);
and U4366 (N_4366,N_3992,N_3951);
nand U4367 (N_4367,N_3716,N_3709);
or U4368 (N_4368,N_3601,N_3931);
and U4369 (N_4369,N_3985,N_3888);
or U4370 (N_4370,N_3658,N_3695);
xor U4371 (N_4371,N_3679,N_3776);
and U4372 (N_4372,N_3923,N_3686);
and U4373 (N_4373,N_3986,N_3880);
nor U4374 (N_4374,N_3725,N_3623);
or U4375 (N_4375,N_3773,N_3744);
or U4376 (N_4376,N_3845,N_3909);
and U4377 (N_4377,N_3774,N_3847);
or U4378 (N_4378,N_3915,N_3870);
or U4379 (N_4379,N_3942,N_3664);
nor U4380 (N_4380,N_3914,N_3605);
and U4381 (N_4381,N_3999,N_3972);
or U4382 (N_4382,N_3899,N_3600);
and U4383 (N_4383,N_3741,N_3815);
nor U4384 (N_4384,N_3645,N_3958);
nand U4385 (N_4385,N_3777,N_3917);
nand U4386 (N_4386,N_3873,N_3808);
and U4387 (N_4387,N_3974,N_3649);
xnor U4388 (N_4388,N_3790,N_3888);
nor U4389 (N_4389,N_3658,N_3955);
and U4390 (N_4390,N_3840,N_3992);
nand U4391 (N_4391,N_3630,N_3708);
nand U4392 (N_4392,N_3832,N_3656);
or U4393 (N_4393,N_3873,N_3779);
xnor U4394 (N_4394,N_3934,N_3746);
nand U4395 (N_4395,N_3934,N_3611);
nor U4396 (N_4396,N_3788,N_3612);
and U4397 (N_4397,N_3897,N_3845);
or U4398 (N_4398,N_3940,N_3892);
and U4399 (N_4399,N_3917,N_3955);
nor U4400 (N_4400,N_4207,N_4064);
nand U4401 (N_4401,N_4023,N_4013);
or U4402 (N_4402,N_4169,N_4165);
nor U4403 (N_4403,N_4311,N_4332);
nand U4404 (N_4404,N_4349,N_4137);
nor U4405 (N_4405,N_4095,N_4235);
or U4406 (N_4406,N_4290,N_4082);
or U4407 (N_4407,N_4373,N_4166);
xnor U4408 (N_4408,N_4371,N_4282);
or U4409 (N_4409,N_4139,N_4018);
nand U4410 (N_4410,N_4008,N_4090);
nand U4411 (N_4411,N_4312,N_4193);
xor U4412 (N_4412,N_4375,N_4047);
and U4413 (N_4413,N_4131,N_4032);
or U4414 (N_4414,N_4102,N_4106);
and U4415 (N_4415,N_4045,N_4093);
or U4416 (N_4416,N_4211,N_4161);
nor U4417 (N_4417,N_4264,N_4391);
nand U4418 (N_4418,N_4026,N_4124);
and U4419 (N_4419,N_4267,N_4020);
nor U4420 (N_4420,N_4393,N_4172);
and U4421 (N_4421,N_4119,N_4170);
or U4422 (N_4422,N_4078,N_4292);
or U4423 (N_4423,N_4209,N_4244);
nand U4424 (N_4424,N_4107,N_4214);
and U4425 (N_4425,N_4315,N_4146);
and U4426 (N_4426,N_4188,N_4380);
or U4427 (N_4427,N_4043,N_4343);
xnor U4428 (N_4428,N_4329,N_4101);
xnor U4429 (N_4429,N_4058,N_4310);
and U4430 (N_4430,N_4255,N_4394);
nor U4431 (N_4431,N_4365,N_4024);
xor U4432 (N_4432,N_4361,N_4044);
nor U4433 (N_4433,N_4347,N_4357);
nor U4434 (N_4434,N_4396,N_4189);
xnor U4435 (N_4435,N_4298,N_4208);
or U4436 (N_4436,N_4109,N_4002);
and U4437 (N_4437,N_4204,N_4021);
nor U4438 (N_4438,N_4274,N_4398);
xor U4439 (N_4439,N_4324,N_4356);
xor U4440 (N_4440,N_4141,N_4163);
and U4441 (N_4441,N_4280,N_4336);
nand U4442 (N_4442,N_4351,N_4127);
or U4443 (N_4443,N_4118,N_4073);
nor U4444 (N_4444,N_4114,N_4168);
xnor U4445 (N_4445,N_4157,N_4149);
and U4446 (N_4446,N_4245,N_4092);
or U4447 (N_4447,N_4259,N_4272);
and U4448 (N_4448,N_4216,N_4056);
xnor U4449 (N_4449,N_4300,N_4307);
and U4450 (N_4450,N_4096,N_4254);
nand U4451 (N_4451,N_4003,N_4246);
nand U4452 (N_4452,N_4194,N_4134);
nand U4453 (N_4453,N_4320,N_4089);
and U4454 (N_4454,N_4116,N_4328);
nor U4455 (N_4455,N_4221,N_4341);
xnor U4456 (N_4456,N_4293,N_4145);
nor U4457 (N_4457,N_4387,N_4385);
nand U4458 (N_4458,N_4034,N_4382);
and U4459 (N_4459,N_4010,N_4305);
nor U4460 (N_4460,N_4289,N_4130);
and U4461 (N_4461,N_4117,N_4180);
or U4462 (N_4462,N_4379,N_4253);
nand U4463 (N_4463,N_4276,N_4278);
nor U4464 (N_4464,N_4065,N_4182);
and U4465 (N_4465,N_4030,N_4012);
or U4466 (N_4466,N_4074,N_4353);
or U4467 (N_4467,N_4025,N_4242);
xor U4468 (N_4468,N_4152,N_4059);
and U4469 (N_4469,N_4196,N_4147);
nand U4470 (N_4470,N_4048,N_4346);
and U4471 (N_4471,N_4266,N_4288);
and U4472 (N_4472,N_4317,N_4386);
or U4473 (N_4473,N_4151,N_4053);
nand U4474 (N_4474,N_4110,N_4179);
nand U4475 (N_4475,N_4006,N_4279);
xor U4476 (N_4476,N_4183,N_4258);
nand U4477 (N_4477,N_4138,N_4017);
and U4478 (N_4478,N_4205,N_4212);
or U4479 (N_4479,N_4286,N_4055);
nor U4480 (N_4480,N_4173,N_4014);
nor U4481 (N_4481,N_4036,N_4140);
xor U4482 (N_4482,N_4222,N_4233);
nand U4483 (N_4483,N_4041,N_4031);
and U4484 (N_4484,N_4178,N_4142);
xnor U4485 (N_4485,N_4084,N_4094);
nand U4486 (N_4486,N_4303,N_4306);
nand U4487 (N_4487,N_4304,N_4384);
xor U4488 (N_4488,N_4285,N_4225);
nand U4489 (N_4489,N_4228,N_4085);
xnor U4490 (N_4490,N_4252,N_4129);
or U4491 (N_4491,N_4348,N_4372);
nand U4492 (N_4492,N_4144,N_4389);
or U4493 (N_4493,N_4067,N_4281);
nand U4494 (N_4494,N_4011,N_4197);
xnor U4495 (N_4495,N_4227,N_4123);
nand U4496 (N_4496,N_4277,N_4294);
and U4497 (N_4497,N_4072,N_4184);
or U4498 (N_4498,N_4087,N_4162);
nand U4499 (N_4499,N_4241,N_4200);
nand U4500 (N_4500,N_4007,N_4358);
and U4501 (N_4501,N_4381,N_4001);
nor U4502 (N_4502,N_4220,N_4181);
or U4503 (N_4503,N_4238,N_4125);
nand U4504 (N_4504,N_4248,N_4203);
nor U4505 (N_4505,N_4399,N_4037);
and U4506 (N_4506,N_4344,N_4360);
and U4507 (N_4507,N_4316,N_4345);
nand U4508 (N_4508,N_4273,N_4370);
or U4509 (N_4509,N_4326,N_4148);
nor U4510 (N_4510,N_4230,N_4236);
and U4511 (N_4511,N_4318,N_4201);
and U4512 (N_4512,N_4088,N_4283);
and U4513 (N_4513,N_4042,N_4190);
xnor U4514 (N_4514,N_4263,N_4378);
and U4515 (N_4515,N_4052,N_4257);
and U4516 (N_4516,N_4135,N_4340);
nand U4517 (N_4517,N_4120,N_4261);
nand U4518 (N_4518,N_4226,N_4070);
xnor U4519 (N_4519,N_4249,N_4210);
nand U4520 (N_4520,N_4362,N_4066);
nand U4521 (N_4521,N_4218,N_4076);
nor U4522 (N_4522,N_4260,N_4080);
or U4523 (N_4523,N_4251,N_4167);
or U4524 (N_4524,N_4097,N_4215);
nand U4525 (N_4525,N_4035,N_4395);
and U4526 (N_4526,N_4219,N_4327);
nor U4527 (N_4527,N_4105,N_4319);
or U4528 (N_4528,N_4158,N_4313);
or U4529 (N_4529,N_4062,N_4295);
nand U4530 (N_4530,N_4213,N_4038);
or U4531 (N_4531,N_4126,N_4063);
nand U4532 (N_4532,N_4268,N_4022);
nor U4533 (N_4533,N_4359,N_4027);
nand U4534 (N_4534,N_4186,N_4104);
and U4535 (N_4535,N_4330,N_4150);
nor U4536 (N_4536,N_4176,N_4355);
and U4537 (N_4537,N_4171,N_4217);
nor U4538 (N_4538,N_4061,N_4111);
nand U4539 (N_4539,N_4103,N_4051);
nand U4540 (N_4540,N_4206,N_4185);
or U4541 (N_4541,N_4247,N_4291);
nor U4542 (N_4542,N_4079,N_4337);
xnor U4543 (N_4543,N_4029,N_4335);
xor U4544 (N_4544,N_4367,N_4083);
nor U4545 (N_4545,N_4374,N_4269);
nand U4546 (N_4546,N_4239,N_4050);
and U4547 (N_4547,N_4339,N_4308);
nor U4548 (N_4548,N_4069,N_4377);
and U4549 (N_4549,N_4071,N_4115);
and U4550 (N_4550,N_4302,N_4363);
and U4551 (N_4551,N_4091,N_4271);
nor U4552 (N_4552,N_4350,N_4231);
or U4553 (N_4553,N_4174,N_4077);
and U4554 (N_4554,N_4270,N_4392);
xnor U4555 (N_4555,N_4331,N_4364);
and U4556 (N_4556,N_4376,N_4046);
nor U4557 (N_4557,N_4195,N_4160);
and U4558 (N_4558,N_4154,N_4342);
nor U4559 (N_4559,N_4287,N_4301);
and U4560 (N_4560,N_4175,N_4250);
and U4561 (N_4561,N_4132,N_4325);
nor U4562 (N_4562,N_4243,N_4033);
xnor U4563 (N_4563,N_4297,N_4128);
nand U4564 (N_4564,N_4322,N_4296);
nand U4565 (N_4565,N_4019,N_4314);
or U4566 (N_4566,N_4198,N_4000);
or U4567 (N_4567,N_4122,N_4005);
or U4568 (N_4568,N_4156,N_4113);
or U4569 (N_4569,N_4309,N_4199);
and U4570 (N_4570,N_4323,N_4112);
and U4571 (N_4571,N_4159,N_4040);
xnor U4572 (N_4572,N_4081,N_4098);
nor U4573 (N_4573,N_4368,N_4155);
nor U4574 (N_4574,N_4334,N_4234);
nor U4575 (N_4575,N_4192,N_4240);
and U4576 (N_4576,N_4100,N_4237);
and U4577 (N_4577,N_4153,N_4039);
nor U4578 (N_4578,N_4229,N_4054);
xor U4579 (N_4579,N_4202,N_4338);
nand U4580 (N_4580,N_4369,N_4028);
and U4581 (N_4581,N_4224,N_4354);
nor U4582 (N_4582,N_4352,N_4015);
or U4583 (N_4583,N_4133,N_4086);
nor U4584 (N_4584,N_4136,N_4121);
or U4585 (N_4585,N_4388,N_4223);
nand U4586 (N_4586,N_4321,N_4060);
nand U4587 (N_4587,N_4390,N_4383);
nor U4588 (N_4588,N_4299,N_4187);
xor U4589 (N_4589,N_4108,N_4397);
and U4590 (N_4590,N_4284,N_4164);
xnor U4591 (N_4591,N_4099,N_4256);
nand U4592 (N_4592,N_4275,N_4177);
nand U4593 (N_4593,N_4143,N_4009);
xnor U4594 (N_4594,N_4265,N_4068);
xor U4595 (N_4595,N_4191,N_4016);
nor U4596 (N_4596,N_4232,N_4262);
xor U4597 (N_4597,N_4049,N_4366);
xnor U4598 (N_4598,N_4004,N_4057);
and U4599 (N_4599,N_4333,N_4075);
nor U4600 (N_4600,N_4212,N_4091);
or U4601 (N_4601,N_4319,N_4037);
xor U4602 (N_4602,N_4165,N_4261);
or U4603 (N_4603,N_4312,N_4135);
or U4604 (N_4604,N_4193,N_4059);
nand U4605 (N_4605,N_4034,N_4241);
and U4606 (N_4606,N_4284,N_4136);
and U4607 (N_4607,N_4315,N_4393);
and U4608 (N_4608,N_4060,N_4279);
or U4609 (N_4609,N_4004,N_4141);
and U4610 (N_4610,N_4131,N_4224);
and U4611 (N_4611,N_4147,N_4088);
and U4612 (N_4612,N_4098,N_4339);
nand U4613 (N_4613,N_4306,N_4199);
or U4614 (N_4614,N_4232,N_4282);
nor U4615 (N_4615,N_4150,N_4384);
xnor U4616 (N_4616,N_4083,N_4375);
or U4617 (N_4617,N_4075,N_4310);
nor U4618 (N_4618,N_4151,N_4169);
nand U4619 (N_4619,N_4316,N_4135);
nor U4620 (N_4620,N_4235,N_4375);
nor U4621 (N_4621,N_4283,N_4037);
and U4622 (N_4622,N_4216,N_4290);
xor U4623 (N_4623,N_4093,N_4357);
nand U4624 (N_4624,N_4217,N_4225);
nand U4625 (N_4625,N_4015,N_4182);
and U4626 (N_4626,N_4248,N_4191);
or U4627 (N_4627,N_4317,N_4102);
nor U4628 (N_4628,N_4071,N_4133);
or U4629 (N_4629,N_4291,N_4200);
xnor U4630 (N_4630,N_4141,N_4181);
xor U4631 (N_4631,N_4240,N_4293);
xnor U4632 (N_4632,N_4383,N_4109);
xor U4633 (N_4633,N_4184,N_4183);
or U4634 (N_4634,N_4130,N_4057);
nor U4635 (N_4635,N_4227,N_4064);
nand U4636 (N_4636,N_4325,N_4116);
nand U4637 (N_4637,N_4143,N_4261);
nor U4638 (N_4638,N_4349,N_4387);
nand U4639 (N_4639,N_4176,N_4293);
nor U4640 (N_4640,N_4107,N_4339);
or U4641 (N_4641,N_4133,N_4132);
xnor U4642 (N_4642,N_4103,N_4054);
nor U4643 (N_4643,N_4081,N_4361);
nor U4644 (N_4644,N_4148,N_4329);
nor U4645 (N_4645,N_4064,N_4055);
nor U4646 (N_4646,N_4123,N_4362);
or U4647 (N_4647,N_4226,N_4177);
or U4648 (N_4648,N_4041,N_4085);
and U4649 (N_4649,N_4100,N_4088);
xnor U4650 (N_4650,N_4034,N_4143);
nand U4651 (N_4651,N_4037,N_4121);
and U4652 (N_4652,N_4341,N_4020);
nor U4653 (N_4653,N_4327,N_4248);
or U4654 (N_4654,N_4344,N_4220);
or U4655 (N_4655,N_4015,N_4202);
and U4656 (N_4656,N_4354,N_4063);
nor U4657 (N_4657,N_4096,N_4297);
nor U4658 (N_4658,N_4029,N_4220);
nand U4659 (N_4659,N_4103,N_4023);
or U4660 (N_4660,N_4266,N_4066);
or U4661 (N_4661,N_4384,N_4113);
and U4662 (N_4662,N_4114,N_4052);
and U4663 (N_4663,N_4028,N_4029);
nor U4664 (N_4664,N_4285,N_4384);
xor U4665 (N_4665,N_4351,N_4092);
nand U4666 (N_4666,N_4370,N_4241);
and U4667 (N_4667,N_4202,N_4356);
nand U4668 (N_4668,N_4297,N_4292);
or U4669 (N_4669,N_4389,N_4048);
xnor U4670 (N_4670,N_4191,N_4372);
and U4671 (N_4671,N_4246,N_4099);
nand U4672 (N_4672,N_4060,N_4288);
nand U4673 (N_4673,N_4133,N_4310);
xnor U4674 (N_4674,N_4029,N_4249);
xor U4675 (N_4675,N_4131,N_4203);
or U4676 (N_4676,N_4330,N_4196);
nand U4677 (N_4677,N_4074,N_4047);
and U4678 (N_4678,N_4277,N_4093);
xnor U4679 (N_4679,N_4282,N_4005);
or U4680 (N_4680,N_4323,N_4322);
nor U4681 (N_4681,N_4194,N_4298);
nand U4682 (N_4682,N_4360,N_4063);
xor U4683 (N_4683,N_4140,N_4136);
and U4684 (N_4684,N_4080,N_4290);
and U4685 (N_4685,N_4056,N_4201);
nor U4686 (N_4686,N_4368,N_4032);
nor U4687 (N_4687,N_4264,N_4357);
and U4688 (N_4688,N_4010,N_4324);
xnor U4689 (N_4689,N_4153,N_4176);
xor U4690 (N_4690,N_4268,N_4290);
or U4691 (N_4691,N_4296,N_4139);
or U4692 (N_4692,N_4044,N_4240);
nand U4693 (N_4693,N_4206,N_4313);
nor U4694 (N_4694,N_4082,N_4354);
nor U4695 (N_4695,N_4131,N_4098);
or U4696 (N_4696,N_4050,N_4228);
or U4697 (N_4697,N_4044,N_4253);
and U4698 (N_4698,N_4364,N_4168);
xnor U4699 (N_4699,N_4245,N_4108);
nand U4700 (N_4700,N_4158,N_4078);
or U4701 (N_4701,N_4049,N_4299);
nand U4702 (N_4702,N_4340,N_4363);
nand U4703 (N_4703,N_4168,N_4176);
nor U4704 (N_4704,N_4373,N_4380);
or U4705 (N_4705,N_4372,N_4168);
or U4706 (N_4706,N_4208,N_4078);
xnor U4707 (N_4707,N_4035,N_4163);
nand U4708 (N_4708,N_4360,N_4267);
and U4709 (N_4709,N_4280,N_4192);
nand U4710 (N_4710,N_4183,N_4341);
and U4711 (N_4711,N_4077,N_4293);
nor U4712 (N_4712,N_4020,N_4241);
or U4713 (N_4713,N_4095,N_4246);
or U4714 (N_4714,N_4222,N_4309);
xnor U4715 (N_4715,N_4011,N_4357);
and U4716 (N_4716,N_4362,N_4234);
or U4717 (N_4717,N_4207,N_4196);
nand U4718 (N_4718,N_4105,N_4000);
nor U4719 (N_4719,N_4064,N_4146);
or U4720 (N_4720,N_4085,N_4120);
or U4721 (N_4721,N_4190,N_4179);
nor U4722 (N_4722,N_4006,N_4098);
nand U4723 (N_4723,N_4088,N_4154);
or U4724 (N_4724,N_4006,N_4138);
nand U4725 (N_4725,N_4287,N_4356);
xor U4726 (N_4726,N_4328,N_4337);
and U4727 (N_4727,N_4144,N_4209);
xnor U4728 (N_4728,N_4369,N_4398);
or U4729 (N_4729,N_4088,N_4135);
nor U4730 (N_4730,N_4170,N_4265);
xor U4731 (N_4731,N_4123,N_4266);
xnor U4732 (N_4732,N_4121,N_4193);
nand U4733 (N_4733,N_4349,N_4212);
and U4734 (N_4734,N_4047,N_4162);
xor U4735 (N_4735,N_4269,N_4050);
and U4736 (N_4736,N_4272,N_4075);
nor U4737 (N_4737,N_4129,N_4118);
nand U4738 (N_4738,N_4161,N_4128);
nor U4739 (N_4739,N_4039,N_4332);
or U4740 (N_4740,N_4019,N_4058);
nor U4741 (N_4741,N_4006,N_4296);
xor U4742 (N_4742,N_4097,N_4230);
and U4743 (N_4743,N_4162,N_4398);
xor U4744 (N_4744,N_4375,N_4131);
or U4745 (N_4745,N_4025,N_4174);
nand U4746 (N_4746,N_4289,N_4194);
or U4747 (N_4747,N_4396,N_4043);
nor U4748 (N_4748,N_4196,N_4237);
and U4749 (N_4749,N_4057,N_4285);
nor U4750 (N_4750,N_4316,N_4121);
xnor U4751 (N_4751,N_4156,N_4105);
nand U4752 (N_4752,N_4081,N_4315);
and U4753 (N_4753,N_4355,N_4190);
nand U4754 (N_4754,N_4330,N_4139);
and U4755 (N_4755,N_4059,N_4249);
nand U4756 (N_4756,N_4393,N_4372);
nor U4757 (N_4757,N_4010,N_4005);
nor U4758 (N_4758,N_4239,N_4001);
nand U4759 (N_4759,N_4191,N_4249);
nand U4760 (N_4760,N_4255,N_4178);
xor U4761 (N_4761,N_4221,N_4002);
nor U4762 (N_4762,N_4090,N_4030);
and U4763 (N_4763,N_4363,N_4190);
or U4764 (N_4764,N_4103,N_4028);
and U4765 (N_4765,N_4044,N_4048);
nor U4766 (N_4766,N_4276,N_4051);
and U4767 (N_4767,N_4047,N_4365);
nand U4768 (N_4768,N_4293,N_4378);
and U4769 (N_4769,N_4261,N_4025);
or U4770 (N_4770,N_4058,N_4105);
nor U4771 (N_4771,N_4062,N_4041);
or U4772 (N_4772,N_4190,N_4116);
nand U4773 (N_4773,N_4076,N_4181);
or U4774 (N_4774,N_4390,N_4009);
nor U4775 (N_4775,N_4195,N_4031);
or U4776 (N_4776,N_4372,N_4121);
nand U4777 (N_4777,N_4344,N_4160);
nand U4778 (N_4778,N_4252,N_4083);
nor U4779 (N_4779,N_4233,N_4057);
or U4780 (N_4780,N_4151,N_4321);
nand U4781 (N_4781,N_4382,N_4243);
nand U4782 (N_4782,N_4165,N_4128);
or U4783 (N_4783,N_4385,N_4094);
or U4784 (N_4784,N_4389,N_4170);
nor U4785 (N_4785,N_4112,N_4203);
xnor U4786 (N_4786,N_4089,N_4145);
or U4787 (N_4787,N_4079,N_4197);
xor U4788 (N_4788,N_4344,N_4224);
nand U4789 (N_4789,N_4090,N_4074);
xnor U4790 (N_4790,N_4368,N_4078);
or U4791 (N_4791,N_4333,N_4134);
xnor U4792 (N_4792,N_4339,N_4342);
nand U4793 (N_4793,N_4203,N_4146);
nor U4794 (N_4794,N_4267,N_4110);
or U4795 (N_4795,N_4177,N_4332);
xnor U4796 (N_4796,N_4164,N_4111);
and U4797 (N_4797,N_4288,N_4360);
nor U4798 (N_4798,N_4207,N_4186);
nand U4799 (N_4799,N_4123,N_4337);
xor U4800 (N_4800,N_4400,N_4736);
or U4801 (N_4801,N_4459,N_4746);
and U4802 (N_4802,N_4521,N_4714);
xor U4803 (N_4803,N_4616,N_4756);
nor U4804 (N_4804,N_4611,N_4495);
nand U4805 (N_4805,N_4791,N_4608);
nor U4806 (N_4806,N_4769,N_4476);
nand U4807 (N_4807,N_4457,N_4525);
and U4808 (N_4808,N_4653,N_4477);
or U4809 (N_4809,N_4593,N_4543);
xnor U4810 (N_4810,N_4579,N_4681);
or U4811 (N_4811,N_4700,N_4526);
and U4812 (N_4812,N_4581,N_4564);
nor U4813 (N_4813,N_4503,N_4505);
nor U4814 (N_4814,N_4677,N_4698);
and U4815 (N_4815,N_4435,N_4721);
nor U4816 (N_4816,N_4654,N_4410);
nor U4817 (N_4817,N_4604,N_4491);
nand U4818 (N_4818,N_4662,N_4461);
xor U4819 (N_4819,N_4790,N_4587);
and U4820 (N_4820,N_4530,N_4730);
nor U4821 (N_4821,N_4613,N_4414);
xnor U4822 (N_4822,N_4742,N_4538);
or U4823 (N_4823,N_4515,N_4633);
nand U4824 (N_4824,N_4501,N_4462);
xnor U4825 (N_4825,N_4549,N_4446);
and U4826 (N_4826,N_4518,N_4404);
and U4827 (N_4827,N_4517,N_4552);
xnor U4828 (N_4828,N_4561,N_4719);
nand U4829 (N_4829,N_4559,N_4431);
nand U4830 (N_4830,N_4718,N_4738);
nand U4831 (N_4831,N_4488,N_4539);
xnor U4832 (N_4832,N_4733,N_4689);
nor U4833 (N_4833,N_4782,N_4522);
xnor U4834 (N_4834,N_4666,N_4475);
nand U4835 (N_4835,N_4694,N_4785);
nand U4836 (N_4836,N_4486,N_4553);
or U4837 (N_4837,N_4743,N_4565);
or U4838 (N_4838,N_4695,N_4487);
and U4839 (N_4839,N_4720,N_4766);
and U4840 (N_4840,N_4643,N_4509);
and U4841 (N_4841,N_4418,N_4607);
or U4842 (N_4842,N_4433,N_4444);
xor U4843 (N_4843,N_4734,N_4612);
or U4844 (N_4844,N_4661,N_4499);
nand U4845 (N_4845,N_4760,N_4532);
nor U4846 (N_4846,N_4649,N_4603);
and U4847 (N_4847,N_4678,N_4508);
or U4848 (N_4848,N_4440,N_4696);
or U4849 (N_4849,N_4586,N_4797);
or U4850 (N_4850,N_4659,N_4513);
xor U4851 (N_4851,N_4590,N_4749);
or U4852 (N_4852,N_4629,N_4597);
nor U4853 (N_4853,N_4789,N_4709);
and U4854 (N_4854,N_4644,N_4614);
xnor U4855 (N_4855,N_4415,N_4550);
or U4856 (N_4856,N_4413,N_4407);
and U4857 (N_4857,N_4554,N_4573);
nand U4858 (N_4858,N_4627,N_4527);
nand U4859 (N_4859,N_4406,N_4767);
and U4860 (N_4860,N_4711,N_4679);
xnor U4861 (N_4861,N_4422,N_4483);
and U4862 (N_4862,N_4596,N_4704);
and U4863 (N_4863,N_4795,N_4442);
or U4864 (N_4864,N_4408,N_4715);
or U4865 (N_4865,N_4453,N_4670);
nand U4866 (N_4866,N_4636,N_4702);
and U4867 (N_4867,N_4683,N_4535);
and U4868 (N_4868,N_4658,N_4548);
nor U4869 (N_4869,N_4570,N_4490);
and U4870 (N_4870,N_4722,N_4606);
nand U4871 (N_4871,N_4595,N_4560);
or U4872 (N_4872,N_4610,N_4676);
or U4873 (N_4873,N_4635,N_4728);
nor U4874 (N_4874,N_4656,N_4437);
nor U4875 (N_4875,N_4484,N_4725);
or U4876 (N_4876,N_4741,N_4474);
nor U4877 (N_4877,N_4545,N_4753);
or U4878 (N_4878,N_4764,N_4687);
nand U4879 (N_4879,N_4451,N_4434);
and U4880 (N_4880,N_4669,N_4726);
or U4881 (N_4881,N_4419,N_4626);
and U4882 (N_4882,N_4450,N_4786);
nand U4883 (N_4883,N_4497,N_4599);
xor U4884 (N_4884,N_4628,N_4572);
and U4885 (N_4885,N_4529,N_4655);
xnor U4886 (N_4886,N_4680,N_4426);
xor U4887 (N_4887,N_4737,N_4480);
or U4888 (N_4888,N_4438,N_4660);
nand U4889 (N_4889,N_4631,N_4624);
nor U4890 (N_4890,N_4759,N_4510);
or U4891 (N_4891,N_4690,N_4744);
xor U4892 (N_4892,N_4710,N_4411);
nor U4893 (N_4893,N_4427,N_4519);
nor U4894 (N_4894,N_4536,N_4402);
nand U4895 (N_4895,N_4555,N_4639);
and U4896 (N_4896,N_4420,N_4778);
nor U4897 (N_4897,N_4443,N_4546);
and U4898 (N_4898,N_4506,N_4657);
nand U4899 (N_4899,N_4494,N_4688);
xnor U4900 (N_4900,N_4664,N_4429);
or U4901 (N_4901,N_4470,N_4675);
xor U4902 (N_4902,N_4432,N_4617);
or U4903 (N_4903,N_4638,N_4412);
xor U4904 (N_4904,N_4605,N_4747);
nor U4905 (N_4905,N_4481,N_4699);
and U4906 (N_4906,N_4707,N_4697);
nor U4907 (N_4907,N_4528,N_4752);
nand U4908 (N_4908,N_4472,N_4641);
nand U4909 (N_4909,N_4602,N_4489);
or U4910 (N_4910,N_4534,N_4609);
nor U4911 (N_4911,N_4458,N_4703);
or U4912 (N_4912,N_4772,N_4421);
or U4913 (N_4913,N_4779,N_4493);
nor U4914 (N_4914,N_4571,N_4739);
xnor U4915 (N_4915,N_4424,N_4540);
nor U4916 (N_4916,N_4448,N_4674);
nor U4917 (N_4917,N_4511,N_4773);
or U4918 (N_4918,N_4642,N_4646);
xnor U4919 (N_4919,N_4479,N_4621);
xnor U4920 (N_4920,N_4425,N_4516);
and U4921 (N_4921,N_4682,N_4583);
nor U4922 (N_4922,N_4794,N_4575);
nor U4923 (N_4923,N_4651,N_4648);
nand U4924 (N_4924,N_4466,N_4562);
nand U4925 (N_4925,N_4547,N_4500);
nor U4926 (N_4926,N_4594,N_4632);
or U4927 (N_4927,N_4783,N_4645);
xnor U4928 (N_4928,N_4625,N_4650);
nor U4929 (N_4929,N_4622,N_4558);
nand U4930 (N_4930,N_4585,N_4598);
nor U4931 (N_4931,N_4568,N_4708);
xnor U4932 (N_4932,N_4799,N_4401);
or U4933 (N_4933,N_4620,N_4647);
xor U4934 (N_4934,N_4777,N_4724);
nor U4935 (N_4935,N_4445,N_4436);
nor U4936 (N_4936,N_4567,N_4460);
nor U4937 (N_4937,N_4672,N_4580);
nor U4938 (N_4938,N_4692,N_4531);
xor U4939 (N_4939,N_4485,N_4447);
nand U4940 (N_4940,N_4512,N_4492);
nand U4941 (N_4941,N_4471,N_4551);
nor U4942 (N_4942,N_4740,N_4478);
xor U4943 (N_4943,N_4671,N_4623);
nor U4944 (N_4944,N_4723,N_4750);
nor U4945 (N_4945,N_4463,N_4524);
nand U4946 (N_4946,N_4452,N_4667);
xnor U4947 (N_4947,N_4507,N_4589);
nor U4948 (N_4948,N_4757,N_4409);
or U4949 (N_4949,N_4751,N_4618);
or U4950 (N_4950,N_4788,N_4775);
nand U4951 (N_4951,N_4566,N_4793);
nor U4952 (N_4952,N_4584,N_4706);
nor U4953 (N_4953,N_4712,N_4504);
nand U4954 (N_4954,N_4592,N_4691);
nand U4955 (N_4955,N_4755,N_4762);
or U4956 (N_4956,N_4577,N_4533);
xor U4957 (N_4957,N_4615,N_4441);
nand U4958 (N_4958,N_4665,N_4765);
nand U4959 (N_4959,N_4482,N_4403);
xnor U4960 (N_4960,N_4473,N_4569);
nand U4961 (N_4961,N_4405,N_4582);
or U4962 (N_4962,N_4630,N_4563);
or U4963 (N_4963,N_4686,N_4784);
and U4964 (N_4964,N_4705,N_4428);
xnor U4965 (N_4965,N_4763,N_4792);
xnor U4966 (N_4966,N_4498,N_4576);
and U4967 (N_4967,N_4600,N_4557);
xor U4968 (N_4968,N_4423,N_4732);
and U4969 (N_4969,N_4717,N_4663);
or U4970 (N_4970,N_4684,N_4652);
or U4971 (N_4971,N_4464,N_4776);
and U4972 (N_4972,N_4748,N_4693);
and U4973 (N_4973,N_4601,N_4634);
nor U4974 (N_4974,N_4496,N_4640);
or U4975 (N_4975,N_4544,N_4745);
and U4976 (N_4976,N_4798,N_4465);
xnor U4977 (N_4977,N_4574,N_4469);
nor U4978 (N_4978,N_4774,N_4770);
nand U4979 (N_4979,N_4591,N_4556);
nor U4980 (N_4980,N_4619,N_4713);
or U4981 (N_4981,N_4430,N_4729);
or U4982 (N_4982,N_4754,N_4716);
nand U4983 (N_4983,N_4417,N_4456);
nand U4984 (N_4984,N_4537,N_4502);
or U4985 (N_4985,N_4588,N_4514);
and U4986 (N_4986,N_4541,N_4449);
nand U4987 (N_4987,N_4467,N_4685);
nand U4988 (N_4988,N_4701,N_4454);
nand U4989 (N_4989,N_4468,N_4758);
nand U4990 (N_4990,N_4578,N_4637);
or U4991 (N_4991,N_4523,N_4520);
or U4992 (N_4992,N_4735,N_4731);
nor U4993 (N_4993,N_4416,N_4796);
and U4994 (N_4994,N_4787,N_4761);
and U4995 (N_4995,N_4668,N_4781);
and U4996 (N_4996,N_4727,N_4455);
and U4997 (N_4997,N_4768,N_4542);
and U4998 (N_4998,N_4673,N_4780);
xor U4999 (N_4999,N_4439,N_4771);
xor U5000 (N_5000,N_4588,N_4643);
and U5001 (N_5001,N_4638,N_4494);
nand U5002 (N_5002,N_4417,N_4475);
and U5003 (N_5003,N_4425,N_4797);
xnor U5004 (N_5004,N_4506,N_4594);
xor U5005 (N_5005,N_4779,N_4744);
and U5006 (N_5006,N_4679,N_4433);
nor U5007 (N_5007,N_4418,N_4630);
or U5008 (N_5008,N_4400,N_4534);
and U5009 (N_5009,N_4410,N_4686);
xor U5010 (N_5010,N_4798,N_4505);
or U5011 (N_5011,N_4579,N_4470);
nor U5012 (N_5012,N_4411,N_4727);
and U5013 (N_5013,N_4616,N_4663);
or U5014 (N_5014,N_4680,N_4580);
xor U5015 (N_5015,N_4564,N_4721);
xnor U5016 (N_5016,N_4521,N_4411);
nand U5017 (N_5017,N_4481,N_4555);
and U5018 (N_5018,N_4503,N_4504);
nor U5019 (N_5019,N_4709,N_4706);
nand U5020 (N_5020,N_4464,N_4411);
or U5021 (N_5021,N_4468,N_4409);
xnor U5022 (N_5022,N_4744,N_4424);
nand U5023 (N_5023,N_4440,N_4780);
or U5024 (N_5024,N_4759,N_4452);
nor U5025 (N_5025,N_4546,N_4706);
nand U5026 (N_5026,N_4754,N_4798);
xor U5027 (N_5027,N_4508,N_4556);
nand U5028 (N_5028,N_4441,N_4781);
and U5029 (N_5029,N_4502,N_4521);
and U5030 (N_5030,N_4626,N_4561);
nor U5031 (N_5031,N_4723,N_4650);
and U5032 (N_5032,N_4699,N_4478);
and U5033 (N_5033,N_4607,N_4434);
xnor U5034 (N_5034,N_4771,N_4642);
nor U5035 (N_5035,N_4582,N_4780);
nor U5036 (N_5036,N_4713,N_4524);
nor U5037 (N_5037,N_4787,N_4519);
nand U5038 (N_5038,N_4575,N_4423);
and U5039 (N_5039,N_4487,N_4404);
nor U5040 (N_5040,N_4656,N_4463);
and U5041 (N_5041,N_4734,N_4552);
nor U5042 (N_5042,N_4783,N_4709);
and U5043 (N_5043,N_4659,N_4576);
or U5044 (N_5044,N_4431,N_4765);
xnor U5045 (N_5045,N_4461,N_4649);
nor U5046 (N_5046,N_4760,N_4743);
nor U5047 (N_5047,N_4527,N_4778);
or U5048 (N_5048,N_4471,N_4632);
xnor U5049 (N_5049,N_4552,N_4574);
or U5050 (N_5050,N_4493,N_4653);
and U5051 (N_5051,N_4793,N_4481);
and U5052 (N_5052,N_4684,N_4672);
and U5053 (N_5053,N_4572,N_4443);
nand U5054 (N_5054,N_4576,N_4686);
nor U5055 (N_5055,N_4424,N_4707);
nand U5056 (N_5056,N_4491,N_4472);
and U5057 (N_5057,N_4594,N_4720);
nor U5058 (N_5058,N_4687,N_4681);
nand U5059 (N_5059,N_4722,N_4745);
xnor U5060 (N_5060,N_4614,N_4578);
xor U5061 (N_5061,N_4585,N_4591);
nand U5062 (N_5062,N_4649,N_4729);
nand U5063 (N_5063,N_4674,N_4413);
and U5064 (N_5064,N_4592,N_4686);
or U5065 (N_5065,N_4796,N_4702);
and U5066 (N_5066,N_4761,N_4583);
and U5067 (N_5067,N_4711,N_4428);
xnor U5068 (N_5068,N_4659,N_4548);
nor U5069 (N_5069,N_4710,N_4555);
and U5070 (N_5070,N_4797,N_4423);
or U5071 (N_5071,N_4664,N_4469);
and U5072 (N_5072,N_4438,N_4506);
xnor U5073 (N_5073,N_4538,N_4502);
xnor U5074 (N_5074,N_4615,N_4710);
or U5075 (N_5075,N_4451,N_4688);
or U5076 (N_5076,N_4413,N_4411);
nand U5077 (N_5077,N_4620,N_4456);
nor U5078 (N_5078,N_4592,N_4439);
and U5079 (N_5079,N_4682,N_4447);
or U5080 (N_5080,N_4644,N_4415);
or U5081 (N_5081,N_4606,N_4508);
nor U5082 (N_5082,N_4772,N_4789);
nand U5083 (N_5083,N_4757,N_4494);
xor U5084 (N_5084,N_4748,N_4452);
nand U5085 (N_5085,N_4600,N_4690);
or U5086 (N_5086,N_4607,N_4683);
or U5087 (N_5087,N_4432,N_4573);
xnor U5088 (N_5088,N_4601,N_4505);
nand U5089 (N_5089,N_4446,N_4703);
xor U5090 (N_5090,N_4757,N_4724);
or U5091 (N_5091,N_4734,N_4748);
nor U5092 (N_5092,N_4544,N_4475);
nor U5093 (N_5093,N_4406,N_4673);
nor U5094 (N_5094,N_4496,N_4668);
or U5095 (N_5095,N_4632,N_4497);
or U5096 (N_5096,N_4595,N_4442);
nor U5097 (N_5097,N_4521,N_4663);
xor U5098 (N_5098,N_4781,N_4660);
nand U5099 (N_5099,N_4605,N_4435);
nand U5100 (N_5100,N_4745,N_4673);
nand U5101 (N_5101,N_4767,N_4799);
nand U5102 (N_5102,N_4601,N_4550);
nand U5103 (N_5103,N_4696,N_4785);
nand U5104 (N_5104,N_4461,N_4787);
xnor U5105 (N_5105,N_4519,N_4712);
nand U5106 (N_5106,N_4731,N_4626);
nor U5107 (N_5107,N_4504,N_4459);
nor U5108 (N_5108,N_4662,N_4783);
xor U5109 (N_5109,N_4660,N_4507);
and U5110 (N_5110,N_4657,N_4739);
or U5111 (N_5111,N_4460,N_4647);
or U5112 (N_5112,N_4717,N_4597);
nand U5113 (N_5113,N_4639,N_4439);
or U5114 (N_5114,N_4512,N_4472);
and U5115 (N_5115,N_4531,N_4671);
and U5116 (N_5116,N_4763,N_4419);
xnor U5117 (N_5117,N_4711,N_4570);
and U5118 (N_5118,N_4700,N_4745);
nand U5119 (N_5119,N_4635,N_4498);
nor U5120 (N_5120,N_4739,N_4430);
nand U5121 (N_5121,N_4719,N_4677);
nor U5122 (N_5122,N_4719,N_4479);
nor U5123 (N_5123,N_4725,N_4601);
and U5124 (N_5124,N_4751,N_4717);
or U5125 (N_5125,N_4546,N_4681);
nor U5126 (N_5126,N_4615,N_4453);
nand U5127 (N_5127,N_4520,N_4589);
nor U5128 (N_5128,N_4624,N_4460);
and U5129 (N_5129,N_4555,N_4784);
and U5130 (N_5130,N_4637,N_4495);
or U5131 (N_5131,N_4703,N_4638);
xnor U5132 (N_5132,N_4642,N_4533);
nand U5133 (N_5133,N_4726,N_4406);
xor U5134 (N_5134,N_4407,N_4714);
xor U5135 (N_5135,N_4612,N_4639);
xnor U5136 (N_5136,N_4527,N_4585);
and U5137 (N_5137,N_4491,N_4692);
and U5138 (N_5138,N_4508,N_4716);
nor U5139 (N_5139,N_4519,N_4560);
and U5140 (N_5140,N_4543,N_4526);
or U5141 (N_5141,N_4752,N_4779);
xnor U5142 (N_5142,N_4574,N_4654);
or U5143 (N_5143,N_4543,N_4538);
xnor U5144 (N_5144,N_4789,N_4581);
or U5145 (N_5145,N_4521,N_4742);
or U5146 (N_5146,N_4646,N_4695);
nor U5147 (N_5147,N_4646,N_4606);
and U5148 (N_5148,N_4415,N_4719);
or U5149 (N_5149,N_4488,N_4684);
nor U5150 (N_5150,N_4636,N_4626);
xnor U5151 (N_5151,N_4645,N_4481);
and U5152 (N_5152,N_4508,N_4707);
nand U5153 (N_5153,N_4470,N_4533);
or U5154 (N_5154,N_4622,N_4431);
xnor U5155 (N_5155,N_4785,N_4488);
and U5156 (N_5156,N_4712,N_4693);
nand U5157 (N_5157,N_4513,N_4515);
or U5158 (N_5158,N_4503,N_4436);
nand U5159 (N_5159,N_4648,N_4609);
and U5160 (N_5160,N_4647,N_4793);
xnor U5161 (N_5161,N_4698,N_4797);
nand U5162 (N_5162,N_4531,N_4419);
nand U5163 (N_5163,N_4507,N_4596);
nand U5164 (N_5164,N_4667,N_4686);
and U5165 (N_5165,N_4457,N_4678);
and U5166 (N_5166,N_4696,N_4414);
nand U5167 (N_5167,N_4734,N_4578);
and U5168 (N_5168,N_4710,N_4729);
xnor U5169 (N_5169,N_4739,N_4680);
nand U5170 (N_5170,N_4571,N_4563);
xnor U5171 (N_5171,N_4521,N_4459);
and U5172 (N_5172,N_4597,N_4645);
nand U5173 (N_5173,N_4468,N_4510);
nor U5174 (N_5174,N_4465,N_4450);
or U5175 (N_5175,N_4528,N_4580);
or U5176 (N_5176,N_4740,N_4730);
nand U5177 (N_5177,N_4542,N_4567);
or U5178 (N_5178,N_4599,N_4441);
and U5179 (N_5179,N_4571,N_4548);
nand U5180 (N_5180,N_4748,N_4621);
nor U5181 (N_5181,N_4633,N_4435);
nor U5182 (N_5182,N_4498,N_4568);
nand U5183 (N_5183,N_4444,N_4672);
nand U5184 (N_5184,N_4404,N_4634);
nand U5185 (N_5185,N_4619,N_4465);
xnor U5186 (N_5186,N_4713,N_4621);
nand U5187 (N_5187,N_4446,N_4535);
nand U5188 (N_5188,N_4629,N_4661);
nand U5189 (N_5189,N_4511,N_4687);
or U5190 (N_5190,N_4673,N_4590);
nor U5191 (N_5191,N_4607,N_4494);
nor U5192 (N_5192,N_4540,N_4486);
or U5193 (N_5193,N_4444,N_4754);
nor U5194 (N_5194,N_4600,N_4466);
nor U5195 (N_5195,N_4563,N_4475);
nand U5196 (N_5196,N_4737,N_4571);
or U5197 (N_5197,N_4575,N_4576);
and U5198 (N_5198,N_4647,N_4661);
xor U5199 (N_5199,N_4478,N_4600);
or U5200 (N_5200,N_5014,N_5116);
nand U5201 (N_5201,N_5131,N_4824);
or U5202 (N_5202,N_5135,N_5149);
nor U5203 (N_5203,N_5099,N_4840);
or U5204 (N_5204,N_5119,N_5081);
and U5205 (N_5205,N_5147,N_4977);
and U5206 (N_5206,N_4879,N_4914);
or U5207 (N_5207,N_5185,N_4911);
xnor U5208 (N_5208,N_5106,N_5006);
nor U5209 (N_5209,N_5065,N_5176);
and U5210 (N_5210,N_5007,N_4934);
nand U5211 (N_5211,N_5017,N_4995);
nor U5212 (N_5212,N_5186,N_4820);
nand U5213 (N_5213,N_5151,N_5000);
nand U5214 (N_5214,N_5023,N_4945);
nor U5215 (N_5215,N_5002,N_5182);
nor U5216 (N_5216,N_4916,N_4936);
and U5217 (N_5217,N_4876,N_5127);
or U5218 (N_5218,N_4954,N_5087);
nor U5219 (N_5219,N_4851,N_5112);
or U5220 (N_5220,N_5097,N_5180);
or U5221 (N_5221,N_4984,N_5100);
or U5222 (N_5222,N_4882,N_5168);
xor U5223 (N_5223,N_5030,N_4816);
and U5224 (N_5224,N_5189,N_4947);
and U5225 (N_5225,N_5161,N_4929);
nor U5226 (N_5226,N_5059,N_4933);
or U5227 (N_5227,N_4819,N_4969);
nand U5228 (N_5228,N_5040,N_4894);
or U5229 (N_5229,N_4861,N_4839);
and U5230 (N_5230,N_5067,N_5073);
and U5231 (N_5231,N_4921,N_5029);
and U5232 (N_5232,N_5039,N_4843);
nor U5233 (N_5233,N_5034,N_5046);
and U5234 (N_5234,N_4932,N_5193);
or U5235 (N_5235,N_5041,N_4910);
or U5236 (N_5236,N_4973,N_5146);
nand U5237 (N_5237,N_5120,N_5139);
and U5238 (N_5238,N_5062,N_4908);
xor U5239 (N_5239,N_4983,N_4884);
nand U5240 (N_5240,N_5092,N_4847);
or U5241 (N_5241,N_4918,N_4880);
nor U5242 (N_5242,N_5128,N_5166);
or U5243 (N_5243,N_5118,N_4842);
or U5244 (N_5244,N_5078,N_5110);
nand U5245 (N_5245,N_5152,N_5033);
or U5246 (N_5246,N_5077,N_4868);
and U5247 (N_5247,N_5082,N_5058);
xor U5248 (N_5248,N_5187,N_5133);
xnor U5249 (N_5249,N_5153,N_4896);
xor U5250 (N_5250,N_4900,N_4972);
or U5251 (N_5251,N_5072,N_5107);
or U5252 (N_5252,N_5155,N_5032);
or U5253 (N_5253,N_5143,N_4986);
nor U5254 (N_5254,N_4808,N_4817);
nor U5255 (N_5255,N_5194,N_5031);
nand U5256 (N_5256,N_4885,N_4821);
or U5257 (N_5257,N_4804,N_4965);
nor U5258 (N_5258,N_5080,N_5096);
and U5259 (N_5259,N_4962,N_4993);
and U5260 (N_5260,N_5008,N_4828);
or U5261 (N_5261,N_4811,N_4987);
nor U5262 (N_5262,N_5057,N_4889);
or U5263 (N_5263,N_5148,N_4937);
nand U5264 (N_5264,N_4991,N_4940);
or U5265 (N_5265,N_5113,N_4800);
or U5266 (N_5266,N_4836,N_5157);
and U5267 (N_5267,N_5095,N_4814);
nor U5268 (N_5268,N_5083,N_4830);
nand U5269 (N_5269,N_5132,N_5156);
xnor U5270 (N_5270,N_5124,N_4812);
nor U5271 (N_5271,N_4938,N_4871);
or U5272 (N_5272,N_4975,N_4943);
nand U5273 (N_5273,N_5011,N_5198);
and U5274 (N_5274,N_5104,N_4873);
or U5275 (N_5275,N_4810,N_4970);
or U5276 (N_5276,N_4854,N_4905);
or U5277 (N_5277,N_4951,N_4849);
nand U5278 (N_5278,N_4961,N_5145);
xnor U5279 (N_5279,N_5190,N_5012);
nand U5280 (N_5280,N_5136,N_5159);
nand U5281 (N_5281,N_4834,N_5121);
nand U5282 (N_5282,N_5044,N_4858);
nor U5283 (N_5283,N_5084,N_5091);
xnor U5284 (N_5284,N_5004,N_5009);
nand U5285 (N_5285,N_5089,N_5027);
and U5286 (N_5286,N_4890,N_5042);
and U5287 (N_5287,N_5137,N_4926);
or U5288 (N_5288,N_5043,N_5162);
or U5289 (N_5289,N_5129,N_4928);
nor U5290 (N_5290,N_5010,N_5169);
and U5291 (N_5291,N_4907,N_5050);
xor U5292 (N_5292,N_5098,N_4815);
nand U5293 (N_5293,N_5158,N_5114);
xnor U5294 (N_5294,N_5045,N_4952);
xor U5295 (N_5295,N_5024,N_4957);
or U5296 (N_5296,N_4902,N_4872);
nand U5297 (N_5297,N_5195,N_4801);
and U5298 (N_5298,N_5049,N_4992);
nor U5299 (N_5299,N_5142,N_5115);
or U5300 (N_5300,N_4831,N_4924);
xor U5301 (N_5301,N_5074,N_5093);
nand U5302 (N_5302,N_4895,N_5102);
xnor U5303 (N_5303,N_4838,N_4920);
or U5304 (N_5304,N_4856,N_5015);
or U5305 (N_5305,N_5079,N_5154);
nand U5306 (N_5306,N_5150,N_5177);
nor U5307 (N_5307,N_4837,N_4866);
nor U5308 (N_5308,N_5060,N_4930);
nor U5309 (N_5309,N_4967,N_4877);
nor U5310 (N_5310,N_5160,N_4848);
and U5311 (N_5311,N_4950,N_5178);
xor U5312 (N_5312,N_5140,N_4845);
and U5313 (N_5313,N_4818,N_5013);
xor U5314 (N_5314,N_5164,N_4974);
or U5315 (N_5315,N_4982,N_5105);
xor U5316 (N_5316,N_4979,N_4886);
xor U5317 (N_5317,N_5175,N_5076);
xor U5318 (N_5318,N_5064,N_4941);
nand U5319 (N_5319,N_5191,N_4939);
nand U5320 (N_5320,N_4852,N_5141);
xor U5321 (N_5321,N_5163,N_4988);
nor U5322 (N_5322,N_4917,N_4953);
nand U5323 (N_5323,N_5019,N_5199);
xor U5324 (N_5324,N_4981,N_5184);
and U5325 (N_5325,N_4963,N_4985);
or U5326 (N_5326,N_5109,N_4809);
and U5327 (N_5327,N_4825,N_4935);
nand U5328 (N_5328,N_4862,N_4925);
and U5329 (N_5329,N_5101,N_4959);
xor U5330 (N_5330,N_5181,N_4853);
xnor U5331 (N_5331,N_4922,N_4878);
or U5332 (N_5332,N_4826,N_4960);
or U5333 (N_5333,N_4802,N_4913);
xor U5334 (N_5334,N_5111,N_4841);
xor U5335 (N_5335,N_4996,N_5068);
or U5336 (N_5336,N_5167,N_5171);
or U5337 (N_5337,N_5056,N_4846);
and U5338 (N_5338,N_5173,N_4906);
nand U5339 (N_5339,N_4942,N_5170);
nor U5340 (N_5340,N_5090,N_5126);
or U5341 (N_5341,N_5052,N_5048);
nand U5342 (N_5342,N_5053,N_5003);
nand U5343 (N_5343,N_4860,N_4859);
xor U5344 (N_5344,N_5108,N_4844);
and U5345 (N_5345,N_4897,N_5016);
or U5346 (N_5346,N_4822,N_4813);
nor U5347 (N_5347,N_5134,N_4833);
and U5348 (N_5348,N_5138,N_4999);
xnor U5349 (N_5349,N_5086,N_4806);
xor U5350 (N_5350,N_5021,N_4971);
nand U5351 (N_5351,N_4870,N_4887);
or U5352 (N_5352,N_5103,N_4998);
xor U5353 (N_5353,N_5066,N_4874);
xnor U5354 (N_5354,N_4966,N_4903);
nor U5355 (N_5355,N_5125,N_4956);
nor U5356 (N_5356,N_4955,N_4835);
nand U5357 (N_5357,N_4915,N_4865);
nand U5358 (N_5358,N_5085,N_5005);
nor U5359 (N_5359,N_4948,N_5188);
and U5360 (N_5360,N_4823,N_4864);
or U5361 (N_5361,N_5020,N_5071);
or U5362 (N_5362,N_5037,N_5130);
nor U5363 (N_5363,N_5088,N_5075);
nor U5364 (N_5364,N_5094,N_4989);
or U5365 (N_5365,N_5069,N_5122);
nand U5366 (N_5366,N_5051,N_4893);
nor U5367 (N_5367,N_5063,N_4881);
nand U5368 (N_5368,N_5196,N_4899);
and U5369 (N_5369,N_5192,N_4931);
and U5370 (N_5370,N_4869,N_5183);
nor U5371 (N_5371,N_4863,N_5117);
or U5372 (N_5372,N_4912,N_4832);
nor U5373 (N_5373,N_4946,N_4997);
nand U5374 (N_5374,N_5055,N_4949);
xnor U5375 (N_5375,N_4976,N_4964);
xnor U5376 (N_5376,N_5179,N_5165);
nand U5377 (N_5377,N_4805,N_5047);
or U5378 (N_5378,N_4923,N_4909);
xor U5379 (N_5379,N_4867,N_4807);
nor U5380 (N_5380,N_4855,N_5018);
xor U5381 (N_5381,N_4829,N_4827);
or U5382 (N_5382,N_4892,N_4904);
and U5383 (N_5383,N_4968,N_5035);
xor U5384 (N_5384,N_5070,N_5038);
nor U5385 (N_5385,N_5036,N_5174);
nor U5386 (N_5386,N_4901,N_4803);
nor U5387 (N_5387,N_4898,N_4919);
xnor U5388 (N_5388,N_5144,N_5001);
and U5389 (N_5389,N_5123,N_4980);
xor U5390 (N_5390,N_5172,N_5022);
nand U5391 (N_5391,N_4978,N_4888);
xor U5392 (N_5392,N_5061,N_5197);
and U5393 (N_5393,N_4857,N_5025);
nand U5394 (N_5394,N_5054,N_4994);
nor U5395 (N_5395,N_5026,N_4850);
nand U5396 (N_5396,N_4891,N_4883);
and U5397 (N_5397,N_4990,N_5028);
xor U5398 (N_5398,N_4944,N_4927);
xor U5399 (N_5399,N_4958,N_4875);
nor U5400 (N_5400,N_4913,N_5112);
and U5401 (N_5401,N_4917,N_4815);
or U5402 (N_5402,N_4822,N_4949);
and U5403 (N_5403,N_5072,N_5145);
nand U5404 (N_5404,N_5028,N_4947);
xor U5405 (N_5405,N_4950,N_4965);
nand U5406 (N_5406,N_4834,N_5123);
or U5407 (N_5407,N_5113,N_5061);
and U5408 (N_5408,N_5127,N_5055);
or U5409 (N_5409,N_4841,N_5021);
and U5410 (N_5410,N_4957,N_5197);
nor U5411 (N_5411,N_5146,N_5157);
xor U5412 (N_5412,N_5156,N_4984);
nor U5413 (N_5413,N_4925,N_5175);
or U5414 (N_5414,N_4859,N_5077);
nor U5415 (N_5415,N_5030,N_4909);
nand U5416 (N_5416,N_5091,N_4974);
nor U5417 (N_5417,N_4901,N_4834);
xor U5418 (N_5418,N_4862,N_5102);
and U5419 (N_5419,N_4801,N_5073);
nor U5420 (N_5420,N_4864,N_4987);
and U5421 (N_5421,N_4992,N_4881);
xnor U5422 (N_5422,N_5083,N_4892);
nor U5423 (N_5423,N_4857,N_5096);
nand U5424 (N_5424,N_5153,N_5084);
nor U5425 (N_5425,N_4936,N_5112);
or U5426 (N_5426,N_4811,N_5070);
nor U5427 (N_5427,N_5148,N_5013);
and U5428 (N_5428,N_4804,N_5011);
and U5429 (N_5429,N_4813,N_5098);
nor U5430 (N_5430,N_4892,N_4886);
nand U5431 (N_5431,N_4981,N_4987);
nand U5432 (N_5432,N_5039,N_5034);
and U5433 (N_5433,N_4949,N_5106);
and U5434 (N_5434,N_5068,N_4902);
and U5435 (N_5435,N_5003,N_4834);
or U5436 (N_5436,N_4853,N_5125);
nor U5437 (N_5437,N_4977,N_5174);
nor U5438 (N_5438,N_5078,N_5196);
xor U5439 (N_5439,N_5119,N_4832);
xnor U5440 (N_5440,N_5194,N_4847);
and U5441 (N_5441,N_5165,N_5194);
xnor U5442 (N_5442,N_5004,N_5041);
xor U5443 (N_5443,N_5027,N_5199);
nand U5444 (N_5444,N_4802,N_4956);
nor U5445 (N_5445,N_5013,N_5184);
or U5446 (N_5446,N_4803,N_5067);
xor U5447 (N_5447,N_4990,N_5130);
nor U5448 (N_5448,N_4905,N_4968);
and U5449 (N_5449,N_4967,N_5012);
and U5450 (N_5450,N_5157,N_5172);
xnor U5451 (N_5451,N_4855,N_4963);
and U5452 (N_5452,N_4917,N_5112);
and U5453 (N_5453,N_5032,N_4985);
or U5454 (N_5454,N_4807,N_5093);
and U5455 (N_5455,N_5132,N_4927);
and U5456 (N_5456,N_5118,N_4861);
xnor U5457 (N_5457,N_5183,N_5047);
nor U5458 (N_5458,N_4988,N_4939);
or U5459 (N_5459,N_5118,N_4925);
or U5460 (N_5460,N_4810,N_5167);
nand U5461 (N_5461,N_4827,N_4943);
nor U5462 (N_5462,N_4922,N_5082);
nand U5463 (N_5463,N_4937,N_5161);
xnor U5464 (N_5464,N_5125,N_5167);
or U5465 (N_5465,N_4952,N_4994);
nand U5466 (N_5466,N_5140,N_5072);
nor U5467 (N_5467,N_4851,N_5145);
nor U5468 (N_5468,N_5099,N_4839);
and U5469 (N_5469,N_5123,N_4988);
or U5470 (N_5470,N_4800,N_4835);
and U5471 (N_5471,N_4961,N_4846);
nor U5472 (N_5472,N_4914,N_4961);
xor U5473 (N_5473,N_5170,N_4812);
and U5474 (N_5474,N_5177,N_5020);
or U5475 (N_5475,N_5122,N_5083);
nand U5476 (N_5476,N_5169,N_4832);
or U5477 (N_5477,N_4929,N_4892);
nor U5478 (N_5478,N_5091,N_4884);
nor U5479 (N_5479,N_4866,N_4831);
or U5480 (N_5480,N_5131,N_4947);
and U5481 (N_5481,N_5153,N_5131);
xor U5482 (N_5482,N_4996,N_5000);
nor U5483 (N_5483,N_4907,N_5056);
and U5484 (N_5484,N_5091,N_4811);
nor U5485 (N_5485,N_4871,N_4887);
and U5486 (N_5486,N_4989,N_4876);
xnor U5487 (N_5487,N_5004,N_4949);
nor U5488 (N_5488,N_4951,N_4979);
xnor U5489 (N_5489,N_4881,N_4886);
and U5490 (N_5490,N_5152,N_4801);
xnor U5491 (N_5491,N_4826,N_5055);
xor U5492 (N_5492,N_5175,N_4825);
nor U5493 (N_5493,N_5016,N_4875);
nor U5494 (N_5494,N_4998,N_4881);
and U5495 (N_5495,N_4995,N_5006);
xor U5496 (N_5496,N_4821,N_5162);
nand U5497 (N_5497,N_4891,N_4952);
or U5498 (N_5498,N_5080,N_4954);
xnor U5499 (N_5499,N_4968,N_4944);
xor U5500 (N_5500,N_5085,N_5186);
xor U5501 (N_5501,N_4807,N_5045);
xor U5502 (N_5502,N_4910,N_4854);
nor U5503 (N_5503,N_4829,N_5043);
nand U5504 (N_5504,N_4820,N_4909);
nand U5505 (N_5505,N_4872,N_5058);
nand U5506 (N_5506,N_5171,N_5094);
and U5507 (N_5507,N_4868,N_5170);
nand U5508 (N_5508,N_5039,N_5092);
nor U5509 (N_5509,N_4992,N_5129);
xnor U5510 (N_5510,N_5126,N_5061);
and U5511 (N_5511,N_5084,N_5077);
nand U5512 (N_5512,N_4841,N_5134);
nor U5513 (N_5513,N_4937,N_5100);
nand U5514 (N_5514,N_4846,N_5051);
nor U5515 (N_5515,N_4947,N_5198);
xor U5516 (N_5516,N_5052,N_4808);
nand U5517 (N_5517,N_5114,N_4835);
and U5518 (N_5518,N_5199,N_4902);
or U5519 (N_5519,N_4903,N_4854);
xor U5520 (N_5520,N_5130,N_5036);
nand U5521 (N_5521,N_4822,N_4948);
nand U5522 (N_5522,N_4963,N_5162);
and U5523 (N_5523,N_4959,N_4973);
nand U5524 (N_5524,N_4894,N_5115);
or U5525 (N_5525,N_4858,N_5147);
nor U5526 (N_5526,N_4933,N_5128);
xor U5527 (N_5527,N_5161,N_4862);
nor U5528 (N_5528,N_5130,N_4972);
and U5529 (N_5529,N_5062,N_5104);
nand U5530 (N_5530,N_5142,N_4905);
xor U5531 (N_5531,N_5178,N_4872);
nand U5532 (N_5532,N_4974,N_4848);
and U5533 (N_5533,N_4839,N_5065);
and U5534 (N_5534,N_5069,N_4947);
nor U5535 (N_5535,N_5166,N_4890);
or U5536 (N_5536,N_5116,N_5186);
nor U5537 (N_5537,N_5135,N_4876);
and U5538 (N_5538,N_4924,N_5182);
nand U5539 (N_5539,N_4833,N_4841);
nor U5540 (N_5540,N_4912,N_5108);
and U5541 (N_5541,N_5130,N_5149);
nor U5542 (N_5542,N_5026,N_5156);
nor U5543 (N_5543,N_4990,N_5193);
or U5544 (N_5544,N_4879,N_4866);
xnor U5545 (N_5545,N_4832,N_5091);
and U5546 (N_5546,N_4817,N_5184);
and U5547 (N_5547,N_5101,N_5078);
xor U5548 (N_5548,N_5098,N_5034);
or U5549 (N_5549,N_4846,N_4991);
and U5550 (N_5550,N_4846,N_4894);
nor U5551 (N_5551,N_5140,N_4933);
or U5552 (N_5552,N_4823,N_4822);
or U5553 (N_5553,N_4851,N_4918);
xor U5554 (N_5554,N_5159,N_5116);
nand U5555 (N_5555,N_5059,N_4944);
nand U5556 (N_5556,N_4979,N_5118);
nor U5557 (N_5557,N_4949,N_4903);
nand U5558 (N_5558,N_4910,N_4980);
nor U5559 (N_5559,N_4954,N_5181);
xnor U5560 (N_5560,N_4801,N_4822);
and U5561 (N_5561,N_5055,N_4828);
xnor U5562 (N_5562,N_5124,N_4975);
or U5563 (N_5563,N_5026,N_4870);
or U5564 (N_5564,N_5027,N_4878);
or U5565 (N_5565,N_5060,N_4956);
or U5566 (N_5566,N_4800,N_4864);
or U5567 (N_5567,N_4883,N_5136);
and U5568 (N_5568,N_4852,N_5143);
nand U5569 (N_5569,N_5128,N_4924);
or U5570 (N_5570,N_5157,N_5131);
xor U5571 (N_5571,N_5125,N_5086);
xor U5572 (N_5572,N_5012,N_4818);
nand U5573 (N_5573,N_4822,N_5051);
and U5574 (N_5574,N_5040,N_4906);
nand U5575 (N_5575,N_5006,N_4881);
nor U5576 (N_5576,N_5096,N_4864);
nand U5577 (N_5577,N_4810,N_5039);
nand U5578 (N_5578,N_5008,N_4917);
nor U5579 (N_5579,N_5196,N_4815);
or U5580 (N_5580,N_4856,N_4976);
nor U5581 (N_5581,N_4961,N_5142);
and U5582 (N_5582,N_5094,N_5095);
nand U5583 (N_5583,N_4963,N_5177);
and U5584 (N_5584,N_5048,N_5060);
and U5585 (N_5585,N_4857,N_4845);
and U5586 (N_5586,N_5067,N_5138);
and U5587 (N_5587,N_5135,N_5068);
and U5588 (N_5588,N_5076,N_5068);
or U5589 (N_5589,N_5183,N_4822);
nor U5590 (N_5590,N_4812,N_4878);
nand U5591 (N_5591,N_5170,N_5125);
or U5592 (N_5592,N_4852,N_4859);
or U5593 (N_5593,N_5139,N_4940);
and U5594 (N_5594,N_5155,N_4905);
nand U5595 (N_5595,N_5021,N_4869);
nor U5596 (N_5596,N_5079,N_4840);
nor U5597 (N_5597,N_5134,N_4984);
nand U5598 (N_5598,N_5072,N_5033);
xor U5599 (N_5599,N_5196,N_5157);
nand U5600 (N_5600,N_5315,N_5204);
nand U5601 (N_5601,N_5376,N_5219);
xnor U5602 (N_5602,N_5276,N_5464);
nor U5603 (N_5603,N_5586,N_5458);
nand U5604 (N_5604,N_5431,N_5591);
or U5605 (N_5605,N_5382,N_5371);
nor U5606 (N_5606,N_5213,N_5413);
xor U5607 (N_5607,N_5257,N_5465);
nor U5608 (N_5608,N_5383,N_5225);
xnor U5609 (N_5609,N_5261,N_5317);
and U5610 (N_5610,N_5461,N_5214);
nor U5611 (N_5611,N_5342,N_5491);
or U5612 (N_5612,N_5557,N_5263);
and U5613 (N_5613,N_5594,N_5248);
and U5614 (N_5614,N_5488,N_5212);
xor U5615 (N_5615,N_5512,N_5332);
nor U5616 (N_5616,N_5550,N_5532);
xnor U5617 (N_5617,N_5411,N_5243);
and U5618 (N_5618,N_5242,N_5322);
xnor U5619 (N_5619,N_5504,N_5318);
nand U5620 (N_5620,N_5453,N_5426);
nand U5621 (N_5621,N_5267,N_5517);
and U5622 (N_5622,N_5279,N_5485);
and U5623 (N_5623,N_5387,N_5561);
or U5624 (N_5624,N_5294,N_5283);
and U5625 (N_5625,N_5339,N_5568);
and U5626 (N_5626,N_5447,N_5576);
nor U5627 (N_5627,N_5303,N_5200);
nor U5628 (N_5628,N_5296,N_5246);
and U5629 (N_5629,N_5285,N_5506);
or U5630 (N_5630,N_5524,N_5421);
or U5631 (N_5631,N_5265,N_5529);
xor U5632 (N_5632,N_5450,N_5521);
or U5633 (N_5633,N_5388,N_5579);
and U5634 (N_5634,N_5587,N_5410);
xor U5635 (N_5635,N_5327,N_5203);
xor U5636 (N_5636,N_5354,N_5456);
and U5637 (N_5637,N_5329,N_5425);
nand U5638 (N_5638,N_5287,N_5364);
nand U5639 (N_5639,N_5330,N_5370);
nand U5640 (N_5640,N_5406,N_5311);
or U5641 (N_5641,N_5422,N_5556);
or U5642 (N_5642,N_5384,N_5574);
and U5643 (N_5643,N_5271,N_5323);
nand U5644 (N_5644,N_5564,N_5566);
nor U5645 (N_5645,N_5588,N_5525);
nor U5646 (N_5646,N_5580,N_5560);
nor U5647 (N_5647,N_5501,N_5362);
xor U5648 (N_5648,N_5502,N_5375);
nand U5649 (N_5649,N_5215,N_5496);
and U5650 (N_5650,N_5514,N_5490);
or U5651 (N_5651,N_5221,N_5526);
nor U5652 (N_5652,N_5286,N_5408);
nor U5653 (N_5653,N_5513,N_5348);
and U5654 (N_5654,N_5433,N_5483);
or U5655 (N_5655,N_5241,N_5438);
and U5656 (N_5656,N_5310,N_5328);
or U5657 (N_5657,N_5418,N_5455);
nand U5658 (N_5658,N_5335,N_5238);
and U5659 (N_5659,N_5443,N_5533);
nand U5660 (N_5660,N_5343,N_5280);
or U5661 (N_5661,N_5227,N_5356);
xnor U5662 (N_5662,N_5585,N_5407);
nand U5663 (N_5663,N_5385,N_5252);
xnor U5664 (N_5664,N_5442,N_5218);
xor U5665 (N_5665,N_5543,N_5262);
nor U5666 (N_5666,N_5349,N_5597);
nand U5667 (N_5667,N_5309,N_5559);
or U5668 (N_5668,N_5545,N_5272);
nor U5669 (N_5669,N_5207,N_5575);
nand U5670 (N_5670,N_5444,N_5558);
and U5671 (N_5671,N_5540,N_5359);
nor U5672 (N_5672,N_5333,N_5393);
nand U5673 (N_5673,N_5487,N_5582);
xnor U5674 (N_5674,N_5222,N_5592);
or U5675 (N_5675,N_5548,N_5552);
nand U5676 (N_5676,N_5305,N_5472);
xnor U5677 (N_5677,N_5462,N_5389);
xnor U5678 (N_5678,N_5497,N_5473);
nor U5679 (N_5679,N_5205,N_5297);
nor U5680 (N_5680,N_5549,N_5381);
and U5681 (N_5681,N_5495,N_5367);
xnor U5682 (N_5682,N_5386,N_5351);
xor U5683 (N_5683,N_5350,N_5581);
xor U5684 (N_5684,N_5471,N_5454);
nand U5685 (N_5685,N_5353,N_5522);
nor U5686 (N_5686,N_5479,N_5236);
nor U5687 (N_5687,N_5520,N_5395);
and U5688 (N_5688,N_5571,N_5448);
and U5689 (N_5689,N_5449,N_5527);
or U5690 (N_5690,N_5542,N_5554);
or U5691 (N_5691,N_5292,N_5427);
and U5692 (N_5692,N_5429,N_5233);
nor U5693 (N_5693,N_5217,N_5291);
nor U5694 (N_5694,N_5230,N_5440);
xor U5695 (N_5695,N_5598,N_5331);
nor U5696 (N_5696,N_5569,N_5451);
nand U5697 (N_5697,N_5477,N_5363);
or U5698 (N_5698,N_5469,N_5249);
nor U5699 (N_5699,N_5360,N_5298);
xor U5700 (N_5700,N_5336,N_5377);
nor U5701 (N_5701,N_5255,N_5369);
xnor U5702 (N_5702,N_5211,N_5402);
and U5703 (N_5703,N_5256,N_5417);
nand U5704 (N_5704,N_5304,N_5535);
nand U5705 (N_5705,N_5264,N_5567);
and U5706 (N_5706,N_5489,N_5539);
and U5707 (N_5707,N_5345,N_5206);
and U5708 (N_5708,N_5577,N_5326);
nor U5709 (N_5709,N_5368,N_5240);
nand U5710 (N_5710,N_5401,N_5397);
xnor U5711 (N_5711,N_5480,N_5253);
or U5712 (N_5712,N_5380,N_5570);
nor U5713 (N_5713,N_5302,N_5482);
nand U5714 (N_5714,N_5234,N_5226);
xor U5715 (N_5715,N_5589,N_5365);
or U5716 (N_5716,N_5546,N_5289);
and U5717 (N_5717,N_5301,N_5424);
xor U5718 (N_5718,N_5509,N_5404);
xor U5719 (N_5719,N_5361,N_5499);
xnor U5720 (N_5720,N_5414,N_5284);
nand U5721 (N_5721,N_5434,N_5282);
nor U5722 (N_5722,N_5324,N_5593);
nor U5723 (N_5723,N_5531,N_5201);
nor U5724 (N_5724,N_5275,N_5295);
xnor U5725 (N_5725,N_5536,N_5321);
or U5726 (N_5726,N_5224,N_5366);
xor U5727 (N_5727,N_5555,N_5439);
xnor U5728 (N_5728,N_5374,N_5312);
or U5729 (N_5729,N_5270,N_5583);
nor U5730 (N_5730,N_5254,N_5538);
and U5731 (N_5731,N_5346,N_5396);
nor U5732 (N_5732,N_5416,N_5319);
and U5733 (N_5733,N_5510,N_5358);
and U5734 (N_5734,N_5278,N_5266);
and U5735 (N_5735,N_5338,N_5290);
or U5736 (N_5736,N_5306,N_5373);
xor U5737 (N_5737,N_5247,N_5273);
or U5738 (N_5738,N_5528,N_5435);
xor U5739 (N_5739,N_5596,N_5340);
and U5740 (N_5740,N_5399,N_5223);
nor U5741 (N_5741,N_5378,N_5220);
xor U5742 (N_5742,N_5511,N_5423);
nand U5743 (N_5743,N_5235,N_5352);
or U5744 (N_5744,N_5544,N_5503);
xnor U5745 (N_5745,N_5415,N_5478);
or U5746 (N_5746,N_5498,N_5379);
nor U5747 (N_5747,N_5430,N_5209);
or U5748 (N_5748,N_5541,N_5484);
xnor U5749 (N_5749,N_5460,N_5505);
xor U5750 (N_5750,N_5584,N_5563);
or U5751 (N_5751,N_5508,N_5400);
and U5752 (N_5752,N_5412,N_5258);
nor U5753 (N_5753,N_5562,N_5537);
or U5754 (N_5754,N_5534,N_5515);
nand U5755 (N_5755,N_5251,N_5507);
or U5756 (N_5756,N_5237,N_5269);
xor U5757 (N_5757,N_5347,N_5229);
nor U5758 (N_5758,N_5405,N_5551);
and U5759 (N_5759,N_5239,N_5320);
and U5760 (N_5760,N_5573,N_5578);
xnor U5761 (N_5761,N_5519,N_5516);
nor U5762 (N_5762,N_5436,N_5392);
or U5763 (N_5763,N_5390,N_5446);
and U5764 (N_5764,N_5599,N_5493);
and U5765 (N_5765,N_5547,N_5288);
nand U5766 (N_5766,N_5481,N_5409);
and U5767 (N_5767,N_5394,N_5210);
xnor U5768 (N_5768,N_5523,N_5590);
nor U5769 (N_5769,N_5277,N_5441);
nand U5770 (N_5770,N_5344,N_5391);
xnor U5771 (N_5771,N_5300,N_5403);
and U5772 (N_5772,N_5565,N_5250);
nor U5773 (N_5773,N_5445,N_5281);
and U5774 (N_5774,N_5470,N_5299);
xor U5775 (N_5775,N_5466,N_5372);
and U5776 (N_5776,N_5313,N_5492);
and U5777 (N_5777,N_5245,N_5293);
and U5778 (N_5778,N_5518,N_5231);
nor U5779 (N_5779,N_5337,N_5334);
and U5780 (N_5780,N_5457,N_5316);
xor U5781 (N_5781,N_5341,N_5474);
nor U5782 (N_5782,N_5357,N_5428);
and U5783 (N_5783,N_5398,N_5325);
and U5784 (N_5784,N_5307,N_5244);
nor U5785 (N_5785,N_5260,N_5595);
and U5786 (N_5786,N_5208,N_5216);
nand U5787 (N_5787,N_5432,N_5232);
nand U5788 (N_5788,N_5486,N_5530);
nor U5789 (N_5789,N_5468,N_5494);
nand U5790 (N_5790,N_5467,N_5475);
xor U5791 (N_5791,N_5202,N_5459);
xor U5792 (N_5792,N_5314,N_5553);
and U5793 (N_5793,N_5463,N_5420);
nand U5794 (N_5794,N_5437,N_5268);
nor U5795 (N_5795,N_5452,N_5355);
nand U5796 (N_5796,N_5259,N_5572);
or U5797 (N_5797,N_5274,N_5228);
xor U5798 (N_5798,N_5419,N_5308);
nand U5799 (N_5799,N_5500,N_5476);
nand U5800 (N_5800,N_5434,N_5413);
xor U5801 (N_5801,N_5268,N_5453);
xor U5802 (N_5802,N_5568,N_5575);
nor U5803 (N_5803,N_5254,N_5324);
nand U5804 (N_5804,N_5510,N_5235);
nor U5805 (N_5805,N_5293,N_5432);
nor U5806 (N_5806,N_5420,N_5356);
xnor U5807 (N_5807,N_5306,N_5276);
nor U5808 (N_5808,N_5248,N_5412);
nor U5809 (N_5809,N_5242,N_5249);
and U5810 (N_5810,N_5231,N_5386);
and U5811 (N_5811,N_5535,N_5377);
and U5812 (N_5812,N_5253,N_5581);
and U5813 (N_5813,N_5341,N_5422);
nand U5814 (N_5814,N_5223,N_5323);
or U5815 (N_5815,N_5298,N_5319);
nand U5816 (N_5816,N_5307,N_5227);
xor U5817 (N_5817,N_5372,N_5577);
xor U5818 (N_5818,N_5502,N_5329);
xnor U5819 (N_5819,N_5427,N_5294);
nand U5820 (N_5820,N_5304,N_5278);
nor U5821 (N_5821,N_5526,N_5425);
nor U5822 (N_5822,N_5234,N_5310);
xnor U5823 (N_5823,N_5228,N_5266);
xor U5824 (N_5824,N_5482,N_5322);
and U5825 (N_5825,N_5469,N_5538);
or U5826 (N_5826,N_5318,N_5419);
or U5827 (N_5827,N_5360,N_5248);
or U5828 (N_5828,N_5301,N_5226);
or U5829 (N_5829,N_5598,N_5373);
and U5830 (N_5830,N_5507,N_5505);
nand U5831 (N_5831,N_5297,N_5427);
and U5832 (N_5832,N_5571,N_5225);
nand U5833 (N_5833,N_5233,N_5368);
nand U5834 (N_5834,N_5297,N_5359);
nand U5835 (N_5835,N_5415,N_5457);
or U5836 (N_5836,N_5289,N_5533);
nor U5837 (N_5837,N_5215,N_5347);
xor U5838 (N_5838,N_5549,N_5258);
and U5839 (N_5839,N_5454,N_5456);
nand U5840 (N_5840,N_5552,N_5453);
and U5841 (N_5841,N_5389,N_5281);
nor U5842 (N_5842,N_5436,N_5205);
nand U5843 (N_5843,N_5478,N_5299);
and U5844 (N_5844,N_5444,N_5580);
and U5845 (N_5845,N_5594,N_5533);
nand U5846 (N_5846,N_5586,N_5221);
xor U5847 (N_5847,N_5546,N_5221);
or U5848 (N_5848,N_5204,N_5268);
and U5849 (N_5849,N_5564,N_5270);
xor U5850 (N_5850,N_5476,N_5324);
nand U5851 (N_5851,N_5393,N_5409);
xor U5852 (N_5852,N_5397,N_5247);
or U5853 (N_5853,N_5501,N_5297);
nor U5854 (N_5854,N_5372,N_5339);
or U5855 (N_5855,N_5235,N_5207);
or U5856 (N_5856,N_5435,N_5296);
and U5857 (N_5857,N_5334,N_5553);
xnor U5858 (N_5858,N_5598,N_5504);
or U5859 (N_5859,N_5516,N_5557);
or U5860 (N_5860,N_5484,N_5432);
xnor U5861 (N_5861,N_5563,N_5573);
and U5862 (N_5862,N_5218,N_5412);
and U5863 (N_5863,N_5468,N_5404);
or U5864 (N_5864,N_5598,N_5502);
nor U5865 (N_5865,N_5428,N_5324);
nor U5866 (N_5866,N_5449,N_5466);
or U5867 (N_5867,N_5408,N_5235);
and U5868 (N_5868,N_5283,N_5430);
nor U5869 (N_5869,N_5459,N_5458);
nand U5870 (N_5870,N_5482,N_5508);
or U5871 (N_5871,N_5456,N_5510);
or U5872 (N_5872,N_5289,N_5220);
or U5873 (N_5873,N_5349,N_5373);
nand U5874 (N_5874,N_5504,N_5227);
nand U5875 (N_5875,N_5524,N_5564);
and U5876 (N_5876,N_5334,N_5360);
nor U5877 (N_5877,N_5444,N_5587);
and U5878 (N_5878,N_5572,N_5203);
and U5879 (N_5879,N_5498,N_5243);
nand U5880 (N_5880,N_5356,N_5258);
nor U5881 (N_5881,N_5253,N_5475);
nand U5882 (N_5882,N_5517,N_5521);
nand U5883 (N_5883,N_5379,N_5588);
xor U5884 (N_5884,N_5587,N_5561);
xnor U5885 (N_5885,N_5218,N_5335);
or U5886 (N_5886,N_5496,N_5277);
or U5887 (N_5887,N_5369,N_5386);
or U5888 (N_5888,N_5483,N_5566);
or U5889 (N_5889,N_5532,N_5490);
and U5890 (N_5890,N_5515,N_5553);
and U5891 (N_5891,N_5312,N_5367);
nand U5892 (N_5892,N_5393,N_5477);
xnor U5893 (N_5893,N_5409,N_5531);
or U5894 (N_5894,N_5472,N_5239);
or U5895 (N_5895,N_5336,N_5580);
or U5896 (N_5896,N_5344,N_5556);
nor U5897 (N_5897,N_5490,N_5574);
nand U5898 (N_5898,N_5287,N_5248);
or U5899 (N_5899,N_5255,N_5493);
xor U5900 (N_5900,N_5207,N_5439);
and U5901 (N_5901,N_5280,N_5442);
nor U5902 (N_5902,N_5569,N_5374);
and U5903 (N_5903,N_5580,N_5542);
and U5904 (N_5904,N_5393,N_5239);
nor U5905 (N_5905,N_5546,N_5243);
xnor U5906 (N_5906,N_5351,N_5518);
nor U5907 (N_5907,N_5416,N_5216);
or U5908 (N_5908,N_5421,N_5591);
and U5909 (N_5909,N_5543,N_5555);
or U5910 (N_5910,N_5311,N_5420);
and U5911 (N_5911,N_5571,N_5369);
or U5912 (N_5912,N_5357,N_5505);
or U5913 (N_5913,N_5587,N_5203);
and U5914 (N_5914,N_5209,N_5506);
nand U5915 (N_5915,N_5289,N_5365);
and U5916 (N_5916,N_5266,N_5535);
xor U5917 (N_5917,N_5433,N_5269);
and U5918 (N_5918,N_5268,N_5425);
and U5919 (N_5919,N_5350,N_5563);
or U5920 (N_5920,N_5330,N_5416);
or U5921 (N_5921,N_5251,N_5520);
xor U5922 (N_5922,N_5253,N_5357);
nand U5923 (N_5923,N_5313,N_5528);
or U5924 (N_5924,N_5272,N_5415);
xor U5925 (N_5925,N_5469,N_5595);
nor U5926 (N_5926,N_5281,N_5311);
xnor U5927 (N_5927,N_5300,N_5387);
nor U5928 (N_5928,N_5213,N_5543);
or U5929 (N_5929,N_5206,N_5512);
xor U5930 (N_5930,N_5391,N_5332);
or U5931 (N_5931,N_5429,N_5313);
xnor U5932 (N_5932,N_5587,N_5354);
xor U5933 (N_5933,N_5347,N_5500);
or U5934 (N_5934,N_5454,N_5369);
xnor U5935 (N_5935,N_5415,N_5598);
xor U5936 (N_5936,N_5467,N_5500);
xnor U5937 (N_5937,N_5493,N_5524);
or U5938 (N_5938,N_5470,N_5573);
nand U5939 (N_5939,N_5459,N_5292);
and U5940 (N_5940,N_5357,N_5538);
or U5941 (N_5941,N_5532,N_5515);
xor U5942 (N_5942,N_5474,N_5348);
xor U5943 (N_5943,N_5330,N_5563);
xor U5944 (N_5944,N_5248,N_5213);
nor U5945 (N_5945,N_5392,N_5210);
xor U5946 (N_5946,N_5417,N_5238);
and U5947 (N_5947,N_5388,N_5371);
and U5948 (N_5948,N_5538,N_5493);
xnor U5949 (N_5949,N_5516,N_5445);
and U5950 (N_5950,N_5475,N_5418);
nand U5951 (N_5951,N_5333,N_5448);
and U5952 (N_5952,N_5327,N_5252);
or U5953 (N_5953,N_5517,N_5306);
nor U5954 (N_5954,N_5493,N_5565);
or U5955 (N_5955,N_5256,N_5392);
or U5956 (N_5956,N_5574,N_5304);
or U5957 (N_5957,N_5599,N_5315);
nand U5958 (N_5958,N_5319,N_5557);
nor U5959 (N_5959,N_5321,N_5574);
and U5960 (N_5960,N_5492,N_5229);
and U5961 (N_5961,N_5569,N_5335);
nor U5962 (N_5962,N_5495,N_5498);
or U5963 (N_5963,N_5378,N_5223);
or U5964 (N_5964,N_5353,N_5591);
or U5965 (N_5965,N_5559,N_5334);
nor U5966 (N_5966,N_5479,N_5592);
or U5967 (N_5967,N_5331,N_5479);
xnor U5968 (N_5968,N_5424,N_5330);
nor U5969 (N_5969,N_5270,N_5579);
nand U5970 (N_5970,N_5564,N_5254);
nor U5971 (N_5971,N_5453,N_5228);
nor U5972 (N_5972,N_5364,N_5432);
or U5973 (N_5973,N_5217,N_5223);
nor U5974 (N_5974,N_5396,N_5235);
and U5975 (N_5975,N_5485,N_5389);
nand U5976 (N_5976,N_5430,N_5323);
nor U5977 (N_5977,N_5524,N_5473);
xnor U5978 (N_5978,N_5342,N_5358);
or U5979 (N_5979,N_5573,N_5576);
or U5980 (N_5980,N_5432,N_5483);
xor U5981 (N_5981,N_5290,N_5313);
xnor U5982 (N_5982,N_5585,N_5421);
and U5983 (N_5983,N_5241,N_5487);
xnor U5984 (N_5984,N_5567,N_5273);
and U5985 (N_5985,N_5211,N_5200);
nand U5986 (N_5986,N_5552,N_5289);
nand U5987 (N_5987,N_5201,N_5504);
xor U5988 (N_5988,N_5242,N_5287);
and U5989 (N_5989,N_5273,N_5537);
nor U5990 (N_5990,N_5308,N_5532);
and U5991 (N_5991,N_5282,N_5361);
nand U5992 (N_5992,N_5468,N_5590);
nor U5993 (N_5993,N_5524,N_5541);
and U5994 (N_5994,N_5447,N_5313);
nor U5995 (N_5995,N_5220,N_5459);
nor U5996 (N_5996,N_5392,N_5521);
or U5997 (N_5997,N_5388,N_5464);
nor U5998 (N_5998,N_5394,N_5253);
nor U5999 (N_5999,N_5384,N_5298);
or U6000 (N_6000,N_5669,N_5636);
nand U6001 (N_6001,N_5869,N_5897);
nor U6002 (N_6002,N_5876,N_5964);
xor U6003 (N_6003,N_5944,N_5602);
xor U6004 (N_6004,N_5683,N_5812);
or U6005 (N_6005,N_5634,N_5953);
and U6006 (N_6006,N_5748,N_5714);
xor U6007 (N_6007,N_5810,N_5735);
or U6008 (N_6008,N_5777,N_5823);
xnor U6009 (N_6009,N_5643,N_5638);
or U6010 (N_6010,N_5607,N_5807);
xnor U6011 (N_6011,N_5806,N_5771);
xor U6012 (N_6012,N_5605,N_5639);
nor U6013 (N_6013,N_5838,N_5940);
or U6014 (N_6014,N_5664,N_5929);
nor U6015 (N_6015,N_5744,N_5673);
nor U6016 (N_6016,N_5918,N_5752);
xnor U6017 (N_6017,N_5841,N_5705);
and U6018 (N_6018,N_5661,N_5837);
nand U6019 (N_6019,N_5935,N_5955);
xnor U6020 (N_6020,N_5926,N_5952);
and U6021 (N_6021,N_5624,N_5846);
or U6022 (N_6022,N_5941,N_5724);
nor U6023 (N_6023,N_5736,N_5785);
or U6024 (N_6024,N_5832,N_5781);
or U6025 (N_6025,N_5879,N_5890);
nor U6026 (N_6026,N_5889,N_5622);
and U6027 (N_6027,N_5932,N_5662);
xnor U6028 (N_6028,N_5829,N_5697);
or U6029 (N_6029,N_5759,N_5958);
nor U6030 (N_6030,N_5718,N_5779);
or U6031 (N_6031,N_5737,N_5687);
nor U6032 (N_6032,N_5977,N_5672);
or U6033 (N_6033,N_5776,N_5690);
and U6034 (N_6034,N_5853,N_5808);
or U6035 (N_6035,N_5657,N_5968);
or U6036 (N_6036,N_5908,N_5680);
or U6037 (N_6037,N_5973,N_5709);
or U6038 (N_6038,N_5763,N_5674);
nand U6039 (N_6039,N_5809,N_5725);
xor U6040 (N_6040,N_5604,N_5775);
nor U6041 (N_6041,N_5849,N_5619);
xor U6042 (N_6042,N_5970,N_5830);
xor U6043 (N_6043,N_5923,N_5706);
xnor U6044 (N_6044,N_5868,N_5627);
and U6045 (N_6045,N_5710,N_5653);
nor U6046 (N_6046,N_5915,N_5800);
and U6047 (N_6047,N_5728,N_5720);
nand U6048 (N_6048,N_5729,N_5982);
nor U6049 (N_6049,N_5787,N_5772);
nor U6050 (N_6050,N_5803,N_5642);
xor U6051 (N_6051,N_5871,N_5942);
nand U6052 (N_6052,N_5797,N_5618);
or U6053 (N_6053,N_5865,N_5962);
xnor U6054 (N_6054,N_5992,N_5663);
xnor U6055 (N_6055,N_5770,N_5997);
xnor U6056 (N_6056,N_5948,N_5640);
and U6057 (N_6057,N_5760,N_5665);
or U6058 (N_6058,N_5886,N_5991);
nor U6059 (N_6059,N_5647,N_5901);
xnor U6060 (N_6060,N_5917,N_5993);
xnor U6061 (N_6061,N_5825,N_5788);
and U6062 (N_6062,N_5857,N_5692);
and U6063 (N_6063,N_5911,N_5633);
or U6064 (N_6064,N_5701,N_5861);
nand U6065 (N_6065,N_5855,N_5954);
xnor U6066 (N_6066,N_5816,N_5924);
nor U6067 (N_6067,N_5767,N_5696);
or U6068 (N_6068,N_5721,N_5712);
or U6069 (N_6069,N_5927,N_5758);
or U6070 (N_6070,N_5761,N_5906);
nand U6071 (N_6071,N_5757,N_5983);
nand U6072 (N_6072,N_5799,N_5920);
xnor U6073 (N_6073,N_5742,N_5693);
and U6074 (N_6074,N_5684,N_5603);
xor U6075 (N_6075,N_5987,N_5996);
xnor U6076 (N_6076,N_5978,N_5883);
and U6077 (N_6077,N_5798,N_5834);
nand U6078 (N_6078,N_5668,N_5630);
nor U6079 (N_6079,N_5727,N_5854);
nor U6080 (N_6080,N_5990,N_5786);
or U6081 (N_6081,N_5621,N_5723);
nand U6082 (N_6082,N_5822,N_5681);
nor U6083 (N_6083,N_5804,N_5629);
or U6084 (N_6084,N_5717,N_5914);
and U6085 (N_6085,N_5769,N_5999);
nand U6086 (N_6086,N_5874,N_5732);
nand U6087 (N_6087,N_5998,N_5862);
nor U6088 (N_6088,N_5877,N_5780);
and U6089 (N_6089,N_5863,N_5715);
nor U6090 (N_6090,N_5898,N_5976);
nand U6091 (N_6091,N_5951,N_5766);
and U6092 (N_6092,N_5891,N_5625);
xnor U6093 (N_6093,N_5704,N_5845);
nand U6094 (N_6094,N_5824,N_5652);
or U6095 (N_6095,N_5608,N_5892);
or U6096 (N_6096,N_5610,N_5887);
and U6097 (N_6097,N_5971,N_5682);
nand U6098 (N_6098,N_5945,N_5654);
and U6099 (N_6099,N_5819,N_5694);
nand U6100 (N_6100,N_5894,N_5745);
nor U6101 (N_6101,N_5873,N_5912);
nand U6102 (N_6102,N_5677,N_5730);
xor U6103 (N_6103,N_5773,N_5922);
xnor U6104 (N_6104,N_5820,N_5979);
xnor U6105 (N_6105,N_5864,N_5660);
nor U6106 (N_6106,N_5835,N_5956);
nand U6107 (N_6107,N_5635,N_5859);
nor U6108 (N_6108,N_5994,N_5617);
nor U6109 (N_6109,N_5933,N_5880);
and U6110 (N_6110,N_5765,N_5641);
xnor U6111 (N_6111,N_5756,N_5930);
nor U6112 (N_6112,N_5826,N_5980);
or U6113 (N_6113,N_5601,N_5778);
xor U6114 (N_6114,N_5784,N_5843);
xor U6115 (N_6115,N_5811,N_5878);
nor U6116 (N_6116,N_5750,N_5919);
and U6117 (N_6117,N_5893,N_5836);
and U6118 (N_6118,N_5839,N_5913);
xor U6119 (N_6119,N_5733,N_5858);
xnor U6120 (N_6120,N_5670,N_5722);
or U6121 (N_6121,N_5972,N_5813);
xnor U6122 (N_6122,N_5910,N_5774);
xnor U6123 (N_6123,N_5611,N_5679);
or U6124 (N_6124,N_5795,N_5899);
nand U6125 (N_6125,N_5989,N_5957);
and U6126 (N_6126,N_5981,N_5632);
and U6127 (N_6127,N_5731,N_5882);
xor U6128 (N_6128,N_5699,N_5848);
and U6129 (N_6129,N_5842,N_5716);
xor U6130 (N_6130,N_5768,N_5961);
nor U6131 (N_6131,N_5614,N_5719);
nor U6132 (N_6132,N_5686,N_5844);
and U6133 (N_6133,N_5646,N_5833);
or U6134 (N_6134,N_5762,N_5792);
nand U6135 (N_6135,N_5749,N_5711);
nor U6136 (N_6136,N_5726,N_5666);
nor U6137 (N_6137,N_5675,N_5740);
xor U6138 (N_6138,N_5651,N_5609);
xor U6139 (N_6139,N_5902,N_5909);
or U6140 (N_6140,N_5975,N_5904);
or U6141 (N_6141,N_5685,N_5695);
and U6142 (N_6142,N_5995,N_5827);
nand U6143 (N_6143,N_5688,N_5631);
nand U6144 (N_6144,N_5676,N_5938);
nand U6145 (N_6145,N_5885,N_5888);
or U6146 (N_6146,N_5851,N_5821);
and U6147 (N_6147,N_5986,N_5656);
xor U6148 (N_6148,N_5649,N_5928);
nor U6149 (N_6149,N_5814,N_5950);
and U6150 (N_6150,N_5984,N_5905);
and U6151 (N_6151,N_5628,N_5739);
xor U6152 (N_6152,N_5793,N_5648);
xor U6153 (N_6153,N_5818,N_5794);
nor U6154 (N_6154,N_5671,N_5659);
nor U6155 (N_6155,N_5623,N_5626);
or U6156 (N_6156,N_5852,N_5934);
nand U6157 (N_6157,N_5612,N_5707);
nor U6158 (N_6158,N_5801,N_5616);
nor U6159 (N_6159,N_5743,N_5866);
nor U6160 (N_6160,N_5949,N_5741);
nand U6161 (N_6161,N_5700,N_5703);
xor U6162 (N_6162,N_5966,N_5606);
and U6163 (N_6163,N_5637,N_5907);
nand U6164 (N_6164,N_5734,N_5985);
nand U6165 (N_6165,N_5974,N_5847);
nand U6166 (N_6166,N_5805,N_5840);
nor U6167 (N_6167,N_5738,N_5782);
nor U6168 (N_6168,N_5791,N_5753);
xnor U6169 (N_6169,N_5796,N_5959);
xnor U6170 (N_6170,N_5658,N_5691);
or U6171 (N_6171,N_5931,N_5960);
nor U6172 (N_6172,N_5713,N_5870);
or U6173 (N_6173,N_5667,N_5947);
nand U6174 (N_6174,N_5678,N_5969);
xnor U6175 (N_6175,N_5754,N_5875);
and U6176 (N_6176,N_5815,N_5895);
xor U6177 (N_6177,N_5867,N_5689);
nand U6178 (N_6178,N_5988,N_5746);
or U6179 (N_6179,N_5620,N_5965);
and U6180 (N_6180,N_5613,N_5783);
xnor U6181 (N_6181,N_5872,N_5615);
xor U6182 (N_6182,N_5802,N_5881);
xor U6183 (N_6183,N_5790,N_5789);
nand U6184 (N_6184,N_5896,N_5764);
nor U6185 (N_6185,N_5708,N_5967);
nor U6186 (N_6186,N_5937,N_5828);
xor U6187 (N_6187,N_5946,N_5644);
or U6188 (N_6188,N_5860,N_5650);
nor U6189 (N_6189,N_5600,N_5831);
and U6190 (N_6190,N_5963,N_5916);
xnor U6191 (N_6191,N_5850,N_5936);
xor U6192 (N_6192,N_5939,N_5856);
nor U6193 (N_6193,N_5698,N_5702);
or U6194 (N_6194,N_5755,N_5655);
nand U6195 (N_6195,N_5884,N_5751);
or U6196 (N_6196,N_5817,N_5645);
or U6197 (N_6197,N_5900,N_5921);
nand U6198 (N_6198,N_5747,N_5943);
and U6199 (N_6199,N_5925,N_5903);
nor U6200 (N_6200,N_5869,N_5770);
nor U6201 (N_6201,N_5982,N_5989);
xor U6202 (N_6202,N_5609,N_5964);
xnor U6203 (N_6203,N_5971,N_5876);
nor U6204 (N_6204,N_5636,N_5962);
nor U6205 (N_6205,N_5634,N_5794);
or U6206 (N_6206,N_5721,N_5988);
nor U6207 (N_6207,N_5752,N_5757);
and U6208 (N_6208,N_5799,N_5728);
or U6209 (N_6209,N_5782,N_5828);
nand U6210 (N_6210,N_5711,N_5621);
xor U6211 (N_6211,N_5833,N_5919);
nand U6212 (N_6212,N_5723,N_5665);
and U6213 (N_6213,N_5940,N_5986);
nand U6214 (N_6214,N_5811,N_5983);
nor U6215 (N_6215,N_5876,N_5785);
and U6216 (N_6216,N_5692,N_5948);
nor U6217 (N_6217,N_5664,N_5620);
nand U6218 (N_6218,N_5639,N_5787);
xnor U6219 (N_6219,N_5870,N_5621);
xnor U6220 (N_6220,N_5708,N_5989);
and U6221 (N_6221,N_5713,N_5736);
and U6222 (N_6222,N_5945,N_5617);
or U6223 (N_6223,N_5813,N_5922);
nor U6224 (N_6224,N_5965,N_5903);
or U6225 (N_6225,N_5671,N_5769);
xnor U6226 (N_6226,N_5909,N_5840);
xnor U6227 (N_6227,N_5953,N_5927);
and U6228 (N_6228,N_5977,N_5605);
nor U6229 (N_6229,N_5772,N_5684);
or U6230 (N_6230,N_5802,N_5749);
nor U6231 (N_6231,N_5718,N_5930);
and U6232 (N_6232,N_5686,N_5765);
nor U6233 (N_6233,N_5706,N_5775);
nand U6234 (N_6234,N_5817,N_5976);
and U6235 (N_6235,N_5955,N_5872);
or U6236 (N_6236,N_5792,N_5743);
xor U6237 (N_6237,N_5818,N_5937);
nor U6238 (N_6238,N_5676,N_5685);
or U6239 (N_6239,N_5676,N_5749);
xor U6240 (N_6240,N_5835,N_5641);
xnor U6241 (N_6241,N_5972,N_5610);
xor U6242 (N_6242,N_5782,N_5986);
and U6243 (N_6243,N_5660,N_5961);
and U6244 (N_6244,N_5626,N_5644);
xor U6245 (N_6245,N_5922,N_5736);
and U6246 (N_6246,N_5713,N_5891);
xnor U6247 (N_6247,N_5905,N_5810);
xor U6248 (N_6248,N_5681,N_5858);
and U6249 (N_6249,N_5954,N_5965);
xnor U6250 (N_6250,N_5672,N_5793);
or U6251 (N_6251,N_5808,N_5718);
and U6252 (N_6252,N_5915,N_5660);
nand U6253 (N_6253,N_5952,N_5835);
nor U6254 (N_6254,N_5627,N_5672);
xnor U6255 (N_6255,N_5850,N_5869);
and U6256 (N_6256,N_5713,N_5624);
nand U6257 (N_6257,N_5691,N_5653);
or U6258 (N_6258,N_5779,N_5817);
nand U6259 (N_6259,N_5981,N_5833);
or U6260 (N_6260,N_5725,N_5701);
xor U6261 (N_6261,N_5919,N_5902);
nor U6262 (N_6262,N_5627,N_5648);
nor U6263 (N_6263,N_5708,N_5917);
and U6264 (N_6264,N_5933,N_5658);
or U6265 (N_6265,N_5694,N_5612);
nand U6266 (N_6266,N_5993,N_5675);
nor U6267 (N_6267,N_5891,N_5726);
nand U6268 (N_6268,N_5630,N_5831);
nand U6269 (N_6269,N_5903,N_5766);
nor U6270 (N_6270,N_5693,N_5904);
nand U6271 (N_6271,N_5628,N_5686);
xnor U6272 (N_6272,N_5785,N_5853);
and U6273 (N_6273,N_5623,N_5978);
and U6274 (N_6274,N_5922,N_5981);
or U6275 (N_6275,N_5847,N_5774);
or U6276 (N_6276,N_5707,N_5998);
or U6277 (N_6277,N_5951,N_5813);
nor U6278 (N_6278,N_5704,N_5705);
and U6279 (N_6279,N_5976,N_5823);
nor U6280 (N_6280,N_5798,N_5777);
or U6281 (N_6281,N_5935,N_5617);
nor U6282 (N_6282,N_5948,N_5903);
nor U6283 (N_6283,N_5828,N_5971);
or U6284 (N_6284,N_5740,N_5990);
nand U6285 (N_6285,N_5850,N_5956);
nor U6286 (N_6286,N_5654,N_5882);
or U6287 (N_6287,N_5898,N_5620);
nor U6288 (N_6288,N_5959,N_5843);
nand U6289 (N_6289,N_5986,N_5918);
or U6290 (N_6290,N_5740,N_5659);
nor U6291 (N_6291,N_5604,N_5706);
and U6292 (N_6292,N_5707,N_5628);
nor U6293 (N_6293,N_5656,N_5992);
xor U6294 (N_6294,N_5612,N_5840);
nor U6295 (N_6295,N_5629,N_5706);
or U6296 (N_6296,N_5818,N_5859);
nand U6297 (N_6297,N_5641,N_5908);
nand U6298 (N_6298,N_5980,N_5666);
or U6299 (N_6299,N_5703,N_5705);
and U6300 (N_6300,N_5850,N_5989);
xor U6301 (N_6301,N_5721,N_5899);
and U6302 (N_6302,N_5868,N_5871);
nand U6303 (N_6303,N_5688,N_5832);
nand U6304 (N_6304,N_5899,N_5857);
and U6305 (N_6305,N_5707,N_5627);
and U6306 (N_6306,N_5803,N_5962);
or U6307 (N_6307,N_5988,N_5761);
xor U6308 (N_6308,N_5622,N_5954);
or U6309 (N_6309,N_5914,N_5691);
or U6310 (N_6310,N_5765,N_5689);
and U6311 (N_6311,N_5755,N_5606);
nand U6312 (N_6312,N_5801,N_5805);
nand U6313 (N_6313,N_5912,N_5962);
nand U6314 (N_6314,N_5741,N_5701);
or U6315 (N_6315,N_5992,N_5880);
xor U6316 (N_6316,N_5712,N_5734);
xor U6317 (N_6317,N_5968,N_5771);
nand U6318 (N_6318,N_5957,N_5882);
and U6319 (N_6319,N_5655,N_5981);
nand U6320 (N_6320,N_5964,N_5939);
or U6321 (N_6321,N_5946,N_5749);
and U6322 (N_6322,N_5784,N_5938);
or U6323 (N_6323,N_5977,N_5713);
and U6324 (N_6324,N_5928,N_5973);
and U6325 (N_6325,N_5756,N_5952);
and U6326 (N_6326,N_5656,N_5847);
nor U6327 (N_6327,N_5831,N_5776);
nand U6328 (N_6328,N_5963,N_5637);
nor U6329 (N_6329,N_5959,N_5641);
nand U6330 (N_6330,N_5602,N_5900);
xor U6331 (N_6331,N_5601,N_5957);
nand U6332 (N_6332,N_5926,N_5987);
or U6333 (N_6333,N_5821,N_5990);
and U6334 (N_6334,N_5992,N_5816);
and U6335 (N_6335,N_5657,N_5868);
nor U6336 (N_6336,N_5707,N_5855);
or U6337 (N_6337,N_5602,N_5982);
xnor U6338 (N_6338,N_5743,N_5682);
and U6339 (N_6339,N_5988,N_5668);
and U6340 (N_6340,N_5713,N_5682);
or U6341 (N_6341,N_5928,N_5724);
nor U6342 (N_6342,N_5867,N_5862);
xor U6343 (N_6343,N_5834,N_5763);
or U6344 (N_6344,N_5880,N_5821);
nand U6345 (N_6345,N_5924,N_5780);
or U6346 (N_6346,N_5708,N_5769);
nor U6347 (N_6347,N_5956,N_5667);
nor U6348 (N_6348,N_5877,N_5652);
xnor U6349 (N_6349,N_5700,N_5777);
and U6350 (N_6350,N_5871,N_5748);
or U6351 (N_6351,N_5640,N_5884);
nor U6352 (N_6352,N_5892,N_5977);
xor U6353 (N_6353,N_5891,N_5649);
nor U6354 (N_6354,N_5820,N_5949);
nand U6355 (N_6355,N_5968,N_5644);
nor U6356 (N_6356,N_5907,N_5875);
xnor U6357 (N_6357,N_5876,N_5960);
or U6358 (N_6358,N_5703,N_5980);
nand U6359 (N_6359,N_5934,N_5866);
xnor U6360 (N_6360,N_5912,N_5713);
and U6361 (N_6361,N_5626,N_5662);
or U6362 (N_6362,N_5679,N_5990);
nor U6363 (N_6363,N_5892,N_5993);
or U6364 (N_6364,N_5647,N_5737);
nand U6365 (N_6365,N_5729,N_5669);
nand U6366 (N_6366,N_5717,N_5815);
or U6367 (N_6367,N_5903,N_5682);
xor U6368 (N_6368,N_5866,N_5637);
nand U6369 (N_6369,N_5857,N_5930);
or U6370 (N_6370,N_5903,N_5697);
nor U6371 (N_6371,N_5680,N_5779);
and U6372 (N_6372,N_5909,N_5664);
or U6373 (N_6373,N_5848,N_5864);
nand U6374 (N_6374,N_5704,N_5882);
nand U6375 (N_6375,N_5814,N_5651);
xor U6376 (N_6376,N_5639,N_5773);
or U6377 (N_6377,N_5795,N_5896);
and U6378 (N_6378,N_5691,N_5787);
xnor U6379 (N_6379,N_5804,N_5838);
nor U6380 (N_6380,N_5830,N_5660);
xnor U6381 (N_6381,N_5972,N_5838);
and U6382 (N_6382,N_5851,N_5987);
xor U6383 (N_6383,N_5607,N_5935);
xnor U6384 (N_6384,N_5741,N_5889);
and U6385 (N_6385,N_5768,N_5798);
and U6386 (N_6386,N_5851,N_5800);
or U6387 (N_6387,N_5775,N_5779);
nand U6388 (N_6388,N_5735,N_5779);
nor U6389 (N_6389,N_5998,N_5718);
or U6390 (N_6390,N_5785,N_5934);
nor U6391 (N_6391,N_5752,N_5833);
nor U6392 (N_6392,N_5836,N_5843);
xnor U6393 (N_6393,N_5616,N_5944);
nand U6394 (N_6394,N_5631,N_5681);
nor U6395 (N_6395,N_5931,N_5732);
or U6396 (N_6396,N_5709,N_5883);
or U6397 (N_6397,N_5952,N_5864);
nor U6398 (N_6398,N_5810,N_5715);
xor U6399 (N_6399,N_5675,N_5814);
or U6400 (N_6400,N_6394,N_6241);
xnor U6401 (N_6401,N_6151,N_6100);
xnor U6402 (N_6402,N_6179,N_6190);
or U6403 (N_6403,N_6320,N_6333);
and U6404 (N_6404,N_6214,N_6073);
xor U6405 (N_6405,N_6153,N_6075);
or U6406 (N_6406,N_6194,N_6276);
and U6407 (N_6407,N_6306,N_6165);
xor U6408 (N_6408,N_6095,N_6208);
xor U6409 (N_6409,N_6132,N_6036);
or U6410 (N_6410,N_6014,N_6027);
or U6411 (N_6411,N_6347,N_6029);
nor U6412 (N_6412,N_6023,N_6217);
nor U6413 (N_6413,N_6051,N_6229);
nor U6414 (N_6414,N_6334,N_6041);
nor U6415 (N_6415,N_6396,N_6129);
and U6416 (N_6416,N_6032,N_6285);
xnor U6417 (N_6417,N_6008,N_6260);
nand U6418 (N_6418,N_6055,N_6018);
xor U6419 (N_6419,N_6300,N_6031);
xor U6420 (N_6420,N_6067,N_6056);
xnor U6421 (N_6421,N_6133,N_6355);
or U6422 (N_6422,N_6150,N_6262);
nor U6423 (N_6423,N_6188,N_6220);
xor U6424 (N_6424,N_6038,N_6119);
or U6425 (N_6425,N_6127,N_6037);
nand U6426 (N_6426,N_6392,N_6203);
nor U6427 (N_6427,N_6328,N_6135);
or U6428 (N_6428,N_6216,N_6022);
nand U6429 (N_6429,N_6069,N_6357);
nand U6430 (N_6430,N_6389,N_6168);
or U6431 (N_6431,N_6265,N_6263);
or U6432 (N_6432,N_6379,N_6255);
nand U6433 (N_6433,N_6227,N_6221);
or U6434 (N_6434,N_6293,N_6068);
xnor U6435 (N_6435,N_6324,N_6259);
and U6436 (N_6436,N_6232,N_6278);
nor U6437 (N_6437,N_6313,N_6269);
xor U6438 (N_6438,N_6024,N_6351);
nand U6439 (N_6439,N_6287,N_6273);
nand U6440 (N_6440,N_6286,N_6366);
nand U6441 (N_6441,N_6201,N_6044);
xor U6442 (N_6442,N_6280,N_6172);
xnor U6443 (N_6443,N_6114,N_6159);
xor U6444 (N_6444,N_6195,N_6021);
xor U6445 (N_6445,N_6146,N_6378);
xnor U6446 (N_6446,N_6141,N_6242);
xnor U6447 (N_6447,N_6131,N_6149);
or U6448 (N_6448,N_6384,N_6171);
nor U6449 (N_6449,N_6012,N_6152);
and U6450 (N_6450,N_6167,N_6289);
nor U6451 (N_6451,N_6381,N_6015);
nand U6452 (N_6452,N_6202,N_6019);
xnor U6453 (N_6453,N_6175,N_6110);
xnor U6454 (N_6454,N_6092,N_6145);
xnor U6455 (N_6455,N_6047,N_6206);
or U6456 (N_6456,N_6016,N_6377);
nand U6457 (N_6457,N_6388,N_6139);
or U6458 (N_6458,N_6246,N_6084);
or U6459 (N_6459,N_6080,N_6117);
or U6460 (N_6460,N_6143,N_6148);
xnor U6461 (N_6461,N_6089,N_6130);
nor U6462 (N_6462,N_6372,N_6296);
nand U6463 (N_6463,N_6233,N_6050);
and U6464 (N_6464,N_6118,N_6025);
nand U6465 (N_6465,N_6197,N_6310);
nor U6466 (N_6466,N_6222,N_6213);
and U6467 (N_6467,N_6006,N_6077);
nand U6468 (N_6468,N_6272,N_6251);
nor U6469 (N_6469,N_6048,N_6199);
and U6470 (N_6470,N_6316,N_6070);
and U6471 (N_6471,N_6196,N_6001);
and U6472 (N_6472,N_6277,N_6111);
xor U6473 (N_6473,N_6356,N_6256);
xnor U6474 (N_6474,N_6099,N_6354);
nand U6475 (N_6475,N_6370,N_6049);
and U6476 (N_6476,N_6395,N_6339);
and U6477 (N_6477,N_6093,N_6258);
nand U6478 (N_6478,N_6128,N_6076);
nor U6479 (N_6479,N_6043,N_6304);
xor U6480 (N_6480,N_6173,N_6218);
or U6481 (N_6481,N_6108,N_6361);
and U6482 (N_6482,N_6398,N_6071);
nand U6483 (N_6483,N_6298,N_6096);
nor U6484 (N_6484,N_6061,N_6267);
and U6485 (N_6485,N_6236,N_6030);
xor U6486 (N_6486,N_6302,N_6033);
and U6487 (N_6487,N_6137,N_6109);
nor U6488 (N_6488,N_6375,N_6340);
or U6489 (N_6489,N_6112,N_6097);
xnor U6490 (N_6490,N_6091,N_6281);
nand U6491 (N_6491,N_6087,N_6059);
nand U6492 (N_6492,N_6138,N_6326);
and U6493 (N_6493,N_6226,N_6397);
and U6494 (N_6494,N_6297,N_6261);
or U6495 (N_6495,N_6387,N_6166);
nor U6496 (N_6496,N_6086,N_6363);
and U6497 (N_6497,N_6185,N_6243);
nor U6498 (N_6498,N_6360,N_6386);
and U6499 (N_6499,N_6140,N_6292);
xnor U6500 (N_6500,N_6072,N_6101);
nand U6501 (N_6501,N_6184,N_6104);
nor U6502 (N_6502,N_6391,N_6342);
or U6503 (N_6503,N_6182,N_6090);
xor U6504 (N_6504,N_6329,N_6115);
and U6505 (N_6505,N_6039,N_6215);
xor U6506 (N_6506,N_6063,N_6368);
nor U6507 (N_6507,N_6349,N_6317);
and U6508 (N_6508,N_6335,N_6125);
nor U6509 (N_6509,N_6078,N_6332);
nand U6510 (N_6510,N_6373,N_6126);
and U6511 (N_6511,N_6338,N_6007);
or U6512 (N_6512,N_6345,N_6209);
xor U6513 (N_6513,N_6299,N_6295);
nor U6514 (N_6514,N_6249,N_6374);
nand U6515 (N_6515,N_6106,N_6352);
and U6516 (N_6516,N_6311,N_6219);
nor U6517 (N_6517,N_6189,N_6094);
nand U6518 (N_6518,N_6283,N_6026);
xnor U6519 (N_6519,N_6383,N_6376);
xnor U6520 (N_6520,N_6010,N_6186);
xnor U6521 (N_6521,N_6393,N_6231);
nand U6522 (N_6522,N_6122,N_6123);
and U6523 (N_6523,N_6204,N_6239);
nand U6524 (N_6524,N_6382,N_6230);
xor U6525 (N_6525,N_6211,N_6271);
xor U6526 (N_6526,N_6004,N_6181);
or U6527 (N_6527,N_6319,N_6013);
or U6528 (N_6528,N_6344,N_6074);
and U6529 (N_6529,N_6113,N_6142);
nor U6530 (N_6530,N_6079,N_6088);
and U6531 (N_6531,N_6169,N_6158);
nand U6532 (N_6532,N_6144,N_6358);
nand U6533 (N_6533,N_6341,N_6365);
nand U6534 (N_6534,N_6224,N_6052);
and U6535 (N_6535,N_6157,N_6098);
or U6536 (N_6536,N_6028,N_6294);
and U6537 (N_6537,N_6264,N_6060);
and U6538 (N_6538,N_6385,N_6275);
nand U6539 (N_6539,N_6081,N_6228);
xnor U6540 (N_6540,N_6318,N_6066);
nand U6541 (N_6541,N_6134,N_6200);
and U6542 (N_6542,N_6178,N_6322);
nand U6543 (N_6543,N_6331,N_6058);
and U6544 (N_6544,N_6234,N_6210);
or U6545 (N_6545,N_6042,N_6225);
and U6546 (N_6546,N_6174,N_6223);
nor U6547 (N_6547,N_6017,N_6160);
nand U6548 (N_6548,N_6301,N_6336);
xor U6549 (N_6549,N_6003,N_6235);
nor U6550 (N_6550,N_6082,N_6253);
xor U6551 (N_6551,N_6162,N_6274);
and U6552 (N_6552,N_6353,N_6367);
or U6553 (N_6553,N_6191,N_6252);
and U6554 (N_6554,N_6268,N_6245);
and U6555 (N_6555,N_6282,N_6116);
and U6556 (N_6556,N_6020,N_6207);
nor U6557 (N_6557,N_6315,N_6161);
xnor U6558 (N_6558,N_6187,N_6350);
xor U6559 (N_6559,N_6240,N_6290);
nor U6560 (N_6560,N_6284,N_6000);
xor U6561 (N_6561,N_6279,N_6257);
or U6562 (N_6562,N_6247,N_6053);
and U6563 (N_6563,N_6399,N_6064);
nor U6564 (N_6564,N_6359,N_6046);
xor U6565 (N_6565,N_6205,N_6321);
and U6566 (N_6566,N_6040,N_6248);
xor U6567 (N_6567,N_6192,N_6380);
or U6568 (N_6568,N_6054,N_6183);
nor U6569 (N_6569,N_6198,N_6156);
and U6570 (N_6570,N_6120,N_6034);
xnor U6571 (N_6571,N_6103,N_6348);
or U6572 (N_6572,N_6362,N_6154);
or U6573 (N_6573,N_6121,N_6346);
xor U6574 (N_6574,N_6193,N_6107);
nand U6575 (N_6575,N_6266,N_6057);
nand U6576 (N_6576,N_6005,N_6180);
xor U6577 (N_6577,N_6305,N_6102);
or U6578 (N_6578,N_6212,N_6237);
or U6579 (N_6579,N_6011,N_6170);
and U6580 (N_6580,N_6083,N_6250);
nand U6581 (N_6581,N_6062,N_6288);
xnor U6582 (N_6582,N_6065,N_6105);
and U6583 (N_6583,N_6308,N_6136);
nand U6584 (N_6584,N_6270,N_6303);
nand U6585 (N_6585,N_6312,N_6009);
and U6586 (N_6586,N_6238,N_6163);
or U6587 (N_6587,N_6369,N_6343);
and U6588 (N_6588,N_6327,N_6291);
xor U6589 (N_6589,N_6155,N_6045);
and U6590 (N_6590,N_6147,N_6124);
xnor U6591 (N_6591,N_6330,N_6254);
and U6592 (N_6592,N_6371,N_6176);
nand U6593 (N_6593,N_6390,N_6325);
nand U6594 (N_6594,N_6307,N_6309);
nor U6595 (N_6595,N_6177,N_6164);
or U6596 (N_6596,N_6314,N_6323);
nor U6597 (N_6597,N_6364,N_6002);
or U6598 (N_6598,N_6035,N_6085);
xor U6599 (N_6599,N_6337,N_6244);
xnor U6600 (N_6600,N_6002,N_6229);
nor U6601 (N_6601,N_6001,N_6079);
or U6602 (N_6602,N_6019,N_6237);
or U6603 (N_6603,N_6264,N_6053);
nor U6604 (N_6604,N_6224,N_6146);
nand U6605 (N_6605,N_6217,N_6304);
or U6606 (N_6606,N_6247,N_6277);
nand U6607 (N_6607,N_6284,N_6097);
nand U6608 (N_6608,N_6125,N_6080);
nand U6609 (N_6609,N_6012,N_6092);
xor U6610 (N_6610,N_6366,N_6120);
nor U6611 (N_6611,N_6152,N_6021);
nor U6612 (N_6612,N_6075,N_6295);
nand U6613 (N_6613,N_6151,N_6309);
or U6614 (N_6614,N_6357,N_6273);
or U6615 (N_6615,N_6205,N_6070);
nor U6616 (N_6616,N_6087,N_6246);
nor U6617 (N_6617,N_6317,N_6219);
nor U6618 (N_6618,N_6333,N_6171);
nand U6619 (N_6619,N_6063,N_6220);
or U6620 (N_6620,N_6104,N_6330);
xor U6621 (N_6621,N_6324,N_6336);
xor U6622 (N_6622,N_6358,N_6128);
nor U6623 (N_6623,N_6323,N_6158);
or U6624 (N_6624,N_6286,N_6363);
nor U6625 (N_6625,N_6250,N_6349);
xnor U6626 (N_6626,N_6162,N_6007);
nor U6627 (N_6627,N_6010,N_6264);
or U6628 (N_6628,N_6257,N_6324);
xnor U6629 (N_6629,N_6210,N_6107);
or U6630 (N_6630,N_6326,N_6230);
nand U6631 (N_6631,N_6123,N_6063);
or U6632 (N_6632,N_6354,N_6215);
and U6633 (N_6633,N_6051,N_6334);
and U6634 (N_6634,N_6141,N_6052);
and U6635 (N_6635,N_6036,N_6151);
nor U6636 (N_6636,N_6040,N_6184);
xnor U6637 (N_6637,N_6256,N_6281);
and U6638 (N_6638,N_6377,N_6077);
nor U6639 (N_6639,N_6398,N_6022);
nor U6640 (N_6640,N_6237,N_6221);
or U6641 (N_6641,N_6087,N_6222);
xnor U6642 (N_6642,N_6275,N_6258);
nor U6643 (N_6643,N_6317,N_6008);
nand U6644 (N_6644,N_6199,N_6358);
or U6645 (N_6645,N_6278,N_6341);
and U6646 (N_6646,N_6210,N_6176);
nand U6647 (N_6647,N_6397,N_6389);
nor U6648 (N_6648,N_6042,N_6052);
nor U6649 (N_6649,N_6089,N_6287);
nand U6650 (N_6650,N_6273,N_6345);
xnor U6651 (N_6651,N_6017,N_6234);
and U6652 (N_6652,N_6165,N_6348);
and U6653 (N_6653,N_6042,N_6357);
nor U6654 (N_6654,N_6039,N_6160);
nor U6655 (N_6655,N_6102,N_6230);
nor U6656 (N_6656,N_6227,N_6344);
and U6657 (N_6657,N_6115,N_6137);
nor U6658 (N_6658,N_6107,N_6062);
and U6659 (N_6659,N_6059,N_6053);
nor U6660 (N_6660,N_6004,N_6232);
and U6661 (N_6661,N_6123,N_6209);
and U6662 (N_6662,N_6371,N_6075);
or U6663 (N_6663,N_6026,N_6028);
or U6664 (N_6664,N_6272,N_6181);
nor U6665 (N_6665,N_6188,N_6095);
and U6666 (N_6666,N_6337,N_6307);
and U6667 (N_6667,N_6163,N_6237);
xor U6668 (N_6668,N_6270,N_6188);
xor U6669 (N_6669,N_6012,N_6023);
xnor U6670 (N_6670,N_6168,N_6270);
xnor U6671 (N_6671,N_6227,N_6361);
or U6672 (N_6672,N_6183,N_6219);
and U6673 (N_6673,N_6025,N_6310);
nand U6674 (N_6674,N_6117,N_6366);
xnor U6675 (N_6675,N_6153,N_6304);
nand U6676 (N_6676,N_6290,N_6352);
nor U6677 (N_6677,N_6040,N_6189);
nor U6678 (N_6678,N_6241,N_6276);
xor U6679 (N_6679,N_6011,N_6377);
nor U6680 (N_6680,N_6194,N_6046);
xnor U6681 (N_6681,N_6019,N_6337);
and U6682 (N_6682,N_6127,N_6154);
nand U6683 (N_6683,N_6288,N_6341);
and U6684 (N_6684,N_6369,N_6334);
nor U6685 (N_6685,N_6133,N_6089);
nor U6686 (N_6686,N_6119,N_6026);
xor U6687 (N_6687,N_6174,N_6127);
or U6688 (N_6688,N_6347,N_6238);
nor U6689 (N_6689,N_6238,N_6373);
nand U6690 (N_6690,N_6233,N_6044);
or U6691 (N_6691,N_6054,N_6023);
nor U6692 (N_6692,N_6353,N_6294);
and U6693 (N_6693,N_6268,N_6359);
nor U6694 (N_6694,N_6342,N_6386);
nor U6695 (N_6695,N_6012,N_6080);
and U6696 (N_6696,N_6310,N_6295);
xor U6697 (N_6697,N_6207,N_6313);
and U6698 (N_6698,N_6114,N_6161);
nor U6699 (N_6699,N_6061,N_6228);
and U6700 (N_6700,N_6143,N_6214);
xnor U6701 (N_6701,N_6090,N_6335);
and U6702 (N_6702,N_6131,N_6309);
nand U6703 (N_6703,N_6304,N_6236);
nand U6704 (N_6704,N_6365,N_6391);
nand U6705 (N_6705,N_6175,N_6012);
or U6706 (N_6706,N_6270,N_6335);
or U6707 (N_6707,N_6292,N_6313);
xnor U6708 (N_6708,N_6238,N_6222);
xor U6709 (N_6709,N_6315,N_6253);
and U6710 (N_6710,N_6062,N_6105);
nand U6711 (N_6711,N_6255,N_6178);
nand U6712 (N_6712,N_6271,N_6335);
xor U6713 (N_6713,N_6076,N_6329);
and U6714 (N_6714,N_6149,N_6138);
nor U6715 (N_6715,N_6199,N_6058);
xnor U6716 (N_6716,N_6391,N_6055);
xnor U6717 (N_6717,N_6205,N_6341);
xnor U6718 (N_6718,N_6071,N_6043);
xor U6719 (N_6719,N_6110,N_6370);
nor U6720 (N_6720,N_6006,N_6075);
nor U6721 (N_6721,N_6144,N_6222);
nand U6722 (N_6722,N_6252,N_6303);
nand U6723 (N_6723,N_6061,N_6093);
nand U6724 (N_6724,N_6248,N_6134);
and U6725 (N_6725,N_6029,N_6291);
and U6726 (N_6726,N_6314,N_6236);
xnor U6727 (N_6727,N_6093,N_6070);
nand U6728 (N_6728,N_6265,N_6325);
nand U6729 (N_6729,N_6134,N_6046);
nand U6730 (N_6730,N_6193,N_6067);
and U6731 (N_6731,N_6166,N_6074);
xnor U6732 (N_6732,N_6092,N_6132);
nand U6733 (N_6733,N_6319,N_6109);
nand U6734 (N_6734,N_6188,N_6298);
and U6735 (N_6735,N_6076,N_6134);
and U6736 (N_6736,N_6008,N_6177);
or U6737 (N_6737,N_6343,N_6052);
or U6738 (N_6738,N_6317,N_6057);
nor U6739 (N_6739,N_6038,N_6118);
nor U6740 (N_6740,N_6063,N_6184);
and U6741 (N_6741,N_6391,N_6258);
nor U6742 (N_6742,N_6019,N_6384);
nand U6743 (N_6743,N_6265,N_6270);
or U6744 (N_6744,N_6112,N_6091);
xor U6745 (N_6745,N_6310,N_6265);
nand U6746 (N_6746,N_6183,N_6151);
nor U6747 (N_6747,N_6173,N_6187);
xor U6748 (N_6748,N_6069,N_6370);
xor U6749 (N_6749,N_6120,N_6232);
or U6750 (N_6750,N_6261,N_6117);
nand U6751 (N_6751,N_6377,N_6327);
xor U6752 (N_6752,N_6238,N_6096);
xnor U6753 (N_6753,N_6244,N_6391);
nor U6754 (N_6754,N_6141,N_6306);
or U6755 (N_6755,N_6086,N_6191);
nor U6756 (N_6756,N_6130,N_6292);
and U6757 (N_6757,N_6392,N_6045);
and U6758 (N_6758,N_6356,N_6224);
nor U6759 (N_6759,N_6114,N_6009);
or U6760 (N_6760,N_6076,N_6370);
and U6761 (N_6761,N_6391,N_6291);
xnor U6762 (N_6762,N_6138,N_6105);
or U6763 (N_6763,N_6162,N_6066);
nor U6764 (N_6764,N_6264,N_6331);
xor U6765 (N_6765,N_6004,N_6352);
nand U6766 (N_6766,N_6284,N_6241);
nor U6767 (N_6767,N_6277,N_6109);
nor U6768 (N_6768,N_6005,N_6164);
xor U6769 (N_6769,N_6241,N_6188);
and U6770 (N_6770,N_6322,N_6084);
and U6771 (N_6771,N_6324,N_6208);
or U6772 (N_6772,N_6077,N_6202);
nor U6773 (N_6773,N_6392,N_6055);
and U6774 (N_6774,N_6328,N_6031);
nor U6775 (N_6775,N_6302,N_6225);
or U6776 (N_6776,N_6387,N_6249);
nor U6777 (N_6777,N_6281,N_6263);
and U6778 (N_6778,N_6396,N_6037);
or U6779 (N_6779,N_6054,N_6185);
nand U6780 (N_6780,N_6366,N_6367);
or U6781 (N_6781,N_6089,N_6361);
nand U6782 (N_6782,N_6163,N_6219);
nor U6783 (N_6783,N_6060,N_6037);
nor U6784 (N_6784,N_6365,N_6113);
or U6785 (N_6785,N_6046,N_6345);
and U6786 (N_6786,N_6134,N_6102);
and U6787 (N_6787,N_6049,N_6162);
and U6788 (N_6788,N_6144,N_6171);
xnor U6789 (N_6789,N_6210,N_6396);
nor U6790 (N_6790,N_6062,N_6143);
nand U6791 (N_6791,N_6117,N_6266);
xor U6792 (N_6792,N_6180,N_6133);
xnor U6793 (N_6793,N_6082,N_6186);
nand U6794 (N_6794,N_6371,N_6262);
xnor U6795 (N_6795,N_6216,N_6372);
xor U6796 (N_6796,N_6234,N_6164);
xor U6797 (N_6797,N_6146,N_6123);
or U6798 (N_6798,N_6379,N_6362);
nor U6799 (N_6799,N_6355,N_6206);
nor U6800 (N_6800,N_6594,N_6571);
and U6801 (N_6801,N_6583,N_6563);
and U6802 (N_6802,N_6514,N_6742);
or U6803 (N_6803,N_6499,N_6758);
or U6804 (N_6804,N_6430,N_6556);
nor U6805 (N_6805,N_6605,N_6738);
nand U6806 (N_6806,N_6592,N_6727);
nand U6807 (N_6807,N_6585,N_6717);
nor U6808 (N_6808,N_6636,N_6584);
and U6809 (N_6809,N_6622,N_6716);
or U6810 (N_6810,N_6435,N_6692);
or U6811 (N_6811,N_6537,N_6502);
nand U6812 (N_6812,N_6478,N_6641);
nand U6813 (N_6813,N_6560,N_6721);
and U6814 (N_6814,N_6649,N_6658);
nor U6815 (N_6815,N_6558,N_6755);
and U6816 (N_6816,N_6796,N_6667);
and U6817 (N_6817,N_6718,N_6714);
xnor U6818 (N_6818,N_6523,N_6766);
and U6819 (N_6819,N_6790,N_6688);
and U6820 (N_6820,N_6544,N_6413);
and U6821 (N_6821,N_6724,N_6771);
nand U6822 (N_6822,N_6473,N_6606);
nand U6823 (N_6823,N_6572,N_6446);
nor U6824 (N_6824,N_6479,N_6640);
nor U6825 (N_6825,N_6775,N_6533);
nand U6826 (N_6826,N_6565,N_6626);
xor U6827 (N_6827,N_6722,N_6557);
nor U6828 (N_6828,N_6400,N_6728);
nand U6829 (N_6829,N_6483,N_6554);
or U6830 (N_6830,N_6778,N_6534);
xnor U6831 (N_6831,N_6675,N_6782);
nor U6832 (N_6832,N_6451,N_6509);
and U6833 (N_6833,N_6507,N_6603);
xor U6834 (N_6834,N_6673,N_6672);
xnor U6835 (N_6835,N_6547,N_6769);
nand U6836 (N_6836,N_6639,N_6518);
nand U6837 (N_6837,N_6500,N_6632);
and U6838 (N_6838,N_6657,N_6700);
or U6839 (N_6839,N_6598,N_6419);
nand U6840 (N_6840,N_6732,N_6741);
nor U6841 (N_6841,N_6408,N_6531);
xor U6842 (N_6842,N_6498,N_6420);
or U6843 (N_6843,N_6783,N_6638);
nor U6844 (N_6844,N_6651,N_6734);
or U6845 (N_6845,N_6645,N_6450);
nor U6846 (N_6846,N_6614,N_6600);
or U6847 (N_6847,N_6505,N_6597);
or U6848 (N_6848,N_6511,N_6476);
nor U6849 (N_6849,N_6752,N_6454);
or U6850 (N_6850,N_6604,N_6480);
nor U6851 (N_6851,N_6616,N_6449);
nor U6852 (N_6852,N_6481,N_6617);
nor U6853 (N_6853,N_6684,N_6411);
xor U6854 (N_6854,N_6553,N_6494);
and U6855 (N_6855,N_6461,N_6540);
and U6856 (N_6856,N_6417,N_6767);
nand U6857 (N_6857,N_6660,N_6777);
nor U6858 (N_6858,N_6631,N_6624);
or U6859 (N_6859,N_6542,N_6409);
xnor U6860 (N_6860,N_6635,N_6410);
xor U6861 (N_6861,N_6762,N_6780);
or U6862 (N_6862,N_6686,N_6510);
and U6863 (N_6863,N_6418,N_6564);
or U6864 (N_6864,N_6754,N_6576);
nand U6865 (N_6865,N_6559,N_6730);
nor U6866 (N_6866,N_6665,N_6466);
and U6867 (N_6867,N_6587,N_6527);
or U6868 (N_6868,N_6415,N_6432);
and U6869 (N_6869,N_6590,N_6562);
nor U6870 (N_6870,N_6412,N_6611);
xor U6871 (N_6871,N_6702,N_6647);
nor U6872 (N_6872,N_6669,N_6713);
nor U6873 (N_6873,N_6630,N_6524);
and U6874 (N_6874,N_6776,N_6452);
nor U6875 (N_6875,N_6488,N_6586);
or U6876 (N_6876,N_6792,N_6575);
and U6877 (N_6877,N_6462,N_6751);
xnor U6878 (N_6878,N_6487,N_6519);
and U6879 (N_6879,N_6723,N_6791);
and U6880 (N_6880,N_6512,N_6472);
and U6881 (N_6881,N_6474,N_6753);
nor U6882 (N_6882,N_6469,N_6619);
nand U6883 (N_6883,N_6555,N_6642);
nor U6884 (N_6884,N_6529,N_6689);
nor U6885 (N_6885,N_6793,N_6679);
and U6886 (N_6886,N_6425,N_6629);
nor U6887 (N_6887,N_6666,N_6460);
or U6888 (N_6888,N_6489,N_6661);
or U6889 (N_6889,N_6463,N_6426);
or U6890 (N_6890,N_6467,N_6433);
xnor U6891 (N_6891,N_6668,N_6595);
xor U6892 (N_6892,N_6715,N_6704);
nor U6893 (N_6893,N_6455,N_6427);
nor U6894 (N_6894,N_6726,N_6516);
xor U6895 (N_6895,N_6404,N_6736);
xor U6896 (N_6896,N_6610,N_6422);
nand U6897 (N_6897,N_6545,N_6677);
nand U6898 (N_6898,N_6464,N_6477);
xnor U6899 (N_6899,N_6773,N_6761);
nand U6900 (N_6900,N_6593,N_6765);
and U6901 (N_6901,N_6705,N_6437);
xnor U6902 (N_6902,N_6628,N_6764);
nand U6903 (N_6903,N_6681,N_6744);
nand U6904 (N_6904,N_6613,N_6567);
or U6905 (N_6905,N_6486,N_6401);
or U6906 (N_6906,N_6618,N_6698);
nor U6907 (N_6907,N_6579,N_6407);
xnor U6908 (N_6908,N_6709,N_6470);
nor U6909 (N_6909,N_6503,N_6615);
nor U6910 (N_6910,N_6710,N_6599);
nand U6911 (N_6911,N_6442,N_6772);
and U6912 (N_6912,N_6458,N_6694);
and U6913 (N_6913,N_6546,N_6440);
nand U6914 (N_6914,N_6438,N_6530);
and U6915 (N_6915,N_6747,N_6428);
or U6916 (N_6916,N_6431,N_6471);
nor U6917 (N_6917,N_6561,N_6746);
nor U6918 (N_6918,N_6457,N_6490);
xor U6919 (N_6919,N_6646,N_6441);
nand U6920 (N_6920,N_6712,N_6749);
or U6921 (N_6921,N_6569,N_6685);
and U6922 (N_6922,N_6608,N_6508);
nand U6923 (N_6923,N_6696,N_6623);
or U6924 (N_6924,N_6528,N_6740);
and U6925 (N_6925,N_6570,N_6515);
nand U6926 (N_6926,N_6612,N_6731);
nand U6927 (N_6927,N_6743,N_6525);
or U6928 (N_6928,N_6539,N_6785);
and U6929 (N_6929,N_6797,N_6699);
nand U6930 (N_6930,N_6653,N_6779);
and U6931 (N_6931,N_6548,N_6453);
xor U6932 (N_6932,N_6707,N_6670);
nor U6933 (N_6933,N_6621,N_6549);
and U6934 (N_6934,N_6609,N_6627);
and U6935 (N_6935,N_6482,N_6448);
nor U6936 (N_6936,N_6532,N_6729);
nand U6937 (N_6937,N_6795,N_6521);
and U6938 (N_6938,N_6706,N_6475);
nand U6939 (N_6939,N_6701,N_6620);
or U6940 (N_6940,N_6650,N_6648);
xnor U6941 (N_6941,N_6687,N_6535);
nand U6942 (N_6942,N_6787,N_6637);
and U6943 (N_6943,N_6403,N_6484);
nand U6944 (N_6944,N_6725,N_6703);
xnor U6945 (N_6945,N_6578,N_6662);
xor U6946 (N_6946,N_6443,N_6436);
and U6947 (N_6947,N_6682,N_6550);
xor U6948 (N_6948,N_6759,N_6424);
xor U6949 (N_6949,N_6497,N_6633);
nor U6950 (N_6950,N_6551,N_6693);
nand U6951 (N_6951,N_6581,N_6748);
xnor U6952 (N_6952,N_6774,N_6421);
nor U6953 (N_6953,N_6799,N_6652);
and U6954 (N_6954,N_6735,N_6444);
nand U6955 (N_6955,N_6406,N_6784);
or U6956 (N_6956,N_6697,N_6739);
nand U6957 (N_6957,N_6520,N_6459);
nand U6958 (N_6958,N_6589,N_6745);
and U6959 (N_6959,N_6504,N_6405);
or U6960 (N_6960,N_6678,N_6492);
or U6961 (N_6961,N_6763,N_6485);
nand U6962 (N_6962,N_6607,N_6695);
nor U6963 (N_6963,N_6552,N_6543);
nor U6964 (N_6964,N_6574,N_6445);
nand U6965 (N_6965,N_6691,N_6634);
xnor U6966 (N_6966,N_6596,N_6416);
and U6967 (N_6967,N_6654,N_6496);
nor U6968 (N_6968,N_6536,N_6733);
and U6969 (N_6969,N_6671,N_6756);
nor U6970 (N_6970,N_6768,N_6788);
nor U6971 (N_6971,N_6708,N_6541);
nor U6972 (N_6972,N_6465,N_6798);
nor U6973 (N_6973,N_6402,N_6750);
nor U6974 (N_6974,N_6760,N_6781);
or U6975 (N_6975,N_6495,N_6737);
or U6976 (N_6976,N_6644,N_6588);
xor U6977 (N_6977,N_6429,N_6577);
nand U6978 (N_6978,N_6456,N_6789);
nand U6979 (N_6979,N_6526,N_6517);
nor U6980 (N_6980,N_6680,N_6423);
nor U6981 (N_6981,N_6757,N_6711);
nor U6982 (N_6982,N_6468,N_6656);
xnor U6983 (N_6983,N_6601,N_6794);
and U6984 (N_6984,N_6655,N_6538);
or U6985 (N_6985,N_6591,N_6719);
xnor U6986 (N_6986,N_6522,N_6683);
nor U6987 (N_6987,N_6663,N_6720);
and U6988 (N_6988,N_6506,N_6568);
xor U6989 (N_6989,N_6513,N_6674);
and U6990 (N_6990,N_6493,N_6580);
xor U6991 (N_6991,N_6434,N_6566);
nor U6992 (N_6992,N_6770,N_6786);
xnor U6993 (N_6993,N_6625,N_6602);
or U6994 (N_6994,N_6501,N_6690);
and U6995 (N_6995,N_6582,N_6447);
and U6996 (N_6996,N_6491,N_6643);
or U6997 (N_6997,N_6414,N_6659);
nor U6998 (N_6998,N_6573,N_6664);
xnor U6999 (N_6999,N_6439,N_6676);
or U7000 (N_7000,N_6772,N_6664);
nand U7001 (N_7001,N_6796,N_6696);
nor U7002 (N_7002,N_6706,N_6700);
nor U7003 (N_7003,N_6533,N_6476);
xnor U7004 (N_7004,N_6683,N_6714);
xnor U7005 (N_7005,N_6406,N_6553);
nor U7006 (N_7006,N_6682,N_6709);
nor U7007 (N_7007,N_6777,N_6554);
nand U7008 (N_7008,N_6404,N_6619);
or U7009 (N_7009,N_6573,N_6497);
or U7010 (N_7010,N_6754,N_6742);
xnor U7011 (N_7011,N_6639,N_6561);
nor U7012 (N_7012,N_6447,N_6792);
and U7013 (N_7013,N_6705,N_6404);
and U7014 (N_7014,N_6562,N_6597);
and U7015 (N_7015,N_6537,N_6672);
or U7016 (N_7016,N_6644,N_6715);
and U7017 (N_7017,N_6405,N_6495);
nand U7018 (N_7018,N_6537,N_6416);
and U7019 (N_7019,N_6639,N_6736);
nand U7020 (N_7020,N_6618,N_6473);
and U7021 (N_7021,N_6497,N_6671);
nor U7022 (N_7022,N_6689,N_6701);
or U7023 (N_7023,N_6639,N_6595);
or U7024 (N_7024,N_6624,N_6718);
nand U7025 (N_7025,N_6659,N_6491);
nand U7026 (N_7026,N_6458,N_6528);
nand U7027 (N_7027,N_6643,N_6589);
xor U7028 (N_7028,N_6768,N_6441);
and U7029 (N_7029,N_6695,N_6788);
or U7030 (N_7030,N_6792,N_6669);
and U7031 (N_7031,N_6512,N_6651);
xnor U7032 (N_7032,N_6487,N_6773);
nand U7033 (N_7033,N_6584,N_6787);
and U7034 (N_7034,N_6679,N_6738);
xor U7035 (N_7035,N_6650,N_6451);
nand U7036 (N_7036,N_6562,N_6641);
nor U7037 (N_7037,N_6450,N_6552);
xor U7038 (N_7038,N_6763,N_6790);
xnor U7039 (N_7039,N_6656,N_6541);
nand U7040 (N_7040,N_6446,N_6540);
nand U7041 (N_7041,N_6713,N_6769);
xnor U7042 (N_7042,N_6477,N_6522);
xor U7043 (N_7043,N_6729,N_6423);
xor U7044 (N_7044,N_6724,N_6567);
xnor U7045 (N_7045,N_6524,N_6747);
and U7046 (N_7046,N_6406,N_6699);
and U7047 (N_7047,N_6616,N_6462);
nand U7048 (N_7048,N_6694,N_6534);
and U7049 (N_7049,N_6693,N_6604);
and U7050 (N_7050,N_6437,N_6696);
or U7051 (N_7051,N_6727,N_6432);
nand U7052 (N_7052,N_6720,N_6474);
or U7053 (N_7053,N_6425,N_6743);
xnor U7054 (N_7054,N_6489,N_6637);
xnor U7055 (N_7055,N_6659,N_6613);
nand U7056 (N_7056,N_6453,N_6443);
xnor U7057 (N_7057,N_6466,N_6558);
xnor U7058 (N_7058,N_6667,N_6471);
xnor U7059 (N_7059,N_6743,N_6459);
nand U7060 (N_7060,N_6585,N_6483);
nand U7061 (N_7061,N_6524,N_6558);
nand U7062 (N_7062,N_6444,N_6508);
and U7063 (N_7063,N_6725,N_6673);
nand U7064 (N_7064,N_6401,N_6751);
nand U7065 (N_7065,N_6756,N_6419);
nor U7066 (N_7066,N_6779,N_6758);
or U7067 (N_7067,N_6554,N_6427);
or U7068 (N_7068,N_6444,N_6697);
and U7069 (N_7069,N_6697,N_6575);
or U7070 (N_7070,N_6737,N_6594);
nand U7071 (N_7071,N_6638,N_6730);
xor U7072 (N_7072,N_6670,N_6480);
or U7073 (N_7073,N_6436,N_6528);
xnor U7074 (N_7074,N_6705,N_6599);
xnor U7075 (N_7075,N_6430,N_6498);
nor U7076 (N_7076,N_6504,N_6732);
xnor U7077 (N_7077,N_6442,N_6411);
xor U7078 (N_7078,N_6505,N_6516);
or U7079 (N_7079,N_6637,N_6669);
and U7080 (N_7080,N_6597,N_6714);
xor U7081 (N_7081,N_6727,N_6643);
nor U7082 (N_7082,N_6500,N_6624);
nand U7083 (N_7083,N_6526,N_6444);
nor U7084 (N_7084,N_6494,N_6466);
xnor U7085 (N_7085,N_6555,N_6612);
xnor U7086 (N_7086,N_6495,N_6492);
and U7087 (N_7087,N_6466,N_6526);
or U7088 (N_7088,N_6464,N_6572);
or U7089 (N_7089,N_6471,N_6611);
or U7090 (N_7090,N_6780,N_6525);
nor U7091 (N_7091,N_6689,N_6421);
nand U7092 (N_7092,N_6545,N_6616);
and U7093 (N_7093,N_6429,N_6788);
nand U7094 (N_7094,N_6401,N_6527);
or U7095 (N_7095,N_6612,N_6738);
nand U7096 (N_7096,N_6442,N_6446);
or U7097 (N_7097,N_6737,N_6759);
and U7098 (N_7098,N_6604,N_6484);
and U7099 (N_7099,N_6749,N_6421);
or U7100 (N_7100,N_6407,N_6469);
nand U7101 (N_7101,N_6663,N_6547);
nand U7102 (N_7102,N_6780,N_6733);
xnor U7103 (N_7103,N_6633,N_6728);
nor U7104 (N_7104,N_6434,N_6767);
or U7105 (N_7105,N_6585,N_6613);
or U7106 (N_7106,N_6499,N_6672);
nor U7107 (N_7107,N_6542,N_6660);
xor U7108 (N_7108,N_6715,N_6672);
nand U7109 (N_7109,N_6432,N_6506);
and U7110 (N_7110,N_6454,N_6420);
nand U7111 (N_7111,N_6479,N_6718);
nand U7112 (N_7112,N_6569,N_6734);
xor U7113 (N_7113,N_6676,N_6421);
xnor U7114 (N_7114,N_6674,N_6501);
xnor U7115 (N_7115,N_6653,N_6520);
or U7116 (N_7116,N_6522,N_6685);
xor U7117 (N_7117,N_6684,N_6534);
and U7118 (N_7118,N_6672,N_6567);
or U7119 (N_7119,N_6668,N_6561);
nor U7120 (N_7120,N_6573,N_6482);
xor U7121 (N_7121,N_6654,N_6793);
or U7122 (N_7122,N_6796,N_6624);
xor U7123 (N_7123,N_6475,N_6526);
nor U7124 (N_7124,N_6528,N_6588);
or U7125 (N_7125,N_6568,N_6449);
and U7126 (N_7126,N_6416,N_6782);
xnor U7127 (N_7127,N_6760,N_6445);
and U7128 (N_7128,N_6535,N_6550);
nand U7129 (N_7129,N_6676,N_6440);
or U7130 (N_7130,N_6430,N_6758);
nand U7131 (N_7131,N_6754,N_6729);
nor U7132 (N_7132,N_6626,N_6413);
xnor U7133 (N_7133,N_6552,N_6797);
nand U7134 (N_7134,N_6532,N_6626);
nand U7135 (N_7135,N_6592,N_6722);
nor U7136 (N_7136,N_6726,N_6581);
nand U7137 (N_7137,N_6602,N_6434);
xor U7138 (N_7138,N_6705,N_6709);
and U7139 (N_7139,N_6770,N_6600);
nor U7140 (N_7140,N_6764,N_6726);
and U7141 (N_7141,N_6489,N_6793);
xor U7142 (N_7142,N_6434,N_6635);
xor U7143 (N_7143,N_6532,N_6606);
or U7144 (N_7144,N_6626,N_6664);
xnor U7145 (N_7145,N_6793,N_6796);
nand U7146 (N_7146,N_6711,N_6775);
nor U7147 (N_7147,N_6473,N_6783);
nand U7148 (N_7148,N_6629,N_6614);
or U7149 (N_7149,N_6434,N_6704);
nand U7150 (N_7150,N_6598,N_6482);
nor U7151 (N_7151,N_6654,N_6571);
or U7152 (N_7152,N_6407,N_6404);
nor U7153 (N_7153,N_6741,N_6689);
and U7154 (N_7154,N_6759,N_6417);
xnor U7155 (N_7155,N_6677,N_6505);
xor U7156 (N_7156,N_6671,N_6669);
nor U7157 (N_7157,N_6699,N_6410);
and U7158 (N_7158,N_6745,N_6565);
xnor U7159 (N_7159,N_6505,N_6763);
and U7160 (N_7160,N_6560,N_6672);
nor U7161 (N_7161,N_6547,N_6780);
and U7162 (N_7162,N_6465,N_6505);
and U7163 (N_7163,N_6774,N_6531);
and U7164 (N_7164,N_6458,N_6751);
nor U7165 (N_7165,N_6715,N_6578);
or U7166 (N_7166,N_6669,N_6672);
nor U7167 (N_7167,N_6543,N_6577);
or U7168 (N_7168,N_6539,N_6706);
and U7169 (N_7169,N_6585,N_6599);
and U7170 (N_7170,N_6444,N_6740);
xor U7171 (N_7171,N_6483,N_6463);
nand U7172 (N_7172,N_6733,N_6503);
xor U7173 (N_7173,N_6737,N_6703);
and U7174 (N_7174,N_6423,N_6431);
nand U7175 (N_7175,N_6683,N_6472);
or U7176 (N_7176,N_6753,N_6502);
nor U7177 (N_7177,N_6543,N_6615);
and U7178 (N_7178,N_6460,N_6741);
and U7179 (N_7179,N_6780,N_6608);
and U7180 (N_7180,N_6587,N_6671);
nor U7181 (N_7181,N_6510,N_6410);
nand U7182 (N_7182,N_6596,N_6756);
nand U7183 (N_7183,N_6797,N_6795);
nand U7184 (N_7184,N_6413,N_6431);
xnor U7185 (N_7185,N_6759,N_6468);
xnor U7186 (N_7186,N_6566,N_6570);
or U7187 (N_7187,N_6501,N_6795);
and U7188 (N_7188,N_6580,N_6741);
nand U7189 (N_7189,N_6751,N_6689);
xnor U7190 (N_7190,N_6455,N_6581);
nand U7191 (N_7191,N_6622,N_6431);
or U7192 (N_7192,N_6730,N_6442);
xor U7193 (N_7193,N_6717,N_6780);
nor U7194 (N_7194,N_6649,N_6483);
and U7195 (N_7195,N_6679,N_6534);
nand U7196 (N_7196,N_6675,N_6572);
nand U7197 (N_7197,N_6612,N_6799);
and U7198 (N_7198,N_6514,N_6587);
nor U7199 (N_7199,N_6670,N_6437);
nand U7200 (N_7200,N_6801,N_7015);
xnor U7201 (N_7201,N_7080,N_7154);
xnor U7202 (N_7202,N_6956,N_7062);
nand U7203 (N_7203,N_7039,N_7020);
or U7204 (N_7204,N_6996,N_6984);
or U7205 (N_7205,N_7097,N_6883);
nand U7206 (N_7206,N_7198,N_7042);
or U7207 (N_7207,N_6986,N_7123);
nand U7208 (N_7208,N_7094,N_7130);
nand U7209 (N_7209,N_6937,N_7182);
and U7210 (N_7210,N_7171,N_6850);
xor U7211 (N_7211,N_7108,N_6953);
nor U7212 (N_7212,N_7081,N_6822);
or U7213 (N_7213,N_6949,N_7115);
or U7214 (N_7214,N_7033,N_7059);
nor U7215 (N_7215,N_6889,N_7045);
nor U7216 (N_7216,N_6805,N_7168);
xor U7217 (N_7217,N_7193,N_6854);
and U7218 (N_7218,N_7110,N_6947);
and U7219 (N_7219,N_7172,N_6964);
xnor U7220 (N_7220,N_6867,N_7014);
nand U7221 (N_7221,N_6933,N_7149);
or U7222 (N_7222,N_6969,N_7137);
xor U7223 (N_7223,N_7052,N_6966);
nand U7224 (N_7224,N_6897,N_6981);
and U7225 (N_7225,N_7019,N_7109);
or U7226 (N_7226,N_7105,N_6960);
nand U7227 (N_7227,N_6988,N_6987);
xor U7228 (N_7228,N_7099,N_6998);
xor U7229 (N_7229,N_7101,N_6908);
xnor U7230 (N_7230,N_7083,N_6989);
and U7231 (N_7231,N_7030,N_7167);
or U7232 (N_7232,N_7012,N_6838);
or U7233 (N_7233,N_7162,N_6861);
and U7234 (N_7234,N_7046,N_6837);
or U7235 (N_7235,N_7116,N_6863);
and U7236 (N_7236,N_6895,N_6948);
nand U7237 (N_7237,N_6851,N_6823);
nand U7238 (N_7238,N_7128,N_7117);
and U7239 (N_7239,N_7184,N_6979);
nand U7240 (N_7240,N_6888,N_6935);
or U7241 (N_7241,N_6857,N_6971);
nand U7242 (N_7242,N_6865,N_7032);
xnor U7243 (N_7243,N_6923,N_7063);
and U7244 (N_7244,N_7022,N_7009);
and U7245 (N_7245,N_6840,N_6808);
nand U7246 (N_7246,N_6951,N_6967);
nand U7247 (N_7247,N_7164,N_7034);
and U7248 (N_7248,N_6932,N_7112);
nand U7249 (N_7249,N_7031,N_6855);
nand U7250 (N_7250,N_6885,N_6862);
nor U7251 (N_7251,N_7125,N_6802);
nand U7252 (N_7252,N_7102,N_6970);
xor U7253 (N_7253,N_6955,N_7174);
xnor U7254 (N_7254,N_6902,N_6818);
xnor U7255 (N_7255,N_6978,N_6939);
nand U7256 (N_7256,N_6848,N_7160);
nor U7257 (N_7257,N_6982,N_6812);
nor U7258 (N_7258,N_6945,N_6807);
and U7259 (N_7259,N_6990,N_6866);
or U7260 (N_7260,N_7189,N_7197);
or U7261 (N_7261,N_7005,N_6874);
or U7262 (N_7262,N_7138,N_6803);
or U7263 (N_7263,N_6877,N_7131);
nor U7264 (N_7264,N_6907,N_7017);
or U7265 (N_7265,N_7004,N_7175);
xnor U7266 (N_7266,N_6906,N_7078);
xnor U7267 (N_7267,N_6929,N_7120);
xnor U7268 (N_7268,N_6890,N_6963);
or U7269 (N_7269,N_7040,N_6813);
xor U7270 (N_7270,N_7041,N_6809);
nand U7271 (N_7271,N_7106,N_7107);
and U7272 (N_7272,N_7150,N_7098);
xnor U7273 (N_7273,N_7090,N_7181);
nand U7274 (N_7274,N_7087,N_7057);
and U7275 (N_7275,N_6976,N_6903);
or U7276 (N_7276,N_6910,N_6962);
xor U7277 (N_7277,N_6958,N_7124);
nand U7278 (N_7278,N_7143,N_6905);
and U7279 (N_7279,N_7024,N_7023);
nand U7280 (N_7280,N_6881,N_6878);
nor U7281 (N_7281,N_7194,N_6873);
nor U7282 (N_7282,N_6841,N_6849);
and U7283 (N_7283,N_6800,N_6891);
xor U7284 (N_7284,N_7077,N_6938);
nor U7285 (N_7285,N_7111,N_7145);
nor U7286 (N_7286,N_7146,N_6957);
or U7287 (N_7287,N_6968,N_7191);
and U7288 (N_7288,N_7199,N_7163);
nand U7289 (N_7289,N_7104,N_6853);
nor U7290 (N_7290,N_6924,N_6806);
nand U7291 (N_7291,N_7073,N_7076);
xnor U7292 (N_7292,N_7007,N_6992);
xnor U7293 (N_7293,N_6829,N_7096);
nor U7294 (N_7294,N_7066,N_6901);
or U7295 (N_7295,N_6983,N_6927);
nand U7296 (N_7296,N_7013,N_6917);
nor U7297 (N_7297,N_7103,N_6997);
or U7298 (N_7298,N_6920,N_7196);
nor U7299 (N_7299,N_7000,N_7038);
and U7300 (N_7300,N_7173,N_6887);
and U7301 (N_7301,N_7085,N_6961);
nand U7302 (N_7302,N_6944,N_7190);
nand U7303 (N_7303,N_7006,N_6975);
xnor U7304 (N_7304,N_6824,N_7010);
xnor U7305 (N_7305,N_6973,N_7061);
or U7306 (N_7306,N_6959,N_7050);
nor U7307 (N_7307,N_7133,N_6833);
xor U7308 (N_7308,N_7165,N_6814);
nand U7309 (N_7309,N_6915,N_6900);
nor U7310 (N_7310,N_6993,N_7129);
nor U7311 (N_7311,N_7091,N_7113);
and U7312 (N_7312,N_7088,N_7161);
and U7313 (N_7313,N_6875,N_7192);
xnor U7314 (N_7314,N_6804,N_7092);
nor U7315 (N_7315,N_6918,N_7188);
and U7316 (N_7316,N_6810,N_6847);
xor U7317 (N_7317,N_7027,N_6872);
and U7318 (N_7318,N_7127,N_6826);
and U7319 (N_7319,N_7064,N_7028);
and U7320 (N_7320,N_6913,N_7079);
nand U7321 (N_7321,N_6852,N_7074);
and U7322 (N_7322,N_6870,N_6882);
xor U7323 (N_7323,N_6940,N_7100);
nand U7324 (N_7324,N_7089,N_7003);
nor U7325 (N_7325,N_6994,N_7048);
nor U7326 (N_7326,N_7195,N_6842);
and U7327 (N_7327,N_6869,N_6820);
and U7328 (N_7328,N_6819,N_6868);
and U7329 (N_7329,N_7072,N_7139);
xor U7330 (N_7330,N_6934,N_7021);
nand U7331 (N_7331,N_7156,N_7068);
or U7332 (N_7332,N_6928,N_7153);
and U7333 (N_7333,N_7158,N_6912);
xor U7334 (N_7334,N_7086,N_7144);
nand U7335 (N_7335,N_7095,N_6941);
nand U7336 (N_7336,N_7016,N_7141);
nand U7337 (N_7337,N_7140,N_6844);
nor U7338 (N_7338,N_6816,N_6916);
nor U7339 (N_7339,N_7135,N_7037);
nor U7340 (N_7340,N_6950,N_7183);
xnor U7341 (N_7341,N_6884,N_6817);
nand U7342 (N_7342,N_6922,N_7053);
xor U7343 (N_7343,N_6880,N_6921);
nor U7344 (N_7344,N_7029,N_6896);
nand U7345 (N_7345,N_7178,N_7134);
and U7346 (N_7346,N_7049,N_7093);
or U7347 (N_7347,N_6974,N_6836);
nand U7348 (N_7348,N_7122,N_6972);
nor U7349 (N_7349,N_7177,N_6919);
nor U7350 (N_7350,N_6843,N_7008);
nor U7351 (N_7351,N_7114,N_7002);
xnor U7352 (N_7352,N_6835,N_7047);
and U7353 (N_7353,N_7056,N_7155);
and U7354 (N_7354,N_6926,N_6930);
nor U7355 (N_7355,N_7148,N_6943);
xor U7356 (N_7356,N_6931,N_7186);
xor U7357 (N_7357,N_6991,N_7055);
nand U7358 (N_7358,N_6845,N_6898);
and U7359 (N_7359,N_6860,N_6828);
nor U7360 (N_7360,N_7069,N_6980);
nand U7361 (N_7361,N_7170,N_6871);
and U7362 (N_7362,N_6815,N_7018);
and U7363 (N_7363,N_7036,N_7152);
or U7364 (N_7364,N_6894,N_7185);
xnor U7365 (N_7365,N_6831,N_6821);
xnor U7366 (N_7366,N_7157,N_7060);
nor U7367 (N_7367,N_7187,N_6825);
nor U7368 (N_7368,N_7118,N_7082);
nand U7369 (N_7369,N_7179,N_7180);
or U7370 (N_7370,N_6830,N_7065);
nand U7371 (N_7371,N_6954,N_6834);
and U7372 (N_7372,N_6914,N_6859);
and U7373 (N_7373,N_7044,N_7126);
and U7374 (N_7374,N_7121,N_6886);
or U7375 (N_7375,N_7166,N_7119);
nor U7376 (N_7376,N_6925,N_7001);
xor U7377 (N_7377,N_6999,N_7136);
xnor U7378 (N_7378,N_6811,N_6858);
nand U7379 (N_7379,N_6952,N_6936);
xnor U7380 (N_7380,N_7067,N_7025);
xnor U7381 (N_7381,N_6892,N_7151);
and U7382 (N_7382,N_6846,N_6946);
or U7383 (N_7383,N_6899,N_7058);
and U7384 (N_7384,N_7035,N_7142);
or U7385 (N_7385,N_6965,N_7169);
nor U7386 (N_7386,N_6839,N_6985);
xnor U7387 (N_7387,N_7071,N_7011);
and U7388 (N_7388,N_6893,N_6832);
xor U7389 (N_7389,N_7070,N_7159);
or U7390 (N_7390,N_7054,N_6909);
nand U7391 (N_7391,N_6995,N_6879);
and U7392 (N_7392,N_7147,N_6864);
xnor U7393 (N_7393,N_7075,N_7043);
nand U7394 (N_7394,N_6904,N_7176);
or U7395 (N_7395,N_6911,N_6977);
or U7396 (N_7396,N_7026,N_6827);
and U7397 (N_7397,N_7051,N_6876);
nor U7398 (N_7398,N_6942,N_7132);
and U7399 (N_7399,N_7084,N_6856);
xor U7400 (N_7400,N_7051,N_7056);
and U7401 (N_7401,N_6849,N_7041);
nand U7402 (N_7402,N_7132,N_6975);
and U7403 (N_7403,N_7070,N_7101);
nor U7404 (N_7404,N_7136,N_7158);
xnor U7405 (N_7405,N_7153,N_7040);
and U7406 (N_7406,N_6988,N_6817);
nor U7407 (N_7407,N_6923,N_6827);
nand U7408 (N_7408,N_7188,N_7151);
and U7409 (N_7409,N_6983,N_6965);
xor U7410 (N_7410,N_7037,N_6924);
or U7411 (N_7411,N_7102,N_7139);
xor U7412 (N_7412,N_7155,N_6907);
nor U7413 (N_7413,N_7145,N_7158);
nor U7414 (N_7414,N_6979,N_7109);
nor U7415 (N_7415,N_7072,N_6847);
nand U7416 (N_7416,N_7074,N_6866);
and U7417 (N_7417,N_6963,N_7159);
nor U7418 (N_7418,N_7092,N_7021);
nor U7419 (N_7419,N_7017,N_7097);
nand U7420 (N_7420,N_6848,N_7061);
and U7421 (N_7421,N_7097,N_6813);
and U7422 (N_7422,N_6916,N_6865);
and U7423 (N_7423,N_6955,N_6909);
and U7424 (N_7424,N_6917,N_6914);
xnor U7425 (N_7425,N_7107,N_6857);
xnor U7426 (N_7426,N_6923,N_6931);
and U7427 (N_7427,N_7110,N_7183);
or U7428 (N_7428,N_6997,N_7022);
xor U7429 (N_7429,N_6824,N_7089);
nand U7430 (N_7430,N_7168,N_7022);
or U7431 (N_7431,N_6985,N_6909);
nand U7432 (N_7432,N_7094,N_6869);
xnor U7433 (N_7433,N_7014,N_7114);
nor U7434 (N_7434,N_7192,N_7094);
and U7435 (N_7435,N_6923,N_7175);
and U7436 (N_7436,N_6822,N_7110);
nor U7437 (N_7437,N_6886,N_6824);
or U7438 (N_7438,N_6961,N_7100);
nand U7439 (N_7439,N_6911,N_6903);
nand U7440 (N_7440,N_6953,N_7067);
or U7441 (N_7441,N_6955,N_7060);
and U7442 (N_7442,N_7034,N_7112);
nand U7443 (N_7443,N_6825,N_6945);
and U7444 (N_7444,N_6897,N_6960);
xnor U7445 (N_7445,N_7139,N_7130);
nand U7446 (N_7446,N_7043,N_6918);
xnor U7447 (N_7447,N_6828,N_6994);
nor U7448 (N_7448,N_7140,N_6823);
xor U7449 (N_7449,N_6834,N_7138);
nand U7450 (N_7450,N_7187,N_7134);
nor U7451 (N_7451,N_6851,N_7021);
nand U7452 (N_7452,N_7146,N_6840);
or U7453 (N_7453,N_7151,N_6852);
nor U7454 (N_7454,N_7143,N_6869);
nand U7455 (N_7455,N_7046,N_7140);
or U7456 (N_7456,N_6994,N_6972);
nor U7457 (N_7457,N_6990,N_6999);
xor U7458 (N_7458,N_7134,N_7045);
nand U7459 (N_7459,N_6999,N_7158);
xor U7460 (N_7460,N_7021,N_7148);
xnor U7461 (N_7461,N_7121,N_6903);
nand U7462 (N_7462,N_6817,N_6869);
xor U7463 (N_7463,N_7100,N_6959);
or U7464 (N_7464,N_7108,N_7142);
nand U7465 (N_7465,N_6989,N_6966);
xnor U7466 (N_7466,N_7096,N_7000);
and U7467 (N_7467,N_7026,N_7062);
nand U7468 (N_7468,N_6853,N_6955);
nor U7469 (N_7469,N_6829,N_7055);
or U7470 (N_7470,N_7092,N_7127);
xnor U7471 (N_7471,N_6801,N_6964);
and U7472 (N_7472,N_7172,N_7118);
nor U7473 (N_7473,N_7142,N_7152);
xor U7474 (N_7474,N_6877,N_6829);
xnor U7475 (N_7475,N_6993,N_6898);
or U7476 (N_7476,N_7097,N_7133);
and U7477 (N_7477,N_6856,N_6900);
nor U7478 (N_7478,N_6849,N_7136);
nor U7479 (N_7479,N_6850,N_6916);
xor U7480 (N_7480,N_6934,N_7060);
nor U7481 (N_7481,N_7133,N_7186);
or U7482 (N_7482,N_7111,N_7194);
and U7483 (N_7483,N_6819,N_6848);
nor U7484 (N_7484,N_7018,N_7073);
xor U7485 (N_7485,N_7175,N_7135);
or U7486 (N_7486,N_7035,N_6974);
and U7487 (N_7487,N_6931,N_6818);
nor U7488 (N_7488,N_7172,N_7024);
nand U7489 (N_7489,N_7107,N_7032);
nor U7490 (N_7490,N_7060,N_6839);
and U7491 (N_7491,N_7138,N_6827);
or U7492 (N_7492,N_7142,N_7016);
and U7493 (N_7493,N_6814,N_6971);
nand U7494 (N_7494,N_7171,N_6937);
nand U7495 (N_7495,N_7036,N_7039);
nor U7496 (N_7496,N_6949,N_7181);
nand U7497 (N_7497,N_7015,N_7181);
xnor U7498 (N_7498,N_6975,N_7012);
or U7499 (N_7499,N_6920,N_7047);
nand U7500 (N_7500,N_6935,N_7113);
or U7501 (N_7501,N_6823,N_7055);
or U7502 (N_7502,N_6888,N_6841);
nor U7503 (N_7503,N_6800,N_6833);
nand U7504 (N_7504,N_6855,N_6806);
xor U7505 (N_7505,N_7039,N_6837);
and U7506 (N_7506,N_6955,N_7172);
or U7507 (N_7507,N_6885,N_7131);
nand U7508 (N_7508,N_7175,N_7132);
nor U7509 (N_7509,N_6881,N_6814);
and U7510 (N_7510,N_7040,N_6900);
nor U7511 (N_7511,N_6871,N_6925);
and U7512 (N_7512,N_6804,N_6969);
and U7513 (N_7513,N_6804,N_7109);
and U7514 (N_7514,N_7110,N_6974);
nand U7515 (N_7515,N_7180,N_7111);
nand U7516 (N_7516,N_7039,N_6817);
xnor U7517 (N_7517,N_6875,N_6958);
or U7518 (N_7518,N_6841,N_6945);
nor U7519 (N_7519,N_6934,N_6999);
xnor U7520 (N_7520,N_7137,N_7057);
xor U7521 (N_7521,N_6952,N_7109);
nand U7522 (N_7522,N_7157,N_7102);
nor U7523 (N_7523,N_7033,N_6804);
nor U7524 (N_7524,N_7107,N_7020);
and U7525 (N_7525,N_6928,N_6828);
xor U7526 (N_7526,N_6991,N_6904);
and U7527 (N_7527,N_7143,N_6902);
nand U7528 (N_7528,N_6901,N_6980);
and U7529 (N_7529,N_7003,N_7166);
nor U7530 (N_7530,N_6956,N_6993);
xor U7531 (N_7531,N_6978,N_7125);
or U7532 (N_7532,N_7038,N_6928);
nor U7533 (N_7533,N_7012,N_6806);
or U7534 (N_7534,N_6963,N_6969);
or U7535 (N_7535,N_7194,N_7120);
or U7536 (N_7536,N_7153,N_7194);
nor U7537 (N_7537,N_7001,N_7185);
nand U7538 (N_7538,N_6902,N_6850);
nor U7539 (N_7539,N_7044,N_6919);
nor U7540 (N_7540,N_7073,N_6801);
nor U7541 (N_7541,N_6921,N_6905);
xnor U7542 (N_7542,N_6809,N_7030);
or U7543 (N_7543,N_7168,N_7086);
nor U7544 (N_7544,N_6998,N_7122);
nor U7545 (N_7545,N_7132,N_7062);
nand U7546 (N_7546,N_6974,N_6940);
nand U7547 (N_7547,N_6838,N_7035);
xor U7548 (N_7548,N_7059,N_6817);
or U7549 (N_7549,N_6801,N_7022);
or U7550 (N_7550,N_7151,N_7170);
xnor U7551 (N_7551,N_6944,N_7134);
nand U7552 (N_7552,N_7037,N_7170);
or U7553 (N_7553,N_6856,N_6941);
or U7554 (N_7554,N_6984,N_7170);
or U7555 (N_7555,N_6991,N_7024);
nor U7556 (N_7556,N_6992,N_7171);
nand U7557 (N_7557,N_7171,N_7199);
nor U7558 (N_7558,N_6820,N_6874);
and U7559 (N_7559,N_6837,N_6917);
nand U7560 (N_7560,N_6957,N_7094);
nand U7561 (N_7561,N_7047,N_6960);
nand U7562 (N_7562,N_7096,N_7178);
and U7563 (N_7563,N_7076,N_6996);
nor U7564 (N_7564,N_6928,N_6913);
and U7565 (N_7565,N_7180,N_6994);
nand U7566 (N_7566,N_7028,N_7038);
or U7567 (N_7567,N_6912,N_7192);
nand U7568 (N_7568,N_6950,N_7175);
xor U7569 (N_7569,N_6948,N_6854);
xor U7570 (N_7570,N_6836,N_6853);
xnor U7571 (N_7571,N_6932,N_6930);
nand U7572 (N_7572,N_6830,N_6829);
or U7573 (N_7573,N_6816,N_6957);
or U7574 (N_7574,N_6856,N_6871);
or U7575 (N_7575,N_6810,N_6895);
and U7576 (N_7576,N_7035,N_7076);
and U7577 (N_7577,N_6964,N_7117);
and U7578 (N_7578,N_6896,N_7126);
and U7579 (N_7579,N_6801,N_6840);
nand U7580 (N_7580,N_7045,N_6955);
nor U7581 (N_7581,N_7028,N_6910);
nor U7582 (N_7582,N_7111,N_6944);
nor U7583 (N_7583,N_6889,N_6974);
xnor U7584 (N_7584,N_7161,N_6803);
xnor U7585 (N_7585,N_7007,N_7154);
or U7586 (N_7586,N_7139,N_7191);
or U7587 (N_7587,N_6875,N_7060);
and U7588 (N_7588,N_7010,N_7198);
nor U7589 (N_7589,N_7112,N_6838);
xnor U7590 (N_7590,N_7150,N_7036);
xnor U7591 (N_7591,N_7133,N_6901);
nor U7592 (N_7592,N_7044,N_6881);
and U7593 (N_7593,N_7090,N_6950);
xor U7594 (N_7594,N_7059,N_6970);
and U7595 (N_7595,N_6922,N_7155);
xor U7596 (N_7596,N_7038,N_7036);
and U7597 (N_7597,N_6989,N_6955);
and U7598 (N_7598,N_6812,N_7087);
and U7599 (N_7599,N_7133,N_7043);
or U7600 (N_7600,N_7474,N_7343);
nor U7601 (N_7601,N_7454,N_7419);
nor U7602 (N_7602,N_7416,N_7405);
nor U7603 (N_7603,N_7308,N_7272);
and U7604 (N_7604,N_7337,N_7313);
nor U7605 (N_7605,N_7213,N_7373);
or U7606 (N_7606,N_7513,N_7567);
and U7607 (N_7607,N_7459,N_7326);
and U7608 (N_7608,N_7336,N_7374);
nand U7609 (N_7609,N_7330,N_7526);
or U7610 (N_7610,N_7582,N_7576);
and U7611 (N_7611,N_7312,N_7227);
nor U7612 (N_7612,N_7387,N_7208);
and U7613 (N_7613,N_7475,N_7569);
and U7614 (N_7614,N_7445,N_7452);
and U7615 (N_7615,N_7252,N_7578);
and U7616 (N_7616,N_7339,N_7575);
xnor U7617 (N_7617,N_7568,N_7270);
nor U7618 (N_7618,N_7243,N_7372);
or U7619 (N_7619,N_7542,N_7429);
nor U7620 (N_7620,N_7306,N_7255);
xor U7621 (N_7621,N_7344,N_7433);
nor U7622 (N_7622,N_7586,N_7281);
xnor U7623 (N_7623,N_7523,N_7477);
or U7624 (N_7624,N_7497,N_7489);
nor U7625 (N_7625,N_7555,N_7463);
or U7626 (N_7626,N_7359,N_7241);
or U7627 (N_7627,N_7515,N_7324);
xnor U7628 (N_7628,N_7398,N_7464);
or U7629 (N_7629,N_7540,N_7534);
or U7630 (N_7630,N_7351,N_7211);
nor U7631 (N_7631,N_7260,N_7558);
or U7632 (N_7632,N_7520,N_7266);
and U7633 (N_7633,N_7277,N_7380);
and U7634 (N_7634,N_7206,N_7212);
nand U7635 (N_7635,N_7573,N_7323);
nand U7636 (N_7636,N_7299,N_7381);
xor U7637 (N_7637,N_7476,N_7244);
nor U7638 (N_7638,N_7462,N_7483);
nor U7639 (N_7639,N_7551,N_7508);
or U7640 (N_7640,N_7317,N_7396);
nor U7641 (N_7641,N_7221,N_7570);
xnor U7642 (N_7642,N_7547,N_7450);
or U7643 (N_7643,N_7358,N_7302);
nor U7644 (N_7644,N_7493,N_7298);
and U7645 (N_7645,N_7512,N_7559);
nand U7646 (N_7646,N_7203,N_7538);
nand U7647 (N_7647,N_7282,N_7407);
nand U7648 (N_7648,N_7517,N_7552);
and U7649 (N_7649,N_7492,N_7403);
nor U7650 (N_7650,N_7311,N_7253);
or U7651 (N_7651,N_7451,N_7401);
and U7652 (N_7652,N_7283,N_7356);
or U7653 (N_7653,N_7516,N_7415);
nand U7654 (N_7654,N_7402,N_7362);
or U7655 (N_7655,N_7305,N_7245);
or U7656 (N_7656,N_7292,N_7329);
nor U7657 (N_7657,N_7465,N_7242);
nand U7658 (N_7658,N_7502,N_7393);
nor U7659 (N_7659,N_7361,N_7310);
xor U7660 (N_7660,N_7456,N_7335);
nand U7661 (N_7661,N_7406,N_7368);
and U7662 (N_7662,N_7594,N_7455);
and U7663 (N_7663,N_7511,N_7446);
nand U7664 (N_7664,N_7322,N_7333);
xor U7665 (N_7665,N_7434,N_7400);
xnor U7666 (N_7666,N_7413,N_7467);
xor U7667 (N_7667,N_7224,N_7265);
nor U7668 (N_7668,N_7522,N_7580);
nand U7669 (N_7669,N_7409,N_7458);
nand U7670 (N_7670,N_7595,N_7593);
or U7671 (N_7671,N_7423,N_7314);
nor U7672 (N_7672,N_7514,N_7490);
xnor U7673 (N_7673,N_7519,N_7363);
nand U7674 (N_7674,N_7597,N_7447);
xor U7675 (N_7675,N_7531,N_7325);
nand U7676 (N_7676,N_7533,N_7591);
nand U7677 (N_7677,N_7436,N_7529);
or U7678 (N_7678,N_7544,N_7566);
nand U7679 (N_7679,N_7438,N_7577);
nor U7680 (N_7680,N_7288,N_7411);
nand U7681 (N_7681,N_7205,N_7556);
or U7682 (N_7682,N_7262,N_7285);
and U7683 (N_7683,N_7386,N_7294);
or U7684 (N_7684,N_7496,N_7259);
and U7685 (N_7685,N_7439,N_7318);
nand U7686 (N_7686,N_7261,N_7300);
nand U7687 (N_7687,N_7448,N_7338);
xor U7688 (N_7688,N_7367,N_7412);
xnor U7689 (N_7689,N_7204,N_7371);
and U7690 (N_7690,N_7506,N_7315);
nor U7691 (N_7691,N_7369,N_7341);
nand U7692 (N_7692,N_7440,N_7479);
nand U7693 (N_7693,N_7276,N_7420);
and U7694 (N_7694,N_7596,N_7530);
and U7695 (N_7695,N_7414,N_7364);
nand U7696 (N_7696,N_7236,N_7257);
and U7697 (N_7697,N_7388,N_7494);
nand U7698 (N_7698,N_7256,N_7360);
or U7699 (N_7699,N_7349,N_7537);
or U7700 (N_7700,N_7268,N_7543);
xnor U7701 (N_7701,N_7382,N_7592);
and U7702 (N_7702,N_7331,N_7353);
xnor U7703 (N_7703,N_7421,N_7482);
and U7704 (N_7704,N_7327,N_7307);
xnor U7705 (N_7705,N_7539,N_7428);
and U7706 (N_7706,N_7304,N_7215);
nand U7707 (N_7707,N_7491,N_7470);
nor U7708 (N_7708,N_7488,N_7549);
nand U7709 (N_7709,N_7233,N_7425);
xor U7710 (N_7710,N_7590,N_7460);
or U7711 (N_7711,N_7354,N_7525);
nand U7712 (N_7712,N_7218,N_7340);
xor U7713 (N_7713,N_7246,N_7478);
nand U7714 (N_7714,N_7527,N_7541);
or U7715 (N_7715,N_7395,N_7202);
nand U7716 (N_7716,N_7442,N_7279);
xor U7717 (N_7717,N_7426,N_7377);
and U7718 (N_7718,N_7225,N_7301);
nor U7719 (N_7719,N_7507,N_7210);
nand U7720 (N_7720,N_7437,N_7303);
nand U7721 (N_7721,N_7269,N_7365);
and U7722 (N_7722,N_7278,N_7319);
nor U7723 (N_7723,N_7498,N_7274);
and U7724 (N_7724,N_7471,N_7287);
nand U7725 (N_7725,N_7200,N_7560);
xnor U7726 (N_7726,N_7226,N_7286);
nand U7727 (N_7727,N_7275,N_7391);
xnor U7728 (N_7728,N_7589,N_7528);
and U7729 (N_7729,N_7410,N_7284);
nand U7730 (N_7730,N_7342,N_7431);
or U7731 (N_7731,N_7532,N_7487);
or U7732 (N_7732,N_7267,N_7562);
nand U7733 (N_7733,N_7444,N_7348);
or U7734 (N_7734,N_7584,N_7320);
nor U7735 (N_7735,N_7316,N_7554);
xnor U7736 (N_7736,N_7404,N_7220);
nor U7737 (N_7737,N_7505,N_7378);
nor U7738 (N_7738,N_7214,N_7545);
nor U7739 (N_7739,N_7232,N_7328);
nor U7740 (N_7740,N_7443,N_7290);
and U7741 (N_7741,N_7579,N_7352);
and U7742 (N_7742,N_7418,N_7536);
nand U7743 (N_7743,N_7397,N_7469);
xor U7744 (N_7744,N_7441,N_7231);
or U7745 (N_7745,N_7346,N_7557);
and U7746 (N_7746,N_7384,N_7435);
and U7747 (N_7747,N_7501,N_7553);
or U7748 (N_7748,N_7347,N_7563);
xnor U7749 (N_7749,N_7295,N_7357);
or U7750 (N_7750,N_7366,N_7289);
and U7751 (N_7751,N_7585,N_7237);
nor U7752 (N_7752,N_7535,N_7238);
and U7753 (N_7753,N_7422,N_7217);
or U7754 (N_7754,N_7332,N_7546);
xnor U7755 (N_7755,N_7223,N_7499);
or U7756 (N_7756,N_7263,N_7375);
or U7757 (N_7757,N_7510,N_7249);
nor U7758 (N_7758,N_7430,N_7209);
nor U7759 (N_7759,N_7258,N_7548);
nor U7760 (N_7760,N_7500,N_7355);
nand U7761 (N_7761,N_7234,N_7229);
nor U7762 (N_7762,N_7504,N_7427);
xnor U7763 (N_7763,N_7503,N_7222);
nand U7764 (N_7764,N_7370,N_7457);
nor U7765 (N_7765,N_7432,N_7468);
xor U7766 (N_7766,N_7207,N_7296);
and U7767 (N_7767,N_7521,N_7385);
nor U7768 (N_7768,N_7550,N_7473);
xor U7769 (N_7769,N_7309,N_7219);
xnor U7770 (N_7770,N_7581,N_7564);
nand U7771 (N_7771,N_7273,N_7518);
nor U7772 (N_7772,N_7389,N_7571);
or U7773 (N_7773,N_7399,N_7588);
nand U7774 (N_7774,N_7583,N_7250);
and U7775 (N_7775,N_7481,N_7264);
xor U7776 (N_7776,N_7247,N_7461);
nand U7777 (N_7777,N_7392,N_7321);
and U7778 (N_7778,N_7472,N_7254);
or U7779 (N_7779,N_7291,N_7235);
or U7780 (N_7780,N_7293,N_7248);
nand U7781 (N_7781,N_7383,N_7201);
nand U7782 (N_7782,N_7376,N_7280);
nand U7783 (N_7783,N_7572,N_7598);
xnor U7784 (N_7784,N_7449,N_7524);
or U7785 (N_7785,N_7350,N_7509);
and U7786 (N_7786,N_7239,N_7453);
nor U7787 (N_7787,N_7561,N_7230);
nor U7788 (N_7788,N_7271,N_7574);
xor U7789 (N_7789,N_7486,N_7228);
or U7790 (N_7790,N_7345,N_7297);
and U7791 (N_7791,N_7408,N_7394);
and U7792 (N_7792,N_7424,N_7485);
or U7793 (N_7793,N_7216,N_7379);
or U7794 (N_7794,N_7334,N_7599);
and U7795 (N_7795,N_7390,N_7565);
and U7796 (N_7796,N_7240,N_7495);
or U7797 (N_7797,N_7480,N_7466);
nand U7798 (N_7798,N_7587,N_7484);
or U7799 (N_7799,N_7417,N_7251);
and U7800 (N_7800,N_7249,N_7524);
nand U7801 (N_7801,N_7543,N_7219);
nor U7802 (N_7802,N_7507,N_7475);
and U7803 (N_7803,N_7556,N_7315);
nand U7804 (N_7804,N_7564,N_7327);
nor U7805 (N_7805,N_7475,N_7547);
nand U7806 (N_7806,N_7568,N_7359);
xor U7807 (N_7807,N_7536,N_7538);
nand U7808 (N_7808,N_7471,N_7313);
or U7809 (N_7809,N_7271,N_7303);
or U7810 (N_7810,N_7392,N_7278);
nand U7811 (N_7811,N_7232,N_7264);
nor U7812 (N_7812,N_7427,N_7428);
nor U7813 (N_7813,N_7282,N_7250);
and U7814 (N_7814,N_7244,N_7262);
nor U7815 (N_7815,N_7586,N_7576);
or U7816 (N_7816,N_7378,N_7514);
xnor U7817 (N_7817,N_7396,N_7437);
xor U7818 (N_7818,N_7513,N_7287);
and U7819 (N_7819,N_7335,N_7415);
xor U7820 (N_7820,N_7201,N_7252);
nand U7821 (N_7821,N_7292,N_7333);
nor U7822 (N_7822,N_7249,N_7459);
xor U7823 (N_7823,N_7389,N_7309);
or U7824 (N_7824,N_7529,N_7453);
nor U7825 (N_7825,N_7323,N_7264);
or U7826 (N_7826,N_7233,N_7232);
and U7827 (N_7827,N_7364,N_7528);
xor U7828 (N_7828,N_7243,N_7584);
nand U7829 (N_7829,N_7421,N_7334);
nor U7830 (N_7830,N_7508,N_7366);
xnor U7831 (N_7831,N_7452,N_7377);
xor U7832 (N_7832,N_7255,N_7456);
nor U7833 (N_7833,N_7291,N_7389);
or U7834 (N_7834,N_7219,N_7204);
nand U7835 (N_7835,N_7523,N_7451);
xor U7836 (N_7836,N_7545,N_7252);
nand U7837 (N_7837,N_7473,N_7552);
nand U7838 (N_7838,N_7499,N_7284);
nor U7839 (N_7839,N_7264,N_7421);
nand U7840 (N_7840,N_7453,N_7216);
nand U7841 (N_7841,N_7425,N_7565);
nor U7842 (N_7842,N_7510,N_7563);
xor U7843 (N_7843,N_7452,N_7592);
or U7844 (N_7844,N_7413,N_7395);
and U7845 (N_7845,N_7364,N_7527);
nand U7846 (N_7846,N_7320,N_7293);
xor U7847 (N_7847,N_7445,N_7549);
nor U7848 (N_7848,N_7490,N_7533);
and U7849 (N_7849,N_7294,N_7222);
nor U7850 (N_7850,N_7401,N_7326);
nand U7851 (N_7851,N_7583,N_7561);
and U7852 (N_7852,N_7271,N_7352);
nor U7853 (N_7853,N_7418,N_7224);
or U7854 (N_7854,N_7230,N_7389);
nand U7855 (N_7855,N_7252,N_7416);
or U7856 (N_7856,N_7406,N_7216);
and U7857 (N_7857,N_7322,N_7283);
and U7858 (N_7858,N_7299,N_7380);
or U7859 (N_7859,N_7365,N_7248);
or U7860 (N_7860,N_7245,N_7241);
or U7861 (N_7861,N_7464,N_7518);
or U7862 (N_7862,N_7595,N_7271);
nand U7863 (N_7863,N_7598,N_7336);
and U7864 (N_7864,N_7497,N_7316);
nor U7865 (N_7865,N_7323,N_7349);
nand U7866 (N_7866,N_7439,N_7492);
nand U7867 (N_7867,N_7210,N_7434);
and U7868 (N_7868,N_7247,N_7221);
nand U7869 (N_7869,N_7497,N_7230);
or U7870 (N_7870,N_7522,N_7508);
or U7871 (N_7871,N_7455,N_7519);
and U7872 (N_7872,N_7407,N_7207);
xnor U7873 (N_7873,N_7467,N_7556);
nor U7874 (N_7874,N_7462,N_7578);
xor U7875 (N_7875,N_7270,N_7292);
or U7876 (N_7876,N_7259,N_7284);
nor U7877 (N_7877,N_7308,N_7596);
and U7878 (N_7878,N_7570,N_7573);
xnor U7879 (N_7879,N_7474,N_7414);
nor U7880 (N_7880,N_7400,N_7257);
nor U7881 (N_7881,N_7582,N_7446);
nand U7882 (N_7882,N_7371,N_7486);
and U7883 (N_7883,N_7394,N_7533);
or U7884 (N_7884,N_7466,N_7587);
xor U7885 (N_7885,N_7217,N_7479);
nor U7886 (N_7886,N_7223,N_7303);
nand U7887 (N_7887,N_7580,N_7298);
nand U7888 (N_7888,N_7448,N_7233);
nand U7889 (N_7889,N_7335,N_7292);
or U7890 (N_7890,N_7231,N_7552);
nand U7891 (N_7891,N_7584,N_7270);
nand U7892 (N_7892,N_7239,N_7489);
nand U7893 (N_7893,N_7522,N_7390);
and U7894 (N_7894,N_7203,N_7238);
xor U7895 (N_7895,N_7598,N_7587);
nand U7896 (N_7896,N_7458,N_7235);
nand U7897 (N_7897,N_7467,N_7262);
and U7898 (N_7898,N_7214,N_7250);
or U7899 (N_7899,N_7491,N_7333);
and U7900 (N_7900,N_7587,N_7581);
or U7901 (N_7901,N_7537,N_7576);
and U7902 (N_7902,N_7293,N_7478);
or U7903 (N_7903,N_7398,N_7449);
xor U7904 (N_7904,N_7384,N_7596);
and U7905 (N_7905,N_7200,N_7452);
nor U7906 (N_7906,N_7589,N_7240);
or U7907 (N_7907,N_7336,N_7248);
nand U7908 (N_7908,N_7429,N_7488);
or U7909 (N_7909,N_7396,N_7292);
nor U7910 (N_7910,N_7261,N_7580);
or U7911 (N_7911,N_7523,N_7273);
and U7912 (N_7912,N_7322,N_7469);
nor U7913 (N_7913,N_7490,N_7487);
and U7914 (N_7914,N_7543,N_7591);
nand U7915 (N_7915,N_7448,N_7240);
and U7916 (N_7916,N_7221,N_7524);
or U7917 (N_7917,N_7463,N_7383);
or U7918 (N_7918,N_7427,N_7279);
and U7919 (N_7919,N_7390,N_7575);
nand U7920 (N_7920,N_7287,N_7413);
nor U7921 (N_7921,N_7247,N_7553);
or U7922 (N_7922,N_7337,N_7459);
and U7923 (N_7923,N_7240,N_7344);
nor U7924 (N_7924,N_7578,N_7395);
xor U7925 (N_7925,N_7469,N_7276);
xnor U7926 (N_7926,N_7537,N_7201);
nand U7927 (N_7927,N_7555,N_7580);
xnor U7928 (N_7928,N_7289,N_7515);
xor U7929 (N_7929,N_7598,N_7484);
nand U7930 (N_7930,N_7535,N_7250);
or U7931 (N_7931,N_7518,N_7205);
nand U7932 (N_7932,N_7559,N_7572);
or U7933 (N_7933,N_7558,N_7253);
xnor U7934 (N_7934,N_7530,N_7583);
and U7935 (N_7935,N_7487,N_7365);
and U7936 (N_7936,N_7206,N_7445);
nor U7937 (N_7937,N_7597,N_7410);
nor U7938 (N_7938,N_7310,N_7529);
nand U7939 (N_7939,N_7499,N_7368);
or U7940 (N_7940,N_7420,N_7584);
nor U7941 (N_7941,N_7473,N_7409);
xnor U7942 (N_7942,N_7321,N_7305);
nand U7943 (N_7943,N_7277,N_7587);
nor U7944 (N_7944,N_7272,N_7493);
xnor U7945 (N_7945,N_7408,N_7346);
xnor U7946 (N_7946,N_7467,N_7512);
nor U7947 (N_7947,N_7329,N_7525);
xnor U7948 (N_7948,N_7218,N_7227);
nand U7949 (N_7949,N_7449,N_7241);
nand U7950 (N_7950,N_7585,N_7333);
xor U7951 (N_7951,N_7411,N_7502);
nand U7952 (N_7952,N_7210,N_7411);
and U7953 (N_7953,N_7463,N_7350);
xor U7954 (N_7954,N_7293,N_7249);
nand U7955 (N_7955,N_7594,N_7225);
or U7956 (N_7956,N_7348,N_7434);
nor U7957 (N_7957,N_7502,N_7463);
xnor U7958 (N_7958,N_7242,N_7584);
and U7959 (N_7959,N_7325,N_7495);
nor U7960 (N_7960,N_7290,N_7532);
nor U7961 (N_7961,N_7449,N_7573);
xor U7962 (N_7962,N_7487,N_7374);
and U7963 (N_7963,N_7494,N_7414);
nor U7964 (N_7964,N_7379,N_7275);
xnor U7965 (N_7965,N_7351,N_7253);
or U7966 (N_7966,N_7578,N_7452);
and U7967 (N_7967,N_7351,N_7305);
nor U7968 (N_7968,N_7251,N_7441);
nor U7969 (N_7969,N_7286,N_7550);
nand U7970 (N_7970,N_7362,N_7305);
and U7971 (N_7971,N_7516,N_7228);
xor U7972 (N_7972,N_7481,N_7550);
nor U7973 (N_7973,N_7233,N_7487);
nand U7974 (N_7974,N_7582,N_7381);
nand U7975 (N_7975,N_7263,N_7388);
or U7976 (N_7976,N_7353,N_7576);
and U7977 (N_7977,N_7473,N_7271);
and U7978 (N_7978,N_7527,N_7315);
and U7979 (N_7979,N_7343,N_7425);
nand U7980 (N_7980,N_7582,N_7424);
nor U7981 (N_7981,N_7354,N_7580);
or U7982 (N_7982,N_7439,N_7265);
or U7983 (N_7983,N_7216,N_7205);
xnor U7984 (N_7984,N_7547,N_7323);
and U7985 (N_7985,N_7222,N_7269);
xnor U7986 (N_7986,N_7406,N_7551);
nand U7987 (N_7987,N_7468,N_7247);
xnor U7988 (N_7988,N_7261,N_7382);
or U7989 (N_7989,N_7380,N_7585);
xor U7990 (N_7990,N_7263,N_7562);
nand U7991 (N_7991,N_7352,N_7230);
and U7992 (N_7992,N_7355,N_7257);
and U7993 (N_7993,N_7503,N_7324);
nand U7994 (N_7994,N_7313,N_7388);
nand U7995 (N_7995,N_7333,N_7279);
and U7996 (N_7996,N_7557,N_7295);
xor U7997 (N_7997,N_7347,N_7486);
or U7998 (N_7998,N_7231,N_7224);
nor U7999 (N_7999,N_7253,N_7448);
nor U8000 (N_8000,N_7723,N_7714);
xor U8001 (N_8001,N_7809,N_7676);
or U8002 (N_8002,N_7709,N_7825);
xor U8003 (N_8003,N_7936,N_7941);
xnor U8004 (N_8004,N_7786,N_7744);
xor U8005 (N_8005,N_7696,N_7679);
nand U8006 (N_8006,N_7707,N_7962);
or U8007 (N_8007,N_7894,N_7717);
xor U8008 (N_8008,N_7913,N_7953);
and U8009 (N_8009,N_7779,N_7728);
xor U8010 (N_8010,N_7831,N_7955);
or U8011 (N_8011,N_7691,N_7908);
and U8012 (N_8012,N_7887,N_7731);
or U8013 (N_8013,N_7802,N_7788);
and U8014 (N_8014,N_7920,N_7938);
or U8015 (N_8015,N_7946,N_7862);
or U8016 (N_8016,N_7857,N_7973);
xnor U8017 (N_8017,N_7865,N_7641);
and U8018 (N_8018,N_7890,N_7912);
nor U8019 (N_8019,N_7740,N_7984);
and U8020 (N_8020,N_7943,N_7839);
or U8021 (N_8021,N_7932,N_7898);
or U8022 (N_8022,N_7929,N_7643);
or U8023 (N_8023,N_7860,N_7609);
nand U8024 (N_8024,N_7937,N_7636);
or U8025 (N_8025,N_7949,N_7611);
nand U8026 (N_8026,N_7896,N_7944);
nor U8027 (N_8027,N_7652,N_7852);
nor U8028 (N_8028,N_7766,N_7735);
or U8029 (N_8029,N_7759,N_7749);
and U8030 (N_8030,N_7686,N_7859);
or U8031 (N_8031,N_7764,N_7746);
nand U8032 (N_8032,N_7952,N_7732);
nand U8033 (N_8033,N_7800,N_7876);
and U8034 (N_8034,N_7813,N_7902);
and U8035 (N_8035,N_7635,N_7989);
or U8036 (N_8036,N_7789,N_7905);
nor U8037 (N_8037,N_7924,N_7725);
or U8038 (N_8038,N_7647,N_7660);
nand U8039 (N_8039,N_7910,N_7903);
or U8040 (N_8040,N_7971,N_7982);
nor U8041 (N_8041,N_7607,N_7718);
nor U8042 (N_8042,N_7904,N_7730);
and U8043 (N_8043,N_7870,N_7947);
or U8044 (N_8044,N_7666,N_7968);
xor U8045 (N_8045,N_7958,N_7794);
and U8046 (N_8046,N_7710,N_7754);
nand U8047 (N_8047,N_7604,N_7790);
and U8048 (N_8048,N_7842,N_7621);
xnor U8049 (N_8049,N_7614,N_7770);
nand U8050 (N_8050,N_7922,N_7995);
or U8051 (N_8051,N_7771,N_7806);
and U8052 (N_8052,N_7617,N_7756);
and U8053 (N_8053,N_7954,N_7654);
nor U8054 (N_8054,N_7655,N_7827);
or U8055 (N_8055,N_7692,N_7942);
or U8056 (N_8056,N_7748,N_7868);
nand U8057 (N_8057,N_7664,N_7830);
and U8058 (N_8058,N_7872,N_7861);
xor U8059 (N_8059,N_7638,N_7757);
and U8060 (N_8060,N_7671,N_7773);
and U8061 (N_8061,N_7612,N_7640);
nor U8062 (N_8062,N_7911,N_7627);
and U8063 (N_8063,N_7822,N_7633);
xor U8064 (N_8064,N_7608,N_7618);
nor U8065 (N_8065,N_7705,N_7854);
or U8066 (N_8066,N_7834,N_7927);
xor U8067 (N_8067,N_7787,N_7866);
xnor U8068 (N_8068,N_7919,N_7644);
xnor U8069 (N_8069,N_7605,N_7776);
xor U8070 (N_8070,N_7739,N_7657);
nor U8071 (N_8071,N_7950,N_7993);
or U8072 (N_8072,N_7697,N_7703);
nor U8073 (N_8073,N_7682,N_7634);
and U8074 (N_8074,N_7965,N_7616);
or U8075 (N_8075,N_7819,N_7975);
nor U8076 (N_8076,N_7838,N_7632);
nor U8077 (N_8077,N_7677,N_7818);
nor U8078 (N_8078,N_7716,N_7669);
and U8079 (N_8079,N_7845,N_7791);
or U8080 (N_8080,N_7877,N_7829);
nand U8081 (N_8081,N_7805,N_7969);
nand U8082 (N_8082,N_7662,N_7712);
nor U8083 (N_8083,N_7864,N_7940);
and U8084 (N_8084,N_7782,N_7629);
and U8085 (N_8085,N_7630,N_7978);
xor U8086 (N_8086,N_7923,N_7899);
or U8087 (N_8087,N_7994,N_7815);
and U8088 (N_8088,N_7752,N_7847);
nor U8089 (N_8089,N_7761,N_7972);
or U8090 (N_8090,N_7882,N_7698);
and U8091 (N_8091,N_7933,N_7893);
nor U8092 (N_8092,N_7951,N_7663);
nor U8093 (N_8093,N_7821,N_7701);
nor U8094 (N_8094,N_7863,N_7992);
or U8095 (N_8095,N_7767,N_7850);
nor U8096 (N_8096,N_7785,N_7720);
nor U8097 (N_8097,N_7848,N_7751);
or U8098 (N_8098,N_7892,N_7816);
nand U8099 (N_8099,N_7656,N_7836);
and U8100 (N_8100,N_7959,N_7916);
and U8101 (N_8101,N_7706,N_7930);
xor U8102 (N_8102,N_7700,N_7810);
and U8103 (N_8103,N_7981,N_7807);
nor U8104 (N_8104,N_7755,N_7774);
nor U8105 (N_8105,N_7835,N_7826);
nand U8106 (N_8106,N_7760,N_7727);
and U8107 (N_8107,N_7708,N_7606);
and U8108 (N_8108,N_7880,N_7685);
nand U8109 (N_8109,N_7853,N_7622);
nand U8110 (N_8110,N_7832,N_7624);
nor U8111 (N_8111,N_7777,N_7948);
nand U8112 (N_8112,N_7999,N_7673);
nor U8113 (N_8113,N_7990,N_7983);
and U8114 (N_8114,N_7695,N_7693);
and U8115 (N_8115,N_7909,N_7623);
nand U8116 (N_8116,N_7799,N_7688);
nor U8117 (N_8117,N_7957,N_7721);
or U8118 (N_8118,N_7658,N_7798);
and U8119 (N_8119,N_7670,N_7665);
or U8120 (N_8120,N_7886,N_7625);
or U8121 (N_8121,N_7897,N_7795);
xor U8122 (N_8122,N_7977,N_7747);
and U8123 (N_8123,N_7750,N_7917);
nand U8124 (N_8124,N_7793,N_7684);
nor U8125 (N_8125,N_7762,N_7823);
nor U8126 (N_8126,N_7915,N_7681);
and U8127 (N_8127,N_7934,N_7653);
xnor U8128 (N_8128,N_7869,N_7996);
xor U8129 (N_8129,N_7758,N_7711);
nand U8130 (N_8130,N_7997,N_7814);
nor U8131 (N_8131,N_7874,N_7926);
and U8132 (N_8132,N_7768,N_7987);
nor U8133 (N_8133,N_7600,N_7907);
xnor U8134 (N_8134,N_7737,N_7840);
or U8135 (N_8135,N_7719,N_7763);
and U8136 (N_8136,N_7648,N_7667);
and U8137 (N_8137,N_7906,N_7833);
nor U8138 (N_8138,N_7856,N_7858);
nand U8139 (N_8139,N_7742,N_7797);
xnor U8140 (N_8140,N_7675,N_7772);
xor U8141 (N_8141,N_7646,N_7745);
nand U8142 (N_8142,N_7784,N_7991);
nor U8143 (N_8143,N_7775,N_7846);
and U8144 (N_8144,N_7736,N_7986);
nor U8145 (N_8145,N_7715,N_7921);
xor U8146 (N_8146,N_7734,N_7649);
nand U8147 (N_8147,N_7824,N_7871);
and U8148 (N_8148,N_7626,N_7939);
and U8149 (N_8149,N_7873,N_7704);
and U8150 (N_8150,N_7998,N_7650);
nand U8151 (N_8151,N_7843,N_7603);
nand U8152 (N_8152,N_7931,N_7674);
xor U8153 (N_8153,N_7837,N_7765);
nor U8154 (N_8154,N_7960,N_7900);
nor U8155 (N_8155,N_7945,N_7672);
nor U8156 (N_8156,N_7889,N_7741);
or U8157 (N_8157,N_7613,N_7970);
nand U8158 (N_8158,N_7628,N_7988);
nor U8159 (N_8159,N_7642,N_7668);
or U8160 (N_8160,N_7888,N_7974);
and U8161 (N_8161,N_7733,N_7610);
and U8162 (N_8162,N_7867,N_7792);
or U8163 (N_8163,N_7935,N_7964);
or U8164 (N_8164,N_7601,N_7783);
xor U8165 (N_8165,N_7689,N_7680);
and U8166 (N_8166,N_7820,N_7753);
xnor U8167 (N_8167,N_7678,N_7967);
nor U8168 (N_8168,N_7690,N_7659);
nand U8169 (N_8169,N_7637,N_7729);
and U8170 (N_8170,N_7702,N_7683);
nand U8171 (N_8171,N_7743,N_7841);
nand U8172 (N_8172,N_7781,N_7817);
or U8173 (N_8173,N_7963,N_7661);
or U8174 (N_8174,N_7602,N_7619);
or U8175 (N_8175,N_7956,N_7879);
nand U8176 (N_8176,N_7828,N_7812);
nand U8177 (N_8177,N_7875,N_7980);
or U8178 (N_8178,N_7801,N_7796);
and U8179 (N_8179,N_7804,N_7769);
xor U8180 (N_8180,N_7699,N_7891);
xor U8181 (N_8181,N_7808,N_7849);
nor U8182 (N_8182,N_7901,N_7687);
or U8183 (N_8183,N_7883,N_7615);
xor U8184 (N_8184,N_7811,N_7878);
or U8185 (N_8185,N_7713,N_7803);
or U8186 (N_8186,N_7620,N_7925);
nand U8187 (N_8187,N_7724,N_7694);
nor U8188 (N_8188,N_7855,N_7639);
nand U8189 (N_8189,N_7651,N_7914);
and U8190 (N_8190,N_7961,N_7918);
nor U8191 (N_8191,N_7985,N_7928);
and U8192 (N_8192,N_7780,N_7895);
or U8193 (N_8193,N_7851,N_7884);
nor U8194 (N_8194,N_7722,N_7979);
xnor U8195 (N_8195,N_7738,N_7966);
and U8196 (N_8196,N_7844,N_7631);
xor U8197 (N_8197,N_7885,N_7726);
xnor U8198 (N_8198,N_7881,N_7778);
nand U8199 (N_8199,N_7976,N_7645);
and U8200 (N_8200,N_7656,N_7906);
and U8201 (N_8201,N_7822,N_7854);
or U8202 (N_8202,N_7709,N_7643);
or U8203 (N_8203,N_7837,N_7610);
or U8204 (N_8204,N_7978,N_7826);
or U8205 (N_8205,N_7671,N_7836);
and U8206 (N_8206,N_7780,N_7740);
nor U8207 (N_8207,N_7789,N_7699);
and U8208 (N_8208,N_7897,N_7900);
and U8209 (N_8209,N_7649,N_7985);
or U8210 (N_8210,N_7629,N_7977);
xor U8211 (N_8211,N_7984,N_7785);
and U8212 (N_8212,N_7699,N_7728);
or U8213 (N_8213,N_7827,N_7910);
and U8214 (N_8214,N_7964,N_7988);
nand U8215 (N_8215,N_7625,N_7742);
nand U8216 (N_8216,N_7693,N_7849);
nor U8217 (N_8217,N_7815,N_7892);
or U8218 (N_8218,N_7733,N_7741);
or U8219 (N_8219,N_7854,N_7987);
nor U8220 (N_8220,N_7628,N_7674);
or U8221 (N_8221,N_7942,N_7706);
and U8222 (N_8222,N_7967,N_7695);
nand U8223 (N_8223,N_7836,N_7711);
and U8224 (N_8224,N_7769,N_7900);
nor U8225 (N_8225,N_7850,N_7978);
or U8226 (N_8226,N_7683,N_7778);
xnor U8227 (N_8227,N_7853,N_7871);
nor U8228 (N_8228,N_7775,N_7740);
or U8229 (N_8229,N_7644,N_7727);
or U8230 (N_8230,N_7772,N_7819);
xnor U8231 (N_8231,N_7826,N_7700);
nor U8232 (N_8232,N_7764,N_7700);
and U8233 (N_8233,N_7843,N_7879);
nand U8234 (N_8234,N_7734,N_7932);
or U8235 (N_8235,N_7767,N_7636);
or U8236 (N_8236,N_7843,N_7887);
nor U8237 (N_8237,N_7637,N_7772);
nand U8238 (N_8238,N_7842,N_7638);
xnor U8239 (N_8239,N_7680,N_7783);
nor U8240 (N_8240,N_7996,N_7910);
or U8241 (N_8241,N_7713,N_7839);
nor U8242 (N_8242,N_7735,N_7738);
nor U8243 (N_8243,N_7653,N_7869);
nand U8244 (N_8244,N_7624,N_7690);
xnor U8245 (N_8245,N_7870,N_7986);
and U8246 (N_8246,N_7934,N_7860);
nor U8247 (N_8247,N_7778,N_7756);
xnor U8248 (N_8248,N_7995,N_7904);
nor U8249 (N_8249,N_7757,N_7736);
and U8250 (N_8250,N_7970,N_7645);
or U8251 (N_8251,N_7624,N_7969);
nand U8252 (N_8252,N_7986,N_7872);
nor U8253 (N_8253,N_7981,N_7681);
and U8254 (N_8254,N_7943,N_7763);
or U8255 (N_8255,N_7666,N_7868);
and U8256 (N_8256,N_7837,N_7668);
nor U8257 (N_8257,N_7955,N_7752);
nand U8258 (N_8258,N_7991,N_7647);
and U8259 (N_8259,N_7727,N_7722);
nor U8260 (N_8260,N_7961,N_7902);
nor U8261 (N_8261,N_7604,N_7855);
and U8262 (N_8262,N_7938,N_7768);
or U8263 (N_8263,N_7735,N_7932);
nor U8264 (N_8264,N_7970,N_7702);
nor U8265 (N_8265,N_7862,N_7914);
and U8266 (N_8266,N_7992,N_7983);
nand U8267 (N_8267,N_7649,N_7773);
xnor U8268 (N_8268,N_7968,N_7911);
or U8269 (N_8269,N_7817,N_7974);
nor U8270 (N_8270,N_7726,N_7681);
xor U8271 (N_8271,N_7839,N_7634);
or U8272 (N_8272,N_7771,N_7615);
xnor U8273 (N_8273,N_7631,N_7889);
nor U8274 (N_8274,N_7682,N_7759);
nand U8275 (N_8275,N_7836,N_7894);
or U8276 (N_8276,N_7723,N_7984);
and U8277 (N_8277,N_7911,N_7954);
and U8278 (N_8278,N_7918,N_7992);
nand U8279 (N_8279,N_7970,N_7979);
nand U8280 (N_8280,N_7718,N_7692);
nor U8281 (N_8281,N_7993,N_7622);
or U8282 (N_8282,N_7643,N_7685);
or U8283 (N_8283,N_7747,N_7691);
nor U8284 (N_8284,N_7782,N_7970);
nand U8285 (N_8285,N_7671,N_7976);
nand U8286 (N_8286,N_7831,N_7825);
nand U8287 (N_8287,N_7869,N_7894);
nand U8288 (N_8288,N_7669,N_7819);
nand U8289 (N_8289,N_7929,N_7756);
xnor U8290 (N_8290,N_7704,N_7670);
or U8291 (N_8291,N_7779,N_7684);
and U8292 (N_8292,N_7990,N_7619);
nand U8293 (N_8293,N_7925,N_7983);
nand U8294 (N_8294,N_7938,N_7869);
xor U8295 (N_8295,N_7867,N_7769);
nor U8296 (N_8296,N_7868,N_7957);
xnor U8297 (N_8297,N_7806,N_7800);
or U8298 (N_8298,N_7623,N_7732);
xor U8299 (N_8299,N_7747,N_7781);
and U8300 (N_8300,N_7703,N_7848);
or U8301 (N_8301,N_7698,N_7891);
nand U8302 (N_8302,N_7890,N_7624);
xor U8303 (N_8303,N_7601,N_7612);
and U8304 (N_8304,N_7734,N_7742);
or U8305 (N_8305,N_7923,N_7694);
or U8306 (N_8306,N_7745,N_7965);
nand U8307 (N_8307,N_7837,N_7921);
and U8308 (N_8308,N_7933,N_7791);
nand U8309 (N_8309,N_7712,N_7981);
nand U8310 (N_8310,N_7941,N_7713);
nand U8311 (N_8311,N_7808,N_7612);
nor U8312 (N_8312,N_7799,N_7765);
xor U8313 (N_8313,N_7772,N_7867);
or U8314 (N_8314,N_7965,N_7935);
or U8315 (N_8315,N_7771,N_7814);
or U8316 (N_8316,N_7930,N_7788);
and U8317 (N_8317,N_7943,N_7931);
nand U8318 (N_8318,N_7884,N_7883);
nor U8319 (N_8319,N_7688,N_7675);
nor U8320 (N_8320,N_7722,N_7808);
or U8321 (N_8321,N_7862,N_7653);
or U8322 (N_8322,N_7681,N_7801);
and U8323 (N_8323,N_7733,N_7952);
nor U8324 (N_8324,N_7727,N_7778);
xnor U8325 (N_8325,N_7883,N_7755);
nand U8326 (N_8326,N_7847,N_7967);
nor U8327 (N_8327,N_7748,N_7780);
and U8328 (N_8328,N_7724,N_7627);
xnor U8329 (N_8329,N_7976,N_7746);
xnor U8330 (N_8330,N_7753,N_7962);
nand U8331 (N_8331,N_7617,N_7755);
nand U8332 (N_8332,N_7666,N_7763);
xor U8333 (N_8333,N_7962,N_7689);
and U8334 (N_8334,N_7818,N_7838);
xnor U8335 (N_8335,N_7878,N_7774);
nor U8336 (N_8336,N_7870,N_7871);
nand U8337 (N_8337,N_7849,N_7697);
xor U8338 (N_8338,N_7888,N_7780);
and U8339 (N_8339,N_7877,N_7610);
and U8340 (N_8340,N_7882,N_7964);
nand U8341 (N_8341,N_7857,N_7608);
nor U8342 (N_8342,N_7667,N_7760);
nand U8343 (N_8343,N_7607,N_7621);
xnor U8344 (N_8344,N_7824,N_7787);
xnor U8345 (N_8345,N_7750,N_7857);
xnor U8346 (N_8346,N_7948,N_7696);
nor U8347 (N_8347,N_7939,N_7912);
or U8348 (N_8348,N_7926,N_7634);
nand U8349 (N_8349,N_7905,N_7909);
or U8350 (N_8350,N_7694,N_7827);
nand U8351 (N_8351,N_7772,N_7750);
nand U8352 (N_8352,N_7705,N_7971);
nand U8353 (N_8353,N_7985,N_7881);
nand U8354 (N_8354,N_7905,N_7748);
or U8355 (N_8355,N_7905,N_7670);
nor U8356 (N_8356,N_7925,N_7997);
and U8357 (N_8357,N_7936,N_7759);
and U8358 (N_8358,N_7925,N_7602);
xnor U8359 (N_8359,N_7952,N_7683);
nand U8360 (N_8360,N_7916,N_7913);
nand U8361 (N_8361,N_7670,N_7696);
nand U8362 (N_8362,N_7620,N_7704);
nor U8363 (N_8363,N_7821,N_7771);
and U8364 (N_8364,N_7765,N_7728);
or U8365 (N_8365,N_7919,N_7869);
nand U8366 (N_8366,N_7728,N_7965);
nand U8367 (N_8367,N_7995,N_7929);
nand U8368 (N_8368,N_7784,N_7979);
xnor U8369 (N_8369,N_7827,N_7664);
and U8370 (N_8370,N_7622,N_7692);
or U8371 (N_8371,N_7752,N_7788);
or U8372 (N_8372,N_7649,N_7666);
nand U8373 (N_8373,N_7964,N_7867);
nand U8374 (N_8374,N_7870,N_7975);
or U8375 (N_8375,N_7958,N_7814);
or U8376 (N_8376,N_7633,N_7614);
nor U8377 (N_8377,N_7882,N_7621);
nand U8378 (N_8378,N_7784,N_7849);
and U8379 (N_8379,N_7727,N_7844);
and U8380 (N_8380,N_7953,N_7751);
xor U8381 (N_8381,N_7845,N_7725);
and U8382 (N_8382,N_7806,N_7772);
and U8383 (N_8383,N_7663,N_7824);
and U8384 (N_8384,N_7765,N_7747);
xor U8385 (N_8385,N_7670,N_7657);
or U8386 (N_8386,N_7765,N_7767);
nand U8387 (N_8387,N_7634,N_7981);
nand U8388 (N_8388,N_7783,N_7642);
nor U8389 (N_8389,N_7780,N_7622);
or U8390 (N_8390,N_7651,N_7968);
xor U8391 (N_8391,N_7692,N_7868);
nand U8392 (N_8392,N_7919,N_7667);
and U8393 (N_8393,N_7671,N_7932);
xor U8394 (N_8394,N_7910,N_7848);
or U8395 (N_8395,N_7815,N_7810);
nor U8396 (N_8396,N_7653,N_7897);
xnor U8397 (N_8397,N_7864,N_7635);
nor U8398 (N_8398,N_7897,N_7690);
and U8399 (N_8399,N_7788,N_7837);
nand U8400 (N_8400,N_8167,N_8141);
xor U8401 (N_8401,N_8058,N_8086);
nor U8402 (N_8402,N_8063,N_8396);
nand U8403 (N_8403,N_8270,N_8202);
xnor U8404 (N_8404,N_8189,N_8066);
or U8405 (N_8405,N_8161,N_8077);
nand U8406 (N_8406,N_8187,N_8144);
and U8407 (N_8407,N_8069,N_8256);
and U8408 (N_8408,N_8268,N_8055);
nand U8409 (N_8409,N_8290,N_8262);
xor U8410 (N_8410,N_8044,N_8240);
and U8411 (N_8411,N_8029,N_8281);
or U8412 (N_8412,N_8383,N_8070);
xnor U8413 (N_8413,N_8180,N_8230);
and U8414 (N_8414,N_8001,N_8027);
or U8415 (N_8415,N_8079,N_8047);
nor U8416 (N_8416,N_8274,N_8165);
nand U8417 (N_8417,N_8163,N_8030);
or U8418 (N_8418,N_8105,N_8379);
nor U8419 (N_8419,N_8038,N_8152);
xor U8420 (N_8420,N_8217,N_8172);
xnor U8421 (N_8421,N_8157,N_8036);
and U8422 (N_8422,N_8394,N_8385);
and U8423 (N_8423,N_8326,N_8068);
and U8424 (N_8424,N_8158,N_8249);
and U8425 (N_8425,N_8022,N_8175);
and U8426 (N_8426,N_8159,N_8129);
xor U8427 (N_8427,N_8072,N_8366);
nand U8428 (N_8428,N_8247,N_8201);
xnor U8429 (N_8429,N_8088,N_8284);
nand U8430 (N_8430,N_8288,N_8314);
or U8431 (N_8431,N_8050,N_8118);
nor U8432 (N_8432,N_8294,N_8322);
xor U8433 (N_8433,N_8233,N_8358);
xor U8434 (N_8434,N_8226,N_8090);
nand U8435 (N_8435,N_8215,N_8133);
and U8436 (N_8436,N_8252,N_8039);
or U8437 (N_8437,N_8271,N_8287);
nand U8438 (N_8438,N_8190,N_8193);
and U8439 (N_8439,N_8232,N_8355);
and U8440 (N_8440,N_8034,N_8128);
nor U8441 (N_8441,N_8289,N_8346);
nor U8442 (N_8442,N_8208,N_8220);
xnor U8443 (N_8443,N_8302,N_8388);
nand U8444 (N_8444,N_8299,N_8026);
nand U8445 (N_8445,N_8285,N_8196);
xor U8446 (N_8446,N_8258,N_8378);
and U8447 (N_8447,N_8339,N_8253);
nor U8448 (N_8448,N_8259,N_8041);
xnor U8449 (N_8449,N_8124,N_8060);
xnor U8450 (N_8450,N_8049,N_8057);
xor U8451 (N_8451,N_8316,N_8371);
nand U8452 (N_8452,N_8370,N_8365);
nand U8453 (N_8453,N_8145,N_8183);
nand U8454 (N_8454,N_8359,N_8037);
nor U8455 (N_8455,N_8243,N_8176);
nor U8456 (N_8456,N_8238,N_8012);
xnor U8457 (N_8457,N_8195,N_8239);
nand U8458 (N_8458,N_8059,N_8228);
and U8459 (N_8459,N_8021,N_8260);
and U8460 (N_8460,N_8218,N_8344);
and U8461 (N_8461,N_8368,N_8219);
and U8462 (N_8462,N_8315,N_8397);
nand U8463 (N_8463,N_8122,N_8130);
or U8464 (N_8464,N_8225,N_8235);
nand U8465 (N_8465,N_8301,N_8361);
nor U8466 (N_8466,N_8283,N_8182);
xnor U8467 (N_8467,N_8064,N_8376);
and U8468 (N_8468,N_8179,N_8393);
xor U8469 (N_8469,N_8310,N_8053);
xnor U8470 (N_8470,N_8280,N_8317);
nand U8471 (N_8471,N_8108,N_8292);
nand U8472 (N_8472,N_8237,N_8076);
xor U8473 (N_8473,N_8153,N_8333);
or U8474 (N_8474,N_8051,N_8251);
xor U8475 (N_8475,N_8277,N_8092);
nor U8476 (N_8476,N_8296,N_8033);
and U8477 (N_8477,N_8348,N_8123);
nor U8478 (N_8478,N_8173,N_8156);
nor U8479 (N_8479,N_8148,N_8095);
nand U8480 (N_8480,N_8342,N_8354);
xnor U8481 (N_8481,N_8046,N_8200);
or U8482 (N_8482,N_8045,N_8330);
and U8483 (N_8483,N_8003,N_8194);
nor U8484 (N_8484,N_8276,N_8389);
nand U8485 (N_8485,N_8328,N_8116);
nand U8486 (N_8486,N_8007,N_8131);
or U8487 (N_8487,N_8162,N_8140);
or U8488 (N_8488,N_8099,N_8155);
and U8489 (N_8489,N_8340,N_8320);
nor U8490 (N_8490,N_8255,N_8094);
or U8491 (N_8491,N_8335,N_8000);
and U8492 (N_8492,N_8171,N_8040);
nand U8493 (N_8493,N_8343,N_8221);
and U8494 (N_8494,N_8132,N_8298);
nand U8495 (N_8495,N_8244,N_8367);
nand U8496 (N_8496,N_8127,N_8091);
nor U8497 (N_8497,N_8282,N_8236);
nand U8498 (N_8498,N_8224,N_8143);
nor U8499 (N_8499,N_8360,N_8111);
nand U8500 (N_8500,N_8363,N_8178);
and U8501 (N_8501,N_8013,N_8192);
xor U8502 (N_8502,N_8211,N_8386);
xnor U8503 (N_8503,N_8151,N_8364);
and U8504 (N_8504,N_8186,N_8010);
or U8505 (N_8505,N_8074,N_8149);
and U8506 (N_8506,N_8185,N_8168);
and U8507 (N_8507,N_8032,N_8214);
and U8508 (N_8508,N_8392,N_8031);
xor U8509 (N_8509,N_8234,N_8071);
nor U8510 (N_8510,N_8206,N_8223);
and U8511 (N_8511,N_8293,N_8341);
and U8512 (N_8512,N_8222,N_8126);
nand U8513 (N_8513,N_8350,N_8164);
xnor U8514 (N_8514,N_8197,N_8306);
nand U8515 (N_8515,N_8107,N_8177);
nor U8516 (N_8516,N_8267,N_8075);
and U8517 (N_8517,N_8054,N_8275);
nand U8518 (N_8518,N_8269,N_8257);
xnor U8519 (N_8519,N_8097,N_8254);
nor U8520 (N_8520,N_8345,N_8005);
nor U8521 (N_8521,N_8093,N_8203);
and U8522 (N_8522,N_8205,N_8369);
xnor U8523 (N_8523,N_8014,N_8242);
nor U8524 (N_8524,N_8198,N_8078);
nand U8525 (N_8525,N_8381,N_8263);
xnor U8526 (N_8526,N_8147,N_8150);
nand U8527 (N_8527,N_8025,N_8102);
xor U8528 (N_8528,N_8043,N_8020);
xor U8529 (N_8529,N_8017,N_8035);
nand U8530 (N_8530,N_8391,N_8272);
xor U8531 (N_8531,N_8023,N_8347);
or U8532 (N_8532,N_8120,N_8184);
or U8533 (N_8533,N_8297,N_8137);
or U8534 (N_8534,N_8212,N_8134);
nor U8535 (N_8535,N_8336,N_8015);
xnor U8536 (N_8536,N_8216,N_8323);
nand U8537 (N_8537,N_8080,N_8313);
or U8538 (N_8538,N_8207,N_8109);
nand U8539 (N_8539,N_8204,N_8384);
or U8540 (N_8540,N_8209,N_8387);
xor U8541 (N_8541,N_8169,N_8114);
nor U8542 (N_8542,N_8113,N_8304);
nand U8543 (N_8543,N_8227,N_8117);
nand U8544 (N_8544,N_8191,N_8112);
nand U8545 (N_8545,N_8087,N_8353);
nor U8546 (N_8546,N_8352,N_8338);
nor U8547 (N_8547,N_8098,N_8011);
nand U8548 (N_8548,N_8291,N_8002);
and U8549 (N_8549,N_8100,N_8009);
nand U8550 (N_8550,N_8018,N_8265);
nand U8551 (N_8551,N_8006,N_8067);
nor U8552 (N_8552,N_8199,N_8308);
nand U8553 (N_8553,N_8082,N_8125);
or U8554 (N_8554,N_8300,N_8154);
nand U8555 (N_8555,N_8321,N_8318);
or U8556 (N_8556,N_8229,N_8286);
nand U8557 (N_8557,N_8052,N_8062);
nor U8558 (N_8558,N_8377,N_8081);
and U8559 (N_8559,N_8231,N_8349);
nand U8560 (N_8560,N_8398,N_8374);
or U8561 (N_8561,N_8261,N_8372);
or U8562 (N_8562,N_8115,N_8136);
nand U8563 (N_8563,N_8278,N_8264);
or U8564 (N_8564,N_8016,N_8273);
and U8565 (N_8565,N_8142,N_8028);
xor U8566 (N_8566,N_8135,N_8170);
xor U8567 (N_8567,N_8337,N_8073);
and U8568 (N_8568,N_8083,N_8279);
or U8569 (N_8569,N_8241,N_8309);
nand U8570 (N_8570,N_8210,N_8061);
nor U8571 (N_8571,N_8375,N_8246);
nor U8572 (N_8572,N_8019,N_8042);
nor U8573 (N_8573,N_8362,N_8103);
nand U8574 (N_8574,N_8104,N_8213);
nor U8575 (N_8575,N_8084,N_8351);
nand U8576 (N_8576,N_8248,N_8312);
nand U8577 (N_8577,N_8146,N_8089);
or U8578 (N_8578,N_8139,N_8266);
nor U8579 (N_8579,N_8324,N_8008);
nor U8580 (N_8580,N_8110,N_8096);
or U8581 (N_8581,N_8356,N_8399);
nand U8582 (N_8582,N_8303,N_8395);
nor U8583 (N_8583,N_8181,N_8332);
or U8584 (N_8584,N_8160,N_8024);
and U8585 (N_8585,N_8380,N_8250);
and U8586 (N_8586,N_8382,N_8101);
nand U8587 (N_8587,N_8319,N_8311);
and U8588 (N_8588,N_8188,N_8106);
nor U8589 (N_8589,N_8331,N_8295);
nand U8590 (N_8590,N_8334,N_8119);
and U8591 (N_8591,N_8373,N_8329);
and U8592 (N_8592,N_8048,N_8056);
nor U8593 (N_8593,N_8307,N_8085);
or U8594 (N_8594,N_8245,N_8325);
nor U8595 (N_8595,N_8065,N_8357);
xor U8596 (N_8596,N_8004,N_8305);
xor U8597 (N_8597,N_8138,N_8390);
and U8598 (N_8598,N_8121,N_8174);
nor U8599 (N_8599,N_8166,N_8327);
nand U8600 (N_8600,N_8302,N_8165);
xnor U8601 (N_8601,N_8243,N_8041);
or U8602 (N_8602,N_8143,N_8034);
and U8603 (N_8603,N_8367,N_8038);
xor U8604 (N_8604,N_8283,N_8006);
nor U8605 (N_8605,N_8321,N_8024);
nand U8606 (N_8606,N_8383,N_8382);
nand U8607 (N_8607,N_8238,N_8009);
nand U8608 (N_8608,N_8194,N_8374);
or U8609 (N_8609,N_8333,N_8171);
nor U8610 (N_8610,N_8177,N_8053);
and U8611 (N_8611,N_8180,N_8338);
nor U8612 (N_8612,N_8071,N_8376);
xnor U8613 (N_8613,N_8247,N_8305);
xnor U8614 (N_8614,N_8375,N_8204);
or U8615 (N_8615,N_8363,N_8081);
nor U8616 (N_8616,N_8337,N_8155);
or U8617 (N_8617,N_8300,N_8256);
or U8618 (N_8618,N_8338,N_8193);
or U8619 (N_8619,N_8253,N_8246);
xnor U8620 (N_8620,N_8020,N_8164);
nor U8621 (N_8621,N_8331,N_8374);
and U8622 (N_8622,N_8105,N_8371);
or U8623 (N_8623,N_8079,N_8262);
and U8624 (N_8624,N_8381,N_8154);
or U8625 (N_8625,N_8042,N_8326);
and U8626 (N_8626,N_8140,N_8121);
nor U8627 (N_8627,N_8161,N_8261);
xor U8628 (N_8628,N_8032,N_8010);
xor U8629 (N_8629,N_8131,N_8072);
nand U8630 (N_8630,N_8212,N_8295);
nand U8631 (N_8631,N_8134,N_8094);
and U8632 (N_8632,N_8216,N_8391);
nand U8633 (N_8633,N_8066,N_8218);
or U8634 (N_8634,N_8067,N_8245);
xor U8635 (N_8635,N_8386,N_8255);
xnor U8636 (N_8636,N_8110,N_8040);
nor U8637 (N_8637,N_8049,N_8069);
nor U8638 (N_8638,N_8256,N_8210);
xor U8639 (N_8639,N_8314,N_8251);
nor U8640 (N_8640,N_8219,N_8034);
xor U8641 (N_8641,N_8037,N_8067);
or U8642 (N_8642,N_8277,N_8322);
xor U8643 (N_8643,N_8243,N_8333);
and U8644 (N_8644,N_8210,N_8216);
nor U8645 (N_8645,N_8070,N_8384);
nor U8646 (N_8646,N_8197,N_8192);
and U8647 (N_8647,N_8243,N_8093);
nor U8648 (N_8648,N_8106,N_8273);
xor U8649 (N_8649,N_8037,N_8042);
nor U8650 (N_8650,N_8315,N_8104);
xor U8651 (N_8651,N_8192,N_8120);
nand U8652 (N_8652,N_8087,N_8060);
nor U8653 (N_8653,N_8050,N_8098);
and U8654 (N_8654,N_8095,N_8289);
xnor U8655 (N_8655,N_8336,N_8163);
and U8656 (N_8656,N_8238,N_8350);
nand U8657 (N_8657,N_8223,N_8264);
nand U8658 (N_8658,N_8082,N_8120);
and U8659 (N_8659,N_8205,N_8291);
or U8660 (N_8660,N_8076,N_8268);
and U8661 (N_8661,N_8135,N_8106);
xor U8662 (N_8662,N_8314,N_8395);
xor U8663 (N_8663,N_8092,N_8365);
nand U8664 (N_8664,N_8227,N_8286);
xor U8665 (N_8665,N_8023,N_8095);
nor U8666 (N_8666,N_8310,N_8355);
nand U8667 (N_8667,N_8279,N_8121);
xor U8668 (N_8668,N_8205,N_8313);
nor U8669 (N_8669,N_8024,N_8264);
or U8670 (N_8670,N_8327,N_8239);
and U8671 (N_8671,N_8057,N_8228);
or U8672 (N_8672,N_8300,N_8218);
nor U8673 (N_8673,N_8100,N_8362);
nand U8674 (N_8674,N_8125,N_8009);
nand U8675 (N_8675,N_8390,N_8113);
and U8676 (N_8676,N_8275,N_8347);
and U8677 (N_8677,N_8235,N_8035);
nand U8678 (N_8678,N_8385,N_8204);
or U8679 (N_8679,N_8086,N_8343);
and U8680 (N_8680,N_8092,N_8187);
nand U8681 (N_8681,N_8351,N_8244);
xnor U8682 (N_8682,N_8134,N_8244);
nand U8683 (N_8683,N_8162,N_8245);
or U8684 (N_8684,N_8395,N_8145);
nor U8685 (N_8685,N_8030,N_8338);
xnor U8686 (N_8686,N_8221,N_8341);
nand U8687 (N_8687,N_8188,N_8161);
or U8688 (N_8688,N_8007,N_8348);
and U8689 (N_8689,N_8347,N_8147);
nand U8690 (N_8690,N_8302,N_8155);
nand U8691 (N_8691,N_8240,N_8293);
or U8692 (N_8692,N_8374,N_8205);
nand U8693 (N_8693,N_8055,N_8144);
xor U8694 (N_8694,N_8031,N_8255);
nand U8695 (N_8695,N_8014,N_8023);
nor U8696 (N_8696,N_8157,N_8274);
nand U8697 (N_8697,N_8321,N_8111);
or U8698 (N_8698,N_8279,N_8338);
nand U8699 (N_8699,N_8326,N_8024);
nand U8700 (N_8700,N_8212,N_8261);
nand U8701 (N_8701,N_8262,N_8387);
nand U8702 (N_8702,N_8355,N_8371);
nand U8703 (N_8703,N_8381,N_8229);
nor U8704 (N_8704,N_8186,N_8119);
nor U8705 (N_8705,N_8263,N_8338);
and U8706 (N_8706,N_8188,N_8191);
nand U8707 (N_8707,N_8221,N_8007);
nand U8708 (N_8708,N_8216,N_8142);
or U8709 (N_8709,N_8067,N_8066);
nand U8710 (N_8710,N_8361,N_8009);
nand U8711 (N_8711,N_8327,N_8195);
nor U8712 (N_8712,N_8341,N_8357);
or U8713 (N_8713,N_8312,N_8372);
or U8714 (N_8714,N_8208,N_8240);
xor U8715 (N_8715,N_8306,N_8136);
xnor U8716 (N_8716,N_8070,N_8161);
xor U8717 (N_8717,N_8213,N_8360);
or U8718 (N_8718,N_8381,N_8291);
xnor U8719 (N_8719,N_8333,N_8113);
and U8720 (N_8720,N_8049,N_8011);
nand U8721 (N_8721,N_8368,N_8256);
nand U8722 (N_8722,N_8073,N_8289);
nor U8723 (N_8723,N_8385,N_8143);
nand U8724 (N_8724,N_8168,N_8175);
and U8725 (N_8725,N_8121,N_8006);
and U8726 (N_8726,N_8147,N_8124);
xnor U8727 (N_8727,N_8262,N_8126);
or U8728 (N_8728,N_8266,N_8027);
or U8729 (N_8729,N_8063,N_8083);
nor U8730 (N_8730,N_8090,N_8068);
nor U8731 (N_8731,N_8082,N_8284);
and U8732 (N_8732,N_8193,N_8148);
or U8733 (N_8733,N_8371,N_8315);
nor U8734 (N_8734,N_8065,N_8275);
and U8735 (N_8735,N_8027,N_8253);
nand U8736 (N_8736,N_8215,N_8395);
and U8737 (N_8737,N_8032,N_8107);
nor U8738 (N_8738,N_8283,N_8335);
xor U8739 (N_8739,N_8028,N_8229);
nand U8740 (N_8740,N_8045,N_8073);
and U8741 (N_8741,N_8244,N_8081);
or U8742 (N_8742,N_8039,N_8352);
and U8743 (N_8743,N_8205,N_8140);
or U8744 (N_8744,N_8210,N_8303);
nor U8745 (N_8745,N_8079,N_8349);
or U8746 (N_8746,N_8139,N_8242);
or U8747 (N_8747,N_8309,N_8143);
nor U8748 (N_8748,N_8340,N_8107);
xor U8749 (N_8749,N_8056,N_8341);
nor U8750 (N_8750,N_8118,N_8026);
nand U8751 (N_8751,N_8002,N_8313);
xnor U8752 (N_8752,N_8157,N_8111);
and U8753 (N_8753,N_8061,N_8108);
xor U8754 (N_8754,N_8265,N_8155);
nor U8755 (N_8755,N_8233,N_8253);
or U8756 (N_8756,N_8095,N_8158);
nor U8757 (N_8757,N_8186,N_8120);
or U8758 (N_8758,N_8185,N_8214);
nor U8759 (N_8759,N_8048,N_8347);
nand U8760 (N_8760,N_8317,N_8066);
nor U8761 (N_8761,N_8254,N_8282);
xor U8762 (N_8762,N_8179,N_8113);
nor U8763 (N_8763,N_8176,N_8156);
nor U8764 (N_8764,N_8272,N_8207);
and U8765 (N_8765,N_8074,N_8301);
nor U8766 (N_8766,N_8252,N_8228);
xor U8767 (N_8767,N_8338,N_8371);
xor U8768 (N_8768,N_8131,N_8146);
or U8769 (N_8769,N_8254,N_8339);
nand U8770 (N_8770,N_8078,N_8089);
or U8771 (N_8771,N_8354,N_8321);
nand U8772 (N_8772,N_8135,N_8281);
nor U8773 (N_8773,N_8189,N_8258);
and U8774 (N_8774,N_8173,N_8311);
and U8775 (N_8775,N_8289,N_8328);
and U8776 (N_8776,N_8305,N_8024);
nand U8777 (N_8777,N_8236,N_8016);
nor U8778 (N_8778,N_8152,N_8299);
xnor U8779 (N_8779,N_8196,N_8056);
nor U8780 (N_8780,N_8249,N_8198);
nand U8781 (N_8781,N_8282,N_8206);
nand U8782 (N_8782,N_8174,N_8380);
and U8783 (N_8783,N_8268,N_8299);
nand U8784 (N_8784,N_8119,N_8298);
nor U8785 (N_8785,N_8106,N_8105);
nand U8786 (N_8786,N_8393,N_8329);
and U8787 (N_8787,N_8064,N_8257);
nor U8788 (N_8788,N_8349,N_8243);
nor U8789 (N_8789,N_8140,N_8075);
xor U8790 (N_8790,N_8196,N_8163);
xor U8791 (N_8791,N_8300,N_8158);
xnor U8792 (N_8792,N_8015,N_8122);
and U8793 (N_8793,N_8220,N_8165);
xor U8794 (N_8794,N_8235,N_8017);
nand U8795 (N_8795,N_8272,N_8049);
and U8796 (N_8796,N_8347,N_8128);
xor U8797 (N_8797,N_8123,N_8086);
nand U8798 (N_8798,N_8389,N_8375);
xnor U8799 (N_8799,N_8394,N_8308);
xnor U8800 (N_8800,N_8569,N_8785);
nor U8801 (N_8801,N_8603,N_8768);
xnor U8802 (N_8802,N_8675,N_8550);
nor U8803 (N_8803,N_8470,N_8698);
nor U8804 (N_8804,N_8437,N_8485);
nor U8805 (N_8805,N_8405,N_8460);
nand U8806 (N_8806,N_8631,N_8677);
nand U8807 (N_8807,N_8628,N_8772);
nand U8808 (N_8808,N_8536,N_8749);
nand U8809 (N_8809,N_8425,N_8672);
and U8810 (N_8810,N_8649,N_8546);
nor U8811 (N_8811,N_8403,N_8618);
nand U8812 (N_8812,N_8673,N_8765);
xnor U8813 (N_8813,N_8617,N_8430);
or U8814 (N_8814,N_8761,N_8688);
xor U8815 (N_8815,N_8750,N_8453);
xnor U8816 (N_8816,N_8442,N_8757);
xnor U8817 (N_8817,N_8520,N_8682);
nor U8818 (N_8818,N_8481,N_8690);
nor U8819 (N_8819,N_8473,N_8566);
nand U8820 (N_8820,N_8633,N_8693);
nand U8821 (N_8821,N_8674,N_8576);
or U8822 (N_8822,N_8584,N_8630);
or U8823 (N_8823,N_8668,N_8592);
nor U8824 (N_8824,N_8515,N_8614);
and U8825 (N_8825,N_8454,N_8663);
and U8826 (N_8826,N_8594,N_8639);
or U8827 (N_8827,N_8486,N_8711);
and U8828 (N_8828,N_8725,N_8604);
nor U8829 (N_8829,N_8789,N_8570);
and U8830 (N_8830,N_8792,N_8527);
xnor U8831 (N_8831,N_8737,N_8606);
nand U8832 (N_8832,N_8538,N_8544);
nand U8833 (N_8833,N_8552,N_8565);
nor U8834 (N_8834,N_8703,N_8714);
nor U8835 (N_8835,N_8678,N_8531);
and U8836 (N_8836,N_8601,N_8529);
and U8837 (N_8837,N_8502,N_8627);
xor U8838 (N_8838,N_8581,N_8448);
nand U8839 (N_8839,N_8426,N_8595);
or U8840 (N_8840,N_8503,N_8653);
nor U8841 (N_8841,N_8452,N_8559);
and U8842 (N_8842,N_8717,N_8652);
xor U8843 (N_8843,N_8716,N_8778);
and U8844 (N_8844,N_8608,N_8651);
nor U8845 (N_8845,N_8758,N_8622);
nand U8846 (N_8846,N_8548,N_8457);
xnor U8847 (N_8847,N_8766,N_8522);
and U8848 (N_8848,N_8476,N_8401);
xnor U8849 (N_8849,N_8477,N_8610);
nand U8850 (N_8850,N_8773,N_8459);
nor U8851 (N_8851,N_8720,N_8721);
nor U8852 (N_8852,N_8433,N_8466);
nand U8853 (N_8853,N_8530,N_8635);
nand U8854 (N_8854,N_8474,N_8769);
nand U8855 (N_8855,N_8469,N_8794);
and U8856 (N_8856,N_8472,N_8694);
nor U8857 (N_8857,N_8767,N_8461);
and U8858 (N_8858,N_8752,N_8499);
and U8859 (N_8859,N_8587,N_8620);
and U8860 (N_8860,N_8407,N_8704);
nand U8861 (N_8861,N_8458,N_8751);
nand U8862 (N_8862,N_8419,N_8662);
xnor U8863 (N_8863,N_8744,N_8621);
and U8864 (N_8864,N_8555,N_8701);
or U8865 (N_8865,N_8414,N_8739);
and U8866 (N_8866,N_8488,N_8416);
xor U8867 (N_8867,N_8432,N_8764);
nand U8868 (N_8868,N_8611,N_8541);
nand U8869 (N_8869,N_8615,N_8423);
and U8870 (N_8870,N_8676,N_8483);
or U8871 (N_8871,N_8753,N_8738);
nand U8872 (N_8872,N_8523,N_8556);
or U8873 (N_8873,N_8686,N_8699);
or U8874 (N_8874,N_8647,N_8504);
or U8875 (N_8875,N_8718,N_8511);
and U8876 (N_8876,N_8726,N_8429);
and U8877 (N_8877,N_8687,N_8787);
xor U8878 (N_8878,N_8642,N_8696);
and U8879 (N_8879,N_8444,N_8786);
and U8880 (N_8880,N_8634,N_8733);
nor U8881 (N_8881,N_8435,N_8625);
nor U8882 (N_8882,N_8605,N_8549);
nor U8883 (N_8883,N_8497,N_8700);
and U8884 (N_8884,N_8648,N_8557);
or U8885 (N_8885,N_8567,N_8406);
nand U8886 (N_8886,N_8748,N_8783);
nand U8887 (N_8887,N_8456,N_8415);
and U8888 (N_8888,N_8585,N_8422);
and U8889 (N_8889,N_8440,N_8526);
nand U8890 (N_8890,N_8417,N_8708);
nand U8891 (N_8891,N_8543,N_8712);
xor U8892 (N_8892,N_8754,N_8586);
or U8893 (N_8893,N_8702,N_8600);
nor U8894 (N_8894,N_8508,N_8547);
and U8895 (N_8895,N_8759,N_8501);
and U8896 (N_8896,N_8695,N_8684);
or U8897 (N_8897,N_8577,N_8528);
and U8898 (N_8898,N_8667,N_8658);
or U8899 (N_8899,N_8514,N_8609);
and U8900 (N_8900,N_8740,N_8496);
xnor U8901 (N_8901,N_8760,N_8478);
nor U8902 (N_8902,N_8644,N_8660);
nand U8903 (N_8903,N_8728,N_8413);
nor U8904 (N_8904,N_8624,N_8747);
or U8905 (N_8905,N_8500,N_8495);
xor U8906 (N_8906,N_8692,N_8774);
nand U8907 (N_8907,N_8591,N_8561);
nor U8908 (N_8908,N_8468,N_8475);
xor U8909 (N_8909,N_8575,N_8731);
xnor U8910 (N_8910,N_8664,N_8408);
or U8911 (N_8911,N_8705,N_8613);
nand U8912 (N_8912,N_8713,N_8580);
nor U8913 (N_8913,N_8681,N_8428);
nor U8914 (N_8914,N_8404,N_8629);
or U8915 (N_8915,N_8697,N_8619);
and U8916 (N_8916,N_8492,N_8411);
nor U8917 (N_8917,N_8519,N_8489);
and U8918 (N_8918,N_8562,N_8539);
or U8919 (N_8919,N_8599,N_8517);
nor U8920 (N_8920,N_8588,N_8509);
and U8921 (N_8921,N_8724,N_8507);
and U8922 (N_8922,N_8480,N_8579);
nor U8923 (N_8923,N_8597,N_8418);
and U8924 (N_8924,N_8467,N_8636);
nor U8925 (N_8925,N_8650,N_8780);
and U8926 (N_8926,N_8671,N_8494);
and U8927 (N_8927,N_8616,N_8782);
and U8928 (N_8928,N_8572,N_8777);
and U8929 (N_8929,N_8734,N_8771);
or U8930 (N_8930,N_8525,N_8412);
and U8931 (N_8931,N_8596,N_8545);
nand U8932 (N_8932,N_8434,N_8732);
nor U8933 (N_8933,N_8755,N_8455);
xor U8934 (N_8934,N_8735,N_8654);
nand U8935 (N_8935,N_8719,N_8602);
xor U8936 (N_8936,N_8465,N_8449);
and U8937 (N_8937,N_8640,N_8791);
or U8938 (N_8938,N_8558,N_8400);
and U8939 (N_8939,N_8512,N_8762);
and U8940 (N_8940,N_8568,N_8402);
and U8941 (N_8941,N_8779,N_8583);
or U8942 (N_8942,N_8560,N_8438);
or U8943 (N_8943,N_8554,N_8745);
xnor U8944 (N_8944,N_8447,N_8729);
nand U8945 (N_8945,N_8775,N_8710);
nand U8946 (N_8946,N_8491,N_8421);
xnor U8947 (N_8947,N_8505,N_8533);
nand U8948 (N_8948,N_8707,N_8424);
nor U8949 (N_8949,N_8510,N_8683);
nor U8950 (N_8950,N_8571,N_8493);
nor U8951 (N_8951,N_8551,N_8706);
or U8952 (N_8952,N_8670,N_8582);
nor U8953 (N_8953,N_8623,N_8564);
nand U8954 (N_8954,N_8490,N_8741);
nor U8955 (N_8955,N_8445,N_8743);
nor U8956 (N_8956,N_8464,N_8763);
or U8957 (N_8957,N_8689,N_8612);
or U8958 (N_8958,N_8709,N_8756);
nor U8959 (N_8959,N_8598,N_8691);
nor U8960 (N_8960,N_8665,N_8790);
and U8961 (N_8961,N_8532,N_8482);
and U8962 (N_8962,N_8513,N_8506);
or U8963 (N_8963,N_8788,N_8542);
or U8964 (N_8964,N_8638,N_8645);
xor U8965 (N_8965,N_8730,N_8573);
and U8966 (N_8966,N_8656,N_8641);
nor U8967 (N_8967,N_8798,N_8516);
nand U8968 (N_8968,N_8646,N_8479);
nand U8969 (N_8969,N_8484,N_8524);
nand U8970 (N_8970,N_8436,N_8471);
nand U8971 (N_8971,N_8799,N_8540);
nand U8972 (N_8972,N_8637,N_8431);
nand U8973 (N_8973,N_8657,N_8487);
xor U8974 (N_8974,N_8722,N_8679);
or U8975 (N_8975,N_8742,N_8518);
nand U8976 (N_8976,N_8685,N_8574);
nand U8977 (N_8977,N_8439,N_8563);
nor U8978 (N_8978,N_8793,N_8521);
or U8979 (N_8979,N_8578,N_8776);
and U8980 (N_8980,N_8446,N_8796);
nor U8981 (N_8981,N_8553,N_8797);
or U8982 (N_8982,N_8441,N_8643);
nor U8983 (N_8983,N_8715,N_8410);
nand U8984 (N_8984,N_8607,N_8659);
and U8985 (N_8985,N_8590,N_8795);
nand U8986 (N_8986,N_8589,N_8498);
nor U8987 (N_8987,N_8409,N_8535);
nor U8988 (N_8988,N_8593,N_8463);
or U8989 (N_8989,N_8781,N_8534);
xor U8990 (N_8990,N_8770,N_8669);
nand U8991 (N_8991,N_8784,N_8420);
nor U8992 (N_8992,N_8537,N_8443);
and U8993 (N_8993,N_8746,N_8680);
or U8994 (N_8994,N_8451,N_8450);
and U8995 (N_8995,N_8661,N_8666);
and U8996 (N_8996,N_8723,N_8727);
nor U8997 (N_8997,N_8427,N_8462);
nand U8998 (N_8998,N_8655,N_8626);
and U8999 (N_8999,N_8736,N_8632);
nor U9000 (N_9000,N_8672,N_8654);
nand U9001 (N_9001,N_8509,N_8710);
or U9002 (N_9002,N_8655,N_8633);
nor U9003 (N_9003,N_8751,N_8553);
and U9004 (N_9004,N_8464,N_8731);
nand U9005 (N_9005,N_8608,N_8790);
and U9006 (N_9006,N_8738,N_8552);
or U9007 (N_9007,N_8615,N_8622);
xor U9008 (N_9008,N_8642,N_8423);
nor U9009 (N_9009,N_8541,N_8473);
and U9010 (N_9010,N_8569,N_8467);
xnor U9011 (N_9011,N_8676,N_8438);
nor U9012 (N_9012,N_8515,N_8751);
xor U9013 (N_9013,N_8568,N_8713);
xnor U9014 (N_9014,N_8686,N_8507);
nor U9015 (N_9015,N_8520,N_8736);
xnor U9016 (N_9016,N_8419,N_8589);
xnor U9017 (N_9017,N_8560,N_8649);
nor U9018 (N_9018,N_8472,N_8761);
xor U9019 (N_9019,N_8619,N_8591);
nor U9020 (N_9020,N_8450,N_8621);
nand U9021 (N_9021,N_8429,N_8794);
xnor U9022 (N_9022,N_8573,N_8536);
xor U9023 (N_9023,N_8418,N_8761);
or U9024 (N_9024,N_8592,N_8769);
and U9025 (N_9025,N_8593,N_8444);
and U9026 (N_9026,N_8680,N_8754);
nor U9027 (N_9027,N_8632,N_8778);
and U9028 (N_9028,N_8548,N_8480);
nand U9029 (N_9029,N_8697,N_8758);
nor U9030 (N_9030,N_8651,N_8615);
xor U9031 (N_9031,N_8751,N_8435);
nor U9032 (N_9032,N_8521,N_8613);
and U9033 (N_9033,N_8426,N_8443);
and U9034 (N_9034,N_8789,N_8658);
nor U9035 (N_9035,N_8689,N_8643);
and U9036 (N_9036,N_8595,N_8786);
nor U9037 (N_9037,N_8540,N_8667);
or U9038 (N_9038,N_8723,N_8711);
and U9039 (N_9039,N_8480,N_8440);
nand U9040 (N_9040,N_8497,N_8650);
and U9041 (N_9041,N_8512,N_8639);
and U9042 (N_9042,N_8501,N_8780);
and U9043 (N_9043,N_8755,N_8583);
or U9044 (N_9044,N_8549,N_8751);
and U9045 (N_9045,N_8612,N_8589);
and U9046 (N_9046,N_8599,N_8513);
xnor U9047 (N_9047,N_8481,N_8604);
nand U9048 (N_9048,N_8441,N_8783);
nand U9049 (N_9049,N_8503,N_8427);
and U9050 (N_9050,N_8788,N_8612);
xor U9051 (N_9051,N_8731,N_8768);
or U9052 (N_9052,N_8555,N_8522);
nand U9053 (N_9053,N_8644,N_8484);
xor U9054 (N_9054,N_8692,N_8665);
and U9055 (N_9055,N_8417,N_8472);
nor U9056 (N_9056,N_8711,N_8703);
nor U9057 (N_9057,N_8626,N_8705);
nor U9058 (N_9058,N_8609,N_8719);
or U9059 (N_9059,N_8443,N_8682);
nor U9060 (N_9060,N_8401,N_8414);
xor U9061 (N_9061,N_8482,N_8589);
nor U9062 (N_9062,N_8576,N_8694);
and U9063 (N_9063,N_8602,N_8648);
nor U9064 (N_9064,N_8598,N_8774);
nand U9065 (N_9065,N_8772,N_8605);
nand U9066 (N_9066,N_8674,N_8416);
xnor U9067 (N_9067,N_8567,N_8711);
and U9068 (N_9068,N_8527,N_8707);
and U9069 (N_9069,N_8442,N_8729);
nand U9070 (N_9070,N_8774,N_8602);
nor U9071 (N_9071,N_8417,N_8457);
nor U9072 (N_9072,N_8561,N_8536);
nand U9073 (N_9073,N_8718,N_8723);
nor U9074 (N_9074,N_8703,N_8503);
and U9075 (N_9075,N_8744,N_8599);
or U9076 (N_9076,N_8536,N_8426);
nor U9077 (N_9077,N_8635,N_8429);
or U9078 (N_9078,N_8557,N_8469);
xor U9079 (N_9079,N_8671,N_8606);
or U9080 (N_9080,N_8499,N_8642);
nor U9081 (N_9081,N_8665,N_8705);
or U9082 (N_9082,N_8741,N_8439);
and U9083 (N_9083,N_8526,N_8637);
nor U9084 (N_9084,N_8436,N_8593);
nand U9085 (N_9085,N_8431,N_8577);
and U9086 (N_9086,N_8640,N_8624);
and U9087 (N_9087,N_8651,N_8791);
nor U9088 (N_9088,N_8656,N_8741);
nand U9089 (N_9089,N_8797,N_8740);
nor U9090 (N_9090,N_8633,N_8546);
and U9091 (N_9091,N_8539,N_8437);
and U9092 (N_9092,N_8439,N_8756);
nand U9093 (N_9093,N_8435,N_8691);
and U9094 (N_9094,N_8579,N_8461);
and U9095 (N_9095,N_8652,N_8657);
xnor U9096 (N_9096,N_8405,N_8721);
nand U9097 (N_9097,N_8645,N_8644);
nor U9098 (N_9098,N_8707,N_8428);
nand U9099 (N_9099,N_8443,N_8716);
xnor U9100 (N_9100,N_8672,N_8484);
xor U9101 (N_9101,N_8527,N_8682);
xor U9102 (N_9102,N_8639,N_8438);
nor U9103 (N_9103,N_8686,N_8646);
and U9104 (N_9104,N_8561,N_8758);
nor U9105 (N_9105,N_8709,N_8627);
or U9106 (N_9106,N_8714,N_8532);
and U9107 (N_9107,N_8784,N_8561);
nor U9108 (N_9108,N_8566,N_8424);
xnor U9109 (N_9109,N_8618,N_8588);
nor U9110 (N_9110,N_8497,N_8633);
nand U9111 (N_9111,N_8460,N_8538);
and U9112 (N_9112,N_8429,N_8775);
xor U9113 (N_9113,N_8675,N_8705);
nor U9114 (N_9114,N_8591,N_8493);
or U9115 (N_9115,N_8498,N_8770);
nor U9116 (N_9116,N_8454,N_8591);
and U9117 (N_9117,N_8541,N_8797);
or U9118 (N_9118,N_8469,N_8651);
or U9119 (N_9119,N_8542,N_8731);
and U9120 (N_9120,N_8509,N_8603);
or U9121 (N_9121,N_8798,N_8613);
nor U9122 (N_9122,N_8477,N_8688);
nand U9123 (N_9123,N_8549,N_8678);
nor U9124 (N_9124,N_8692,N_8449);
nor U9125 (N_9125,N_8430,N_8475);
nor U9126 (N_9126,N_8414,N_8700);
or U9127 (N_9127,N_8652,N_8552);
nor U9128 (N_9128,N_8475,N_8642);
xor U9129 (N_9129,N_8692,N_8536);
nand U9130 (N_9130,N_8719,N_8630);
xnor U9131 (N_9131,N_8609,N_8722);
or U9132 (N_9132,N_8747,N_8402);
nor U9133 (N_9133,N_8641,N_8609);
xnor U9134 (N_9134,N_8612,N_8617);
and U9135 (N_9135,N_8462,N_8775);
and U9136 (N_9136,N_8536,N_8510);
xor U9137 (N_9137,N_8678,N_8574);
and U9138 (N_9138,N_8788,N_8478);
xor U9139 (N_9139,N_8620,N_8664);
nand U9140 (N_9140,N_8591,N_8516);
xor U9141 (N_9141,N_8467,N_8483);
and U9142 (N_9142,N_8568,N_8537);
and U9143 (N_9143,N_8725,N_8530);
xor U9144 (N_9144,N_8625,N_8686);
xnor U9145 (N_9145,N_8406,N_8781);
nand U9146 (N_9146,N_8658,N_8776);
xnor U9147 (N_9147,N_8782,N_8650);
nor U9148 (N_9148,N_8660,N_8404);
and U9149 (N_9149,N_8758,N_8558);
or U9150 (N_9150,N_8796,N_8490);
nand U9151 (N_9151,N_8740,N_8543);
or U9152 (N_9152,N_8504,N_8754);
and U9153 (N_9153,N_8521,N_8759);
nor U9154 (N_9154,N_8508,N_8473);
nor U9155 (N_9155,N_8423,N_8568);
nor U9156 (N_9156,N_8795,N_8615);
or U9157 (N_9157,N_8574,N_8739);
or U9158 (N_9158,N_8764,N_8482);
and U9159 (N_9159,N_8642,N_8582);
and U9160 (N_9160,N_8544,N_8733);
nor U9161 (N_9161,N_8440,N_8455);
or U9162 (N_9162,N_8605,N_8574);
nor U9163 (N_9163,N_8732,N_8635);
xnor U9164 (N_9164,N_8505,N_8658);
nand U9165 (N_9165,N_8744,N_8498);
or U9166 (N_9166,N_8508,N_8697);
nor U9167 (N_9167,N_8456,N_8439);
or U9168 (N_9168,N_8443,N_8611);
nor U9169 (N_9169,N_8457,N_8748);
or U9170 (N_9170,N_8542,N_8677);
or U9171 (N_9171,N_8538,N_8653);
or U9172 (N_9172,N_8761,N_8408);
nand U9173 (N_9173,N_8687,N_8640);
or U9174 (N_9174,N_8632,N_8413);
nor U9175 (N_9175,N_8423,N_8776);
nor U9176 (N_9176,N_8716,N_8610);
nor U9177 (N_9177,N_8687,N_8499);
nand U9178 (N_9178,N_8571,N_8562);
nor U9179 (N_9179,N_8455,N_8674);
or U9180 (N_9180,N_8459,N_8582);
nand U9181 (N_9181,N_8550,N_8793);
nor U9182 (N_9182,N_8626,N_8622);
nor U9183 (N_9183,N_8731,N_8771);
or U9184 (N_9184,N_8487,N_8463);
nand U9185 (N_9185,N_8656,N_8460);
nor U9186 (N_9186,N_8424,N_8531);
nand U9187 (N_9187,N_8797,N_8628);
or U9188 (N_9188,N_8705,N_8481);
xnor U9189 (N_9189,N_8626,N_8729);
and U9190 (N_9190,N_8520,N_8729);
xor U9191 (N_9191,N_8686,N_8739);
or U9192 (N_9192,N_8494,N_8695);
xnor U9193 (N_9193,N_8763,N_8568);
nor U9194 (N_9194,N_8464,N_8756);
or U9195 (N_9195,N_8612,N_8605);
nand U9196 (N_9196,N_8523,N_8482);
nand U9197 (N_9197,N_8402,N_8603);
nand U9198 (N_9198,N_8624,N_8492);
and U9199 (N_9199,N_8457,N_8491);
nand U9200 (N_9200,N_8833,N_9018);
xor U9201 (N_9201,N_8902,N_9075);
nor U9202 (N_9202,N_8858,N_8993);
or U9203 (N_9203,N_8989,N_8957);
xnor U9204 (N_9204,N_9175,N_9125);
and U9205 (N_9205,N_9156,N_9133);
and U9206 (N_9206,N_8882,N_8804);
or U9207 (N_9207,N_9083,N_9136);
nor U9208 (N_9208,N_8958,N_9068);
or U9209 (N_9209,N_9062,N_8938);
nor U9210 (N_9210,N_9003,N_9045);
xor U9211 (N_9211,N_8814,N_8840);
and U9212 (N_9212,N_9076,N_9043);
and U9213 (N_9213,N_8931,N_8849);
xnor U9214 (N_9214,N_8848,N_9177);
nor U9215 (N_9215,N_8866,N_9154);
and U9216 (N_9216,N_9072,N_9058);
or U9217 (N_9217,N_8865,N_8888);
xor U9218 (N_9218,N_9039,N_9164);
or U9219 (N_9219,N_8868,N_9168);
xor U9220 (N_9220,N_9195,N_9052);
nand U9221 (N_9221,N_9189,N_9187);
nand U9222 (N_9222,N_9004,N_8801);
xnor U9223 (N_9223,N_8924,N_8992);
nand U9224 (N_9224,N_9126,N_9051);
nand U9225 (N_9225,N_9042,N_8869);
and U9226 (N_9226,N_8816,N_8912);
xor U9227 (N_9227,N_9146,N_8935);
nand U9228 (N_9228,N_8941,N_9163);
and U9229 (N_9229,N_9088,N_8907);
or U9230 (N_9230,N_8963,N_8889);
nor U9231 (N_9231,N_8988,N_8986);
nand U9232 (N_9232,N_9153,N_8911);
xor U9233 (N_9233,N_8925,N_8921);
nor U9234 (N_9234,N_9169,N_9155);
and U9235 (N_9235,N_9198,N_9047);
xor U9236 (N_9236,N_8861,N_9111);
nand U9237 (N_9237,N_8896,N_9055);
or U9238 (N_9238,N_9103,N_9093);
nand U9239 (N_9239,N_9006,N_8817);
nor U9240 (N_9240,N_9184,N_9030);
nor U9241 (N_9241,N_9167,N_8987);
or U9242 (N_9242,N_8829,N_8835);
xor U9243 (N_9243,N_8980,N_9151);
or U9244 (N_9244,N_8850,N_9110);
xor U9245 (N_9245,N_9007,N_8994);
nand U9246 (N_9246,N_9015,N_8903);
and U9247 (N_9247,N_9165,N_8838);
nor U9248 (N_9248,N_8805,N_8942);
nand U9249 (N_9249,N_8825,N_8933);
or U9250 (N_9250,N_9145,N_8873);
xor U9251 (N_9251,N_9056,N_9095);
nand U9252 (N_9252,N_8915,N_8810);
nor U9253 (N_9253,N_8939,N_9158);
xnor U9254 (N_9254,N_9016,N_8955);
nand U9255 (N_9255,N_8839,N_9193);
or U9256 (N_9256,N_8893,N_9149);
xor U9257 (N_9257,N_8842,N_8818);
or U9258 (N_9258,N_8802,N_8975);
and U9259 (N_9259,N_9192,N_8976);
nor U9260 (N_9260,N_9186,N_8920);
and U9261 (N_9261,N_9053,N_8936);
or U9262 (N_9262,N_9002,N_8949);
nand U9263 (N_9263,N_8905,N_8851);
or U9264 (N_9264,N_8983,N_8885);
and U9265 (N_9265,N_9078,N_9080);
xnor U9266 (N_9266,N_8977,N_8813);
nor U9267 (N_9267,N_8826,N_9098);
nor U9268 (N_9268,N_9019,N_9014);
or U9269 (N_9269,N_8972,N_8953);
xor U9270 (N_9270,N_8952,N_9179);
xnor U9271 (N_9271,N_8996,N_9101);
nor U9272 (N_9272,N_8815,N_9024);
or U9273 (N_9273,N_8830,N_9129);
xnor U9274 (N_9274,N_9140,N_9182);
or U9275 (N_9275,N_8960,N_8959);
and U9276 (N_9276,N_8886,N_8926);
or U9277 (N_9277,N_8875,N_8897);
xor U9278 (N_9278,N_8961,N_9054);
and U9279 (N_9279,N_9181,N_9131);
nor U9280 (N_9280,N_8913,N_8978);
xnor U9281 (N_9281,N_9021,N_9170);
nand U9282 (N_9282,N_8895,N_9176);
and U9283 (N_9283,N_9035,N_9026);
xor U9284 (N_9284,N_9123,N_9032);
nor U9285 (N_9285,N_9127,N_8883);
and U9286 (N_9286,N_9008,N_9115);
or U9287 (N_9287,N_9174,N_8821);
and U9288 (N_9288,N_9041,N_9023);
nand U9289 (N_9289,N_9173,N_9084);
nor U9290 (N_9290,N_8854,N_8878);
nand U9291 (N_9291,N_9022,N_8962);
nor U9292 (N_9292,N_8867,N_9074);
xnor U9293 (N_9293,N_9166,N_8954);
xnor U9294 (N_9294,N_8937,N_9104);
nand U9295 (N_9295,N_8844,N_9124);
xnor U9296 (N_9296,N_9094,N_9005);
nand U9297 (N_9297,N_9147,N_8956);
nand U9298 (N_9298,N_9188,N_9141);
and U9299 (N_9299,N_8890,N_9114);
xor U9300 (N_9300,N_9046,N_9096);
xnor U9301 (N_9301,N_8846,N_9120);
and U9302 (N_9302,N_9117,N_9121);
nand U9303 (N_9303,N_8910,N_8820);
or U9304 (N_9304,N_9064,N_9102);
and U9305 (N_9305,N_8836,N_9190);
xor U9306 (N_9306,N_9057,N_8932);
xor U9307 (N_9307,N_9081,N_8917);
or U9308 (N_9308,N_9161,N_8843);
nor U9309 (N_9309,N_9060,N_8891);
nand U9310 (N_9310,N_8807,N_9118);
and U9311 (N_9311,N_9066,N_9135);
or U9312 (N_9312,N_8806,N_8974);
and U9313 (N_9313,N_8997,N_8863);
or U9314 (N_9314,N_9100,N_9112);
nand U9315 (N_9315,N_8968,N_8811);
or U9316 (N_9316,N_8951,N_8950);
xor U9317 (N_9317,N_8832,N_8874);
and U9318 (N_9318,N_9194,N_8995);
and U9319 (N_9319,N_9172,N_8947);
xor U9320 (N_9320,N_8982,N_9113);
nand U9321 (N_9321,N_9157,N_8899);
nand U9322 (N_9322,N_9150,N_8881);
xnor U9323 (N_9323,N_8857,N_8940);
and U9324 (N_9324,N_8856,N_9086);
xnor U9325 (N_9325,N_8930,N_8837);
xnor U9326 (N_9326,N_9106,N_9063);
or U9327 (N_9327,N_9079,N_9049);
xnor U9328 (N_9328,N_9034,N_8864);
and U9329 (N_9329,N_8943,N_9159);
and U9330 (N_9330,N_9142,N_9082);
nand U9331 (N_9331,N_9009,N_8800);
nor U9332 (N_9332,N_9148,N_8908);
xor U9333 (N_9333,N_8823,N_8822);
nor U9334 (N_9334,N_9180,N_8871);
nand U9335 (N_9335,N_8914,N_9162);
or U9336 (N_9336,N_8990,N_9000);
or U9337 (N_9337,N_8870,N_8879);
nand U9338 (N_9338,N_8999,N_9087);
xnor U9339 (N_9339,N_8803,N_9097);
and U9340 (N_9340,N_9013,N_9059);
nand U9341 (N_9341,N_8985,N_8929);
and U9342 (N_9342,N_9197,N_9077);
or U9343 (N_9343,N_8824,N_9128);
or U9344 (N_9344,N_9048,N_9144);
or U9345 (N_9345,N_9071,N_8845);
nand U9346 (N_9346,N_8852,N_8998);
xnor U9347 (N_9347,N_9090,N_8948);
nor U9348 (N_9348,N_8900,N_8966);
or U9349 (N_9349,N_8901,N_9029);
or U9350 (N_9350,N_8991,N_9139);
nand U9351 (N_9351,N_9040,N_9028);
xnor U9352 (N_9352,N_9033,N_9092);
or U9353 (N_9353,N_8809,N_8918);
xnor U9354 (N_9354,N_8841,N_9152);
nand U9355 (N_9355,N_9017,N_8812);
xnor U9356 (N_9356,N_8828,N_9011);
nor U9357 (N_9357,N_8834,N_8880);
or U9358 (N_9358,N_9012,N_9183);
and U9359 (N_9359,N_9160,N_9020);
or U9360 (N_9360,N_8928,N_8981);
or U9361 (N_9361,N_9099,N_9191);
xor U9362 (N_9362,N_9089,N_9037);
or U9363 (N_9363,N_8892,N_9116);
or U9364 (N_9364,N_8855,N_9107);
xor U9365 (N_9365,N_8884,N_9132);
and U9366 (N_9366,N_8923,N_9108);
nor U9367 (N_9367,N_9119,N_9199);
nand U9368 (N_9368,N_9138,N_9171);
xor U9369 (N_9369,N_8862,N_8922);
nand U9370 (N_9370,N_8819,N_9065);
nand U9371 (N_9371,N_8894,N_9031);
nand U9372 (N_9372,N_8944,N_8827);
xor U9373 (N_9373,N_8934,N_9185);
or U9374 (N_9374,N_9010,N_9073);
or U9375 (N_9375,N_9061,N_8853);
nor U9376 (N_9376,N_8927,N_9196);
nand U9377 (N_9377,N_9130,N_8979);
and U9378 (N_9378,N_8860,N_9044);
nand U9379 (N_9379,N_9025,N_9067);
nor U9380 (N_9380,N_8967,N_8971);
nand U9381 (N_9381,N_8859,N_9050);
nand U9382 (N_9382,N_8969,N_8831);
or U9383 (N_9383,N_8872,N_9036);
or U9384 (N_9384,N_8847,N_9134);
nor U9385 (N_9385,N_8898,N_8973);
xnor U9386 (N_9386,N_9069,N_8984);
or U9387 (N_9387,N_8964,N_9070);
xnor U9388 (N_9388,N_8965,N_9027);
or U9389 (N_9389,N_8916,N_8904);
nor U9390 (N_9390,N_9143,N_9109);
xor U9391 (N_9391,N_8945,N_9085);
and U9392 (N_9392,N_8909,N_9122);
nand U9393 (N_9393,N_8970,N_9091);
nand U9394 (N_9394,N_9105,N_8877);
nand U9395 (N_9395,N_9038,N_8808);
or U9396 (N_9396,N_8946,N_9178);
or U9397 (N_9397,N_9137,N_8887);
or U9398 (N_9398,N_8919,N_8906);
nand U9399 (N_9399,N_8876,N_9001);
and U9400 (N_9400,N_8900,N_8800);
and U9401 (N_9401,N_8990,N_9154);
xnor U9402 (N_9402,N_8854,N_8963);
and U9403 (N_9403,N_8896,N_9007);
xnor U9404 (N_9404,N_8942,N_8907);
and U9405 (N_9405,N_9101,N_9075);
and U9406 (N_9406,N_8936,N_9123);
or U9407 (N_9407,N_9005,N_9166);
and U9408 (N_9408,N_9151,N_9182);
nor U9409 (N_9409,N_9124,N_9055);
nor U9410 (N_9410,N_9004,N_8831);
nand U9411 (N_9411,N_8851,N_8939);
nor U9412 (N_9412,N_8865,N_8944);
or U9413 (N_9413,N_8999,N_9018);
or U9414 (N_9414,N_9182,N_9106);
nand U9415 (N_9415,N_9144,N_8977);
or U9416 (N_9416,N_8811,N_8923);
xnor U9417 (N_9417,N_9182,N_9077);
xnor U9418 (N_9418,N_9038,N_9173);
and U9419 (N_9419,N_8951,N_9026);
xnor U9420 (N_9420,N_9048,N_9118);
or U9421 (N_9421,N_8913,N_8919);
xnor U9422 (N_9422,N_9085,N_8875);
nand U9423 (N_9423,N_9085,N_9062);
nor U9424 (N_9424,N_8838,N_9056);
xnor U9425 (N_9425,N_9017,N_8893);
nor U9426 (N_9426,N_9032,N_9034);
and U9427 (N_9427,N_9055,N_8833);
and U9428 (N_9428,N_8839,N_8835);
nand U9429 (N_9429,N_8988,N_9171);
and U9430 (N_9430,N_9101,N_8811);
xor U9431 (N_9431,N_9160,N_8988);
or U9432 (N_9432,N_8840,N_9145);
xnor U9433 (N_9433,N_9006,N_8987);
xnor U9434 (N_9434,N_8839,N_8812);
or U9435 (N_9435,N_9091,N_9138);
or U9436 (N_9436,N_8997,N_9022);
xnor U9437 (N_9437,N_8907,N_9083);
and U9438 (N_9438,N_8965,N_9128);
nor U9439 (N_9439,N_8953,N_9003);
xor U9440 (N_9440,N_9170,N_9099);
nand U9441 (N_9441,N_9158,N_8904);
nand U9442 (N_9442,N_8865,N_8984);
nand U9443 (N_9443,N_9046,N_8921);
and U9444 (N_9444,N_8878,N_8993);
xor U9445 (N_9445,N_8855,N_9110);
and U9446 (N_9446,N_9078,N_9084);
xnor U9447 (N_9447,N_8852,N_8962);
xnor U9448 (N_9448,N_9053,N_8903);
or U9449 (N_9449,N_8811,N_9124);
and U9450 (N_9450,N_9052,N_9062);
nand U9451 (N_9451,N_8994,N_9018);
nand U9452 (N_9452,N_9063,N_8877);
or U9453 (N_9453,N_8829,N_9176);
nor U9454 (N_9454,N_9125,N_9004);
or U9455 (N_9455,N_9175,N_8826);
and U9456 (N_9456,N_9105,N_9096);
xor U9457 (N_9457,N_9067,N_8864);
or U9458 (N_9458,N_9071,N_9001);
nand U9459 (N_9459,N_8844,N_9122);
and U9460 (N_9460,N_8859,N_9196);
xor U9461 (N_9461,N_9032,N_9061);
or U9462 (N_9462,N_8848,N_9016);
or U9463 (N_9463,N_8931,N_8886);
nand U9464 (N_9464,N_8878,N_9002);
nand U9465 (N_9465,N_9022,N_9036);
or U9466 (N_9466,N_8883,N_8999);
xnor U9467 (N_9467,N_9054,N_8879);
nor U9468 (N_9468,N_9078,N_8870);
or U9469 (N_9469,N_9166,N_8821);
xor U9470 (N_9470,N_8904,N_9017);
xor U9471 (N_9471,N_8858,N_9115);
xnor U9472 (N_9472,N_8997,N_9133);
nand U9473 (N_9473,N_9128,N_9111);
xor U9474 (N_9474,N_9143,N_8869);
nor U9475 (N_9475,N_9018,N_8851);
nor U9476 (N_9476,N_8850,N_8963);
xnor U9477 (N_9477,N_9122,N_8962);
and U9478 (N_9478,N_8969,N_9112);
nor U9479 (N_9479,N_9126,N_9034);
nand U9480 (N_9480,N_9017,N_8830);
and U9481 (N_9481,N_8902,N_8873);
or U9482 (N_9482,N_8834,N_8893);
nand U9483 (N_9483,N_9069,N_8848);
and U9484 (N_9484,N_9005,N_9089);
xor U9485 (N_9485,N_8989,N_9083);
or U9486 (N_9486,N_8906,N_8884);
nand U9487 (N_9487,N_8832,N_9043);
and U9488 (N_9488,N_8854,N_8823);
or U9489 (N_9489,N_9061,N_8996);
and U9490 (N_9490,N_8908,N_8907);
nand U9491 (N_9491,N_8893,N_9190);
xnor U9492 (N_9492,N_9173,N_9004);
xnor U9493 (N_9493,N_8986,N_9159);
nand U9494 (N_9494,N_9193,N_8964);
and U9495 (N_9495,N_9076,N_8954);
nand U9496 (N_9496,N_9066,N_9172);
and U9497 (N_9497,N_8950,N_8998);
nor U9498 (N_9498,N_9190,N_8972);
xor U9499 (N_9499,N_9149,N_9066);
nor U9500 (N_9500,N_8878,N_9075);
xnor U9501 (N_9501,N_8968,N_8874);
xnor U9502 (N_9502,N_8955,N_8872);
xor U9503 (N_9503,N_9061,N_9087);
or U9504 (N_9504,N_8947,N_9044);
and U9505 (N_9505,N_8982,N_9059);
nor U9506 (N_9506,N_9065,N_9070);
xor U9507 (N_9507,N_8813,N_9094);
nor U9508 (N_9508,N_9085,N_8868);
nand U9509 (N_9509,N_8825,N_8958);
nand U9510 (N_9510,N_9130,N_9057);
and U9511 (N_9511,N_9046,N_8970);
or U9512 (N_9512,N_9092,N_8805);
xnor U9513 (N_9513,N_9048,N_9042);
or U9514 (N_9514,N_9095,N_9108);
xor U9515 (N_9515,N_9085,N_9119);
or U9516 (N_9516,N_9088,N_9133);
xnor U9517 (N_9517,N_8991,N_9082);
or U9518 (N_9518,N_8853,N_8801);
and U9519 (N_9519,N_9167,N_8834);
nor U9520 (N_9520,N_8875,N_9172);
nor U9521 (N_9521,N_9098,N_8968);
and U9522 (N_9522,N_9049,N_8990);
or U9523 (N_9523,N_8861,N_9173);
and U9524 (N_9524,N_8879,N_9147);
and U9525 (N_9525,N_9004,N_9131);
or U9526 (N_9526,N_9128,N_8868);
xor U9527 (N_9527,N_8877,N_9017);
or U9528 (N_9528,N_8850,N_9063);
and U9529 (N_9529,N_8830,N_9011);
nor U9530 (N_9530,N_9097,N_9188);
or U9531 (N_9531,N_8906,N_9064);
or U9532 (N_9532,N_9066,N_8816);
and U9533 (N_9533,N_9171,N_9197);
xor U9534 (N_9534,N_9044,N_9184);
nor U9535 (N_9535,N_8879,N_8857);
nor U9536 (N_9536,N_9016,N_9099);
or U9537 (N_9537,N_8837,N_8809);
nand U9538 (N_9538,N_9131,N_9076);
xor U9539 (N_9539,N_8960,N_8812);
nand U9540 (N_9540,N_9082,N_9192);
xor U9541 (N_9541,N_8856,N_8969);
xor U9542 (N_9542,N_9105,N_9125);
and U9543 (N_9543,N_9012,N_8878);
nor U9544 (N_9544,N_8961,N_8886);
or U9545 (N_9545,N_9038,N_9144);
nand U9546 (N_9546,N_8808,N_9098);
or U9547 (N_9547,N_9015,N_8853);
and U9548 (N_9548,N_8977,N_9181);
and U9549 (N_9549,N_8933,N_8835);
or U9550 (N_9550,N_9157,N_8920);
and U9551 (N_9551,N_8985,N_8996);
xor U9552 (N_9552,N_8811,N_9193);
and U9553 (N_9553,N_8980,N_8973);
xnor U9554 (N_9554,N_8918,N_9063);
or U9555 (N_9555,N_9157,N_9094);
nor U9556 (N_9556,N_9139,N_9144);
or U9557 (N_9557,N_9175,N_8811);
nor U9558 (N_9558,N_8943,N_8848);
or U9559 (N_9559,N_9051,N_9195);
or U9560 (N_9560,N_8839,N_8836);
nor U9561 (N_9561,N_8827,N_9018);
or U9562 (N_9562,N_8840,N_9117);
xor U9563 (N_9563,N_9104,N_8916);
xnor U9564 (N_9564,N_8910,N_8929);
nor U9565 (N_9565,N_9153,N_9116);
xnor U9566 (N_9566,N_9147,N_9188);
or U9567 (N_9567,N_8847,N_8828);
or U9568 (N_9568,N_8814,N_9071);
nand U9569 (N_9569,N_9160,N_8875);
nor U9570 (N_9570,N_9021,N_9140);
nor U9571 (N_9571,N_9150,N_8843);
and U9572 (N_9572,N_8888,N_8840);
and U9573 (N_9573,N_8965,N_8867);
or U9574 (N_9574,N_9050,N_8945);
nor U9575 (N_9575,N_9141,N_9110);
and U9576 (N_9576,N_9175,N_8992);
and U9577 (N_9577,N_8965,N_9178);
or U9578 (N_9578,N_9071,N_9015);
or U9579 (N_9579,N_9139,N_9077);
xor U9580 (N_9580,N_8988,N_8800);
nand U9581 (N_9581,N_9189,N_9142);
nor U9582 (N_9582,N_8957,N_8806);
or U9583 (N_9583,N_8968,N_9176);
xnor U9584 (N_9584,N_8838,N_8958);
nor U9585 (N_9585,N_8825,N_9006);
or U9586 (N_9586,N_9001,N_9085);
nor U9587 (N_9587,N_8979,N_8878);
nor U9588 (N_9588,N_8921,N_9111);
nor U9589 (N_9589,N_8911,N_9036);
nand U9590 (N_9590,N_8924,N_9100);
xor U9591 (N_9591,N_8846,N_9117);
nor U9592 (N_9592,N_8954,N_9141);
nand U9593 (N_9593,N_9172,N_8910);
and U9594 (N_9594,N_8987,N_8895);
xnor U9595 (N_9595,N_8819,N_8981);
nor U9596 (N_9596,N_8894,N_8924);
nand U9597 (N_9597,N_8859,N_8865);
nor U9598 (N_9598,N_8984,N_8837);
nand U9599 (N_9599,N_9112,N_9037);
or U9600 (N_9600,N_9262,N_9349);
xnor U9601 (N_9601,N_9361,N_9496);
or U9602 (N_9602,N_9317,N_9222);
and U9603 (N_9603,N_9375,N_9246);
xnor U9604 (N_9604,N_9487,N_9280);
and U9605 (N_9605,N_9338,N_9537);
or U9606 (N_9606,N_9323,N_9208);
or U9607 (N_9607,N_9470,N_9324);
nand U9608 (N_9608,N_9386,N_9554);
and U9609 (N_9609,N_9599,N_9326);
or U9610 (N_9610,N_9396,N_9581);
or U9611 (N_9611,N_9411,N_9365);
or U9612 (N_9612,N_9545,N_9254);
and U9613 (N_9613,N_9500,N_9538);
and U9614 (N_9614,N_9418,N_9582);
xor U9615 (N_9615,N_9283,N_9300);
nor U9616 (N_9616,N_9414,N_9216);
nor U9617 (N_9617,N_9557,N_9281);
or U9618 (N_9618,N_9366,N_9372);
and U9619 (N_9619,N_9244,N_9217);
xor U9620 (N_9620,N_9406,N_9401);
xnor U9621 (N_9621,N_9573,N_9436);
and U9622 (N_9622,N_9315,N_9239);
or U9623 (N_9623,N_9202,N_9577);
or U9624 (N_9624,N_9462,N_9343);
and U9625 (N_9625,N_9229,N_9227);
and U9626 (N_9626,N_9336,N_9201);
or U9627 (N_9627,N_9289,N_9446);
nor U9628 (N_9628,N_9410,N_9498);
nand U9629 (N_9629,N_9256,N_9491);
nand U9630 (N_9630,N_9377,N_9364);
nor U9631 (N_9631,N_9433,N_9541);
xor U9632 (N_9632,N_9274,N_9539);
or U9633 (N_9633,N_9242,N_9298);
nand U9634 (N_9634,N_9532,N_9352);
nand U9635 (N_9635,N_9218,N_9568);
nor U9636 (N_9636,N_9385,N_9322);
nor U9637 (N_9637,N_9556,N_9510);
nor U9638 (N_9638,N_9555,N_9203);
nor U9639 (N_9639,N_9574,N_9445);
nand U9640 (N_9640,N_9296,N_9595);
nor U9641 (N_9641,N_9428,N_9469);
xnor U9642 (N_9642,N_9562,N_9519);
xor U9643 (N_9643,N_9509,N_9454);
and U9644 (N_9644,N_9405,N_9378);
xnor U9645 (N_9645,N_9348,N_9358);
nor U9646 (N_9646,N_9589,N_9291);
nand U9647 (N_9647,N_9327,N_9503);
and U9648 (N_9648,N_9467,N_9564);
nor U9649 (N_9649,N_9294,N_9207);
nor U9650 (N_9650,N_9293,N_9442);
nor U9651 (N_9651,N_9457,N_9515);
and U9652 (N_9652,N_9394,N_9382);
nor U9653 (N_9653,N_9416,N_9219);
xor U9654 (N_9654,N_9429,N_9330);
nor U9655 (N_9655,N_9308,N_9404);
or U9656 (N_9656,N_9286,N_9460);
nor U9657 (N_9657,N_9389,N_9521);
xnor U9658 (N_9658,N_9580,N_9591);
nand U9659 (N_9659,N_9369,N_9448);
and U9660 (N_9660,N_9443,N_9463);
nor U9661 (N_9661,N_9360,N_9493);
xor U9662 (N_9662,N_9535,N_9270);
and U9663 (N_9663,N_9261,N_9536);
nor U9664 (N_9664,N_9517,N_9299);
or U9665 (N_9665,N_9211,N_9277);
nand U9666 (N_9666,N_9345,N_9402);
and U9667 (N_9667,N_9456,N_9504);
xnor U9668 (N_9668,N_9533,N_9282);
nand U9669 (N_9669,N_9214,N_9356);
and U9670 (N_9670,N_9459,N_9260);
nand U9671 (N_9671,N_9347,N_9439);
nor U9672 (N_9672,N_9305,N_9426);
xnor U9673 (N_9673,N_9495,N_9257);
and U9674 (N_9674,N_9477,N_9423);
nor U9675 (N_9675,N_9248,N_9512);
nor U9676 (N_9676,N_9398,N_9335);
nor U9677 (N_9677,N_9507,N_9492);
xnor U9678 (N_9678,N_9523,N_9571);
and U9679 (N_9679,N_9221,N_9430);
or U9680 (N_9680,N_9210,N_9321);
or U9681 (N_9681,N_9553,N_9485);
nand U9682 (N_9682,N_9316,N_9351);
xor U9683 (N_9683,N_9466,N_9547);
nor U9684 (N_9684,N_9204,N_9325);
or U9685 (N_9685,N_9403,N_9267);
nor U9686 (N_9686,N_9306,N_9399);
nor U9687 (N_9687,N_9337,N_9569);
nor U9688 (N_9688,N_9563,N_9419);
nand U9689 (N_9689,N_9596,N_9393);
or U9690 (N_9690,N_9455,N_9530);
and U9691 (N_9691,N_9472,N_9284);
xor U9692 (N_9692,N_9479,N_9359);
nor U9693 (N_9693,N_9272,N_9447);
and U9694 (N_9694,N_9520,N_9384);
and U9695 (N_9695,N_9588,N_9292);
nand U9696 (N_9696,N_9407,N_9339);
or U9697 (N_9697,N_9548,N_9587);
xor U9698 (N_9698,N_9237,N_9258);
or U9699 (N_9699,N_9228,N_9527);
and U9700 (N_9700,N_9309,N_9392);
nor U9701 (N_9701,N_9478,N_9451);
nor U9702 (N_9702,N_9307,N_9566);
nand U9703 (N_9703,N_9576,N_9583);
and U9704 (N_9704,N_9531,N_9561);
nand U9705 (N_9705,N_9444,N_9431);
nor U9706 (N_9706,N_9559,N_9200);
nand U9707 (N_9707,N_9434,N_9544);
or U9708 (N_9708,N_9551,N_9209);
and U9709 (N_9709,N_9318,N_9572);
nor U9710 (N_9710,N_9437,N_9474);
nand U9711 (N_9711,N_9508,N_9251);
nor U9712 (N_9712,N_9379,N_9435);
and U9713 (N_9713,N_9499,N_9213);
and U9714 (N_9714,N_9511,N_9471);
nor U9715 (N_9715,N_9301,N_9333);
xor U9716 (N_9716,N_9481,N_9584);
xor U9717 (N_9717,N_9558,N_9247);
xor U9718 (N_9718,N_9413,N_9391);
nor U9719 (N_9719,N_9543,N_9390);
or U9720 (N_9720,N_9220,N_9355);
nand U9721 (N_9721,N_9250,N_9290);
or U9722 (N_9722,N_9236,N_9233);
xor U9723 (N_9723,N_9505,N_9346);
xnor U9724 (N_9724,N_9464,N_9287);
or U9725 (N_9725,N_9524,N_9367);
or U9726 (N_9726,N_9458,N_9354);
nand U9727 (N_9727,N_9238,N_9331);
nand U9728 (N_9728,N_9542,N_9332);
xor U9729 (N_9729,N_9288,N_9226);
and U9730 (N_9730,N_9395,N_9578);
xnor U9731 (N_9731,N_9313,N_9597);
nand U9732 (N_9732,N_9285,N_9314);
or U9733 (N_9733,N_9415,N_9522);
nor U9734 (N_9734,N_9334,N_9560);
and U9735 (N_9735,N_9265,N_9376);
or U9736 (N_9736,N_9480,N_9231);
and U9737 (N_9737,N_9534,N_9525);
xnor U9738 (N_9738,N_9565,N_9380);
nor U9739 (N_9739,N_9234,N_9513);
xor U9740 (N_9740,N_9362,N_9304);
and U9741 (N_9741,N_9488,N_9465);
nor U9742 (N_9742,N_9422,N_9368);
xor U9743 (N_9743,N_9303,N_9585);
and U9744 (N_9744,N_9461,N_9295);
nor U9745 (N_9745,N_9409,N_9567);
nor U9746 (N_9746,N_9357,N_9205);
xnor U9747 (N_9747,N_9417,N_9206);
or U9748 (N_9748,N_9310,N_9526);
xnor U9749 (N_9749,N_9388,N_9381);
and U9750 (N_9750,N_9490,N_9594);
xor U9751 (N_9751,N_9212,N_9271);
nand U9752 (N_9752,N_9516,N_9438);
and U9753 (N_9753,N_9235,N_9240);
nor U9754 (N_9754,N_9412,N_9424);
xnor U9755 (N_9755,N_9263,N_9328);
or U9756 (N_9756,N_9241,N_9232);
and U9757 (N_9757,N_9276,N_9223);
and U9758 (N_9758,N_9540,N_9476);
and U9759 (N_9759,N_9297,N_9353);
and U9760 (N_9760,N_9506,N_9249);
nor U9761 (N_9761,N_9255,N_9514);
nor U9762 (N_9762,N_9273,N_9344);
xnor U9763 (N_9763,N_9486,N_9484);
or U9764 (N_9764,N_9425,N_9528);
or U9765 (N_9765,N_9592,N_9397);
nor U9766 (N_9766,N_9340,N_9598);
and U9767 (N_9767,N_9550,N_9371);
or U9768 (N_9768,N_9502,N_9494);
nand U9769 (N_9769,N_9400,N_9341);
nand U9770 (N_9770,N_9275,N_9575);
nand U9771 (N_9771,N_9373,N_9549);
nand U9772 (N_9772,N_9529,N_9420);
and U9773 (N_9773,N_9452,N_9312);
nand U9774 (N_9774,N_9311,N_9329);
xor U9775 (N_9775,N_9475,N_9579);
or U9776 (N_9776,N_9224,N_9342);
or U9777 (N_9777,N_9374,N_9268);
and U9778 (N_9778,N_9501,N_9468);
and U9779 (N_9779,N_9482,N_9383);
xor U9780 (N_9780,N_9421,N_9243);
and U9781 (N_9781,N_9449,N_9259);
and U9782 (N_9782,N_9450,N_9266);
and U9783 (N_9783,N_9253,N_9320);
nand U9784 (N_9784,N_9570,N_9215);
nand U9785 (N_9785,N_9489,N_9350);
nand U9786 (N_9786,N_9245,N_9252);
or U9787 (N_9787,N_9552,N_9370);
nor U9788 (N_9788,N_9302,N_9440);
nor U9789 (N_9789,N_9363,N_9483);
xnor U9790 (N_9790,N_9546,N_9432);
and U9791 (N_9791,N_9319,N_9269);
xnor U9792 (N_9792,N_9518,N_9441);
or U9793 (N_9793,N_9590,N_9408);
xnor U9794 (N_9794,N_9453,N_9279);
nor U9795 (N_9795,N_9278,N_9497);
and U9796 (N_9796,N_9473,N_9230);
and U9797 (N_9797,N_9225,N_9264);
nand U9798 (N_9798,N_9387,N_9586);
xor U9799 (N_9799,N_9593,N_9427);
xor U9800 (N_9800,N_9521,N_9296);
and U9801 (N_9801,N_9548,N_9526);
nor U9802 (N_9802,N_9591,N_9505);
nand U9803 (N_9803,N_9237,N_9316);
nand U9804 (N_9804,N_9515,N_9514);
or U9805 (N_9805,N_9265,N_9491);
xor U9806 (N_9806,N_9271,N_9312);
nor U9807 (N_9807,N_9230,N_9337);
and U9808 (N_9808,N_9344,N_9214);
or U9809 (N_9809,N_9543,N_9549);
and U9810 (N_9810,N_9264,N_9466);
and U9811 (N_9811,N_9541,N_9339);
or U9812 (N_9812,N_9215,N_9329);
and U9813 (N_9813,N_9372,N_9475);
xor U9814 (N_9814,N_9595,N_9358);
nor U9815 (N_9815,N_9303,N_9592);
nor U9816 (N_9816,N_9343,N_9213);
or U9817 (N_9817,N_9534,N_9491);
and U9818 (N_9818,N_9254,N_9359);
nand U9819 (N_9819,N_9569,N_9219);
and U9820 (N_9820,N_9306,N_9470);
or U9821 (N_9821,N_9362,N_9363);
and U9822 (N_9822,N_9557,N_9278);
nor U9823 (N_9823,N_9506,N_9519);
nor U9824 (N_9824,N_9557,N_9267);
or U9825 (N_9825,N_9447,N_9537);
xor U9826 (N_9826,N_9506,N_9305);
or U9827 (N_9827,N_9404,N_9244);
xor U9828 (N_9828,N_9294,N_9286);
xor U9829 (N_9829,N_9408,N_9221);
xnor U9830 (N_9830,N_9329,N_9221);
xnor U9831 (N_9831,N_9244,N_9255);
or U9832 (N_9832,N_9206,N_9320);
nand U9833 (N_9833,N_9241,N_9352);
and U9834 (N_9834,N_9275,N_9437);
nor U9835 (N_9835,N_9504,N_9535);
xor U9836 (N_9836,N_9459,N_9536);
or U9837 (N_9837,N_9257,N_9249);
nand U9838 (N_9838,N_9412,N_9509);
and U9839 (N_9839,N_9560,N_9365);
or U9840 (N_9840,N_9364,N_9342);
nand U9841 (N_9841,N_9213,N_9231);
xor U9842 (N_9842,N_9507,N_9385);
nor U9843 (N_9843,N_9377,N_9500);
nand U9844 (N_9844,N_9540,N_9510);
or U9845 (N_9845,N_9398,N_9527);
nor U9846 (N_9846,N_9261,N_9301);
and U9847 (N_9847,N_9294,N_9484);
or U9848 (N_9848,N_9240,N_9287);
nand U9849 (N_9849,N_9542,N_9452);
xor U9850 (N_9850,N_9288,N_9446);
or U9851 (N_9851,N_9518,N_9391);
nor U9852 (N_9852,N_9377,N_9553);
nand U9853 (N_9853,N_9423,N_9583);
xnor U9854 (N_9854,N_9539,N_9595);
nor U9855 (N_9855,N_9228,N_9264);
or U9856 (N_9856,N_9440,N_9429);
nor U9857 (N_9857,N_9470,N_9573);
nand U9858 (N_9858,N_9586,N_9570);
xnor U9859 (N_9859,N_9514,N_9323);
or U9860 (N_9860,N_9268,N_9494);
nor U9861 (N_9861,N_9460,N_9434);
and U9862 (N_9862,N_9384,N_9572);
or U9863 (N_9863,N_9375,N_9215);
xnor U9864 (N_9864,N_9502,N_9350);
xor U9865 (N_9865,N_9210,N_9264);
nand U9866 (N_9866,N_9397,N_9342);
or U9867 (N_9867,N_9541,N_9573);
or U9868 (N_9868,N_9439,N_9418);
nand U9869 (N_9869,N_9350,N_9265);
and U9870 (N_9870,N_9530,N_9543);
or U9871 (N_9871,N_9505,N_9469);
and U9872 (N_9872,N_9522,N_9397);
nor U9873 (N_9873,N_9317,N_9265);
or U9874 (N_9874,N_9380,N_9481);
nand U9875 (N_9875,N_9504,N_9200);
nand U9876 (N_9876,N_9252,N_9344);
xor U9877 (N_9877,N_9237,N_9268);
nand U9878 (N_9878,N_9558,N_9238);
nor U9879 (N_9879,N_9217,N_9395);
or U9880 (N_9880,N_9534,N_9368);
xor U9881 (N_9881,N_9537,N_9591);
and U9882 (N_9882,N_9576,N_9456);
nand U9883 (N_9883,N_9374,N_9561);
nor U9884 (N_9884,N_9229,N_9384);
or U9885 (N_9885,N_9436,N_9255);
or U9886 (N_9886,N_9368,N_9494);
or U9887 (N_9887,N_9403,N_9292);
xnor U9888 (N_9888,N_9545,N_9492);
nor U9889 (N_9889,N_9443,N_9455);
nand U9890 (N_9890,N_9350,N_9381);
and U9891 (N_9891,N_9594,N_9241);
and U9892 (N_9892,N_9556,N_9520);
nand U9893 (N_9893,N_9483,N_9411);
nand U9894 (N_9894,N_9390,N_9259);
nand U9895 (N_9895,N_9530,N_9250);
nor U9896 (N_9896,N_9243,N_9367);
and U9897 (N_9897,N_9458,N_9231);
xnor U9898 (N_9898,N_9221,N_9394);
nor U9899 (N_9899,N_9546,N_9466);
xor U9900 (N_9900,N_9267,N_9418);
nor U9901 (N_9901,N_9465,N_9205);
and U9902 (N_9902,N_9411,N_9430);
nor U9903 (N_9903,N_9414,N_9483);
or U9904 (N_9904,N_9392,N_9543);
or U9905 (N_9905,N_9402,N_9368);
xor U9906 (N_9906,N_9568,N_9527);
nor U9907 (N_9907,N_9466,N_9583);
and U9908 (N_9908,N_9211,N_9456);
and U9909 (N_9909,N_9449,N_9232);
and U9910 (N_9910,N_9420,N_9595);
or U9911 (N_9911,N_9223,N_9494);
nor U9912 (N_9912,N_9412,N_9581);
nor U9913 (N_9913,N_9336,N_9541);
and U9914 (N_9914,N_9480,N_9587);
nand U9915 (N_9915,N_9349,N_9244);
and U9916 (N_9916,N_9348,N_9229);
or U9917 (N_9917,N_9491,N_9370);
xor U9918 (N_9918,N_9431,N_9284);
and U9919 (N_9919,N_9212,N_9428);
and U9920 (N_9920,N_9316,N_9329);
nor U9921 (N_9921,N_9316,N_9307);
and U9922 (N_9922,N_9428,N_9318);
and U9923 (N_9923,N_9307,N_9321);
or U9924 (N_9924,N_9438,N_9223);
and U9925 (N_9925,N_9486,N_9228);
or U9926 (N_9926,N_9297,N_9455);
xor U9927 (N_9927,N_9203,N_9254);
nor U9928 (N_9928,N_9588,N_9351);
xor U9929 (N_9929,N_9284,N_9245);
nor U9930 (N_9930,N_9488,N_9422);
and U9931 (N_9931,N_9353,N_9356);
and U9932 (N_9932,N_9364,N_9315);
and U9933 (N_9933,N_9361,N_9321);
and U9934 (N_9934,N_9424,N_9569);
nand U9935 (N_9935,N_9392,N_9207);
nor U9936 (N_9936,N_9465,N_9500);
nor U9937 (N_9937,N_9489,N_9509);
or U9938 (N_9938,N_9260,N_9297);
xor U9939 (N_9939,N_9456,N_9252);
and U9940 (N_9940,N_9504,N_9306);
and U9941 (N_9941,N_9254,N_9318);
or U9942 (N_9942,N_9263,N_9366);
nor U9943 (N_9943,N_9521,N_9532);
or U9944 (N_9944,N_9510,N_9388);
nor U9945 (N_9945,N_9258,N_9517);
nand U9946 (N_9946,N_9247,N_9384);
nor U9947 (N_9947,N_9517,N_9433);
xor U9948 (N_9948,N_9358,N_9534);
or U9949 (N_9949,N_9343,N_9275);
nand U9950 (N_9950,N_9389,N_9372);
or U9951 (N_9951,N_9494,N_9545);
xor U9952 (N_9952,N_9400,N_9482);
nor U9953 (N_9953,N_9355,N_9474);
nor U9954 (N_9954,N_9284,N_9485);
nand U9955 (N_9955,N_9574,N_9586);
xnor U9956 (N_9956,N_9538,N_9366);
and U9957 (N_9957,N_9444,N_9200);
nor U9958 (N_9958,N_9572,N_9417);
xor U9959 (N_9959,N_9484,N_9447);
xor U9960 (N_9960,N_9494,N_9204);
nor U9961 (N_9961,N_9232,N_9300);
nand U9962 (N_9962,N_9419,N_9537);
and U9963 (N_9963,N_9577,N_9592);
or U9964 (N_9964,N_9515,N_9345);
or U9965 (N_9965,N_9396,N_9510);
nor U9966 (N_9966,N_9355,N_9464);
xnor U9967 (N_9967,N_9592,N_9349);
nand U9968 (N_9968,N_9575,N_9502);
xor U9969 (N_9969,N_9488,N_9203);
nand U9970 (N_9970,N_9363,N_9432);
or U9971 (N_9971,N_9323,N_9276);
xnor U9972 (N_9972,N_9226,N_9381);
xor U9973 (N_9973,N_9559,N_9382);
nand U9974 (N_9974,N_9520,N_9251);
xnor U9975 (N_9975,N_9499,N_9311);
xor U9976 (N_9976,N_9537,N_9450);
or U9977 (N_9977,N_9504,N_9466);
and U9978 (N_9978,N_9380,N_9330);
and U9979 (N_9979,N_9438,N_9578);
or U9980 (N_9980,N_9554,N_9580);
and U9981 (N_9981,N_9245,N_9228);
nor U9982 (N_9982,N_9341,N_9283);
nand U9983 (N_9983,N_9574,N_9347);
and U9984 (N_9984,N_9279,N_9414);
nand U9985 (N_9985,N_9260,N_9214);
nor U9986 (N_9986,N_9494,N_9507);
and U9987 (N_9987,N_9463,N_9204);
or U9988 (N_9988,N_9418,N_9276);
or U9989 (N_9989,N_9566,N_9564);
and U9990 (N_9990,N_9474,N_9315);
nand U9991 (N_9991,N_9358,N_9441);
nand U9992 (N_9992,N_9471,N_9276);
nand U9993 (N_9993,N_9324,N_9552);
or U9994 (N_9994,N_9599,N_9204);
and U9995 (N_9995,N_9591,N_9458);
xor U9996 (N_9996,N_9596,N_9287);
nand U9997 (N_9997,N_9236,N_9576);
or U9998 (N_9998,N_9386,N_9457);
nand U9999 (N_9999,N_9351,N_9498);
or U10000 (N_10000,N_9688,N_9879);
nand U10001 (N_10001,N_9780,N_9733);
nor U10002 (N_10002,N_9942,N_9964);
nand U10003 (N_10003,N_9807,N_9700);
nor U10004 (N_10004,N_9954,N_9701);
nand U10005 (N_10005,N_9704,N_9644);
xor U10006 (N_10006,N_9680,N_9927);
or U10007 (N_10007,N_9662,N_9978);
nor U10008 (N_10008,N_9961,N_9721);
nor U10009 (N_10009,N_9606,N_9820);
nor U10010 (N_10010,N_9994,N_9660);
and U10011 (N_10011,N_9819,N_9873);
or U10012 (N_10012,N_9656,N_9811);
xnor U10013 (N_10013,N_9789,N_9816);
nand U10014 (N_10014,N_9950,N_9874);
xor U10015 (N_10015,N_9695,N_9933);
and U10016 (N_10016,N_9792,N_9751);
xnor U10017 (N_10017,N_9777,N_9666);
and U10018 (N_10018,N_9960,N_9831);
nand U10019 (N_10019,N_9737,N_9713);
nor U10020 (N_10020,N_9823,N_9636);
nor U10021 (N_10021,N_9776,N_9650);
xor U10022 (N_10022,N_9817,N_9800);
xor U10023 (N_10023,N_9735,N_9767);
or U10024 (N_10024,N_9798,N_9769);
or U10025 (N_10025,N_9602,N_9901);
nor U10026 (N_10026,N_9959,N_9762);
and U10027 (N_10027,N_9743,N_9795);
nand U10028 (N_10028,N_9752,N_9943);
nor U10029 (N_10029,N_9782,N_9673);
or U10030 (N_10030,N_9870,N_9815);
nand U10031 (N_10031,N_9856,N_9771);
or U10032 (N_10032,N_9672,N_9936);
xnor U10033 (N_10033,N_9890,N_9685);
xnor U10034 (N_10034,N_9615,N_9955);
nand U10035 (N_10035,N_9681,N_9896);
nor U10036 (N_10036,N_9931,N_9854);
nand U10037 (N_10037,N_9640,N_9894);
nand U10038 (N_10038,N_9665,N_9965);
and U10039 (N_10039,N_9711,N_9729);
xor U10040 (N_10040,N_9679,N_9625);
xnor U10041 (N_10041,N_9832,N_9603);
xor U10042 (N_10042,N_9853,N_9757);
nand U10043 (N_10043,N_9750,N_9635);
nor U10044 (N_10044,N_9953,N_9781);
nand U10045 (N_10045,N_9663,N_9710);
xnor U10046 (N_10046,N_9884,N_9814);
or U10047 (N_10047,N_9667,N_9696);
nand U10048 (N_10048,N_9651,N_9984);
nor U10049 (N_10049,N_9813,N_9722);
nand U10050 (N_10050,N_9827,N_9968);
or U10051 (N_10051,N_9639,N_9844);
and U10052 (N_10052,N_9684,N_9718);
or U10053 (N_10053,N_9637,N_9956);
nor U10054 (N_10054,N_9846,N_9694);
or U10055 (N_10055,N_9627,N_9971);
and U10056 (N_10056,N_9612,N_9987);
or U10057 (N_10057,N_9834,N_9728);
nor U10058 (N_10058,N_9826,N_9855);
and U10059 (N_10059,N_9939,N_9706);
nor U10060 (N_10060,N_9726,N_9993);
xnor U10061 (N_10061,N_9716,N_9812);
or U10062 (N_10062,N_9628,N_9608);
xor U10063 (N_10063,N_9766,N_9648);
nor U10064 (N_10064,N_9919,N_9768);
xnor U10065 (N_10065,N_9934,N_9938);
nand U10066 (N_10066,N_9916,N_9881);
nor U10067 (N_10067,N_9828,N_9727);
nor U10068 (N_10068,N_9868,N_9958);
xor U10069 (N_10069,N_9808,N_9617);
or U10070 (N_10070,N_9745,N_9742);
nand U10071 (N_10071,N_9744,N_9730);
and U10072 (N_10072,N_9906,N_9990);
xnor U10073 (N_10073,N_9849,N_9842);
nor U10074 (N_10074,N_9654,N_9822);
nor U10075 (N_10075,N_9880,N_9836);
nand U10076 (N_10076,N_9793,N_9783);
and U10077 (N_10077,N_9758,N_9903);
xnor U10078 (N_10078,N_9765,N_9966);
and U10079 (N_10079,N_9703,N_9979);
or U10080 (N_10080,N_9661,N_9669);
nand U10081 (N_10081,N_9980,N_9804);
and U10082 (N_10082,N_9940,N_9859);
nand U10083 (N_10083,N_9773,N_9611);
and U10084 (N_10084,N_9902,N_9806);
and U10085 (N_10085,N_9788,N_9922);
nor U10086 (N_10086,N_9796,N_9652);
nor U10087 (N_10087,N_9988,N_9801);
xor U10088 (N_10088,N_9653,N_9852);
xor U10089 (N_10089,N_9967,N_9848);
nand U10090 (N_10090,N_9893,N_9837);
xor U10091 (N_10091,N_9920,N_9865);
and U10092 (N_10092,N_9803,N_9835);
xnor U10093 (N_10093,N_9818,N_9671);
nand U10094 (N_10094,N_9618,N_9824);
nor U10095 (N_10095,N_9882,N_9915);
xnor U10096 (N_10096,N_9791,N_9948);
xor U10097 (N_10097,N_9974,N_9887);
and U10098 (N_10098,N_9877,N_9784);
and U10099 (N_10099,N_9851,N_9946);
nor U10100 (N_10100,N_9949,N_9872);
nor U10101 (N_10101,N_9907,N_9712);
nand U10102 (N_10102,N_9682,N_9996);
nor U10103 (N_10103,N_9624,N_9995);
or U10104 (N_10104,N_9962,N_9969);
or U10105 (N_10105,N_9951,N_9763);
and U10106 (N_10106,N_9715,N_9925);
nor U10107 (N_10107,N_9687,N_9862);
nand U10108 (N_10108,N_9697,N_9892);
nand U10109 (N_10109,N_9693,N_9629);
or U10110 (N_10110,N_9747,N_9829);
nor U10111 (N_10111,N_9778,N_9785);
xnor U10112 (N_10112,N_9898,N_9674);
or U10113 (N_10113,N_9690,N_9989);
and U10114 (N_10114,N_9647,N_9719);
nand U10115 (N_10115,N_9913,N_9932);
nand U10116 (N_10116,N_9850,N_9992);
or U10117 (N_10117,N_9634,N_9642);
and U10118 (N_10118,N_9857,N_9866);
nor U10119 (N_10119,N_9912,N_9923);
nand U10120 (N_10120,N_9613,N_9924);
xnor U10121 (N_10121,N_9621,N_9708);
nor U10122 (N_10122,N_9741,N_9875);
nor U10123 (N_10123,N_9734,N_9620);
nor U10124 (N_10124,N_9626,N_9658);
nand U10125 (N_10125,N_9977,N_9957);
and U10126 (N_10126,N_9632,N_9668);
nor U10127 (N_10127,N_9926,N_9645);
or U10128 (N_10128,N_9997,N_9731);
nand U10129 (N_10129,N_9664,N_9619);
nand U10130 (N_10130,N_9952,N_9717);
nand U10131 (N_10131,N_9764,N_9600);
and U10132 (N_10132,N_9963,N_9790);
nor U10133 (N_10133,N_9886,N_9888);
xnor U10134 (N_10134,N_9840,N_9659);
nor U10135 (N_10135,N_9623,N_9909);
and U10136 (N_10136,N_9889,N_9941);
nand U10137 (N_10137,N_9775,N_9843);
xor U10138 (N_10138,N_9676,N_9761);
nor U10139 (N_10139,N_9643,N_9830);
or U10140 (N_10140,N_9723,N_9918);
xnor U10141 (N_10141,N_9641,N_9839);
and U10142 (N_10142,N_9805,N_9675);
and U10143 (N_10143,N_9905,N_9759);
nor U10144 (N_10144,N_9714,N_9770);
nand U10145 (N_10145,N_9895,N_9983);
nand U10146 (N_10146,N_9833,N_9860);
nand U10147 (N_10147,N_9809,N_9885);
xnor U10148 (N_10148,N_9739,N_9947);
nand U10149 (N_10149,N_9930,N_9614);
xnor U10150 (N_10150,N_9655,N_9910);
nand U10151 (N_10151,N_9616,N_9601);
and U10152 (N_10152,N_9698,N_9670);
and U10153 (N_10153,N_9749,N_9883);
nor U10154 (N_10154,N_9867,N_9702);
and U10155 (N_10155,N_9736,N_9631);
and U10156 (N_10156,N_9755,N_9838);
nor U10157 (N_10157,N_9797,N_9861);
nand U10158 (N_10158,N_9756,N_9982);
nand U10159 (N_10159,N_9891,N_9649);
nor U10160 (N_10160,N_9630,N_9707);
nand U10161 (N_10161,N_9917,N_9841);
or U10162 (N_10162,N_9864,N_9802);
nand U10163 (N_10163,N_9604,N_9774);
or U10164 (N_10164,N_9876,N_9858);
or U10165 (N_10165,N_9845,N_9646);
xor U10166 (N_10166,N_9689,N_9760);
nand U10167 (N_10167,N_9657,N_9945);
or U10168 (N_10168,N_9929,N_9677);
and U10169 (N_10169,N_9683,N_9691);
nor U10170 (N_10170,N_9904,N_9976);
nand U10171 (N_10171,N_9732,N_9970);
nand U10172 (N_10172,N_9869,N_9821);
nor U10173 (N_10173,N_9692,N_9738);
nor U10174 (N_10174,N_9638,N_9724);
xor U10175 (N_10175,N_9863,N_9699);
nand U10176 (N_10176,N_9911,N_9985);
nand U10177 (N_10177,N_9779,N_9610);
nand U10178 (N_10178,N_9678,N_9794);
xor U10179 (N_10179,N_9944,N_9825);
xor U10180 (N_10180,N_9753,N_9871);
or U10181 (N_10181,N_9921,N_9786);
nor U10182 (N_10182,N_9937,N_9725);
and U10183 (N_10183,N_9899,N_9975);
or U10184 (N_10184,N_9709,N_9772);
nand U10185 (N_10185,N_9900,N_9981);
and U10186 (N_10186,N_9705,N_9607);
and U10187 (N_10187,N_9847,N_9754);
nor U10188 (N_10188,N_9999,N_9810);
nor U10189 (N_10189,N_9991,N_9928);
xor U10190 (N_10190,N_9740,N_9914);
nand U10191 (N_10191,N_9799,N_9622);
nand U10192 (N_10192,N_9605,N_9998);
xor U10193 (N_10193,N_9935,N_9878);
nor U10194 (N_10194,N_9973,N_9609);
or U10195 (N_10195,N_9897,N_9720);
and U10196 (N_10196,N_9633,N_9748);
and U10197 (N_10197,N_9787,N_9686);
and U10198 (N_10198,N_9746,N_9986);
or U10199 (N_10199,N_9908,N_9972);
nor U10200 (N_10200,N_9982,N_9835);
xor U10201 (N_10201,N_9908,N_9757);
and U10202 (N_10202,N_9799,N_9823);
nand U10203 (N_10203,N_9835,N_9612);
and U10204 (N_10204,N_9624,N_9677);
nand U10205 (N_10205,N_9610,N_9803);
nor U10206 (N_10206,N_9959,N_9726);
nor U10207 (N_10207,N_9903,N_9668);
or U10208 (N_10208,N_9658,N_9794);
nor U10209 (N_10209,N_9798,N_9890);
nor U10210 (N_10210,N_9671,N_9851);
xnor U10211 (N_10211,N_9765,N_9757);
and U10212 (N_10212,N_9723,N_9665);
nand U10213 (N_10213,N_9836,N_9783);
and U10214 (N_10214,N_9806,N_9849);
nand U10215 (N_10215,N_9660,N_9612);
nand U10216 (N_10216,N_9784,N_9737);
or U10217 (N_10217,N_9810,N_9707);
nand U10218 (N_10218,N_9689,N_9920);
xnor U10219 (N_10219,N_9774,N_9962);
and U10220 (N_10220,N_9783,N_9984);
and U10221 (N_10221,N_9948,N_9672);
nand U10222 (N_10222,N_9756,N_9602);
or U10223 (N_10223,N_9671,N_9968);
nand U10224 (N_10224,N_9830,N_9903);
nand U10225 (N_10225,N_9811,N_9665);
xnor U10226 (N_10226,N_9916,N_9781);
xnor U10227 (N_10227,N_9674,N_9651);
and U10228 (N_10228,N_9880,N_9973);
xor U10229 (N_10229,N_9713,N_9805);
xor U10230 (N_10230,N_9797,N_9805);
or U10231 (N_10231,N_9978,N_9960);
and U10232 (N_10232,N_9881,N_9917);
nand U10233 (N_10233,N_9997,N_9681);
nor U10234 (N_10234,N_9989,N_9804);
nor U10235 (N_10235,N_9711,N_9925);
xor U10236 (N_10236,N_9648,N_9821);
nand U10237 (N_10237,N_9812,N_9605);
nand U10238 (N_10238,N_9972,N_9758);
xnor U10239 (N_10239,N_9957,N_9717);
nor U10240 (N_10240,N_9970,N_9679);
nand U10241 (N_10241,N_9899,N_9855);
xnor U10242 (N_10242,N_9799,N_9812);
nand U10243 (N_10243,N_9727,N_9889);
xnor U10244 (N_10244,N_9774,N_9937);
xnor U10245 (N_10245,N_9753,N_9985);
or U10246 (N_10246,N_9933,N_9799);
xor U10247 (N_10247,N_9883,N_9855);
and U10248 (N_10248,N_9739,N_9890);
xnor U10249 (N_10249,N_9920,N_9705);
nand U10250 (N_10250,N_9814,N_9751);
xor U10251 (N_10251,N_9698,N_9683);
nor U10252 (N_10252,N_9805,N_9841);
xor U10253 (N_10253,N_9787,N_9602);
nor U10254 (N_10254,N_9825,N_9700);
nor U10255 (N_10255,N_9993,N_9873);
xnor U10256 (N_10256,N_9697,N_9804);
and U10257 (N_10257,N_9717,N_9715);
or U10258 (N_10258,N_9753,N_9651);
nand U10259 (N_10259,N_9944,N_9727);
and U10260 (N_10260,N_9809,N_9833);
or U10261 (N_10261,N_9649,N_9933);
or U10262 (N_10262,N_9920,N_9812);
and U10263 (N_10263,N_9881,N_9926);
xor U10264 (N_10264,N_9804,N_9858);
nor U10265 (N_10265,N_9974,N_9975);
xnor U10266 (N_10266,N_9612,N_9874);
or U10267 (N_10267,N_9814,N_9984);
and U10268 (N_10268,N_9660,N_9627);
nor U10269 (N_10269,N_9829,N_9798);
nor U10270 (N_10270,N_9931,N_9925);
xnor U10271 (N_10271,N_9935,N_9862);
or U10272 (N_10272,N_9899,N_9639);
and U10273 (N_10273,N_9648,N_9700);
and U10274 (N_10274,N_9767,N_9831);
nor U10275 (N_10275,N_9756,N_9868);
nor U10276 (N_10276,N_9933,N_9693);
nor U10277 (N_10277,N_9891,N_9940);
xnor U10278 (N_10278,N_9725,N_9709);
or U10279 (N_10279,N_9731,N_9689);
and U10280 (N_10280,N_9726,N_9607);
or U10281 (N_10281,N_9914,N_9692);
xor U10282 (N_10282,N_9616,N_9880);
xor U10283 (N_10283,N_9650,N_9759);
or U10284 (N_10284,N_9795,N_9709);
xnor U10285 (N_10285,N_9687,N_9909);
nor U10286 (N_10286,N_9984,N_9953);
nand U10287 (N_10287,N_9890,N_9858);
nor U10288 (N_10288,N_9841,N_9797);
or U10289 (N_10289,N_9938,N_9834);
nand U10290 (N_10290,N_9629,N_9968);
xor U10291 (N_10291,N_9793,N_9808);
or U10292 (N_10292,N_9779,N_9869);
and U10293 (N_10293,N_9931,N_9781);
nand U10294 (N_10294,N_9961,N_9869);
or U10295 (N_10295,N_9836,N_9918);
nor U10296 (N_10296,N_9841,N_9646);
nand U10297 (N_10297,N_9885,N_9991);
nor U10298 (N_10298,N_9873,N_9957);
or U10299 (N_10299,N_9620,N_9763);
xor U10300 (N_10300,N_9726,N_9655);
or U10301 (N_10301,N_9638,N_9951);
xnor U10302 (N_10302,N_9719,N_9841);
xor U10303 (N_10303,N_9705,N_9862);
nor U10304 (N_10304,N_9666,N_9840);
nand U10305 (N_10305,N_9714,N_9769);
or U10306 (N_10306,N_9814,N_9712);
or U10307 (N_10307,N_9799,N_9894);
xnor U10308 (N_10308,N_9747,N_9675);
xor U10309 (N_10309,N_9931,N_9770);
nand U10310 (N_10310,N_9780,N_9911);
nand U10311 (N_10311,N_9769,N_9606);
or U10312 (N_10312,N_9614,N_9624);
nand U10313 (N_10313,N_9792,N_9625);
xor U10314 (N_10314,N_9619,N_9737);
xor U10315 (N_10315,N_9893,N_9937);
nand U10316 (N_10316,N_9616,N_9709);
nor U10317 (N_10317,N_9826,N_9933);
xnor U10318 (N_10318,N_9637,N_9817);
nand U10319 (N_10319,N_9797,N_9967);
nor U10320 (N_10320,N_9782,N_9715);
xor U10321 (N_10321,N_9607,N_9716);
nand U10322 (N_10322,N_9839,N_9673);
or U10323 (N_10323,N_9882,N_9707);
nor U10324 (N_10324,N_9835,N_9702);
nor U10325 (N_10325,N_9823,N_9976);
nor U10326 (N_10326,N_9656,N_9662);
or U10327 (N_10327,N_9838,N_9805);
nand U10328 (N_10328,N_9640,N_9863);
xor U10329 (N_10329,N_9815,N_9911);
or U10330 (N_10330,N_9633,N_9833);
and U10331 (N_10331,N_9767,N_9855);
nor U10332 (N_10332,N_9954,N_9647);
nand U10333 (N_10333,N_9605,N_9911);
and U10334 (N_10334,N_9859,N_9899);
nand U10335 (N_10335,N_9829,N_9938);
nand U10336 (N_10336,N_9625,N_9899);
xnor U10337 (N_10337,N_9763,N_9760);
nor U10338 (N_10338,N_9701,N_9820);
nand U10339 (N_10339,N_9696,N_9726);
or U10340 (N_10340,N_9806,N_9959);
nor U10341 (N_10341,N_9647,N_9827);
nor U10342 (N_10342,N_9778,N_9832);
and U10343 (N_10343,N_9989,N_9806);
nand U10344 (N_10344,N_9670,N_9944);
or U10345 (N_10345,N_9776,N_9703);
xnor U10346 (N_10346,N_9932,N_9844);
xor U10347 (N_10347,N_9737,N_9608);
nand U10348 (N_10348,N_9866,N_9638);
nor U10349 (N_10349,N_9855,N_9809);
xor U10350 (N_10350,N_9700,N_9917);
xnor U10351 (N_10351,N_9664,N_9869);
nor U10352 (N_10352,N_9801,N_9993);
nand U10353 (N_10353,N_9784,N_9835);
and U10354 (N_10354,N_9844,N_9668);
and U10355 (N_10355,N_9759,N_9901);
nor U10356 (N_10356,N_9871,N_9731);
or U10357 (N_10357,N_9655,N_9611);
nor U10358 (N_10358,N_9984,N_9658);
xnor U10359 (N_10359,N_9889,N_9830);
nor U10360 (N_10360,N_9609,N_9863);
nand U10361 (N_10361,N_9996,N_9742);
xnor U10362 (N_10362,N_9855,N_9784);
or U10363 (N_10363,N_9945,N_9831);
or U10364 (N_10364,N_9752,N_9920);
or U10365 (N_10365,N_9988,N_9673);
xor U10366 (N_10366,N_9769,N_9748);
nor U10367 (N_10367,N_9743,N_9998);
and U10368 (N_10368,N_9768,N_9618);
xor U10369 (N_10369,N_9812,N_9997);
and U10370 (N_10370,N_9958,N_9605);
xnor U10371 (N_10371,N_9859,N_9700);
nand U10372 (N_10372,N_9873,N_9931);
nand U10373 (N_10373,N_9655,N_9799);
xor U10374 (N_10374,N_9616,N_9906);
or U10375 (N_10375,N_9608,N_9860);
xnor U10376 (N_10376,N_9735,N_9682);
xor U10377 (N_10377,N_9774,N_9691);
xor U10378 (N_10378,N_9814,N_9876);
and U10379 (N_10379,N_9643,N_9967);
xor U10380 (N_10380,N_9971,N_9769);
and U10381 (N_10381,N_9652,N_9757);
and U10382 (N_10382,N_9601,N_9830);
nor U10383 (N_10383,N_9719,N_9616);
and U10384 (N_10384,N_9995,N_9741);
or U10385 (N_10385,N_9898,N_9695);
and U10386 (N_10386,N_9886,N_9885);
nor U10387 (N_10387,N_9946,N_9945);
and U10388 (N_10388,N_9764,N_9765);
nor U10389 (N_10389,N_9840,N_9887);
xnor U10390 (N_10390,N_9817,N_9786);
nor U10391 (N_10391,N_9812,N_9835);
nor U10392 (N_10392,N_9982,N_9725);
or U10393 (N_10393,N_9652,N_9995);
nand U10394 (N_10394,N_9917,N_9644);
and U10395 (N_10395,N_9935,N_9860);
xor U10396 (N_10396,N_9841,N_9839);
and U10397 (N_10397,N_9935,N_9813);
or U10398 (N_10398,N_9920,N_9639);
or U10399 (N_10399,N_9939,N_9870);
xor U10400 (N_10400,N_10080,N_10300);
xnor U10401 (N_10401,N_10067,N_10139);
xor U10402 (N_10402,N_10182,N_10278);
nand U10403 (N_10403,N_10190,N_10172);
or U10404 (N_10404,N_10052,N_10030);
nor U10405 (N_10405,N_10089,N_10377);
xnor U10406 (N_10406,N_10072,N_10218);
and U10407 (N_10407,N_10081,N_10101);
nand U10408 (N_10408,N_10287,N_10000);
nor U10409 (N_10409,N_10198,N_10233);
xor U10410 (N_10410,N_10009,N_10196);
nor U10411 (N_10411,N_10303,N_10284);
or U10412 (N_10412,N_10168,N_10290);
and U10413 (N_10413,N_10097,N_10316);
or U10414 (N_10414,N_10350,N_10297);
nor U10415 (N_10415,N_10184,N_10147);
nor U10416 (N_10416,N_10028,N_10324);
or U10417 (N_10417,N_10262,N_10112);
xor U10418 (N_10418,N_10209,N_10063);
or U10419 (N_10419,N_10007,N_10044);
and U10420 (N_10420,N_10326,N_10189);
nor U10421 (N_10421,N_10347,N_10335);
xor U10422 (N_10422,N_10373,N_10006);
or U10423 (N_10423,N_10064,N_10179);
nor U10424 (N_10424,N_10046,N_10259);
or U10425 (N_10425,N_10175,N_10123);
xor U10426 (N_10426,N_10340,N_10034);
or U10427 (N_10427,N_10236,N_10227);
nor U10428 (N_10428,N_10294,N_10301);
nand U10429 (N_10429,N_10231,N_10383);
xor U10430 (N_10430,N_10291,N_10137);
xnor U10431 (N_10431,N_10153,N_10221);
and U10432 (N_10432,N_10048,N_10352);
xor U10433 (N_10433,N_10387,N_10271);
xor U10434 (N_10434,N_10128,N_10166);
or U10435 (N_10435,N_10029,N_10215);
and U10436 (N_10436,N_10167,N_10171);
or U10437 (N_10437,N_10267,N_10117);
nand U10438 (N_10438,N_10041,N_10228);
xnor U10439 (N_10439,N_10155,N_10132);
nand U10440 (N_10440,N_10138,N_10314);
nor U10441 (N_10441,N_10111,N_10275);
nand U10442 (N_10442,N_10238,N_10277);
and U10443 (N_10443,N_10393,N_10254);
or U10444 (N_10444,N_10252,N_10071);
or U10445 (N_10445,N_10346,N_10143);
or U10446 (N_10446,N_10388,N_10016);
nor U10447 (N_10447,N_10160,N_10364);
nand U10448 (N_10448,N_10152,N_10018);
or U10449 (N_10449,N_10251,N_10205);
nand U10450 (N_10450,N_10313,N_10317);
nor U10451 (N_10451,N_10305,N_10157);
xor U10452 (N_10452,N_10075,N_10201);
or U10453 (N_10453,N_10253,N_10362);
and U10454 (N_10454,N_10116,N_10114);
nand U10455 (N_10455,N_10079,N_10154);
or U10456 (N_10456,N_10134,N_10105);
and U10457 (N_10457,N_10107,N_10069);
xor U10458 (N_10458,N_10269,N_10381);
nor U10459 (N_10459,N_10359,N_10035);
or U10460 (N_10460,N_10082,N_10051);
xnor U10461 (N_10461,N_10203,N_10037);
and U10462 (N_10462,N_10242,N_10012);
nand U10463 (N_10463,N_10149,N_10165);
nor U10464 (N_10464,N_10004,N_10309);
nand U10465 (N_10465,N_10308,N_10281);
or U10466 (N_10466,N_10380,N_10087);
or U10467 (N_10467,N_10243,N_10050);
and U10468 (N_10468,N_10136,N_10120);
xor U10469 (N_10469,N_10397,N_10365);
and U10470 (N_10470,N_10022,N_10174);
nor U10471 (N_10471,N_10333,N_10239);
nand U10472 (N_10472,N_10360,N_10031);
nor U10473 (N_10473,N_10357,N_10370);
nor U10474 (N_10474,N_10199,N_10158);
or U10475 (N_10475,N_10255,N_10283);
xnor U10476 (N_10476,N_10096,N_10320);
or U10477 (N_10477,N_10056,N_10059);
or U10478 (N_10478,N_10321,N_10235);
and U10479 (N_10479,N_10003,N_10135);
nor U10480 (N_10480,N_10109,N_10204);
nand U10481 (N_10481,N_10263,N_10306);
xor U10482 (N_10482,N_10224,N_10240);
xor U10483 (N_10483,N_10200,N_10376);
xor U10484 (N_10484,N_10328,N_10285);
xnor U10485 (N_10485,N_10021,N_10040);
or U10486 (N_10486,N_10094,N_10057);
nor U10487 (N_10487,N_10104,N_10348);
and U10488 (N_10488,N_10384,N_10361);
nand U10489 (N_10489,N_10025,N_10342);
nand U10490 (N_10490,N_10173,N_10020);
and U10491 (N_10491,N_10011,N_10344);
or U10492 (N_10492,N_10163,N_10332);
nand U10493 (N_10493,N_10141,N_10245);
and U10494 (N_10494,N_10256,N_10207);
and U10495 (N_10495,N_10077,N_10178);
xnor U10496 (N_10496,N_10142,N_10296);
or U10497 (N_10497,N_10014,N_10232);
nand U10498 (N_10498,N_10001,N_10086);
nor U10499 (N_10499,N_10208,N_10268);
nor U10500 (N_10500,N_10356,N_10090);
and U10501 (N_10501,N_10131,N_10144);
or U10502 (N_10502,N_10118,N_10185);
or U10503 (N_10503,N_10156,N_10358);
or U10504 (N_10504,N_10013,N_10108);
xor U10505 (N_10505,N_10274,N_10330);
nand U10506 (N_10506,N_10076,N_10193);
nand U10507 (N_10507,N_10113,N_10053);
or U10508 (N_10508,N_10394,N_10258);
nor U10509 (N_10509,N_10244,N_10095);
nand U10510 (N_10510,N_10026,N_10270);
nor U10511 (N_10511,N_10150,N_10299);
nor U10512 (N_10512,N_10216,N_10129);
or U10513 (N_10513,N_10148,N_10264);
nand U10514 (N_10514,N_10043,N_10345);
or U10515 (N_10515,N_10382,N_10246);
and U10516 (N_10516,N_10169,N_10125);
nor U10517 (N_10517,N_10307,N_10389);
and U10518 (N_10518,N_10015,N_10042);
xor U10519 (N_10519,N_10372,N_10222);
nand U10520 (N_10520,N_10170,N_10247);
xnor U10521 (N_10521,N_10093,N_10180);
xnor U10522 (N_10522,N_10212,N_10146);
xnor U10523 (N_10523,N_10033,N_10351);
nand U10524 (N_10524,N_10127,N_10337);
nor U10525 (N_10525,N_10186,N_10088);
xor U10526 (N_10526,N_10273,N_10368);
nor U10527 (N_10527,N_10045,N_10391);
and U10528 (N_10528,N_10084,N_10280);
nand U10529 (N_10529,N_10065,N_10323);
and U10530 (N_10530,N_10214,N_10266);
and U10531 (N_10531,N_10140,N_10295);
nand U10532 (N_10532,N_10197,N_10399);
xor U10533 (N_10533,N_10145,N_10126);
or U10534 (N_10534,N_10047,N_10103);
xor U10535 (N_10535,N_10195,N_10331);
xnor U10536 (N_10536,N_10177,N_10100);
xnor U10537 (N_10537,N_10005,N_10036);
nor U10538 (N_10538,N_10371,N_10133);
and U10539 (N_10539,N_10191,N_10312);
or U10540 (N_10540,N_10188,N_10322);
xor U10541 (N_10541,N_10398,N_10343);
xnor U10542 (N_10542,N_10083,N_10265);
xor U10543 (N_10543,N_10392,N_10099);
nor U10544 (N_10544,N_10039,N_10092);
or U10545 (N_10545,N_10319,N_10237);
or U10546 (N_10546,N_10353,N_10363);
nor U10547 (N_10547,N_10032,N_10329);
xor U10548 (N_10548,N_10049,N_10282);
nor U10549 (N_10549,N_10375,N_10257);
xnor U10550 (N_10550,N_10106,N_10260);
xnor U10551 (N_10551,N_10334,N_10002);
xnor U10552 (N_10552,N_10395,N_10181);
or U10553 (N_10553,N_10293,N_10219);
or U10554 (N_10554,N_10085,N_10379);
nor U10555 (N_10555,N_10369,N_10378);
nand U10556 (N_10556,N_10017,N_10302);
or U10557 (N_10557,N_10230,N_10292);
or U10558 (N_10558,N_10192,N_10229);
or U10559 (N_10559,N_10289,N_10070);
xnor U10560 (N_10560,N_10311,N_10024);
nor U10561 (N_10561,N_10038,N_10159);
nor U10562 (N_10562,N_10091,N_10023);
and U10563 (N_10563,N_10286,N_10327);
xor U10564 (N_10564,N_10220,N_10121);
nand U10565 (N_10565,N_10058,N_10130);
xor U10566 (N_10566,N_10396,N_10054);
nor U10567 (N_10567,N_10339,N_10176);
and U10568 (N_10568,N_10060,N_10183);
nand U10569 (N_10569,N_10062,N_10349);
or U10570 (N_10570,N_10122,N_10304);
nand U10571 (N_10571,N_10225,N_10213);
xnor U10572 (N_10572,N_10374,N_10194);
or U10573 (N_10573,N_10336,N_10010);
nand U10574 (N_10574,N_10318,N_10124);
or U10575 (N_10575,N_10367,N_10241);
nand U10576 (N_10576,N_10390,N_10223);
or U10577 (N_10577,N_10310,N_10206);
nand U10578 (N_10578,N_10276,N_10068);
nor U10579 (N_10579,N_10098,N_10073);
nor U10580 (N_10580,N_10074,N_10164);
xor U10581 (N_10581,N_10250,N_10110);
and U10582 (N_10582,N_10078,N_10279);
nor U10583 (N_10583,N_10151,N_10027);
and U10584 (N_10584,N_10019,N_10226);
xor U10585 (N_10585,N_10161,N_10272);
nand U10586 (N_10586,N_10210,N_10261);
and U10587 (N_10587,N_10341,N_10187);
xnor U10588 (N_10588,N_10102,N_10061);
nor U10589 (N_10589,N_10217,N_10288);
and U10590 (N_10590,N_10386,N_10315);
and U10591 (N_10591,N_10325,N_10248);
nand U10592 (N_10592,N_10008,N_10355);
or U10593 (N_10593,N_10211,N_10115);
or U10594 (N_10594,N_10055,N_10234);
xor U10595 (N_10595,N_10119,N_10298);
xnor U10596 (N_10596,N_10066,N_10385);
nand U10597 (N_10597,N_10249,N_10162);
nand U10598 (N_10598,N_10366,N_10338);
nor U10599 (N_10599,N_10202,N_10354);
or U10600 (N_10600,N_10341,N_10015);
nor U10601 (N_10601,N_10245,N_10009);
xnor U10602 (N_10602,N_10209,N_10004);
and U10603 (N_10603,N_10152,N_10379);
xnor U10604 (N_10604,N_10216,N_10192);
and U10605 (N_10605,N_10034,N_10170);
nor U10606 (N_10606,N_10039,N_10267);
xor U10607 (N_10607,N_10113,N_10003);
or U10608 (N_10608,N_10085,N_10303);
xnor U10609 (N_10609,N_10368,N_10215);
or U10610 (N_10610,N_10191,N_10157);
or U10611 (N_10611,N_10136,N_10259);
nand U10612 (N_10612,N_10271,N_10304);
or U10613 (N_10613,N_10295,N_10288);
xnor U10614 (N_10614,N_10145,N_10380);
or U10615 (N_10615,N_10295,N_10197);
and U10616 (N_10616,N_10209,N_10300);
xor U10617 (N_10617,N_10283,N_10293);
or U10618 (N_10618,N_10141,N_10012);
nor U10619 (N_10619,N_10294,N_10061);
and U10620 (N_10620,N_10365,N_10071);
nand U10621 (N_10621,N_10351,N_10318);
and U10622 (N_10622,N_10357,N_10130);
nand U10623 (N_10623,N_10093,N_10007);
and U10624 (N_10624,N_10167,N_10042);
or U10625 (N_10625,N_10217,N_10377);
and U10626 (N_10626,N_10241,N_10256);
or U10627 (N_10627,N_10009,N_10207);
and U10628 (N_10628,N_10020,N_10087);
and U10629 (N_10629,N_10221,N_10040);
or U10630 (N_10630,N_10341,N_10124);
nor U10631 (N_10631,N_10123,N_10189);
nor U10632 (N_10632,N_10325,N_10026);
and U10633 (N_10633,N_10180,N_10222);
and U10634 (N_10634,N_10201,N_10087);
or U10635 (N_10635,N_10346,N_10009);
nor U10636 (N_10636,N_10097,N_10235);
nand U10637 (N_10637,N_10213,N_10341);
nand U10638 (N_10638,N_10035,N_10123);
or U10639 (N_10639,N_10348,N_10158);
nand U10640 (N_10640,N_10179,N_10183);
and U10641 (N_10641,N_10281,N_10278);
or U10642 (N_10642,N_10129,N_10254);
or U10643 (N_10643,N_10025,N_10026);
nand U10644 (N_10644,N_10123,N_10254);
nor U10645 (N_10645,N_10238,N_10272);
and U10646 (N_10646,N_10065,N_10206);
or U10647 (N_10647,N_10189,N_10383);
nand U10648 (N_10648,N_10010,N_10123);
nor U10649 (N_10649,N_10383,N_10089);
nand U10650 (N_10650,N_10039,N_10041);
xnor U10651 (N_10651,N_10207,N_10005);
nor U10652 (N_10652,N_10142,N_10224);
xor U10653 (N_10653,N_10057,N_10055);
nor U10654 (N_10654,N_10034,N_10317);
or U10655 (N_10655,N_10046,N_10044);
and U10656 (N_10656,N_10336,N_10033);
or U10657 (N_10657,N_10119,N_10334);
or U10658 (N_10658,N_10060,N_10240);
and U10659 (N_10659,N_10214,N_10096);
nor U10660 (N_10660,N_10355,N_10003);
nor U10661 (N_10661,N_10032,N_10305);
nand U10662 (N_10662,N_10160,N_10069);
nor U10663 (N_10663,N_10280,N_10087);
and U10664 (N_10664,N_10170,N_10193);
and U10665 (N_10665,N_10172,N_10378);
and U10666 (N_10666,N_10065,N_10225);
xnor U10667 (N_10667,N_10118,N_10347);
nor U10668 (N_10668,N_10088,N_10349);
and U10669 (N_10669,N_10325,N_10039);
nor U10670 (N_10670,N_10150,N_10207);
nor U10671 (N_10671,N_10142,N_10213);
xnor U10672 (N_10672,N_10306,N_10172);
xor U10673 (N_10673,N_10105,N_10077);
xor U10674 (N_10674,N_10041,N_10006);
and U10675 (N_10675,N_10299,N_10240);
or U10676 (N_10676,N_10227,N_10004);
xor U10677 (N_10677,N_10065,N_10060);
nand U10678 (N_10678,N_10124,N_10291);
and U10679 (N_10679,N_10385,N_10171);
xnor U10680 (N_10680,N_10219,N_10377);
nand U10681 (N_10681,N_10350,N_10370);
or U10682 (N_10682,N_10176,N_10079);
and U10683 (N_10683,N_10004,N_10161);
xor U10684 (N_10684,N_10107,N_10146);
xnor U10685 (N_10685,N_10139,N_10077);
or U10686 (N_10686,N_10179,N_10275);
nand U10687 (N_10687,N_10123,N_10156);
and U10688 (N_10688,N_10090,N_10156);
or U10689 (N_10689,N_10152,N_10181);
or U10690 (N_10690,N_10089,N_10229);
nor U10691 (N_10691,N_10023,N_10074);
xnor U10692 (N_10692,N_10294,N_10097);
or U10693 (N_10693,N_10289,N_10311);
nor U10694 (N_10694,N_10285,N_10274);
nand U10695 (N_10695,N_10197,N_10262);
and U10696 (N_10696,N_10065,N_10283);
nor U10697 (N_10697,N_10014,N_10361);
xor U10698 (N_10698,N_10111,N_10186);
or U10699 (N_10699,N_10356,N_10145);
xor U10700 (N_10700,N_10171,N_10235);
and U10701 (N_10701,N_10340,N_10284);
or U10702 (N_10702,N_10123,N_10158);
or U10703 (N_10703,N_10188,N_10303);
and U10704 (N_10704,N_10362,N_10011);
nand U10705 (N_10705,N_10247,N_10114);
xnor U10706 (N_10706,N_10054,N_10125);
xor U10707 (N_10707,N_10124,N_10280);
and U10708 (N_10708,N_10280,N_10020);
and U10709 (N_10709,N_10366,N_10297);
nor U10710 (N_10710,N_10124,N_10335);
nor U10711 (N_10711,N_10137,N_10098);
or U10712 (N_10712,N_10140,N_10391);
nor U10713 (N_10713,N_10073,N_10216);
xnor U10714 (N_10714,N_10123,N_10213);
nand U10715 (N_10715,N_10345,N_10331);
and U10716 (N_10716,N_10319,N_10330);
nand U10717 (N_10717,N_10394,N_10197);
or U10718 (N_10718,N_10380,N_10103);
nor U10719 (N_10719,N_10314,N_10140);
and U10720 (N_10720,N_10338,N_10199);
xor U10721 (N_10721,N_10277,N_10268);
nand U10722 (N_10722,N_10050,N_10267);
nand U10723 (N_10723,N_10379,N_10246);
nand U10724 (N_10724,N_10246,N_10086);
xnor U10725 (N_10725,N_10291,N_10077);
xnor U10726 (N_10726,N_10063,N_10378);
and U10727 (N_10727,N_10047,N_10237);
or U10728 (N_10728,N_10072,N_10252);
nand U10729 (N_10729,N_10161,N_10253);
or U10730 (N_10730,N_10084,N_10041);
xnor U10731 (N_10731,N_10092,N_10169);
nand U10732 (N_10732,N_10082,N_10360);
and U10733 (N_10733,N_10015,N_10040);
or U10734 (N_10734,N_10172,N_10309);
nand U10735 (N_10735,N_10136,N_10258);
nor U10736 (N_10736,N_10315,N_10364);
nand U10737 (N_10737,N_10038,N_10091);
nand U10738 (N_10738,N_10340,N_10165);
and U10739 (N_10739,N_10383,N_10396);
and U10740 (N_10740,N_10108,N_10074);
xor U10741 (N_10741,N_10117,N_10020);
xnor U10742 (N_10742,N_10323,N_10389);
or U10743 (N_10743,N_10052,N_10373);
and U10744 (N_10744,N_10367,N_10107);
xor U10745 (N_10745,N_10312,N_10217);
and U10746 (N_10746,N_10141,N_10365);
xnor U10747 (N_10747,N_10138,N_10100);
nor U10748 (N_10748,N_10286,N_10058);
and U10749 (N_10749,N_10379,N_10201);
xor U10750 (N_10750,N_10207,N_10017);
or U10751 (N_10751,N_10117,N_10256);
nand U10752 (N_10752,N_10133,N_10248);
and U10753 (N_10753,N_10214,N_10222);
nand U10754 (N_10754,N_10316,N_10108);
xor U10755 (N_10755,N_10192,N_10235);
nor U10756 (N_10756,N_10390,N_10271);
and U10757 (N_10757,N_10331,N_10051);
xnor U10758 (N_10758,N_10309,N_10174);
nor U10759 (N_10759,N_10057,N_10225);
xnor U10760 (N_10760,N_10018,N_10110);
nand U10761 (N_10761,N_10189,N_10355);
or U10762 (N_10762,N_10371,N_10119);
or U10763 (N_10763,N_10276,N_10298);
or U10764 (N_10764,N_10259,N_10010);
or U10765 (N_10765,N_10187,N_10134);
or U10766 (N_10766,N_10366,N_10313);
nand U10767 (N_10767,N_10056,N_10183);
nor U10768 (N_10768,N_10326,N_10387);
nor U10769 (N_10769,N_10302,N_10201);
nand U10770 (N_10770,N_10371,N_10312);
nand U10771 (N_10771,N_10304,N_10121);
xor U10772 (N_10772,N_10183,N_10340);
and U10773 (N_10773,N_10297,N_10282);
xor U10774 (N_10774,N_10369,N_10181);
and U10775 (N_10775,N_10110,N_10003);
xor U10776 (N_10776,N_10065,N_10024);
xnor U10777 (N_10777,N_10336,N_10250);
and U10778 (N_10778,N_10156,N_10227);
or U10779 (N_10779,N_10018,N_10209);
nand U10780 (N_10780,N_10310,N_10287);
nand U10781 (N_10781,N_10390,N_10161);
nor U10782 (N_10782,N_10000,N_10076);
xnor U10783 (N_10783,N_10197,N_10204);
or U10784 (N_10784,N_10120,N_10391);
xor U10785 (N_10785,N_10125,N_10136);
nor U10786 (N_10786,N_10316,N_10293);
xnor U10787 (N_10787,N_10364,N_10288);
and U10788 (N_10788,N_10160,N_10108);
nand U10789 (N_10789,N_10038,N_10191);
xor U10790 (N_10790,N_10033,N_10207);
nand U10791 (N_10791,N_10011,N_10130);
or U10792 (N_10792,N_10321,N_10037);
xnor U10793 (N_10793,N_10293,N_10339);
or U10794 (N_10794,N_10231,N_10155);
xnor U10795 (N_10795,N_10035,N_10259);
xnor U10796 (N_10796,N_10149,N_10131);
xor U10797 (N_10797,N_10089,N_10197);
nand U10798 (N_10798,N_10052,N_10240);
xor U10799 (N_10799,N_10135,N_10318);
and U10800 (N_10800,N_10759,N_10663);
nand U10801 (N_10801,N_10538,N_10769);
and U10802 (N_10802,N_10442,N_10683);
nand U10803 (N_10803,N_10501,N_10526);
nor U10804 (N_10804,N_10672,N_10601);
nor U10805 (N_10805,N_10569,N_10778);
nor U10806 (N_10806,N_10704,N_10647);
nand U10807 (N_10807,N_10689,N_10434);
and U10808 (N_10808,N_10564,N_10447);
xnor U10809 (N_10809,N_10755,N_10636);
xor U10810 (N_10810,N_10504,N_10761);
and U10811 (N_10811,N_10468,N_10618);
and U10812 (N_10812,N_10760,N_10664);
xor U10813 (N_10813,N_10763,N_10791);
and U10814 (N_10814,N_10448,N_10550);
nor U10815 (N_10815,N_10716,N_10457);
or U10816 (N_10816,N_10431,N_10451);
or U10817 (N_10817,N_10418,N_10466);
and U10818 (N_10818,N_10687,N_10721);
nor U10819 (N_10819,N_10630,N_10532);
or U10820 (N_10820,N_10509,N_10789);
nor U10821 (N_10821,N_10407,N_10596);
or U10822 (N_10822,N_10472,N_10606);
or U10823 (N_10823,N_10503,N_10638);
nand U10824 (N_10824,N_10793,N_10548);
and U10825 (N_10825,N_10456,N_10698);
nand U10826 (N_10826,N_10561,N_10541);
nand U10827 (N_10827,N_10489,N_10792);
xor U10828 (N_10828,N_10681,N_10747);
nor U10829 (N_10829,N_10494,N_10549);
nor U10830 (N_10830,N_10637,N_10745);
and U10831 (N_10831,N_10514,N_10496);
nor U10832 (N_10832,N_10517,N_10610);
nor U10833 (N_10833,N_10487,N_10720);
or U10834 (N_10834,N_10593,N_10677);
or U10835 (N_10835,N_10400,N_10497);
nor U10836 (N_10836,N_10483,N_10575);
nand U10837 (N_10837,N_10511,N_10612);
or U10838 (N_10838,N_10770,N_10626);
xnor U10839 (N_10839,N_10507,N_10686);
and U10840 (N_10840,N_10600,N_10421);
or U10841 (N_10841,N_10658,N_10542);
nand U10842 (N_10842,N_10777,N_10665);
nor U10843 (N_10843,N_10765,N_10555);
and U10844 (N_10844,N_10422,N_10408);
and U10845 (N_10845,N_10639,N_10694);
and U10846 (N_10846,N_10751,N_10752);
and U10847 (N_10847,N_10565,N_10558);
xnor U10848 (N_10848,N_10474,N_10490);
or U10849 (N_10849,N_10591,N_10557);
nor U10850 (N_10850,N_10404,N_10732);
and U10851 (N_10851,N_10736,N_10411);
xnor U10852 (N_10852,N_10520,N_10657);
nand U10853 (N_10853,N_10633,N_10594);
nor U10854 (N_10854,N_10534,N_10644);
nand U10855 (N_10855,N_10785,N_10790);
nor U10856 (N_10856,N_10676,N_10794);
xor U10857 (N_10857,N_10592,N_10443);
or U10858 (N_10858,N_10423,N_10729);
nor U10859 (N_10859,N_10481,N_10695);
and U10860 (N_10860,N_10462,N_10512);
and U10861 (N_10861,N_10605,N_10525);
nand U10862 (N_10862,N_10762,N_10484);
xor U10863 (N_10863,N_10797,N_10631);
xor U10864 (N_10864,N_10754,N_10660);
xnor U10865 (N_10865,N_10486,N_10653);
xor U10866 (N_10866,N_10479,N_10623);
xor U10867 (N_10867,N_10563,N_10670);
xnor U10868 (N_10868,N_10620,N_10455);
xnor U10869 (N_10869,N_10554,N_10572);
nand U10870 (N_10870,N_10774,N_10533);
nor U10871 (N_10871,N_10654,N_10491);
nor U10872 (N_10872,N_10570,N_10562);
and U10873 (N_10873,N_10559,N_10666);
or U10874 (N_10874,N_10444,N_10615);
and U10875 (N_10875,N_10750,N_10599);
nand U10876 (N_10876,N_10645,N_10693);
or U10877 (N_10877,N_10413,N_10619);
nor U10878 (N_10878,N_10604,N_10682);
or U10879 (N_10879,N_10656,N_10627);
or U10880 (N_10880,N_10467,N_10705);
and U10881 (N_10881,N_10401,N_10624);
or U10882 (N_10882,N_10417,N_10643);
and U10883 (N_10883,N_10579,N_10427);
xor U10884 (N_10884,N_10724,N_10632);
nor U10885 (N_10885,N_10758,N_10518);
nand U10886 (N_10886,N_10781,N_10609);
and U10887 (N_10887,N_10582,N_10586);
nor U10888 (N_10888,N_10524,N_10416);
and U10889 (N_10889,N_10535,N_10515);
nor U10890 (N_10890,N_10607,N_10674);
and U10891 (N_10891,N_10784,N_10488);
and U10892 (N_10892,N_10419,N_10722);
nor U10893 (N_10893,N_10767,N_10414);
and U10894 (N_10894,N_10473,N_10587);
nand U10895 (N_10895,N_10679,N_10475);
or U10896 (N_10896,N_10588,N_10782);
nor U10897 (N_10897,N_10478,N_10734);
or U10898 (N_10898,N_10748,N_10611);
nand U10899 (N_10899,N_10715,N_10780);
nor U10900 (N_10900,N_10669,N_10634);
nand U10901 (N_10901,N_10614,N_10420);
nor U10902 (N_10902,N_10690,N_10508);
and U10903 (N_10903,N_10405,N_10471);
and U10904 (N_10904,N_10652,N_10498);
xnor U10905 (N_10905,N_10493,N_10712);
and U10906 (N_10906,N_10566,N_10437);
xor U10907 (N_10907,N_10616,N_10661);
and U10908 (N_10908,N_10551,N_10523);
xnor U10909 (N_10909,N_10540,N_10560);
xnor U10910 (N_10910,N_10465,N_10766);
and U10911 (N_10911,N_10463,N_10458);
nand U10912 (N_10912,N_10460,N_10703);
xor U10913 (N_10913,N_10459,N_10415);
xnor U10914 (N_10914,N_10642,N_10406);
nand U10915 (N_10915,N_10519,N_10678);
nand U10916 (N_10916,N_10753,N_10505);
xnor U10917 (N_10917,N_10675,N_10454);
xnor U10918 (N_10918,N_10556,N_10544);
xor U10919 (N_10919,N_10739,N_10700);
or U10920 (N_10920,N_10684,N_10757);
nand U10921 (N_10921,N_10441,N_10726);
and U10922 (N_10922,N_10590,N_10725);
and U10923 (N_10923,N_10659,N_10673);
xor U10924 (N_10924,N_10527,N_10480);
and U10925 (N_10925,N_10640,N_10603);
or U10926 (N_10926,N_10680,N_10744);
xnor U10927 (N_10927,N_10410,N_10438);
nor U10928 (N_10928,N_10702,N_10799);
nor U10929 (N_10929,N_10688,N_10409);
and U10930 (N_10930,N_10783,N_10585);
or U10931 (N_10931,N_10798,N_10733);
and U10932 (N_10932,N_10506,N_10452);
nor U10933 (N_10933,N_10552,N_10502);
xnor U10934 (N_10934,N_10696,N_10731);
or U10935 (N_10935,N_10589,N_10461);
xor U10936 (N_10936,N_10646,N_10613);
nor U10937 (N_10937,N_10635,N_10573);
or U10938 (N_10938,N_10433,N_10628);
and U10939 (N_10939,N_10795,N_10788);
nand U10940 (N_10940,N_10553,N_10771);
nand U10941 (N_10941,N_10701,N_10727);
and U10942 (N_10942,N_10692,N_10741);
nand U10943 (N_10943,N_10697,N_10671);
nor U10944 (N_10944,N_10598,N_10709);
nand U10945 (N_10945,N_10629,N_10436);
nand U10946 (N_10946,N_10685,N_10723);
nor U10947 (N_10947,N_10691,N_10429);
nor U10948 (N_10948,N_10500,N_10786);
xor U10949 (N_10949,N_10470,N_10521);
or U10950 (N_10950,N_10730,N_10776);
xnor U10951 (N_10951,N_10516,N_10648);
or U10952 (N_10952,N_10655,N_10428);
nand U10953 (N_10953,N_10580,N_10649);
nor U10954 (N_10954,N_10710,N_10536);
or U10955 (N_10955,N_10522,N_10787);
nand U10956 (N_10956,N_10583,N_10531);
nor U10957 (N_10957,N_10749,N_10738);
nand U10958 (N_10958,N_10768,N_10584);
nand U10959 (N_10959,N_10699,N_10432);
nand U10960 (N_10960,N_10425,N_10568);
and U10961 (N_10961,N_10773,N_10424);
and U10962 (N_10962,N_10426,N_10597);
nand U10963 (N_10963,N_10641,N_10707);
nor U10964 (N_10964,N_10485,N_10439);
nor U10965 (N_10965,N_10625,N_10719);
and U10966 (N_10966,N_10528,N_10430);
xor U10967 (N_10967,N_10403,N_10576);
nor U10968 (N_10968,N_10543,N_10714);
xor U10969 (N_10969,N_10450,N_10706);
nand U10970 (N_10970,N_10440,N_10622);
and U10971 (N_10971,N_10482,N_10510);
nor U10972 (N_10972,N_10621,N_10530);
nor U10973 (N_10973,N_10718,N_10469);
or U10974 (N_10974,N_10595,N_10708);
nand U10975 (N_10975,N_10537,N_10435);
nor U10976 (N_10976,N_10711,N_10402);
and U10977 (N_10977,N_10713,N_10651);
nand U10978 (N_10978,N_10464,N_10662);
and U10979 (N_10979,N_10667,N_10717);
xor U10980 (N_10980,N_10668,N_10574);
nand U10981 (N_10981,N_10779,N_10449);
and U10982 (N_10982,N_10476,N_10772);
or U10983 (N_10983,N_10577,N_10539);
xor U10984 (N_10984,N_10775,N_10546);
nor U10985 (N_10985,N_10578,N_10495);
xnor U10986 (N_10986,N_10453,N_10617);
and U10987 (N_10987,N_10547,N_10735);
xor U10988 (N_10988,N_10743,N_10608);
nand U10989 (N_10989,N_10412,N_10545);
nor U10990 (N_10990,N_10740,N_10737);
and U10991 (N_10991,N_10746,N_10796);
xor U10992 (N_10992,N_10571,N_10445);
nand U10993 (N_10993,N_10513,N_10446);
nand U10994 (N_10994,N_10529,N_10742);
xnor U10995 (N_10995,N_10728,N_10764);
nor U10996 (N_10996,N_10499,N_10756);
and U10997 (N_10997,N_10492,N_10477);
or U10998 (N_10998,N_10567,N_10602);
or U10999 (N_10999,N_10581,N_10650);
xnor U11000 (N_11000,N_10702,N_10600);
nor U11001 (N_11001,N_10615,N_10759);
xnor U11002 (N_11002,N_10679,N_10656);
nand U11003 (N_11003,N_10723,N_10494);
or U11004 (N_11004,N_10715,N_10570);
xor U11005 (N_11005,N_10601,N_10590);
or U11006 (N_11006,N_10497,N_10647);
nand U11007 (N_11007,N_10749,N_10572);
nor U11008 (N_11008,N_10608,N_10647);
nor U11009 (N_11009,N_10703,N_10554);
nor U11010 (N_11010,N_10515,N_10676);
and U11011 (N_11011,N_10492,N_10720);
xnor U11012 (N_11012,N_10721,N_10650);
nor U11013 (N_11013,N_10697,N_10483);
nand U11014 (N_11014,N_10583,N_10446);
nand U11015 (N_11015,N_10669,N_10601);
or U11016 (N_11016,N_10753,N_10771);
or U11017 (N_11017,N_10763,N_10619);
nand U11018 (N_11018,N_10737,N_10709);
xor U11019 (N_11019,N_10697,N_10578);
and U11020 (N_11020,N_10453,N_10573);
and U11021 (N_11021,N_10655,N_10589);
nor U11022 (N_11022,N_10680,N_10738);
nor U11023 (N_11023,N_10674,N_10707);
and U11024 (N_11024,N_10451,N_10582);
and U11025 (N_11025,N_10793,N_10438);
nor U11026 (N_11026,N_10560,N_10791);
nand U11027 (N_11027,N_10447,N_10646);
nor U11028 (N_11028,N_10481,N_10754);
nand U11029 (N_11029,N_10590,N_10406);
nand U11030 (N_11030,N_10466,N_10437);
and U11031 (N_11031,N_10425,N_10551);
xnor U11032 (N_11032,N_10504,N_10690);
or U11033 (N_11033,N_10612,N_10403);
xnor U11034 (N_11034,N_10523,N_10634);
or U11035 (N_11035,N_10557,N_10542);
or U11036 (N_11036,N_10610,N_10731);
nor U11037 (N_11037,N_10439,N_10759);
nand U11038 (N_11038,N_10416,N_10564);
xnor U11039 (N_11039,N_10640,N_10455);
xnor U11040 (N_11040,N_10603,N_10509);
xnor U11041 (N_11041,N_10724,N_10519);
or U11042 (N_11042,N_10683,N_10490);
or U11043 (N_11043,N_10534,N_10499);
and U11044 (N_11044,N_10695,N_10644);
xor U11045 (N_11045,N_10697,N_10541);
xnor U11046 (N_11046,N_10752,N_10544);
or U11047 (N_11047,N_10597,N_10669);
and U11048 (N_11048,N_10627,N_10541);
and U11049 (N_11049,N_10714,N_10623);
or U11050 (N_11050,N_10707,N_10485);
and U11051 (N_11051,N_10564,N_10747);
or U11052 (N_11052,N_10770,N_10783);
or U11053 (N_11053,N_10406,N_10614);
and U11054 (N_11054,N_10487,N_10633);
nand U11055 (N_11055,N_10495,N_10463);
or U11056 (N_11056,N_10776,N_10795);
or U11057 (N_11057,N_10434,N_10574);
or U11058 (N_11058,N_10614,N_10422);
nor U11059 (N_11059,N_10490,N_10647);
and U11060 (N_11060,N_10664,N_10745);
nand U11061 (N_11061,N_10712,N_10443);
nor U11062 (N_11062,N_10572,N_10614);
xor U11063 (N_11063,N_10579,N_10671);
xnor U11064 (N_11064,N_10463,N_10707);
or U11065 (N_11065,N_10518,N_10619);
or U11066 (N_11066,N_10760,N_10530);
and U11067 (N_11067,N_10474,N_10735);
xnor U11068 (N_11068,N_10641,N_10589);
nor U11069 (N_11069,N_10493,N_10415);
nand U11070 (N_11070,N_10480,N_10759);
xnor U11071 (N_11071,N_10761,N_10631);
nor U11072 (N_11072,N_10617,N_10587);
xor U11073 (N_11073,N_10614,N_10595);
nand U11074 (N_11074,N_10694,N_10699);
and U11075 (N_11075,N_10441,N_10631);
and U11076 (N_11076,N_10650,N_10488);
or U11077 (N_11077,N_10768,N_10562);
or U11078 (N_11078,N_10571,N_10781);
xor U11079 (N_11079,N_10697,N_10762);
xnor U11080 (N_11080,N_10567,N_10425);
or U11081 (N_11081,N_10526,N_10449);
nand U11082 (N_11082,N_10635,N_10550);
xnor U11083 (N_11083,N_10487,N_10779);
nor U11084 (N_11084,N_10684,N_10532);
xor U11085 (N_11085,N_10452,N_10536);
and U11086 (N_11086,N_10634,N_10420);
and U11087 (N_11087,N_10537,N_10568);
xor U11088 (N_11088,N_10410,N_10717);
or U11089 (N_11089,N_10430,N_10563);
xnor U11090 (N_11090,N_10496,N_10726);
nand U11091 (N_11091,N_10618,N_10760);
xor U11092 (N_11092,N_10484,N_10768);
xnor U11093 (N_11093,N_10456,N_10448);
nand U11094 (N_11094,N_10537,N_10530);
xor U11095 (N_11095,N_10400,N_10414);
nor U11096 (N_11096,N_10487,N_10739);
and U11097 (N_11097,N_10734,N_10721);
xnor U11098 (N_11098,N_10410,N_10668);
and U11099 (N_11099,N_10701,N_10403);
nand U11100 (N_11100,N_10778,N_10760);
nand U11101 (N_11101,N_10580,N_10421);
xor U11102 (N_11102,N_10691,N_10795);
or U11103 (N_11103,N_10795,N_10796);
xnor U11104 (N_11104,N_10706,N_10447);
xor U11105 (N_11105,N_10585,N_10503);
xor U11106 (N_11106,N_10465,N_10712);
nand U11107 (N_11107,N_10567,N_10661);
and U11108 (N_11108,N_10449,N_10619);
nor U11109 (N_11109,N_10424,N_10575);
nand U11110 (N_11110,N_10558,N_10528);
xor U11111 (N_11111,N_10536,N_10438);
nand U11112 (N_11112,N_10706,N_10762);
and U11113 (N_11113,N_10400,N_10644);
xor U11114 (N_11114,N_10773,N_10796);
or U11115 (N_11115,N_10729,N_10409);
nand U11116 (N_11116,N_10514,N_10638);
and U11117 (N_11117,N_10516,N_10652);
xor U11118 (N_11118,N_10652,N_10648);
and U11119 (N_11119,N_10520,N_10491);
nand U11120 (N_11120,N_10667,N_10453);
xnor U11121 (N_11121,N_10702,N_10620);
nor U11122 (N_11122,N_10671,N_10456);
xnor U11123 (N_11123,N_10641,N_10762);
nor U11124 (N_11124,N_10538,N_10441);
and U11125 (N_11125,N_10779,N_10684);
and U11126 (N_11126,N_10582,N_10660);
xor U11127 (N_11127,N_10703,N_10706);
or U11128 (N_11128,N_10642,N_10465);
nor U11129 (N_11129,N_10760,N_10687);
nor U11130 (N_11130,N_10439,N_10631);
xnor U11131 (N_11131,N_10678,N_10501);
xor U11132 (N_11132,N_10570,N_10596);
or U11133 (N_11133,N_10798,N_10440);
xnor U11134 (N_11134,N_10766,N_10537);
nor U11135 (N_11135,N_10719,N_10451);
nor U11136 (N_11136,N_10775,N_10740);
and U11137 (N_11137,N_10563,N_10706);
nand U11138 (N_11138,N_10591,N_10480);
and U11139 (N_11139,N_10677,N_10751);
nor U11140 (N_11140,N_10670,N_10799);
xnor U11141 (N_11141,N_10502,N_10585);
xor U11142 (N_11142,N_10541,N_10542);
nor U11143 (N_11143,N_10716,N_10580);
and U11144 (N_11144,N_10682,N_10537);
nor U11145 (N_11145,N_10649,N_10746);
and U11146 (N_11146,N_10648,N_10418);
nor U11147 (N_11147,N_10726,N_10425);
nor U11148 (N_11148,N_10676,N_10411);
nor U11149 (N_11149,N_10664,N_10539);
nor U11150 (N_11150,N_10474,N_10574);
nor U11151 (N_11151,N_10759,N_10419);
nand U11152 (N_11152,N_10674,N_10465);
nor U11153 (N_11153,N_10711,N_10689);
or U11154 (N_11154,N_10790,N_10539);
or U11155 (N_11155,N_10440,N_10644);
nand U11156 (N_11156,N_10615,N_10640);
xnor U11157 (N_11157,N_10400,N_10598);
or U11158 (N_11158,N_10777,N_10581);
nand U11159 (N_11159,N_10731,N_10549);
nor U11160 (N_11160,N_10481,N_10589);
xnor U11161 (N_11161,N_10500,N_10677);
nand U11162 (N_11162,N_10698,N_10679);
xnor U11163 (N_11163,N_10682,N_10649);
xnor U11164 (N_11164,N_10492,N_10601);
or U11165 (N_11165,N_10493,N_10717);
nand U11166 (N_11166,N_10422,N_10477);
and U11167 (N_11167,N_10729,N_10622);
nand U11168 (N_11168,N_10435,N_10711);
and U11169 (N_11169,N_10456,N_10650);
nor U11170 (N_11170,N_10515,N_10678);
or U11171 (N_11171,N_10612,N_10716);
and U11172 (N_11172,N_10768,N_10580);
and U11173 (N_11173,N_10423,N_10570);
and U11174 (N_11174,N_10405,N_10768);
and U11175 (N_11175,N_10630,N_10540);
and U11176 (N_11176,N_10611,N_10618);
nor U11177 (N_11177,N_10597,N_10536);
and U11178 (N_11178,N_10490,N_10420);
or U11179 (N_11179,N_10463,N_10423);
or U11180 (N_11180,N_10723,N_10769);
or U11181 (N_11181,N_10575,N_10619);
and U11182 (N_11182,N_10495,N_10749);
or U11183 (N_11183,N_10443,N_10651);
and U11184 (N_11184,N_10696,N_10458);
xor U11185 (N_11185,N_10684,N_10623);
nor U11186 (N_11186,N_10602,N_10784);
nand U11187 (N_11187,N_10659,N_10724);
and U11188 (N_11188,N_10679,N_10524);
and U11189 (N_11189,N_10789,N_10493);
nor U11190 (N_11190,N_10709,N_10643);
and U11191 (N_11191,N_10538,N_10703);
nor U11192 (N_11192,N_10798,N_10794);
nor U11193 (N_11193,N_10577,N_10707);
and U11194 (N_11194,N_10767,N_10615);
and U11195 (N_11195,N_10628,N_10659);
nand U11196 (N_11196,N_10632,N_10720);
xnor U11197 (N_11197,N_10554,N_10437);
xor U11198 (N_11198,N_10486,N_10638);
nand U11199 (N_11199,N_10432,N_10561);
nand U11200 (N_11200,N_10903,N_10919);
and U11201 (N_11201,N_10810,N_11036);
nand U11202 (N_11202,N_10920,N_11140);
nor U11203 (N_11203,N_11138,N_11197);
or U11204 (N_11204,N_10902,N_11075);
nor U11205 (N_11205,N_10884,N_11032);
or U11206 (N_11206,N_11184,N_10921);
nand U11207 (N_11207,N_11183,N_11050);
or U11208 (N_11208,N_10971,N_11073);
nand U11209 (N_11209,N_10930,N_10857);
nor U11210 (N_11210,N_10897,N_10898);
nor U11211 (N_11211,N_10937,N_11131);
or U11212 (N_11212,N_11026,N_10832);
nor U11213 (N_11213,N_10833,N_10865);
nor U11214 (N_11214,N_11024,N_10992);
and U11215 (N_11215,N_10942,N_11031);
xnor U11216 (N_11216,N_10945,N_11079);
or U11217 (N_11217,N_10831,N_10905);
and U11218 (N_11218,N_11002,N_11025);
or U11219 (N_11219,N_10841,N_10870);
nand U11220 (N_11220,N_11174,N_11055);
nand U11221 (N_11221,N_11132,N_11185);
and U11222 (N_11222,N_10805,N_10838);
nand U11223 (N_11223,N_10852,N_10887);
xor U11224 (N_11224,N_11192,N_10860);
nor U11225 (N_11225,N_10856,N_11144);
or U11226 (N_11226,N_11124,N_10961);
xnor U11227 (N_11227,N_11083,N_11013);
or U11228 (N_11228,N_10806,N_10990);
nor U11229 (N_11229,N_10951,N_10842);
and U11230 (N_11230,N_11118,N_11194);
xnor U11231 (N_11231,N_11141,N_11097);
xor U11232 (N_11232,N_11170,N_10809);
or U11233 (N_11233,N_11049,N_11051);
or U11234 (N_11234,N_10802,N_11136);
xor U11235 (N_11235,N_10888,N_11101);
nand U11236 (N_11236,N_10949,N_11180);
nor U11237 (N_11237,N_11146,N_11047);
or U11238 (N_11238,N_10984,N_10918);
nor U11239 (N_11239,N_10892,N_10877);
nor U11240 (N_11240,N_10952,N_10871);
nand U11241 (N_11241,N_11195,N_10824);
xnor U11242 (N_11242,N_10851,N_10943);
and U11243 (N_11243,N_10886,N_11166);
nand U11244 (N_11244,N_11151,N_11048);
nand U11245 (N_11245,N_11057,N_11092);
nor U11246 (N_11246,N_11099,N_10885);
nand U11247 (N_11247,N_11125,N_11068);
and U11248 (N_11248,N_11107,N_11177);
and U11249 (N_11249,N_11155,N_11030);
and U11250 (N_11250,N_10813,N_10853);
and U11251 (N_11251,N_10959,N_11081);
or U11252 (N_11252,N_10933,N_10932);
nand U11253 (N_11253,N_11196,N_10991);
nor U11254 (N_11254,N_10967,N_10958);
xnor U11255 (N_11255,N_10963,N_10881);
xnor U11256 (N_11256,N_11028,N_10934);
xnor U11257 (N_11257,N_11113,N_10988);
nand U11258 (N_11258,N_11006,N_11104);
and U11259 (N_11259,N_10849,N_10972);
or U11260 (N_11260,N_10906,N_11128);
nand U11261 (N_11261,N_10976,N_11114);
or U11262 (N_11262,N_11149,N_11089);
xor U11263 (N_11263,N_10830,N_10968);
xor U11264 (N_11264,N_10873,N_11198);
xnor U11265 (N_11265,N_11112,N_10985);
nor U11266 (N_11266,N_11018,N_11066);
and U11267 (N_11267,N_11193,N_10820);
and U11268 (N_11268,N_10896,N_11163);
and U11269 (N_11269,N_10875,N_11148);
nor U11270 (N_11270,N_11115,N_10823);
nor U11271 (N_11271,N_11060,N_11065);
or U11272 (N_11272,N_11181,N_10995);
nand U11273 (N_11273,N_10863,N_11012);
xor U11274 (N_11274,N_11077,N_10844);
xor U11275 (N_11275,N_11017,N_11190);
xnor U11276 (N_11276,N_11009,N_10843);
nor U11277 (N_11277,N_11103,N_11142);
nor U11278 (N_11278,N_10862,N_10814);
or U11279 (N_11279,N_11072,N_10821);
nor U11280 (N_11280,N_11059,N_11035);
nor U11281 (N_11281,N_10882,N_10822);
nor U11282 (N_11282,N_11110,N_10941);
nand U11283 (N_11283,N_11127,N_11123);
or U11284 (N_11284,N_11062,N_10987);
nand U11285 (N_11285,N_10954,N_11011);
and U11286 (N_11286,N_10812,N_11045);
nor U11287 (N_11287,N_10962,N_10931);
and U11288 (N_11288,N_10986,N_11167);
xor U11289 (N_11289,N_11046,N_10926);
and U11290 (N_11290,N_10974,N_11119);
xnor U11291 (N_11291,N_11179,N_10913);
nand U11292 (N_11292,N_11095,N_10893);
and U11293 (N_11293,N_11150,N_10876);
or U11294 (N_11294,N_10929,N_10953);
or U11295 (N_11295,N_10911,N_10878);
xor U11296 (N_11296,N_11037,N_11082);
nand U11297 (N_11297,N_10835,N_10904);
xor U11298 (N_11298,N_10804,N_11000);
xor U11299 (N_11299,N_11085,N_11019);
nand U11300 (N_11300,N_11008,N_10845);
nor U11301 (N_11301,N_10922,N_11105);
and U11302 (N_11302,N_10816,N_10955);
nor U11303 (N_11303,N_10997,N_10939);
nand U11304 (N_11304,N_10989,N_11109);
nor U11305 (N_11305,N_11084,N_11005);
or U11306 (N_11306,N_10828,N_10975);
and U11307 (N_11307,N_10983,N_10811);
xor U11308 (N_11308,N_11122,N_10827);
nand U11309 (N_11309,N_11106,N_11076);
xor U11310 (N_11310,N_11086,N_10998);
or U11311 (N_11311,N_11022,N_11001);
and U11312 (N_11312,N_10969,N_10917);
nor U11313 (N_11313,N_11038,N_10839);
nand U11314 (N_11314,N_11069,N_10973);
and U11315 (N_11315,N_11171,N_10928);
or U11316 (N_11316,N_11121,N_10848);
nor U11317 (N_11317,N_10915,N_11043);
or U11318 (N_11318,N_11165,N_10817);
xor U11319 (N_11319,N_11040,N_11056);
or U11320 (N_11320,N_10996,N_11015);
nand U11321 (N_11321,N_11090,N_11116);
and U11322 (N_11322,N_11172,N_10825);
and U11323 (N_11323,N_10891,N_11133);
or U11324 (N_11324,N_11029,N_11058);
nand U11325 (N_11325,N_11088,N_11159);
nor U11326 (N_11326,N_11186,N_10808);
nor U11327 (N_11327,N_10979,N_10889);
nand U11328 (N_11328,N_10840,N_10899);
xor U11329 (N_11329,N_10826,N_11199);
xnor U11330 (N_11330,N_10994,N_11158);
xor U11331 (N_11331,N_11129,N_10855);
and U11332 (N_11332,N_10815,N_11041);
nor U11333 (N_11333,N_10850,N_11096);
or U11334 (N_11334,N_10940,N_11143);
or U11335 (N_11335,N_11070,N_11023);
or U11336 (N_11336,N_11137,N_11126);
or U11337 (N_11337,N_10901,N_11188);
nor U11338 (N_11338,N_10819,N_11016);
and U11339 (N_11339,N_10868,N_10982);
or U11340 (N_11340,N_10960,N_10859);
nor U11341 (N_11341,N_10880,N_11111);
or U11342 (N_11342,N_10883,N_10947);
nor U11343 (N_11343,N_10935,N_11074);
or U11344 (N_11344,N_10908,N_11087);
nand U11345 (N_11345,N_10803,N_11169);
nand U11346 (N_11346,N_10890,N_10924);
nand U11347 (N_11347,N_11153,N_10944);
nand U11348 (N_11348,N_11027,N_11100);
nor U11349 (N_11349,N_11175,N_11007);
nand U11350 (N_11350,N_10956,N_10801);
and U11351 (N_11351,N_10981,N_11162);
nand U11352 (N_11352,N_10866,N_10869);
nor U11353 (N_11353,N_11093,N_11152);
nand U11354 (N_11354,N_10957,N_11071);
nor U11355 (N_11355,N_10927,N_11053);
nand U11356 (N_11356,N_11154,N_11067);
xnor U11357 (N_11357,N_11063,N_10864);
and U11358 (N_11358,N_10894,N_10909);
or U11359 (N_11359,N_11134,N_10895);
nor U11360 (N_11360,N_10948,N_11034);
nand U11361 (N_11361,N_11120,N_11052);
or U11362 (N_11362,N_11020,N_10916);
xor U11363 (N_11363,N_11091,N_10836);
xor U11364 (N_11364,N_11078,N_11094);
nor U11365 (N_11365,N_11098,N_10999);
or U11366 (N_11366,N_10818,N_10837);
and U11367 (N_11367,N_11156,N_11168);
nand U11368 (N_11368,N_10936,N_10800);
and U11369 (N_11369,N_11108,N_10874);
nor U11370 (N_11370,N_10993,N_10970);
and U11371 (N_11371,N_11182,N_10861);
nor U11372 (N_11372,N_11164,N_10914);
nor U11373 (N_11373,N_10807,N_11191);
or U11374 (N_11374,N_11102,N_10854);
nand U11375 (N_11375,N_10964,N_10965);
and U11376 (N_11376,N_10977,N_11061);
nor U11377 (N_11377,N_11139,N_11157);
or U11378 (N_11378,N_11042,N_11178);
or U11379 (N_11379,N_10925,N_11189);
xnor U11380 (N_11380,N_11080,N_11033);
xor U11381 (N_11381,N_10879,N_11173);
nor U11382 (N_11382,N_11160,N_11064);
and U11383 (N_11383,N_11004,N_11014);
nor U11384 (N_11384,N_11117,N_11010);
nor U11385 (N_11385,N_10858,N_10867);
nand U11386 (N_11386,N_10912,N_10846);
nand U11387 (N_11387,N_10978,N_11135);
and U11388 (N_11388,N_10980,N_10966);
and U11389 (N_11389,N_10910,N_10923);
nand U11390 (N_11390,N_11039,N_11176);
nand U11391 (N_11391,N_10847,N_11145);
nor U11392 (N_11392,N_10907,N_10872);
xor U11393 (N_11393,N_10946,N_11147);
nor U11394 (N_11394,N_11021,N_11187);
xnor U11395 (N_11395,N_11003,N_10829);
nor U11396 (N_11396,N_11161,N_10900);
and U11397 (N_11397,N_11044,N_11130);
and U11398 (N_11398,N_11054,N_10950);
and U11399 (N_11399,N_10938,N_10834);
nand U11400 (N_11400,N_10927,N_10818);
nor U11401 (N_11401,N_11074,N_10951);
xor U11402 (N_11402,N_11116,N_10967);
and U11403 (N_11403,N_11059,N_10960);
and U11404 (N_11404,N_10855,N_11090);
or U11405 (N_11405,N_10930,N_11183);
xnor U11406 (N_11406,N_10925,N_11039);
xor U11407 (N_11407,N_10821,N_11153);
nor U11408 (N_11408,N_10886,N_10903);
nor U11409 (N_11409,N_10971,N_10980);
or U11410 (N_11410,N_11044,N_10848);
nand U11411 (N_11411,N_10863,N_11183);
or U11412 (N_11412,N_11043,N_11080);
nand U11413 (N_11413,N_10973,N_10962);
nor U11414 (N_11414,N_10929,N_10845);
and U11415 (N_11415,N_10816,N_11139);
nor U11416 (N_11416,N_11036,N_10907);
xnor U11417 (N_11417,N_11134,N_11185);
and U11418 (N_11418,N_10885,N_10869);
and U11419 (N_11419,N_10939,N_11129);
nand U11420 (N_11420,N_10998,N_11112);
nand U11421 (N_11421,N_11020,N_10973);
xnor U11422 (N_11422,N_10897,N_10893);
xnor U11423 (N_11423,N_10875,N_10985);
nor U11424 (N_11424,N_10877,N_10907);
or U11425 (N_11425,N_10975,N_11043);
and U11426 (N_11426,N_11061,N_11174);
nand U11427 (N_11427,N_10860,N_10948);
xor U11428 (N_11428,N_10815,N_11105);
and U11429 (N_11429,N_11144,N_10917);
xor U11430 (N_11430,N_11187,N_10817);
nand U11431 (N_11431,N_10994,N_11185);
and U11432 (N_11432,N_11169,N_10985);
or U11433 (N_11433,N_10910,N_10889);
xor U11434 (N_11434,N_11135,N_10839);
nand U11435 (N_11435,N_10822,N_10961);
xor U11436 (N_11436,N_11041,N_10967);
and U11437 (N_11437,N_10816,N_11110);
nor U11438 (N_11438,N_10933,N_11198);
or U11439 (N_11439,N_11119,N_10853);
or U11440 (N_11440,N_11152,N_11158);
xnor U11441 (N_11441,N_10859,N_11171);
and U11442 (N_11442,N_10802,N_11003);
nand U11443 (N_11443,N_11130,N_11194);
nor U11444 (N_11444,N_10851,N_11095);
xnor U11445 (N_11445,N_10804,N_10962);
and U11446 (N_11446,N_11084,N_10812);
nand U11447 (N_11447,N_11116,N_10805);
and U11448 (N_11448,N_10973,N_11056);
or U11449 (N_11449,N_11161,N_10834);
nand U11450 (N_11450,N_11009,N_10996);
xnor U11451 (N_11451,N_10824,N_10981);
nor U11452 (N_11452,N_10880,N_11002);
nand U11453 (N_11453,N_11158,N_10969);
xnor U11454 (N_11454,N_11003,N_10895);
xnor U11455 (N_11455,N_11051,N_10931);
nand U11456 (N_11456,N_10806,N_11135);
or U11457 (N_11457,N_11061,N_10975);
or U11458 (N_11458,N_11033,N_11184);
nor U11459 (N_11459,N_10803,N_11030);
or U11460 (N_11460,N_10970,N_10928);
xor U11461 (N_11461,N_10816,N_10846);
and U11462 (N_11462,N_10992,N_10872);
and U11463 (N_11463,N_10903,N_11026);
nand U11464 (N_11464,N_10869,N_10892);
and U11465 (N_11465,N_11070,N_11021);
nor U11466 (N_11466,N_10938,N_10999);
and U11467 (N_11467,N_10903,N_10837);
or U11468 (N_11468,N_10844,N_10841);
xnor U11469 (N_11469,N_10896,N_11070);
nor U11470 (N_11470,N_10865,N_11033);
xnor U11471 (N_11471,N_10956,N_11175);
nand U11472 (N_11472,N_10874,N_10992);
and U11473 (N_11473,N_10903,N_10842);
and U11474 (N_11474,N_10806,N_10901);
and U11475 (N_11475,N_11096,N_10957);
or U11476 (N_11476,N_10905,N_10833);
and U11477 (N_11477,N_11026,N_10997);
or U11478 (N_11478,N_10863,N_10933);
xnor U11479 (N_11479,N_10960,N_10884);
and U11480 (N_11480,N_11077,N_10970);
nor U11481 (N_11481,N_11167,N_11186);
nor U11482 (N_11482,N_10844,N_11113);
or U11483 (N_11483,N_11127,N_11023);
nor U11484 (N_11484,N_11060,N_11043);
xnor U11485 (N_11485,N_10995,N_10978);
nor U11486 (N_11486,N_11109,N_10870);
and U11487 (N_11487,N_11191,N_11105);
and U11488 (N_11488,N_11142,N_11014);
or U11489 (N_11489,N_11022,N_11107);
and U11490 (N_11490,N_10944,N_10820);
or U11491 (N_11491,N_11009,N_11173);
or U11492 (N_11492,N_10924,N_10932);
nand U11493 (N_11493,N_10963,N_10847);
xor U11494 (N_11494,N_11161,N_11089);
and U11495 (N_11495,N_10974,N_10804);
nor U11496 (N_11496,N_11115,N_10860);
nand U11497 (N_11497,N_11044,N_10802);
nor U11498 (N_11498,N_10940,N_10934);
xnor U11499 (N_11499,N_11004,N_10947);
or U11500 (N_11500,N_11039,N_10869);
nand U11501 (N_11501,N_10958,N_10969);
nor U11502 (N_11502,N_11186,N_10970);
or U11503 (N_11503,N_11065,N_11059);
nand U11504 (N_11504,N_10972,N_10897);
xor U11505 (N_11505,N_10962,N_10877);
nand U11506 (N_11506,N_11118,N_10826);
nor U11507 (N_11507,N_10940,N_11147);
nor U11508 (N_11508,N_10846,N_10835);
xor U11509 (N_11509,N_11055,N_10923);
and U11510 (N_11510,N_11167,N_11055);
or U11511 (N_11511,N_10978,N_10906);
and U11512 (N_11512,N_10897,N_11193);
xor U11513 (N_11513,N_10835,N_11011);
and U11514 (N_11514,N_10885,N_11167);
xor U11515 (N_11515,N_10939,N_10843);
or U11516 (N_11516,N_10921,N_10999);
or U11517 (N_11517,N_10844,N_11012);
or U11518 (N_11518,N_11059,N_10977);
or U11519 (N_11519,N_11035,N_11106);
and U11520 (N_11520,N_10833,N_11183);
nand U11521 (N_11521,N_10848,N_10987);
nor U11522 (N_11522,N_10910,N_10807);
and U11523 (N_11523,N_10805,N_11130);
nor U11524 (N_11524,N_10880,N_11159);
xnor U11525 (N_11525,N_11106,N_10867);
and U11526 (N_11526,N_10911,N_11006);
or U11527 (N_11527,N_11156,N_11188);
nor U11528 (N_11528,N_10814,N_10835);
nand U11529 (N_11529,N_11028,N_10894);
nor U11530 (N_11530,N_10821,N_11162);
nand U11531 (N_11531,N_11014,N_10930);
and U11532 (N_11532,N_10902,N_11047);
xnor U11533 (N_11533,N_10830,N_11132);
nand U11534 (N_11534,N_10815,N_11034);
nand U11535 (N_11535,N_10863,N_11085);
xnor U11536 (N_11536,N_10843,N_10908);
and U11537 (N_11537,N_10889,N_10940);
nor U11538 (N_11538,N_10981,N_10831);
and U11539 (N_11539,N_11144,N_10899);
or U11540 (N_11540,N_10839,N_11125);
or U11541 (N_11541,N_11185,N_11060);
and U11542 (N_11542,N_11005,N_10815);
nor U11543 (N_11543,N_10854,N_10845);
or U11544 (N_11544,N_11045,N_10990);
nand U11545 (N_11545,N_10982,N_11123);
xnor U11546 (N_11546,N_10887,N_10821);
nor U11547 (N_11547,N_11116,N_10944);
and U11548 (N_11548,N_10959,N_11156);
nand U11549 (N_11549,N_10859,N_11161);
nor U11550 (N_11550,N_11178,N_10832);
xnor U11551 (N_11551,N_11196,N_11026);
nand U11552 (N_11552,N_10854,N_10883);
nand U11553 (N_11553,N_11109,N_11126);
nor U11554 (N_11554,N_10977,N_10812);
and U11555 (N_11555,N_10923,N_11146);
nor U11556 (N_11556,N_11124,N_10984);
nand U11557 (N_11557,N_11088,N_10944);
and U11558 (N_11558,N_11023,N_11199);
nor U11559 (N_11559,N_10976,N_10840);
nor U11560 (N_11560,N_11123,N_11138);
nor U11561 (N_11561,N_10926,N_10868);
nand U11562 (N_11562,N_10807,N_11194);
xnor U11563 (N_11563,N_10900,N_10810);
and U11564 (N_11564,N_10878,N_10924);
xor U11565 (N_11565,N_10912,N_11158);
or U11566 (N_11566,N_11027,N_11038);
and U11567 (N_11567,N_11006,N_10877);
or U11568 (N_11568,N_11138,N_11092);
nand U11569 (N_11569,N_10868,N_11192);
xnor U11570 (N_11570,N_10984,N_11058);
nand U11571 (N_11571,N_10948,N_11099);
xor U11572 (N_11572,N_11044,N_10815);
nor U11573 (N_11573,N_11034,N_11197);
nand U11574 (N_11574,N_11114,N_11184);
and U11575 (N_11575,N_10878,N_10931);
nand U11576 (N_11576,N_10824,N_11027);
nand U11577 (N_11577,N_10949,N_10854);
xor U11578 (N_11578,N_11077,N_11090);
or U11579 (N_11579,N_10819,N_11129);
nand U11580 (N_11580,N_11025,N_11199);
nor U11581 (N_11581,N_10991,N_10813);
or U11582 (N_11582,N_11065,N_11030);
xnor U11583 (N_11583,N_11039,N_11005);
xnor U11584 (N_11584,N_10823,N_10900);
nand U11585 (N_11585,N_10929,N_10854);
or U11586 (N_11586,N_11051,N_10841);
and U11587 (N_11587,N_10878,N_11001);
nand U11588 (N_11588,N_11026,N_10866);
nor U11589 (N_11589,N_11037,N_10818);
nand U11590 (N_11590,N_11132,N_11047);
nand U11591 (N_11591,N_10935,N_11027);
xnor U11592 (N_11592,N_11043,N_11142);
or U11593 (N_11593,N_10848,N_11052);
and U11594 (N_11594,N_11143,N_10949);
nand U11595 (N_11595,N_11047,N_11105);
xor U11596 (N_11596,N_11099,N_11057);
nand U11597 (N_11597,N_10961,N_11132);
or U11598 (N_11598,N_11094,N_11044);
nand U11599 (N_11599,N_11195,N_10801);
nand U11600 (N_11600,N_11252,N_11224);
nand U11601 (N_11601,N_11484,N_11255);
or U11602 (N_11602,N_11253,N_11515);
xor U11603 (N_11603,N_11431,N_11341);
or U11604 (N_11604,N_11398,N_11483);
nor U11605 (N_11605,N_11239,N_11569);
nor U11606 (N_11606,N_11283,N_11510);
or U11607 (N_11607,N_11392,N_11373);
nor U11608 (N_11608,N_11383,N_11324);
and U11609 (N_11609,N_11216,N_11347);
or U11610 (N_11610,N_11335,N_11272);
and U11611 (N_11611,N_11466,N_11560);
and U11612 (N_11612,N_11501,N_11305);
xor U11613 (N_11613,N_11280,N_11288);
nand U11614 (N_11614,N_11217,N_11410);
xnor U11615 (N_11615,N_11480,N_11325);
nand U11616 (N_11616,N_11586,N_11476);
nand U11617 (N_11617,N_11457,N_11320);
xnor U11618 (N_11618,N_11414,N_11459);
xnor U11619 (N_11619,N_11573,N_11578);
xor U11620 (N_11620,N_11566,N_11267);
xnor U11621 (N_11621,N_11428,N_11424);
or U11622 (N_11622,N_11562,N_11449);
nand U11623 (N_11623,N_11526,N_11319);
xor U11624 (N_11624,N_11505,N_11437);
xnor U11625 (N_11625,N_11295,N_11380);
and U11626 (N_11626,N_11208,N_11277);
or U11627 (N_11627,N_11390,N_11436);
and U11628 (N_11628,N_11502,N_11202);
nor U11629 (N_11629,N_11420,N_11386);
or U11630 (N_11630,N_11470,N_11258);
nand U11631 (N_11631,N_11469,N_11337);
or U11632 (N_11632,N_11233,N_11353);
and U11633 (N_11633,N_11399,N_11238);
and U11634 (N_11634,N_11475,N_11473);
and U11635 (N_11635,N_11522,N_11456);
nand U11636 (N_11636,N_11525,N_11210);
nor U11637 (N_11637,N_11517,N_11381);
and U11638 (N_11638,N_11362,N_11550);
and U11639 (N_11639,N_11364,N_11508);
and U11640 (N_11640,N_11260,N_11306);
nand U11641 (N_11641,N_11318,N_11450);
xor U11642 (N_11642,N_11453,N_11412);
xnor U11643 (N_11643,N_11552,N_11571);
xor U11644 (N_11644,N_11230,N_11557);
nand U11645 (N_11645,N_11554,N_11518);
or U11646 (N_11646,N_11213,N_11312);
xor U11647 (N_11647,N_11395,N_11532);
nor U11648 (N_11648,N_11326,N_11530);
nor U11649 (N_11649,N_11598,N_11268);
and U11650 (N_11650,N_11223,N_11355);
nor U11651 (N_11651,N_11350,N_11561);
and U11652 (N_11652,N_11316,N_11374);
or U11653 (N_11653,N_11235,N_11504);
or U11654 (N_11654,N_11568,N_11265);
xor U11655 (N_11655,N_11489,N_11580);
nand U11656 (N_11656,N_11538,N_11313);
xnor U11657 (N_11657,N_11241,N_11503);
nand U11658 (N_11658,N_11291,N_11487);
nor U11659 (N_11659,N_11274,N_11369);
and U11660 (N_11660,N_11592,N_11345);
nor U11661 (N_11661,N_11323,N_11559);
nor U11662 (N_11662,N_11472,N_11418);
nand U11663 (N_11663,N_11528,N_11303);
xnor U11664 (N_11664,N_11356,N_11371);
nand U11665 (N_11665,N_11259,N_11546);
and U11666 (N_11666,N_11273,N_11269);
nor U11667 (N_11667,N_11296,N_11376);
nand U11668 (N_11668,N_11458,N_11464);
and U11669 (N_11669,N_11226,N_11520);
nand U11670 (N_11670,N_11279,N_11556);
and U11671 (N_11671,N_11465,N_11594);
or U11672 (N_11672,N_11361,N_11521);
and U11673 (N_11673,N_11330,N_11408);
nor U11674 (N_11674,N_11462,N_11354);
nand U11675 (N_11675,N_11551,N_11553);
nand U11676 (N_11676,N_11490,N_11493);
nor U11677 (N_11677,N_11447,N_11486);
xnor U11678 (N_11678,N_11596,N_11468);
nand U11679 (N_11679,N_11271,N_11506);
nand U11680 (N_11680,N_11200,N_11382);
nor U11681 (N_11681,N_11509,N_11227);
and U11682 (N_11682,N_11264,N_11523);
nand U11683 (N_11683,N_11293,N_11589);
xnor U11684 (N_11684,N_11240,N_11304);
or U11685 (N_11685,N_11276,N_11375);
nor U11686 (N_11686,N_11218,N_11467);
nor U11687 (N_11687,N_11455,N_11315);
or U11688 (N_11688,N_11360,N_11359);
nor U11689 (N_11689,N_11294,N_11488);
or U11690 (N_11690,N_11593,N_11211);
nor U11691 (N_11691,N_11421,N_11401);
nor U11692 (N_11692,N_11249,N_11242);
xnor U11693 (N_11693,N_11286,N_11220);
nand U11694 (N_11694,N_11494,N_11368);
or U11695 (N_11695,N_11426,N_11496);
nand U11696 (N_11696,N_11314,N_11278);
nor U11697 (N_11697,N_11405,N_11251);
xor U11698 (N_11698,N_11535,N_11246);
nand U11699 (N_11699,N_11244,N_11367);
and U11700 (N_11700,N_11377,N_11282);
nand U11701 (N_11701,N_11474,N_11477);
nor U11702 (N_11702,N_11558,N_11400);
or U11703 (N_11703,N_11429,N_11397);
xnor U11704 (N_11704,N_11581,N_11454);
nor U11705 (N_11705,N_11500,N_11292);
and U11706 (N_11706,N_11433,N_11463);
nand U11707 (N_11707,N_11221,N_11229);
xnor U11708 (N_11708,N_11519,N_11411);
nand U11709 (N_11709,N_11302,N_11555);
nor U11710 (N_11710,N_11572,N_11537);
nand U11711 (N_11711,N_11591,N_11570);
nor U11712 (N_11712,N_11225,N_11387);
and U11713 (N_11713,N_11284,N_11346);
nor U11714 (N_11714,N_11232,N_11434);
nor U11715 (N_11715,N_11334,N_11539);
or U11716 (N_11716,N_11497,N_11404);
and U11717 (N_11717,N_11287,N_11451);
or U11718 (N_11718,N_11297,N_11243);
and U11719 (N_11719,N_11406,N_11247);
or U11720 (N_11720,N_11513,N_11416);
or U11721 (N_11721,N_11435,N_11511);
nand U11722 (N_11722,N_11499,N_11385);
xor U11723 (N_11723,N_11485,N_11575);
and U11724 (N_11724,N_11516,N_11492);
nor U11725 (N_11725,N_11425,N_11236);
xor U11726 (N_11726,N_11542,N_11394);
and U11727 (N_11727,N_11479,N_11384);
and U11728 (N_11728,N_11270,N_11442);
nor U11729 (N_11729,N_11328,N_11263);
or U11730 (N_11730,N_11372,N_11254);
and U11731 (N_11731,N_11512,N_11402);
nand U11732 (N_11732,N_11219,N_11438);
and U11733 (N_11733,N_11257,N_11444);
nand U11734 (N_11734,N_11262,N_11440);
nand U11735 (N_11735,N_11298,N_11333);
nor U11736 (N_11736,N_11524,N_11363);
xnor U11737 (N_11737,N_11482,N_11419);
xor U11738 (N_11738,N_11340,N_11234);
and U11739 (N_11739,N_11309,N_11527);
nand U11740 (N_11740,N_11228,N_11543);
xor U11741 (N_11741,N_11595,N_11514);
nor U11742 (N_11742,N_11307,N_11478);
nand U11743 (N_11743,N_11203,N_11248);
or U11744 (N_11744,N_11365,N_11544);
or U11745 (N_11745,N_11388,N_11245);
nand U11746 (N_11746,N_11461,N_11391);
nand U11747 (N_11747,N_11417,N_11205);
nor U11748 (N_11748,N_11222,N_11332);
or U11749 (N_11749,N_11409,N_11256);
nor U11750 (N_11750,N_11310,N_11201);
xnor U11751 (N_11751,N_11507,N_11351);
nand U11752 (N_11752,N_11577,N_11261);
nand U11753 (N_11753,N_11413,N_11357);
xnor U11754 (N_11754,N_11549,N_11352);
xor U11755 (N_11755,N_11582,N_11545);
and U11756 (N_11756,N_11331,N_11299);
nor U11757 (N_11757,N_11441,N_11567);
xor U11758 (N_11758,N_11336,N_11423);
or U11759 (N_11759,N_11548,N_11498);
nor U11760 (N_11760,N_11533,N_11393);
nor U11761 (N_11761,N_11321,N_11481);
nand U11762 (N_11762,N_11290,N_11491);
and U11763 (N_11763,N_11452,N_11531);
or U11764 (N_11764,N_11275,N_11446);
or U11765 (N_11765,N_11301,N_11237);
xnor U11766 (N_11766,N_11212,N_11427);
and U11767 (N_11767,N_11266,N_11563);
and U11768 (N_11768,N_11378,N_11327);
nand U11769 (N_11769,N_11432,N_11448);
and U11770 (N_11770,N_11585,N_11206);
and U11771 (N_11771,N_11389,N_11460);
and U11772 (N_11772,N_11343,N_11587);
xor U11773 (N_11773,N_11342,N_11445);
xnor U11774 (N_11774,N_11308,N_11564);
nand U11775 (N_11775,N_11407,N_11231);
or U11776 (N_11776,N_11322,N_11536);
nand U11777 (N_11777,N_11344,N_11396);
xor U11778 (N_11778,N_11370,N_11430);
xnor U11779 (N_11779,N_11250,N_11289);
or U11780 (N_11780,N_11207,N_11338);
nor U11781 (N_11781,N_11588,N_11329);
or U11782 (N_11782,N_11439,N_11540);
nor U11783 (N_11783,N_11471,N_11415);
nor U11784 (N_11784,N_11529,N_11215);
or U11785 (N_11785,N_11285,N_11311);
or U11786 (N_11786,N_11204,N_11317);
nor U11787 (N_11787,N_11300,N_11214);
and U11788 (N_11788,N_11495,N_11209);
or U11789 (N_11789,N_11348,N_11590);
and U11790 (N_11790,N_11379,N_11366);
nor U11791 (N_11791,N_11443,N_11565);
nand U11792 (N_11792,N_11579,N_11574);
and U11793 (N_11793,N_11583,N_11422);
xor U11794 (N_11794,N_11339,N_11597);
or U11795 (N_11795,N_11584,N_11576);
nand U11796 (N_11796,N_11349,N_11541);
xor U11797 (N_11797,N_11547,N_11281);
or U11798 (N_11798,N_11403,N_11534);
nand U11799 (N_11799,N_11358,N_11599);
and U11800 (N_11800,N_11470,N_11543);
nor U11801 (N_11801,N_11215,N_11387);
nor U11802 (N_11802,N_11575,N_11328);
and U11803 (N_11803,N_11370,N_11335);
or U11804 (N_11804,N_11594,N_11398);
nor U11805 (N_11805,N_11547,N_11352);
nand U11806 (N_11806,N_11460,N_11306);
or U11807 (N_11807,N_11245,N_11556);
nor U11808 (N_11808,N_11549,N_11479);
or U11809 (N_11809,N_11426,N_11484);
xnor U11810 (N_11810,N_11495,N_11484);
xor U11811 (N_11811,N_11419,N_11280);
or U11812 (N_11812,N_11320,N_11486);
xor U11813 (N_11813,N_11520,N_11586);
nand U11814 (N_11814,N_11574,N_11325);
and U11815 (N_11815,N_11262,N_11517);
nor U11816 (N_11816,N_11554,N_11361);
and U11817 (N_11817,N_11485,N_11270);
xor U11818 (N_11818,N_11255,N_11440);
xor U11819 (N_11819,N_11430,N_11234);
or U11820 (N_11820,N_11463,N_11313);
or U11821 (N_11821,N_11569,N_11245);
nand U11822 (N_11822,N_11379,N_11521);
nor U11823 (N_11823,N_11532,N_11219);
or U11824 (N_11824,N_11525,N_11313);
nor U11825 (N_11825,N_11216,N_11358);
or U11826 (N_11826,N_11547,N_11201);
or U11827 (N_11827,N_11391,N_11336);
nand U11828 (N_11828,N_11375,N_11284);
xnor U11829 (N_11829,N_11278,N_11529);
xnor U11830 (N_11830,N_11388,N_11340);
nand U11831 (N_11831,N_11485,N_11593);
xnor U11832 (N_11832,N_11219,N_11368);
and U11833 (N_11833,N_11241,N_11330);
and U11834 (N_11834,N_11214,N_11598);
and U11835 (N_11835,N_11376,N_11204);
or U11836 (N_11836,N_11450,N_11483);
and U11837 (N_11837,N_11342,N_11201);
and U11838 (N_11838,N_11598,N_11556);
or U11839 (N_11839,N_11576,N_11299);
nand U11840 (N_11840,N_11324,N_11281);
nand U11841 (N_11841,N_11287,N_11459);
nand U11842 (N_11842,N_11228,N_11454);
and U11843 (N_11843,N_11484,N_11239);
or U11844 (N_11844,N_11517,N_11536);
xor U11845 (N_11845,N_11484,N_11345);
and U11846 (N_11846,N_11556,N_11360);
or U11847 (N_11847,N_11438,N_11360);
nand U11848 (N_11848,N_11454,N_11261);
nand U11849 (N_11849,N_11432,N_11469);
xnor U11850 (N_11850,N_11375,N_11395);
xnor U11851 (N_11851,N_11338,N_11584);
xor U11852 (N_11852,N_11426,N_11361);
nor U11853 (N_11853,N_11317,N_11372);
nand U11854 (N_11854,N_11415,N_11350);
or U11855 (N_11855,N_11244,N_11526);
xnor U11856 (N_11856,N_11546,N_11284);
nand U11857 (N_11857,N_11534,N_11598);
xor U11858 (N_11858,N_11462,N_11408);
and U11859 (N_11859,N_11331,N_11459);
and U11860 (N_11860,N_11273,N_11411);
xnor U11861 (N_11861,N_11531,N_11568);
or U11862 (N_11862,N_11513,N_11586);
xor U11863 (N_11863,N_11315,N_11545);
xor U11864 (N_11864,N_11320,N_11285);
nor U11865 (N_11865,N_11558,N_11459);
nor U11866 (N_11866,N_11384,N_11295);
xnor U11867 (N_11867,N_11468,N_11295);
xor U11868 (N_11868,N_11230,N_11536);
xnor U11869 (N_11869,N_11587,N_11465);
or U11870 (N_11870,N_11270,N_11430);
and U11871 (N_11871,N_11508,N_11294);
nand U11872 (N_11872,N_11354,N_11226);
and U11873 (N_11873,N_11585,N_11497);
and U11874 (N_11874,N_11552,N_11215);
xor U11875 (N_11875,N_11426,N_11433);
or U11876 (N_11876,N_11563,N_11577);
and U11877 (N_11877,N_11376,N_11253);
nor U11878 (N_11878,N_11211,N_11467);
and U11879 (N_11879,N_11214,N_11281);
or U11880 (N_11880,N_11494,N_11410);
nand U11881 (N_11881,N_11400,N_11208);
nor U11882 (N_11882,N_11553,N_11326);
or U11883 (N_11883,N_11420,N_11222);
or U11884 (N_11884,N_11482,N_11545);
and U11885 (N_11885,N_11230,N_11439);
nand U11886 (N_11886,N_11514,N_11403);
nor U11887 (N_11887,N_11321,N_11515);
nor U11888 (N_11888,N_11446,N_11321);
nor U11889 (N_11889,N_11409,N_11416);
or U11890 (N_11890,N_11373,N_11324);
nor U11891 (N_11891,N_11273,N_11421);
and U11892 (N_11892,N_11582,N_11477);
and U11893 (N_11893,N_11386,N_11390);
and U11894 (N_11894,N_11398,N_11204);
xnor U11895 (N_11895,N_11584,N_11499);
and U11896 (N_11896,N_11310,N_11392);
or U11897 (N_11897,N_11321,N_11535);
nand U11898 (N_11898,N_11537,N_11274);
or U11899 (N_11899,N_11243,N_11556);
nand U11900 (N_11900,N_11444,N_11372);
xnor U11901 (N_11901,N_11529,N_11353);
xor U11902 (N_11902,N_11232,N_11400);
nor U11903 (N_11903,N_11302,N_11586);
xor U11904 (N_11904,N_11586,N_11501);
or U11905 (N_11905,N_11256,N_11462);
nor U11906 (N_11906,N_11360,N_11378);
or U11907 (N_11907,N_11517,N_11368);
or U11908 (N_11908,N_11366,N_11226);
nor U11909 (N_11909,N_11264,N_11481);
or U11910 (N_11910,N_11562,N_11347);
and U11911 (N_11911,N_11299,N_11227);
xor U11912 (N_11912,N_11518,N_11370);
nor U11913 (N_11913,N_11449,N_11432);
nand U11914 (N_11914,N_11531,N_11519);
xnor U11915 (N_11915,N_11357,N_11308);
and U11916 (N_11916,N_11245,N_11534);
and U11917 (N_11917,N_11389,N_11469);
xnor U11918 (N_11918,N_11283,N_11545);
nor U11919 (N_11919,N_11211,N_11452);
and U11920 (N_11920,N_11471,N_11483);
nor U11921 (N_11921,N_11452,N_11540);
nand U11922 (N_11922,N_11201,N_11579);
or U11923 (N_11923,N_11309,N_11567);
and U11924 (N_11924,N_11270,N_11595);
nor U11925 (N_11925,N_11436,N_11352);
nor U11926 (N_11926,N_11433,N_11474);
nor U11927 (N_11927,N_11326,N_11201);
or U11928 (N_11928,N_11327,N_11356);
and U11929 (N_11929,N_11331,N_11494);
or U11930 (N_11930,N_11447,N_11200);
nand U11931 (N_11931,N_11440,N_11393);
or U11932 (N_11932,N_11269,N_11278);
xor U11933 (N_11933,N_11595,N_11472);
nand U11934 (N_11934,N_11594,N_11239);
xor U11935 (N_11935,N_11587,N_11365);
nand U11936 (N_11936,N_11409,N_11228);
nor U11937 (N_11937,N_11404,N_11478);
nor U11938 (N_11938,N_11596,N_11370);
or U11939 (N_11939,N_11377,N_11205);
nor U11940 (N_11940,N_11208,N_11388);
and U11941 (N_11941,N_11554,N_11489);
and U11942 (N_11942,N_11307,N_11499);
nor U11943 (N_11943,N_11200,N_11457);
nor U11944 (N_11944,N_11508,N_11450);
xor U11945 (N_11945,N_11548,N_11502);
and U11946 (N_11946,N_11542,N_11565);
nor U11947 (N_11947,N_11304,N_11498);
nor U11948 (N_11948,N_11327,N_11531);
nand U11949 (N_11949,N_11385,N_11488);
or U11950 (N_11950,N_11516,N_11524);
nor U11951 (N_11951,N_11283,N_11493);
nor U11952 (N_11952,N_11363,N_11395);
nand U11953 (N_11953,N_11476,N_11223);
nand U11954 (N_11954,N_11461,N_11479);
nor U11955 (N_11955,N_11260,N_11562);
and U11956 (N_11956,N_11384,N_11273);
nor U11957 (N_11957,N_11308,N_11432);
and U11958 (N_11958,N_11506,N_11474);
xor U11959 (N_11959,N_11496,N_11586);
or U11960 (N_11960,N_11487,N_11475);
and U11961 (N_11961,N_11576,N_11497);
nand U11962 (N_11962,N_11260,N_11274);
nor U11963 (N_11963,N_11476,N_11419);
and U11964 (N_11964,N_11303,N_11217);
or U11965 (N_11965,N_11223,N_11262);
nand U11966 (N_11966,N_11551,N_11349);
nand U11967 (N_11967,N_11245,N_11384);
and U11968 (N_11968,N_11544,N_11419);
nand U11969 (N_11969,N_11266,N_11598);
and U11970 (N_11970,N_11216,N_11568);
nand U11971 (N_11971,N_11435,N_11512);
or U11972 (N_11972,N_11375,N_11496);
and U11973 (N_11973,N_11520,N_11396);
or U11974 (N_11974,N_11230,N_11268);
nor U11975 (N_11975,N_11496,N_11482);
xor U11976 (N_11976,N_11270,N_11231);
nor U11977 (N_11977,N_11581,N_11519);
nand U11978 (N_11978,N_11418,N_11450);
and U11979 (N_11979,N_11471,N_11212);
xor U11980 (N_11980,N_11428,N_11254);
and U11981 (N_11981,N_11210,N_11300);
nand U11982 (N_11982,N_11282,N_11400);
nand U11983 (N_11983,N_11569,N_11219);
xor U11984 (N_11984,N_11534,N_11270);
nor U11985 (N_11985,N_11310,N_11406);
xnor U11986 (N_11986,N_11203,N_11560);
and U11987 (N_11987,N_11220,N_11545);
nand U11988 (N_11988,N_11307,N_11249);
and U11989 (N_11989,N_11486,N_11490);
xor U11990 (N_11990,N_11299,N_11375);
xor U11991 (N_11991,N_11343,N_11425);
nor U11992 (N_11992,N_11560,N_11404);
nor U11993 (N_11993,N_11572,N_11551);
xnor U11994 (N_11994,N_11581,N_11377);
nand U11995 (N_11995,N_11469,N_11585);
and U11996 (N_11996,N_11395,N_11208);
nor U11997 (N_11997,N_11580,N_11385);
xor U11998 (N_11998,N_11550,N_11513);
nand U11999 (N_11999,N_11412,N_11313);
or U12000 (N_12000,N_11693,N_11602);
and U12001 (N_12001,N_11617,N_11868);
nor U12002 (N_12002,N_11755,N_11870);
and U12003 (N_12003,N_11985,N_11747);
nand U12004 (N_12004,N_11927,N_11765);
and U12005 (N_12005,N_11713,N_11632);
nand U12006 (N_12006,N_11790,N_11768);
and U12007 (N_12007,N_11802,N_11879);
and U12008 (N_12008,N_11669,N_11795);
nand U12009 (N_12009,N_11645,N_11851);
xor U12010 (N_12010,N_11909,N_11697);
and U12011 (N_12011,N_11857,N_11903);
xnor U12012 (N_12012,N_11630,N_11629);
or U12013 (N_12013,N_11968,N_11711);
xor U12014 (N_12014,N_11971,N_11840);
xnor U12015 (N_12015,N_11935,N_11732);
and U12016 (N_12016,N_11875,N_11637);
and U12017 (N_12017,N_11657,N_11804);
or U12018 (N_12018,N_11845,N_11627);
and U12019 (N_12019,N_11715,N_11818);
and U12020 (N_12020,N_11685,N_11690);
nor U12021 (N_12021,N_11731,N_11744);
or U12022 (N_12022,N_11673,N_11972);
and U12023 (N_12023,N_11740,N_11932);
nor U12024 (N_12024,N_11862,N_11962);
and U12025 (N_12025,N_11748,N_11853);
nor U12026 (N_12026,N_11953,N_11904);
or U12027 (N_12027,N_11681,N_11781);
nor U12028 (N_12028,N_11808,N_11915);
xnor U12029 (N_12029,N_11722,N_11729);
and U12030 (N_12030,N_11736,N_11982);
nand U12031 (N_12031,N_11674,N_11896);
xor U12032 (N_12032,N_11905,N_11668);
or U12033 (N_12033,N_11821,N_11803);
xnor U12034 (N_12034,N_11825,N_11965);
and U12035 (N_12035,N_11719,N_11882);
or U12036 (N_12036,N_11837,N_11652);
xor U12037 (N_12037,N_11753,N_11976);
or U12038 (N_12038,N_11923,N_11613);
xor U12039 (N_12039,N_11937,N_11767);
xnor U12040 (N_12040,N_11786,N_11716);
and U12041 (N_12041,N_11960,N_11607);
nand U12042 (N_12042,N_11757,N_11936);
nand U12043 (N_12043,N_11819,N_11728);
nand U12044 (N_12044,N_11720,N_11707);
nor U12045 (N_12045,N_11718,N_11634);
xor U12046 (N_12046,N_11631,N_11611);
or U12047 (N_12047,N_11815,N_11626);
xor U12048 (N_12048,N_11799,N_11969);
and U12049 (N_12049,N_11788,N_11725);
nor U12050 (N_12050,N_11745,N_11770);
xor U12051 (N_12051,N_11908,N_11890);
nand U12052 (N_12052,N_11616,N_11911);
and U12053 (N_12053,N_11996,N_11615);
or U12054 (N_12054,N_11894,N_11966);
and U12055 (N_12055,N_11625,N_11689);
xor U12056 (N_12056,N_11672,N_11656);
xor U12057 (N_12057,N_11761,N_11798);
and U12058 (N_12058,N_11628,N_11891);
and U12059 (N_12059,N_11604,N_11942);
or U12060 (N_12060,N_11900,N_11858);
xnor U12061 (N_12061,N_11874,N_11924);
nor U12062 (N_12062,N_11662,N_11785);
nand U12063 (N_12063,N_11764,N_11940);
or U12064 (N_12064,N_11961,N_11843);
xor U12065 (N_12065,N_11792,N_11827);
nor U12066 (N_12066,N_11738,N_11991);
and U12067 (N_12067,N_11665,N_11778);
xnor U12068 (N_12068,N_11947,N_11609);
nor U12069 (N_12069,N_11925,N_11601);
nand U12070 (N_12070,N_11897,N_11649);
nand U12071 (N_12071,N_11832,N_11952);
and U12072 (N_12072,N_11812,N_11641);
and U12073 (N_12073,N_11885,N_11756);
and U12074 (N_12074,N_11763,N_11855);
or U12075 (N_12075,N_11854,N_11724);
nor U12076 (N_12076,N_11954,N_11823);
xnor U12077 (N_12077,N_11998,N_11774);
xor U12078 (N_12078,N_11675,N_11898);
nor U12079 (N_12079,N_11635,N_11886);
and U12080 (N_12080,N_11796,N_11640);
nand U12081 (N_12081,N_11918,N_11957);
or U12082 (N_12082,N_11861,N_11852);
and U12083 (N_12083,N_11844,N_11906);
or U12084 (N_12084,N_11679,N_11913);
xor U12085 (N_12085,N_11916,N_11987);
nand U12086 (N_12086,N_11734,N_11794);
nor U12087 (N_12087,N_11723,N_11981);
xnor U12088 (N_12088,N_11610,N_11813);
nand U12089 (N_12089,N_11780,N_11783);
or U12090 (N_12090,N_11977,N_11810);
or U12091 (N_12091,N_11699,N_11730);
or U12092 (N_12092,N_11789,N_11647);
nor U12093 (N_12093,N_11816,N_11726);
nor U12094 (N_12094,N_11926,N_11817);
or U12095 (N_12095,N_11620,N_11989);
or U12096 (N_12096,N_11691,N_11717);
and U12097 (N_12097,N_11603,N_11850);
xnor U12098 (N_12098,N_11921,N_11992);
and U12099 (N_12099,N_11702,N_11979);
or U12100 (N_12100,N_11871,N_11907);
or U12101 (N_12101,N_11828,N_11983);
or U12102 (N_12102,N_11865,N_11883);
nor U12103 (N_12103,N_11791,N_11706);
nand U12104 (N_12104,N_11737,N_11650);
xor U12105 (N_12105,N_11990,N_11614);
or U12106 (N_12106,N_11884,N_11950);
or U12107 (N_12107,N_11750,N_11931);
or U12108 (N_12108,N_11683,N_11880);
and U12109 (N_12109,N_11671,N_11914);
xor U12110 (N_12110,N_11997,N_11695);
and U12111 (N_12111,N_11866,N_11608);
xnor U12112 (N_12112,N_11687,N_11754);
nand U12113 (N_12113,N_11970,N_11860);
nand U12114 (N_12114,N_11784,N_11876);
or U12115 (N_12115,N_11948,N_11878);
xor U12116 (N_12116,N_11988,N_11856);
or U12117 (N_12117,N_11655,N_11956);
nor U12118 (N_12118,N_11618,N_11877);
and U12119 (N_12119,N_11994,N_11704);
xnor U12120 (N_12120,N_11949,N_11801);
xor U12121 (N_12121,N_11666,N_11873);
nand U12122 (N_12122,N_11887,N_11814);
nand U12123 (N_12123,N_11773,N_11696);
and U12124 (N_12124,N_11946,N_11644);
or U12125 (N_12125,N_11933,N_11912);
or U12126 (N_12126,N_11619,N_11945);
and U12127 (N_12127,N_11864,N_11708);
or U12128 (N_12128,N_11643,N_11677);
and U12129 (N_12129,N_11701,N_11959);
nand U12130 (N_12130,N_11901,N_11746);
nor U12131 (N_12131,N_11951,N_11848);
or U12132 (N_12132,N_11973,N_11639);
xnor U12133 (N_12133,N_11661,N_11698);
nand U12134 (N_12134,N_11721,N_11606);
xor U12135 (N_12135,N_11842,N_11777);
and U12136 (N_12136,N_11749,N_11703);
and U12137 (N_12137,N_11760,N_11809);
nand U12138 (N_12138,N_11667,N_11984);
xnor U12139 (N_12139,N_11838,N_11600);
nand U12140 (N_12140,N_11967,N_11869);
xor U12141 (N_12141,N_11779,N_11772);
or U12142 (N_12142,N_11660,N_11752);
or U12143 (N_12143,N_11975,N_11682);
nor U12144 (N_12144,N_11742,N_11920);
nand U12145 (N_12145,N_11980,N_11705);
nand U12146 (N_12146,N_11974,N_11684);
and U12147 (N_12147,N_11692,N_11955);
nor U12148 (N_12148,N_11826,N_11714);
nor U12149 (N_12149,N_11612,N_11811);
and U12150 (N_12150,N_11733,N_11758);
or U12151 (N_12151,N_11849,N_11922);
xnor U12152 (N_12152,N_11782,N_11646);
nand U12153 (N_12153,N_11664,N_11839);
and U12154 (N_12154,N_11622,N_11895);
xor U12155 (N_12155,N_11686,N_11636);
or U12156 (N_12156,N_11943,N_11800);
and U12157 (N_12157,N_11917,N_11700);
and U12158 (N_12158,N_11889,N_11964);
nor U12159 (N_12159,N_11993,N_11944);
nor U12160 (N_12160,N_11712,N_11978);
nor U12161 (N_12161,N_11929,N_11659);
nor U12162 (N_12162,N_11727,N_11995);
and U12163 (N_12163,N_11824,N_11776);
xor U12164 (N_12164,N_11709,N_11678);
nand U12165 (N_12165,N_11751,N_11771);
nor U12166 (N_12166,N_11658,N_11833);
nor U12167 (N_12167,N_11892,N_11934);
nor U12168 (N_12168,N_11775,N_11863);
xnor U12169 (N_12169,N_11899,N_11938);
nand U12170 (N_12170,N_11766,N_11902);
nand U12171 (N_12171,N_11654,N_11605);
xnor U12172 (N_12172,N_11919,N_11836);
nand U12173 (N_12173,N_11638,N_11910);
and U12174 (N_12174,N_11762,N_11741);
nand U12175 (N_12175,N_11710,N_11653);
nand U12176 (N_12176,N_11663,N_11835);
xor U12177 (N_12177,N_11881,N_11888);
xnor U12178 (N_12178,N_11787,N_11822);
or U12179 (N_12179,N_11820,N_11651);
xor U12180 (N_12180,N_11841,N_11670);
nand U12181 (N_12181,N_11829,N_11986);
nand U12182 (N_12182,N_11676,N_11797);
or U12183 (N_12183,N_11807,N_11963);
xor U12184 (N_12184,N_11806,N_11621);
and U12185 (N_12185,N_11939,N_11624);
and U12186 (N_12186,N_11846,N_11805);
xor U12187 (N_12187,N_11623,N_11859);
nor U12188 (N_12188,N_11831,N_11958);
or U12189 (N_12189,N_11648,N_11680);
xnor U12190 (N_12190,N_11769,N_11688);
and U12191 (N_12191,N_11893,N_11872);
and U12192 (N_12192,N_11759,N_11941);
and U12193 (N_12193,N_11642,N_11633);
and U12194 (N_12194,N_11867,N_11930);
nor U12195 (N_12195,N_11793,N_11830);
xor U12196 (N_12196,N_11743,N_11834);
nand U12197 (N_12197,N_11735,N_11694);
or U12198 (N_12198,N_11999,N_11928);
nor U12199 (N_12199,N_11739,N_11847);
or U12200 (N_12200,N_11682,N_11605);
xnor U12201 (N_12201,N_11771,N_11990);
nand U12202 (N_12202,N_11793,N_11712);
nor U12203 (N_12203,N_11673,N_11615);
xor U12204 (N_12204,N_11737,N_11662);
nand U12205 (N_12205,N_11835,N_11803);
nand U12206 (N_12206,N_11915,N_11906);
and U12207 (N_12207,N_11749,N_11940);
xnor U12208 (N_12208,N_11783,N_11815);
nor U12209 (N_12209,N_11650,N_11860);
xnor U12210 (N_12210,N_11900,N_11665);
nor U12211 (N_12211,N_11914,N_11990);
and U12212 (N_12212,N_11745,N_11874);
nor U12213 (N_12213,N_11946,N_11936);
nor U12214 (N_12214,N_11827,N_11965);
nor U12215 (N_12215,N_11965,N_11867);
nand U12216 (N_12216,N_11746,N_11823);
nand U12217 (N_12217,N_11635,N_11888);
nand U12218 (N_12218,N_11801,N_11813);
nor U12219 (N_12219,N_11843,N_11711);
and U12220 (N_12220,N_11801,N_11824);
or U12221 (N_12221,N_11994,N_11821);
xnor U12222 (N_12222,N_11684,N_11871);
nand U12223 (N_12223,N_11868,N_11685);
xnor U12224 (N_12224,N_11647,N_11745);
or U12225 (N_12225,N_11919,N_11746);
nand U12226 (N_12226,N_11634,N_11731);
or U12227 (N_12227,N_11731,N_11996);
and U12228 (N_12228,N_11751,N_11621);
nand U12229 (N_12229,N_11847,N_11692);
xnor U12230 (N_12230,N_11939,N_11694);
or U12231 (N_12231,N_11727,N_11904);
nand U12232 (N_12232,N_11963,N_11670);
or U12233 (N_12233,N_11607,N_11952);
and U12234 (N_12234,N_11897,N_11920);
or U12235 (N_12235,N_11890,N_11808);
nor U12236 (N_12236,N_11743,N_11932);
and U12237 (N_12237,N_11921,N_11685);
and U12238 (N_12238,N_11625,N_11601);
and U12239 (N_12239,N_11898,N_11962);
xor U12240 (N_12240,N_11889,N_11603);
nand U12241 (N_12241,N_11955,N_11666);
xnor U12242 (N_12242,N_11682,N_11928);
nor U12243 (N_12243,N_11633,N_11704);
and U12244 (N_12244,N_11602,N_11643);
nand U12245 (N_12245,N_11679,N_11934);
or U12246 (N_12246,N_11757,N_11676);
nor U12247 (N_12247,N_11841,N_11788);
nand U12248 (N_12248,N_11956,N_11891);
nand U12249 (N_12249,N_11916,N_11698);
or U12250 (N_12250,N_11668,N_11968);
or U12251 (N_12251,N_11971,N_11730);
nand U12252 (N_12252,N_11703,N_11693);
xor U12253 (N_12253,N_11910,N_11908);
and U12254 (N_12254,N_11946,N_11721);
nor U12255 (N_12255,N_11916,N_11659);
xnor U12256 (N_12256,N_11601,N_11705);
and U12257 (N_12257,N_11889,N_11769);
nand U12258 (N_12258,N_11738,N_11999);
nor U12259 (N_12259,N_11663,N_11745);
nor U12260 (N_12260,N_11768,N_11862);
nand U12261 (N_12261,N_11911,N_11998);
or U12262 (N_12262,N_11618,N_11670);
and U12263 (N_12263,N_11953,N_11983);
and U12264 (N_12264,N_11645,N_11940);
or U12265 (N_12265,N_11963,N_11678);
xor U12266 (N_12266,N_11965,N_11893);
nand U12267 (N_12267,N_11701,N_11660);
nand U12268 (N_12268,N_11817,N_11785);
and U12269 (N_12269,N_11917,N_11775);
and U12270 (N_12270,N_11955,N_11663);
nand U12271 (N_12271,N_11893,N_11941);
or U12272 (N_12272,N_11816,N_11687);
or U12273 (N_12273,N_11701,N_11940);
and U12274 (N_12274,N_11630,N_11874);
xor U12275 (N_12275,N_11715,N_11921);
xnor U12276 (N_12276,N_11655,N_11619);
and U12277 (N_12277,N_11858,N_11957);
or U12278 (N_12278,N_11656,N_11869);
and U12279 (N_12279,N_11691,N_11645);
or U12280 (N_12280,N_11932,N_11817);
or U12281 (N_12281,N_11952,N_11872);
xor U12282 (N_12282,N_11816,N_11710);
or U12283 (N_12283,N_11934,N_11654);
and U12284 (N_12284,N_11877,N_11746);
and U12285 (N_12285,N_11628,N_11848);
and U12286 (N_12286,N_11908,N_11887);
xnor U12287 (N_12287,N_11602,N_11870);
or U12288 (N_12288,N_11944,N_11889);
and U12289 (N_12289,N_11985,N_11969);
nor U12290 (N_12290,N_11948,N_11678);
xnor U12291 (N_12291,N_11616,N_11652);
xnor U12292 (N_12292,N_11614,N_11611);
nor U12293 (N_12293,N_11717,N_11873);
and U12294 (N_12294,N_11816,N_11889);
xnor U12295 (N_12295,N_11656,N_11894);
nor U12296 (N_12296,N_11763,N_11968);
nand U12297 (N_12297,N_11666,N_11743);
and U12298 (N_12298,N_11689,N_11871);
and U12299 (N_12299,N_11992,N_11672);
nand U12300 (N_12300,N_11718,N_11769);
nor U12301 (N_12301,N_11833,N_11789);
or U12302 (N_12302,N_11730,N_11840);
nor U12303 (N_12303,N_11993,N_11941);
or U12304 (N_12304,N_11761,N_11782);
or U12305 (N_12305,N_11816,N_11602);
nand U12306 (N_12306,N_11916,N_11867);
or U12307 (N_12307,N_11949,N_11737);
nor U12308 (N_12308,N_11850,N_11629);
xnor U12309 (N_12309,N_11914,N_11779);
nor U12310 (N_12310,N_11890,N_11931);
nand U12311 (N_12311,N_11619,N_11707);
xnor U12312 (N_12312,N_11878,N_11867);
or U12313 (N_12313,N_11682,N_11755);
or U12314 (N_12314,N_11884,N_11808);
nand U12315 (N_12315,N_11746,N_11938);
nand U12316 (N_12316,N_11979,N_11704);
or U12317 (N_12317,N_11971,N_11624);
and U12318 (N_12318,N_11845,N_11700);
nand U12319 (N_12319,N_11900,N_11910);
nor U12320 (N_12320,N_11702,N_11833);
or U12321 (N_12321,N_11995,N_11676);
nor U12322 (N_12322,N_11973,N_11670);
nor U12323 (N_12323,N_11844,N_11714);
nor U12324 (N_12324,N_11669,N_11695);
nor U12325 (N_12325,N_11863,N_11664);
xnor U12326 (N_12326,N_11907,N_11749);
and U12327 (N_12327,N_11685,N_11934);
xnor U12328 (N_12328,N_11891,N_11986);
nand U12329 (N_12329,N_11685,N_11624);
nor U12330 (N_12330,N_11750,N_11705);
nor U12331 (N_12331,N_11822,N_11716);
xnor U12332 (N_12332,N_11997,N_11993);
xor U12333 (N_12333,N_11862,N_11696);
xor U12334 (N_12334,N_11808,N_11969);
and U12335 (N_12335,N_11733,N_11848);
xnor U12336 (N_12336,N_11724,N_11860);
xor U12337 (N_12337,N_11640,N_11621);
nor U12338 (N_12338,N_11737,N_11880);
nor U12339 (N_12339,N_11736,N_11977);
or U12340 (N_12340,N_11926,N_11769);
or U12341 (N_12341,N_11746,N_11611);
nor U12342 (N_12342,N_11980,N_11931);
xnor U12343 (N_12343,N_11676,N_11783);
and U12344 (N_12344,N_11652,N_11781);
nand U12345 (N_12345,N_11890,N_11876);
or U12346 (N_12346,N_11859,N_11608);
nor U12347 (N_12347,N_11938,N_11912);
nand U12348 (N_12348,N_11775,N_11673);
xor U12349 (N_12349,N_11761,N_11973);
or U12350 (N_12350,N_11908,N_11699);
and U12351 (N_12351,N_11742,N_11644);
and U12352 (N_12352,N_11685,N_11951);
nor U12353 (N_12353,N_11992,N_11656);
and U12354 (N_12354,N_11611,N_11643);
xnor U12355 (N_12355,N_11631,N_11824);
nand U12356 (N_12356,N_11771,N_11883);
and U12357 (N_12357,N_11710,N_11934);
xnor U12358 (N_12358,N_11708,N_11945);
and U12359 (N_12359,N_11817,N_11774);
and U12360 (N_12360,N_11997,N_11799);
or U12361 (N_12361,N_11856,N_11818);
nor U12362 (N_12362,N_11764,N_11953);
nor U12363 (N_12363,N_11716,N_11793);
nand U12364 (N_12364,N_11768,N_11758);
nor U12365 (N_12365,N_11786,N_11614);
xnor U12366 (N_12366,N_11859,N_11855);
nand U12367 (N_12367,N_11871,N_11686);
or U12368 (N_12368,N_11988,N_11725);
and U12369 (N_12369,N_11856,N_11755);
and U12370 (N_12370,N_11693,N_11879);
or U12371 (N_12371,N_11881,N_11781);
or U12372 (N_12372,N_11721,N_11959);
nor U12373 (N_12373,N_11886,N_11881);
nor U12374 (N_12374,N_11798,N_11887);
nand U12375 (N_12375,N_11859,N_11983);
nand U12376 (N_12376,N_11926,N_11951);
and U12377 (N_12377,N_11725,N_11938);
nor U12378 (N_12378,N_11931,N_11942);
or U12379 (N_12379,N_11685,N_11771);
or U12380 (N_12380,N_11666,N_11692);
nand U12381 (N_12381,N_11681,N_11932);
nand U12382 (N_12382,N_11752,N_11680);
or U12383 (N_12383,N_11783,N_11975);
nand U12384 (N_12384,N_11953,N_11688);
or U12385 (N_12385,N_11866,N_11625);
or U12386 (N_12386,N_11883,N_11744);
or U12387 (N_12387,N_11893,N_11878);
or U12388 (N_12388,N_11756,N_11632);
xnor U12389 (N_12389,N_11955,N_11772);
and U12390 (N_12390,N_11660,N_11976);
or U12391 (N_12391,N_11992,N_11860);
xor U12392 (N_12392,N_11834,N_11785);
or U12393 (N_12393,N_11851,N_11765);
nand U12394 (N_12394,N_11675,N_11833);
and U12395 (N_12395,N_11681,N_11827);
xor U12396 (N_12396,N_11835,N_11837);
and U12397 (N_12397,N_11722,N_11874);
nor U12398 (N_12398,N_11990,N_11819);
nor U12399 (N_12399,N_11673,N_11850);
and U12400 (N_12400,N_12339,N_12350);
and U12401 (N_12401,N_12148,N_12247);
xnor U12402 (N_12402,N_12143,N_12399);
or U12403 (N_12403,N_12056,N_12286);
xnor U12404 (N_12404,N_12235,N_12153);
nand U12405 (N_12405,N_12150,N_12037);
nor U12406 (N_12406,N_12346,N_12043);
and U12407 (N_12407,N_12135,N_12053);
nor U12408 (N_12408,N_12371,N_12079);
xor U12409 (N_12409,N_12106,N_12035);
xor U12410 (N_12410,N_12029,N_12131);
or U12411 (N_12411,N_12267,N_12138);
xor U12412 (N_12412,N_12326,N_12117);
or U12413 (N_12413,N_12128,N_12384);
and U12414 (N_12414,N_12118,N_12170);
xnor U12415 (N_12415,N_12007,N_12041);
nand U12416 (N_12416,N_12217,N_12026);
nand U12417 (N_12417,N_12008,N_12067);
and U12418 (N_12418,N_12299,N_12162);
nor U12419 (N_12419,N_12264,N_12307);
or U12420 (N_12420,N_12182,N_12277);
or U12421 (N_12421,N_12000,N_12179);
xor U12422 (N_12422,N_12266,N_12392);
xor U12423 (N_12423,N_12361,N_12057);
and U12424 (N_12424,N_12039,N_12227);
xor U12425 (N_12425,N_12362,N_12329);
and U12426 (N_12426,N_12136,N_12382);
xor U12427 (N_12427,N_12220,N_12322);
nand U12428 (N_12428,N_12111,N_12042);
nand U12429 (N_12429,N_12281,N_12199);
and U12430 (N_12430,N_12192,N_12188);
nor U12431 (N_12431,N_12107,N_12250);
nand U12432 (N_12432,N_12103,N_12232);
xor U12433 (N_12433,N_12157,N_12300);
nor U12434 (N_12434,N_12075,N_12085);
nand U12435 (N_12435,N_12115,N_12330);
nor U12436 (N_12436,N_12314,N_12102);
or U12437 (N_12437,N_12292,N_12032);
and U12438 (N_12438,N_12351,N_12325);
and U12439 (N_12439,N_12181,N_12210);
or U12440 (N_12440,N_12254,N_12205);
or U12441 (N_12441,N_12175,N_12271);
nor U12442 (N_12442,N_12078,N_12347);
xor U12443 (N_12443,N_12069,N_12064);
or U12444 (N_12444,N_12087,N_12386);
xor U12445 (N_12445,N_12076,N_12296);
nor U12446 (N_12446,N_12302,N_12385);
xor U12447 (N_12447,N_12327,N_12173);
nor U12448 (N_12448,N_12212,N_12383);
or U12449 (N_12449,N_12003,N_12354);
or U12450 (N_12450,N_12391,N_12313);
or U12451 (N_12451,N_12185,N_12348);
or U12452 (N_12452,N_12082,N_12092);
nor U12453 (N_12453,N_12015,N_12163);
nor U12454 (N_12454,N_12013,N_12226);
xnor U12455 (N_12455,N_12114,N_12086);
xor U12456 (N_12456,N_12344,N_12225);
or U12457 (N_12457,N_12331,N_12309);
or U12458 (N_12458,N_12071,N_12018);
or U12459 (N_12459,N_12252,N_12228);
or U12460 (N_12460,N_12245,N_12258);
nand U12461 (N_12461,N_12262,N_12219);
nand U12462 (N_12462,N_12398,N_12378);
xor U12463 (N_12463,N_12184,N_12036);
or U12464 (N_12464,N_12001,N_12390);
nand U12465 (N_12465,N_12012,N_12165);
and U12466 (N_12466,N_12233,N_12388);
nor U12467 (N_12467,N_12169,N_12268);
nor U12468 (N_12468,N_12062,N_12146);
xnor U12469 (N_12469,N_12260,N_12206);
nor U12470 (N_12470,N_12202,N_12280);
nor U12471 (N_12471,N_12224,N_12288);
nor U12472 (N_12472,N_12019,N_12108);
nor U12473 (N_12473,N_12272,N_12270);
xor U12474 (N_12474,N_12174,N_12316);
and U12475 (N_12475,N_12073,N_12360);
and U12476 (N_12476,N_12077,N_12010);
or U12477 (N_12477,N_12089,N_12161);
nand U12478 (N_12478,N_12207,N_12093);
and U12479 (N_12479,N_12095,N_12023);
nor U12480 (N_12480,N_12060,N_12369);
nor U12481 (N_12481,N_12144,N_12194);
and U12482 (N_12482,N_12024,N_12047);
and U12483 (N_12483,N_12241,N_12176);
nor U12484 (N_12484,N_12234,N_12155);
nor U12485 (N_12485,N_12223,N_12028);
xnor U12486 (N_12486,N_12290,N_12249);
nand U12487 (N_12487,N_12246,N_12049);
or U12488 (N_12488,N_12372,N_12259);
and U12489 (N_12489,N_12311,N_12198);
nor U12490 (N_12490,N_12341,N_12335);
or U12491 (N_12491,N_12139,N_12231);
or U12492 (N_12492,N_12213,N_12381);
nor U12493 (N_12493,N_12253,N_12190);
nand U12494 (N_12494,N_12125,N_12183);
nor U12495 (N_12495,N_12298,N_12303);
nor U12496 (N_12496,N_12321,N_12261);
or U12497 (N_12497,N_12284,N_12195);
nor U12498 (N_12498,N_12317,N_12011);
nand U12499 (N_12499,N_12145,N_12373);
and U12500 (N_12500,N_12178,N_12294);
and U12501 (N_12501,N_12243,N_12209);
or U12502 (N_12502,N_12295,N_12230);
nand U12503 (N_12503,N_12091,N_12034);
nand U12504 (N_12504,N_12353,N_12142);
nor U12505 (N_12505,N_12127,N_12364);
or U12506 (N_12506,N_12248,N_12375);
nand U12507 (N_12507,N_12074,N_12070);
or U12508 (N_12508,N_12025,N_12002);
nand U12509 (N_12509,N_12265,N_12164);
or U12510 (N_12510,N_12200,N_12216);
xor U12511 (N_12511,N_12120,N_12318);
nor U12512 (N_12512,N_12044,N_12154);
or U12513 (N_12513,N_12357,N_12061);
nand U12514 (N_12514,N_12275,N_12149);
nand U12515 (N_12515,N_12126,N_12158);
xor U12516 (N_12516,N_12359,N_12196);
and U12517 (N_12517,N_12203,N_12097);
and U12518 (N_12518,N_12285,N_12104);
or U12519 (N_12519,N_12387,N_12063);
nand U12520 (N_12520,N_12276,N_12094);
and U12521 (N_12521,N_12160,N_12096);
nand U12522 (N_12522,N_12394,N_12211);
or U12523 (N_12523,N_12137,N_12374);
nor U12524 (N_12524,N_12050,N_12167);
xor U12525 (N_12525,N_12263,N_12279);
nor U12526 (N_12526,N_12177,N_12052);
nor U12527 (N_12527,N_12308,N_12014);
xor U12528 (N_12528,N_12201,N_12187);
or U12529 (N_12529,N_12365,N_12324);
xor U12530 (N_12530,N_12040,N_12191);
nand U12531 (N_12531,N_12215,N_12134);
nand U12532 (N_12532,N_12081,N_12363);
xnor U12533 (N_12533,N_12343,N_12328);
nor U12534 (N_12534,N_12033,N_12389);
nor U12535 (N_12535,N_12278,N_12379);
nand U12536 (N_12536,N_12315,N_12274);
nor U12537 (N_12537,N_12323,N_12340);
or U12538 (N_12538,N_12204,N_12214);
and U12539 (N_12539,N_12171,N_12397);
or U12540 (N_12540,N_12306,N_12240);
or U12541 (N_12541,N_12244,N_12159);
nor U12542 (N_12542,N_12345,N_12312);
xnor U12543 (N_12543,N_12380,N_12109);
xnor U12544 (N_12544,N_12256,N_12046);
xor U12545 (N_12545,N_12016,N_12186);
xor U12546 (N_12546,N_12297,N_12273);
xnor U12547 (N_12547,N_12080,N_12289);
xor U12548 (N_12548,N_12006,N_12320);
or U12549 (N_12549,N_12342,N_12237);
and U12550 (N_12550,N_12366,N_12238);
nand U12551 (N_12551,N_12110,N_12090);
and U12552 (N_12552,N_12377,N_12055);
nand U12553 (N_12553,N_12287,N_12132);
and U12554 (N_12554,N_12283,N_12368);
nor U12555 (N_12555,N_12156,N_12239);
and U12556 (N_12556,N_12084,N_12152);
nor U12557 (N_12557,N_12083,N_12255);
and U12558 (N_12558,N_12101,N_12395);
nand U12559 (N_12559,N_12349,N_12310);
and U12560 (N_12560,N_12133,N_12021);
nand U12561 (N_12561,N_12121,N_12269);
nand U12562 (N_12562,N_12236,N_12242);
nand U12563 (N_12563,N_12396,N_12337);
nor U12564 (N_12564,N_12058,N_12022);
or U12565 (N_12565,N_12304,N_12367);
xnor U12566 (N_12566,N_12122,N_12119);
nand U12567 (N_12567,N_12113,N_12229);
or U12568 (N_12568,N_12336,N_12293);
and U12569 (N_12569,N_12051,N_12112);
xor U12570 (N_12570,N_12065,N_12370);
and U12571 (N_12571,N_12072,N_12116);
and U12572 (N_12572,N_12088,N_12393);
or U12573 (N_12573,N_12100,N_12105);
nand U12574 (N_12574,N_12166,N_12301);
xor U12575 (N_12575,N_12291,N_12358);
and U12576 (N_12576,N_12045,N_12352);
xor U12577 (N_12577,N_12004,N_12319);
nor U12578 (N_12578,N_12027,N_12066);
nor U12579 (N_12579,N_12005,N_12030);
nand U12580 (N_12580,N_12098,N_12130);
or U12581 (N_12581,N_12257,N_12189);
or U12582 (N_12582,N_12282,N_12208);
nand U12583 (N_12583,N_12356,N_12222);
or U12584 (N_12584,N_12338,N_12168);
nand U12585 (N_12585,N_12151,N_12197);
and U12586 (N_12586,N_12172,N_12376);
nand U12587 (N_12587,N_12020,N_12334);
nor U12588 (N_12588,N_12140,N_12333);
nand U12589 (N_12589,N_12332,N_12068);
and U12590 (N_12590,N_12099,N_12305);
or U12591 (N_12591,N_12129,N_12355);
nor U12592 (N_12592,N_12221,N_12180);
or U12593 (N_12593,N_12251,N_12017);
or U12594 (N_12594,N_12031,N_12141);
nand U12595 (N_12595,N_12048,N_12123);
nor U12596 (N_12596,N_12059,N_12038);
or U12597 (N_12597,N_12009,N_12147);
or U12598 (N_12598,N_12218,N_12054);
and U12599 (N_12599,N_12124,N_12193);
nand U12600 (N_12600,N_12078,N_12062);
and U12601 (N_12601,N_12197,N_12115);
xor U12602 (N_12602,N_12092,N_12085);
nand U12603 (N_12603,N_12344,N_12294);
nand U12604 (N_12604,N_12399,N_12185);
or U12605 (N_12605,N_12214,N_12083);
or U12606 (N_12606,N_12362,N_12052);
or U12607 (N_12607,N_12238,N_12061);
and U12608 (N_12608,N_12026,N_12175);
nor U12609 (N_12609,N_12280,N_12357);
xnor U12610 (N_12610,N_12214,N_12376);
or U12611 (N_12611,N_12314,N_12008);
nand U12612 (N_12612,N_12110,N_12375);
nor U12613 (N_12613,N_12135,N_12018);
xor U12614 (N_12614,N_12154,N_12354);
xnor U12615 (N_12615,N_12103,N_12177);
xor U12616 (N_12616,N_12291,N_12036);
or U12617 (N_12617,N_12096,N_12094);
nand U12618 (N_12618,N_12227,N_12035);
or U12619 (N_12619,N_12247,N_12299);
and U12620 (N_12620,N_12042,N_12235);
xor U12621 (N_12621,N_12384,N_12347);
nand U12622 (N_12622,N_12208,N_12388);
or U12623 (N_12623,N_12197,N_12052);
nor U12624 (N_12624,N_12304,N_12243);
and U12625 (N_12625,N_12282,N_12111);
nand U12626 (N_12626,N_12325,N_12373);
nand U12627 (N_12627,N_12241,N_12117);
nor U12628 (N_12628,N_12154,N_12386);
nand U12629 (N_12629,N_12193,N_12132);
nor U12630 (N_12630,N_12067,N_12249);
or U12631 (N_12631,N_12180,N_12214);
and U12632 (N_12632,N_12307,N_12348);
or U12633 (N_12633,N_12203,N_12020);
nor U12634 (N_12634,N_12011,N_12149);
or U12635 (N_12635,N_12126,N_12128);
or U12636 (N_12636,N_12333,N_12256);
nor U12637 (N_12637,N_12316,N_12009);
or U12638 (N_12638,N_12361,N_12375);
xnor U12639 (N_12639,N_12357,N_12339);
xor U12640 (N_12640,N_12182,N_12252);
or U12641 (N_12641,N_12141,N_12208);
and U12642 (N_12642,N_12317,N_12253);
or U12643 (N_12643,N_12141,N_12043);
xnor U12644 (N_12644,N_12219,N_12096);
xnor U12645 (N_12645,N_12250,N_12220);
or U12646 (N_12646,N_12066,N_12098);
or U12647 (N_12647,N_12116,N_12099);
xor U12648 (N_12648,N_12156,N_12040);
nand U12649 (N_12649,N_12257,N_12284);
nor U12650 (N_12650,N_12154,N_12116);
xnor U12651 (N_12651,N_12035,N_12188);
or U12652 (N_12652,N_12030,N_12047);
or U12653 (N_12653,N_12369,N_12324);
and U12654 (N_12654,N_12174,N_12279);
and U12655 (N_12655,N_12114,N_12395);
nand U12656 (N_12656,N_12381,N_12234);
xor U12657 (N_12657,N_12171,N_12386);
and U12658 (N_12658,N_12321,N_12097);
xnor U12659 (N_12659,N_12018,N_12307);
nand U12660 (N_12660,N_12080,N_12144);
nand U12661 (N_12661,N_12009,N_12380);
xor U12662 (N_12662,N_12204,N_12093);
xnor U12663 (N_12663,N_12001,N_12033);
xnor U12664 (N_12664,N_12056,N_12084);
nor U12665 (N_12665,N_12327,N_12168);
nor U12666 (N_12666,N_12038,N_12384);
or U12667 (N_12667,N_12356,N_12121);
and U12668 (N_12668,N_12280,N_12362);
and U12669 (N_12669,N_12111,N_12137);
xor U12670 (N_12670,N_12369,N_12138);
xor U12671 (N_12671,N_12211,N_12129);
and U12672 (N_12672,N_12272,N_12202);
nand U12673 (N_12673,N_12368,N_12277);
nand U12674 (N_12674,N_12273,N_12244);
or U12675 (N_12675,N_12322,N_12166);
and U12676 (N_12676,N_12159,N_12114);
nor U12677 (N_12677,N_12246,N_12174);
or U12678 (N_12678,N_12110,N_12392);
nand U12679 (N_12679,N_12291,N_12278);
xor U12680 (N_12680,N_12101,N_12169);
or U12681 (N_12681,N_12094,N_12231);
nand U12682 (N_12682,N_12085,N_12005);
xnor U12683 (N_12683,N_12348,N_12073);
and U12684 (N_12684,N_12199,N_12161);
xor U12685 (N_12685,N_12076,N_12063);
or U12686 (N_12686,N_12105,N_12377);
nor U12687 (N_12687,N_12346,N_12263);
or U12688 (N_12688,N_12298,N_12141);
or U12689 (N_12689,N_12000,N_12097);
and U12690 (N_12690,N_12322,N_12117);
xnor U12691 (N_12691,N_12080,N_12069);
and U12692 (N_12692,N_12028,N_12316);
and U12693 (N_12693,N_12322,N_12134);
xnor U12694 (N_12694,N_12036,N_12220);
nor U12695 (N_12695,N_12120,N_12383);
nand U12696 (N_12696,N_12081,N_12385);
nor U12697 (N_12697,N_12007,N_12229);
or U12698 (N_12698,N_12142,N_12187);
and U12699 (N_12699,N_12115,N_12123);
nand U12700 (N_12700,N_12277,N_12012);
and U12701 (N_12701,N_12211,N_12167);
nor U12702 (N_12702,N_12376,N_12333);
xor U12703 (N_12703,N_12178,N_12390);
and U12704 (N_12704,N_12357,N_12177);
xor U12705 (N_12705,N_12202,N_12376);
nor U12706 (N_12706,N_12048,N_12169);
or U12707 (N_12707,N_12080,N_12093);
nor U12708 (N_12708,N_12223,N_12107);
nor U12709 (N_12709,N_12114,N_12099);
and U12710 (N_12710,N_12354,N_12089);
and U12711 (N_12711,N_12298,N_12045);
or U12712 (N_12712,N_12137,N_12274);
xor U12713 (N_12713,N_12054,N_12354);
and U12714 (N_12714,N_12286,N_12068);
nor U12715 (N_12715,N_12275,N_12276);
and U12716 (N_12716,N_12167,N_12288);
or U12717 (N_12717,N_12072,N_12296);
nand U12718 (N_12718,N_12137,N_12268);
xnor U12719 (N_12719,N_12343,N_12302);
nor U12720 (N_12720,N_12023,N_12185);
or U12721 (N_12721,N_12020,N_12048);
xor U12722 (N_12722,N_12102,N_12208);
xor U12723 (N_12723,N_12318,N_12132);
nand U12724 (N_12724,N_12102,N_12210);
or U12725 (N_12725,N_12159,N_12397);
nand U12726 (N_12726,N_12169,N_12373);
nor U12727 (N_12727,N_12163,N_12216);
nor U12728 (N_12728,N_12106,N_12043);
or U12729 (N_12729,N_12175,N_12282);
xor U12730 (N_12730,N_12029,N_12233);
or U12731 (N_12731,N_12213,N_12388);
nand U12732 (N_12732,N_12179,N_12019);
and U12733 (N_12733,N_12208,N_12015);
or U12734 (N_12734,N_12012,N_12181);
and U12735 (N_12735,N_12168,N_12365);
xor U12736 (N_12736,N_12380,N_12357);
and U12737 (N_12737,N_12031,N_12054);
or U12738 (N_12738,N_12251,N_12009);
or U12739 (N_12739,N_12012,N_12066);
and U12740 (N_12740,N_12052,N_12260);
or U12741 (N_12741,N_12034,N_12051);
xnor U12742 (N_12742,N_12016,N_12337);
nand U12743 (N_12743,N_12059,N_12332);
or U12744 (N_12744,N_12397,N_12200);
xnor U12745 (N_12745,N_12293,N_12364);
or U12746 (N_12746,N_12397,N_12348);
nand U12747 (N_12747,N_12252,N_12314);
xnor U12748 (N_12748,N_12152,N_12180);
xnor U12749 (N_12749,N_12056,N_12159);
xor U12750 (N_12750,N_12074,N_12094);
xor U12751 (N_12751,N_12020,N_12258);
and U12752 (N_12752,N_12164,N_12222);
xor U12753 (N_12753,N_12246,N_12164);
or U12754 (N_12754,N_12182,N_12218);
nand U12755 (N_12755,N_12114,N_12140);
nand U12756 (N_12756,N_12116,N_12212);
nand U12757 (N_12757,N_12215,N_12068);
or U12758 (N_12758,N_12042,N_12095);
or U12759 (N_12759,N_12097,N_12324);
and U12760 (N_12760,N_12372,N_12183);
xor U12761 (N_12761,N_12277,N_12188);
xor U12762 (N_12762,N_12177,N_12188);
nor U12763 (N_12763,N_12053,N_12064);
and U12764 (N_12764,N_12232,N_12035);
and U12765 (N_12765,N_12109,N_12030);
xnor U12766 (N_12766,N_12199,N_12219);
and U12767 (N_12767,N_12358,N_12164);
and U12768 (N_12768,N_12006,N_12280);
nor U12769 (N_12769,N_12024,N_12209);
or U12770 (N_12770,N_12038,N_12023);
nand U12771 (N_12771,N_12323,N_12373);
or U12772 (N_12772,N_12370,N_12173);
and U12773 (N_12773,N_12379,N_12151);
nand U12774 (N_12774,N_12201,N_12290);
nand U12775 (N_12775,N_12269,N_12258);
nand U12776 (N_12776,N_12112,N_12029);
nand U12777 (N_12777,N_12023,N_12186);
xor U12778 (N_12778,N_12041,N_12087);
xnor U12779 (N_12779,N_12295,N_12053);
or U12780 (N_12780,N_12185,N_12320);
and U12781 (N_12781,N_12285,N_12086);
nor U12782 (N_12782,N_12099,N_12146);
and U12783 (N_12783,N_12280,N_12353);
xor U12784 (N_12784,N_12197,N_12154);
or U12785 (N_12785,N_12140,N_12349);
or U12786 (N_12786,N_12095,N_12163);
and U12787 (N_12787,N_12298,N_12059);
or U12788 (N_12788,N_12079,N_12319);
nor U12789 (N_12789,N_12191,N_12131);
nor U12790 (N_12790,N_12102,N_12180);
and U12791 (N_12791,N_12351,N_12314);
nand U12792 (N_12792,N_12316,N_12265);
nand U12793 (N_12793,N_12030,N_12018);
nor U12794 (N_12794,N_12396,N_12036);
xnor U12795 (N_12795,N_12158,N_12043);
xnor U12796 (N_12796,N_12318,N_12354);
nand U12797 (N_12797,N_12370,N_12013);
nand U12798 (N_12798,N_12344,N_12064);
nand U12799 (N_12799,N_12250,N_12222);
nor U12800 (N_12800,N_12746,N_12596);
nand U12801 (N_12801,N_12646,N_12573);
nor U12802 (N_12802,N_12575,N_12693);
nor U12803 (N_12803,N_12579,N_12439);
xor U12804 (N_12804,N_12773,N_12780);
nand U12805 (N_12805,N_12584,N_12753);
xnor U12806 (N_12806,N_12466,N_12588);
xor U12807 (N_12807,N_12651,N_12440);
nand U12808 (N_12808,N_12473,N_12770);
and U12809 (N_12809,N_12538,N_12748);
nor U12810 (N_12810,N_12406,N_12716);
xnor U12811 (N_12811,N_12593,N_12709);
xnor U12812 (N_12812,N_12465,N_12551);
xor U12813 (N_12813,N_12694,N_12408);
and U12814 (N_12814,N_12454,N_12720);
or U12815 (N_12815,N_12699,N_12405);
nand U12816 (N_12816,N_12497,N_12647);
or U12817 (N_12817,N_12479,N_12796);
nand U12818 (N_12818,N_12562,N_12578);
nand U12819 (N_12819,N_12704,N_12754);
and U12820 (N_12820,N_12603,N_12416);
nor U12821 (N_12821,N_12652,N_12536);
xor U12822 (N_12822,N_12418,N_12555);
and U12823 (N_12823,N_12580,N_12758);
and U12824 (N_12824,N_12427,N_12494);
and U12825 (N_12825,N_12400,N_12790);
xor U12826 (N_12826,N_12544,N_12769);
xnor U12827 (N_12827,N_12657,N_12730);
or U12828 (N_12828,N_12421,N_12686);
and U12829 (N_12829,N_12673,N_12464);
nand U12830 (N_12830,N_12715,N_12508);
nor U12831 (N_12831,N_12460,N_12581);
nor U12832 (N_12832,N_12543,N_12455);
xor U12833 (N_12833,N_12449,N_12711);
nand U12834 (N_12834,N_12582,N_12425);
nand U12835 (N_12835,N_12710,N_12437);
nor U12836 (N_12836,N_12597,N_12432);
nand U12837 (N_12837,N_12447,N_12637);
nor U12838 (N_12838,N_12500,N_12781);
nand U12839 (N_12839,N_12535,N_12409);
xor U12840 (N_12840,N_12797,N_12613);
and U12841 (N_12841,N_12752,N_12666);
and U12842 (N_12842,N_12412,N_12749);
and U12843 (N_12843,N_12481,N_12532);
or U12844 (N_12844,N_12482,N_12677);
or U12845 (N_12845,N_12629,N_12772);
xnor U12846 (N_12846,N_12734,N_12798);
nand U12847 (N_12847,N_12702,N_12624);
nand U12848 (N_12848,N_12736,N_12788);
xor U12849 (N_12849,N_12552,N_12679);
or U12850 (N_12850,N_12598,N_12442);
nand U12851 (N_12851,N_12470,N_12766);
or U12852 (N_12852,N_12478,N_12712);
xor U12853 (N_12853,N_12518,N_12407);
and U12854 (N_12854,N_12533,N_12743);
or U12855 (N_12855,N_12641,N_12690);
nand U12856 (N_12856,N_12682,N_12531);
or U12857 (N_12857,N_12521,N_12695);
nand U12858 (N_12858,N_12502,N_12496);
nor U12859 (N_12859,N_12608,N_12491);
and U12860 (N_12860,N_12745,N_12461);
or U12861 (N_12861,N_12669,N_12763);
and U12862 (N_12862,N_12643,N_12732);
and U12863 (N_12863,N_12495,N_12723);
or U12864 (N_12864,N_12751,N_12403);
and U12865 (N_12865,N_12504,N_12477);
xnor U12866 (N_12866,N_12565,N_12660);
nand U12867 (N_12867,N_12675,N_12556);
nor U12868 (N_12868,N_12762,N_12576);
and U12869 (N_12869,N_12501,N_12661);
xnor U12870 (N_12870,N_12512,N_12431);
and U12871 (N_12871,N_12618,N_12450);
xnor U12872 (N_12872,N_12413,N_12714);
xor U12873 (N_12873,N_12719,N_12701);
nand U12874 (N_12874,N_12786,N_12606);
xnor U12875 (N_12875,N_12604,N_12795);
xor U12876 (N_12876,N_12537,N_12724);
xor U12877 (N_12877,N_12778,N_12735);
xor U12878 (N_12878,N_12612,N_12767);
xor U12879 (N_12879,N_12434,N_12506);
nor U12880 (N_12880,N_12609,N_12415);
and U12881 (N_12881,N_12728,N_12436);
or U12882 (N_12882,N_12451,N_12667);
xor U12883 (N_12883,N_12605,N_12642);
xor U12884 (N_12884,N_12463,N_12511);
and U12885 (N_12885,N_12446,N_12600);
or U12886 (N_12886,N_12785,N_12731);
and U12887 (N_12887,N_12665,N_12692);
nor U12888 (N_12888,N_12622,N_12649);
nor U12889 (N_12889,N_12632,N_12586);
xnor U12890 (N_12890,N_12727,N_12640);
or U12891 (N_12891,N_12420,N_12475);
or U12892 (N_12892,N_12700,N_12733);
or U12893 (N_12893,N_12678,N_12570);
and U12894 (N_12894,N_12611,N_12591);
xnor U12895 (N_12895,N_12659,N_12545);
nor U12896 (N_12896,N_12505,N_12784);
xnor U12897 (N_12897,N_12410,N_12487);
nor U12898 (N_12898,N_12423,N_12468);
nand U12899 (N_12899,N_12697,N_12779);
nor U12900 (N_12900,N_12787,N_12634);
xnor U12901 (N_12901,N_12486,N_12499);
or U12902 (N_12902,N_12539,N_12590);
xor U12903 (N_12903,N_12703,N_12617);
and U12904 (N_12904,N_12404,N_12757);
xnor U12905 (N_12905,N_12483,N_12515);
and U12906 (N_12906,N_12509,N_12644);
xnor U12907 (N_12907,N_12658,N_12696);
nand U12908 (N_12908,N_12650,N_12639);
or U12909 (N_12909,N_12592,N_12526);
nand U12910 (N_12910,N_12474,N_12636);
or U12911 (N_12911,N_12540,N_12589);
or U12912 (N_12912,N_12534,N_12510);
xnor U12913 (N_12913,N_12574,N_12523);
and U12914 (N_12914,N_12623,N_12648);
or U12915 (N_12915,N_12519,N_12681);
nor U12916 (N_12916,N_12616,N_12627);
xor U12917 (N_12917,N_12443,N_12654);
nand U12918 (N_12918,N_12708,N_12670);
nor U12919 (N_12919,N_12656,N_12740);
or U12920 (N_12920,N_12774,N_12680);
nor U12921 (N_12921,N_12776,N_12467);
xnor U12922 (N_12922,N_12553,N_12633);
or U12923 (N_12923,N_12563,N_12718);
or U12924 (N_12924,N_12620,N_12583);
and U12925 (N_12925,N_12564,N_12530);
or U12926 (N_12926,N_12554,N_12765);
and U12927 (N_12927,N_12768,N_12602);
and U12928 (N_12928,N_12594,N_12655);
nor U12929 (N_12929,N_12422,N_12462);
nor U12930 (N_12930,N_12614,N_12668);
or U12931 (N_12931,N_12472,N_12717);
and U12932 (N_12932,N_12683,N_12610);
xnor U12933 (N_12933,N_12782,N_12527);
xor U12934 (N_12934,N_12448,N_12428);
xor U12935 (N_12935,N_12729,N_12503);
nor U12936 (N_12936,N_12663,N_12755);
nor U12937 (N_12937,N_12524,N_12764);
or U12938 (N_12938,N_12726,N_12548);
nand U12939 (N_12939,N_12571,N_12417);
nand U12940 (N_12940,N_12783,N_12684);
or U12941 (N_12941,N_12628,N_12747);
xor U12942 (N_12942,N_12713,N_12559);
xnor U12943 (N_12943,N_12799,N_12572);
and U12944 (N_12944,N_12471,N_12687);
and U12945 (N_12945,N_12426,N_12541);
nor U12946 (N_12946,N_12759,N_12607);
xor U12947 (N_12947,N_12685,N_12619);
xnor U12948 (N_12948,N_12793,N_12411);
nor U12949 (N_12949,N_12750,N_12676);
nand U12950 (N_12950,N_12469,N_12560);
nor U12951 (N_12951,N_12621,N_12631);
nand U12952 (N_12952,N_12688,N_12698);
nand U12953 (N_12953,N_12480,N_12485);
nand U12954 (N_12954,N_12438,N_12638);
and U12955 (N_12955,N_12626,N_12689);
or U12956 (N_12956,N_12528,N_12595);
and U12957 (N_12957,N_12792,N_12635);
xnor U12958 (N_12958,N_12671,N_12722);
nand U12959 (N_12959,N_12498,N_12741);
and U12960 (N_12960,N_12645,N_12569);
nor U12961 (N_12961,N_12705,N_12419);
or U12962 (N_12962,N_12615,N_12653);
and U12963 (N_12963,N_12529,N_12738);
nor U12964 (N_12964,N_12401,N_12547);
and U12965 (N_12965,N_12775,N_12585);
nand U12966 (N_12966,N_12546,N_12476);
nand U12967 (N_12967,N_12457,N_12549);
and U12968 (N_12968,N_12672,N_12459);
and U12969 (N_12969,N_12706,N_12525);
nand U12970 (N_12970,N_12568,N_12691);
nor U12971 (N_12971,N_12453,N_12517);
xnor U12972 (N_12972,N_12433,N_12761);
xor U12973 (N_12973,N_12489,N_12742);
or U12974 (N_12974,N_12513,N_12587);
nand U12975 (N_12975,N_12522,N_12542);
nand U12976 (N_12976,N_12760,N_12744);
or U12977 (N_12977,N_12777,N_12557);
or U12978 (N_12978,N_12445,N_12725);
nand U12979 (N_12979,N_12558,N_12625);
or U12980 (N_12980,N_12599,N_12550);
or U12981 (N_12981,N_12514,N_12456);
and U12982 (N_12982,N_12662,N_12424);
nand U12983 (N_12983,N_12520,N_12737);
or U12984 (N_12984,N_12435,N_12507);
xor U12985 (N_12985,N_12429,N_12561);
and U12986 (N_12986,N_12721,N_12493);
or U12987 (N_12987,N_12488,N_12452);
xor U12988 (N_12988,N_12791,N_12756);
nor U12989 (N_12989,N_12630,N_12441);
nor U12990 (N_12990,N_12674,N_12794);
and U12991 (N_12991,N_12444,N_12402);
xnor U12992 (N_12992,N_12516,N_12430);
nand U12993 (N_12993,N_12490,N_12707);
nor U12994 (N_12994,N_12414,N_12458);
and U12995 (N_12995,N_12771,N_12601);
xnor U12996 (N_12996,N_12739,N_12789);
xor U12997 (N_12997,N_12492,N_12577);
or U12998 (N_12998,N_12566,N_12567);
nand U12999 (N_12999,N_12484,N_12664);
nand U13000 (N_13000,N_12793,N_12556);
or U13001 (N_13001,N_12459,N_12620);
nor U13002 (N_13002,N_12731,N_12746);
xor U13003 (N_13003,N_12650,N_12730);
nand U13004 (N_13004,N_12555,N_12402);
or U13005 (N_13005,N_12740,N_12453);
nand U13006 (N_13006,N_12513,N_12736);
nor U13007 (N_13007,N_12667,N_12498);
nor U13008 (N_13008,N_12438,N_12554);
or U13009 (N_13009,N_12666,N_12465);
or U13010 (N_13010,N_12566,N_12694);
nor U13011 (N_13011,N_12692,N_12676);
xnor U13012 (N_13012,N_12554,N_12627);
xnor U13013 (N_13013,N_12614,N_12626);
nor U13014 (N_13014,N_12414,N_12694);
nand U13015 (N_13015,N_12741,N_12619);
nand U13016 (N_13016,N_12766,N_12731);
or U13017 (N_13017,N_12420,N_12744);
or U13018 (N_13018,N_12471,N_12549);
and U13019 (N_13019,N_12578,N_12746);
and U13020 (N_13020,N_12653,N_12464);
nand U13021 (N_13021,N_12587,N_12772);
nand U13022 (N_13022,N_12599,N_12464);
nand U13023 (N_13023,N_12713,N_12611);
or U13024 (N_13024,N_12761,N_12477);
nor U13025 (N_13025,N_12514,N_12543);
nand U13026 (N_13026,N_12440,N_12783);
or U13027 (N_13027,N_12763,N_12466);
nand U13028 (N_13028,N_12606,N_12575);
and U13029 (N_13029,N_12519,N_12567);
nand U13030 (N_13030,N_12485,N_12753);
or U13031 (N_13031,N_12532,N_12487);
nor U13032 (N_13032,N_12544,N_12543);
xnor U13033 (N_13033,N_12478,N_12785);
and U13034 (N_13034,N_12646,N_12783);
or U13035 (N_13035,N_12576,N_12545);
nand U13036 (N_13036,N_12779,N_12519);
and U13037 (N_13037,N_12695,N_12622);
nor U13038 (N_13038,N_12507,N_12735);
nor U13039 (N_13039,N_12778,N_12698);
nand U13040 (N_13040,N_12512,N_12792);
and U13041 (N_13041,N_12542,N_12575);
xor U13042 (N_13042,N_12588,N_12612);
and U13043 (N_13043,N_12677,N_12678);
or U13044 (N_13044,N_12703,N_12713);
and U13045 (N_13045,N_12431,N_12568);
xnor U13046 (N_13046,N_12694,N_12412);
and U13047 (N_13047,N_12793,N_12752);
nand U13048 (N_13048,N_12426,N_12754);
nand U13049 (N_13049,N_12516,N_12437);
or U13050 (N_13050,N_12628,N_12565);
xor U13051 (N_13051,N_12571,N_12757);
nor U13052 (N_13052,N_12690,N_12702);
and U13053 (N_13053,N_12426,N_12687);
nand U13054 (N_13054,N_12659,N_12671);
nand U13055 (N_13055,N_12556,N_12687);
or U13056 (N_13056,N_12400,N_12635);
and U13057 (N_13057,N_12535,N_12581);
nand U13058 (N_13058,N_12460,N_12663);
or U13059 (N_13059,N_12622,N_12464);
nor U13060 (N_13060,N_12738,N_12576);
nor U13061 (N_13061,N_12724,N_12719);
nand U13062 (N_13062,N_12777,N_12791);
xnor U13063 (N_13063,N_12630,N_12702);
xor U13064 (N_13064,N_12779,N_12676);
or U13065 (N_13065,N_12752,N_12463);
nor U13066 (N_13066,N_12763,N_12615);
nor U13067 (N_13067,N_12713,N_12670);
nor U13068 (N_13068,N_12615,N_12505);
nor U13069 (N_13069,N_12627,N_12733);
or U13070 (N_13070,N_12649,N_12693);
and U13071 (N_13071,N_12483,N_12731);
nor U13072 (N_13072,N_12797,N_12501);
or U13073 (N_13073,N_12747,N_12683);
nor U13074 (N_13074,N_12542,N_12780);
and U13075 (N_13075,N_12654,N_12667);
and U13076 (N_13076,N_12462,N_12436);
or U13077 (N_13077,N_12463,N_12617);
or U13078 (N_13078,N_12769,N_12570);
or U13079 (N_13079,N_12491,N_12674);
and U13080 (N_13080,N_12723,N_12646);
nor U13081 (N_13081,N_12655,N_12505);
nor U13082 (N_13082,N_12673,N_12609);
nand U13083 (N_13083,N_12604,N_12506);
nor U13084 (N_13084,N_12639,N_12604);
nand U13085 (N_13085,N_12761,N_12773);
and U13086 (N_13086,N_12598,N_12508);
and U13087 (N_13087,N_12460,N_12731);
and U13088 (N_13088,N_12587,N_12536);
nand U13089 (N_13089,N_12517,N_12602);
nand U13090 (N_13090,N_12696,N_12445);
xor U13091 (N_13091,N_12487,N_12585);
nand U13092 (N_13092,N_12640,N_12588);
xnor U13093 (N_13093,N_12477,N_12740);
nor U13094 (N_13094,N_12587,N_12550);
nand U13095 (N_13095,N_12744,N_12587);
nand U13096 (N_13096,N_12734,N_12669);
nor U13097 (N_13097,N_12680,N_12400);
nand U13098 (N_13098,N_12729,N_12455);
nand U13099 (N_13099,N_12442,N_12623);
nor U13100 (N_13100,N_12422,N_12418);
xor U13101 (N_13101,N_12516,N_12543);
and U13102 (N_13102,N_12736,N_12477);
xor U13103 (N_13103,N_12722,N_12524);
or U13104 (N_13104,N_12599,N_12734);
nand U13105 (N_13105,N_12538,N_12548);
and U13106 (N_13106,N_12678,N_12627);
nor U13107 (N_13107,N_12470,N_12625);
nand U13108 (N_13108,N_12515,N_12488);
or U13109 (N_13109,N_12569,N_12673);
nor U13110 (N_13110,N_12794,N_12479);
and U13111 (N_13111,N_12708,N_12523);
xor U13112 (N_13112,N_12413,N_12725);
or U13113 (N_13113,N_12448,N_12647);
or U13114 (N_13114,N_12565,N_12650);
xor U13115 (N_13115,N_12673,N_12699);
nand U13116 (N_13116,N_12655,N_12578);
nand U13117 (N_13117,N_12573,N_12432);
and U13118 (N_13118,N_12689,N_12677);
and U13119 (N_13119,N_12646,N_12492);
xnor U13120 (N_13120,N_12401,N_12473);
or U13121 (N_13121,N_12423,N_12527);
nand U13122 (N_13122,N_12694,N_12542);
nand U13123 (N_13123,N_12781,N_12732);
or U13124 (N_13124,N_12732,N_12535);
nand U13125 (N_13125,N_12662,N_12784);
or U13126 (N_13126,N_12588,N_12733);
or U13127 (N_13127,N_12496,N_12469);
xor U13128 (N_13128,N_12464,N_12444);
or U13129 (N_13129,N_12785,N_12627);
nand U13130 (N_13130,N_12697,N_12530);
xor U13131 (N_13131,N_12528,N_12772);
xor U13132 (N_13132,N_12732,N_12756);
nor U13133 (N_13133,N_12730,N_12723);
nor U13134 (N_13134,N_12795,N_12585);
nor U13135 (N_13135,N_12693,N_12494);
or U13136 (N_13136,N_12490,N_12436);
and U13137 (N_13137,N_12479,N_12675);
nor U13138 (N_13138,N_12508,N_12591);
xor U13139 (N_13139,N_12623,N_12505);
and U13140 (N_13140,N_12777,N_12768);
and U13141 (N_13141,N_12622,N_12582);
and U13142 (N_13142,N_12553,N_12799);
and U13143 (N_13143,N_12685,N_12491);
or U13144 (N_13144,N_12534,N_12573);
xor U13145 (N_13145,N_12715,N_12667);
nand U13146 (N_13146,N_12690,N_12741);
nor U13147 (N_13147,N_12678,N_12411);
or U13148 (N_13148,N_12400,N_12606);
nor U13149 (N_13149,N_12429,N_12784);
nor U13150 (N_13150,N_12628,N_12798);
or U13151 (N_13151,N_12670,N_12781);
xnor U13152 (N_13152,N_12741,N_12780);
xnor U13153 (N_13153,N_12601,N_12529);
or U13154 (N_13154,N_12579,N_12471);
and U13155 (N_13155,N_12697,N_12474);
xnor U13156 (N_13156,N_12502,N_12553);
and U13157 (N_13157,N_12762,N_12713);
and U13158 (N_13158,N_12636,N_12419);
nor U13159 (N_13159,N_12616,N_12443);
nand U13160 (N_13160,N_12615,N_12631);
and U13161 (N_13161,N_12403,N_12446);
or U13162 (N_13162,N_12451,N_12602);
and U13163 (N_13163,N_12516,N_12529);
or U13164 (N_13164,N_12594,N_12620);
xnor U13165 (N_13165,N_12593,N_12730);
and U13166 (N_13166,N_12428,N_12463);
xnor U13167 (N_13167,N_12517,N_12549);
and U13168 (N_13168,N_12781,N_12708);
and U13169 (N_13169,N_12704,N_12772);
and U13170 (N_13170,N_12537,N_12607);
xor U13171 (N_13171,N_12732,N_12713);
xnor U13172 (N_13172,N_12410,N_12783);
or U13173 (N_13173,N_12429,N_12637);
nand U13174 (N_13174,N_12455,N_12578);
or U13175 (N_13175,N_12481,N_12592);
xor U13176 (N_13176,N_12766,N_12561);
nand U13177 (N_13177,N_12532,N_12524);
nor U13178 (N_13178,N_12782,N_12688);
and U13179 (N_13179,N_12649,N_12487);
nor U13180 (N_13180,N_12521,N_12555);
or U13181 (N_13181,N_12405,N_12475);
nor U13182 (N_13182,N_12503,N_12755);
nand U13183 (N_13183,N_12505,N_12520);
nor U13184 (N_13184,N_12516,N_12561);
or U13185 (N_13185,N_12630,N_12657);
nor U13186 (N_13186,N_12548,N_12665);
xnor U13187 (N_13187,N_12710,N_12666);
and U13188 (N_13188,N_12733,N_12612);
and U13189 (N_13189,N_12577,N_12737);
nand U13190 (N_13190,N_12704,N_12588);
or U13191 (N_13191,N_12797,N_12483);
nand U13192 (N_13192,N_12422,N_12759);
nor U13193 (N_13193,N_12751,N_12585);
nor U13194 (N_13194,N_12464,N_12496);
or U13195 (N_13195,N_12430,N_12527);
xnor U13196 (N_13196,N_12564,N_12626);
nor U13197 (N_13197,N_12709,N_12442);
xnor U13198 (N_13198,N_12699,N_12404);
or U13199 (N_13199,N_12439,N_12796);
nand U13200 (N_13200,N_12808,N_12828);
xor U13201 (N_13201,N_12922,N_13196);
or U13202 (N_13202,N_13030,N_13151);
or U13203 (N_13203,N_12829,N_12891);
and U13204 (N_13204,N_12976,N_13009);
and U13205 (N_13205,N_12839,N_13168);
and U13206 (N_13206,N_13101,N_13185);
nand U13207 (N_13207,N_13111,N_12858);
xnor U13208 (N_13208,N_13034,N_13124);
and U13209 (N_13209,N_13190,N_13110);
and U13210 (N_13210,N_13028,N_12871);
xor U13211 (N_13211,N_13036,N_13115);
nor U13212 (N_13212,N_13086,N_12855);
nor U13213 (N_13213,N_12833,N_13037);
or U13214 (N_13214,N_13018,N_12819);
and U13215 (N_13215,N_13020,N_13155);
and U13216 (N_13216,N_13065,N_12892);
and U13217 (N_13217,N_12893,N_12914);
nand U13218 (N_13218,N_13123,N_13054);
or U13219 (N_13219,N_12873,N_12803);
and U13220 (N_13220,N_12864,N_13008);
xnor U13221 (N_13221,N_12806,N_13173);
or U13222 (N_13222,N_13141,N_13074);
nand U13223 (N_13223,N_12986,N_13084);
xor U13224 (N_13224,N_12877,N_12822);
nor U13225 (N_13225,N_13023,N_13144);
nand U13226 (N_13226,N_12905,N_13147);
or U13227 (N_13227,N_12980,N_12811);
nand U13228 (N_13228,N_12946,N_13114);
xor U13229 (N_13229,N_12928,N_13029);
nor U13230 (N_13230,N_13135,N_12944);
and U13231 (N_13231,N_12912,N_12959);
xor U13232 (N_13232,N_13098,N_13100);
and U13233 (N_13233,N_13094,N_13143);
or U13234 (N_13234,N_12883,N_13104);
and U13235 (N_13235,N_13152,N_12967);
and U13236 (N_13236,N_12996,N_12801);
xor U13237 (N_13237,N_12863,N_13193);
and U13238 (N_13238,N_12911,N_12963);
nor U13239 (N_13239,N_12993,N_13085);
and U13240 (N_13240,N_12961,N_13072);
and U13241 (N_13241,N_13088,N_12949);
xor U13242 (N_13242,N_12882,N_13099);
and U13243 (N_13243,N_13195,N_13081);
or U13244 (N_13244,N_12902,N_12969);
xnor U13245 (N_13245,N_13004,N_12934);
nor U13246 (N_13246,N_12999,N_13077);
or U13247 (N_13247,N_13162,N_13040);
or U13248 (N_13248,N_12945,N_12805);
or U13249 (N_13249,N_13015,N_13022);
nor U13250 (N_13250,N_12895,N_13116);
and U13251 (N_13251,N_13106,N_12920);
nor U13252 (N_13252,N_12926,N_13049);
and U13253 (N_13253,N_12830,N_13070);
nor U13254 (N_13254,N_13156,N_13131);
or U13255 (N_13255,N_12867,N_13003);
nor U13256 (N_13256,N_13064,N_13026);
or U13257 (N_13257,N_12865,N_12852);
and U13258 (N_13258,N_13073,N_12832);
xnor U13259 (N_13259,N_12915,N_12816);
xor U13260 (N_13260,N_12994,N_12971);
nand U13261 (N_13261,N_13157,N_13118);
and U13262 (N_13262,N_12958,N_13062);
or U13263 (N_13263,N_13090,N_12941);
nand U13264 (N_13264,N_12988,N_13165);
nand U13265 (N_13265,N_13044,N_12856);
and U13266 (N_13266,N_12973,N_13133);
nor U13267 (N_13267,N_12826,N_12862);
and U13268 (N_13268,N_13191,N_12880);
and U13269 (N_13269,N_13045,N_13175);
and U13270 (N_13270,N_13102,N_12807);
and U13271 (N_13271,N_12979,N_13132);
nand U13272 (N_13272,N_13182,N_12935);
nand U13273 (N_13273,N_12917,N_12929);
and U13274 (N_13274,N_13061,N_13186);
xnor U13275 (N_13275,N_13059,N_13035);
nand U13276 (N_13276,N_12872,N_13161);
or U13277 (N_13277,N_13112,N_12870);
and U13278 (N_13278,N_13007,N_13171);
nor U13279 (N_13279,N_12851,N_13056);
or U13280 (N_13280,N_13148,N_12853);
nor U13281 (N_13281,N_13113,N_13105);
or U13282 (N_13282,N_13129,N_12940);
or U13283 (N_13283,N_13067,N_12901);
nand U13284 (N_13284,N_13117,N_12972);
or U13285 (N_13285,N_13192,N_13046);
and U13286 (N_13286,N_12962,N_13032);
nor U13287 (N_13287,N_12874,N_13000);
and U13288 (N_13288,N_13093,N_13174);
nor U13289 (N_13289,N_12974,N_13006);
nand U13290 (N_13290,N_13134,N_13199);
or U13291 (N_13291,N_12981,N_12925);
and U13292 (N_13292,N_13096,N_13089);
or U13293 (N_13293,N_12906,N_13146);
nand U13294 (N_13294,N_13047,N_12978);
and U13295 (N_13295,N_12800,N_13137);
or U13296 (N_13296,N_12834,N_12936);
nor U13297 (N_13297,N_12836,N_13198);
xor U13298 (N_13298,N_12846,N_12884);
and U13299 (N_13299,N_12885,N_12982);
nor U13300 (N_13300,N_13158,N_13033);
xor U13301 (N_13301,N_12859,N_13001);
or U13302 (N_13302,N_13082,N_12931);
xor U13303 (N_13303,N_12907,N_13055);
or U13304 (N_13304,N_12909,N_12923);
nor U13305 (N_13305,N_13140,N_13197);
or U13306 (N_13306,N_13012,N_12990);
nor U13307 (N_13307,N_12814,N_13016);
nand U13308 (N_13308,N_13017,N_12987);
nand U13309 (N_13309,N_13019,N_12841);
and U13310 (N_13310,N_13176,N_13014);
nand U13311 (N_13311,N_13002,N_13095);
nor U13312 (N_13312,N_13080,N_12954);
and U13313 (N_13313,N_12964,N_12998);
nand U13314 (N_13314,N_12838,N_13178);
xor U13315 (N_13315,N_13060,N_13125);
nor U13316 (N_13316,N_12854,N_13087);
xor U13317 (N_13317,N_13139,N_13160);
or U13318 (N_13318,N_12983,N_13024);
xor U13319 (N_13319,N_13068,N_12804);
xnor U13320 (N_13320,N_12835,N_12897);
or U13321 (N_13321,N_12847,N_13188);
nand U13322 (N_13322,N_12843,N_13164);
nor U13323 (N_13323,N_12896,N_12918);
nor U13324 (N_13324,N_12879,N_12878);
xnor U13325 (N_13325,N_12975,N_13092);
nor U13326 (N_13326,N_12930,N_12845);
and U13327 (N_13327,N_13150,N_12957);
nor U13328 (N_13328,N_13128,N_13180);
nand U13329 (N_13329,N_13058,N_13083);
or U13330 (N_13330,N_12844,N_12956);
nor U13331 (N_13331,N_12881,N_12951);
nand U13332 (N_13332,N_12827,N_13179);
xor U13333 (N_13333,N_12989,N_13078);
xor U13334 (N_13334,N_13031,N_13109);
and U13335 (N_13335,N_12985,N_13130);
nor U13336 (N_13336,N_12953,N_12924);
nor U13337 (N_13337,N_13189,N_12916);
nor U13338 (N_13338,N_12888,N_12992);
nand U13339 (N_13339,N_12943,N_12849);
and U13340 (N_13340,N_12960,N_13167);
nor U13341 (N_13341,N_13122,N_13108);
xnor U13342 (N_13342,N_13166,N_13013);
xnor U13343 (N_13343,N_12937,N_13042);
nor U13344 (N_13344,N_13184,N_12886);
and U13345 (N_13345,N_13051,N_12952);
and U13346 (N_13346,N_12821,N_12825);
xnor U13347 (N_13347,N_12942,N_13021);
or U13348 (N_13348,N_13126,N_13107);
xor U13349 (N_13349,N_13005,N_13079);
and U13350 (N_13350,N_12933,N_12875);
and U13351 (N_13351,N_12890,N_13142);
nor U13352 (N_13352,N_12997,N_13053);
or U13353 (N_13353,N_13120,N_12866);
xnor U13354 (N_13354,N_12947,N_12966);
nor U13355 (N_13355,N_13097,N_12889);
nand U13356 (N_13356,N_13181,N_13063);
or U13357 (N_13357,N_12840,N_12908);
nor U13358 (N_13358,N_12948,N_13071);
xor U13359 (N_13359,N_12820,N_13127);
nor U13360 (N_13360,N_13025,N_13170);
xnor U13361 (N_13361,N_12818,N_12837);
nor U13362 (N_13362,N_12876,N_12955);
and U13363 (N_13363,N_13057,N_12887);
xor U13364 (N_13364,N_13010,N_12939);
xor U13365 (N_13365,N_13187,N_13138);
nor U13366 (N_13366,N_13163,N_12848);
xor U13367 (N_13367,N_12913,N_12860);
nor U13368 (N_13368,N_12900,N_12995);
or U13369 (N_13369,N_12938,N_12950);
and U13370 (N_13370,N_12894,N_12868);
nor U13371 (N_13371,N_13103,N_12813);
nand U13372 (N_13372,N_12809,N_12968);
nor U13373 (N_13373,N_12932,N_12927);
or U13374 (N_13374,N_13169,N_12919);
or U13375 (N_13375,N_13076,N_13172);
or U13376 (N_13376,N_13011,N_12898);
or U13377 (N_13377,N_12824,N_13091);
nor U13378 (N_13378,N_13039,N_12965);
and U13379 (N_13379,N_13119,N_12899);
nand U13380 (N_13380,N_12984,N_13075);
or U13381 (N_13381,N_12857,N_13149);
nand U13382 (N_13382,N_12850,N_13069);
nor U13383 (N_13383,N_13183,N_12861);
nand U13384 (N_13384,N_13145,N_13154);
nor U13385 (N_13385,N_12812,N_13041);
and U13386 (N_13386,N_12817,N_12869);
xor U13387 (N_13387,N_12977,N_13136);
and U13388 (N_13388,N_12810,N_12970);
nand U13389 (N_13389,N_12903,N_12842);
nand U13390 (N_13390,N_13043,N_13177);
nand U13391 (N_13391,N_12904,N_12815);
or U13392 (N_13392,N_13153,N_12823);
or U13393 (N_13393,N_13048,N_13050);
nor U13394 (N_13394,N_13159,N_12831);
and U13395 (N_13395,N_13194,N_13027);
xor U13396 (N_13396,N_13052,N_12802);
nand U13397 (N_13397,N_13121,N_13038);
xnor U13398 (N_13398,N_13066,N_12991);
or U13399 (N_13399,N_12910,N_12921);
and U13400 (N_13400,N_13047,N_12808);
and U13401 (N_13401,N_13076,N_12966);
xor U13402 (N_13402,N_13093,N_13041);
nand U13403 (N_13403,N_12868,N_13002);
and U13404 (N_13404,N_13077,N_13054);
or U13405 (N_13405,N_12995,N_13021);
and U13406 (N_13406,N_13184,N_12904);
and U13407 (N_13407,N_13197,N_12894);
or U13408 (N_13408,N_12984,N_13092);
xnor U13409 (N_13409,N_13194,N_13004);
or U13410 (N_13410,N_13031,N_13077);
or U13411 (N_13411,N_13112,N_13021);
and U13412 (N_13412,N_13160,N_12865);
nor U13413 (N_13413,N_12924,N_12800);
xor U13414 (N_13414,N_12914,N_12937);
xor U13415 (N_13415,N_13101,N_12896);
nor U13416 (N_13416,N_12947,N_12996);
nand U13417 (N_13417,N_12932,N_12929);
nand U13418 (N_13418,N_12965,N_12832);
xor U13419 (N_13419,N_13125,N_13127);
nand U13420 (N_13420,N_12894,N_13034);
and U13421 (N_13421,N_12896,N_13090);
or U13422 (N_13422,N_13083,N_13071);
and U13423 (N_13423,N_13006,N_12868);
or U13424 (N_13424,N_13137,N_12837);
nand U13425 (N_13425,N_12936,N_13129);
xor U13426 (N_13426,N_13045,N_12861);
or U13427 (N_13427,N_13074,N_12948);
and U13428 (N_13428,N_12909,N_12938);
and U13429 (N_13429,N_13003,N_13031);
xnor U13430 (N_13430,N_12925,N_13119);
nor U13431 (N_13431,N_13021,N_13067);
or U13432 (N_13432,N_12816,N_13126);
nand U13433 (N_13433,N_13072,N_13147);
or U13434 (N_13434,N_12877,N_13179);
nor U13435 (N_13435,N_12852,N_12812);
nand U13436 (N_13436,N_12838,N_12926);
xor U13437 (N_13437,N_12933,N_12911);
or U13438 (N_13438,N_13060,N_13144);
and U13439 (N_13439,N_13068,N_12802);
nor U13440 (N_13440,N_13064,N_12856);
nand U13441 (N_13441,N_12899,N_13047);
or U13442 (N_13442,N_13181,N_13130);
nand U13443 (N_13443,N_12948,N_12906);
xnor U13444 (N_13444,N_12983,N_12928);
nand U13445 (N_13445,N_13094,N_12941);
nor U13446 (N_13446,N_13142,N_13106);
xnor U13447 (N_13447,N_13166,N_13088);
and U13448 (N_13448,N_12820,N_13043);
xnor U13449 (N_13449,N_13186,N_12887);
or U13450 (N_13450,N_12963,N_13067);
xnor U13451 (N_13451,N_13194,N_13010);
or U13452 (N_13452,N_12833,N_12942);
nor U13453 (N_13453,N_12876,N_12905);
and U13454 (N_13454,N_13079,N_13048);
nor U13455 (N_13455,N_12893,N_12911);
or U13456 (N_13456,N_13073,N_12951);
and U13457 (N_13457,N_13198,N_12953);
and U13458 (N_13458,N_13028,N_13142);
or U13459 (N_13459,N_13183,N_13073);
nor U13460 (N_13460,N_13065,N_12991);
xor U13461 (N_13461,N_13080,N_12861);
and U13462 (N_13462,N_13004,N_12957);
nand U13463 (N_13463,N_12800,N_12859);
nand U13464 (N_13464,N_12995,N_13166);
and U13465 (N_13465,N_13085,N_13128);
nand U13466 (N_13466,N_13094,N_13188);
nand U13467 (N_13467,N_12823,N_12876);
xor U13468 (N_13468,N_12873,N_12840);
xor U13469 (N_13469,N_13164,N_12995);
nor U13470 (N_13470,N_13149,N_12864);
nand U13471 (N_13471,N_12996,N_13000);
nor U13472 (N_13472,N_13002,N_13165);
and U13473 (N_13473,N_12990,N_13007);
or U13474 (N_13474,N_13186,N_12917);
nor U13475 (N_13475,N_12996,N_13155);
nand U13476 (N_13476,N_12811,N_12953);
nor U13477 (N_13477,N_13064,N_13100);
or U13478 (N_13478,N_12812,N_12971);
xor U13479 (N_13479,N_12987,N_13128);
xnor U13480 (N_13480,N_12933,N_12957);
xnor U13481 (N_13481,N_13147,N_13199);
xor U13482 (N_13482,N_13158,N_12998);
nor U13483 (N_13483,N_12932,N_13049);
or U13484 (N_13484,N_13066,N_13037);
and U13485 (N_13485,N_12923,N_12920);
nand U13486 (N_13486,N_13067,N_13162);
xnor U13487 (N_13487,N_13053,N_13108);
or U13488 (N_13488,N_13153,N_12849);
xor U13489 (N_13489,N_13087,N_12992);
nand U13490 (N_13490,N_12878,N_13143);
nand U13491 (N_13491,N_13138,N_13172);
or U13492 (N_13492,N_13033,N_12845);
xor U13493 (N_13493,N_12811,N_13170);
nor U13494 (N_13494,N_12865,N_12866);
and U13495 (N_13495,N_12937,N_13136);
nand U13496 (N_13496,N_12906,N_12874);
nand U13497 (N_13497,N_13114,N_13178);
nor U13498 (N_13498,N_13144,N_13161);
or U13499 (N_13499,N_12864,N_13000);
or U13500 (N_13500,N_12807,N_13118);
or U13501 (N_13501,N_13183,N_13015);
or U13502 (N_13502,N_13132,N_12971);
nor U13503 (N_13503,N_12824,N_13150);
nor U13504 (N_13504,N_12934,N_13183);
or U13505 (N_13505,N_13141,N_13057);
xnor U13506 (N_13506,N_13077,N_13005);
and U13507 (N_13507,N_12850,N_13116);
nor U13508 (N_13508,N_13021,N_12825);
nor U13509 (N_13509,N_13028,N_13132);
nor U13510 (N_13510,N_13197,N_12940);
nor U13511 (N_13511,N_12830,N_12989);
xor U13512 (N_13512,N_12857,N_12843);
or U13513 (N_13513,N_13150,N_13078);
nand U13514 (N_13514,N_12875,N_12910);
or U13515 (N_13515,N_12879,N_13078);
nor U13516 (N_13516,N_13167,N_12899);
and U13517 (N_13517,N_13167,N_12928);
and U13518 (N_13518,N_12836,N_12970);
or U13519 (N_13519,N_12911,N_13093);
nand U13520 (N_13520,N_13165,N_13033);
or U13521 (N_13521,N_12853,N_13197);
nor U13522 (N_13522,N_13146,N_12941);
and U13523 (N_13523,N_12857,N_13094);
nor U13524 (N_13524,N_13061,N_13016);
nor U13525 (N_13525,N_13109,N_13125);
xor U13526 (N_13526,N_13050,N_13091);
nand U13527 (N_13527,N_13146,N_13023);
or U13528 (N_13528,N_13110,N_12890);
nand U13529 (N_13529,N_12950,N_13106);
and U13530 (N_13530,N_12862,N_13197);
xor U13531 (N_13531,N_13065,N_13105);
and U13532 (N_13532,N_13180,N_12924);
xnor U13533 (N_13533,N_12906,N_12956);
nand U13534 (N_13534,N_13039,N_13178);
or U13535 (N_13535,N_13110,N_12835);
nor U13536 (N_13536,N_13031,N_13100);
nand U13537 (N_13537,N_13117,N_13155);
xor U13538 (N_13538,N_12864,N_12909);
or U13539 (N_13539,N_12951,N_13164);
xnor U13540 (N_13540,N_13105,N_12937);
or U13541 (N_13541,N_13189,N_12928);
and U13542 (N_13542,N_13110,N_13106);
nand U13543 (N_13543,N_12877,N_12801);
nor U13544 (N_13544,N_12987,N_12908);
nor U13545 (N_13545,N_13129,N_12974);
nand U13546 (N_13546,N_12977,N_12841);
or U13547 (N_13547,N_13080,N_13062);
xnor U13548 (N_13548,N_13086,N_12816);
xnor U13549 (N_13549,N_13026,N_13009);
nand U13550 (N_13550,N_13155,N_12882);
nor U13551 (N_13551,N_13090,N_13108);
and U13552 (N_13552,N_12843,N_13037);
xor U13553 (N_13553,N_13071,N_12855);
and U13554 (N_13554,N_12946,N_12980);
xor U13555 (N_13555,N_12903,N_12960);
and U13556 (N_13556,N_13181,N_13050);
or U13557 (N_13557,N_12913,N_12824);
xnor U13558 (N_13558,N_12853,N_12962);
xor U13559 (N_13559,N_12942,N_12991);
nand U13560 (N_13560,N_12825,N_12859);
nand U13561 (N_13561,N_13039,N_13084);
and U13562 (N_13562,N_12833,N_13119);
nand U13563 (N_13563,N_12910,N_13103);
or U13564 (N_13564,N_13130,N_12923);
or U13565 (N_13565,N_13087,N_12929);
nand U13566 (N_13566,N_12994,N_12832);
nor U13567 (N_13567,N_13079,N_13027);
nand U13568 (N_13568,N_13182,N_12813);
xor U13569 (N_13569,N_12845,N_12991);
or U13570 (N_13570,N_13010,N_12847);
nand U13571 (N_13571,N_12892,N_13135);
and U13572 (N_13572,N_12939,N_12808);
xnor U13573 (N_13573,N_12854,N_12855);
and U13574 (N_13574,N_13031,N_12988);
xor U13575 (N_13575,N_13053,N_12893);
nand U13576 (N_13576,N_12953,N_13015);
nand U13577 (N_13577,N_12963,N_13114);
nand U13578 (N_13578,N_13079,N_13063);
or U13579 (N_13579,N_12851,N_12802);
and U13580 (N_13580,N_12945,N_13007);
nand U13581 (N_13581,N_12854,N_12833);
and U13582 (N_13582,N_12956,N_13155);
nor U13583 (N_13583,N_12918,N_13117);
and U13584 (N_13584,N_12941,N_12817);
and U13585 (N_13585,N_13155,N_13194);
and U13586 (N_13586,N_13116,N_12830);
xor U13587 (N_13587,N_13170,N_13014);
nand U13588 (N_13588,N_13085,N_13144);
and U13589 (N_13589,N_12890,N_13043);
xnor U13590 (N_13590,N_12903,N_12873);
xor U13591 (N_13591,N_12829,N_13091);
nor U13592 (N_13592,N_12928,N_12817);
nor U13593 (N_13593,N_12863,N_13153);
and U13594 (N_13594,N_13059,N_12973);
and U13595 (N_13595,N_13070,N_13057);
nor U13596 (N_13596,N_12958,N_13044);
and U13597 (N_13597,N_12880,N_12996);
nand U13598 (N_13598,N_13034,N_12929);
xnor U13599 (N_13599,N_13141,N_12928);
nand U13600 (N_13600,N_13359,N_13328);
nor U13601 (N_13601,N_13383,N_13353);
nor U13602 (N_13602,N_13317,N_13387);
xor U13603 (N_13603,N_13203,N_13391);
xnor U13604 (N_13604,N_13447,N_13311);
xor U13605 (N_13605,N_13453,N_13486);
or U13606 (N_13606,N_13440,N_13270);
and U13607 (N_13607,N_13514,N_13573);
or U13608 (N_13608,N_13424,N_13577);
or U13609 (N_13609,N_13288,N_13558);
nor U13610 (N_13610,N_13448,N_13475);
xor U13611 (N_13611,N_13268,N_13471);
and U13612 (N_13612,N_13588,N_13252);
or U13613 (N_13613,N_13239,N_13429);
xnor U13614 (N_13614,N_13456,N_13451);
or U13615 (N_13615,N_13389,N_13274);
and U13616 (N_13616,N_13444,N_13499);
nand U13617 (N_13617,N_13281,N_13264);
nand U13618 (N_13618,N_13404,N_13285);
xor U13619 (N_13619,N_13323,N_13445);
nor U13620 (N_13620,N_13555,N_13282);
and U13621 (N_13621,N_13520,N_13345);
nor U13622 (N_13622,N_13375,N_13489);
xnor U13623 (N_13623,N_13412,N_13421);
and U13624 (N_13624,N_13557,N_13218);
xnor U13625 (N_13625,N_13427,N_13291);
or U13626 (N_13626,N_13518,N_13519);
nand U13627 (N_13627,N_13493,N_13432);
and U13628 (N_13628,N_13305,N_13470);
nor U13629 (N_13629,N_13221,N_13420);
xor U13630 (N_13630,N_13565,N_13572);
or U13631 (N_13631,N_13370,N_13251);
or U13632 (N_13632,N_13243,N_13304);
nand U13633 (N_13633,N_13483,N_13235);
or U13634 (N_13634,N_13594,N_13388);
and U13635 (N_13635,N_13337,N_13494);
xor U13636 (N_13636,N_13552,N_13267);
nor U13637 (N_13637,N_13228,N_13276);
xnor U13638 (N_13638,N_13393,N_13501);
nor U13639 (N_13639,N_13208,N_13576);
or U13640 (N_13640,N_13356,N_13454);
xnor U13641 (N_13641,N_13418,N_13597);
or U13642 (N_13642,N_13488,N_13508);
or U13643 (N_13643,N_13405,N_13461);
xnor U13644 (N_13644,N_13215,N_13322);
xnor U13645 (N_13645,N_13423,N_13502);
and U13646 (N_13646,N_13299,N_13306);
nor U13647 (N_13647,N_13587,N_13240);
xor U13648 (N_13648,N_13210,N_13455);
or U13649 (N_13649,N_13296,N_13211);
xor U13650 (N_13650,N_13439,N_13592);
or U13651 (N_13651,N_13583,N_13544);
or U13652 (N_13652,N_13517,N_13318);
nand U13653 (N_13653,N_13372,N_13524);
or U13654 (N_13654,N_13376,N_13283);
or U13655 (N_13655,N_13233,N_13244);
nand U13656 (N_13656,N_13309,N_13556);
or U13657 (N_13657,N_13255,N_13277);
nor U13658 (N_13658,N_13400,N_13542);
or U13659 (N_13659,N_13348,N_13428);
xnor U13660 (N_13660,N_13509,N_13338);
xor U13661 (N_13661,N_13408,N_13415);
xor U13662 (N_13662,N_13272,N_13549);
or U13663 (N_13663,N_13350,N_13416);
nand U13664 (N_13664,N_13342,N_13574);
nand U13665 (N_13665,N_13580,N_13554);
and U13666 (N_13666,N_13566,N_13452);
and U13667 (N_13667,N_13516,N_13510);
xor U13668 (N_13668,N_13589,N_13246);
nand U13669 (N_13669,N_13327,N_13563);
or U13670 (N_13670,N_13579,N_13598);
or U13671 (N_13671,N_13326,N_13314);
and U13672 (N_13672,N_13414,N_13398);
nand U13673 (N_13673,N_13377,N_13262);
and U13674 (N_13674,N_13530,N_13473);
nor U13675 (N_13675,N_13586,N_13321);
and U13676 (N_13676,N_13310,N_13234);
nor U13677 (N_13677,N_13485,N_13212);
xnor U13678 (N_13678,N_13362,N_13507);
nor U13679 (N_13679,N_13223,N_13320);
nand U13680 (N_13680,N_13490,N_13339);
nand U13681 (N_13681,N_13535,N_13543);
xnor U13682 (N_13682,N_13443,N_13365);
nand U13683 (N_13683,N_13357,N_13332);
nor U13684 (N_13684,N_13459,N_13496);
and U13685 (N_13685,N_13373,N_13546);
xnor U13686 (N_13686,N_13504,N_13380);
nand U13687 (N_13687,N_13249,N_13464);
xor U13688 (N_13688,N_13225,N_13278);
and U13689 (N_13689,N_13351,N_13265);
xnor U13690 (N_13690,N_13495,N_13528);
or U13691 (N_13691,N_13515,N_13430);
nor U13692 (N_13692,N_13275,N_13216);
and U13693 (N_13693,N_13532,N_13472);
or U13694 (N_13694,N_13425,N_13536);
xor U13695 (N_13695,N_13220,N_13341);
nand U13696 (N_13696,N_13319,N_13395);
xnor U13697 (N_13697,N_13273,N_13287);
or U13698 (N_13698,N_13284,N_13333);
and U13699 (N_13699,N_13349,N_13522);
or U13700 (N_13700,N_13300,N_13410);
xor U13701 (N_13701,N_13325,N_13575);
nand U13702 (N_13702,N_13437,N_13254);
nor U13703 (N_13703,N_13492,N_13258);
xnor U13704 (N_13704,N_13385,N_13458);
and U13705 (N_13705,N_13512,N_13417);
nand U13706 (N_13706,N_13201,N_13571);
and U13707 (N_13707,N_13253,N_13467);
or U13708 (N_13708,N_13289,N_13540);
xnor U13709 (N_13709,N_13596,N_13595);
nor U13710 (N_13710,N_13374,N_13537);
nor U13711 (N_13711,N_13476,N_13331);
xor U13712 (N_13712,N_13403,N_13263);
and U13713 (N_13713,N_13336,N_13409);
or U13714 (N_13714,N_13584,N_13346);
xnor U13715 (N_13715,N_13379,N_13550);
and U13716 (N_13716,N_13545,N_13286);
nand U13717 (N_13717,N_13560,N_13355);
and U13718 (N_13718,N_13438,N_13334);
nor U13719 (N_13719,N_13358,N_13590);
nand U13720 (N_13720,N_13581,N_13266);
or U13721 (N_13721,N_13324,N_13271);
nand U13722 (N_13722,N_13247,N_13237);
and U13723 (N_13723,N_13371,N_13585);
and U13724 (N_13724,N_13396,N_13497);
or U13725 (N_13725,N_13312,N_13491);
xor U13726 (N_13726,N_13591,N_13369);
nand U13727 (N_13727,N_13570,N_13361);
xnor U13728 (N_13728,N_13307,N_13433);
xnor U13729 (N_13729,N_13397,N_13513);
and U13730 (N_13730,N_13477,N_13261);
and U13731 (N_13731,N_13578,N_13363);
or U13732 (N_13732,N_13347,N_13561);
or U13733 (N_13733,N_13269,N_13564);
xnor U13734 (N_13734,N_13204,N_13242);
xnor U13735 (N_13735,N_13303,N_13386);
nor U13736 (N_13736,N_13526,N_13413);
xnor U13737 (N_13737,N_13207,N_13360);
xor U13738 (N_13738,N_13406,N_13527);
or U13739 (N_13739,N_13213,N_13506);
nor U13740 (N_13740,N_13538,N_13460);
or U13741 (N_13741,N_13469,N_13498);
nor U13742 (N_13742,N_13279,N_13446);
nand U13743 (N_13743,N_13313,N_13569);
and U13744 (N_13744,N_13250,N_13381);
nand U13745 (N_13745,N_13343,N_13241);
or U13746 (N_13746,N_13434,N_13295);
xnor U13747 (N_13747,N_13230,N_13511);
nand U13748 (N_13748,N_13206,N_13441);
and U13749 (N_13749,N_13294,N_13466);
xnor U13750 (N_13750,N_13582,N_13227);
and U13751 (N_13751,N_13531,N_13481);
nor U13752 (N_13752,N_13390,N_13482);
xnor U13753 (N_13753,N_13248,N_13500);
nand U13754 (N_13754,N_13449,N_13529);
xor U13755 (N_13755,N_13200,N_13226);
and U13756 (N_13756,N_13468,N_13301);
xnor U13757 (N_13757,N_13205,N_13352);
or U13758 (N_13758,N_13367,N_13298);
xnor U13759 (N_13759,N_13539,N_13484);
or U13760 (N_13760,N_13308,N_13260);
or U13761 (N_13761,N_13259,N_13257);
nand U13762 (N_13762,N_13521,N_13431);
nor U13763 (N_13763,N_13422,N_13533);
nand U13764 (N_13764,N_13354,N_13463);
or U13765 (N_13765,N_13302,N_13222);
nor U13766 (N_13766,N_13478,N_13392);
nand U13767 (N_13767,N_13551,N_13547);
nand U13768 (N_13768,N_13442,N_13401);
nor U13769 (N_13769,N_13209,N_13568);
xnor U13770 (N_13770,N_13407,N_13474);
xnor U13771 (N_13771,N_13384,N_13293);
nor U13772 (N_13772,N_13330,N_13525);
and U13773 (N_13773,N_13232,N_13394);
xor U13774 (N_13774,N_13202,N_13435);
xnor U13775 (N_13775,N_13548,N_13436);
nor U13776 (N_13776,N_13224,N_13559);
and U13777 (N_13777,N_13229,N_13236);
xor U13778 (N_13778,N_13562,N_13419);
nor U13779 (N_13779,N_13402,N_13426);
and U13780 (N_13780,N_13366,N_13479);
and U13781 (N_13781,N_13567,N_13256);
xnor U13782 (N_13782,N_13523,N_13329);
or U13783 (N_13783,N_13599,N_13219);
nor U13784 (N_13784,N_13335,N_13534);
nor U13785 (N_13785,N_13231,N_13214);
nor U13786 (N_13786,N_13292,N_13450);
or U13787 (N_13787,N_13465,N_13480);
xor U13788 (N_13788,N_13378,N_13364);
or U13789 (N_13789,N_13487,N_13503);
nand U13790 (N_13790,N_13315,N_13541);
xor U13791 (N_13791,N_13368,N_13411);
or U13792 (N_13792,N_13340,N_13316);
or U13793 (N_13793,N_13593,N_13553);
and U13794 (N_13794,N_13344,N_13297);
nand U13795 (N_13795,N_13280,N_13462);
and U13796 (N_13796,N_13457,N_13290);
nor U13797 (N_13797,N_13382,N_13505);
nor U13798 (N_13798,N_13217,N_13399);
or U13799 (N_13799,N_13245,N_13238);
xor U13800 (N_13800,N_13462,N_13256);
nor U13801 (N_13801,N_13417,N_13354);
nor U13802 (N_13802,N_13210,N_13303);
nor U13803 (N_13803,N_13303,N_13361);
nand U13804 (N_13804,N_13397,N_13452);
or U13805 (N_13805,N_13355,N_13281);
nor U13806 (N_13806,N_13334,N_13300);
and U13807 (N_13807,N_13225,N_13471);
xor U13808 (N_13808,N_13242,N_13462);
and U13809 (N_13809,N_13582,N_13312);
and U13810 (N_13810,N_13513,N_13398);
and U13811 (N_13811,N_13329,N_13404);
and U13812 (N_13812,N_13226,N_13350);
or U13813 (N_13813,N_13441,N_13326);
nand U13814 (N_13814,N_13430,N_13502);
nand U13815 (N_13815,N_13576,N_13308);
or U13816 (N_13816,N_13571,N_13358);
or U13817 (N_13817,N_13397,N_13548);
or U13818 (N_13818,N_13366,N_13295);
nor U13819 (N_13819,N_13211,N_13308);
xor U13820 (N_13820,N_13320,N_13555);
xnor U13821 (N_13821,N_13224,N_13273);
nand U13822 (N_13822,N_13379,N_13454);
or U13823 (N_13823,N_13432,N_13208);
or U13824 (N_13824,N_13379,N_13461);
and U13825 (N_13825,N_13423,N_13398);
or U13826 (N_13826,N_13382,N_13229);
nor U13827 (N_13827,N_13517,N_13476);
nand U13828 (N_13828,N_13409,N_13398);
nor U13829 (N_13829,N_13448,N_13420);
xnor U13830 (N_13830,N_13313,N_13577);
or U13831 (N_13831,N_13539,N_13594);
and U13832 (N_13832,N_13220,N_13431);
or U13833 (N_13833,N_13342,N_13310);
and U13834 (N_13834,N_13394,N_13430);
nor U13835 (N_13835,N_13252,N_13448);
xnor U13836 (N_13836,N_13498,N_13518);
xnor U13837 (N_13837,N_13546,N_13380);
nor U13838 (N_13838,N_13253,N_13314);
xnor U13839 (N_13839,N_13530,N_13293);
nor U13840 (N_13840,N_13590,N_13332);
nor U13841 (N_13841,N_13248,N_13230);
nor U13842 (N_13842,N_13593,N_13242);
nand U13843 (N_13843,N_13338,N_13273);
xor U13844 (N_13844,N_13339,N_13369);
xor U13845 (N_13845,N_13442,N_13311);
nor U13846 (N_13846,N_13373,N_13356);
xor U13847 (N_13847,N_13565,N_13519);
nor U13848 (N_13848,N_13484,N_13406);
and U13849 (N_13849,N_13218,N_13595);
xnor U13850 (N_13850,N_13454,N_13377);
nor U13851 (N_13851,N_13285,N_13282);
xor U13852 (N_13852,N_13546,N_13573);
nand U13853 (N_13853,N_13525,N_13523);
nand U13854 (N_13854,N_13290,N_13211);
xnor U13855 (N_13855,N_13237,N_13297);
xnor U13856 (N_13856,N_13310,N_13293);
and U13857 (N_13857,N_13445,N_13318);
nand U13858 (N_13858,N_13462,N_13512);
or U13859 (N_13859,N_13339,N_13416);
xor U13860 (N_13860,N_13567,N_13437);
xor U13861 (N_13861,N_13369,N_13435);
nor U13862 (N_13862,N_13406,N_13220);
xor U13863 (N_13863,N_13333,N_13355);
nand U13864 (N_13864,N_13318,N_13556);
or U13865 (N_13865,N_13495,N_13321);
and U13866 (N_13866,N_13323,N_13349);
and U13867 (N_13867,N_13479,N_13372);
nand U13868 (N_13868,N_13450,N_13269);
xnor U13869 (N_13869,N_13201,N_13287);
xnor U13870 (N_13870,N_13497,N_13243);
xor U13871 (N_13871,N_13471,N_13503);
and U13872 (N_13872,N_13367,N_13577);
xor U13873 (N_13873,N_13209,N_13232);
and U13874 (N_13874,N_13236,N_13572);
or U13875 (N_13875,N_13257,N_13387);
or U13876 (N_13876,N_13339,N_13308);
and U13877 (N_13877,N_13559,N_13592);
xor U13878 (N_13878,N_13354,N_13561);
xor U13879 (N_13879,N_13577,N_13231);
xnor U13880 (N_13880,N_13524,N_13386);
and U13881 (N_13881,N_13314,N_13274);
xnor U13882 (N_13882,N_13342,N_13546);
nand U13883 (N_13883,N_13277,N_13386);
nand U13884 (N_13884,N_13437,N_13239);
and U13885 (N_13885,N_13528,N_13280);
nand U13886 (N_13886,N_13436,N_13483);
xnor U13887 (N_13887,N_13588,N_13279);
nand U13888 (N_13888,N_13503,N_13349);
nor U13889 (N_13889,N_13369,N_13564);
nor U13890 (N_13890,N_13553,N_13519);
xor U13891 (N_13891,N_13370,N_13298);
xnor U13892 (N_13892,N_13449,N_13499);
and U13893 (N_13893,N_13216,N_13352);
nor U13894 (N_13894,N_13468,N_13230);
nand U13895 (N_13895,N_13555,N_13436);
nand U13896 (N_13896,N_13326,N_13264);
and U13897 (N_13897,N_13286,N_13431);
nand U13898 (N_13898,N_13403,N_13311);
or U13899 (N_13899,N_13394,N_13260);
nand U13900 (N_13900,N_13407,N_13447);
and U13901 (N_13901,N_13326,N_13344);
xor U13902 (N_13902,N_13230,N_13337);
xor U13903 (N_13903,N_13397,N_13492);
xnor U13904 (N_13904,N_13517,N_13538);
xor U13905 (N_13905,N_13325,N_13541);
xnor U13906 (N_13906,N_13491,N_13419);
nand U13907 (N_13907,N_13368,N_13380);
and U13908 (N_13908,N_13425,N_13391);
and U13909 (N_13909,N_13246,N_13349);
nand U13910 (N_13910,N_13598,N_13381);
xnor U13911 (N_13911,N_13504,N_13524);
or U13912 (N_13912,N_13324,N_13596);
or U13913 (N_13913,N_13579,N_13518);
or U13914 (N_13914,N_13325,N_13251);
and U13915 (N_13915,N_13569,N_13429);
nand U13916 (N_13916,N_13413,N_13292);
nor U13917 (N_13917,N_13439,N_13550);
xnor U13918 (N_13918,N_13560,N_13201);
nor U13919 (N_13919,N_13405,N_13442);
nor U13920 (N_13920,N_13266,N_13565);
nor U13921 (N_13921,N_13500,N_13586);
xor U13922 (N_13922,N_13342,N_13594);
and U13923 (N_13923,N_13485,N_13402);
and U13924 (N_13924,N_13493,N_13505);
xor U13925 (N_13925,N_13589,N_13233);
and U13926 (N_13926,N_13223,N_13222);
or U13927 (N_13927,N_13427,N_13287);
nor U13928 (N_13928,N_13587,N_13452);
nor U13929 (N_13929,N_13274,N_13360);
and U13930 (N_13930,N_13572,N_13233);
or U13931 (N_13931,N_13395,N_13552);
xor U13932 (N_13932,N_13402,N_13451);
and U13933 (N_13933,N_13455,N_13312);
nand U13934 (N_13934,N_13557,N_13222);
xor U13935 (N_13935,N_13209,N_13390);
nand U13936 (N_13936,N_13541,N_13204);
nor U13937 (N_13937,N_13379,N_13578);
and U13938 (N_13938,N_13402,N_13237);
or U13939 (N_13939,N_13533,N_13479);
or U13940 (N_13940,N_13528,N_13589);
and U13941 (N_13941,N_13469,N_13205);
nor U13942 (N_13942,N_13289,N_13260);
nor U13943 (N_13943,N_13567,N_13585);
or U13944 (N_13944,N_13485,N_13570);
xnor U13945 (N_13945,N_13252,N_13254);
xor U13946 (N_13946,N_13389,N_13556);
or U13947 (N_13947,N_13332,N_13523);
xnor U13948 (N_13948,N_13571,N_13217);
or U13949 (N_13949,N_13216,N_13365);
xnor U13950 (N_13950,N_13530,N_13378);
xnor U13951 (N_13951,N_13392,N_13528);
nand U13952 (N_13952,N_13489,N_13463);
xor U13953 (N_13953,N_13421,N_13547);
or U13954 (N_13954,N_13570,N_13459);
nor U13955 (N_13955,N_13343,N_13344);
nor U13956 (N_13956,N_13245,N_13350);
and U13957 (N_13957,N_13413,N_13232);
xnor U13958 (N_13958,N_13281,N_13575);
nand U13959 (N_13959,N_13212,N_13384);
and U13960 (N_13960,N_13422,N_13342);
and U13961 (N_13961,N_13261,N_13324);
or U13962 (N_13962,N_13414,N_13520);
xor U13963 (N_13963,N_13339,N_13448);
and U13964 (N_13964,N_13278,N_13555);
nor U13965 (N_13965,N_13274,N_13552);
xnor U13966 (N_13966,N_13215,N_13260);
and U13967 (N_13967,N_13395,N_13385);
nor U13968 (N_13968,N_13590,N_13270);
nor U13969 (N_13969,N_13305,N_13204);
xor U13970 (N_13970,N_13487,N_13561);
xor U13971 (N_13971,N_13344,N_13267);
xnor U13972 (N_13972,N_13384,N_13298);
nand U13973 (N_13973,N_13458,N_13513);
nor U13974 (N_13974,N_13325,N_13271);
and U13975 (N_13975,N_13259,N_13299);
and U13976 (N_13976,N_13213,N_13396);
and U13977 (N_13977,N_13363,N_13330);
nor U13978 (N_13978,N_13357,N_13262);
xnor U13979 (N_13979,N_13211,N_13204);
and U13980 (N_13980,N_13566,N_13310);
nor U13981 (N_13981,N_13351,N_13295);
or U13982 (N_13982,N_13557,N_13473);
nor U13983 (N_13983,N_13317,N_13490);
or U13984 (N_13984,N_13222,N_13208);
and U13985 (N_13985,N_13362,N_13487);
xnor U13986 (N_13986,N_13420,N_13411);
xnor U13987 (N_13987,N_13535,N_13279);
and U13988 (N_13988,N_13544,N_13419);
nor U13989 (N_13989,N_13574,N_13226);
nor U13990 (N_13990,N_13375,N_13490);
nor U13991 (N_13991,N_13566,N_13565);
nand U13992 (N_13992,N_13427,N_13515);
nand U13993 (N_13993,N_13261,N_13400);
nor U13994 (N_13994,N_13561,N_13205);
xnor U13995 (N_13995,N_13524,N_13309);
or U13996 (N_13996,N_13583,N_13257);
nor U13997 (N_13997,N_13329,N_13233);
nand U13998 (N_13998,N_13352,N_13475);
and U13999 (N_13999,N_13338,N_13220);
or U14000 (N_14000,N_13903,N_13688);
and U14001 (N_14001,N_13873,N_13817);
xnor U14002 (N_14002,N_13835,N_13967);
and U14003 (N_14003,N_13821,N_13709);
nor U14004 (N_14004,N_13915,N_13824);
xnor U14005 (N_14005,N_13942,N_13671);
and U14006 (N_14006,N_13697,N_13608);
and U14007 (N_14007,N_13693,N_13989);
nor U14008 (N_14008,N_13675,N_13762);
nand U14009 (N_14009,N_13600,N_13870);
nor U14010 (N_14010,N_13845,N_13815);
nand U14011 (N_14011,N_13722,N_13751);
xor U14012 (N_14012,N_13711,N_13929);
and U14013 (N_14013,N_13670,N_13909);
nand U14014 (N_14014,N_13650,N_13914);
and U14015 (N_14015,N_13640,N_13853);
or U14016 (N_14016,N_13872,N_13962);
and U14017 (N_14017,N_13740,N_13612);
or U14018 (N_14018,N_13772,N_13826);
xor U14019 (N_14019,N_13738,N_13776);
and U14020 (N_14020,N_13764,N_13834);
and U14021 (N_14021,N_13859,N_13829);
nand U14022 (N_14022,N_13951,N_13869);
and U14023 (N_14023,N_13712,N_13863);
or U14024 (N_14024,N_13921,N_13832);
xnor U14025 (N_14025,N_13808,N_13771);
and U14026 (N_14026,N_13926,N_13953);
nor U14027 (N_14027,N_13797,N_13961);
and U14028 (N_14028,N_13878,N_13755);
nor U14029 (N_14029,N_13790,N_13628);
nand U14030 (N_14030,N_13792,N_13736);
nand U14031 (N_14031,N_13976,N_13723);
nand U14032 (N_14032,N_13681,N_13954);
xnor U14033 (N_14033,N_13981,N_13999);
nor U14034 (N_14034,N_13615,N_13818);
nand U14035 (N_14035,N_13918,N_13663);
and U14036 (N_14036,N_13984,N_13925);
xnor U14037 (N_14037,N_13777,N_13644);
or U14038 (N_14038,N_13623,N_13719);
or U14039 (N_14039,N_13964,N_13896);
nor U14040 (N_14040,N_13922,N_13780);
nor U14041 (N_14041,N_13888,N_13674);
or U14042 (N_14042,N_13843,N_13897);
xnor U14043 (N_14043,N_13858,N_13744);
nor U14044 (N_14044,N_13747,N_13759);
nor U14045 (N_14045,N_13960,N_13767);
nor U14046 (N_14046,N_13812,N_13911);
nand U14047 (N_14047,N_13912,N_13654);
nor U14048 (N_14048,N_13643,N_13716);
and U14049 (N_14049,N_13754,N_13703);
nand U14050 (N_14050,N_13705,N_13787);
and U14051 (N_14051,N_13758,N_13837);
nand U14052 (N_14052,N_13864,N_13848);
nor U14053 (N_14053,N_13955,N_13930);
nand U14054 (N_14054,N_13645,N_13778);
and U14055 (N_14055,N_13865,N_13831);
nand U14056 (N_14056,N_13769,N_13957);
and U14057 (N_14057,N_13680,N_13616);
nand U14058 (N_14058,N_13852,N_13701);
nand U14059 (N_14059,N_13673,N_13841);
xnor U14060 (N_14060,N_13983,N_13657);
xor U14061 (N_14061,N_13820,N_13696);
or U14062 (N_14062,N_13613,N_13624);
xor U14063 (N_14063,N_13795,N_13672);
or U14064 (N_14064,N_13940,N_13810);
or U14065 (N_14065,N_13803,N_13879);
nor U14066 (N_14066,N_13713,N_13653);
or U14067 (N_14067,N_13816,N_13760);
or U14068 (N_14068,N_13847,N_13900);
or U14069 (N_14069,N_13796,N_13782);
or U14070 (N_14070,N_13646,N_13811);
and U14071 (N_14071,N_13799,N_13775);
nand U14072 (N_14072,N_13710,N_13655);
xor U14073 (N_14073,N_13849,N_13916);
nand U14074 (N_14074,N_13636,N_13609);
and U14075 (N_14075,N_13979,N_13721);
nand U14076 (N_14076,N_13698,N_13602);
xor U14077 (N_14077,N_13935,N_13883);
and U14078 (N_14078,N_13938,N_13689);
or U14079 (N_14079,N_13913,N_13631);
nand U14080 (N_14080,N_13601,N_13625);
and U14081 (N_14081,N_13948,N_13881);
nor U14082 (N_14082,N_13844,N_13784);
or U14083 (N_14083,N_13980,N_13949);
nor U14084 (N_14084,N_13635,N_13684);
xnor U14085 (N_14085,N_13885,N_13724);
nor U14086 (N_14086,N_13904,N_13910);
or U14087 (N_14087,N_13828,N_13850);
or U14088 (N_14088,N_13669,N_13927);
xnor U14089 (N_14089,N_13814,N_13833);
xor U14090 (N_14090,N_13750,N_13895);
nor U14091 (N_14091,N_13996,N_13614);
nor U14092 (N_14092,N_13765,N_13757);
nor U14093 (N_14093,N_13891,N_13920);
and U14094 (N_14094,N_13768,N_13699);
nor U14095 (N_14095,N_13708,N_13839);
or U14096 (N_14096,N_13685,N_13735);
and U14097 (N_14097,N_13781,N_13854);
nand U14098 (N_14098,N_13667,N_13785);
nor U14099 (N_14099,N_13978,N_13620);
nor U14100 (N_14100,N_13627,N_13855);
or U14101 (N_14101,N_13741,N_13813);
or U14102 (N_14102,N_13846,N_13791);
and U14103 (N_14103,N_13678,N_13793);
or U14104 (N_14104,N_13731,N_13739);
xnor U14105 (N_14105,N_13648,N_13786);
nor U14106 (N_14106,N_13605,N_13867);
nand U14107 (N_14107,N_13958,N_13634);
and U14108 (N_14108,N_13941,N_13714);
nor U14109 (N_14109,N_13973,N_13823);
nor U14110 (N_14110,N_13742,N_13804);
nand U14111 (N_14111,N_13622,N_13905);
and U14112 (N_14112,N_13945,N_13836);
nand U14113 (N_14113,N_13856,N_13977);
nor U14114 (N_14114,N_13652,N_13923);
nor U14115 (N_14115,N_13748,N_13611);
or U14116 (N_14116,N_13687,N_13734);
xnor U14117 (N_14117,N_13950,N_13761);
nor U14118 (N_14118,N_13908,N_13805);
or U14119 (N_14119,N_13756,N_13665);
or U14120 (N_14120,N_13691,N_13919);
and U14121 (N_14121,N_13963,N_13906);
xnor U14122 (N_14122,N_13875,N_13871);
nor U14123 (N_14123,N_13706,N_13683);
nor U14124 (N_14124,N_13662,N_13763);
or U14125 (N_14125,N_13774,N_13874);
and U14126 (N_14126,N_13728,N_13842);
or U14127 (N_14127,N_13966,N_13933);
nor U14128 (N_14128,N_13860,N_13647);
xor U14129 (N_14129,N_13946,N_13857);
nand U14130 (N_14130,N_13800,N_13807);
or U14131 (N_14131,N_13985,N_13656);
and U14132 (N_14132,N_13783,N_13727);
and U14133 (N_14133,N_13991,N_13773);
and U14134 (N_14134,N_13986,N_13629);
xor U14135 (N_14135,N_13664,N_13630);
nor U14136 (N_14136,N_13880,N_13715);
nand U14137 (N_14137,N_13660,N_13690);
xnor U14138 (N_14138,N_13752,N_13937);
nand U14139 (N_14139,N_13982,N_13718);
nor U14140 (N_14140,N_13788,N_13725);
xnor U14141 (N_14141,N_13998,N_13745);
nand U14142 (N_14142,N_13753,N_13947);
or U14143 (N_14143,N_13621,N_13868);
nand U14144 (N_14144,N_13642,N_13668);
or U14145 (N_14145,N_13801,N_13994);
nor U14146 (N_14146,N_13840,N_13892);
or U14147 (N_14147,N_13694,N_13997);
and U14148 (N_14148,N_13968,N_13898);
or U14149 (N_14149,N_13658,N_13877);
xnor U14150 (N_14150,N_13626,N_13944);
nand U14151 (N_14151,N_13819,N_13749);
nor U14152 (N_14152,N_13825,N_13902);
nand U14153 (N_14153,N_13939,N_13641);
and U14154 (N_14154,N_13651,N_13866);
nand U14155 (N_14155,N_13993,N_13726);
or U14156 (N_14156,N_13928,N_13884);
or U14157 (N_14157,N_13838,N_13969);
or U14158 (N_14158,N_13737,N_13932);
nor U14159 (N_14159,N_13861,N_13889);
xor U14160 (N_14160,N_13679,N_13907);
or U14161 (N_14161,N_13633,N_13618);
or U14162 (N_14162,N_13607,N_13830);
and U14163 (N_14163,N_13702,N_13606);
or U14164 (N_14164,N_13936,N_13992);
xnor U14165 (N_14165,N_13610,N_13952);
and U14166 (N_14166,N_13720,N_13965);
xor U14167 (N_14167,N_13729,N_13682);
and U14168 (N_14168,N_13692,N_13639);
or U14169 (N_14169,N_13931,N_13894);
nor U14170 (N_14170,N_13604,N_13827);
or U14171 (N_14171,N_13893,N_13637);
and U14172 (N_14172,N_13603,N_13676);
xor U14173 (N_14173,N_13717,N_13743);
xor U14174 (N_14174,N_13733,N_13924);
or U14175 (N_14175,N_13638,N_13988);
nand U14176 (N_14176,N_13987,N_13730);
nand U14177 (N_14177,N_13882,N_13995);
or U14178 (N_14178,N_13862,N_13704);
xnor U14179 (N_14179,N_13619,N_13649);
or U14180 (N_14180,N_13666,N_13890);
nand U14181 (N_14181,N_13974,N_13809);
xor U14182 (N_14182,N_13746,N_13779);
nand U14183 (N_14183,N_13677,N_13990);
nor U14184 (N_14184,N_13707,N_13917);
nand U14185 (N_14185,N_13972,N_13659);
nand U14186 (N_14186,N_13970,N_13766);
nand U14187 (N_14187,N_13700,N_13789);
and U14188 (N_14188,N_13887,N_13617);
xnor U14189 (N_14189,N_13956,N_13661);
nand U14190 (N_14190,N_13876,N_13732);
nor U14191 (N_14191,N_13934,N_13971);
nand U14192 (N_14192,N_13806,N_13770);
and U14193 (N_14193,N_13798,N_13632);
nand U14194 (N_14194,N_13959,N_13686);
and U14195 (N_14195,N_13695,N_13822);
xnor U14196 (N_14196,N_13899,N_13851);
and U14197 (N_14197,N_13802,N_13886);
and U14198 (N_14198,N_13943,N_13794);
nand U14199 (N_14199,N_13975,N_13901);
nor U14200 (N_14200,N_13804,N_13821);
xor U14201 (N_14201,N_13849,N_13841);
xor U14202 (N_14202,N_13720,N_13856);
or U14203 (N_14203,N_13943,N_13680);
xnor U14204 (N_14204,N_13768,N_13696);
xor U14205 (N_14205,N_13945,N_13650);
nor U14206 (N_14206,N_13995,N_13656);
and U14207 (N_14207,N_13791,N_13620);
and U14208 (N_14208,N_13975,N_13726);
nor U14209 (N_14209,N_13726,N_13881);
and U14210 (N_14210,N_13754,N_13903);
and U14211 (N_14211,N_13608,N_13890);
xor U14212 (N_14212,N_13810,N_13609);
or U14213 (N_14213,N_13934,N_13761);
xor U14214 (N_14214,N_13718,N_13966);
xnor U14215 (N_14215,N_13775,N_13992);
and U14216 (N_14216,N_13648,N_13887);
nor U14217 (N_14217,N_13993,N_13813);
nand U14218 (N_14218,N_13644,N_13694);
and U14219 (N_14219,N_13934,N_13799);
and U14220 (N_14220,N_13868,N_13975);
nor U14221 (N_14221,N_13947,N_13848);
nand U14222 (N_14222,N_13900,N_13944);
nor U14223 (N_14223,N_13891,N_13858);
or U14224 (N_14224,N_13956,N_13776);
nand U14225 (N_14225,N_13775,N_13923);
nand U14226 (N_14226,N_13788,N_13964);
or U14227 (N_14227,N_13718,N_13675);
and U14228 (N_14228,N_13803,N_13992);
and U14229 (N_14229,N_13871,N_13754);
and U14230 (N_14230,N_13964,N_13906);
xor U14231 (N_14231,N_13680,N_13658);
xnor U14232 (N_14232,N_13982,N_13951);
nand U14233 (N_14233,N_13877,N_13825);
nand U14234 (N_14234,N_13841,N_13647);
xnor U14235 (N_14235,N_13815,N_13833);
and U14236 (N_14236,N_13945,N_13851);
nand U14237 (N_14237,N_13736,N_13659);
nor U14238 (N_14238,N_13989,N_13956);
nor U14239 (N_14239,N_13918,N_13626);
and U14240 (N_14240,N_13721,N_13984);
xor U14241 (N_14241,N_13952,N_13741);
or U14242 (N_14242,N_13997,N_13629);
xnor U14243 (N_14243,N_13969,N_13716);
and U14244 (N_14244,N_13686,N_13919);
nand U14245 (N_14245,N_13662,N_13743);
and U14246 (N_14246,N_13970,N_13778);
nor U14247 (N_14247,N_13896,N_13655);
or U14248 (N_14248,N_13777,N_13648);
and U14249 (N_14249,N_13743,N_13850);
nor U14250 (N_14250,N_13963,N_13604);
nand U14251 (N_14251,N_13940,N_13931);
nand U14252 (N_14252,N_13871,N_13634);
nor U14253 (N_14253,N_13621,N_13790);
xnor U14254 (N_14254,N_13906,N_13831);
and U14255 (N_14255,N_13843,N_13921);
nand U14256 (N_14256,N_13907,N_13942);
and U14257 (N_14257,N_13980,N_13837);
nor U14258 (N_14258,N_13984,N_13604);
nor U14259 (N_14259,N_13873,N_13869);
nor U14260 (N_14260,N_13891,N_13618);
or U14261 (N_14261,N_13941,N_13617);
xnor U14262 (N_14262,N_13964,N_13756);
and U14263 (N_14263,N_13870,N_13853);
and U14264 (N_14264,N_13724,N_13634);
and U14265 (N_14265,N_13987,N_13815);
nor U14266 (N_14266,N_13783,N_13893);
nand U14267 (N_14267,N_13769,N_13609);
xor U14268 (N_14268,N_13780,N_13715);
or U14269 (N_14269,N_13715,N_13661);
nor U14270 (N_14270,N_13791,N_13877);
and U14271 (N_14271,N_13603,N_13788);
and U14272 (N_14272,N_13668,N_13682);
and U14273 (N_14273,N_13861,N_13949);
or U14274 (N_14274,N_13811,N_13845);
nor U14275 (N_14275,N_13985,N_13904);
and U14276 (N_14276,N_13922,N_13908);
or U14277 (N_14277,N_13788,N_13740);
nand U14278 (N_14278,N_13749,N_13826);
nand U14279 (N_14279,N_13916,N_13623);
nor U14280 (N_14280,N_13793,N_13702);
or U14281 (N_14281,N_13759,N_13822);
nor U14282 (N_14282,N_13917,N_13868);
xor U14283 (N_14283,N_13845,N_13754);
xnor U14284 (N_14284,N_13962,N_13659);
or U14285 (N_14285,N_13631,N_13790);
xor U14286 (N_14286,N_13966,N_13765);
nor U14287 (N_14287,N_13661,N_13971);
or U14288 (N_14288,N_13933,N_13866);
nand U14289 (N_14289,N_13897,N_13847);
xnor U14290 (N_14290,N_13678,N_13753);
nor U14291 (N_14291,N_13825,N_13713);
and U14292 (N_14292,N_13682,N_13905);
xnor U14293 (N_14293,N_13946,N_13645);
or U14294 (N_14294,N_13989,N_13984);
xor U14295 (N_14295,N_13828,N_13847);
nand U14296 (N_14296,N_13954,N_13765);
xor U14297 (N_14297,N_13935,N_13975);
xnor U14298 (N_14298,N_13725,N_13951);
xnor U14299 (N_14299,N_13823,N_13632);
and U14300 (N_14300,N_13867,N_13895);
xnor U14301 (N_14301,N_13627,N_13841);
and U14302 (N_14302,N_13978,N_13760);
xnor U14303 (N_14303,N_13900,N_13684);
nand U14304 (N_14304,N_13759,N_13996);
or U14305 (N_14305,N_13848,N_13731);
xnor U14306 (N_14306,N_13831,N_13962);
nand U14307 (N_14307,N_13739,N_13916);
or U14308 (N_14308,N_13674,N_13883);
and U14309 (N_14309,N_13769,N_13893);
and U14310 (N_14310,N_13839,N_13711);
xor U14311 (N_14311,N_13786,N_13973);
nand U14312 (N_14312,N_13715,N_13782);
xnor U14313 (N_14313,N_13837,N_13687);
nand U14314 (N_14314,N_13750,N_13715);
and U14315 (N_14315,N_13626,N_13643);
or U14316 (N_14316,N_13612,N_13822);
or U14317 (N_14317,N_13670,N_13967);
nor U14318 (N_14318,N_13702,N_13871);
nor U14319 (N_14319,N_13956,N_13690);
xor U14320 (N_14320,N_13966,N_13751);
nand U14321 (N_14321,N_13938,N_13690);
nor U14322 (N_14322,N_13911,N_13686);
xnor U14323 (N_14323,N_13931,N_13721);
nand U14324 (N_14324,N_13844,N_13923);
nor U14325 (N_14325,N_13913,N_13932);
nor U14326 (N_14326,N_13616,N_13602);
nor U14327 (N_14327,N_13958,N_13635);
xnor U14328 (N_14328,N_13868,N_13858);
nor U14329 (N_14329,N_13930,N_13607);
and U14330 (N_14330,N_13895,N_13672);
nand U14331 (N_14331,N_13874,N_13822);
nand U14332 (N_14332,N_13705,N_13657);
nand U14333 (N_14333,N_13936,N_13887);
nand U14334 (N_14334,N_13771,N_13919);
nor U14335 (N_14335,N_13728,N_13983);
nor U14336 (N_14336,N_13976,N_13890);
xnor U14337 (N_14337,N_13805,N_13998);
nor U14338 (N_14338,N_13919,N_13741);
nand U14339 (N_14339,N_13889,N_13677);
or U14340 (N_14340,N_13929,N_13802);
and U14341 (N_14341,N_13772,N_13899);
or U14342 (N_14342,N_13603,N_13659);
and U14343 (N_14343,N_13739,N_13658);
or U14344 (N_14344,N_13612,N_13929);
and U14345 (N_14345,N_13654,N_13824);
or U14346 (N_14346,N_13888,N_13708);
nor U14347 (N_14347,N_13649,N_13622);
nor U14348 (N_14348,N_13800,N_13919);
nand U14349 (N_14349,N_13607,N_13658);
nand U14350 (N_14350,N_13683,N_13939);
xnor U14351 (N_14351,N_13733,N_13761);
nor U14352 (N_14352,N_13798,N_13626);
xor U14353 (N_14353,N_13669,N_13836);
nand U14354 (N_14354,N_13627,N_13887);
and U14355 (N_14355,N_13706,N_13999);
or U14356 (N_14356,N_13716,N_13914);
nor U14357 (N_14357,N_13689,N_13956);
or U14358 (N_14358,N_13942,N_13817);
xor U14359 (N_14359,N_13847,N_13885);
and U14360 (N_14360,N_13903,N_13778);
nor U14361 (N_14361,N_13835,N_13846);
xnor U14362 (N_14362,N_13783,N_13755);
or U14363 (N_14363,N_13804,N_13858);
nor U14364 (N_14364,N_13954,N_13998);
nor U14365 (N_14365,N_13686,N_13830);
nor U14366 (N_14366,N_13785,N_13747);
xor U14367 (N_14367,N_13927,N_13747);
xor U14368 (N_14368,N_13859,N_13728);
and U14369 (N_14369,N_13719,N_13651);
nand U14370 (N_14370,N_13683,N_13695);
xor U14371 (N_14371,N_13862,N_13924);
nand U14372 (N_14372,N_13922,N_13932);
and U14373 (N_14373,N_13620,N_13921);
and U14374 (N_14374,N_13961,N_13855);
or U14375 (N_14375,N_13747,N_13911);
xor U14376 (N_14376,N_13765,N_13758);
nand U14377 (N_14377,N_13866,N_13610);
and U14378 (N_14378,N_13939,N_13677);
or U14379 (N_14379,N_13963,N_13896);
nand U14380 (N_14380,N_13629,N_13845);
or U14381 (N_14381,N_13663,N_13899);
or U14382 (N_14382,N_13710,N_13606);
nand U14383 (N_14383,N_13675,N_13607);
nor U14384 (N_14384,N_13954,N_13679);
nand U14385 (N_14385,N_13707,N_13696);
and U14386 (N_14386,N_13769,N_13896);
nor U14387 (N_14387,N_13666,N_13904);
and U14388 (N_14388,N_13877,N_13689);
and U14389 (N_14389,N_13939,N_13945);
nand U14390 (N_14390,N_13893,N_13681);
or U14391 (N_14391,N_13981,N_13936);
xor U14392 (N_14392,N_13626,N_13848);
nor U14393 (N_14393,N_13905,N_13890);
nor U14394 (N_14394,N_13664,N_13667);
and U14395 (N_14395,N_13756,N_13842);
nor U14396 (N_14396,N_13810,N_13722);
nand U14397 (N_14397,N_13994,N_13953);
and U14398 (N_14398,N_13869,N_13785);
nor U14399 (N_14399,N_13675,N_13891);
nor U14400 (N_14400,N_14362,N_14242);
nor U14401 (N_14401,N_14035,N_14328);
xnor U14402 (N_14402,N_14376,N_14190);
xnor U14403 (N_14403,N_14293,N_14222);
and U14404 (N_14404,N_14163,N_14147);
nand U14405 (N_14405,N_14036,N_14058);
nand U14406 (N_14406,N_14142,N_14378);
nand U14407 (N_14407,N_14168,N_14339);
xnor U14408 (N_14408,N_14223,N_14234);
nand U14409 (N_14409,N_14249,N_14096);
and U14410 (N_14410,N_14215,N_14026);
nor U14411 (N_14411,N_14108,N_14367);
or U14412 (N_14412,N_14233,N_14299);
nand U14413 (N_14413,N_14310,N_14101);
xor U14414 (N_14414,N_14064,N_14075);
xnor U14415 (N_14415,N_14079,N_14143);
or U14416 (N_14416,N_14010,N_14174);
or U14417 (N_14417,N_14192,N_14271);
xor U14418 (N_14418,N_14393,N_14103);
nor U14419 (N_14419,N_14259,N_14068);
xnor U14420 (N_14420,N_14279,N_14386);
or U14421 (N_14421,N_14349,N_14170);
or U14422 (N_14422,N_14235,N_14106);
nand U14423 (N_14423,N_14003,N_14176);
or U14424 (N_14424,N_14256,N_14304);
or U14425 (N_14425,N_14276,N_14063);
or U14426 (N_14426,N_14301,N_14159);
and U14427 (N_14427,N_14370,N_14098);
and U14428 (N_14428,N_14260,N_14216);
xnor U14429 (N_14429,N_14044,N_14125);
nor U14430 (N_14430,N_14070,N_14381);
nand U14431 (N_14431,N_14004,N_14384);
xor U14432 (N_14432,N_14173,N_14313);
xnor U14433 (N_14433,N_14320,N_14080);
nand U14434 (N_14434,N_14364,N_14206);
nand U14435 (N_14435,N_14205,N_14156);
nand U14436 (N_14436,N_14090,N_14247);
and U14437 (N_14437,N_14257,N_14072);
xor U14438 (N_14438,N_14071,N_14074);
and U14439 (N_14439,N_14111,N_14264);
and U14440 (N_14440,N_14179,N_14254);
nand U14441 (N_14441,N_14104,N_14140);
nand U14442 (N_14442,N_14011,N_14252);
and U14443 (N_14443,N_14099,N_14197);
nor U14444 (N_14444,N_14239,N_14387);
nand U14445 (N_14445,N_14018,N_14088);
xor U14446 (N_14446,N_14228,N_14373);
nand U14447 (N_14447,N_14357,N_14291);
or U14448 (N_14448,N_14059,N_14160);
and U14449 (N_14449,N_14199,N_14014);
and U14450 (N_14450,N_14017,N_14137);
nand U14451 (N_14451,N_14081,N_14269);
xor U14452 (N_14452,N_14396,N_14077);
nand U14453 (N_14453,N_14345,N_14133);
or U14454 (N_14454,N_14078,N_14255);
xnor U14455 (N_14455,N_14231,N_14052);
or U14456 (N_14456,N_14122,N_14283);
nand U14457 (N_14457,N_14214,N_14016);
xnor U14458 (N_14458,N_14353,N_14175);
xor U14459 (N_14459,N_14020,N_14289);
and U14460 (N_14460,N_14038,N_14308);
nand U14461 (N_14461,N_14161,N_14377);
and U14462 (N_14462,N_14209,N_14177);
and U14463 (N_14463,N_14095,N_14251);
nor U14464 (N_14464,N_14180,N_14261);
or U14465 (N_14465,N_14329,N_14287);
and U14466 (N_14466,N_14045,N_14332);
xor U14467 (N_14467,N_14262,N_14397);
nor U14468 (N_14468,N_14278,N_14292);
xor U14469 (N_14469,N_14097,N_14100);
xor U14470 (N_14470,N_14273,N_14398);
nand U14471 (N_14471,N_14050,N_14226);
or U14472 (N_14472,N_14282,N_14340);
nor U14473 (N_14473,N_14363,N_14076);
or U14474 (N_14474,N_14394,N_14007);
and U14475 (N_14475,N_14374,N_14105);
nor U14476 (N_14476,N_14109,N_14126);
nor U14477 (N_14477,N_14132,N_14030);
or U14478 (N_14478,N_14290,N_14224);
xor U14479 (N_14479,N_14022,N_14366);
and U14480 (N_14480,N_14281,N_14047);
nand U14481 (N_14481,N_14110,N_14025);
xor U14482 (N_14482,N_14246,N_14321);
or U14483 (N_14483,N_14388,N_14391);
and U14484 (N_14484,N_14032,N_14189);
nor U14485 (N_14485,N_14024,N_14102);
or U14486 (N_14486,N_14136,N_14371);
and U14487 (N_14487,N_14382,N_14324);
nand U14488 (N_14488,N_14225,N_14083);
nand U14489 (N_14489,N_14297,N_14361);
nand U14490 (N_14490,N_14054,N_14336);
nand U14491 (N_14491,N_14303,N_14187);
and U14492 (N_14492,N_14027,N_14277);
or U14493 (N_14493,N_14375,N_14389);
and U14494 (N_14494,N_14023,N_14243);
nor U14495 (N_14495,N_14322,N_14348);
or U14496 (N_14496,N_14130,N_14157);
nand U14497 (N_14497,N_14129,N_14150);
nand U14498 (N_14498,N_14335,N_14270);
xnor U14499 (N_14499,N_14040,N_14116);
xor U14500 (N_14500,N_14316,N_14155);
and U14501 (N_14501,N_14236,N_14146);
or U14502 (N_14502,N_14358,N_14334);
xor U14503 (N_14503,N_14067,N_14057);
nand U14504 (N_14504,N_14092,N_14201);
nand U14505 (N_14505,N_14148,N_14220);
xnor U14506 (N_14506,N_14268,N_14144);
xor U14507 (N_14507,N_14019,N_14114);
and U14508 (N_14508,N_14238,N_14089);
nand U14509 (N_14509,N_14300,N_14346);
and U14510 (N_14510,N_14048,N_14186);
xnor U14511 (N_14511,N_14341,N_14009);
and U14512 (N_14512,N_14274,N_14240);
xor U14513 (N_14513,N_14219,N_14178);
nor U14514 (N_14514,N_14141,N_14202);
xnor U14515 (N_14515,N_14244,N_14123);
xor U14516 (N_14516,N_14165,N_14149);
nor U14517 (N_14517,N_14284,N_14311);
or U14518 (N_14518,N_14385,N_14093);
xor U14519 (N_14519,N_14194,N_14039);
nand U14520 (N_14520,N_14253,N_14280);
and U14521 (N_14521,N_14086,N_14041);
and U14522 (N_14522,N_14113,N_14356);
or U14523 (N_14523,N_14008,N_14317);
xor U14524 (N_14524,N_14073,N_14285);
nand U14525 (N_14525,N_14182,N_14350);
nor U14526 (N_14526,N_14200,N_14193);
xnor U14527 (N_14527,N_14135,N_14119);
and U14528 (N_14528,N_14213,N_14062);
nand U14529 (N_14529,N_14245,N_14359);
nor U14530 (N_14530,N_14055,N_14368);
or U14531 (N_14531,N_14066,N_14272);
or U14532 (N_14532,N_14087,N_14318);
nor U14533 (N_14533,N_14124,N_14399);
and U14534 (N_14534,N_14028,N_14162);
or U14535 (N_14535,N_14037,N_14001);
xnor U14536 (N_14536,N_14158,N_14208);
xor U14537 (N_14537,N_14217,N_14131);
xor U14538 (N_14538,N_14326,N_14218);
nand U14539 (N_14539,N_14296,N_14085);
nand U14540 (N_14540,N_14115,N_14265);
xnor U14541 (N_14541,N_14395,N_14204);
nor U14542 (N_14542,N_14049,N_14171);
nor U14543 (N_14543,N_14166,N_14331);
xor U14544 (N_14544,N_14307,N_14379);
nor U14545 (N_14545,N_14034,N_14065);
nor U14546 (N_14546,N_14319,N_14365);
and U14547 (N_14547,N_14241,N_14372);
or U14548 (N_14548,N_14330,N_14195);
xor U14549 (N_14549,N_14380,N_14053);
or U14550 (N_14550,N_14043,N_14060);
or U14551 (N_14551,N_14069,N_14061);
and U14552 (N_14552,N_14232,N_14383);
or U14553 (N_14553,N_14390,N_14327);
and U14554 (N_14554,N_14342,N_14112);
xor U14555 (N_14555,N_14188,N_14121);
nand U14556 (N_14556,N_14145,N_14084);
and U14557 (N_14557,N_14056,N_14138);
xnor U14558 (N_14558,N_14139,N_14312);
or U14559 (N_14559,N_14298,N_14012);
nand U14560 (N_14560,N_14351,N_14000);
nor U14561 (N_14561,N_14082,N_14333);
or U14562 (N_14562,N_14306,N_14185);
xor U14563 (N_14563,N_14031,N_14230);
xnor U14564 (N_14564,N_14347,N_14352);
and U14565 (N_14565,N_14275,N_14325);
and U14566 (N_14566,N_14033,N_14127);
or U14567 (N_14567,N_14198,N_14196);
nand U14568 (N_14568,N_14152,N_14302);
or U14569 (N_14569,N_14315,N_14250);
xnor U14570 (N_14570,N_14210,N_14128);
or U14571 (N_14571,N_14183,N_14263);
xnor U14572 (N_14572,N_14323,N_14172);
nand U14573 (N_14573,N_14118,N_14294);
nor U14574 (N_14574,N_14151,N_14344);
or U14575 (N_14575,N_14091,N_14046);
nor U14576 (N_14576,N_14288,N_14153);
or U14577 (N_14577,N_14221,N_14360);
nor U14578 (N_14578,N_14184,N_14164);
nand U14579 (N_14579,N_14369,N_14167);
nand U14580 (N_14580,N_14021,N_14029);
and U14581 (N_14581,N_14203,N_14258);
nand U14582 (N_14582,N_14229,N_14134);
nand U14583 (N_14583,N_14013,N_14343);
and U14584 (N_14584,N_14337,N_14314);
or U14585 (N_14585,N_14107,N_14211);
nand U14586 (N_14586,N_14338,N_14207);
xor U14587 (N_14587,N_14002,N_14094);
xor U14588 (N_14588,N_14051,N_14248);
or U14589 (N_14589,N_14169,N_14117);
or U14590 (N_14590,N_14305,N_14237);
or U14591 (N_14591,N_14005,N_14355);
and U14592 (N_14592,N_14227,N_14286);
xnor U14593 (N_14593,N_14006,N_14015);
or U14594 (N_14594,N_14212,N_14120);
nor U14595 (N_14595,N_14295,N_14309);
xor U14596 (N_14596,N_14154,N_14354);
and U14597 (N_14597,N_14267,N_14392);
or U14598 (N_14598,N_14266,N_14191);
and U14599 (N_14599,N_14042,N_14181);
or U14600 (N_14600,N_14329,N_14000);
nor U14601 (N_14601,N_14180,N_14012);
or U14602 (N_14602,N_14239,N_14357);
nand U14603 (N_14603,N_14161,N_14328);
nor U14604 (N_14604,N_14112,N_14207);
or U14605 (N_14605,N_14381,N_14148);
nand U14606 (N_14606,N_14392,N_14043);
nand U14607 (N_14607,N_14354,N_14237);
or U14608 (N_14608,N_14229,N_14228);
nand U14609 (N_14609,N_14337,N_14322);
nor U14610 (N_14610,N_14090,N_14048);
xnor U14611 (N_14611,N_14130,N_14143);
xor U14612 (N_14612,N_14086,N_14016);
nor U14613 (N_14613,N_14164,N_14249);
nand U14614 (N_14614,N_14224,N_14141);
nand U14615 (N_14615,N_14120,N_14297);
nor U14616 (N_14616,N_14294,N_14124);
nor U14617 (N_14617,N_14319,N_14348);
nand U14618 (N_14618,N_14263,N_14197);
xnor U14619 (N_14619,N_14020,N_14053);
and U14620 (N_14620,N_14214,N_14070);
nand U14621 (N_14621,N_14238,N_14192);
nor U14622 (N_14622,N_14211,N_14296);
xnor U14623 (N_14623,N_14015,N_14343);
and U14624 (N_14624,N_14288,N_14155);
or U14625 (N_14625,N_14149,N_14338);
or U14626 (N_14626,N_14293,N_14215);
or U14627 (N_14627,N_14045,N_14052);
nand U14628 (N_14628,N_14035,N_14177);
or U14629 (N_14629,N_14354,N_14147);
nand U14630 (N_14630,N_14022,N_14347);
xnor U14631 (N_14631,N_14055,N_14179);
xnor U14632 (N_14632,N_14172,N_14383);
or U14633 (N_14633,N_14234,N_14341);
or U14634 (N_14634,N_14354,N_14075);
or U14635 (N_14635,N_14156,N_14332);
nand U14636 (N_14636,N_14171,N_14098);
nand U14637 (N_14637,N_14373,N_14071);
xor U14638 (N_14638,N_14243,N_14116);
nor U14639 (N_14639,N_14269,N_14396);
and U14640 (N_14640,N_14375,N_14316);
and U14641 (N_14641,N_14120,N_14208);
nand U14642 (N_14642,N_14360,N_14180);
nand U14643 (N_14643,N_14249,N_14172);
xnor U14644 (N_14644,N_14078,N_14387);
and U14645 (N_14645,N_14011,N_14187);
or U14646 (N_14646,N_14264,N_14282);
and U14647 (N_14647,N_14177,N_14206);
or U14648 (N_14648,N_14071,N_14225);
or U14649 (N_14649,N_14028,N_14178);
nor U14650 (N_14650,N_14290,N_14119);
nor U14651 (N_14651,N_14351,N_14302);
and U14652 (N_14652,N_14297,N_14101);
nor U14653 (N_14653,N_14353,N_14164);
nand U14654 (N_14654,N_14249,N_14178);
or U14655 (N_14655,N_14270,N_14024);
xnor U14656 (N_14656,N_14105,N_14057);
xnor U14657 (N_14657,N_14315,N_14247);
xor U14658 (N_14658,N_14333,N_14300);
and U14659 (N_14659,N_14270,N_14380);
xnor U14660 (N_14660,N_14271,N_14074);
or U14661 (N_14661,N_14296,N_14398);
nand U14662 (N_14662,N_14379,N_14122);
or U14663 (N_14663,N_14234,N_14153);
xor U14664 (N_14664,N_14118,N_14367);
or U14665 (N_14665,N_14113,N_14387);
nor U14666 (N_14666,N_14276,N_14262);
xnor U14667 (N_14667,N_14191,N_14176);
or U14668 (N_14668,N_14096,N_14346);
and U14669 (N_14669,N_14386,N_14112);
nor U14670 (N_14670,N_14219,N_14321);
or U14671 (N_14671,N_14384,N_14083);
nand U14672 (N_14672,N_14215,N_14104);
and U14673 (N_14673,N_14281,N_14039);
nand U14674 (N_14674,N_14250,N_14090);
nand U14675 (N_14675,N_14320,N_14079);
and U14676 (N_14676,N_14279,N_14382);
and U14677 (N_14677,N_14146,N_14048);
nand U14678 (N_14678,N_14103,N_14289);
or U14679 (N_14679,N_14212,N_14198);
and U14680 (N_14680,N_14097,N_14116);
and U14681 (N_14681,N_14100,N_14383);
or U14682 (N_14682,N_14108,N_14272);
or U14683 (N_14683,N_14392,N_14271);
or U14684 (N_14684,N_14304,N_14236);
xor U14685 (N_14685,N_14127,N_14371);
or U14686 (N_14686,N_14327,N_14381);
nand U14687 (N_14687,N_14179,N_14289);
xor U14688 (N_14688,N_14142,N_14049);
nor U14689 (N_14689,N_14018,N_14019);
nor U14690 (N_14690,N_14052,N_14088);
xnor U14691 (N_14691,N_14168,N_14072);
and U14692 (N_14692,N_14018,N_14221);
and U14693 (N_14693,N_14389,N_14032);
nand U14694 (N_14694,N_14198,N_14219);
nor U14695 (N_14695,N_14001,N_14265);
and U14696 (N_14696,N_14251,N_14126);
or U14697 (N_14697,N_14110,N_14070);
nand U14698 (N_14698,N_14320,N_14226);
xor U14699 (N_14699,N_14315,N_14100);
xor U14700 (N_14700,N_14122,N_14193);
and U14701 (N_14701,N_14101,N_14220);
nor U14702 (N_14702,N_14115,N_14208);
nand U14703 (N_14703,N_14346,N_14282);
nor U14704 (N_14704,N_14259,N_14021);
and U14705 (N_14705,N_14003,N_14263);
nor U14706 (N_14706,N_14139,N_14150);
xor U14707 (N_14707,N_14344,N_14126);
or U14708 (N_14708,N_14300,N_14271);
or U14709 (N_14709,N_14020,N_14047);
nor U14710 (N_14710,N_14129,N_14109);
xor U14711 (N_14711,N_14045,N_14162);
xnor U14712 (N_14712,N_14395,N_14055);
nand U14713 (N_14713,N_14188,N_14300);
and U14714 (N_14714,N_14279,N_14208);
or U14715 (N_14715,N_14099,N_14140);
nor U14716 (N_14716,N_14111,N_14335);
and U14717 (N_14717,N_14325,N_14318);
and U14718 (N_14718,N_14210,N_14107);
nor U14719 (N_14719,N_14250,N_14396);
nand U14720 (N_14720,N_14335,N_14191);
nand U14721 (N_14721,N_14350,N_14336);
xnor U14722 (N_14722,N_14337,N_14343);
nor U14723 (N_14723,N_14041,N_14248);
nand U14724 (N_14724,N_14320,N_14195);
xnor U14725 (N_14725,N_14067,N_14019);
and U14726 (N_14726,N_14258,N_14065);
nor U14727 (N_14727,N_14107,N_14169);
xnor U14728 (N_14728,N_14265,N_14293);
xor U14729 (N_14729,N_14229,N_14221);
nand U14730 (N_14730,N_14345,N_14108);
xor U14731 (N_14731,N_14291,N_14151);
xnor U14732 (N_14732,N_14287,N_14291);
or U14733 (N_14733,N_14166,N_14274);
and U14734 (N_14734,N_14373,N_14236);
nor U14735 (N_14735,N_14168,N_14100);
or U14736 (N_14736,N_14094,N_14292);
xor U14737 (N_14737,N_14170,N_14075);
and U14738 (N_14738,N_14320,N_14382);
nand U14739 (N_14739,N_14034,N_14185);
and U14740 (N_14740,N_14175,N_14257);
nand U14741 (N_14741,N_14036,N_14216);
and U14742 (N_14742,N_14082,N_14270);
nor U14743 (N_14743,N_14261,N_14113);
or U14744 (N_14744,N_14052,N_14195);
and U14745 (N_14745,N_14192,N_14326);
and U14746 (N_14746,N_14050,N_14038);
and U14747 (N_14747,N_14355,N_14047);
and U14748 (N_14748,N_14165,N_14157);
xnor U14749 (N_14749,N_14229,N_14145);
nor U14750 (N_14750,N_14027,N_14162);
nor U14751 (N_14751,N_14104,N_14185);
nand U14752 (N_14752,N_14365,N_14037);
xnor U14753 (N_14753,N_14117,N_14109);
nand U14754 (N_14754,N_14210,N_14019);
xor U14755 (N_14755,N_14367,N_14105);
or U14756 (N_14756,N_14330,N_14303);
nor U14757 (N_14757,N_14354,N_14239);
nand U14758 (N_14758,N_14044,N_14052);
nand U14759 (N_14759,N_14149,N_14122);
xnor U14760 (N_14760,N_14173,N_14136);
nor U14761 (N_14761,N_14343,N_14180);
nor U14762 (N_14762,N_14197,N_14366);
or U14763 (N_14763,N_14334,N_14337);
nor U14764 (N_14764,N_14192,N_14243);
or U14765 (N_14765,N_14086,N_14206);
or U14766 (N_14766,N_14039,N_14135);
or U14767 (N_14767,N_14363,N_14188);
xor U14768 (N_14768,N_14245,N_14244);
nor U14769 (N_14769,N_14082,N_14339);
nor U14770 (N_14770,N_14169,N_14257);
nor U14771 (N_14771,N_14112,N_14074);
xor U14772 (N_14772,N_14345,N_14312);
or U14773 (N_14773,N_14231,N_14054);
or U14774 (N_14774,N_14399,N_14100);
and U14775 (N_14775,N_14192,N_14352);
or U14776 (N_14776,N_14083,N_14184);
and U14777 (N_14777,N_14324,N_14152);
and U14778 (N_14778,N_14269,N_14283);
and U14779 (N_14779,N_14228,N_14301);
nand U14780 (N_14780,N_14277,N_14047);
nand U14781 (N_14781,N_14009,N_14067);
xor U14782 (N_14782,N_14197,N_14034);
nor U14783 (N_14783,N_14053,N_14006);
xnor U14784 (N_14784,N_14127,N_14266);
nor U14785 (N_14785,N_14169,N_14281);
nand U14786 (N_14786,N_14137,N_14366);
and U14787 (N_14787,N_14238,N_14149);
xor U14788 (N_14788,N_14357,N_14170);
or U14789 (N_14789,N_14005,N_14387);
xor U14790 (N_14790,N_14020,N_14229);
nand U14791 (N_14791,N_14199,N_14348);
nand U14792 (N_14792,N_14126,N_14138);
xor U14793 (N_14793,N_14359,N_14022);
xnor U14794 (N_14794,N_14195,N_14291);
nor U14795 (N_14795,N_14120,N_14336);
and U14796 (N_14796,N_14311,N_14190);
and U14797 (N_14797,N_14354,N_14199);
and U14798 (N_14798,N_14375,N_14202);
xor U14799 (N_14799,N_14154,N_14350);
and U14800 (N_14800,N_14593,N_14561);
and U14801 (N_14801,N_14491,N_14746);
or U14802 (N_14802,N_14594,N_14676);
nand U14803 (N_14803,N_14460,N_14513);
nor U14804 (N_14804,N_14642,N_14688);
nor U14805 (N_14805,N_14505,N_14464);
nand U14806 (N_14806,N_14629,N_14651);
or U14807 (N_14807,N_14478,N_14672);
nor U14808 (N_14808,N_14702,N_14736);
or U14809 (N_14809,N_14683,N_14472);
or U14810 (N_14810,N_14426,N_14536);
nor U14811 (N_14811,N_14776,N_14582);
or U14812 (N_14812,N_14681,N_14504);
or U14813 (N_14813,N_14752,N_14555);
or U14814 (N_14814,N_14481,N_14753);
nand U14815 (N_14815,N_14442,N_14645);
nor U14816 (N_14816,N_14525,N_14423);
or U14817 (N_14817,N_14579,N_14732);
xor U14818 (N_14818,N_14503,N_14610);
nor U14819 (N_14819,N_14413,N_14599);
nor U14820 (N_14820,N_14775,N_14737);
or U14821 (N_14821,N_14511,N_14720);
nor U14822 (N_14822,N_14495,N_14425);
xor U14823 (N_14823,N_14741,N_14778);
nor U14824 (N_14824,N_14592,N_14527);
or U14825 (N_14825,N_14714,N_14412);
xor U14826 (N_14826,N_14595,N_14479);
nor U14827 (N_14827,N_14760,N_14493);
or U14828 (N_14828,N_14608,N_14763);
and U14829 (N_14829,N_14439,N_14666);
xor U14830 (N_14830,N_14443,N_14695);
xor U14831 (N_14831,N_14535,N_14449);
and U14832 (N_14832,N_14411,N_14768);
nor U14833 (N_14833,N_14656,N_14545);
nand U14834 (N_14834,N_14745,N_14438);
or U14835 (N_14835,N_14414,N_14719);
nand U14836 (N_14836,N_14793,N_14541);
and U14837 (N_14837,N_14687,N_14771);
nand U14838 (N_14838,N_14617,N_14574);
and U14839 (N_14839,N_14640,N_14606);
and U14840 (N_14840,N_14454,N_14557);
and U14841 (N_14841,N_14416,N_14469);
or U14842 (N_14842,N_14697,N_14609);
nand U14843 (N_14843,N_14616,N_14772);
xor U14844 (N_14844,N_14669,N_14436);
nand U14845 (N_14845,N_14601,N_14529);
nor U14846 (N_14846,N_14713,N_14615);
nor U14847 (N_14847,N_14430,N_14446);
or U14848 (N_14848,N_14770,N_14694);
nor U14849 (N_14849,N_14643,N_14466);
and U14850 (N_14850,N_14739,N_14415);
nor U14851 (N_14851,N_14539,N_14731);
nor U14852 (N_14852,N_14708,N_14665);
nor U14853 (N_14853,N_14647,N_14586);
nor U14854 (N_14854,N_14507,N_14626);
and U14855 (N_14855,N_14791,N_14705);
nand U14856 (N_14856,N_14562,N_14653);
xor U14857 (N_14857,N_14692,N_14649);
nor U14858 (N_14858,N_14754,N_14543);
xor U14859 (N_14859,N_14475,N_14785);
and U14860 (N_14860,N_14497,N_14581);
and U14861 (N_14861,N_14567,N_14409);
nand U14862 (N_14862,N_14554,N_14583);
xnor U14863 (N_14863,N_14747,N_14421);
nor U14864 (N_14864,N_14773,N_14428);
nand U14865 (N_14865,N_14678,N_14646);
nor U14866 (N_14866,N_14765,N_14758);
or U14867 (N_14867,N_14476,N_14769);
and U14868 (N_14868,N_14634,N_14703);
nand U14869 (N_14869,N_14548,N_14575);
xnor U14870 (N_14870,N_14502,N_14509);
and U14871 (N_14871,N_14477,N_14734);
xnor U14872 (N_14872,N_14531,N_14743);
or U14873 (N_14873,N_14447,N_14696);
and U14874 (N_14874,N_14405,N_14499);
nand U14875 (N_14875,N_14777,N_14482);
nor U14876 (N_14876,N_14591,N_14795);
nor U14877 (N_14877,N_14598,N_14794);
nor U14878 (N_14878,N_14709,N_14526);
nand U14879 (N_14879,N_14686,N_14780);
or U14880 (N_14880,N_14455,N_14550);
or U14881 (N_14881,N_14623,N_14500);
xnor U14882 (N_14882,N_14691,N_14418);
or U14883 (N_14883,N_14546,N_14783);
xnor U14884 (N_14884,N_14755,N_14596);
and U14885 (N_14885,N_14799,N_14589);
nor U14886 (N_14886,N_14611,N_14724);
or U14887 (N_14887,N_14667,N_14661);
nor U14888 (N_14888,N_14680,N_14684);
nor U14889 (N_14889,N_14727,N_14718);
and U14890 (N_14890,N_14757,N_14501);
nor U14891 (N_14891,N_14722,N_14587);
nand U14892 (N_14892,N_14624,N_14729);
xor U14893 (N_14893,N_14600,N_14489);
xor U14894 (N_14894,N_14756,N_14534);
xnor U14895 (N_14895,N_14671,N_14796);
and U14896 (N_14896,N_14655,N_14621);
and U14897 (N_14897,N_14564,N_14792);
xor U14898 (N_14898,N_14662,N_14515);
or U14899 (N_14899,N_14588,N_14401);
or U14900 (N_14900,N_14690,N_14612);
or U14901 (N_14901,N_14506,N_14675);
xor U14902 (N_14902,N_14560,N_14700);
xnor U14903 (N_14903,N_14578,N_14622);
and U14904 (N_14904,N_14450,N_14512);
nand U14905 (N_14905,N_14528,N_14432);
and U14906 (N_14906,N_14761,N_14518);
or U14907 (N_14907,N_14551,N_14540);
and U14908 (N_14908,N_14429,N_14523);
or U14909 (N_14909,N_14614,N_14677);
xor U14910 (N_14910,N_14648,N_14427);
and U14911 (N_14911,N_14571,N_14408);
nor U14912 (N_14912,N_14577,N_14419);
or U14913 (N_14913,N_14580,N_14715);
and U14914 (N_14914,N_14701,N_14749);
and U14915 (N_14915,N_14522,N_14635);
nor U14916 (N_14916,N_14462,N_14538);
nand U14917 (N_14917,N_14733,N_14782);
and U14918 (N_14918,N_14572,N_14404);
nand U14919 (N_14919,N_14558,N_14605);
xnor U14920 (N_14920,N_14762,N_14448);
and U14921 (N_14921,N_14748,N_14641);
nor U14922 (N_14922,N_14433,N_14537);
xor U14923 (N_14923,N_14471,N_14553);
nand U14924 (N_14924,N_14636,N_14459);
and U14925 (N_14925,N_14767,N_14682);
and U14926 (N_14926,N_14742,N_14650);
xor U14927 (N_14927,N_14422,N_14652);
nand U14928 (N_14928,N_14585,N_14717);
xnor U14929 (N_14929,N_14547,N_14674);
and U14930 (N_14930,N_14787,N_14565);
and U14931 (N_14931,N_14788,N_14668);
or U14932 (N_14932,N_14552,N_14532);
nor U14933 (N_14933,N_14618,N_14781);
xor U14934 (N_14934,N_14620,N_14723);
and U14935 (N_14935,N_14639,N_14437);
or U14936 (N_14936,N_14638,N_14797);
and U14937 (N_14937,N_14607,N_14420);
and U14938 (N_14938,N_14498,N_14631);
nor U14939 (N_14939,N_14402,N_14519);
nor U14940 (N_14940,N_14710,N_14485);
and U14941 (N_14941,N_14603,N_14698);
nor U14942 (N_14942,N_14467,N_14706);
nor U14943 (N_14943,N_14657,N_14726);
xor U14944 (N_14944,N_14711,N_14590);
xor U14945 (N_14945,N_14625,N_14728);
nor U14946 (N_14946,N_14452,N_14533);
xor U14947 (N_14947,N_14707,N_14451);
xnor U14948 (N_14948,N_14510,N_14453);
nor U14949 (N_14949,N_14759,N_14417);
nand U14950 (N_14950,N_14530,N_14400);
and U14951 (N_14951,N_14632,N_14474);
and U14952 (N_14952,N_14735,N_14434);
or U14953 (N_14953,N_14764,N_14663);
xnor U14954 (N_14954,N_14486,N_14544);
or U14955 (N_14955,N_14689,N_14480);
and U14956 (N_14956,N_14597,N_14604);
or U14957 (N_14957,N_14628,N_14484);
nand U14958 (N_14958,N_14670,N_14660);
nor U14959 (N_14959,N_14570,N_14542);
nor U14960 (N_14960,N_14738,N_14789);
nand U14961 (N_14961,N_14457,N_14798);
xor U14962 (N_14962,N_14627,N_14633);
and U14963 (N_14963,N_14483,N_14613);
nor U14964 (N_14964,N_14431,N_14524);
or U14965 (N_14965,N_14468,N_14549);
xnor U14966 (N_14966,N_14716,N_14630);
nor U14967 (N_14967,N_14712,N_14410);
and U14968 (N_14968,N_14744,N_14556);
nand U14969 (N_14969,N_14568,N_14751);
nor U14970 (N_14970,N_14424,N_14463);
nand U14971 (N_14971,N_14569,N_14573);
nand U14972 (N_14972,N_14784,N_14654);
xnor U14973 (N_14973,N_14786,N_14659);
and U14974 (N_14974,N_14508,N_14465);
and U14975 (N_14975,N_14725,N_14490);
or U14976 (N_14976,N_14441,N_14407);
or U14977 (N_14977,N_14699,N_14487);
and U14978 (N_14978,N_14514,N_14496);
xor U14979 (N_14979,N_14435,N_14521);
xnor U14980 (N_14980,N_14456,N_14461);
and U14981 (N_14981,N_14602,N_14492);
xnor U14982 (N_14982,N_14664,N_14559);
or U14983 (N_14983,N_14566,N_14704);
nand U14984 (N_14984,N_14619,N_14494);
or U14985 (N_14985,N_14693,N_14685);
xnor U14986 (N_14986,N_14721,N_14445);
or U14987 (N_14987,N_14458,N_14774);
or U14988 (N_14988,N_14779,N_14740);
and U14989 (N_14989,N_14406,N_14658);
and U14990 (N_14990,N_14520,N_14730);
and U14991 (N_14991,N_14563,N_14473);
and U14992 (N_14992,N_14488,N_14444);
nand U14993 (N_14993,N_14576,N_14644);
or U14994 (N_14994,N_14790,N_14470);
or U14995 (N_14995,N_14673,N_14750);
and U14996 (N_14996,N_14516,N_14679);
nor U14997 (N_14997,N_14403,N_14637);
xnor U14998 (N_14998,N_14517,N_14766);
or U14999 (N_14999,N_14440,N_14584);
or U15000 (N_15000,N_14569,N_14710);
or U15001 (N_15001,N_14477,N_14468);
or U15002 (N_15002,N_14455,N_14462);
or U15003 (N_15003,N_14469,N_14665);
nor U15004 (N_15004,N_14625,N_14706);
nand U15005 (N_15005,N_14732,N_14607);
nor U15006 (N_15006,N_14713,N_14604);
or U15007 (N_15007,N_14653,N_14711);
or U15008 (N_15008,N_14648,N_14501);
nor U15009 (N_15009,N_14682,N_14508);
nand U15010 (N_15010,N_14666,N_14523);
and U15011 (N_15011,N_14480,N_14799);
nand U15012 (N_15012,N_14519,N_14671);
or U15013 (N_15013,N_14725,N_14776);
nand U15014 (N_15014,N_14442,N_14691);
and U15015 (N_15015,N_14546,N_14583);
and U15016 (N_15016,N_14507,N_14480);
or U15017 (N_15017,N_14622,N_14510);
nand U15018 (N_15018,N_14663,N_14471);
or U15019 (N_15019,N_14522,N_14416);
or U15020 (N_15020,N_14580,N_14767);
nor U15021 (N_15021,N_14718,N_14665);
nand U15022 (N_15022,N_14712,N_14797);
nor U15023 (N_15023,N_14519,N_14633);
or U15024 (N_15024,N_14667,N_14658);
nor U15025 (N_15025,N_14435,N_14491);
and U15026 (N_15026,N_14500,N_14491);
nand U15027 (N_15027,N_14472,N_14741);
and U15028 (N_15028,N_14518,N_14654);
or U15029 (N_15029,N_14570,N_14613);
and U15030 (N_15030,N_14513,N_14588);
nor U15031 (N_15031,N_14573,N_14427);
xor U15032 (N_15032,N_14539,N_14583);
or U15033 (N_15033,N_14736,N_14738);
or U15034 (N_15034,N_14522,N_14458);
or U15035 (N_15035,N_14523,N_14547);
and U15036 (N_15036,N_14552,N_14693);
or U15037 (N_15037,N_14567,N_14757);
nor U15038 (N_15038,N_14642,N_14787);
xnor U15039 (N_15039,N_14497,N_14408);
or U15040 (N_15040,N_14702,N_14529);
and U15041 (N_15041,N_14439,N_14420);
nor U15042 (N_15042,N_14591,N_14607);
or U15043 (N_15043,N_14507,N_14764);
nor U15044 (N_15044,N_14593,N_14518);
and U15045 (N_15045,N_14567,N_14632);
xnor U15046 (N_15046,N_14577,N_14770);
xnor U15047 (N_15047,N_14782,N_14440);
and U15048 (N_15048,N_14710,N_14470);
and U15049 (N_15049,N_14494,N_14401);
or U15050 (N_15050,N_14718,N_14684);
or U15051 (N_15051,N_14742,N_14492);
nor U15052 (N_15052,N_14530,N_14418);
nand U15053 (N_15053,N_14528,N_14522);
or U15054 (N_15054,N_14681,N_14463);
or U15055 (N_15055,N_14406,N_14733);
and U15056 (N_15056,N_14570,N_14643);
and U15057 (N_15057,N_14403,N_14743);
nand U15058 (N_15058,N_14593,N_14731);
and U15059 (N_15059,N_14684,N_14529);
or U15060 (N_15060,N_14769,N_14572);
xor U15061 (N_15061,N_14547,N_14573);
xor U15062 (N_15062,N_14574,N_14591);
nand U15063 (N_15063,N_14561,N_14712);
nand U15064 (N_15064,N_14445,N_14581);
or U15065 (N_15065,N_14469,N_14700);
and U15066 (N_15066,N_14541,N_14538);
or U15067 (N_15067,N_14534,N_14676);
and U15068 (N_15068,N_14712,N_14441);
nand U15069 (N_15069,N_14414,N_14490);
nor U15070 (N_15070,N_14488,N_14552);
nor U15071 (N_15071,N_14687,N_14616);
or U15072 (N_15072,N_14463,N_14699);
xor U15073 (N_15073,N_14790,N_14526);
nor U15074 (N_15074,N_14595,N_14745);
xor U15075 (N_15075,N_14726,N_14430);
nor U15076 (N_15076,N_14753,N_14757);
and U15077 (N_15077,N_14554,N_14755);
nor U15078 (N_15078,N_14575,N_14755);
nor U15079 (N_15079,N_14521,N_14732);
xor U15080 (N_15080,N_14712,N_14620);
xor U15081 (N_15081,N_14773,N_14616);
nand U15082 (N_15082,N_14725,N_14753);
nand U15083 (N_15083,N_14698,N_14651);
and U15084 (N_15084,N_14630,N_14751);
or U15085 (N_15085,N_14412,N_14680);
xnor U15086 (N_15086,N_14479,N_14709);
and U15087 (N_15087,N_14748,N_14658);
nor U15088 (N_15088,N_14682,N_14720);
nor U15089 (N_15089,N_14676,N_14418);
or U15090 (N_15090,N_14701,N_14757);
and U15091 (N_15091,N_14675,N_14498);
and U15092 (N_15092,N_14462,N_14643);
or U15093 (N_15093,N_14775,N_14405);
and U15094 (N_15094,N_14555,N_14589);
xnor U15095 (N_15095,N_14765,N_14428);
xor U15096 (N_15096,N_14506,N_14591);
and U15097 (N_15097,N_14610,N_14772);
xnor U15098 (N_15098,N_14715,N_14471);
and U15099 (N_15099,N_14564,N_14623);
and U15100 (N_15100,N_14685,N_14729);
or U15101 (N_15101,N_14741,N_14529);
xor U15102 (N_15102,N_14627,N_14496);
nand U15103 (N_15103,N_14537,N_14665);
nor U15104 (N_15104,N_14436,N_14733);
nor U15105 (N_15105,N_14700,N_14695);
xor U15106 (N_15106,N_14708,N_14554);
nor U15107 (N_15107,N_14786,N_14482);
and U15108 (N_15108,N_14608,N_14494);
nand U15109 (N_15109,N_14686,N_14677);
and U15110 (N_15110,N_14558,N_14653);
or U15111 (N_15111,N_14790,N_14647);
or U15112 (N_15112,N_14737,N_14752);
nand U15113 (N_15113,N_14568,N_14680);
nand U15114 (N_15114,N_14784,N_14538);
xnor U15115 (N_15115,N_14777,N_14792);
xnor U15116 (N_15116,N_14434,N_14504);
or U15117 (N_15117,N_14543,N_14621);
or U15118 (N_15118,N_14796,N_14623);
xnor U15119 (N_15119,N_14553,N_14770);
nand U15120 (N_15120,N_14565,N_14775);
and U15121 (N_15121,N_14722,N_14741);
xor U15122 (N_15122,N_14433,N_14547);
xor U15123 (N_15123,N_14700,N_14735);
and U15124 (N_15124,N_14517,N_14792);
xnor U15125 (N_15125,N_14466,N_14726);
or U15126 (N_15126,N_14796,N_14660);
nor U15127 (N_15127,N_14509,N_14764);
or U15128 (N_15128,N_14728,N_14578);
nor U15129 (N_15129,N_14478,N_14778);
or U15130 (N_15130,N_14511,N_14494);
nand U15131 (N_15131,N_14731,N_14636);
xor U15132 (N_15132,N_14542,N_14780);
nand U15133 (N_15133,N_14645,N_14501);
nand U15134 (N_15134,N_14472,N_14429);
or U15135 (N_15135,N_14628,N_14792);
nor U15136 (N_15136,N_14550,N_14472);
nand U15137 (N_15137,N_14749,N_14463);
and U15138 (N_15138,N_14457,N_14671);
nand U15139 (N_15139,N_14540,N_14692);
and U15140 (N_15140,N_14765,N_14724);
nor U15141 (N_15141,N_14639,N_14795);
nand U15142 (N_15142,N_14697,N_14519);
or U15143 (N_15143,N_14539,N_14423);
xor U15144 (N_15144,N_14609,N_14706);
xnor U15145 (N_15145,N_14425,N_14601);
and U15146 (N_15146,N_14498,N_14592);
nor U15147 (N_15147,N_14515,N_14619);
nand U15148 (N_15148,N_14492,N_14525);
or U15149 (N_15149,N_14713,N_14445);
nor U15150 (N_15150,N_14466,N_14720);
and U15151 (N_15151,N_14638,N_14677);
or U15152 (N_15152,N_14531,N_14650);
or U15153 (N_15153,N_14533,N_14502);
and U15154 (N_15154,N_14538,N_14430);
nor U15155 (N_15155,N_14719,N_14530);
and U15156 (N_15156,N_14452,N_14698);
xnor U15157 (N_15157,N_14582,N_14617);
and U15158 (N_15158,N_14716,N_14740);
nor U15159 (N_15159,N_14615,N_14728);
nand U15160 (N_15160,N_14604,N_14479);
nor U15161 (N_15161,N_14611,N_14624);
nand U15162 (N_15162,N_14789,N_14724);
xnor U15163 (N_15163,N_14436,N_14483);
nor U15164 (N_15164,N_14714,N_14570);
and U15165 (N_15165,N_14531,N_14413);
and U15166 (N_15166,N_14700,N_14528);
nor U15167 (N_15167,N_14435,N_14594);
and U15168 (N_15168,N_14682,N_14497);
xnor U15169 (N_15169,N_14607,N_14402);
and U15170 (N_15170,N_14622,N_14592);
xnor U15171 (N_15171,N_14595,N_14664);
nand U15172 (N_15172,N_14653,N_14410);
and U15173 (N_15173,N_14459,N_14695);
or U15174 (N_15174,N_14403,N_14626);
nand U15175 (N_15175,N_14527,N_14493);
nand U15176 (N_15176,N_14542,N_14598);
and U15177 (N_15177,N_14797,N_14508);
or U15178 (N_15178,N_14581,N_14741);
xnor U15179 (N_15179,N_14760,N_14460);
nor U15180 (N_15180,N_14628,N_14656);
xor U15181 (N_15181,N_14623,N_14577);
or U15182 (N_15182,N_14604,N_14472);
nor U15183 (N_15183,N_14723,N_14626);
xor U15184 (N_15184,N_14568,N_14410);
and U15185 (N_15185,N_14562,N_14795);
xnor U15186 (N_15186,N_14565,N_14654);
xor U15187 (N_15187,N_14547,N_14476);
or U15188 (N_15188,N_14646,N_14607);
nand U15189 (N_15189,N_14694,N_14477);
and U15190 (N_15190,N_14737,N_14733);
or U15191 (N_15191,N_14553,N_14547);
nor U15192 (N_15192,N_14455,N_14437);
xnor U15193 (N_15193,N_14694,N_14537);
nand U15194 (N_15194,N_14622,N_14413);
nor U15195 (N_15195,N_14783,N_14710);
xnor U15196 (N_15196,N_14403,N_14522);
nor U15197 (N_15197,N_14791,N_14557);
xnor U15198 (N_15198,N_14435,N_14635);
nor U15199 (N_15199,N_14576,N_14440);
or U15200 (N_15200,N_14879,N_15063);
or U15201 (N_15201,N_14875,N_15136);
and U15202 (N_15202,N_14953,N_14916);
or U15203 (N_15203,N_15186,N_14903);
nor U15204 (N_15204,N_14958,N_14828);
or U15205 (N_15205,N_14939,N_14876);
and U15206 (N_15206,N_14938,N_14891);
nand U15207 (N_15207,N_15088,N_14917);
or U15208 (N_15208,N_14895,N_14956);
nand U15209 (N_15209,N_14952,N_14987);
or U15210 (N_15210,N_14954,N_14848);
nand U15211 (N_15211,N_15005,N_15085);
or U15212 (N_15212,N_14979,N_15108);
nand U15213 (N_15213,N_15070,N_15029);
xor U15214 (N_15214,N_14811,N_14959);
and U15215 (N_15215,N_15189,N_14902);
or U15216 (N_15216,N_15192,N_15170);
and U15217 (N_15217,N_15173,N_15093);
nand U15218 (N_15218,N_15117,N_15091);
nor U15219 (N_15219,N_14912,N_14974);
nor U15220 (N_15220,N_15048,N_15002);
or U15221 (N_15221,N_15025,N_15167);
and U15222 (N_15222,N_15134,N_15000);
nor U15223 (N_15223,N_14896,N_15174);
xnor U15224 (N_15224,N_14823,N_15184);
xor U15225 (N_15225,N_15116,N_14863);
or U15226 (N_15226,N_15020,N_14948);
and U15227 (N_15227,N_15130,N_15194);
nand U15228 (N_15228,N_14936,N_14943);
xor U15229 (N_15229,N_14856,N_15142);
or U15230 (N_15230,N_15015,N_15110);
or U15231 (N_15231,N_15171,N_14844);
xnor U15232 (N_15232,N_14925,N_15149);
and U15233 (N_15233,N_15051,N_14807);
xnor U15234 (N_15234,N_15072,N_14949);
nand U15235 (N_15235,N_14818,N_15111);
or U15236 (N_15236,N_15043,N_15079);
or U15237 (N_15237,N_15125,N_15061);
or U15238 (N_15238,N_15081,N_15157);
nand U15239 (N_15239,N_14822,N_15097);
nand U15240 (N_15240,N_15033,N_15104);
xor U15241 (N_15241,N_14834,N_14950);
xor U15242 (N_15242,N_15042,N_15038);
or U15243 (N_15243,N_15036,N_14942);
xor U15244 (N_15244,N_15121,N_14932);
and U15245 (N_15245,N_15016,N_15133);
nor U15246 (N_15246,N_15181,N_15031);
nor U15247 (N_15247,N_14884,N_14857);
and U15248 (N_15248,N_14841,N_15197);
and U15249 (N_15249,N_14931,N_14820);
or U15250 (N_15250,N_15137,N_15163);
nor U15251 (N_15251,N_14843,N_15135);
nor U15252 (N_15252,N_14914,N_14851);
or U15253 (N_15253,N_14800,N_15014);
xor U15254 (N_15254,N_15023,N_15168);
xor U15255 (N_15255,N_15082,N_14824);
xnor U15256 (N_15256,N_15046,N_15004);
xnor U15257 (N_15257,N_14985,N_15177);
or U15258 (N_15258,N_14835,N_15096);
xor U15259 (N_15259,N_14846,N_14996);
nor U15260 (N_15260,N_14816,N_15119);
nand U15261 (N_15261,N_15069,N_14937);
or U15262 (N_15262,N_15109,N_14927);
nand U15263 (N_15263,N_15018,N_15047);
nand U15264 (N_15264,N_14805,N_14836);
nor U15265 (N_15265,N_14999,N_15010);
nor U15266 (N_15266,N_14920,N_15122);
and U15267 (N_15267,N_15074,N_14963);
and U15268 (N_15268,N_15150,N_15003);
nand U15269 (N_15269,N_15052,N_14968);
xor U15270 (N_15270,N_14802,N_15199);
nand U15271 (N_15271,N_14928,N_14915);
or U15272 (N_15272,N_14840,N_15007);
xnor U15273 (N_15273,N_15021,N_15164);
and U15274 (N_15274,N_15161,N_14878);
and U15275 (N_15275,N_14874,N_14966);
nor U15276 (N_15276,N_14908,N_15187);
xnor U15277 (N_15277,N_15127,N_14830);
nor U15278 (N_15278,N_14892,N_15145);
and U15279 (N_15279,N_14962,N_14918);
xor U15280 (N_15280,N_14988,N_14894);
xnor U15281 (N_15281,N_14880,N_15050);
nor U15282 (N_15282,N_14862,N_14855);
or U15283 (N_15283,N_15141,N_14826);
and U15284 (N_15284,N_14955,N_14870);
nor U15285 (N_15285,N_15151,N_15172);
xnor U15286 (N_15286,N_14814,N_15009);
and U15287 (N_15287,N_15089,N_14827);
or U15288 (N_15288,N_14972,N_14813);
nand U15289 (N_15289,N_14930,N_15165);
and U15290 (N_15290,N_14872,N_14873);
or U15291 (N_15291,N_15044,N_14905);
xor U15292 (N_15292,N_15124,N_14989);
and U15293 (N_15293,N_14832,N_15084);
nand U15294 (N_15294,N_15182,N_14801);
and U15295 (N_15295,N_15075,N_14911);
nand U15296 (N_15296,N_14971,N_14815);
nor U15297 (N_15297,N_15160,N_15066);
or U15298 (N_15298,N_15147,N_15083);
nand U15299 (N_15299,N_15059,N_14960);
or U15300 (N_15300,N_14919,N_15011);
nand U15301 (N_15301,N_15178,N_15101);
or U15302 (N_15302,N_15180,N_14946);
nor U15303 (N_15303,N_14913,N_14833);
xor U15304 (N_15304,N_15162,N_15022);
or U15305 (N_15305,N_14993,N_14897);
nor U15306 (N_15306,N_15118,N_14866);
nor U15307 (N_15307,N_15090,N_15132);
nand U15308 (N_15308,N_14983,N_14804);
nor U15309 (N_15309,N_14926,N_15188);
nand U15310 (N_15310,N_15198,N_14973);
xnor U15311 (N_15311,N_14859,N_15140);
or U15312 (N_15312,N_14951,N_15152);
xor U15313 (N_15313,N_15120,N_14860);
and U15314 (N_15314,N_15053,N_15017);
nand U15315 (N_15315,N_14850,N_14961);
or U15316 (N_15316,N_15062,N_14881);
nand U15317 (N_15317,N_15092,N_14901);
nand U15318 (N_15318,N_15030,N_15064);
nor U15319 (N_15319,N_14981,N_14922);
and U15320 (N_15320,N_15102,N_15103);
nand U15321 (N_15321,N_14899,N_15076);
and U15322 (N_15322,N_14871,N_15153);
or U15323 (N_15323,N_14904,N_14831);
xnor U15324 (N_15324,N_15039,N_15049);
and U15325 (N_15325,N_15148,N_14907);
or U15326 (N_15326,N_14933,N_15144);
nand U15327 (N_15327,N_15129,N_14994);
xor U15328 (N_15328,N_15154,N_14829);
nand U15329 (N_15329,N_15073,N_14887);
or U15330 (N_15330,N_14839,N_14852);
and U15331 (N_15331,N_15146,N_14986);
xnor U15332 (N_15332,N_15094,N_15067);
or U15333 (N_15333,N_14825,N_15185);
xor U15334 (N_15334,N_15113,N_14964);
xnor U15335 (N_15335,N_14944,N_15086);
and U15336 (N_15336,N_15183,N_15099);
nand U15337 (N_15337,N_14947,N_14893);
nor U15338 (N_15338,N_14868,N_15054);
xor U15339 (N_15339,N_14889,N_15155);
nor U15340 (N_15340,N_14842,N_14990);
and U15341 (N_15341,N_14883,N_15106);
xnor U15342 (N_15342,N_15001,N_15095);
nor U15343 (N_15343,N_14869,N_15013);
xor U15344 (N_15344,N_15006,N_14861);
nor U15345 (N_15345,N_15158,N_14934);
or U15346 (N_15346,N_15035,N_14984);
nor U15347 (N_15347,N_14998,N_14819);
nor U15348 (N_15348,N_15191,N_14967);
nand U15349 (N_15349,N_15105,N_15026);
or U15350 (N_15350,N_14864,N_15057);
or U15351 (N_15351,N_15045,N_15128);
nand U15352 (N_15352,N_15179,N_15037);
nor U15353 (N_15353,N_14900,N_14812);
and U15354 (N_15354,N_14877,N_14809);
nand U15355 (N_15355,N_14945,N_15131);
or U15356 (N_15356,N_14975,N_15139);
xor U15357 (N_15357,N_14970,N_15034);
nand U15358 (N_15358,N_15098,N_14882);
nand U15359 (N_15359,N_14997,N_14977);
and U15360 (N_15360,N_14906,N_14806);
or U15361 (N_15361,N_15065,N_15041);
or U15362 (N_15362,N_15087,N_15028);
nand U15363 (N_15363,N_14821,N_15166);
nand U15364 (N_15364,N_14923,N_15169);
nor U15365 (N_15365,N_15156,N_15078);
nand U15366 (N_15366,N_14858,N_15123);
and U15367 (N_15367,N_15107,N_14940);
xnor U15368 (N_15368,N_14898,N_15032);
and U15369 (N_15369,N_15195,N_14909);
nand U15370 (N_15370,N_14865,N_15143);
and U15371 (N_15371,N_15024,N_14888);
xor U15372 (N_15372,N_15126,N_14837);
xor U15373 (N_15373,N_15077,N_15055);
or U15374 (N_15374,N_15019,N_14921);
nand U15375 (N_15375,N_14957,N_14980);
xnor U15376 (N_15376,N_15008,N_15193);
xnor U15377 (N_15377,N_14982,N_15040);
xnor U15378 (N_15378,N_14924,N_15027);
xnor U15379 (N_15379,N_14810,N_14886);
xnor U15380 (N_15380,N_15071,N_15176);
nand U15381 (N_15381,N_14976,N_15080);
nand U15382 (N_15382,N_15115,N_15060);
nand U15383 (N_15383,N_15138,N_15058);
xnor U15384 (N_15384,N_15190,N_14817);
xor U15385 (N_15385,N_14978,N_15056);
nor U15386 (N_15386,N_14992,N_14995);
nand U15387 (N_15387,N_14849,N_14965);
xor U15388 (N_15388,N_14991,N_15012);
and U15389 (N_15389,N_14845,N_15196);
or U15390 (N_15390,N_14969,N_15114);
nor U15391 (N_15391,N_15100,N_14808);
nor U15392 (N_15392,N_15112,N_14853);
and U15393 (N_15393,N_14803,N_14935);
xnor U15394 (N_15394,N_15068,N_14847);
and U15395 (N_15395,N_14941,N_14867);
and U15396 (N_15396,N_14929,N_14838);
or U15397 (N_15397,N_14910,N_14890);
xnor U15398 (N_15398,N_15175,N_14885);
and U15399 (N_15399,N_15159,N_14854);
nor U15400 (N_15400,N_14994,N_15075);
or U15401 (N_15401,N_15072,N_15015);
nor U15402 (N_15402,N_14883,N_14817);
nor U15403 (N_15403,N_15001,N_14847);
nand U15404 (N_15404,N_14897,N_15136);
and U15405 (N_15405,N_15153,N_14993);
nand U15406 (N_15406,N_15125,N_14982);
or U15407 (N_15407,N_15011,N_14980);
or U15408 (N_15408,N_15040,N_14856);
nor U15409 (N_15409,N_15146,N_15168);
or U15410 (N_15410,N_15036,N_14901);
or U15411 (N_15411,N_14855,N_15069);
nand U15412 (N_15412,N_14989,N_14806);
nor U15413 (N_15413,N_14866,N_15083);
xnor U15414 (N_15414,N_14879,N_14977);
xor U15415 (N_15415,N_14978,N_14928);
and U15416 (N_15416,N_14897,N_15074);
nor U15417 (N_15417,N_15017,N_15004);
or U15418 (N_15418,N_14870,N_15146);
and U15419 (N_15419,N_14972,N_14882);
and U15420 (N_15420,N_14986,N_14961);
nand U15421 (N_15421,N_15022,N_14812);
xnor U15422 (N_15422,N_14855,N_15072);
and U15423 (N_15423,N_15157,N_15169);
nor U15424 (N_15424,N_15001,N_15105);
nand U15425 (N_15425,N_15071,N_15138);
xnor U15426 (N_15426,N_15083,N_14820);
xnor U15427 (N_15427,N_15040,N_14936);
nand U15428 (N_15428,N_14830,N_15098);
and U15429 (N_15429,N_14910,N_14834);
or U15430 (N_15430,N_14999,N_14913);
nand U15431 (N_15431,N_14857,N_14916);
nor U15432 (N_15432,N_15154,N_14894);
nand U15433 (N_15433,N_15188,N_14839);
nor U15434 (N_15434,N_14842,N_15120);
or U15435 (N_15435,N_14986,N_14892);
and U15436 (N_15436,N_15159,N_14861);
or U15437 (N_15437,N_15185,N_15049);
and U15438 (N_15438,N_15117,N_14861);
or U15439 (N_15439,N_14840,N_14874);
or U15440 (N_15440,N_14911,N_14971);
or U15441 (N_15441,N_15118,N_15158);
or U15442 (N_15442,N_14871,N_15050);
or U15443 (N_15443,N_14827,N_14824);
nand U15444 (N_15444,N_15115,N_14895);
xnor U15445 (N_15445,N_15198,N_15164);
or U15446 (N_15446,N_15197,N_14969);
xor U15447 (N_15447,N_15122,N_14900);
nand U15448 (N_15448,N_14901,N_15148);
xor U15449 (N_15449,N_15010,N_15073);
nand U15450 (N_15450,N_14927,N_14930);
nor U15451 (N_15451,N_14865,N_15006);
nand U15452 (N_15452,N_15147,N_15054);
or U15453 (N_15453,N_15090,N_15188);
or U15454 (N_15454,N_15051,N_14933);
nand U15455 (N_15455,N_14858,N_14857);
and U15456 (N_15456,N_15075,N_14821);
and U15457 (N_15457,N_15002,N_15189);
xor U15458 (N_15458,N_15018,N_14831);
nand U15459 (N_15459,N_15059,N_15134);
xnor U15460 (N_15460,N_14881,N_14872);
nor U15461 (N_15461,N_15108,N_15064);
xnor U15462 (N_15462,N_15004,N_14827);
nand U15463 (N_15463,N_15156,N_15150);
nand U15464 (N_15464,N_14877,N_14989);
nor U15465 (N_15465,N_14946,N_14919);
nand U15466 (N_15466,N_15069,N_15052);
nand U15467 (N_15467,N_14947,N_15061);
or U15468 (N_15468,N_15104,N_14905);
nand U15469 (N_15469,N_14923,N_14980);
nor U15470 (N_15470,N_14908,N_14895);
and U15471 (N_15471,N_15134,N_14835);
nand U15472 (N_15472,N_15103,N_15001);
xor U15473 (N_15473,N_14808,N_15066);
nand U15474 (N_15474,N_15013,N_15067);
nor U15475 (N_15475,N_14920,N_14931);
nand U15476 (N_15476,N_14819,N_14989);
nand U15477 (N_15477,N_14893,N_15140);
nor U15478 (N_15478,N_14935,N_15165);
nor U15479 (N_15479,N_15095,N_15062);
and U15480 (N_15480,N_15116,N_15160);
and U15481 (N_15481,N_14843,N_14991);
nand U15482 (N_15482,N_14918,N_14957);
and U15483 (N_15483,N_15136,N_15154);
xor U15484 (N_15484,N_14903,N_14989);
or U15485 (N_15485,N_14970,N_14863);
or U15486 (N_15486,N_14816,N_14953);
nand U15487 (N_15487,N_15081,N_14875);
xor U15488 (N_15488,N_14996,N_14954);
nor U15489 (N_15489,N_15071,N_14988);
xnor U15490 (N_15490,N_14907,N_14851);
nand U15491 (N_15491,N_14980,N_14907);
nor U15492 (N_15492,N_14902,N_15122);
nand U15493 (N_15493,N_15031,N_14873);
nor U15494 (N_15494,N_15015,N_15024);
nor U15495 (N_15495,N_15145,N_14917);
or U15496 (N_15496,N_15168,N_14880);
and U15497 (N_15497,N_15166,N_15162);
or U15498 (N_15498,N_15023,N_15004);
xor U15499 (N_15499,N_14878,N_14818);
and U15500 (N_15500,N_15124,N_14974);
or U15501 (N_15501,N_15195,N_15019);
nand U15502 (N_15502,N_14909,N_15197);
or U15503 (N_15503,N_14975,N_15053);
nand U15504 (N_15504,N_14994,N_15068);
nand U15505 (N_15505,N_15064,N_15014);
and U15506 (N_15506,N_14874,N_14898);
nand U15507 (N_15507,N_15144,N_15036);
xnor U15508 (N_15508,N_14930,N_15150);
or U15509 (N_15509,N_14879,N_15080);
nor U15510 (N_15510,N_15188,N_14827);
and U15511 (N_15511,N_15066,N_15033);
nor U15512 (N_15512,N_15082,N_14807);
xor U15513 (N_15513,N_14917,N_15052);
or U15514 (N_15514,N_14811,N_15184);
xnor U15515 (N_15515,N_14823,N_15150);
nor U15516 (N_15516,N_14939,N_15092);
nor U15517 (N_15517,N_15087,N_14999);
nor U15518 (N_15518,N_15011,N_15178);
or U15519 (N_15519,N_14802,N_14898);
nor U15520 (N_15520,N_15086,N_15167);
and U15521 (N_15521,N_14875,N_15034);
and U15522 (N_15522,N_15138,N_14823);
xnor U15523 (N_15523,N_14937,N_14995);
and U15524 (N_15524,N_15066,N_15088);
nor U15525 (N_15525,N_15141,N_15125);
or U15526 (N_15526,N_14900,N_14971);
or U15527 (N_15527,N_14843,N_14950);
or U15528 (N_15528,N_15025,N_14959);
xnor U15529 (N_15529,N_14959,N_14885);
nor U15530 (N_15530,N_15150,N_15106);
or U15531 (N_15531,N_14893,N_15016);
xor U15532 (N_15532,N_15014,N_15195);
or U15533 (N_15533,N_15081,N_14984);
nand U15534 (N_15534,N_14888,N_14809);
nand U15535 (N_15535,N_14928,N_14993);
nor U15536 (N_15536,N_14991,N_14979);
nand U15537 (N_15537,N_14815,N_14999);
nor U15538 (N_15538,N_14935,N_14843);
and U15539 (N_15539,N_15009,N_15062);
nor U15540 (N_15540,N_14860,N_15008);
nand U15541 (N_15541,N_15053,N_14883);
xnor U15542 (N_15542,N_14927,N_15149);
nor U15543 (N_15543,N_15118,N_14967);
xor U15544 (N_15544,N_14902,N_15133);
nor U15545 (N_15545,N_14954,N_15096);
xor U15546 (N_15546,N_14890,N_15004);
nor U15547 (N_15547,N_15039,N_15155);
xnor U15548 (N_15548,N_14926,N_14844);
nor U15549 (N_15549,N_14970,N_14809);
nor U15550 (N_15550,N_14882,N_14860);
xor U15551 (N_15551,N_15080,N_14842);
and U15552 (N_15552,N_14927,N_15173);
xor U15553 (N_15553,N_15143,N_14880);
nand U15554 (N_15554,N_15160,N_15159);
nor U15555 (N_15555,N_15169,N_15134);
xor U15556 (N_15556,N_15152,N_14960);
and U15557 (N_15557,N_15179,N_15191);
xor U15558 (N_15558,N_14855,N_15004);
and U15559 (N_15559,N_15079,N_15134);
nand U15560 (N_15560,N_15114,N_15117);
nor U15561 (N_15561,N_14978,N_14992);
xnor U15562 (N_15562,N_14970,N_14922);
nor U15563 (N_15563,N_15043,N_14924);
and U15564 (N_15564,N_14858,N_14807);
or U15565 (N_15565,N_15030,N_15096);
nand U15566 (N_15566,N_15085,N_14979);
or U15567 (N_15567,N_15076,N_15199);
or U15568 (N_15568,N_14932,N_14987);
xor U15569 (N_15569,N_15087,N_15148);
nor U15570 (N_15570,N_14833,N_15033);
or U15571 (N_15571,N_14952,N_15149);
and U15572 (N_15572,N_14838,N_14970);
or U15573 (N_15573,N_15143,N_14891);
and U15574 (N_15574,N_15014,N_14864);
nand U15575 (N_15575,N_15051,N_15118);
nand U15576 (N_15576,N_14817,N_14864);
nand U15577 (N_15577,N_14865,N_14907);
and U15578 (N_15578,N_15007,N_14918);
xnor U15579 (N_15579,N_15066,N_15154);
or U15580 (N_15580,N_15012,N_15060);
and U15581 (N_15581,N_15077,N_15022);
xor U15582 (N_15582,N_14987,N_14827);
and U15583 (N_15583,N_15115,N_15087);
nor U15584 (N_15584,N_14818,N_15189);
and U15585 (N_15585,N_15014,N_14956);
or U15586 (N_15586,N_14938,N_14889);
nand U15587 (N_15587,N_14996,N_14955);
or U15588 (N_15588,N_15075,N_15172);
and U15589 (N_15589,N_15113,N_15197);
xnor U15590 (N_15590,N_14964,N_15152);
xnor U15591 (N_15591,N_14805,N_15084);
nor U15592 (N_15592,N_15001,N_14997);
or U15593 (N_15593,N_15033,N_15180);
or U15594 (N_15594,N_15114,N_14974);
or U15595 (N_15595,N_15101,N_15112);
nor U15596 (N_15596,N_14820,N_14840);
nor U15597 (N_15597,N_14867,N_15008);
nand U15598 (N_15598,N_14991,N_14990);
or U15599 (N_15599,N_15168,N_14854);
or U15600 (N_15600,N_15419,N_15581);
and U15601 (N_15601,N_15381,N_15449);
nand U15602 (N_15602,N_15479,N_15594);
and U15603 (N_15603,N_15266,N_15388);
nor U15604 (N_15604,N_15369,N_15210);
xnor U15605 (N_15605,N_15481,N_15284);
xor U15606 (N_15606,N_15500,N_15376);
or U15607 (N_15607,N_15397,N_15432);
and U15608 (N_15608,N_15561,N_15239);
or U15609 (N_15609,N_15330,N_15331);
nand U15610 (N_15610,N_15454,N_15480);
nor U15611 (N_15611,N_15549,N_15336);
nor U15612 (N_15612,N_15577,N_15238);
or U15613 (N_15613,N_15486,N_15421);
nand U15614 (N_15614,N_15447,N_15555);
nand U15615 (N_15615,N_15539,N_15362);
nand U15616 (N_15616,N_15476,N_15366);
xnor U15617 (N_15617,N_15262,N_15599);
nor U15618 (N_15618,N_15280,N_15588);
or U15619 (N_15619,N_15450,N_15269);
xnor U15620 (N_15620,N_15296,N_15367);
and U15621 (N_15621,N_15440,N_15251);
nor U15622 (N_15622,N_15274,N_15541);
nor U15623 (N_15623,N_15385,N_15329);
nand U15624 (N_15624,N_15278,N_15482);
xnor U15625 (N_15625,N_15435,N_15204);
nor U15626 (N_15626,N_15523,N_15484);
nor U15627 (N_15627,N_15254,N_15398);
and U15628 (N_15628,N_15498,N_15218);
nand U15629 (N_15629,N_15308,N_15404);
and U15630 (N_15630,N_15227,N_15585);
nor U15631 (N_15631,N_15597,N_15221);
nor U15632 (N_15632,N_15340,N_15572);
nand U15633 (N_15633,N_15231,N_15578);
nor U15634 (N_15634,N_15573,N_15433);
xor U15635 (N_15635,N_15423,N_15326);
and U15636 (N_15636,N_15426,N_15311);
or U15637 (N_15637,N_15220,N_15203);
nor U15638 (N_15638,N_15408,N_15503);
xor U15639 (N_15639,N_15424,N_15299);
xnor U15640 (N_15640,N_15209,N_15265);
nand U15641 (N_15641,N_15552,N_15233);
nand U15642 (N_15642,N_15249,N_15228);
nand U15643 (N_15643,N_15442,N_15505);
nand U15644 (N_15644,N_15410,N_15212);
xnor U15645 (N_15645,N_15456,N_15402);
nor U15646 (N_15646,N_15320,N_15226);
and U15647 (N_15647,N_15592,N_15566);
and U15648 (N_15648,N_15443,N_15322);
and U15649 (N_15649,N_15507,N_15593);
or U15650 (N_15650,N_15264,N_15201);
and U15651 (N_15651,N_15488,N_15524);
xor U15652 (N_15652,N_15506,N_15595);
and U15653 (N_15653,N_15387,N_15407);
or U15654 (N_15654,N_15455,N_15237);
nor U15655 (N_15655,N_15353,N_15205);
or U15656 (N_15656,N_15272,N_15465);
nor U15657 (N_15657,N_15316,N_15533);
and U15658 (N_15658,N_15391,N_15222);
nor U15659 (N_15659,N_15317,N_15370);
nand U15660 (N_15660,N_15401,N_15574);
nand U15661 (N_15661,N_15590,N_15303);
and U15662 (N_15662,N_15444,N_15553);
nor U15663 (N_15663,N_15396,N_15342);
nor U15664 (N_15664,N_15289,N_15543);
xnor U15665 (N_15665,N_15348,N_15261);
or U15666 (N_15666,N_15546,N_15495);
or U15667 (N_15667,N_15365,N_15493);
nor U15668 (N_15668,N_15291,N_15386);
nand U15669 (N_15669,N_15300,N_15314);
or U15670 (N_15670,N_15310,N_15516);
nand U15671 (N_15671,N_15530,N_15525);
or U15672 (N_15672,N_15409,N_15207);
nor U15673 (N_15673,N_15313,N_15466);
nand U15674 (N_15674,N_15596,N_15544);
and U15675 (N_15675,N_15517,N_15428);
nand U15676 (N_15676,N_15413,N_15492);
xnor U15677 (N_15677,N_15259,N_15319);
or U15678 (N_15678,N_15451,N_15246);
or U15679 (N_15679,N_15478,N_15436);
nand U15680 (N_15680,N_15315,N_15430);
nor U15681 (N_15681,N_15587,N_15349);
nor U15682 (N_15682,N_15267,N_15345);
xnor U15683 (N_15683,N_15297,N_15235);
and U15684 (N_15684,N_15528,N_15459);
and U15685 (N_15685,N_15475,N_15258);
or U15686 (N_15686,N_15429,N_15302);
nand U15687 (N_15687,N_15354,N_15277);
and U15688 (N_15688,N_15522,N_15242);
nor U15689 (N_15689,N_15583,N_15580);
xor U15690 (N_15690,N_15540,N_15598);
xor U15691 (N_15691,N_15335,N_15438);
or U15692 (N_15692,N_15548,N_15591);
nor U15693 (N_15693,N_15374,N_15257);
nor U15694 (N_15694,N_15281,N_15304);
xnor U15695 (N_15695,N_15357,N_15361);
or U15696 (N_15696,N_15562,N_15453);
and U15697 (N_15697,N_15293,N_15208);
nor U15698 (N_15698,N_15542,N_15567);
or U15699 (N_15699,N_15589,N_15384);
nor U15700 (N_15700,N_15462,N_15347);
nor U15701 (N_15701,N_15383,N_15582);
xor U15702 (N_15702,N_15375,N_15415);
or U15703 (N_15703,N_15346,N_15224);
or U15704 (N_15704,N_15570,N_15371);
nand U15705 (N_15705,N_15301,N_15399);
and U15706 (N_15706,N_15485,N_15448);
nand U15707 (N_15707,N_15324,N_15467);
nand U15708 (N_15708,N_15473,N_15260);
or U15709 (N_15709,N_15321,N_15216);
or U15710 (N_15710,N_15325,N_15200);
nand U15711 (N_15711,N_15377,N_15518);
xor U15712 (N_15712,N_15241,N_15282);
nand U15713 (N_15713,N_15513,N_15286);
xor U15714 (N_15714,N_15306,N_15470);
xnor U15715 (N_15715,N_15350,N_15547);
nand U15716 (N_15716,N_15206,N_15287);
nand U15717 (N_15717,N_15416,N_15468);
or U15718 (N_15718,N_15332,N_15236);
and U15719 (N_15719,N_15271,N_15240);
xnor U15720 (N_15720,N_15352,N_15294);
xnor U15721 (N_15721,N_15250,N_15554);
nand U15722 (N_15722,N_15417,N_15248);
nor U15723 (N_15723,N_15344,N_15538);
nand U15724 (N_15724,N_15234,N_15245);
and U15725 (N_15725,N_15531,N_15521);
nor U15726 (N_15726,N_15328,N_15584);
nand U15727 (N_15727,N_15576,N_15558);
or U15728 (N_15728,N_15202,N_15537);
nor U15729 (N_15729,N_15276,N_15529);
xnor U15730 (N_15730,N_15483,N_15508);
nor U15731 (N_15731,N_15490,N_15363);
and U15732 (N_15732,N_15406,N_15255);
nor U15733 (N_15733,N_15288,N_15312);
xor U15734 (N_15734,N_15405,N_15565);
or U15735 (N_15735,N_15372,N_15489);
and U15736 (N_15736,N_15268,N_15568);
and U15737 (N_15737,N_15411,N_15559);
nand U15738 (N_15738,N_15232,N_15252);
nor U15739 (N_15739,N_15263,N_15339);
nor U15740 (N_15740,N_15532,N_15472);
nor U15741 (N_15741,N_15338,N_15351);
and U15742 (N_15742,N_15400,N_15535);
nand U15743 (N_15743,N_15256,N_15422);
or U15744 (N_15744,N_15536,N_15461);
and U15745 (N_15745,N_15403,N_15318);
nand U15746 (N_15746,N_15334,N_15355);
or U15747 (N_15747,N_15586,N_15360);
and U15748 (N_15748,N_15557,N_15364);
nor U15749 (N_15749,N_15477,N_15215);
nand U15750 (N_15750,N_15273,N_15244);
nand U15751 (N_15751,N_15393,N_15295);
nor U15752 (N_15752,N_15247,N_15458);
xnor U15753 (N_15753,N_15379,N_15520);
and U15754 (N_15754,N_15457,N_15464);
nand U15755 (N_15755,N_15526,N_15283);
and U15756 (N_15756,N_15211,N_15327);
nand U15757 (N_15757,N_15392,N_15560);
nor U15758 (N_15758,N_15441,N_15307);
nand U15759 (N_15759,N_15358,N_15510);
and U15760 (N_15760,N_15298,N_15501);
nand U15761 (N_15761,N_15515,N_15309);
xnor U15762 (N_15762,N_15551,N_15445);
and U15763 (N_15763,N_15446,N_15545);
xor U15764 (N_15764,N_15214,N_15434);
nor U15765 (N_15765,N_15343,N_15534);
nor U15766 (N_15766,N_15356,N_15499);
xnor U15767 (N_15767,N_15509,N_15270);
nand U15768 (N_15768,N_15527,N_15217);
nor U15769 (N_15769,N_15563,N_15556);
nor U15770 (N_15770,N_15579,N_15460);
and U15771 (N_15771,N_15285,N_15219);
nor U15772 (N_15772,N_15223,N_15229);
xnor U15773 (N_15773,N_15230,N_15380);
nor U15774 (N_15774,N_15418,N_15569);
and U15775 (N_15775,N_15390,N_15564);
and U15776 (N_15776,N_15511,N_15279);
xnor U15777 (N_15777,N_15469,N_15494);
nor U15778 (N_15778,N_15333,N_15292);
and U15779 (N_15779,N_15502,N_15382);
xnor U15780 (N_15780,N_15425,N_15323);
and U15781 (N_15781,N_15497,N_15504);
nand U15782 (N_15782,N_15427,N_15378);
nand U15783 (N_15783,N_15253,N_15550);
xnor U15784 (N_15784,N_15431,N_15341);
xor U15785 (N_15785,N_15225,N_15496);
nand U15786 (N_15786,N_15373,N_15437);
nand U15787 (N_15787,N_15337,N_15487);
or U15788 (N_15788,N_15414,N_15395);
nor U15789 (N_15789,N_15359,N_15512);
nand U15790 (N_15790,N_15305,N_15463);
or U15791 (N_15791,N_15575,N_15394);
xnor U15792 (N_15792,N_15420,N_15519);
or U15793 (N_15793,N_15290,N_15474);
and U15794 (N_15794,N_15471,N_15571);
nor U15795 (N_15795,N_15213,N_15243);
or U15796 (N_15796,N_15275,N_15514);
nand U15797 (N_15797,N_15491,N_15412);
nor U15798 (N_15798,N_15452,N_15389);
nand U15799 (N_15799,N_15368,N_15439);
xor U15800 (N_15800,N_15537,N_15225);
and U15801 (N_15801,N_15278,N_15569);
nor U15802 (N_15802,N_15402,N_15266);
nor U15803 (N_15803,N_15530,N_15550);
nand U15804 (N_15804,N_15352,N_15298);
and U15805 (N_15805,N_15557,N_15399);
or U15806 (N_15806,N_15206,N_15379);
nor U15807 (N_15807,N_15467,N_15390);
nand U15808 (N_15808,N_15555,N_15573);
nand U15809 (N_15809,N_15314,N_15432);
and U15810 (N_15810,N_15201,N_15337);
or U15811 (N_15811,N_15446,N_15201);
nand U15812 (N_15812,N_15446,N_15458);
nor U15813 (N_15813,N_15526,N_15224);
nand U15814 (N_15814,N_15218,N_15255);
and U15815 (N_15815,N_15255,N_15387);
nand U15816 (N_15816,N_15410,N_15508);
nor U15817 (N_15817,N_15559,N_15520);
and U15818 (N_15818,N_15257,N_15389);
nand U15819 (N_15819,N_15401,N_15446);
nand U15820 (N_15820,N_15493,N_15341);
xor U15821 (N_15821,N_15362,N_15379);
xor U15822 (N_15822,N_15348,N_15502);
and U15823 (N_15823,N_15438,N_15221);
nor U15824 (N_15824,N_15494,N_15247);
xnor U15825 (N_15825,N_15411,N_15234);
and U15826 (N_15826,N_15269,N_15434);
or U15827 (N_15827,N_15410,N_15431);
and U15828 (N_15828,N_15427,N_15353);
nand U15829 (N_15829,N_15248,N_15261);
nor U15830 (N_15830,N_15279,N_15212);
xor U15831 (N_15831,N_15379,N_15270);
and U15832 (N_15832,N_15396,N_15597);
and U15833 (N_15833,N_15510,N_15433);
nor U15834 (N_15834,N_15552,N_15526);
xnor U15835 (N_15835,N_15543,N_15363);
xor U15836 (N_15836,N_15369,N_15571);
and U15837 (N_15837,N_15456,N_15496);
nand U15838 (N_15838,N_15383,N_15423);
xor U15839 (N_15839,N_15442,N_15264);
nor U15840 (N_15840,N_15504,N_15433);
nor U15841 (N_15841,N_15491,N_15207);
or U15842 (N_15842,N_15578,N_15317);
xnor U15843 (N_15843,N_15510,N_15455);
or U15844 (N_15844,N_15487,N_15365);
xor U15845 (N_15845,N_15464,N_15367);
xor U15846 (N_15846,N_15324,N_15282);
and U15847 (N_15847,N_15218,N_15322);
and U15848 (N_15848,N_15381,N_15535);
xor U15849 (N_15849,N_15260,N_15431);
nand U15850 (N_15850,N_15522,N_15438);
or U15851 (N_15851,N_15340,N_15430);
xnor U15852 (N_15852,N_15329,N_15515);
or U15853 (N_15853,N_15491,N_15326);
or U15854 (N_15854,N_15303,N_15486);
xor U15855 (N_15855,N_15315,N_15551);
and U15856 (N_15856,N_15568,N_15359);
or U15857 (N_15857,N_15434,N_15455);
or U15858 (N_15858,N_15280,N_15591);
or U15859 (N_15859,N_15416,N_15263);
xor U15860 (N_15860,N_15363,N_15564);
and U15861 (N_15861,N_15238,N_15502);
and U15862 (N_15862,N_15281,N_15421);
or U15863 (N_15863,N_15504,N_15444);
nand U15864 (N_15864,N_15518,N_15297);
nand U15865 (N_15865,N_15271,N_15263);
xnor U15866 (N_15866,N_15384,N_15437);
xnor U15867 (N_15867,N_15302,N_15441);
xnor U15868 (N_15868,N_15354,N_15387);
xnor U15869 (N_15869,N_15346,N_15506);
or U15870 (N_15870,N_15261,N_15302);
xnor U15871 (N_15871,N_15350,N_15422);
xor U15872 (N_15872,N_15454,N_15439);
nand U15873 (N_15873,N_15331,N_15215);
nor U15874 (N_15874,N_15471,N_15225);
nor U15875 (N_15875,N_15415,N_15221);
and U15876 (N_15876,N_15557,N_15529);
or U15877 (N_15877,N_15383,N_15385);
nand U15878 (N_15878,N_15224,N_15587);
nor U15879 (N_15879,N_15557,N_15501);
nand U15880 (N_15880,N_15406,N_15240);
nand U15881 (N_15881,N_15266,N_15365);
nor U15882 (N_15882,N_15390,N_15418);
or U15883 (N_15883,N_15278,N_15455);
nand U15884 (N_15884,N_15292,N_15504);
xor U15885 (N_15885,N_15377,N_15416);
and U15886 (N_15886,N_15234,N_15509);
nand U15887 (N_15887,N_15272,N_15350);
nor U15888 (N_15888,N_15461,N_15275);
xor U15889 (N_15889,N_15487,N_15374);
nor U15890 (N_15890,N_15531,N_15564);
or U15891 (N_15891,N_15377,N_15470);
xnor U15892 (N_15892,N_15539,N_15356);
and U15893 (N_15893,N_15510,N_15380);
nand U15894 (N_15894,N_15395,N_15314);
and U15895 (N_15895,N_15235,N_15399);
and U15896 (N_15896,N_15282,N_15574);
nand U15897 (N_15897,N_15401,N_15432);
or U15898 (N_15898,N_15297,N_15452);
nand U15899 (N_15899,N_15217,N_15380);
and U15900 (N_15900,N_15353,N_15227);
xnor U15901 (N_15901,N_15250,N_15462);
xor U15902 (N_15902,N_15524,N_15451);
and U15903 (N_15903,N_15445,N_15273);
nor U15904 (N_15904,N_15219,N_15306);
xnor U15905 (N_15905,N_15466,N_15484);
and U15906 (N_15906,N_15405,N_15506);
nand U15907 (N_15907,N_15367,N_15345);
or U15908 (N_15908,N_15279,N_15327);
nand U15909 (N_15909,N_15506,N_15204);
xnor U15910 (N_15910,N_15498,N_15486);
nand U15911 (N_15911,N_15263,N_15559);
and U15912 (N_15912,N_15448,N_15345);
nor U15913 (N_15913,N_15323,N_15580);
xor U15914 (N_15914,N_15534,N_15402);
and U15915 (N_15915,N_15353,N_15477);
and U15916 (N_15916,N_15410,N_15363);
nand U15917 (N_15917,N_15528,N_15399);
or U15918 (N_15918,N_15368,N_15324);
nor U15919 (N_15919,N_15576,N_15301);
and U15920 (N_15920,N_15484,N_15361);
and U15921 (N_15921,N_15267,N_15355);
or U15922 (N_15922,N_15325,N_15208);
nor U15923 (N_15923,N_15286,N_15524);
and U15924 (N_15924,N_15268,N_15559);
and U15925 (N_15925,N_15345,N_15583);
nand U15926 (N_15926,N_15375,N_15287);
xor U15927 (N_15927,N_15235,N_15238);
and U15928 (N_15928,N_15582,N_15215);
and U15929 (N_15929,N_15489,N_15253);
nor U15930 (N_15930,N_15574,N_15455);
nor U15931 (N_15931,N_15492,N_15582);
and U15932 (N_15932,N_15346,N_15232);
and U15933 (N_15933,N_15269,N_15301);
xnor U15934 (N_15934,N_15244,N_15275);
and U15935 (N_15935,N_15289,N_15253);
and U15936 (N_15936,N_15514,N_15507);
and U15937 (N_15937,N_15389,N_15260);
and U15938 (N_15938,N_15325,N_15426);
nand U15939 (N_15939,N_15399,N_15262);
xnor U15940 (N_15940,N_15380,N_15581);
or U15941 (N_15941,N_15234,N_15416);
xnor U15942 (N_15942,N_15487,N_15251);
and U15943 (N_15943,N_15504,N_15290);
nor U15944 (N_15944,N_15339,N_15318);
or U15945 (N_15945,N_15449,N_15424);
or U15946 (N_15946,N_15531,N_15444);
nor U15947 (N_15947,N_15292,N_15318);
or U15948 (N_15948,N_15247,N_15564);
nand U15949 (N_15949,N_15250,N_15422);
nor U15950 (N_15950,N_15543,N_15455);
nor U15951 (N_15951,N_15334,N_15599);
or U15952 (N_15952,N_15436,N_15253);
nor U15953 (N_15953,N_15467,N_15512);
and U15954 (N_15954,N_15420,N_15329);
or U15955 (N_15955,N_15295,N_15549);
xor U15956 (N_15956,N_15312,N_15239);
xnor U15957 (N_15957,N_15379,N_15352);
or U15958 (N_15958,N_15337,N_15491);
nand U15959 (N_15959,N_15434,N_15208);
xor U15960 (N_15960,N_15294,N_15271);
xnor U15961 (N_15961,N_15542,N_15248);
nand U15962 (N_15962,N_15581,N_15552);
nor U15963 (N_15963,N_15321,N_15560);
nor U15964 (N_15964,N_15450,N_15476);
xor U15965 (N_15965,N_15584,N_15491);
nand U15966 (N_15966,N_15409,N_15258);
and U15967 (N_15967,N_15549,N_15440);
or U15968 (N_15968,N_15353,N_15362);
nand U15969 (N_15969,N_15331,N_15213);
xnor U15970 (N_15970,N_15462,N_15217);
or U15971 (N_15971,N_15313,N_15423);
or U15972 (N_15972,N_15591,N_15488);
nand U15973 (N_15973,N_15368,N_15364);
nand U15974 (N_15974,N_15420,N_15379);
nor U15975 (N_15975,N_15247,N_15351);
and U15976 (N_15976,N_15430,N_15257);
nor U15977 (N_15977,N_15497,N_15511);
and U15978 (N_15978,N_15472,N_15246);
xnor U15979 (N_15979,N_15247,N_15525);
nor U15980 (N_15980,N_15263,N_15497);
nor U15981 (N_15981,N_15280,N_15366);
nand U15982 (N_15982,N_15353,N_15471);
nand U15983 (N_15983,N_15338,N_15260);
and U15984 (N_15984,N_15597,N_15595);
and U15985 (N_15985,N_15270,N_15245);
xnor U15986 (N_15986,N_15323,N_15297);
nand U15987 (N_15987,N_15316,N_15463);
nor U15988 (N_15988,N_15234,N_15253);
nor U15989 (N_15989,N_15426,N_15269);
and U15990 (N_15990,N_15278,N_15380);
nor U15991 (N_15991,N_15410,N_15451);
xor U15992 (N_15992,N_15273,N_15543);
xnor U15993 (N_15993,N_15433,N_15265);
or U15994 (N_15994,N_15204,N_15422);
xnor U15995 (N_15995,N_15290,N_15438);
nor U15996 (N_15996,N_15490,N_15544);
nor U15997 (N_15997,N_15443,N_15522);
nor U15998 (N_15998,N_15406,N_15446);
nor U15999 (N_15999,N_15292,N_15519);
xnor U16000 (N_16000,N_15996,N_15991);
or U16001 (N_16001,N_15754,N_15611);
and U16002 (N_16002,N_15682,N_15861);
nand U16003 (N_16003,N_15707,N_15778);
or U16004 (N_16004,N_15748,N_15776);
nand U16005 (N_16005,N_15954,N_15795);
or U16006 (N_16006,N_15768,N_15946);
and U16007 (N_16007,N_15989,N_15923);
and U16008 (N_16008,N_15812,N_15747);
and U16009 (N_16009,N_15877,N_15709);
nand U16010 (N_16010,N_15876,N_15711);
xnor U16011 (N_16011,N_15679,N_15832);
and U16012 (N_16012,N_15891,N_15645);
xor U16013 (N_16013,N_15608,N_15921);
nor U16014 (N_16014,N_15853,N_15668);
nand U16015 (N_16015,N_15820,N_15654);
xnor U16016 (N_16016,N_15888,N_15883);
nand U16017 (N_16017,N_15676,N_15749);
and U16018 (N_16018,N_15600,N_15935);
nand U16019 (N_16019,N_15648,N_15857);
nand U16020 (N_16020,N_15823,N_15916);
nor U16021 (N_16021,N_15848,N_15933);
nand U16022 (N_16022,N_15995,N_15941);
and U16023 (N_16023,N_15724,N_15693);
nor U16024 (N_16024,N_15801,N_15886);
xnor U16025 (N_16025,N_15810,N_15722);
nand U16026 (N_16026,N_15755,N_15854);
and U16027 (N_16027,N_15792,N_15997);
nor U16028 (N_16028,N_15647,N_15992);
nor U16029 (N_16029,N_15818,N_15742);
and U16030 (N_16030,N_15962,N_15631);
nand U16031 (N_16031,N_15761,N_15976);
or U16032 (N_16032,N_15890,N_15908);
xor U16033 (N_16033,N_15858,N_15912);
nor U16034 (N_16034,N_15753,N_15730);
and U16035 (N_16035,N_15943,N_15957);
nand U16036 (N_16036,N_15688,N_15610);
nor U16037 (N_16037,N_15799,N_15987);
and U16038 (N_16038,N_15703,N_15607);
or U16039 (N_16039,N_15892,N_15663);
xor U16040 (N_16040,N_15691,N_15867);
and U16041 (N_16041,N_15814,N_15665);
nand U16042 (N_16042,N_15796,N_15712);
nand U16043 (N_16043,N_15845,N_15869);
and U16044 (N_16044,N_15966,N_15612);
nor U16045 (N_16045,N_15728,N_15826);
xnor U16046 (N_16046,N_15739,N_15819);
nor U16047 (N_16047,N_15609,N_15903);
nand U16048 (N_16048,N_15838,N_15856);
or U16049 (N_16049,N_15725,N_15917);
xnor U16050 (N_16050,N_15939,N_15690);
xnor U16051 (N_16051,N_15620,N_15827);
or U16052 (N_16052,N_15901,N_15956);
or U16053 (N_16053,N_15919,N_15833);
xor U16054 (N_16054,N_15781,N_15863);
and U16055 (N_16055,N_15619,N_15729);
nor U16056 (N_16056,N_15675,N_15930);
and U16057 (N_16057,N_15671,N_15815);
and U16058 (N_16058,N_15999,N_15623);
nor U16059 (N_16059,N_15803,N_15870);
nand U16060 (N_16060,N_15667,N_15813);
and U16061 (N_16061,N_15882,N_15686);
or U16062 (N_16062,N_15752,N_15840);
and U16063 (N_16063,N_15643,N_15660);
nand U16064 (N_16064,N_15843,N_15622);
or U16065 (N_16065,N_15640,N_15750);
or U16066 (N_16066,N_15603,N_15646);
and U16067 (N_16067,N_15906,N_15634);
and U16068 (N_16068,N_15910,N_15851);
nor U16069 (N_16069,N_15740,N_15914);
and U16070 (N_16070,N_15756,N_15894);
or U16071 (N_16071,N_15928,N_15658);
or U16072 (N_16072,N_15684,N_15633);
and U16073 (N_16073,N_15791,N_15873);
xor U16074 (N_16074,N_15696,N_15708);
nand U16075 (N_16075,N_15889,N_15683);
nor U16076 (N_16076,N_15677,N_15859);
or U16077 (N_16077,N_15950,N_15953);
nand U16078 (N_16078,N_15785,N_15661);
or U16079 (N_16079,N_15850,N_15885);
nand U16080 (N_16080,N_15984,N_15936);
and U16081 (N_16081,N_15628,N_15769);
nor U16082 (N_16082,N_15767,N_15630);
nor U16083 (N_16083,N_15907,N_15716);
nand U16084 (N_16084,N_15672,N_15925);
nand U16085 (N_16085,N_15790,N_15652);
nor U16086 (N_16086,N_15804,N_15821);
xor U16087 (N_16087,N_15932,N_15627);
or U16088 (N_16088,N_15875,N_15723);
nor U16089 (N_16089,N_15940,N_15704);
or U16090 (N_16090,N_15763,N_15642);
xor U16091 (N_16091,N_15687,N_15692);
nand U16092 (N_16092,N_15839,N_15699);
or U16093 (N_16093,N_15605,N_15681);
nand U16094 (N_16094,N_15905,N_15805);
xor U16095 (N_16095,N_15915,N_15811);
nand U16096 (N_16096,N_15817,N_15837);
and U16097 (N_16097,N_15972,N_15779);
or U16098 (N_16098,N_15942,N_15702);
or U16099 (N_16099,N_15897,N_15899);
nand U16100 (N_16100,N_15759,N_15980);
and U16101 (N_16101,N_15637,N_15829);
xor U16102 (N_16102,N_15705,N_15762);
xnor U16103 (N_16103,N_15736,N_15746);
or U16104 (N_16104,N_15664,N_15793);
and U16105 (N_16105,N_15738,N_15893);
nor U16106 (N_16106,N_15629,N_15715);
and U16107 (N_16107,N_15973,N_15994);
nand U16108 (N_16108,N_15808,N_15741);
or U16109 (N_16109,N_15884,N_15695);
or U16110 (N_16110,N_15971,N_15697);
nor U16111 (N_16111,N_15929,N_15952);
nor U16112 (N_16112,N_15993,N_15895);
nor U16113 (N_16113,N_15674,N_15784);
and U16114 (N_16114,N_15635,N_15968);
and U16115 (N_16115,N_15842,N_15836);
nand U16116 (N_16116,N_15911,N_15698);
nand U16117 (N_16117,N_15828,N_15777);
nor U16118 (N_16118,N_15864,N_15731);
nor U16119 (N_16119,N_15868,N_15726);
nor U16120 (N_16120,N_15680,N_15733);
and U16121 (N_16121,N_15872,N_15874);
and U16122 (N_16122,N_15766,N_15831);
nand U16123 (N_16123,N_15770,N_15666);
nor U16124 (N_16124,N_15714,N_15721);
nand U16125 (N_16125,N_15662,N_15949);
or U16126 (N_16126,N_15689,N_15617);
and U16127 (N_16127,N_15719,N_15955);
nand U16128 (N_16128,N_15649,N_15765);
xnor U16129 (N_16129,N_15618,N_15678);
or U16130 (N_16130,N_15694,N_15958);
xor U16131 (N_16131,N_15700,N_15800);
nor U16132 (N_16132,N_15743,N_15615);
nor U16133 (N_16133,N_15951,N_15710);
xor U16134 (N_16134,N_15604,N_15732);
xor U16135 (N_16135,N_15758,N_15802);
nor U16136 (N_16136,N_15865,N_15979);
and U16137 (N_16137,N_15806,N_15986);
xnor U16138 (N_16138,N_15835,N_15744);
or U16139 (N_16139,N_15866,N_15764);
xnor U16140 (N_16140,N_15606,N_15773);
and U16141 (N_16141,N_15922,N_15970);
xor U16142 (N_16142,N_15967,N_15780);
and U16143 (N_16143,N_15847,N_15772);
xor U16144 (N_16144,N_15737,N_15625);
xnor U16145 (N_16145,N_15981,N_15825);
xnor U16146 (N_16146,N_15717,N_15706);
nand U16147 (N_16147,N_15947,N_15844);
and U16148 (N_16148,N_15774,N_15969);
nand U16149 (N_16149,N_15751,N_15926);
nand U16150 (N_16150,N_15846,N_15881);
nand U16151 (N_16151,N_15613,N_15878);
and U16152 (N_16152,N_15797,N_15918);
nor U16153 (N_16153,N_15727,N_15757);
xnor U16154 (N_16154,N_15760,N_15788);
or U16155 (N_16155,N_15786,N_15998);
xnor U16156 (N_16156,N_15860,N_15644);
nor U16157 (N_16157,N_15887,N_15655);
nand U16158 (N_16158,N_15771,N_15775);
nand U16159 (N_16159,N_15639,N_15964);
xor U16160 (N_16160,N_15794,N_15653);
or U16161 (N_16161,N_15657,N_15734);
nand U16162 (N_16162,N_15904,N_15735);
xor U16163 (N_16163,N_15945,N_15937);
or U16164 (N_16164,N_15669,N_15841);
nand U16165 (N_16165,N_15902,N_15960);
and U16166 (N_16166,N_15974,N_15636);
nand U16167 (N_16167,N_15807,N_15624);
nor U16168 (N_16168,N_15977,N_15783);
and U16169 (N_16169,N_15834,N_15959);
or U16170 (N_16170,N_15824,N_15614);
nor U16171 (N_16171,N_15880,N_15809);
xor U16172 (N_16172,N_15626,N_15718);
xnor U16173 (N_16173,N_15948,N_15855);
nand U16174 (N_16174,N_15616,N_15822);
nand U16175 (N_16175,N_15965,N_15670);
and U16176 (N_16176,N_15601,N_15898);
nor U16177 (N_16177,N_15944,N_15931);
and U16178 (N_16178,N_15720,N_15988);
nor U16179 (N_16179,N_15871,N_15602);
or U16180 (N_16180,N_15798,N_15789);
or U16181 (N_16181,N_15849,N_15713);
and U16182 (N_16182,N_15830,N_15816);
nor U16183 (N_16183,N_15650,N_15641);
nor U16184 (N_16184,N_15909,N_15787);
and U16185 (N_16185,N_15656,N_15659);
and U16186 (N_16186,N_15745,N_15985);
xnor U16187 (N_16187,N_15975,N_15632);
or U16188 (N_16188,N_15927,N_15638);
nor U16189 (N_16189,N_15978,N_15920);
nor U16190 (N_16190,N_15961,N_15983);
and U16191 (N_16191,N_15673,N_15934);
nor U16192 (N_16192,N_15651,N_15900);
or U16193 (N_16193,N_15990,N_15879);
xor U16194 (N_16194,N_15685,N_15924);
nand U16195 (N_16195,N_15982,N_15701);
nor U16196 (N_16196,N_15963,N_15852);
or U16197 (N_16197,N_15896,N_15782);
xnor U16198 (N_16198,N_15913,N_15862);
or U16199 (N_16199,N_15621,N_15938);
or U16200 (N_16200,N_15659,N_15950);
xor U16201 (N_16201,N_15796,N_15902);
or U16202 (N_16202,N_15839,N_15663);
and U16203 (N_16203,N_15815,N_15998);
xnor U16204 (N_16204,N_15959,N_15704);
nand U16205 (N_16205,N_15736,N_15929);
xnor U16206 (N_16206,N_15821,N_15824);
xor U16207 (N_16207,N_15826,N_15715);
or U16208 (N_16208,N_15607,N_15622);
or U16209 (N_16209,N_15945,N_15687);
or U16210 (N_16210,N_15727,N_15746);
xnor U16211 (N_16211,N_15912,N_15904);
and U16212 (N_16212,N_15815,N_15648);
nor U16213 (N_16213,N_15615,N_15792);
nor U16214 (N_16214,N_15682,N_15769);
xor U16215 (N_16215,N_15682,N_15814);
nor U16216 (N_16216,N_15920,N_15756);
nand U16217 (N_16217,N_15784,N_15738);
xnor U16218 (N_16218,N_15678,N_15617);
or U16219 (N_16219,N_15820,N_15772);
nor U16220 (N_16220,N_15768,N_15997);
nor U16221 (N_16221,N_15630,N_15684);
nand U16222 (N_16222,N_15796,N_15863);
nor U16223 (N_16223,N_15785,N_15799);
xnor U16224 (N_16224,N_15627,N_15904);
and U16225 (N_16225,N_15901,N_15727);
and U16226 (N_16226,N_15817,N_15797);
xnor U16227 (N_16227,N_15926,N_15614);
xnor U16228 (N_16228,N_15675,N_15912);
and U16229 (N_16229,N_15720,N_15833);
xnor U16230 (N_16230,N_15916,N_15753);
xor U16231 (N_16231,N_15721,N_15823);
or U16232 (N_16232,N_15822,N_15930);
and U16233 (N_16233,N_15770,N_15671);
and U16234 (N_16234,N_15661,N_15942);
nor U16235 (N_16235,N_15930,N_15914);
nor U16236 (N_16236,N_15970,N_15864);
or U16237 (N_16237,N_15801,N_15971);
xor U16238 (N_16238,N_15746,N_15905);
nor U16239 (N_16239,N_15602,N_15696);
nor U16240 (N_16240,N_15613,N_15841);
xnor U16241 (N_16241,N_15656,N_15795);
xnor U16242 (N_16242,N_15626,N_15938);
nand U16243 (N_16243,N_15962,N_15827);
or U16244 (N_16244,N_15948,N_15938);
or U16245 (N_16245,N_15873,N_15917);
and U16246 (N_16246,N_15957,N_15833);
and U16247 (N_16247,N_15981,N_15812);
and U16248 (N_16248,N_15642,N_15896);
and U16249 (N_16249,N_15740,N_15681);
nand U16250 (N_16250,N_15814,N_15622);
and U16251 (N_16251,N_15885,N_15682);
xnor U16252 (N_16252,N_15821,N_15833);
xor U16253 (N_16253,N_15963,N_15629);
and U16254 (N_16254,N_15704,N_15870);
xnor U16255 (N_16255,N_15743,N_15753);
xor U16256 (N_16256,N_15725,N_15909);
nand U16257 (N_16257,N_15636,N_15856);
and U16258 (N_16258,N_15704,N_15819);
xnor U16259 (N_16259,N_15761,N_15723);
nand U16260 (N_16260,N_15721,N_15617);
nor U16261 (N_16261,N_15877,N_15779);
or U16262 (N_16262,N_15989,N_15817);
xnor U16263 (N_16263,N_15984,N_15837);
or U16264 (N_16264,N_15822,N_15987);
or U16265 (N_16265,N_15730,N_15809);
nor U16266 (N_16266,N_15847,N_15960);
and U16267 (N_16267,N_15748,N_15827);
and U16268 (N_16268,N_15952,N_15917);
or U16269 (N_16269,N_15667,N_15635);
and U16270 (N_16270,N_15986,N_15682);
nor U16271 (N_16271,N_15873,N_15600);
xnor U16272 (N_16272,N_15671,N_15734);
and U16273 (N_16273,N_15836,N_15761);
xnor U16274 (N_16274,N_15926,N_15884);
nor U16275 (N_16275,N_15704,N_15898);
and U16276 (N_16276,N_15785,N_15634);
or U16277 (N_16277,N_15865,N_15699);
and U16278 (N_16278,N_15632,N_15801);
xnor U16279 (N_16279,N_15915,N_15740);
xor U16280 (N_16280,N_15601,N_15665);
nand U16281 (N_16281,N_15825,N_15767);
nor U16282 (N_16282,N_15701,N_15977);
xor U16283 (N_16283,N_15751,N_15931);
nand U16284 (N_16284,N_15860,N_15982);
nand U16285 (N_16285,N_15636,N_15820);
xnor U16286 (N_16286,N_15878,N_15786);
or U16287 (N_16287,N_15941,N_15915);
and U16288 (N_16288,N_15775,N_15882);
xor U16289 (N_16289,N_15702,N_15680);
or U16290 (N_16290,N_15966,N_15819);
and U16291 (N_16291,N_15623,N_15844);
xor U16292 (N_16292,N_15832,N_15777);
and U16293 (N_16293,N_15754,N_15841);
or U16294 (N_16294,N_15733,N_15699);
nand U16295 (N_16295,N_15641,N_15890);
and U16296 (N_16296,N_15825,N_15933);
xor U16297 (N_16297,N_15640,N_15965);
nand U16298 (N_16298,N_15615,N_15692);
xor U16299 (N_16299,N_15837,N_15908);
nand U16300 (N_16300,N_15841,N_15693);
and U16301 (N_16301,N_15867,N_15673);
nor U16302 (N_16302,N_15664,N_15710);
and U16303 (N_16303,N_15842,N_15815);
and U16304 (N_16304,N_15942,N_15838);
nand U16305 (N_16305,N_15836,N_15945);
nand U16306 (N_16306,N_15704,N_15687);
nand U16307 (N_16307,N_15687,N_15700);
xnor U16308 (N_16308,N_15759,N_15753);
nor U16309 (N_16309,N_15917,N_15863);
xnor U16310 (N_16310,N_15692,N_15954);
or U16311 (N_16311,N_15893,N_15909);
and U16312 (N_16312,N_15832,N_15627);
xor U16313 (N_16313,N_15649,N_15795);
nand U16314 (N_16314,N_15848,N_15827);
and U16315 (N_16315,N_15891,N_15631);
nor U16316 (N_16316,N_15974,N_15992);
nand U16317 (N_16317,N_15745,N_15713);
and U16318 (N_16318,N_15760,N_15841);
or U16319 (N_16319,N_15822,N_15652);
nor U16320 (N_16320,N_15739,N_15853);
xnor U16321 (N_16321,N_15741,N_15634);
nand U16322 (N_16322,N_15875,N_15930);
nor U16323 (N_16323,N_15639,N_15609);
xnor U16324 (N_16324,N_15939,N_15663);
nor U16325 (N_16325,N_15854,N_15870);
nor U16326 (N_16326,N_15977,N_15932);
or U16327 (N_16327,N_15975,N_15813);
nor U16328 (N_16328,N_15764,N_15975);
or U16329 (N_16329,N_15622,N_15762);
nor U16330 (N_16330,N_15656,N_15602);
nand U16331 (N_16331,N_15971,N_15754);
nand U16332 (N_16332,N_15742,N_15696);
xnor U16333 (N_16333,N_15864,N_15968);
nor U16334 (N_16334,N_15625,N_15778);
xnor U16335 (N_16335,N_15864,N_15602);
xor U16336 (N_16336,N_15994,N_15703);
nor U16337 (N_16337,N_15766,N_15883);
and U16338 (N_16338,N_15718,N_15651);
nor U16339 (N_16339,N_15881,N_15992);
xnor U16340 (N_16340,N_15715,N_15847);
nand U16341 (N_16341,N_15605,N_15807);
and U16342 (N_16342,N_15885,N_15700);
nor U16343 (N_16343,N_15689,N_15616);
and U16344 (N_16344,N_15675,N_15701);
nor U16345 (N_16345,N_15970,N_15787);
and U16346 (N_16346,N_15914,N_15830);
nand U16347 (N_16347,N_15887,N_15727);
nand U16348 (N_16348,N_15885,N_15647);
nand U16349 (N_16349,N_15788,N_15796);
and U16350 (N_16350,N_15831,N_15832);
xnor U16351 (N_16351,N_15682,N_15992);
xor U16352 (N_16352,N_15884,N_15711);
and U16353 (N_16353,N_15970,N_15956);
nand U16354 (N_16354,N_15829,N_15945);
or U16355 (N_16355,N_15726,N_15637);
nor U16356 (N_16356,N_15903,N_15838);
xor U16357 (N_16357,N_15842,N_15637);
and U16358 (N_16358,N_15676,N_15716);
nor U16359 (N_16359,N_15942,N_15997);
or U16360 (N_16360,N_15935,N_15902);
and U16361 (N_16361,N_15631,N_15604);
nand U16362 (N_16362,N_15818,N_15896);
nor U16363 (N_16363,N_15892,N_15830);
nor U16364 (N_16364,N_15806,N_15730);
and U16365 (N_16365,N_15918,N_15686);
nor U16366 (N_16366,N_15712,N_15896);
nor U16367 (N_16367,N_15761,N_15902);
or U16368 (N_16368,N_15844,N_15634);
or U16369 (N_16369,N_15965,N_15756);
nand U16370 (N_16370,N_15786,N_15968);
xnor U16371 (N_16371,N_15998,N_15918);
or U16372 (N_16372,N_15887,N_15754);
nand U16373 (N_16373,N_15766,N_15985);
nor U16374 (N_16374,N_15840,N_15663);
xor U16375 (N_16375,N_15794,N_15940);
or U16376 (N_16376,N_15839,N_15936);
nand U16377 (N_16377,N_15874,N_15651);
nand U16378 (N_16378,N_15915,N_15728);
xor U16379 (N_16379,N_15931,N_15887);
xnor U16380 (N_16380,N_15756,N_15610);
nand U16381 (N_16381,N_15879,N_15998);
xor U16382 (N_16382,N_15717,N_15957);
and U16383 (N_16383,N_15659,N_15785);
or U16384 (N_16384,N_15908,N_15624);
and U16385 (N_16385,N_15695,N_15985);
and U16386 (N_16386,N_15613,N_15914);
and U16387 (N_16387,N_15859,N_15840);
or U16388 (N_16388,N_15754,N_15906);
nand U16389 (N_16389,N_15653,N_15988);
or U16390 (N_16390,N_15689,N_15910);
xor U16391 (N_16391,N_15914,N_15881);
nand U16392 (N_16392,N_15688,N_15898);
xnor U16393 (N_16393,N_15665,N_15840);
xor U16394 (N_16394,N_15760,N_15986);
nor U16395 (N_16395,N_15761,N_15974);
xnor U16396 (N_16396,N_15814,N_15944);
xnor U16397 (N_16397,N_15997,N_15948);
or U16398 (N_16398,N_15763,N_15626);
nor U16399 (N_16399,N_15626,N_15826);
xor U16400 (N_16400,N_16036,N_16386);
or U16401 (N_16401,N_16122,N_16365);
xnor U16402 (N_16402,N_16267,N_16177);
xnor U16403 (N_16403,N_16079,N_16395);
nor U16404 (N_16404,N_16082,N_16352);
xnor U16405 (N_16405,N_16038,N_16102);
nand U16406 (N_16406,N_16289,N_16140);
nand U16407 (N_16407,N_16183,N_16347);
nand U16408 (N_16408,N_16203,N_16327);
nor U16409 (N_16409,N_16174,N_16076);
nor U16410 (N_16410,N_16005,N_16092);
nand U16411 (N_16411,N_16078,N_16053);
xor U16412 (N_16412,N_16153,N_16287);
xnor U16413 (N_16413,N_16108,N_16339);
nand U16414 (N_16414,N_16179,N_16193);
and U16415 (N_16415,N_16201,N_16143);
or U16416 (N_16416,N_16310,N_16228);
or U16417 (N_16417,N_16266,N_16240);
xnor U16418 (N_16418,N_16253,N_16272);
nor U16419 (N_16419,N_16305,N_16090);
and U16420 (N_16420,N_16112,N_16012);
and U16421 (N_16421,N_16060,N_16222);
and U16422 (N_16422,N_16227,N_16202);
xnor U16423 (N_16423,N_16151,N_16009);
or U16424 (N_16424,N_16098,N_16093);
nor U16425 (N_16425,N_16200,N_16084);
or U16426 (N_16426,N_16042,N_16043);
nand U16427 (N_16427,N_16166,N_16110);
nor U16428 (N_16428,N_16070,N_16215);
nor U16429 (N_16429,N_16231,N_16329);
nand U16430 (N_16430,N_16320,N_16398);
or U16431 (N_16431,N_16069,N_16354);
and U16432 (N_16432,N_16191,N_16141);
or U16433 (N_16433,N_16261,N_16360);
nand U16434 (N_16434,N_16382,N_16373);
nor U16435 (N_16435,N_16198,N_16045);
xor U16436 (N_16436,N_16158,N_16099);
or U16437 (N_16437,N_16384,N_16381);
nand U16438 (N_16438,N_16019,N_16323);
and U16439 (N_16439,N_16337,N_16181);
and U16440 (N_16440,N_16243,N_16216);
nor U16441 (N_16441,N_16195,N_16057);
nand U16442 (N_16442,N_16309,N_16107);
xor U16443 (N_16443,N_16233,N_16121);
and U16444 (N_16444,N_16361,N_16212);
or U16445 (N_16445,N_16029,N_16376);
and U16446 (N_16446,N_16031,N_16318);
nor U16447 (N_16447,N_16000,N_16189);
xor U16448 (N_16448,N_16375,N_16250);
xor U16449 (N_16449,N_16213,N_16338);
nand U16450 (N_16450,N_16173,N_16259);
nand U16451 (N_16451,N_16109,N_16255);
nor U16452 (N_16452,N_16378,N_16159);
nand U16453 (N_16453,N_16073,N_16188);
nor U16454 (N_16454,N_16308,N_16163);
or U16455 (N_16455,N_16316,N_16169);
and U16456 (N_16456,N_16097,N_16363);
xnor U16457 (N_16457,N_16142,N_16147);
or U16458 (N_16458,N_16127,N_16358);
nand U16459 (N_16459,N_16370,N_16271);
xnor U16460 (N_16460,N_16154,N_16172);
xor U16461 (N_16461,N_16155,N_16218);
xor U16462 (N_16462,N_16303,N_16364);
and U16463 (N_16463,N_16291,N_16392);
nor U16464 (N_16464,N_16377,N_16088);
xnor U16465 (N_16465,N_16391,N_16044);
nor U16466 (N_16466,N_16294,N_16314);
and U16467 (N_16467,N_16221,N_16219);
or U16468 (N_16468,N_16390,N_16299);
or U16469 (N_16469,N_16171,N_16344);
nor U16470 (N_16470,N_16349,N_16055);
nor U16471 (N_16471,N_16238,N_16257);
nor U16472 (N_16472,N_16254,N_16351);
nand U16473 (N_16473,N_16049,N_16230);
xnor U16474 (N_16474,N_16126,N_16283);
nor U16475 (N_16475,N_16348,N_16023);
or U16476 (N_16476,N_16286,N_16194);
nor U16477 (N_16477,N_16371,N_16260);
nor U16478 (N_16478,N_16342,N_16024);
nor U16479 (N_16479,N_16292,N_16041);
nor U16480 (N_16480,N_16282,N_16379);
or U16481 (N_16481,N_16207,N_16214);
or U16482 (N_16482,N_16116,N_16295);
and U16483 (N_16483,N_16077,N_16011);
nor U16484 (N_16484,N_16085,N_16311);
nor U16485 (N_16485,N_16176,N_16130);
or U16486 (N_16486,N_16313,N_16087);
nor U16487 (N_16487,N_16357,N_16321);
or U16488 (N_16488,N_16333,N_16039);
or U16489 (N_16489,N_16072,N_16026);
or U16490 (N_16490,N_16262,N_16270);
xnor U16491 (N_16491,N_16100,N_16054);
xnor U16492 (N_16492,N_16119,N_16008);
and U16493 (N_16493,N_16325,N_16046);
nand U16494 (N_16494,N_16284,N_16236);
xor U16495 (N_16495,N_16205,N_16035);
and U16496 (N_16496,N_16242,N_16144);
nor U16497 (N_16497,N_16280,N_16341);
or U16498 (N_16498,N_16185,N_16335);
and U16499 (N_16499,N_16014,N_16385);
nor U16500 (N_16500,N_16156,N_16393);
or U16501 (N_16501,N_16106,N_16134);
xnor U16502 (N_16502,N_16224,N_16302);
nor U16503 (N_16503,N_16010,N_16315);
nor U16504 (N_16504,N_16182,N_16372);
and U16505 (N_16505,N_16288,N_16190);
xnor U16506 (N_16506,N_16170,N_16001);
nor U16507 (N_16507,N_16204,N_16160);
and U16508 (N_16508,N_16196,N_16133);
nor U16509 (N_16509,N_16138,N_16276);
or U16510 (N_16510,N_16091,N_16150);
and U16511 (N_16511,N_16317,N_16178);
or U16512 (N_16512,N_16394,N_16388);
nor U16513 (N_16513,N_16269,N_16004);
xor U16514 (N_16514,N_16186,N_16326);
and U16515 (N_16515,N_16152,N_16387);
xor U16516 (N_16516,N_16293,N_16145);
xnor U16517 (N_16517,N_16080,N_16273);
nor U16518 (N_16518,N_16263,N_16033);
or U16519 (N_16519,N_16232,N_16022);
or U16520 (N_16520,N_16247,N_16265);
xnor U16521 (N_16521,N_16050,N_16094);
and U16522 (N_16522,N_16223,N_16075);
xnor U16523 (N_16523,N_16148,N_16345);
or U16524 (N_16524,N_16244,N_16165);
nor U16525 (N_16525,N_16021,N_16251);
xor U16526 (N_16526,N_16312,N_16211);
nand U16527 (N_16527,N_16346,N_16275);
nand U16528 (N_16528,N_16324,N_16331);
nor U16529 (N_16529,N_16047,N_16307);
nor U16530 (N_16530,N_16301,N_16355);
and U16531 (N_16531,N_16383,N_16278);
nand U16532 (N_16532,N_16034,N_16058);
nand U16533 (N_16533,N_16281,N_16131);
nand U16534 (N_16534,N_16086,N_16359);
nand U16535 (N_16535,N_16180,N_16319);
xnor U16536 (N_16536,N_16258,N_16064);
nor U16537 (N_16537,N_16062,N_16128);
xnor U16538 (N_16538,N_16328,N_16268);
xnor U16539 (N_16539,N_16322,N_16210);
nor U16540 (N_16540,N_16399,N_16040);
or U16541 (N_16541,N_16096,N_16113);
or U16542 (N_16542,N_16051,N_16139);
and U16543 (N_16543,N_16118,N_16208);
and U16544 (N_16544,N_16175,N_16095);
or U16545 (N_16545,N_16115,N_16229);
or U16546 (N_16546,N_16380,N_16123);
or U16547 (N_16547,N_16068,N_16157);
nor U16548 (N_16548,N_16374,N_16340);
xor U16549 (N_16549,N_16300,N_16330);
or U16550 (N_16550,N_16016,N_16225);
nor U16551 (N_16551,N_16356,N_16248);
or U16552 (N_16552,N_16239,N_16002);
nand U16553 (N_16553,N_16074,N_16006);
nor U16554 (N_16554,N_16013,N_16350);
nand U16555 (N_16555,N_16264,N_16056);
nand U16556 (N_16556,N_16018,N_16114);
nand U16557 (N_16557,N_16071,N_16162);
and U16558 (N_16558,N_16135,N_16149);
xnor U16559 (N_16559,N_16184,N_16048);
and U16560 (N_16560,N_16111,N_16298);
nor U16561 (N_16561,N_16332,N_16164);
xnor U16562 (N_16562,N_16066,N_16161);
or U16563 (N_16563,N_16199,N_16105);
xnor U16564 (N_16564,N_16396,N_16003);
nor U16565 (N_16565,N_16132,N_16187);
nor U16566 (N_16566,N_16304,N_16030);
or U16567 (N_16567,N_16290,N_16274);
or U16568 (N_16568,N_16343,N_16129);
or U16569 (N_16569,N_16197,N_16025);
or U16570 (N_16570,N_16032,N_16168);
or U16571 (N_16571,N_16277,N_16027);
nand U16572 (N_16572,N_16083,N_16081);
and U16573 (N_16573,N_16124,N_16353);
nor U16574 (N_16574,N_16117,N_16279);
nand U16575 (N_16575,N_16120,N_16146);
or U16576 (N_16576,N_16063,N_16245);
nor U16577 (N_16577,N_16296,N_16028);
xor U16578 (N_16578,N_16235,N_16252);
xor U16579 (N_16579,N_16061,N_16104);
and U16580 (N_16580,N_16241,N_16256);
nand U16581 (N_16581,N_16020,N_16246);
nand U16582 (N_16582,N_16015,N_16067);
or U16583 (N_16583,N_16369,N_16334);
nor U16584 (N_16584,N_16237,N_16397);
and U16585 (N_16585,N_16103,N_16249);
nand U16586 (N_16586,N_16285,N_16368);
xnor U16587 (N_16587,N_16389,N_16125);
xor U16588 (N_16588,N_16234,N_16206);
or U16589 (N_16589,N_16220,N_16217);
or U16590 (N_16590,N_16366,N_16059);
xnor U16591 (N_16591,N_16226,N_16336);
nand U16592 (N_16592,N_16007,N_16101);
xnor U16593 (N_16593,N_16362,N_16137);
nor U16594 (N_16594,N_16017,N_16052);
xor U16595 (N_16595,N_16065,N_16367);
nand U16596 (N_16596,N_16136,N_16297);
nand U16597 (N_16597,N_16167,N_16306);
and U16598 (N_16598,N_16192,N_16209);
or U16599 (N_16599,N_16089,N_16037);
xor U16600 (N_16600,N_16293,N_16047);
or U16601 (N_16601,N_16328,N_16064);
nand U16602 (N_16602,N_16336,N_16114);
and U16603 (N_16603,N_16289,N_16310);
xor U16604 (N_16604,N_16391,N_16302);
and U16605 (N_16605,N_16099,N_16390);
xor U16606 (N_16606,N_16292,N_16035);
or U16607 (N_16607,N_16060,N_16328);
xor U16608 (N_16608,N_16016,N_16078);
and U16609 (N_16609,N_16174,N_16051);
nand U16610 (N_16610,N_16399,N_16349);
xnor U16611 (N_16611,N_16261,N_16061);
xor U16612 (N_16612,N_16010,N_16041);
nor U16613 (N_16613,N_16181,N_16008);
nand U16614 (N_16614,N_16232,N_16369);
nand U16615 (N_16615,N_16240,N_16167);
nor U16616 (N_16616,N_16329,N_16283);
nand U16617 (N_16617,N_16165,N_16228);
or U16618 (N_16618,N_16018,N_16235);
or U16619 (N_16619,N_16367,N_16238);
nor U16620 (N_16620,N_16234,N_16223);
or U16621 (N_16621,N_16018,N_16252);
xnor U16622 (N_16622,N_16367,N_16000);
or U16623 (N_16623,N_16099,N_16313);
xor U16624 (N_16624,N_16322,N_16233);
or U16625 (N_16625,N_16359,N_16158);
and U16626 (N_16626,N_16155,N_16088);
xnor U16627 (N_16627,N_16295,N_16330);
nor U16628 (N_16628,N_16120,N_16370);
nand U16629 (N_16629,N_16282,N_16075);
nor U16630 (N_16630,N_16143,N_16320);
xnor U16631 (N_16631,N_16201,N_16313);
xor U16632 (N_16632,N_16324,N_16084);
xor U16633 (N_16633,N_16082,N_16298);
or U16634 (N_16634,N_16189,N_16100);
nand U16635 (N_16635,N_16030,N_16028);
or U16636 (N_16636,N_16313,N_16154);
nor U16637 (N_16637,N_16307,N_16016);
or U16638 (N_16638,N_16397,N_16091);
xor U16639 (N_16639,N_16247,N_16283);
nand U16640 (N_16640,N_16192,N_16152);
nor U16641 (N_16641,N_16104,N_16339);
nor U16642 (N_16642,N_16082,N_16256);
or U16643 (N_16643,N_16305,N_16284);
xnor U16644 (N_16644,N_16267,N_16115);
and U16645 (N_16645,N_16284,N_16375);
xor U16646 (N_16646,N_16001,N_16084);
xor U16647 (N_16647,N_16031,N_16346);
xor U16648 (N_16648,N_16146,N_16297);
or U16649 (N_16649,N_16133,N_16387);
nand U16650 (N_16650,N_16265,N_16360);
nor U16651 (N_16651,N_16067,N_16138);
nor U16652 (N_16652,N_16217,N_16380);
and U16653 (N_16653,N_16313,N_16121);
nor U16654 (N_16654,N_16236,N_16136);
nor U16655 (N_16655,N_16246,N_16261);
xor U16656 (N_16656,N_16096,N_16026);
or U16657 (N_16657,N_16301,N_16190);
and U16658 (N_16658,N_16003,N_16149);
nor U16659 (N_16659,N_16180,N_16387);
or U16660 (N_16660,N_16320,N_16139);
xor U16661 (N_16661,N_16200,N_16392);
nand U16662 (N_16662,N_16358,N_16131);
and U16663 (N_16663,N_16160,N_16277);
and U16664 (N_16664,N_16018,N_16361);
xor U16665 (N_16665,N_16188,N_16330);
xnor U16666 (N_16666,N_16255,N_16260);
and U16667 (N_16667,N_16109,N_16327);
and U16668 (N_16668,N_16278,N_16314);
nand U16669 (N_16669,N_16160,N_16035);
nand U16670 (N_16670,N_16191,N_16252);
or U16671 (N_16671,N_16313,N_16037);
or U16672 (N_16672,N_16301,N_16296);
or U16673 (N_16673,N_16344,N_16069);
and U16674 (N_16674,N_16158,N_16284);
and U16675 (N_16675,N_16128,N_16327);
xnor U16676 (N_16676,N_16095,N_16036);
xor U16677 (N_16677,N_16209,N_16343);
and U16678 (N_16678,N_16225,N_16361);
and U16679 (N_16679,N_16120,N_16160);
nor U16680 (N_16680,N_16156,N_16034);
nand U16681 (N_16681,N_16185,N_16370);
nor U16682 (N_16682,N_16356,N_16040);
or U16683 (N_16683,N_16213,N_16385);
nor U16684 (N_16684,N_16294,N_16186);
nor U16685 (N_16685,N_16389,N_16286);
xor U16686 (N_16686,N_16281,N_16257);
nor U16687 (N_16687,N_16317,N_16080);
xnor U16688 (N_16688,N_16296,N_16371);
xor U16689 (N_16689,N_16200,N_16305);
xor U16690 (N_16690,N_16379,N_16175);
nand U16691 (N_16691,N_16152,N_16369);
xor U16692 (N_16692,N_16101,N_16295);
and U16693 (N_16693,N_16306,N_16100);
or U16694 (N_16694,N_16170,N_16272);
and U16695 (N_16695,N_16163,N_16327);
nor U16696 (N_16696,N_16204,N_16117);
xor U16697 (N_16697,N_16240,N_16232);
and U16698 (N_16698,N_16365,N_16248);
nand U16699 (N_16699,N_16216,N_16347);
nand U16700 (N_16700,N_16135,N_16195);
and U16701 (N_16701,N_16030,N_16262);
nand U16702 (N_16702,N_16388,N_16385);
and U16703 (N_16703,N_16156,N_16378);
or U16704 (N_16704,N_16088,N_16244);
and U16705 (N_16705,N_16064,N_16034);
and U16706 (N_16706,N_16255,N_16137);
nand U16707 (N_16707,N_16261,N_16280);
xor U16708 (N_16708,N_16354,N_16356);
or U16709 (N_16709,N_16318,N_16289);
or U16710 (N_16710,N_16069,N_16047);
nand U16711 (N_16711,N_16304,N_16034);
xnor U16712 (N_16712,N_16184,N_16270);
and U16713 (N_16713,N_16395,N_16026);
nand U16714 (N_16714,N_16004,N_16113);
xor U16715 (N_16715,N_16300,N_16285);
nor U16716 (N_16716,N_16315,N_16015);
or U16717 (N_16717,N_16159,N_16033);
nand U16718 (N_16718,N_16054,N_16007);
and U16719 (N_16719,N_16009,N_16136);
nand U16720 (N_16720,N_16292,N_16177);
xor U16721 (N_16721,N_16095,N_16301);
or U16722 (N_16722,N_16318,N_16050);
nand U16723 (N_16723,N_16038,N_16349);
nand U16724 (N_16724,N_16144,N_16325);
and U16725 (N_16725,N_16185,N_16197);
and U16726 (N_16726,N_16098,N_16104);
and U16727 (N_16727,N_16063,N_16036);
xor U16728 (N_16728,N_16206,N_16319);
nor U16729 (N_16729,N_16325,N_16374);
or U16730 (N_16730,N_16045,N_16073);
nor U16731 (N_16731,N_16057,N_16100);
and U16732 (N_16732,N_16017,N_16356);
and U16733 (N_16733,N_16296,N_16211);
xor U16734 (N_16734,N_16256,N_16270);
xnor U16735 (N_16735,N_16022,N_16160);
nand U16736 (N_16736,N_16016,N_16035);
xnor U16737 (N_16737,N_16014,N_16329);
nand U16738 (N_16738,N_16044,N_16200);
or U16739 (N_16739,N_16121,N_16193);
xnor U16740 (N_16740,N_16324,N_16254);
nor U16741 (N_16741,N_16041,N_16253);
or U16742 (N_16742,N_16051,N_16310);
and U16743 (N_16743,N_16183,N_16186);
or U16744 (N_16744,N_16019,N_16351);
nand U16745 (N_16745,N_16398,N_16111);
or U16746 (N_16746,N_16313,N_16004);
nand U16747 (N_16747,N_16186,N_16181);
nor U16748 (N_16748,N_16248,N_16068);
nand U16749 (N_16749,N_16282,N_16328);
or U16750 (N_16750,N_16161,N_16352);
nand U16751 (N_16751,N_16362,N_16230);
or U16752 (N_16752,N_16295,N_16034);
xor U16753 (N_16753,N_16230,N_16373);
xnor U16754 (N_16754,N_16284,N_16041);
or U16755 (N_16755,N_16194,N_16128);
nand U16756 (N_16756,N_16091,N_16278);
and U16757 (N_16757,N_16000,N_16248);
nand U16758 (N_16758,N_16082,N_16239);
nand U16759 (N_16759,N_16212,N_16021);
xnor U16760 (N_16760,N_16117,N_16284);
or U16761 (N_16761,N_16145,N_16137);
nand U16762 (N_16762,N_16117,N_16250);
nor U16763 (N_16763,N_16123,N_16350);
nand U16764 (N_16764,N_16281,N_16158);
nor U16765 (N_16765,N_16148,N_16353);
or U16766 (N_16766,N_16023,N_16181);
xor U16767 (N_16767,N_16302,N_16184);
xor U16768 (N_16768,N_16321,N_16196);
nand U16769 (N_16769,N_16199,N_16280);
xnor U16770 (N_16770,N_16086,N_16127);
nor U16771 (N_16771,N_16385,N_16155);
or U16772 (N_16772,N_16352,N_16177);
or U16773 (N_16773,N_16102,N_16320);
and U16774 (N_16774,N_16009,N_16086);
nand U16775 (N_16775,N_16055,N_16259);
or U16776 (N_16776,N_16064,N_16338);
nand U16777 (N_16777,N_16354,N_16278);
xor U16778 (N_16778,N_16296,N_16120);
nor U16779 (N_16779,N_16279,N_16357);
xnor U16780 (N_16780,N_16085,N_16008);
nor U16781 (N_16781,N_16040,N_16353);
and U16782 (N_16782,N_16253,N_16019);
xnor U16783 (N_16783,N_16234,N_16368);
xnor U16784 (N_16784,N_16033,N_16068);
xnor U16785 (N_16785,N_16397,N_16383);
and U16786 (N_16786,N_16172,N_16127);
and U16787 (N_16787,N_16215,N_16342);
nor U16788 (N_16788,N_16308,N_16092);
nand U16789 (N_16789,N_16139,N_16059);
nor U16790 (N_16790,N_16102,N_16304);
or U16791 (N_16791,N_16032,N_16118);
and U16792 (N_16792,N_16255,N_16225);
or U16793 (N_16793,N_16307,N_16006);
or U16794 (N_16794,N_16317,N_16279);
or U16795 (N_16795,N_16081,N_16108);
xor U16796 (N_16796,N_16300,N_16365);
nor U16797 (N_16797,N_16092,N_16030);
nand U16798 (N_16798,N_16145,N_16302);
nor U16799 (N_16799,N_16357,N_16059);
or U16800 (N_16800,N_16417,N_16522);
nor U16801 (N_16801,N_16600,N_16794);
xor U16802 (N_16802,N_16619,N_16785);
nand U16803 (N_16803,N_16639,N_16728);
xnor U16804 (N_16804,N_16671,N_16769);
and U16805 (N_16805,N_16450,N_16451);
or U16806 (N_16806,N_16673,N_16449);
or U16807 (N_16807,N_16573,N_16756);
or U16808 (N_16808,N_16462,N_16496);
nor U16809 (N_16809,N_16730,N_16706);
nor U16810 (N_16810,N_16430,N_16718);
and U16811 (N_16811,N_16568,N_16519);
or U16812 (N_16812,N_16667,N_16615);
and U16813 (N_16813,N_16588,N_16646);
xor U16814 (N_16814,N_16484,N_16739);
xor U16815 (N_16815,N_16799,N_16777);
nor U16816 (N_16816,N_16761,N_16481);
nand U16817 (N_16817,N_16716,N_16796);
or U16818 (N_16818,N_16703,N_16604);
and U16819 (N_16819,N_16411,N_16784);
nor U16820 (N_16820,N_16658,N_16627);
or U16821 (N_16821,N_16712,N_16510);
xnor U16822 (N_16822,N_16578,N_16687);
or U16823 (N_16823,N_16762,N_16598);
nor U16824 (N_16824,N_16776,N_16743);
and U16825 (N_16825,N_16734,N_16680);
xnor U16826 (N_16826,N_16668,N_16518);
nor U16827 (N_16827,N_16798,N_16726);
and U16828 (N_16828,N_16638,N_16745);
or U16829 (N_16829,N_16684,N_16460);
nor U16830 (N_16830,N_16436,N_16714);
nand U16831 (N_16831,N_16674,N_16479);
nor U16832 (N_16832,N_16764,N_16515);
and U16833 (N_16833,N_16742,N_16523);
and U16834 (N_16834,N_16514,N_16421);
nand U16835 (N_16835,N_16640,N_16482);
nor U16836 (N_16836,N_16635,N_16404);
nor U16837 (N_16837,N_16550,N_16402);
xor U16838 (N_16838,N_16651,N_16786);
or U16839 (N_16839,N_16551,N_16661);
or U16840 (N_16840,N_16512,N_16401);
nor U16841 (N_16841,N_16704,N_16747);
nor U16842 (N_16842,N_16446,N_16613);
xor U16843 (N_16843,N_16771,N_16412);
nand U16844 (N_16844,N_16427,N_16746);
nand U16845 (N_16845,N_16547,N_16791);
and U16846 (N_16846,N_16490,N_16483);
and U16847 (N_16847,N_16531,N_16789);
or U16848 (N_16848,N_16538,N_16770);
xor U16849 (N_16849,N_16607,N_16763);
xnor U16850 (N_16850,N_16440,N_16662);
nor U16851 (N_16851,N_16602,N_16637);
nor U16852 (N_16852,N_16719,N_16526);
or U16853 (N_16853,N_16603,N_16608);
and U16854 (N_16854,N_16700,N_16583);
nand U16855 (N_16855,N_16541,N_16740);
xor U16856 (N_16856,N_16433,N_16609);
and U16857 (N_16857,N_16413,N_16783);
nand U16858 (N_16858,N_16597,N_16697);
xnor U16859 (N_16859,N_16779,N_16735);
xor U16860 (N_16860,N_16552,N_16408);
or U16861 (N_16861,N_16469,N_16498);
nand U16862 (N_16862,N_16790,N_16620);
or U16863 (N_16863,N_16675,N_16549);
nor U16864 (N_16864,N_16444,N_16470);
xor U16865 (N_16865,N_16766,N_16435);
nand U16866 (N_16866,N_16476,N_16400);
nor U16867 (N_16867,N_16618,N_16407);
nand U16868 (N_16868,N_16636,N_16591);
and U16869 (N_16869,N_16690,N_16467);
or U16870 (N_16870,N_16424,N_16774);
and U16871 (N_16871,N_16472,N_16453);
nand U16872 (N_16872,N_16447,N_16434);
nor U16873 (N_16873,N_16555,N_16582);
nor U16874 (N_16874,N_16775,N_16524);
nand U16875 (N_16875,N_16767,N_16688);
and U16876 (N_16876,N_16737,N_16557);
nor U16877 (N_16877,N_16452,N_16727);
nor U16878 (N_16878,N_16694,N_16581);
and U16879 (N_16879,N_16645,N_16669);
nand U16880 (N_16880,N_16649,N_16652);
nor U16881 (N_16881,N_16558,N_16681);
and U16882 (N_16882,N_16491,N_16502);
or U16883 (N_16883,N_16554,N_16773);
nand U16884 (N_16884,N_16748,N_16729);
xnor U16885 (N_16885,N_16660,N_16692);
xor U16886 (N_16886,N_16656,N_16503);
nor U16887 (N_16887,N_16702,N_16563);
nor U16888 (N_16888,N_16715,N_16647);
nor U16889 (N_16889,N_16631,N_16621);
or U16890 (N_16890,N_16448,N_16534);
or U16891 (N_16891,N_16527,N_16693);
nor U16892 (N_16892,N_16711,N_16787);
xnor U16893 (N_16893,N_16405,N_16439);
or U16894 (N_16894,N_16585,N_16454);
nor U16895 (N_16895,N_16612,N_16516);
xnor U16896 (N_16896,N_16504,N_16601);
or U16897 (N_16897,N_16574,N_16577);
or U16898 (N_16898,N_16463,N_16457);
xor U16899 (N_16899,N_16657,N_16626);
nor U16900 (N_16900,N_16713,N_16617);
nand U16901 (N_16901,N_16556,N_16757);
nand U16902 (N_16902,N_16717,N_16586);
and U16903 (N_16903,N_16486,N_16750);
nor U16904 (N_16904,N_16736,N_16533);
or U16905 (N_16905,N_16487,N_16493);
nor U16906 (N_16906,N_16576,N_16782);
and U16907 (N_16907,N_16724,N_16758);
nand U16908 (N_16908,N_16419,N_16642);
xnor U16909 (N_16909,N_16623,N_16501);
nand U16910 (N_16910,N_16475,N_16593);
xnor U16911 (N_16911,N_16422,N_16441);
nand U16912 (N_16912,N_16506,N_16723);
nand U16913 (N_16913,N_16543,N_16725);
nor U16914 (N_16914,N_16616,N_16478);
and U16915 (N_16915,N_16477,N_16529);
xor U16916 (N_16916,N_16664,N_16464);
nand U16917 (N_16917,N_16548,N_16732);
xnor U16918 (N_16918,N_16489,N_16511);
nor U16919 (N_16919,N_16553,N_16641);
nor U16920 (N_16920,N_16685,N_16765);
xor U16921 (N_16921,N_16753,N_16749);
xor U16922 (N_16922,N_16686,N_16471);
or U16923 (N_16923,N_16542,N_16629);
or U16924 (N_16924,N_16566,N_16455);
xnor U16925 (N_16925,N_16565,N_16445);
nor U16926 (N_16926,N_16569,N_16410);
and U16927 (N_16927,N_16517,N_16530);
nor U16928 (N_16928,N_16473,N_16691);
or U16929 (N_16929,N_16781,N_16495);
or U16930 (N_16930,N_16738,N_16525);
and U16931 (N_16931,N_16759,N_16420);
or U16932 (N_16932,N_16643,N_16676);
nand U16933 (N_16933,N_16438,N_16679);
xor U16934 (N_16934,N_16634,N_16611);
nand U16935 (N_16935,N_16442,N_16768);
xnor U16936 (N_16936,N_16705,N_16653);
and U16937 (N_16937,N_16429,N_16707);
and U16938 (N_16938,N_16494,N_16570);
and U16939 (N_16939,N_16710,N_16741);
and U16940 (N_16940,N_16605,N_16521);
or U16941 (N_16941,N_16670,N_16539);
nor U16942 (N_16942,N_16425,N_16468);
nor U16943 (N_16943,N_16443,N_16535);
xor U16944 (N_16944,N_16708,N_16579);
or U16945 (N_16945,N_16625,N_16701);
and U16946 (N_16946,N_16508,N_16428);
nand U16947 (N_16947,N_16650,N_16731);
nor U16948 (N_16948,N_16622,N_16423);
nand U16949 (N_16949,N_16696,N_16414);
nand U16950 (N_16950,N_16614,N_16461);
and U16951 (N_16951,N_16465,N_16418);
nand U16952 (N_16952,N_16666,N_16722);
xor U16953 (N_16953,N_16632,N_16561);
xor U16954 (N_16954,N_16540,N_16744);
or U16955 (N_16955,N_16683,N_16567);
or U16956 (N_16956,N_16572,N_16780);
nand U16957 (N_16957,N_16480,N_16492);
and U16958 (N_16958,N_16564,N_16596);
nand U16959 (N_16959,N_16456,N_16795);
or U16960 (N_16960,N_16584,N_16559);
xnor U16961 (N_16961,N_16532,N_16432);
or U16962 (N_16962,N_16590,N_16409);
nor U16963 (N_16963,N_16546,N_16458);
nor U16964 (N_16964,N_16499,N_16778);
xor U16965 (N_16965,N_16772,N_16474);
nand U16966 (N_16966,N_16431,N_16633);
nand U16967 (N_16967,N_16760,N_16695);
or U16968 (N_16968,N_16606,N_16507);
nor U16969 (N_16969,N_16665,N_16751);
xor U16970 (N_16970,N_16580,N_16406);
xor U16971 (N_16971,N_16720,N_16537);
xor U16972 (N_16972,N_16644,N_16677);
and U16973 (N_16973,N_16689,N_16509);
nor U16974 (N_16974,N_16466,N_16672);
or U16975 (N_16975,N_16416,N_16505);
or U16976 (N_16976,N_16793,N_16797);
and U16977 (N_16977,N_16699,N_16528);
and U16978 (N_16978,N_16698,N_16575);
nor U16979 (N_16979,N_16415,N_16500);
and U16980 (N_16980,N_16520,N_16513);
and U16981 (N_16981,N_16571,N_16709);
nand U16982 (N_16982,N_16426,N_16497);
nand U16983 (N_16983,N_16624,N_16792);
and U16984 (N_16984,N_16592,N_16536);
or U16985 (N_16985,N_16599,N_16587);
nor U16986 (N_16986,N_16721,N_16659);
or U16987 (N_16987,N_16545,N_16755);
or U16988 (N_16988,N_16610,N_16682);
nand U16989 (N_16989,N_16733,N_16663);
or U16990 (N_16990,N_16628,N_16560);
nand U16991 (N_16991,N_16459,N_16754);
xnor U16992 (N_16992,N_16544,N_16594);
and U16993 (N_16993,N_16562,N_16589);
nand U16994 (N_16994,N_16488,N_16655);
nand U16995 (N_16995,N_16630,N_16788);
or U16996 (N_16996,N_16485,N_16752);
and U16997 (N_16997,N_16403,N_16654);
nand U16998 (N_16998,N_16678,N_16648);
nand U16999 (N_16999,N_16437,N_16595);
nand U17000 (N_17000,N_16437,N_16428);
nor U17001 (N_17001,N_16655,N_16711);
nor U17002 (N_17002,N_16459,N_16464);
or U17003 (N_17003,N_16683,N_16410);
xor U17004 (N_17004,N_16427,N_16783);
or U17005 (N_17005,N_16798,N_16793);
nand U17006 (N_17006,N_16412,N_16433);
nand U17007 (N_17007,N_16536,N_16628);
and U17008 (N_17008,N_16680,N_16550);
and U17009 (N_17009,N_16564,N_16541);
nand U17010 (N_17010,N_16523,N_16658);
nor U17011 (N_17011,N_16787,N_16643);
nor U17012 (N_17012,N_16669,N_16601);
and U17013 (N_17013,N_16464,N_16515);
and U17014 (N_17014,N_16691,N_16746);
xnor U17015 (N_17015,N_16615,N_16581);
or U17016 (N_17016,N_16686,N_16696);
nand U17017 (N_17017,N_16415,N_16648);
nor U17018 (N_17018,N_16491,N_16410);
and U17019 (N_17019,N_16504,N_16668);
xor U17020 (N_17020,N_16720,N_16404);
nand U17021 (N_17021,N_16458,N_16669);
and U17022 (N_17022,N_16596,N_16533);
nand U17023 (N_17023,N_16495,N_16732);
and U17024 (N_17024,N_16766,N_16429);
or U17025 (N_17025,N_16550,N_16430);
and U17026 (N_17026,N_16520,N_16538);
xnor U17027 (N_17027,N_16739,N_16512);
and U17028 (N_17028,N_16444,N_16667);
and U17029 (N_17029,N_16479,N_16526);
nand U17030 (N_17030,N_16699,N_16525);
xor U17031 (N_17031,N_16756,N_16402);
or U17032 (N_17032,N_16682,N_16674);
and U17033 (N_17033,N_16648,N_16459);
nor U17034 (N_17034,N_16649,N_16411);
xnor U17035 (N_17035,N_16492,N_16789);
nor U17036 (N_17036,N_16506,N_16675);
nor U17037 (N_17037,N_16591,N_16703);
and U17038 (N_17038,N_16555,N_16461);
xnor U17039 (N_17039,N_16726,N_16767);
and U17040 (N_17040,N_16762,N_16508);
nand U17041 (N_17041,N_16736,N_16681);
and U17042 (N_17042,N_16450,N_16621);
or U17043 (N_17043,N_16723,N_16777);
or U17044 (N_17044,N_16770,N_16485);
xnor U17045 (N_17045,N_16507,N_16521);
or U17046 (N_17046,N_16419,N_16646);
xnor U17047 (N_17047,N_16773,N_16523);
or U17048 (N_17048,N_16471,N_16694);
nor U17049 (N_17049,N_16605,N_16608);
or U17050 (N_17050,N_16775,N_16650);
xor U17051 (N_17051,N_16532,N_16728);
nand U17052 (N_17052,N_16419,N_16613);
nor U17053 (N_17053,N_16488,N_16669);
and U17054 (N_17054,N_16799,N_16655);
nand U17055 (N_17055,N_16443,N_16689);
or U17056 (N_17056,N_16514,N_16656);
xnor U17057 (N_17057,N_16691,N_16744);
or U17058 (N_17058,N_16771,N_16521);
and U17059 (N_17059,N_16422,N_16491);
xor U17060 (N_17060,N_16701,N_16441);
xor U17061 (N_17061,N_16502,N_16521);
nor U17062 (N_17062,N_16407,N_16613);
and U17063 (N_17063,N_16521,N_16428);
or U17064 (N_17064,N_16537,N_16684);
or U17065 (N_17065,N_16446,N_16760);
nor U17066 (N_17066,N_16746,N_16457);
or U17067 (N_17067,N_16787,N_16573);
xnor U17068 (N_17068,N_16576,N_16664);
xnor U17069 (N_17069,N_16741,N_16667);
and U17070 (N_17070,N_16436,N_16547);
and U17071 (N_17071,N_16482,N_16669);
or U17072 (N_17072,N_16453,N_16581);
nand U17073 (N_17073,N_16488,N_16740);
and U17074 (N_17074,N_16759,N_16466);
nand U17075 (N_17075,N_16515,N_16435);
nor U17076 (N_17076,N_16706,N_16735);
xor U17077 (N_17077,N_16701,N_16605);
or U17078 (N_17078,N_16437,N_16542);
or U17079 (N_17079,N_16455,N_16644);
nand U17080 (N_17080,N_16664,N_16759);
and U17081 (N_17081,N_16653,N_16494);
and U17082 (N_17082,N_16631,N_16760);
or U17083 (N_17083,N_16648,N_16785);
and U17084 (N_17084,N_16729,N_16523);
or U17085 (N_17085,N_16719,N_16657);
or U17086 (N_17086,N_16627,N_16592);
nor U17087 (N_17087,N_16426,N_16554);
and U17088 (N_17088,N_16486,N_16716);
nand U17089 (N_17089,N_16577,N_16600);
or U17090 (N_17090,N_16701,N_16717);
or U17091 (N_17091,N_16690,N_16575);
nor U17092 (N_17092,N_16767,N_16732);
or U17093 (N_17093,N_16651,N_16625);
nor U17094 (N_17094,N_16687,N_16450);
xnor U17095 (N_17095,N_16677,N_16739);
nor U17096 (N_17096,N_16529,N_16407);
and U17097 (N_17097,N_16408,N_16487);
and U17098 (N_17098,N_16464,N_16791);
or U17099 (N_17099,N_16631,N_16679);
and U17100 (N_17100,N_16519,N_16650);
nor U17101 (N_17101,N_16591,N_16666);
xor U17102 (N_17102,N_16567,N_16698);
xor U17103 (N_17103,N_16730,N_16675);
and U17104 (N_17104,N_16694,N_16745);
and U17105 (N_17105,N_16560,N_16652);
or U17106 (N_17106,N_16754,N_16476);
nand U17107 (N_17107,N_16776,N_16618);
and U17108 (N_17108,N_16434,N_16475);
or U17109 (N_17109,N_16423,N_16689);
or U17110 (N_17110,N_16545,N_16732);
nand U17111 (N_17111,N_16479,N_16723);
or U17112 (N_17112,N_16510,N_16632);
and U17113 (N_17113,N_16599,N_16660);
xor U17114 (N_17114,N_16790,N_16450);
xor U17115 (N_17115,N_16756,N_16553);
nand U17116 (N_17116,N_16408,N_16532);
nand U17117 (N_17117,N_16594,N_16513);
or U17118 (N_17118,N_16472,N_16624);
and U17119 (N_17119,N_16474,N_16663);
nor U17120 (N_17120,N_16557,N_16602);
nand U17121 (N_17121,N_16402,N_16653);
and U17122 (N_17122,N_16791,N_16530);
nor U17123 (N_17123,N_16582,N_16463);
and U17124 (N_17124,N_16485,N_16535);
xnor U17125 (N_17125,N_16791,N_16402);
or U17126 (N_17126,N_16697,N_16502);
and U17127 (N_17127,N_16602,N_16430);
xor U17128 (N_17128,N_16431,N_16407);
or U17129 (N_17129,N_16469,N_16673);
xnor U17130 (N_17130,N_16546,N_16446);
and U17131 (N_17131,N_16593,N_16418);
and U17132 (N_17132,N_16672,N_16634);
or U17133 (N_17133,N_16769,N_16564);
and U17134 (N_17134,N_16554,N_16434);
xnor U17135 (N_17135,N_16729,N_16518);
and U17136 (N_17136,N_16527,N_16765);
and U17137 (N_17137,N_16669,N_16558);
nand U17138 (N_17138,N_16794,N_16483);
and U17139 (N_17139,N_16465,N_16597);
nor U17140 (N_17140,N_16657,N_16625);
xnor U17141 (N_17141,N_16544,N_16580);
or U17142 (N_17142,N_16406,N_16752);
and U17143 (N_17143,N_16644,N_16439);
or U17144 (N_17144,N_16525,N_16677);
or U17145 (N_17145,N_16474,N_16555);
xor U17146 (N_17146,N_16450,N_16772);
and U17147 (N_17147,N_16559,N_16752);
and U17148 (N_17148,N_16402,N_16454);
and U17149 (N_17149,N_16574,N_16407);
nand U17150 (N_17150,N_16788,N_16669);
xnor U17151 (N_17151,N_16797,N_16633);
and U17152 (N_17152,N_16689,N_16714);
nand U17153 (N_17153,N_16756,N_16647);
and U17154 (N_17154,N_16426,N_16679);
nand U17155 (N_17155,N_16495,N_16561);
xnor U17156 (N_17156,N_16631,N_16589);
nor U17157 (N_17157,N_16682,N_16617);
nand U17158 (N_17158,N_16771,N_16787);
nand U17159 (N_17159,N_16705,N_16404);
xnor U17160 (N_17160,N_16491,N_16705);
nor U17161 (N_17161,N_16652,N_16740);
or U17162 (N_17162,N_16737,N_16558);
and U17163 (N_17163,N_16562,N_16638);
and U17164 (N_17164,N_16676,N_16498);
and U17165 (N_17165,N_16780,N_16523);
xor U17166 (N_17166,N_16715,N_16586);
nand U17167 (N_17167,N_16662,N_16446);
nor U17168 (N_17168,N_16488,N_16737);
and U17169 (N_17169,N_16562,N_16750);
or U17170 (N_17170,N_16731,N_16537);
nor U17171 (N_17171,N_16511,N_16647);
or U17172 (N_17172,N_16710,N_16586);
or U17173 (N_17173,N_16650,N_16402);
nand U17174 (N_17174,N_16627,N_16437);
or U17175 (N_17175,N_16629,N_16687);
nor U17176 (N_17176,N_16636,N_16619);
or U17177 (N_17177,N_16465,N_16752);
nand U17178 (N_17178,N_16678,N_16596);
nor U17179 (N_17179,N_16718,N_16501);
and U17180 (N_17180,N_16405,N_16650);
and U17181 (N_17181,N_16539,N_16644);
nand U17182 (N_17182,N_16611,N_16553);
and U17183 (N_17183,N_16622,N_16401);
nor U17184 (N_17184,N_16580,N_16618);
or U17185 (N_17185,N_16694,N_16585);
or U17186 (N_17186,N_16733,N_16665);
nor U17187 (N_17187,N_16782,N_16683);
and U17188 (N_17188,N_16604,N_16455);
xor U17189 (N_17189,N_16495,N_16579);
or U17190 (N_17190,N_16666,N_16500);
and U17191 (N_17191,N_16440,N_16564);
or U17192 (N_17192,N_16758,N_16503);
nor U17193 (N_17193,N_16494,N_16527);
and U17194 (N_17194,N_16667,N_16540);
and U17195 (N_17195,N_16407,N_16608);
or U17196 (N_17196,N_16600,N_16777);
xnor U17197 (N_17197,N_16643,N_16683);
xnor U17198 (N_17198,N_16559,N_16577);
xor U17199 (N_17199,N_16597,N_16500);
xnor U17200 (N_17200,N_17049,N_17123);
nand U17201 (N_17201,N_16855,N_16888);
nand U17202 (N_17202,N_16837,N_17189);
nand U17203 (N_17203,N_17036,N_17090);
xnor U17204 (N_17204,N_17060,N_17161);
xor U17205 (N_17205,N_16939,N_17001);
nor U17206 (N_17206,N_16988,N_16981);
xor U17207 (N_17207,N_17014,N_17163);
and U17208 (N_17208,N_16938,N_16989);
or U17209 (N_17209,N_16918,N_17113);
or U17210 (N_17210,N_17187,N_17127);
and U17211 (N_17211,N_17107,N_17000);
nand U17212 (N_17212,N_17009,N_16943);
or U17213 (N_17213,N_16917,N_17152);
or U17214 (N_17214,N_17028,N_16949);
or U17215 (N_17215,N_16993,N_17166);
xnor U17216 (N_17216,N_17063,N_17101);
or U17217 (N_17217,N_17160,N_16903);
and U17218 (N_17218,N_16894,N_17093);
or U17219 (N_17219,N_17013,N_17147);
nor U17220 (N_17220,N_16992,N_16986);
nor U17221 (N_17221,N_17156,N_16942);
xor U17222 (N_17222,N_16835,N_16915);
or U17223 (N_17223,N_17146,N_17135);
or U17224 (N_17224,N_17109,N_16996);
nand U17225 (N_17225,N_16991,N_17121);
and U17226 (N_17226,N_16818,N_16969);
and U17227 (N_17227,N_16919,N_17124);
nand U17228 (N_17228,N_17175,N_16862);
and U17229 (N_17229,N_16987,N_17106);
and U17230 (N_17230,N_17038,N_16847);
nor U17231 (N_17231,N_17142,N_16970);
nor U17232 (N_17232,N_17194,N_17172);
nor U17233 (N_17233,N_17035,N_17033);
xor U17234 (N_17234,N_17017,N_17164);
xnor U17235 (N_17235,N_16930,N_17149);
nor U17236 (N_17236,N_16931,N_16841);
nor U17237 (N_17237,N_17116,N_16832);
or U17238 (N_17238,N_17139,N_16901);
nand U17239 (N_17239,N_16833,N_17077);
xnor U17240 (N_17240,N_17057,N_17007);
nor U17241 (N_17241,N_16854,N_17074);
and U17242 (N_17242,N_17162,N_16946);
or U17243 (N_17243,N_16817,N_17064);
nand U17244 (N_17244,N_17171,N_17059);
nor U17245 (N_17245,N_16821,N_17183);
nor U17246 (N_17246,N_17006,N_17032);
nor U17247 (N_17247,N_17125,N_16829);
xor U17248 (N_17248,N_17176,N_16964);
or U17249 (N_17249,N_17119,N_17167);
and U17250 (N_17250,N_17177,N_17196);
and U17251 (N_17251,N_16904,N_16960);
or U17252 (N_17252,N_16913,N_16826);
nand U17253 (N_17253,N_16984,N_16911);
xnor U17254 (N_17254,N_17094,N_17058);
or U17255 (N_17255,N_16853,N_17184);
nor U17256 (N_17256,N_16838,N_17092);
nand U17257 (N_17257,N_16952,N_17165);
nor U17258 (N_17258,N_16924,N_16910);
nand U17259 (N_17259,N_16885,N_17054);
nand U17260 (N_17260,N_17132,N_17065);
xor U17261 (N_17261,N_16998,N_17078);
and U17262 (N_17262,N_17003,N_16807);
xnor U17263 (N_17263,N_16951,N_16929);
xnor U17264 (N_17264,N_17181,N_17055);
nor U17265 (N_17265,N_16805,N_16857);
nor U17266 (N_17266,N_16925,N_16831);
xor U17267 (N_17267,N_17042,N_16806);
nand U17268 (N_17268,N_16870,N_17131);
xnor U17269 (N_17269,N_16985,N_16965);
nand U17270 (N_17270,N_17004,N_16908);
and U17271 (N_17271,N_17070,N_16804);
and U17272 (N_17272,N_16900,N_16936);
nand U17273 (N_17273,N_16814,N_16926);
xor U17274 (N_17274,N_17072,N_17067);
xnor U17275 (N_17275,N_17129,N_17045);
nor U17276 (N_17276,N_16836,N_17041);
or U17277 (N_17277,N_17178,N_16916);
nor U17278 (N_17278,N_16852,N_17023);
and U17279 (N_17279,N_17144,N_17188);
or U17280 (N_17280,N_16834,N_16954);
xnor U17281 (N_17281,N_16809,N_17046);
nand U17282 (N_17282,N_17192,N_17170);
or U17283 (N_17283,N_17148,N_16874);
nor U17284 (N_17284,N_17044,N_16948);
nand U17285 (N_17285,N_16887,N_16890);
xnor U17286 (N_17286,N_16895,N_16978);
nand U17287 (N_17287,N_17140,N_17011);
nor U17288 (N_17288,N_17138,N_16893);
xnor U17289 (N_17289,N_17086,N_16827);
nand U17290 (N_17290,N_17020,N_17158);
xor U17291 (N_17291,N_16921,N_17111);
nand U17292 (N_17292,N_16845,N_16851);
nor U17293 (N_17293,N_17179,N_16859);
nor U17294 (N_17294,N_16802,N_16820);
and U17295 (N_17295,N_17019,N_16906);
nand U17296 (N_17296,N_17073,N_16933);
or U17297 (N_17297,N_17076,N_16977);
nand U17298 (N_17298,N_16897,N_17137);
nand U17299 (N_17299,N_16849,N_17145);
nor U17300 (N_17300,N_17002,N_17102);
and U17301 (N_17301,N_17141,N_17084);
nand U17302 (N_17302,N_17182,N_17199);
nand U17303 (N_17303,N_16990,N_17027);
nor U17304 (N_17304,N_17190,N_16958);
and U17305 (N_17305,N_16968,N_16879);
nor U17306 (N_17306,N_16994,N_17126);
nor U17307 (N_17307,N_17168,N_16881);
and U17308 (N_17308,N_17180,N_16914);
and U17309 (N_17309,N_17193,N_17155);
xnor U17310 (N_17310,N_17089,N_16982);
nor U17311 (N_17311,N_16875,N_17122);
nor U17312 (N_17312,N_17066,N_16896);
nand U17313 (N_17313,N_17030,N_17085);
and U17314 (N_17314,N_16825,N_17117);
and U17315 (N_17315,N_16898,N_16975);
and U17316 (N_17316,N_16962,N_17097);
xnor U17317 (N_17317,N_17191,N_16800);
nor U17318 (N_17318,N_16819,N_16997);
and U17319 (N_17319,N_16803,N_17143);
xor U17320 (N_17320,N_16844,N_17198);
and U17321 (N_17321,N_17025,N_16950);
or U17322 (N_17322,N_17088,N_17173);
and U17323 (N_17323,N_17134,N_17026);
xnor U17324 (N_17324,N_16983,N_17037);
or U17325 (N_17325,N_16877,N_17069);
or U17326 (N_17326,N_16876,N_16973);
and U17327 (N_17327,N_16909,N_16860);
or U17328 (N_17328,N_16922,N_16810);
nor U17329 (N_17329,N_16867,N_16892);
xor U17330 (N_17330,N_16808,N_16813);
nor U17331 (N_17331,N_17039,N_17010);
xnor U17332 (N_17332,N_17047,N_17112);
nor U17333 (N_17333,N_16999,N_16940);
nor U17334 (N_17334,N_17022,N_17108);
xor U17335 (N_17335,N_16882,N_16866);
and U17336 (N_17336,N_16966,N_17104);
xnor U17337 (N_17337,N_16883,N_16976);
and U17338 (N_17338,N_17082,N_16934);
or U17339 (N_17339,N_17015,N_17031);
and U17340 (N_17340,N_17133,N_16905);
xor U17341 (N_17341,N_17105,N_17005);
xor U17342 (N_17342,N_16873,N_16861);
xnor U17343 (N_17343,N_16932,N_17185);
nor U17344 (N_17344,N_16871,N_17195);
and U17345 (N_17345,N_17048,N_17056);
or U17346 (N_17346,N_17068,N_16801);
or U17347 (N_17347,N_16907,N_16972);
and U17348 (N_17348,N_16974,N_17029);
nor U17349 (N_17349,N_16995,N_17114);
xor U17350 (N_17350,N_16935,N_16945);
xor U17351 (N_17351,N_17062,N_17153);
or U17352 (N_17352,N_16912,N_17115);
nand U17353 (N_17353,N_17012,N_17040);
nand U17354 (N_17354,N_17087,N_16884);
and U17355 (N_17355,N_17120,N_16953);
and U17356 (N_17356,N_16865,N_17157);
xnor U17357 (N_17357,N_17150,N_16941);
nand U17358 (N_17358,N_17053,N_16944);
nor U17359 (N_17359,N_17016,N_17154);
or U17360 (N_17360,N_16823,N_16889);
and U17361 (N_17361,N_16878,N_17197);
nand U17362 (N_17362,N_16961,N_16843);
and U17363 (N_17363,N_17159,N_17080);
nand U17364 (N_17364,N_16868,N_16816);
nor U17365 (N_17365,N_16822,N_17008);
xnor U17366 (N_17366,N_17128,N_17043);
and U17367 (N_17367,N_17061,N_17130);
nand U17368 (N_17368,N_16956,N_16811);
xor U17369 (N_17369,N_17099,N_16971);
and U17370 (N_17370,N_16856,N_16850);
and U17371 (N_17371,N_16959,N_17095);
xnor U17372 (N_17372,N_16864,N_16920);
or U17373 (N_17373,N_17110,N_16872);
or U17374 (N_17374,N_16886,N_17034);
nand U17375 (N_17375,N_16891,N_16880);
or U17376 (N_17376,N_17079,N_16824);
xnor U17377 (N_17377,N_16846,N_16858);
nor U17378 (N_17378,N_16967,N_16828);
and U17379 (N_17379,N_16980,N_16863);
nand U17380 (N_17380,N_17174,N_17169);
nand U17381 (N_17381,N_17081,N_17098);
nor U17382 (N_17382,N_16899,N_17071);
nand U17383 (N_17383,N_17151,N_17118);
and U17384 (N_17384,N_17051,N_17075);
xnor U17385 (N_17385,N_16848,N_16955);
xor U17386 (N_17386,N_16842,N_16830);
nor U17387 (N_17387,N_17083,N_16840);
or U17388 (N_17388,N_17096,N_16957);
nor U17389 (N_17389,N_16963,N_17052);
nand U17390 (N_17390,N_16902,N_17186);
or U17391 (N_17391,N_16947,N_16923);
or U17392 (N_17392,N_16927,N_16869);
or U17393 (N_17393,N_17100,N_17021);
xnor U17394 (N_17394,N_17136,N_16937);
nand U17395 (N_17395,N_16979,N_17050);
xnor U17396 (N_17396,N_16839,N_16815);
nand U17397 (N_17397,N_16812,N_17018);
xor U17398 (N_17398,N_17024,N_16928);
nand U17399 (N_17399,N_17091,N_17103);
and U17400 (N_17400,N_16970,N_17162);
or U17401 (N_17401,N_17014,N_16853);
nand U17402 (N_17402,N_17174,N_17135);
nand U17403 (N_17403,N_16926,N_16930);
xnor U17404 (N_17404,N_16891,N_17182);
nand U17405 (N_17405,N_17053,N_17039);
or U17406 (N_17406,N_16978,N_16822);
nor U17407 (N_17407,N_17195,N_17191);
nand U17408 (N_17408,N_17054,N_16931);
or U17409 (N_17409,N_17009,N_17160);
nand U17410 (N_17410,N_16820,N_17121);
or U17411 (N_17411,N_17158,N_16945);
xor U17412 (N_17412,N_16813,N_17046);
nor U17413 (N_17413,N_17046,N_17048);
and U17414 (N_17414,N_16905,N_17022);
or U17415 (N_17415,N_17097,N_16813);
nor U17416 (N_17416,N_17188,N_17076);
nand U17417 (N_17417,N_17123,N_16958);
and U17418 (N_17418,N_17041,N_17012);
nand U17419 (N_17419,N_17134,N_17124);
xor U17420 (N_17420,N_17190,N_17068);
xor U17421 (N_17421,N_17188,N_16861);
nand U17422 (N_17422,N_17173,N_16867);
xor U17423 (N_17423,N_16870,N_16833);
nand U17424 (N_17424,N_16890,N_16800);
and U17425 (N_17425,N_17138,N_17022);
or U17426 (N_17426,N_16891,N_17006);
nand U17427 (N_17427,N_16995,N_17075);
xor U17428 (N_17428,N_16991,N_16885);
nand U17429 (N_17429,N_16881,N_17127);
and U17430 (N_17430,N_17134,N_16881);
nor U17431 (N_17431,N_17191,N_17045);
and U17432 (N_17432,N_16883,N_16879);
nand U17433 (N_17433,N_17141,N_17058);
and U17434 (N_17434,N_17134,N_17127);
xnor U17435 (N_17435,N_16871,N_16956);
or U17436 (N_17436,N_17064,N_16878);
nand U17437 (N_17437,N_17121,N_16997);
nor U17438 (N_17438,N_17058,N_16835);
and U17439 (N_17439,N_16885,N_17112);
xnor U17440 (N_17440,N_16806,N_17004);
or U17441 (N_17441,N_17065,N_16854);
nor U17442 (N_17442,N_17041,N_16980);
and U17443 (N_17443,N_17104,N_17143);
nor U17444 (N_17444,N_17112,N_17059);
and U17445 (N_17445,N_16963,N_17039);
or U17446 (N_17446,N_17004,N_16854);
nor U17447 (N_17447,N_16913,N_17075);
nor U17448 (N_17448,N_16841,N_17186);
nand U17449 (N_17449,N_16839,N_16951);
xnor U17450 (N_17450,N_17137,N_17100);
nor U17451 (N_17451,N_17135,N_17198);
nor U17452 (N_17452,N_16896,N_17014);
nor U17453 (N_17453,N_16850,N_17132);
nand U17454 (N_17454,N_17045,N_17107);
and U17455 (N_17455,N_16903,N_17056);
nor U17456 (N_17456,N_16823,N_16816);
nor U17457 (N_17457,N_16808,N_16925);
or U17458 (N_17458,N_17058,N_17029);
and U17459 (N_17459,N_17110,N_17160);
or U17460 (N_17460,N_17052,N_17174);
nand U17461 (N_17461,N_17170,N_17033);
or U17462 (N_17462,N_17133,N_17098);
xor U17463 (N_17463,N_17093,N_16972);
or U17464 (N_17464,N_17188,N_16937);
and U17465 (N_17465,N_17077,N_17107);
nor U17466 (N_17466,N_17026,N_16880);
or U17467 (N_17467,N_16825,N_17147);
nand U17468 (N_17468,N_17001,N_17099);
xnor U17469 (N_17469,N_17032,N_17056);
nand U17470 (N_17470,N_17119,N_17090);
or U17471 (N_17471,N_16903,N_16873);
and U17472 (N_17472,N_17026,N_16828);
nor U17473 (N_17473,N_16869,N_16998);
or U17474 (N_17474,N_17094,N_16898);
nor U17475 (N_17475,N_16939,N_17035);
and U17476 (N_17476,N_16815,N_17196);
or U17477 (N_17477,N_16807,N_16838);
or U17478 (N_17478,N_16948,N_17060);
xor U17479 (N_17479,N_17074,N_16925);
nor U17480 (N_17480,N_16928,N_17048);
and U17481 (N_17481,N_16940,N_16809);
xor U17482 (N_17482,N_17010,N_17069);
or U17483 (N_17483,N_16835,N_16811);
and U17484 (N_17484,N_17106,N_16840);
xnor U17485 (N_17485,N_17178,N_17067);
and U17486 (N_17486,N_17075,N_17053);
and U17487 (N_17487,N_17187,N_17044);
nor U17488 (N_17488,N_16834,N_17197);
xnor U17489 (N_17489,N_17176,N_16880);
and U17490 (N_17490,N_16992,N_16912);
nand U17491 (N_17491,N_17035,N_17114);
or U17492 (N_17492,N_17032,N_17071);
nand U17493 (N_17493,N_16994,N_16821);
nor U17494 (N_17494,N_16886,N_17185);
and U17495 (N_17495,N_17183,N_16950);
or U17496 (N_17496,N_17054,N_17138);
xor U17497 (N_17497,N_16931,N_17003);
nor U17498 (N_17498,N_16970,N_16918);
nand U17499 (N_17499,N_16971,N_17173);
nand U17500 (N_17500,N_16903,N_16926);
xnor U17501 (N_17501,N_16816,N_17167);
xor U17502 (N_17502,N_16938,N_17108);
and U17503 (N_17503,N_17075,N_16908);
or U17504 (N_17504,N_17158,N_16966);
and U17505 (N_17505,N_17161,N_16912);
or U17506 (N_17506,N_16895,N_16852);
nor U17507 (N_17507,N_16812,N_17086);
or U17508 (N_17508,N_17148,N_16842);
and U17509 (N_17509,N_17180,N_16806);
nor U17510 (N_17510,N_17077,N_16938);
or U17511 (N_17511,N_16922,N_17123);
nor U17512 (N_17512,N_17100,N_16982);
or U17513 (N_17513,N_17004,N_16871);
or U17514 (N_17514,N_16856,N_17076);
and U17515 (N_17515,N_16907,N_16983);
xor U17516 (N_17516,N_17010,N_17063);
and U17517 (N_17517,N_16906,N_17047);
and U17518 (N_17518,N_16992,N_17177);
and U17519 (N_17519,N_16957,N_17152);
and U17520 (N_17520,N_16990,N_16954);
xnor U17521 (N_17521,N_16987,N_17054);
and U17522 (N_17522,N_17139,N_17157);
xor U17523 (N_17523,N_16812,N_17098);
or U17524 (N_17524,N_17084,N_17130);
nand U17525 (N_17525,N_16926,N_17073);
nand U17526 (N_17526,N_16860,N_17185);
and U17527 (N_17527,N_16891,N_16860);
nor U17528 (N_17528,N_16972,N_17184);
xor U17529 (N_17529,N_16916,N_16805);
or U17530 (N_17530,N_16801,N_16966);
or U17531 (N_17531,N_16955,N_17175);
xor U17532 (N_17532,N_16895,N_16938);
or U17533 (N_17533,N_17182,N_17006);
and U17534 (N_17534,N_17114,N_16877);
and U17535 (N_17535,N_16835,N_16947);
nand U17536 (N_17536,N_17008,N_17026);
nor U17537 (N_17537,N_16855,N_16862);
or U17538 (N_17538,N_16946,N_17176);
nor U17539 (N_17539,N_17049,N_16889);
or U17540 (N_17540,N_16877,N_16864);
nand U17541 (N_17541,N_16989,N_17167);
nand U17542 (N_17542,N_16945,N_16908);
and U17543 (N_17543,N_17161,N_17031);
nor U17544 (N_17544,N_17089,N_17183);
or U17545 (N_17545,N_17130,N_16984);
and U17546 (N_17546,N_16832,N_16807);
or U17547 (N_17547,N_17147,N_16887);
and U17548 (N_17548,N_17177,N_17099);
nor U17549 (N_17549,N_17058,N_16860);
xnor U17550 (N_17550,N_16887,N_17099);
nor U17551 (N_17551,N_16821,N_16953);
or U17552 (N_17552,N_16948,N_16898);
and U17553 (N_17553,N_17024,N_16953);
nor U17554 (N_17554,N_16838,N_17139);
xnor U17555 (N_17555,N_17008,N_16856);
xnor U17556 (N_17556,N_17157,N_16895);
nand U17557 (N_17557,N_17081,N_17096);
nand U17558 (N_17558,N_17036,N_17075);
nand U17559 (N_17559,N_16968,N_17000);
nand U17560 (N_17560,N_16989,N_16939);
or U17561 (N_17561,N_16957,N_17194);
nand U17562 (N_17562,N_17130,N_16819);
nand U17563 (N_17563,N_16935,N_16871);
nand U17564 (N_17564,N_16856,N_16980);
and U17565 (N_17565,N_16854,N_16920);
or U17566 (N_17566,N_16951,N_16856);
and U17567 (N_17567,N_16879,N_17155);
and U17568 (N_17568,N_16830,N_16990);
nor U17569 (N_17569,N_17198,N_17161);
and U17570 (N_17570,N_16951,N_17063);
or U17571 (N_17571,N_17116,N_17009);
nand U17572 (N_17572,N_17155,N_17096);
or U17573 (N_17573,N_16924,N_16974);
nand U17574 (N_17574,N_17172,N_16899);
xnor U17575 (N_17575,N_16829,N_17066);
nand U17576 (N_17576,N_17067,N_16846);
and U17577 (N_17577,N_17046,N_17007);
xnor U17578 (N_17578,N_16940,N_16951);
or U17579 (N_17579,N_17165,N_17017);
xor U17580 (N_17580,N_16944,N_16953);
and U17581 (N_17581,N_16808,N_16918);
and U17582 (N_17582,N_16874,N_17022);
nor U17583 (N_17583,N_16862,N_16941);
and U17584 (N_17584,N_17031,N_17080);
nand U17585 (N_17585,N_17078,N_17161);
xor U17586 (N_17586,N_17025,N_16801);
and U17587 (N_17587,N_16803,N_17137);
nor U17588 (N_17588,N_16879,N_16859);
nor U17589 (N_17589,N_16867,N_17012);
or U17590 (N_17590,N_16897,N_16810);
nor U17591 (N_17591,N_17025,N_16901);
and U17592 (N_17592,N_16939,N_17191);
xor U17593 (N_17593,N_17156,N_17063);
nor U17594 (N_17594,N_16939,N_16953);
nor U17595 (N_17595,N_17126,N_16873);
or U17596 (N_17596,N_16932,N_17037);
nor U17597 (N_17597,N_17156,N_17132);
xnor U17598 (N_17598,N_17002,N_16993);
nor U17599 (N_17599,N_16861,N_16921);
xnor U17600 (N_17600,N_17576,N_17445);
or U17601 (N_17601,N_17587,N_17297);
or U17602 (N_17602,N_17301,N_17333);
and U17603 (N_17603,N_17397,N_17219);
or U17604 (N_17604,N_17457,N_17235);
or U17605 (N_17605,N_17415,N_17325);
xnor U17606 (N_17606,N_17409,N_17387);
or U17607 (N_17607,N_17341,N_17550);
or U17608 (N_17608,N_17476,N_17386);
xnor U17609 (N_17609,N_17347,N_17281);
nand U17610 (N_17610,N_17444,N_17303);
nor U17611 (N_17611,N_17588,N_17460);
and U17612 (N_17612,N_17299,N_17533);
nand U17613 (N_17613,N_17215,N_17529);
or U17614 (N_17614,N_17352,N_17450);
nor U17615 (N_17615,N_17406,N_17586);
xnor U17616 (N_17616,N_17288,N_17481);
and U17617 (N_17617,N_17443,N_17575);
and U17618 (N_17618,N_17572,N_17551);
nand U17619 (N_17619,N_17338,N_17535);
xnor U17620 (N_17620,N_17280,N_17374);
nor U17621 (N_17621,N_17417,N_17350);
or U17622 (N_17622,N_17380,N_17391);
and U17623 (N_17623,N_17218,N_17569);
nor U17624 (N_17624,N_17354,N_17423);
nand U17625 (N_17625,N_17359,N_17238);
nor U17626 (N_17626,N_17453,N_17441);
xor U17627 (N_17627,N_17237,N_17547);
nor U17628 (N_17628,N_17577,N_17536);
nand U17629 (N_17629,N_17447,N_17385);
nand U17630 (N_17630,N_17532,N_17541);
or U17631 (N_17631,N_17442,N_17309);
and U17632 (N_17632,N_17567,N_17452);
or U17633 (N_17633,N_17228,N_17468);
or U17634 (N_17634,N_17383,N_17257);
and U17635 (N_17635,N_17434,N_17498);
or U17636 (N_17636,N_17505,N_17201);
and U17637 (N_17637,N_17462,N_17310);
and U17638 (N_17638,N_17418,N_17390);
xnor U17639 (N_17639,N_17360,N_17488);
nor U17640 (N_17640,N_17348,N_17363);
xnor U17641 (N_17641,N_17477,N_17455);
xor U17642 (N_17642,N_17479,N_17224);
nor U17643 (N_17643,N_17540,N_17463);
xnor U17644 (N_17644,N_17419,N_17272);
or U17645 (N_17645,N_17290,N_17332);
and U17646 (N_17646,N_17340,N_17521);
and U17647 (N_17647,N_17568,N_17578);
nor U17648 (N_17648,N_17292,N_17519);
nand U17649 (N_17649,N_17379,N_17208);
or U17650 (N_17650,N_17286,N_17355);
nand U17651 (N_17651,N_17400,N_17432);
or U17652 (N_17652,N_17508,N_17207);
nor U17653 (N_17653,N_17261,N_17405);
and U17654 (N_17654,N_17378,N_17456);
and U17655 (N_17655,N_17459,N_17315);
xor U17656 (N_17656,N_17525,N_17407);
nand U17657 (N_17657,N_17253,N_17546);
and U17658 (N_17658,N_17252,N_17230);
xor U17659 (N_17659,N_17205,N_17414);
nor U17660 (N_17660,N_17200,N_17268);
nor U17661 (N_17661,N_17236,N_17499);
nor U17662 (N_17662,N_17279,N_17322);
nand U17663 (N_17663,N_17507,N_17313);
and U17664 (N_17664,N_17538,N_17269);
nor U17665 (N_17665,N_17283,N_17307);
and U17666 (N_17666,N_17579,N_17502);
or U17667 (N_17667,N_17544,N_17573);
xnor U17668 (N_17668,N_17597,N_17312);
xnor U17669 (N_17669,N_17308,N_17509);
nor U17670 (N_17670,N_17306,N_17356);
nand U17671 (N_17671,N_17361,N_17248);
or U17672 (N_17672,N_17470,N_17574);
and U17673 (N_17673,N_17478,N_17204);
and U17674 (N_17674,N_17480,N_17277);
nor U17675 (N_17675,N_17593,N_17467);
nor U17676 (N_17676,N_17223,N_17506);
xnor U17677 (N_17677,N_17559,N_17486);
nor U17678 (N_17678,N_17446,N_17565);
nor U17679 (N_17679,N_17398,N_17513);
nor U17680 (N_17680,N_17203,N_17585);
nor U17681 (N_17681,N_17458,N_17330);
nor U17682 (N_17682,N_17430,N_17489);
nand U17683 (N_17683,N_17394,N_17275);
or U17684 (N_17684,N_17410,N_17284);
xor U17685 (N_17685,N_17485,N_17264);
nand U17686 (N_17686,N_17493,N_17501);
nand U17687 (N_17687,N_17583,N_17490);
or U17688 (N_17688,N_17426,N_17367);
or U17689 (N_17689,N_17466,N_17598);
or U17690 (N_17690,N_17554,N_17305);
nand U17691 (N_17691,N_17395,N_17265);
nand U17692 (N_17692,N_17263,N_17451);
and U17693 (N_17693,N_17371,N_17475);
nor U17694 (N_17694,N_17548,N_17590);
or U17695 (N_17695,N_17384,N_17411);
and U17696 (N_17696,N_17408,N_17300);
nand U17697 (N_17697,N_17549,N_17461);
xnor U17698 (N_17698,N_17302,N_17589);
xor U17699 (N_17699,N_17524,N_17247);
xnor U17700 (N_17700,N_17229,N_17249);
nor U17701 (N_17701,N_17210,N_17241);
xor U17702 (N_17702,N_17436,N_17316);
or U17703 (N_17703,N_17329,N_17472);
nand U17704 (N_17704,N_17366,N_17388);
nand U17705 (N_17705,N_17560,N_17404);
nor U17706 (N_17706,N_17471,N_17267);
or U17707 (N_17707,N_17328,N_17276);
xor U17708 (N_17708,N_17530,N_17331);
or U17709 (N_17709,N_17421,N_17433);
nand U17710 (N_17710,N_17562,N_17339);
nor U17711 (N_17711,N_17357,N_17571);
or U17712 (N_17712,N_17424,N_17527);
nand U17713 (N_17713,N_17317,N_17537);
nand U17714 (N_17714,N_17542,N_17254);
nor U17715 (N_17715,N_17381,N_17209);
nand U17716 (N_17716,N_17496,N_17311);
xor U17717 (N_17717,N_17222,N_17427);
nand U17718 (N_17718,N_17438,N_17491);
nor U17719 (N_17719,N_17517,N_17595);
and U17720 (N_17720,N_17246,N_17344);
nand U17721 (N_17721,N_17429,N_17227);
and U17722 (N_17722,N_17392,N_17484);
nand U17723 (N_17723,N_17522,N_17351);
or U17724 (N_17724,N_17528,N_17258);
nand U17725 (N_17725,N_17564,N_17212);
or U17726 (N_17726,N_17206,N_17375);
xnor U17727 (N_17727,N_17543,N_17555);
xnor U17728 (N_17728,N_17231,N_17233);
xnor U17729 (N_17729,N_17566,N_17428);
and U17730 (N_17730,N_17483,N_17250);
and U17731 (N_17731,N_17435,N_17345);
or U17732 (N_17732,N_17323,N_17294);
xnor U17733 (N_17733,N_17422,N_17582);
or U17734 (N_17734,N_17262,N_17511);
nand U17735 (N_17735,N_17495,N_17278);
and U17736 (N_17736,N_17291,N_17221);
xor U17737 (N_17737,N_17469,N_17596);
nand U17738 (N_17738,N_17557,N_17296);
and U17739 (N_17739,N_17592,N_17474);
or U17740 (N_17740,N_17287,N_17396);
nor U17741 (N_17741,N_17599,N_17211);
xor U17742 (N_17742,N_17362,N_17217);
or U17743 (N_17743,N_17584,N_17304);
or U17744 (N_17744,N_17244,N_17449);
nor U17745 (N_17745,N_17413,N_17370);
xnor U17746 (N_17746,N_17558,N_17318);
and U17747 (N_17747,N_17349,N_17274);
nand U17748 (N_17748,N_17497,N_17526);
nor U17749 (N_17749,N_17465,N_17232);
and U17750 (N_17750,N_17270,N_17520);
nor U17751 (N_17751,N_17285,N_17591);
nor U17752 (N_17752,N_17448,N_17372);
xnor U17753 (N_17753,N_17342,N_17260);
nand U17754 (N_17754,N_17334,N_17266);
or U17755 (N_17755,N_17389,N_17214);
nor U17756 (N_17756,N_17382,N_17225);
nor U17757 (N_17757,N_17298,N_17531);
xor U17758 (N_17758,N_17282,N_17202);
and U17759 (N_17759,N_17369,N_17234);
or U17760 (N_17760,N_17368,N_17243);
nand U17761 (N_17761,N_17464,N_17220);
nor U17762 (N_17762,N_17539,N_17420);
nand U17763 (N_17763,N_17346,N_17255);
nor U17764 (N_17764,N_17293,N_17515);
nor U17765 (N_17765,N_17273,N_17320);
and U17766 (N_17766,N_17516,N_17570);
and U17767 (N_17767,N_17343,N_17364);
nor U17768 (N_17768,N_17552,N_17416);
nor U17769 (N_17769,N_17337,N_17271);
or U17770 (N_17770,N_17440,N_17454);
nor U17771 (N_17771,N_17437,N_17377);
nor U17772 (N_17772,N_17245,N_17431);
or U17773 (N_17773,N_17376,N_17594);
and U17774 (N_17774,N_17503,N_17494);
or U17775 (N_17775,N_17399,N_17556);
nand U17776 (N_17776,N_17239,N_17393);
and U17777 (N_17777,N_17514,N_17327);
nand U17778 (N_17778,N_17326,N_17259);
and U17779 (N_17779,N_17226,N_17500);
xor U17780 (N_17780,N_17295,N_17581);
or U17781 (N_17781,N_17353,N_17358);
nor U17782 (N_17782,N_17289,N_17335);
xnor U17783 (N_17783,N_17373,N_17482);
or U17784 (N_17784,N_17473,N_17545);
nor U17785 (N_17785,N_17321,N_17401);
or U17786 (N_17786,N_17518,N_17523);
and U17787 (N_17787,N_17240,N_17487);
or U17788 (N_17788,N_17510,N_17439);
nand U17789 (N_17789,N_17251,N_17365);
nand U17790 (N_17790,N_17504,N_17213);
nor U17791 (N_17791,N_17314,N_17402);
and U17792 (N_17792,N_17319,N_17492);
or U17793 (N_17793,N_17336,N_17534);
nor U17794 (N_17794,N_17580,N_17242);
nand U17795 (N_17795,N_17561,N_17324);
nand U17796 (N_17796,N_17425,N_17256);
or U17797 (N_17797,N_17553,N_17403);
nand U17798 (N_17798,N_17563,N_17512);
nor U17799 (N_17799,N_17216,N_17412);
xnor U17800 (N_17800,N_17305,N_17250);
nand U17801 (N_17801,N_17202,N_17488);
or U17802 (N_17802,N_17393,N_17496);
nand U17803 (N_17803,N_17448,N_17340);
xor U17804 (N_17804,N_17232,N_17261);
nor U17805 (N_17805,N_17444,N_17464);
or U17806 (N_17806,N_17556,N_17559);
xor U17807 (N_17807,N_17391,N_17337);
nor U17808 (N_17808,N_17473,N_17430);
nand U17809 (N_17809,N_17588,N_17207);
nor U17810 (N_17810,N_17241,N_17269);
or U17811 (N_17811,N_17442,N_17509);
nor U17812 (N_17812,N_17564,N_17385);
and U17813 (N_17813,N_17307,N_17424);
and U17814 (N_17814,N_17546,N_17458);
nand U17815 (N_17815,N_17214,N_17413);
nor U17816 (N_17816,N_17355,N_17589);
nand U17817 (N_17817,N_17301,N_17208);
nor U17818 (N_17818,N_17550,N_17417);
xor U17819 (N_17819,N_17451,N_17577);
xnor U17820 (N_17820,N_17468,N_17485);
or U17821 (N_17821,N_17291,N_17594);
or U17822 (N_17822,N_17317,N_17360);
or U17823 (N_17823,N_17455,N_17254);
xor U17824 (N_17824,N_17228,N_17281);
and U17825 (N_17825,N_17209,N_17238);
xnor U17826 (N_17826,N_17294,N_17436);
xor U17827 (N_17827,N_17227,N_17370);
nand U17828 (N_17828,N_17491,N_17347);
and U17829 (N_17829,N_17435,N_17289);
and U17830 (N_17830,N_17206,N_17472);
nand U17831 (N_17831,N_17443,N_17392);
and U17832 (N_17832,N_17366,N_17202);
nand U17833 (N_17833,N_17543,N_17424);
nor U17834 (N_17834,N_17394,N_17363);
nor U17835 (N_17835,N_17333,N_17502);
and U17836 (N_17836,N_17400,N_17467);
or U17837 (N_17837,N_17515,N_17414);
nor U17838 (N_17838,N_17262,N_17410);
or U17839 (N_17839,N_17284,N_17235);
nand U17840 (N_17840,N_17483,N_17321);
xor U17841 (N_17841,N_17500,N_17585);
nand U17842 (N_17842,N_17453,N_17212);
xnor U17843 (N_17843,N_17214,N_17366);
and U17844 (N_17844,N_17523,N_17317);
or U17845 (N_17845,N_17223,N_17374);
nand U17846 (N_17846,N_17548,N_17521);
nor U17847 (N_17847,N_17313,N_17555);
xor U17848 (N_17848,N_17264,N_17353);
or U17849 (N_17849,N_17342,N_17332);
xor U17850 (N_17850,N_17293,N_17505);
nand U17851 (N_17851,N_17579,N_17234);
or U17852 (N_17852,N_17379,N_17461);
nand U17853 (N_17853,N_17565,N_17466);
xnor U17854 (N_17854,N_17338,N_17246);
nor U17855 (N_17855,N_17346,N_17510);
nor U17856 (N_17856,N_17529,N_17297);
and U17857 (N_17857,N_17381,N_17360);
nor U17858 (N_17858,N_17505,N_17532);
or U17859 (N_17859,N_17373,N_17376);
xnor U17860 (N_17860,N_17302,N_17408);
nor U17861 (N_17861,N_17252,N_17207);
or U17862 (N_17862,N_17518,N_17208);
xor U17863 (N_17863,N_17439,N_17435);
xor U17864 (N_17864,N_17580,N_17454);
xor U17865 (N_17865,N_17301,N_17212);
xnor U17866 (N_17866,N_17291,N_17262);
or U17867 (N_17867,N_17470,N_17530);
or U17868 (N_17868,N_17212,N_17238);
xnor U17869 (N_17869,N_17549,N_17210);
xnor U17870 (N_17870,N_17551,N_17374);
or U17871 (N_17871,N_17456,N_17259);
xor U17872 (N_17872,N_17382,N_17462);
or U17873 (N_17873,N_17359,N_17251);
nand U17874 (N_17874,N_17466,N_17407);
nor U17875 (N_17875,N_17500,N_17535);
nand U17876 (N_17876,N_17227,N_17307);
nor U17877 (N_17877,N_17396,N_17494);
xor U17878 (N_17878,N_17426,N_17589);
xor U17879 (N_17879,N_17321,N_17585);
xor U17880 (N_17880,N_17449,N_17590);
or U17881 (N_17881,N_17225,N_17588);
and U17882 (N_17882,N_17346,N_17321);
or U17883 (N_17883,N_17337,N_17468);
nor U17884 (N_17884,N_17319,N_17229);
nor U17885 (N_17885,N_17322,N_17325);
or U17886 (N_17886,N_17388,N_17243);
and U17887 (N_17887,N_17288,N_17422);
xnor U17888 (N_17888,N_17254,N_17319);
nand U17889 (N_17889,N_17351,N_17260);
nor U17890 (N_17890,N_17282,N_17558);
and U17891 (N_17891,N_17358,N_17465);
nor U17892 (N_17892,N_17294,N_17242);
nand U17893 (N_17893,N_17420,N_17436);
xnor U17894 (N_17894,N_17356,N_17532);
nand U17895 (N_17895,N_17386,N_17499);
nand U17896 (N_17896,N_17311,N_17465);
and U17897 (N_17897,N_17555,N_17539);
nor U17898 (N_17898,N_17399,N_17563);
nand U17899 (N_17899,N_17386,N_17401);
or U17900 (N_17900,N_17361,N_17497);
xor U17901 (N_17901,N_17453,N_17552);
or U17902 (N_17902,N_17247,N_17418);
xor U17903 (N_17903,N_17291,N_17280);
or U17904 (N_17904,N_17390,N_17284);
nand U17905 (N_17905,N_17542,N_17591);
xor U17906 (N_17906,N_17260,N_17441);
nor U17907 (N_17907,N_17210,N_17304);
xnor U17908 (N_17908,N_17302,N_17384);
nand U17909 (N_17909,N_17230,N_17504);
nor U17910 (N_17910,N_17380,N_17546);
nand U17911 (N_17911,N_17502,N_17568);
nor U17912 (N_17912,N_17329,N_17301);
nor U17913 (N_17913,N_17314,N_17347);
nand U17914 (N_17914,N_17472,N_17514);
xor U17915 (N_17915,N_17502,N_17265);
xor U17916 (N_17916,N_17451,N_17541);
and U17917 (N_17917,N_17270,N_17482);
and U17918 (N_17918,N_17522,N_17217);
or U17919 (N_17919,N_17427,N_17541);
and U17920 (N_17920,N_17293,N_17232);
and U17921 (N_17921,N_17404,N_17515);
nor U17922 (N_17922,N_17454,N_17547);
and U17923 (N_17923,N_17586,N_17523);
nor U17924 (N_17924,N_17424,N_17299);
and U17925 (N_17925,N_17444,N_17517);
and U17926 (N_17926,N_17548,N_17597);
or U17927 (N_17927,N_17419,N_17568);
or U17928 (N_17928,N_17559,N_17492);
and U17929 (N_17929,N_17383,N_17426);
or U17930 (N_17930,N_17249,N_17571);
nor U17931 (N_17931,N_17401,N_17443);
xnor U17932 (N_17932,N_17365,N_17422);
or U17933 (N_17933,N_17481,N_17423);
and U17934 (N_17934,N_17244,N_17502);
or U17935 (N_17935,N_17240,N_17498);
nand U17936 (N_17936,N_17259,N_17591);
or U17937 (N_17937,N_17532,N_17226);
xor U17938 (N_17938,N_17505,N_17316);
nor U17939 (N_17939,N_17595,N_17578);
xnor U17940 (N_17940,N_17419,N_17323);
or U17941 (N_17941,N_17387,N_17425);
nand U17942 (N_17942,N_17432,N_17391);
nand U17943 (N_17943,N_17515,N_17287);
or U17944 (N_17944,N_17375,N_17353);
nor U17945 (N_17945,N_17260,N_17408);
xnor U17946 (N_17946,N_17357,N_17499);
xnor U17947 (N_17947,N_17484,N_17218);
nor U17948 (N_17948,N_17309,N_17250);
nor U17949 (N_17949,N_17547,N_17311);
xor U17950 (N_17950,N_17576,N_17421);
and U17951 (N_17951,N_17367,N_17498);
nor U17952 (N_17952,N_17589,N_17263);
and U17953 (N_17953,N_17215,N_17267);
or U17954 (N_17954,N_17401,N_17414);
nor U17955 (N_17955,N_17588,N_17379);
nor U17956 (N_17956,N_17335,N_17552);
xor U17957 (N_17957,N_17346,N_17377);
xor U17958 (N_17958,N_17300,N_17271);
xnor U17959 (N_17959,N_17267,N_17351);
or U17960 (N_17960,N_17590,N_17567);
and U17961 (N_17961,N_17479,N_17524);
and U17962 (N_17962,N_17595,N_17540);
or U17963 (N_17963,N_17515,N_17373);
and U17964 (N_17964,N_17546,N_17550);
or U17965 (N_17965,N_17406,N_17426);
or U17966 (N_17966,N_17507,N_17462);
or U17967 (N_17967,N_17315,N_17373);
nand U17968 (N_17968,N_17360,N_17322);
nor U17969 (N_17969,N_17500,N_17530);
or U17970 (N_17970,N_17465,N_17343);
xor U17971 (N_17971,N_17316,N_17585);
and U17972 (N_17972,N_17588,N_17368);
xnor U17973 (N_17973,N_17496,N_17499);
xnor U17974 (N_17974,N_17232,N_17480);
xnor U17975 (N_17975,N_17482,N_17395);
nor U17976 (N_17976,N_17277,N_17409);
nand U17977 (N_17977,N_17487,N_17257);
nand U17978 (N_17978,N_17362,N_17422);
and U17979 (N_17979,N_17543,N_17455);
or U17980 (N_17980,N_17325,N_17416);
nor U17981 (N_17981,N_17356,N_17401);
nand U17982 (N_17982,N_17563,N_17532);
nor U17983 (N_17983,N_17364,N_17223);
xnor U17984 (N_17984,N_17541,N_17294);
nand U17985 (N_17985,N_17560,N_17365);
or U17986 (N_17986,N_17200,N_17283);
nand U17987 (N_17987,N_17376,N_17474);
and U17988 (N_17988,N_17232,N_17264);
xnor U17989 (N_17989,N_17430,N_17388);
nor U17990 (N_17990,N_17205,N_17372);
nand U17991 (N_17991,N_17476,N_17290);
and U17992 (N_17992,N_17328,N_17418);
and U17993 (N_17993,N_17274,N_17511);
and U17994 (N_17994,N_17393,N_17412);
xnor U17995 (N_17995,N_17392,N_17510);
nand U17996 (N_17996,N_17591,N_17241);
and U17997 (N_17997,N_17466,N_17573);
nor U17998 (N_17998,N_17399,N_17221);
xnor U17999 (N_17999,N_17521,N_17221);
nand U18000 (N_18000,N_17956,N_17901);
or U18001 (N_18001,N_17715,N_17896);
and U18002 (N_18002,N_17740,N_17762);
nor U18003 (N_18003,N_17641,N_17951);
nand U18004 (N_18004,N_17710,N_17622);
and U18005 (N_18005,N_17849,N_17938);
or U18006 (N_18006,N_17820,N_17916);
xor U18007 (N_18007,N_17758,N_17795);
or U18008 (N_18008,N_17858,N_17685);
xor U18009 (N_18009,N_17825,N_17962);
nor U18010 (N_18010,N_17712,N_17805);
and U18011 (N_18011,N_17647,N_17929);
and U18012 (N_18012,N_17733,N_17888);
nor U18013 (N_18013,N_17871,N_17719);
xnor U18014 (N_18014,N_17934,N_17626);
nand U18015 (N_18015,N_17772,N_17989);
xor U18016 (N_18016,N_17753,N_17732);
and U18017 (N_18017,N_17664,N_17633);
nor U18018 (N_18018,N_17717,N_17637);
nand U18019 (N_18019,N_17774,N_17747);
or U18020 (N_18020,N_17998,N_17859);
and U18021 (N_18021,N_17670,N_17912);
and U18022 (N_18022,N_17668,N_17894);
and U18023 (N_18023,N_17699,N_17937);
xnor U18024 (N_18024,N_17639,N_17952);
or U18025 (N_18025,N_17659,N_17706);
nor U18026 (N_18026,N_17756,N_17707);
nand U18027 (N_18027,N_17605,N_17686);
nor U18028 (N_18028,N_17971,N_17614);
nor U18029 (N_18029,N_17864,N_17744);
and U18030 (N_18030,N_17680,N_17848);
nor U18031 (N_18031,N_17883,N_17746);
nand U18032 (N_18032,N_17988,N_17850);
or U18033 (N_18033,N_17797,N_17812);
or U18034 (N_18034,N_17767,N_17855);
xnor U18035 (N_18035,N_17972,N_17765);
and U18036 (N_18036,N_17970,N_17757);
or U18037 (N_18037,N_17914,N_17936);
and U18038 (N_18038,N_17611,N_17694);
xor U18039 (N_18039,N_17730,N_17763);
xnor U18040 (N_18040,N_17928,N_17727);
xnor U18041 (N_18041,N_17677,N_17766);
or U18042 (N_18042,N_17913,N_17983);
nand U18043 (N_18043,N_17806,N_17651);
nand U18044 (N_18044,N_17866,N_17803);
or U18045 (N_18045,N_17905,N_17689);
or U18046 (N_18046,N_17656,N_17910);
nor U18047 (N_18047,N_17985,N_17868);
and U18048 (N_18048,N_17721,N_17827);
xnor U18049 (N_18049,N_17926,N_17663);
and U18050 (N_18050,N_17886,N_17839);
nor U18051 (N_18051,N_17602,N_17921);
and U18052 (N_18052,N_17658,N_17648);
or U18053 (N_18053,N_17846,N_17950);
xor U18054 (N_18054,N_17743,N_17613);
and U18055 (N_18055,N_17644,N_17778);
or U18056 (N_18056,N_17815,N_17675);
nor U18057 (N_18057,N_17861,N_17742);
or U18058 (N_18058,N_17674,N_17948);
xnor U18059 (N_18059,N_17904,N_17957);
xor U18060 (N_18060,N_17898,N_17636);
or U18061 (N_18061,N_17939,N_17922);
or U18062 (N_18062,N_17760,N_17666);
and U18063 (N_18063,N_17638,N_17807);
or U18064 (N_18064,N_17683,N_17881);
nand U18065 (N_18065,N_17933,N_17729);
and U18066 (N_18066,N_17695,N_17672);
xnor U18067 (N_18067,N_17703,N_17750);
xnor U18068 (N_18068,N_17783,N_17769);
nand U18069 (N_18069,N_17734,N_17811);
nor U18070 (N_18070,N_17640,N_17645);
nor U18071 (N_18071,N_17691,N_17918);
or U18072 (N_18072,N_17995,N_17963);
or U18073 (N_18073,N_17851,N_17808);
or U18074 (N_18074,N_17779,N_17816);
nand U18075 (N_18075,N_17893,N_17690);
nand U18076 (N_18076,N_17736,N_17661);
and U18077 (N_18077,N_17984,N_17852);
or U18078 (N_18078,N_17857,N_17990);
and U18079 (N_18079,N_17947,N_17773);
and U18080 (N_18080,N_17931,N_17927);
xor U18081 (N_18081,N_17873,N_17788);
nor U18082 (N_18082,N_17775,N_17776);
and U18083 (N_18083,N_17792,N_17999);
nor U18084 (N_18084,N_17841,N_17771);
and U18085 (N_18085,N_17653,N_17973);
or U18086 (N_18086,N_17652,N_17814);
or U18087 (N_18087,N_17798,N_17623);
xnor U18088 (N_18088,N_17960,N_17630);
xnor U18089 (N_18089,N_17780,N_17925);
nor U18090 (N_18090,N_17649,N_17612);
or U18091 (N_18091,N_17911,N_17624);
or U18092 (N_18092,N_17824,N_17946);
nand U18093 (N_18093,N_17632,N_17606);
xnor U18094 (N_18094,N_17616,N_17979);
and U18095 (N_18095,N_17600,N_17909);
xnor U18096 (N_18096,N_17789,N_17897);
nand U18097 (N_18097,N_17688,N_17978);
xnor U18098 (N_18098,N_17784,N_17980);
and U18099 (N_18099,N_17754,N_17945);
and U18100 (N_18100,N_17768,N_17832);
nand U18101 (N_18101,N_17802,N_17704);
nand U18102 (N_18102,N_17974,N_17823);
nand U18103 (N_18103,N_17804,N_17671);
xor U18104 (N_18104,N_17799,N_17697);
nor U18105 (N_18105,N_17696,N_17830);
or U18106 (N_18106,N_17955,N_17887);
nor U18107 (N_18107,N_17711,N_17860);
nor U18108 (N_18108,N_17738,N_17634);
and U18109 (N_18109,N_17728,N_17976);
or U18110 (N_18110,N_17865,N_17603);
or U18111 (N_18111,N_17895,N_17882);
nor U18112 (N_18112,N_17629,N_17987);
and U18113 (N_18113,N_17643,N_17902);
or U18114 (N_18114,N_17739,N_17785);
nor U18115 (N_18115,N_17619,N_17845);
nor U18116 (N_18116,N_17854,N_17818);
or U18117 (N_18117,N_17907,N_17941);
nand U18118 (N_18118,N_17810,N_17713);
or U18119 (N_18119,N_17836,N_17878);
nor U18120 (N_18120,N_17847,N_17700);
or U18121 (N_18121,N_17964,N_17891);
nand U18122 (N_18122,N_17809,N_17764);
or U18123 (N_18123,N_17726,N_17833);
nand U18124 (N_18124,N_17840,N_17996);
xnor U18125 (N_18125,N_17635,N_17967);
nor U18126 (N_18126,N_17838,N_17953);
nand U18127 (N_18127,N_17662,N_17958);
nand U18128 (N_18128,N_17618,N_17819);
nor U18129 (N_18129,N_17642,N_17698);
or U18130 (N_18130,N_17676,N_17646);
nor U18131 (N_18131,N_17787,N_17981);
nor U18132 (N_18132,N_17822,N_17908);
and U18133 (N_18133,N_17994,N_17631);
or U18134 (N_18134,N_17826,N_17885);
nand U18135 (N_18135,N_17800,N_17915);
nor U18136 (N_18136,N_17835,N_17853);
and U18137 (N_18137,N_17761,N_17880);
and U18138 (N_18138,N_17997,N_17705);
and U18139 (N_18139,N_17844,N_17975);
xnor U18140 (N_18140,N_17870,N_17660);
or U18141 (N_18141,N_17617,N_17949);
or U18142 (N_18142,N_17607,N_17770);
nor U18143 (N_18143,N_17889,N_17935);
or U18144 (N_18144,N_17966,N_17917);
nand U18145 (N_18145,N_17609,N_17745);
or U18146 (N_18146,N_17831,N_17991);
nor U18147 (N_18147,N_17687,N_17782);
nor U18148 (N_18148,N_17723,N_17665);
or U18149 (N_18149,N_17725,N_17759);
or U18150 (N_18150,N_17667,N_17801);
nand U18151 (N_18151,N_17993,N_17702);
or U18152 (N_18152,N_17879,N_17610);
and U18153 (N_18153,N_17735,N_17986);
or U18154 (N_18154,N_17874,N_17718);
nor U18155 (N_18155,N_17716,N_17737);
nor U18156 (N_18156,N_17920,N_17693);
and U18157 (N_18157,N_17714,N_17786);
or U18158 (N_18158,N_17752,N_17932);
xor U18159 (N_18159,N_17708,N_17969);
xor U18160 (N_18160,N_17903,N_17625);
and U18161 (N_18161,N_17959,N_17722);
and U18162 (N_18162,N_17930,N_17781);
or U18163 (N_18163,N_17791,N_17842);
xor U18164 (N_18164,N_17682,N_17890);
nand U18165 (N_18165,N_17982,N_17615);
nor U18166 (N_18166,N_17654,N_17884);
nand U18167 (N_18167,N_17793,N_17621);
xor U18168 (N_18168,N_17919,N_17790);
or U18169 (N_18169,N_17650,N_17751);
nand U18170 (N_18170,N_17777,N_17924);
and U18171 (N_18171,N_17892,N_17748);
nor U18172 (N_18172,N_17940,N_17942);
or U18173 (N_18173,N_17679,N_17837);
or U18174 (N_18174,N_17965,N_17794);
nor U18175 (N_18175,N_17655,N_17943);
xnor U18176 (N_18176,N_17720,N_17741);
nand U18177 (N_18177,N_17876,N_17875);
or U18178 (N_18178,N_17709,N_17620);
or U18179 (N_18179,N_17856,N_17724);
nor U18180 (N_18180,N_17684,N_17968);
xor U18181 (N_18181,N_17899,N_17992);
nor U18182 (N_18182,N_17669,N_17961);
nand U18183 (N_18183,N_17906,N_17701);
nand U18184 (N_18184,N_17829,N_17869);
xnor U18185 (N_18185,N_17817,N_17749);
xnor U18186 (N_18186,N_17678,N_17862);
and U18187 (N_18187,N_17601,N_17692);
nor U18188 (N_18188,N_17628,N_17877);
or U18189 (N_18189,N_17872,N_17604);
nor U18190 (N_18190,N_17923,N_17944);
nor U18191 (N_18191,N_17821,N_17863);
and U18192 (N_18192,N_17867,N_17843);
or U18193 (N_18193,N_17954,N_17673);
and U18194 (N_18194,N_17900,N_17977);
xor U18195 (N_18195,N_17796,N_17834);
or U18196 (N_18196,N_17657,N_17731);
nand U18197 (N_18197,N_17755,N_17813);
and U18198 (N_18198,N_17828,N_17627);
nand U18199 (N_18199,N_17608,N_17681);
nand U18200 (N_18200,N_17666,N_17851);
xor U18201 (N_18201,N_17636,N_17986);
nand U18202 (N_18202,N_17941,N_17723);
and U18203 (N_18203,N_17907,N_17964);
nor U18204 (N_18204,N_17936,N_17702);
nor U18205 (N_18205,N_17779,N_17661);
and U18206 (N_18206,N_17974,N_17618);
nor U18207 (N_18207,N_17778,N_17642);
nor U18208 (N_18208,N_17689,N_17729);
nand U18209 (N_18209,N_17934,N_17792);
or U18210 (N_18210,N_17829,N_17900);
and U18211 (N_18211,N_17707,N_17600);
nand U18212 (N_18212,N_17725,N_17872);
xnor U18213 (N_18213,N_17967,N_17666);
xor U18214 (N_18214,N_17998,N_17942);
xnor U18215 (N_18215,N_17720,N_17996);
and U18216 (N_18216,N_17729,N_17798);
nand U18217 (N_18217,N_17760,N_17759);
nor U18218 (N_18218,N_17910,N_17692);
or U18219 (N_18219,N_17727,N_17814);
nor U18220 (N_18220,N_17735,N_17665);
xnor U18221 (N_18221,N_17957,N_17625);
and U18222 (N_18222,N_17889,N_17863);
nand U18223 (N_18223,N_17800,N_17671);
nor U18224 (N_18224,N_17848,N_17859);
nor U18225 (N_18225,N_17884,N_17857);
and U18226 (N_18226,N_17735,N_17625);
nand U18227 (N_18227,N_17803,N_17831);
nand U18228 (N_18228,N_17701,N_17799);
xor U18229 (N_18229,N_17893,N_17726);
or U18230 (N_18230,N_17781,N_17836);
xor U18231 (N_18231,N_17729,N_17804);
or U18232 (N_18232,N_17615,N_17836);
and U18233 (N_18233,N_17731,N_17805);
or U18234 (N_18234,N_17748,N_17629);
xor U18235 (N_18235,N_17889,N_17880);
nor U18236 (N_18236,N_17804,N_17641);
or U18237 (N_18237,N_17825,N_17602);
xnor U18238 (N_18238,N_17838,N_17861);
nor U18239 (N_18239,N_17604,N_17729);
xor U18240 (N_18240,N_17966,N_17949);
nor U18241 (N_18241,N_17950,N_17912);
xor U18242 (N_18242,N_17739,N_17974);
nor U18243 (N_18243,N_17861,N_17764);
nand U18244 (N_18244,N_17925,N_17758);
nand U18245 (N_18245,N_17824,N_17826);
or U18246 (N_18246,N_17796,N_17622);
and U18247 (N_18247,N_17683,N_17894);
or U18248 (N_18248,N_17723,N_17954);
xor U18249 (N_18249,N_17908,N_17738);
xnor U18250 (N_18250,N_17918,N_17824);
or U18251 (N_18251,N_17732,N_17841);
xnor U18252 (N_18252,N_17684,N_17784);
or U18253 (N_18253,N_17750,N_17630);
nand U18254 (N_18254,N_17910,N_17853);
and U18255 (N_18255,N_17932,N_17756);
xnor U18256 (N_18256,N_17676,N_17761);
nand U18257 (N_18257,N_17968,N_17993);
or U18258 (N_18258,N_17655,N_17931);
or U18259 (N_18259,N_17992,N_17931);
nor U18260 (N_18260,N_17821,N_17737);
xnor U18261 (N_18261,N_17600,N_17637);
xor U18262 (N_18262,N_17773,N_17926);
and U18263 (N_18263,N_17903,N_17963);
and U18264 (N_18264,N_17860,N_17994);
and U18265 (N_18265,N_17985,N_17601);
nand U18266 (N_18266,N_17657,N_17938);
xnor U18267 (N_18267,N_17861,N_17957);
or U18268 (N_18268,N_17828,N_17710);
and U18269 (N_18269,N_17923,N_17751);
nand U18270 (N_18270,N_17889,N_17790);
xnor U18271 (N_18271,N_17953,N_17632);
xnor U18272 (N_18272,N_17900,N_17614);
and U18273 (N_18273,N_17871,N_17979);
nand U18274 (N_18274,N_17742,N_17970);
nand U18275 (N_18275,N_17749,N_17973);
nor U18276 (N_18276,N_17788,N_17976);
nand U18277 (N_18277,N_17996,N_17745);
nand U18278 (N_18278,N_17756,N_17826);
xnor U18279 (N_18279,N_17709,N_17685);
or U18280 (N_18280,N_17909,N_17792);
xnor U18281 (N_18281,N_17783,N_17630);
nor U18282 (N_18282,N_17676,N_17763);
nor U18283 (N_18283,N_17881,N_17730);
or U18284 (N_18284,N_17763,N_17891);
nand U18285 (N_18285,N_17606,N_17721);
and U18286 (N_18286,N_17911,N_17859);
nand U18287 (N_18287,N_17767,N_17776);
and U18288 (N_18288,N_17674,N_17722);
nand U18289 (N_18289,N_17902,N_17870);
xnor U18290 (N_18290,N_17656,N_17704);
and U18291 (N_18291,N_17711,N_17865);
nor U18292 (N_18292,N_17746,N_17962);
and U18293 (N_18293,N_17782,N_17769);
nand U18294 (N_18294,N_17901,N_17689);
and U18295 (N_18295,N_17752,N_17970);
nor U18296 (N_18296,N_17725,N_17903);
nor U18297 (N_18297,N_17787,N_17752);
xor U18298 (N_18298,N_17667,N_17707);
and U18299 (N_18299,N_17752,N_17958);
and U18300 (N_18300,N_17847,N_17760);
xnor U18301 (N_18301,N_17685,N_17723);
nor U18302 (N_18302,N_17807,N_17955);
nor U18303 (N_18303,N_17911,N_17713);
xnor U18304 (N_18304,N_17904,N_17672);
nand U18305 (N_18305,N_17821,N_17649);
xnor U18306 (N_18306,N_17951,N_17793);
xor U18307 (N_18307,N_17896,N_17850);
xor U18308 (N_18308,N_17987,N_17621);
or U18309 (N_18309,N_17925,N_17957);
xnor U18310 (N_18310,N_17721,N_17944);
or U18311 (N_18311,N_17931,N_17823);
and U18312 (N_18312,N_17698,N_17952);
or U18313 (N_18313,N_17740,N_17874);
or U18314 (N_18314,N_17805,N_17670);
nand U18315 (N_18315,N_17921,N_17829);
xor U18316 (N_18316,N_17887,N_17899);
nand U18317 (N_18317,N_17839,N_17691);
or U18318 (N_18318,N_17856,N_17754);
nand U18319 (N_18319,N_17607,N_17717);
nor U18320 (N_18320,N_17864,N_17758);
xnor U18321 (N_18321,N_17646,N_17631);
nor U18322 (N_18322,N_17748,N_17993);
and U18323 (N_18323,N_17999,N_17789);
nand U18324 (N_18324,N_17640,N_17711);
xor U18325 (N_18325,N_17774,N_17763);
nor U18326 (N_18326,N_17896,N_17952);
or U18327 (N_18327,N_17963,N_17797);
xnor U18328 (N_18328,N_17696,N_17784);
nand U18329 (N_18329,N_17783,N_17885);
nand U18330 (N_18330,N_17834,N_17676);
nand U18331 (N_18331,N_17667,N_17735);
nand U18332 (N_18332,N_17907,N_17606);
nor U18333 (N_18333,N_17907,N_17677);
and U18334 (N_18334,N_17998,N_17645);
xnor U18335 (N_18335,N_17687,N_17748);
and U18336 (N_18336,N_17750,N_17695);
or U18337 (N_18337,N_17806,N_17859);
and U18338 (N_18338,N_17971,N_17864);
nor U18339 (N_18339,N_17719,N_17790);
nand U18340 (N_18340,N_17685,N_17662);
nand U18341 (N_18341,N_17733,N_17701);
xor U18342 (N_18342,N_17997,N_17876);
nand U18343 (N_18343,N_17853,N_17719);
xnor U18344 (N_18344,N_17825,N_17796);
and U18345 (N_18345,N_17740,N_17654);
xnor U18346 (N_18346,N_17720,N_17735);
nor U18347 (N_18347,N_17620,N_17949);
and U18348 (N_18348,N_17908,N_17973);
nand U18349 (N_18349,N_17802,N_17949);
and U18350 (N_18350,N_17936,N_17606);
and U18351 (N_18351,N_17847,N_17968);
nor U18352 (N_18352,N_17674,N_17864);
and U18353 (N_18353,N_17662,N_17902);
or U18354 (N_18354,N_17793,N_17928);
nand U18355 (N_18355,N_17813,N_17699);
nand U18356 (N_18356,N_17836,N_17815);
or U18357 (N_18357,N_17640,N_17880);
xnor U18358 (N_18358,N_17872,N_17944);
nor U18359 (N_18359,N_17652,N_17607);
or U18360 (N_18360,N_17690,N_17752);
and U18361 (N_18361,N_17909,N_17783);
nor U18362 (N_18362,N_17945,N_17924);
nand U18363 (N_18363,N_17991,N_17644);
nand U18364 (N_18364,N_17810,N_17729);
nand U18365 (N_18365,N_17776,N_17788);
and U18366 (N_18366,N_17989,N_17607);
and U18367 (N_18367,N_17699,N_17760);
and U18368 (N_18368,N_17982,N_17685);
nand U18369 (N_18369,N_17888,N_17859);
or U18370 (N_18370,N_17736,N_17887);
and U18371 (N_18371,N_17993,N_17737);
xor U18372 (N_18372,N_17830,N_17833);
xor U18373 (N_18373,N_17624,N_17909);
or U18374 (N_18374,N_17775,N_17636);
nand U18375 (N_18375,N_17982,N_17600);
nor U18376 (N_18376,N_17629,N_17734);
nand U18377 (N_18377,N_17827,N_17994);
xor U18378 (N_18378,N_17634,N_17685);
or U18379 (N_18379,N_17630,N_17934);
nand U18380 (N_18380,N_17784,N_17715);
xor U18381 (N_18381,N_17710,N_17737);
xor U18382 (N_18382,N_17796,N_17958);
xor U18383 (N_18383,N_17973,N_17638);
nand U18384 (N_18384,N_17643,N_17623);
and U18385 (N_18385,N_17684,N_17770);
or U18386 (N_18386,N_17857,N_17733);
and U18387 (N_18387,N_17868,N_17636);
nand U18388 (N_18388,N_17676,N_17847);
xor U18389 (N_18389,N_17930,N_17901);
or U18390 (N_18390,N_17960,N_17896);
or U18391 (N_18391,N_17941,N_17902);
nand U18392 (N_18392,N_17689,N_17703);
nand U18393 (N_18393,N_17947,N_17868);
and U18394 (N_18394,N_17985,N_17855);
nor U18395 (N_18395,N_17970,N_17991);
xnor U18396 (N_18396,N_17799,N_17648);
or U18397 (N_18397,N_17920,N_17912);
nor U18398 (N_18398,N_17840,N_17970);
and U18399 (N_18399,N_17663,N_17907);
and U18400 (N_18400,N_18205,N_18341);
and U18401 (N_18401,N_18044,N_18294);
xor U18402 (N_18402,N_18351,N_18189);
nor U18403 (N_18403,N_18290,N_18169);
nand U18404 (N_18404,N_18021,N_18061);
or U18405 (N_18405,N_18122,N_18299);
nor U18406 (N_18406,N_18355,N_18014);
nor U18407 (N_18407,N_18292,N_18396);
or U18408 (N_18408,N_18243,N_18229);
nor U18409 (N_18409,N_18285,N_18007);
and U18410 (N_18410,N_18356,N_18390);
nand U18411 (N_18411,N_18043,N_18391);
nand U18412 (N_18412,N_18184,N_18198);
xor U18413 (N_18413,N_18002,N_18338);
and U18414 (N_18414,N_18112,N_18016);
and U18415 (N_18415,N_18067,N_18028);
or U18416 (N_18416,N_18042,N_18328);
nand U18417 (N_18417,N_18045,N_18340);
or U18418 (N_18418,N_18160,N_18202);
or U18419 (N_18419,N_18135,N_18240);
or U18420 (N_18420,N_18241,N_18245);
nor U18421 (N_18421,N_18050,N_18327);
nand U18422 (N_18422,N_18360,N_18389);
nand U18423 (N_18423,N_18309,N_18102);
or U18424 (N_18424,N_18176,N_18171);
or U18425 (N_18425,N_18000,N_18380);
nand U18426 (N_18426,N_18316,N_18311);
nor U18427 (N_18427,N_18395,N_18153);
or U18428 (N_18428,N_18190,N_18249);
and U18429 (N_18429,N_18293,N_18058);
xor U18430 (N_18430,N_18110,N_18098);
and U18431 (N_18431,N_18142,N_18362);
nand U18432 (N_18432,N_18247,N_18074);
xnor U18433 (N_18433,N_18126,N_18315);
and U18434 (N_18434,N_18257,N_18099);
nor U18435 (N_18435,N_18371,N_18270);
xnor U18436 (N_18436,N_18048,N_18230);
xnor U18437 (N_18437,N_18124,N_18162);
and U18438 (N_18438,N_18232,N_18200);
nand U18439 (N_18439,N_18023,N_18064);
nand U18440 (N_18440,N_18033,N_18031);
and U18441 (N_18441,N_18361,N_18280);
xnor U18442 (N_18442,N_18121,N_18339);
and U18443 (N_18443,N_18182,N_18310);
and U18444 (N_18444,N_18273,N_18348);
nand U18445 (N_18445,N_18363,N_18368);
and U18446 (N_18446,N_18277,N_18196);
or U18447 (N_18447,N_18019,N_18344);
nand U18448 (N_18448,N_18386,N_18265);
xor U18449 (N_18449,N_18313,N_18013);
or U18450 (N_18450,N_18103,N_18178);
and U18451 (N_18451,N_18003,N_18300);
and U18452 (N_18452,N_18051,N_18111);
or U18453 (N_18453,N_18125,N_18226);
or U18454 (N_18454,N_18185,N_18297);
nand U18455 (N_18455,N_18094,N_18318);
and U18456 (N_18456,N_18131,N_18161);
nand U18457 (N_18457,N_18156,N_18377);
nor U18458 (N_18458,N_18283,N_18133);
xnor U18459 (N_18459,N_18070,N_18063);
nand U18460 (N_18460,N_18254,N_18199);
xnor U18461 (N_18461,N_18213,N_18286);
and U18462 (N_18462,N_18253,N_18250);
nand U18463 (N_18463,N_18365,N_18062);
nor U18464 (N_18464,N_18346,N_18271);
nor U18465 (N_18465,N_18352,N_18109);
and U18466 (N_18466,N_18204,N_18137);
and U18467 (N_18467,N_18218,N_18015);
nor U18468 (N_18468,N_18095,N_18321);
and U18469 (N_18469,N_18179,N_18319);
or U18470 (N_18470,N_18260,N_18130);
or U18471 (N_18471,N_18100,N_18382);
nor U18472 (N_18472,N_18214,N_18276);
xnor U18473 (N_18473,N_18069,N_18312);
nor U18474 (N_18474,N_18008,N_18248);
and U18475 (N_18475,N_18080,N_18372);
or U18476 (N_18476,N_18084,N_18275);
xor U18477 (N_18477,N_18223,N_18017);
nor U18478 (N_18478,N_18056,N_18059);
or U18479 (N_18479,N_18193,N_18195);
nand U18480 (N_18480,N_18295,N_18366);
and U18481 (N_18481,N_18227,N_18188);
or U18482 (N_18482,N_18082,N_18136);
or U18483 (N_18483,N_18030,N_18272);
nand U18484 (N_18484,N_18212,N_18376);
xnor U18485 (N_18485,N_18224,N_18107);
nand U18486 (N_18486,N_18337,N_18177);
nand U18487 (N_18487,N_18055,N_18369);
or U18488 (N_18488,N_18251,N_18047);
and U18489 (N_18489,N_18113,N_18208);
xor U18490 (N_18490,N_18163,N_18284);
or U18491 (N_18491,N_18154,N_18262);
nand U18492 (N_18492,N_18018,N_18012);
or U18493 (N_18493,N_18001,N_18020);
or U18494 (N_18494,N_18073,N_18239);
nor U18495 (N_18495,N_18215,N_18237);
or U18496 (N_18496,N_18106,N_18201);
or U18497 (N_18497,N_18090,N_18168);
and U18498 (N_18498,N_18308,N_18374);
or U18499 (N_18499,N_18378,N_18332);
and U18500 (N_18500,N_18035,N_18221);
or U18501 (N_18501,N_18115,N_18025);
xor U18502 (N_18502,N_18225,N_18333);
or U18503 (N_18503,N_18342,N_18258);
xor U18504 (N_18504,N_18298,N_18141);
nor U18505 (N_18505,N_18246,N_18139);
or U18506 (N_18506,N_18120,N_18116);
and U18507 (N_18507,N_18104,N_18037);
or U18508 (N_18508,N_18194,N_18119);
and U18509 (N_18509,N_18167,N_18370);
nor U18510 (N_18510,N_18092,N_18173);
nor U18511 (N_18511,N_18353,N_18005);
and U18512 (N_18512,N_18029,N_18235);
xnor U18513 (N_18513,N_18083,N_18209);
nor U18514 (N_18514,N_18326,N_18128);
xor U18515 (N_18515,N_18259,N_18296);
nand U18516 (N_18516,N_18117,N_18279);
and U18517 (N_18517,N_18036,N_18041);
xor U18518 (N_18518,N_18192,N_18317);
xnor U18519 (N_18519,N_18206,N_18373);
or U18520 (N_18520,N_18207,N_18076);
and U18521 (N_18521,N_18088,N_18320);
and U18522 (N_18522,N_18152,N_18331);
or U18523 (N_18523,N_18278,N_18175);
or U18524 (N_18524,N_18144,N_18097);
nor U18525 (N_18525,N_18281,N_18387);
or U18526 (N_18526,N_18228,N_18096);
xnor U18527 (N_18527,N_18040,N_18211);
nand U18528 (N_18528,N_18306,N_18345);
nand U18529 (N_18529,N_18398,N_18089);
and U18530 (N_18530,N_18108,N_18138);
xnor U18531 (N_18531,N_18392,N_18384);
nand U18532 (N_18532,N_18264,N_18336);
or U18533 (N_18533,N_18079,N_18255);
xnor U18534 (N_18534,N_18009,N_18054);
and U18535 (N_18535,N_18081,N_18305);
and U18536 (N_18536,N_18129,N_18216);
and U18537 (N_18537,N_18314,N_18354);
nand U18538 (N_18538,N_18350,N_18191);
nor U18539 (N_18539,N_18397,N_18078);
and U18540 (N_18540,N_18269,N_18220);
and U18541 (N_18541,N_18166,N_18071);
or U18542 (N_18542,N_18375,N_18066);
or U18543 (N_18543,N_18266,N_18263);
nand U18544 (N_18544,N_18261,N_18186);
or U18545 (N_18545,N_18150,N_18157);
xor U18546 (N_18546,N_18301,N_18335);
xor U18547 (N_18547,N_18343,N_18307);
nor U18548 (N_18548,N_18087,N_18038);
and U18549 (N_18549,N_18183,N_18347);
xnor U18550 (N_18550,N_18222,N_18134);
or U18551 (N_18551,N_18385,N_18236);
nand U18552 (N_18552,N_18151,N_18143);
nand U18553 (N_18553,N_18057,N_18118);
nor U18554 (N_18554,N_18091,N_18068);
and U18555 (N_18555,N_18197,N_18114);
and U18556 (N_18556,N_18325,N_18304);
nand U18557 (N_18557,N_18274,N_18324);
and U18558 (N_18558,N_18077,N_18252);
xor U18559 (N_18559,N_18123,N_18242);
nand U18560 (N_18560,N_18367,N_18004);
nand U18561 (N_18561,N_18145,N_18388);
xor U18562 (N_18562,N_18359,N_18268);
xor U18563 (N_18563,N_18233,N_18394);
xnor U18564 (N_18564,N_18231,N_18244);
xnor U18565 (N_18565,N_18149,N_18155);
nor U18566 (N_18566,N_18302,N_18364);
and U18567 (N_18567,N_18219,N_18234);
xor U18568 (N_18568,N_18101,N_18267);
or U18569 (N_18569,N_18011,N_18010);
nor U18570 (N_18570,N_18381,N_18127);
and U18571 (N_18571,N_18032,N_18075);
nand U18572 (N_18572,N_18132,N_18060);
nor U18573 (N_18573,N_18148,N_18203);
nand U18574 (N_18574,N_18334,N_18383);
xor U18575 (N_18575,N_18323,N_18399);
nor U18576 (N_18576,N_18322,N_18358);
xnor U18577 (N_18577,N_18034,N_18164);
and U18578 (N_18578,N_18181,N_18086);
or U18579 (N_18579,N_18165,N_18026);
or U18580 (N_18580,N_18330,N_18174);
or U18581 (N_18581,N_18187,N_18147);
and U18582 (N_18582,N_18393,N_18024);
nor U18583 (N_18583,N_18210,N_18291);
xor U18584 (N_18584,N_18140,N_18238);
nand U18585 (N_18585,N_18046,N_18085);
nor U18586 (N_18586,N_18329,N_18172);
or U18587 (N_18587,N_18049,N_18282);
or U18588 (N_18588,N_18093,N_18217);
xnor U18589 (N_18589,N_18288,N_18052);
and U18590 (N_18590,N_18303,N_18158);
nor U18591 (N_18591,N_18159,N_18053);
nor U18592 (N_18592,N_18170,N_18146);
or U18593 (N_18593,N_18357,N_18105);
and U18594 (N_18594,N_18349,N_18256);
and U18595 (N_18595,N_18180,N_18027);
and U18596 (N_18596,N_18006,N_18072);
xor U18597 (N_18597,N_18065,N_18379);
and U18598 (N_18598,N_18022,N_18287);
or U18599 (N_18599,N_18039,N_18289);
nor U18600 (N_18600,N_18085,N_18395);
or U18601 (N_18601,N_18010,N_18112);
or U18602 (N_18602,N_18025,N_18032);
nand U18603 (N_18603,N_18279,N_18322);
nand U18604 (N_18604,N_18376,N_18173);
xnor U18605 (N_18605,N_18379,N_18384);
nor U18606 (N_18606,N_18199,N_18304);
or U18607 (N_18607,N_18121,N_18311);
nand U18608 (N_18608,N_18068,N_18220);
xnor U18609 (N_18609,N_18279,N_18184);
and U18610 (N_18610,N_18292,N_18087);
nand U18611 (N_18611,N_18232,N_18297);
nand U18612 (N_18612,N_18242,N_18124);
nor U18613 (N_18613,N_18269,N_18166);
xnor U18614 (N_18614,N_18038,N_18335);
nor U18615 (N_18615,N_18187,N_18061);
nor U18616 (N_18616,N_18002,N_18391);
nor U18617 (N_18617,N_18223,N_18107);
xor U18618 (N_18618,N_18307,N_18212);
nor U18619 (N_18619,N_18051,N_18152);
nor U18620 (N_18620,N_18215,N_18158);
nor U18621 (N_18621,N_18353,N_18198);
nor U18622 (N_18622,N_18180,N_18138);
nand U18623 (N_18623,N_18261,N_18077);
and U18624 (N_18624,N_18238,N_18233);
nand U18625 (N_18625,N_18252,N_18012);
nor U18626 (N_18626,N_18331,N_18073);
nand U18627 (N_18627,N_18396,N_18348);
nand U18628 (N_18628,N_18253,N_18143);
nand U18629 (N_18629,N_18395,N_18239);
nor U18630 (N_18630,N_18084,N_18263);
or U18631 (N_18631,N_18263,N_18127);
and U18632 (N_18632,N_18276,N_18018);
nand U18633 (N_18633,N_18195,N_18277);
and U18634 (N_18634,N_18035,N_18075);
nor U18635 (N_18635,N_18300,N_18370);
nand U18636 (N_18636,N_18071,N_18061);
and U18637 (N_18637,N_18355,N_18231);
or U18638 (N_18638,N_18378,N_18228);
or U18639 (N_18639,N_18220,N_18289);
nor U18640 (N_18640,N_18368,N_18021);
xnor U18641 (N_18641,N_18299,N_18349);
nand U18642 (N_18642,N_18122,N_18374);
nor U18643 (N_18643,N_18268,N_18017);
nand U18644 (N_18644,N_18266,N_18265);
xor U18645 (N_18645,N_18230,N_18395);
xor U18646 (N_18646,N_18170,N_18337);
or U18647 (N_18647,N_18358,N_18026);
and U18648 (N_18648,N_18032,N_18058);
nor U18649 (N_18649,N_18222,N_18099);
xnor U18650 (N_18650,N_18279,N_18363);
or U18651 (N_18651,N_18327,N_18171);
or U18652 (N_18652,N_18142,N_18347);
xor U18653 (N_18653,N_18017,N_18288);
and U18654 (N_18654,N_18357,N_18160);
nor U18655 (N_18655,N_18155,N_18367);
and U18656 (N_18656,N_18051,N_18233);
nand U18657 (N_18657,N_18377,N_18152);
or U18658 (N_18658,N_18100,N_18155);
and U18659 (N_18659,N_18110,N_18320);
xnor U18660 (N_18660,N_18338,N_18104);
nor U18661 (N_18661,N_18114,N_18202);
xnor U18662 (N_18662,N_18376,N_18321);
or U18663 (N_18663,N_18307,N_18162);
or U18664 (N_18664,N_18246,N_18184);
or U18665 (N_18665,N_18223,N_18327);
nor U18666 (N_18666,N_18337,N_18075);
or U18667 (N_18667,N_18270,N_18133);
nor U18668 (N_18668,N_18169,N_18202);
nor U18669 (N_18669,N_18029,N_18150);
and U18670 (N_18670,N_18356,N_18199);
or U18671 (N_18671,N_18214,N_18140);
and U18672 (N_18672,N_18383,N_18230);
or U18673 (N_18673,N_18214,N_18320);
xnor U18674 (N_18674,N_18207,N_18206);
and U18675 (N_18675,N_18257,N_18175);
and U18676 (N_18676,N_18162,N_18333);
nor U18677 (N_18677,N_18315,N_18125);
and U18678 (N_18678,N_18336,N_18073);
xor U18679 (N_18679,N_18093,N_18109);
nor U18680 (N_18680,N_18359,N_18339);
nor U18681 (N_18681,N_18116,N_18062);
and U18682 (N_18682,N_18312,N_18199);
and U18683 (N_18683,N_18063,N_18083);
xnor U18684 (N_18684,N_18382,N_18282);
nand U18685 (N_18685,N_18245,N_18361);
or U18686 (N_18686,N_18122,N_18381);
or U18687 (N_18687,N_18181,N_18044);
nor U18688 (N_18688,N_18036,N_18035);
nand U18689 (N_18689,N_18300,N_18340);
xor U18690 (N_18690,N_18087,N_18073);
nand U18691 (N_18691,N_18206,N_18122);
xnor U18692 (N_18692,N_18294,N_18214);
or U18693 (N_18693,N_18139,N_18304);
nor U18694 (N_18694,N_18106,N_18147);
nand U18695 (N_18695,N_18005,N_18015);
nor U18696 (N_18696,N_18129,N_18053);
xnor U18697 (N_18697,N_18386,N_18379);
xor U18698 (N_18698,N_18082,N_18220);
or U18699 (N_18699,N_18004,N_18117);
or U18700 (N_18700,N_18386,N_18030);
xor U18701 (N_18701,N_18271,N_18064);
nor U18702 (N_18702,N_18162,N_18199);
or U18703 (N_18703,N_18356,N_18313);
nor U18704 (N_18704,N_18314,N_18089);
and U18705 (N_18705,N_18261,N_18300);
nand U18706 (N_18706,N_18310,N_18398);
or U18707 (N_18707,N_18221,N_18247);
nor U18708 (N_18708,N_18054,N_18339);
and U18709 (N_18709,N_18185,N_18245);
or U18710 (N_18710,N_18183,N_18231);
or U18711 (N_18711,N_18137,N_18171);
or U18712 (N_18712,N_18278,N_18398);
or U18713 (N_18713,N_18393,N_18232);
nand U18714 (N_18714,N_18186,N_18120);
and U18715 (N_18715,N_18380,N_18264);
and U18716 (N_18716,N_18244,N_18316);
or U18717 (N_18717,N_18397,N_18092);
and U18718 (N_18718,N_18045,N_18212);
or U18719 (N_18719,N_18189,N_18044);
or U18720 (N_18720,N_18148,N_18174);
or U18721 (N_18721,N_18166,N_18262);
or U18722 (N_18722,N_18125,N_18372);
xor U18723 (N_18723,N_18198,N_18299);
xnor U18724 (N_18724,N_18068,N_18398);
nor U18725 (N_18725,N_18341,N_18222);
xnor U18726 (N_18726,N_18392,N_18058);
nor U18727 (N_18727,N_18382,N_18059);
or U18728 (N_18728,N_18124,N_18055);
xnor U18729 (N_18729,N_18136,N_18228);
or U18730 (N_18730,N_18289,N_18237);
nor U18731 (N_18731,N_18152,N_18374);
nor U18732 (N_18732,N_18103,N_18312);
nor U18733 (N_18733,N_18125,N_18336);
or U18734 (N_18734,N_18028,N_18318);
and U18735 (N_18735,N_18047,N_18050);
xor U18736 (N_18736,N_18010,N_18266);
xor U18737 (N_18737,N_18106,N_18008);
nor U18738 (N_18738,N_18399,N_18343);
and U18739 (N_18739,N_18035,N_18003);
nand U18740 (N_18740,N_18016,N_18321);
and U18741 (N_18741,N_18168,N_18182);
and U18742 (N_18742,N_18016,N_18343);
nor U18743 (N_18743,N_18242,N_18252);
xor U18744 (N_18744,N_18134,N_18083);
xor U18745 (N_18745,N_18263,N_18251);
nand U18746 (N_18746,N_18167,N_18089);
and U18747 (N_18747,N_18360,N_18230);
xor U18748 (N_18748,N_18153,N_18151);
or U18749 (N_18749,N_18030,N_18352);
nor U18750 (N_18750,N_18268,N_18228);
or U18751 (N_18751,N_18027,N_18185);
and U18752 (N_18752,N_18024,N_18161);
nor U18753 (N_18753,N_18393,N_18305);
xor U18754 (N_18754,N_18338,N_18009);
nand U18755 (N_18755,N_18325,N_18132);
nand U18756 (N_18756,N_18386,N_18281);
nand U18757 (N_18757,N_18297,N_18325);
or U18758 (N_18758,N_18216,N_18094);
and U18759 (N_18759,N_18150,N_18358);
xor U18760 (N_18760,N_18334,N_18260);
nand U18761 (N_18761,N_18190,N_18036);
nor U18762 (N_18762,N_18170,N_18320);
nand U18763 (N_18763,N_18189,N_18128);
or U18764 (N_18764,N_18359,N_18077);
and U18765 (N_18765,N_18236,N_18239);
nor U18766 (N_18766,N_18230,N_18086);
nor U18767 (N_18767,N_18273,N_18184);
nand U18768 (N_18768,N_18342,N_18269);
or U18769 (N_18769,N_18014,N_18100);
or U18770 (N_18770,N_18183,N_18265);
or U18771 (N_18771,N_18023,N_18212);
and U18772 (N_18772,N_18015,N_18378);
or U18773 (N_18773,N_18275,N_18270);
or U18774 (N_18774,N_18243,N_18024);
nor U18775 (N_18775,N_18079,N_18114);
or U18776 (N_18776,N_18221,N_18399);
nor U18777 (N_18777,N_18085,N_18397);
and U18778 (N_18778,N_18211,N_18172);
nor U18779 (N_18779,N_18213,N_18122);
or U18780 (N_18780,N_18053,N_18175);
nor U18781 (N_18781,N_18023,N_18323);
xnor U18782 (N_18782,N_18298,N_18142);
nand U18783 (N_18783,N_18313,N_18353);
nand U18784 (N_18784,N_18210,N_18006);
nand U18785 (N_18785,N_18234,N_18181);
and U18786 (N_18786,N_18261,N_18346);
or U18787 (N_18787,N_18036,N_18115);
and U18788 (N_18788,N_18011,N_18245);
or U18789 (N_18789,N_18091,N_18080);
or U18790 (N_18790,N_18360,N_18353);
nand U18791 (N_18791,N_18201,N_18174);
and U18792 (N_18792,N_18005,N_18155);
nand U18793 (N_18793,N_18377,N_18238);
xor U18794 (N_18794,N_18381,N_18273);
and U18795 (N_18795,N_18074,N_18262);
nand U18796 (N_18796,N_18314,N_18307);
and U18797 (N_18797,N_18378,N_18157);
and U18798 (N_18798,N_18371,N_18106);
nor U18799 (N_18799,N_18053,N_18217);
and U18800 (N_18800,N_18722,N_18443);
and U18801 (N_18801,N_18473,N_18735);
or U18802 (N_18802,N_18749,N_18419);
and U18803 (N_18803,N_18799,N_18734);
and U18804 (N_18804,N_18669,N_18501);
nor U18805 (N_18805,N_18630,N_18724);
xnor U18806 (N_18806,N_18467,N_18449);
and U18807 (N_18807,N_18486,N_18521);
xnor U18808 (N_18808,N_18791,N_18575);
and U18809 (N_18809,N_18779,N_18455);
and U18810 (N_18810,N_18661,N_18423);
or U18811 (N_18811,N_18551,N_18634);
xor U18812 (N_18812,N_18565,N_18556);
or U18813 (N_18813,N_18766,N_18579);
nand U18814 (N_18814,N_18441,N_18445);
nand U18815 (N_18815,N_18499,N_18746);
nand U18816 (N_18816,N_18438,N_18797);
xnor U18817 (N_18817,N_18462,N_18554);
xnor U18818 (N_18818,N_18402,N_18726);
nand U18819 (N_18819,N_18586,N_18437);
nand U18820 (N_18820,N_18733,N_18631);
nor U18821 (N_18821,N_18622,N_18720);
and U18822 (N_18822,N_18715,N_18599);
or U18823 (N_18823,N_18525,N_18745);
nor U18824 (N_18824,N_18689,N_18500);
and U18825 (N_18825,N_18415,N_18721);
nor U18826 (N_18826,N_18601,N_18616);
nor U18827 (N_18827,N_18709,N_18483);
nor U18828 (N_18828,N_18686,N_18585);
xnor U18829 (N_18829,N_18422,N_18411);
or U18830 (N_18830,N_18490,N_18566);
nand U18831 (N_18831,N_18608,N_18667);
nor U18832 (N_18832,N_18613,N_18489);
nand U18833 (N_18833,N_18407,N_18729);
and U18834 (N_18834,N_18447,N_18503);
nor U18835 (N_18835,N_18452,N_18536);
nor U18836 (N_18836,N_18756,N_18493);
and U18837 (N_18837,N_18535,N_18658);
nand U18838 (N_18838,N_18714,N_18642);
xnor U18839 (N_18839,N_18614,N_18646);
and U18840 (N_18840,N_18540,N_18636);
nor U18841 (N_18841,N_18748,N_18428);
xor U18842 (N_18842,N_18728,N_18479);
or U18843 (N_18843,N_18727,N_18533);
xnor U18844 (N_18844,N_18659,N_18460);
or U18845 (N_18845,N_18628,N_18522);
xor U18846 (N_18846,N_18760,N_18773);
nor U18847 (N_18847,N_18676,N_18732);
nor U18848 (N_18848,N_18534,N_18738);
or U18849 (N_18849,N_18708,N_18641);
nor U18850 (N_18850,N_18427,N_18516);
or U18851 (N_18851,N_18764,N_18456);
nor U18852 (N_18852,N_18504,N_18581);
xor U18853 (N_18853,N_18767,N_18472);
nand U18854 (N_18854,N_18731,N_18719);
xnor U18855 (N_18855,N_18528,N_18584);
nand U18856 (N_18856,N_18673,N_18702);
or U18857 (N_18857,N_18555,N_18648);
nor U18858 (N_18858,N_18795,N_18712);
nor U18859 (N_18859,N_18587,N_18704);
nor U18860 (N_18860,N_18538,N_18639);
and U18861 (N_18861,N_18753,N_18537);
and U18862 (N_18862,N_18482,N_18693);
or U18863 (N_18863,N_18792,N_18434);
nand U18864 (N_18864,N_18511,N_18796);
and U18865 (N_18865,N_18624,N_18692);
and U18866 (N_18866,N_18530,N_18591);
xnor U18867 (N_18867,N_18562,N_18776);
xor U18868 (N_18868,N_18426,N_18671);
nor U18869 (N_18869,N_18644,N_18739);
nand U18870 (N_18870,N_18632,N_18758);
and U18871 (N_18871,N_18546,N_18410);
and U18872 (N_18872,N_18783,N_18424);
or U18873 (N_18873,N_18457,N_18408);
nor U18874 (N_18874,N_18544,N_18567);
nand U18875 (N_18875,N_18588,N_18403);
or U18876 (N_18876,N_18435,N_18469);
nand U18877 (N_18877,N_18744,N_18543);
xor U18878 (N_18878,N_18515,N_18468);
nor U18879 (N_18879,N_18514,N_18774);
and U18880 (N_18880,N_18763,N_18524);
or U18881 (N_18881,N_18418,N_18694);
nor U18882 (N_18882,N_18578,N_18505);
or U18883 (N_18883,N_18770,N_18723);
nor U18884 (N_18884,N_18655,N_18713);
xor U18885 (N_18885,N_18737,N_18409);
xnor U18886 (N_18886,N_18789,N_18668);
xor U18887 (N_18887,N_18548,N_18561);
nor U18888 (N_18888,N_18609,N_18549);
xnor U18889 (N_18889,N_18681,N_18518);
and U18890 (N_18890,N_18442,N_18627);
nor U18891 (N_18891,N_18782,N_18621);
nor U18892 (N_18892,N_18401,N_18510);
and U18893 (N_18893,N_18698,N_18463);
and U18894 (N_18894,N_18492,N_18574);
or U18895 (N_18895,N_18421,N_18718);
or U18896 (N_18896,N_18666,N_18663);
xnor U18897 (N_18897,N_18619,N_18559);
nand U18898 (N_18898,N_18761,N_18598);
nand U18899 (N_18899,N_18592,N_18605);
or U18900 (N_18900,N_18612,N_18496);
nor U18901 (N_18901,N_18684,N_18470);
nand U18902 (N_18902,N_18725,N_18454);
or U18903 (N_18903,N_18741,N_18705);
and U18904 (N_18904,N_18520,N_18414);
nor U18905 (N_18905,N_18425,N_18651);
or U18906 (N_18906,N_18593,N_18664);
and U18907 (N_18907,N_18772,N_18784);
xnor U18908 (N_18908,N_18440,N_18485);
xor U18909 (N_18909,N_18637,N_18618);
or U18910 (N_18910,N_18602,N_18610);
xor U18911 (N_18911,N_18620,N_18570);
nand U18912 (N_18912,N_18569,N_18711);
nand U18913 (N_18913,N_18786,N_18560);
nand U18914 (N_18914,N_18446,N_18458);
and U18915 (N_18915,N_18706,N_18696);
nor U18916 (N_18916,N_18640,N_18406);
nand U18917 (N_18917,N_18471,N_18682);
nor U18918 (N_18918,N_18430,N_18436);
or U18919 (N_18919,N_18769,N_18701);
or U18920 (N_18920,N_18573,N_18757);
xor U18921 (N_18921,N_18781,N_18547);
and U18922 (N_18922,N_18459,N_18649);
nand U18923 (N_18923,N_18710,N_18539);
nor U18924 (N_18924,N_18572,N_18771);
and U18925 (N_18925,N_18595,N_18527);
nor U18926 (N_18926,N_18506,N_18662);
xor U18927 (N_18927,N_18798,N_18400);
xnor U18928 (N_18928,N_18563,N_18532);
and U18929 (N_18929,N_18589,N_18477);
nor U18930 (N_18930,N_18747,N_18451);
or U18931 (N_18931,N_18793,N_18432);
nand U18932 (N_18932,N_18507,N_18464);
nor U18933 (N_18933,N_18583,N_18775);
nand U18934 (N_18934,N_18635,N_18420);
xnor U18935 (N_18935,N_18652,N_18759);
nand U18936 (N_18936,N_18794,N_18582);
nor U18937 (N_18937,N_18703,N_18476);
nor U18938 (N_18938,N_18596,N_18778);
xnor U18939 (N_18939,N_18675,N_18580);
xor U18940 (N_18940,N_18558,N_18431);
and U18941 (N_18941,N_18626,N_18541);
xnor U18942 (N_18942,N_18475,N_18752);
or U18943 (N_18943,N_18404,N_18685);
nor U18944 (N_18944,N_18638,N_18577);
or U18945 (N_18945,N_18754,N_18680);
and U18946 (N_18946,N_18512,N_18590);
or U18947 (N_18947,N_18660,N_18683);
nand U18948 (N_18948,N_18607,N_18755);
and U18949 (N_18949,N_18450,N_18617);
nand U18950 (N_18950,N_18699,N_18571);
xnor U18951 (N_18951,N_18788,N_18597);
nor U18952 (N_18952,N_18513,N_18790);
or U18953 (N_18953,N_18768,N_18780);
or U18954 (N_18954,N_18487,N_18629);
nand U18955 (N_18955,N_18785,N_18656);
or U18956 (N_18956,N_18679,N_18695);
xnor U18957 (N_18957,N_18657,N_18448);
and U18958 (N_18958,N_18765,N_18466);
or U18959 (N_18959,N_18716,N_18568);
xnor U18960 (N_18960,N_18481,N_18542);
nor U18961 (N_18961,N_18461,N_18650);
or U18962 (N_18962,N_18416,N_18654);
or U18963 (N_18963,N_18526,N_18550);
xor U18964 (N_18964,N_18643,N_18484);
and U18965 (N_18965,N_18751,N_18633);
xor U18966 (N_18966,N_18413,N_18677);
or U18967 (N_18967,N_18678,N_18687);
or U18968 (N_18968,N_18611,N_18730);
nand U18969 (N_18969,N_18498,N_18743);
nand U18970 (N_18970,N_18519,N_18552);
nor U18971 (N_18971,N_18576,N_18502);
nand U18972 (N_18972,N_18508,N_18529);
nor U18973 (N_18973,N_18750,N_18688);
nand U18974 (N_18974,N_18777,N_18736);
and U18975 (N_18975,N_18697,N_18417);
nand U18976 (N_18976,N_18523,N_18707);
nor U18977 (N_18977,N_18531,N_18478);
or U18978 (N_18978,N_18488,N_18604);
or U18979 (N_18979,N_18740,N_18545);
and U18980 (N_18980,N_18700,N_18494);
and U18981 (N_18981,N_18495,N_18474);
nand U18982 (N_18982,N_18465,N_18670);
nor U18983 (N_18983,N_18564,N_18625);
nor U18984 (N_18984,N_18517,N_18674);
nor U18985 (N_18985,N_18787,N_18480);
nand U18986 (N_18986,N_18429,N_18491);
nand U18987 (N_18987,N_18412,N_18453);
and U18988 (N_18988,N_18645,N_18606);
xnor U18989 (N_18989,N_18497,N_18653);
or U18990 (N_18990,N_18603,N_18557);
nand U18991 (N_18991,N_18690,N_18433);
and U18992 (N_18992,N_18439,N_18600);
xor U18993 (N_18993,N_18717,N_18623);
nand U18994 (N_18994,N_18509,N_18691);
and U18995 (N_18995,N_18405,N_18762);
or U18996 (N_18996,N_18647,N_18665);
or U18997 (N_18997,N_18444,N_18553);
and U18998 (N_18998,N_18672,N_18594);
or U18999 (N_18999,N_18615,N_18742);
or U19000 (N_19000,N_18584,N_18611);
nor U19001 (N_19001,N_18754,N_18658);
xnor U19002 (N_19002,N_18778,N_18727);
nand U19003 (N_19003,N_18712,N_18667);
or U19004 (N_19004,N_18607,N_18596);
and U19005 (N_19005,N_18436,N_18633);
nand U19006 (N_19006,N_18595,N_18565);
or U19007 (N_19007,N_18699,N_18566);
or U19008 (N_19008,N_18702,N_18439);
xnor U19009 (N_19009,N_18427,N_18584);
nor U19010 (N_19010,N_18501,N_18640);
xnor U19011 (N_19011,N_18766,N_18642);
xor U19012 (N_19012,N_18429,N_18592);
or U19013 (N_19013,N_18702,N_18762);
nand U19014 (N_19014,N_18774,N_18685);
nor U19015 (N_19015,N_18509,N_18731);
and U19016 (N_19016,N_18757,N_18428);
xor U19017 (N_19017,N_18556,N_18569);
nor U19018 (N_19018,N_18596,N_18563);
and U19019 (N_19019,N_18725,N_18670);
and U19020 (N_19020,N_18537,N_18591);
xor U19021 (N_19021,N_18406,N_18506);
nand U19022 (N_19022,N_18735,N_18612);
nor U19023 (N_19023,N_18471,N_18560);
nor U19024 (N_19024,N_18524,N_18653);
nand U19025 (N_19025,N_18751,N_18470);
nand U19026 (N_19026,N_18739,N_18715);
and U19027 (N_19027,N_18682,N_18754);
nor U19028 (N_19028,N_18775,N_18515);
nor U19029 (N_19029,N_18630,N_18458);
or U19030 (N_19030,N_18623,N_18732);
and U19031 (N_19031,N_18499,N_18753);
nor U19032 (N_19032,N_18756,N_18450);
or U19033 (N_19033,N_18497,N_18768);
nor U19034 (N_19034,N_18687,N_18733);
nor U19035 (N_19035,N_18594,N_18425);
nor U19036 (N_19036,N_18553,N_18638);
or U19037 (N_19037,N_18425,N_18740);
xor U19038 (N_19038,N_18725,N_18775);
nand U19039 (N_19039,N_18672,N_18582);
and U19040 (N_19040,N_18655,N_18568);
nor U19041 (N_19041,N_18596,N_18652);
nand U19042 (N_19042,N_18424,N_18736);
nand U19043 (N_19043,N_18713,N_18543);
nor U19044 (N_19044,N_18737,N_18583);
xor U19045 (N_19045,N_18524,N_18753);
nand U19046 (N_19046,N_18513,N_18724);
or U19047 (N_19047,N_18504,N_18472);
or U19048 (N_19048,N_18501,N_18403);
and U19049 (N_19049,N_18417,N_18423);
and U19050 (N_19050,N_18618,N_18720);
nand U19051 (N_19051,N_18434,N_18525);
or U19052 (N_19052,N_18569,N_18453);
xnor U19053 (N_19053,N_18758,N_18606);
and U19054 (N_19054,N_18492,N_18470);
and U19055 (N_19055,N_18723,N_18673);
nand U19056 (N_19056,N_18516,N_18755);
and U19057 (N_19057,N_18473,N_18616);
nand U19058 (N_19058,N_18427,N_18698);
xnor U19059 (N_19059,N_18525,N_18661);
nor U19060 (N_19060,N_18767,N_18780);
nor U19061 (N_19061,N_18790,N_18472);
nand U19062 (N_19062,N_18495,N_18750);
nor U19063 (N_19063,N_18648,N_18749);
nor U19064 (N_19064,N_18773,N_18557);
xor U19065 (N_19065,N_18731,N_18685);
and U19066 (N_19066,N_18459,N_18623);
nor U19067 (N_19067,N_18748,N_18646);
and U19068 (N_19068,N_18759,N_18502);
xor U19069 (N_19069,N_18755,N_18552);
nand U19070 (N_19070,N_18468,N_18693);
and U19071 (N_19071,N_18712,N_18736);
nor U19072 (N_19072,N_18437,N_18429);
nor U19073 (N_19073,N_18607,N_18548);
or U19074 (N_19074,N_18751,N_18654);
nand U19075 (N_19075,N_18680,N_18745);
nand U19076 (N_19076,N_18744,N_18753);
and U19077 (N_19077,N_18564,N_18553);
nor U19078 (N_19078,N_18549,N_18484);
xor U19079 (N_19079,N_18730,N_18629);
or U19080 (N_19080,N_18750,N_18570);
nand U19081 (N_19081,N_18523,N_18562);
nor U19082 (N_19082,N_18731,N_18581);
and U19083 (N_19083,N_18548,N_18708);
xor U19084 (N_19084,N_18774,N_18443);
and U19085 (N_19085,N_18562,N_18599);
nor U19086 (N_19086,N_18458,N_18571);
xnor U19087 (N_19087,N_18574,N_18552);
nand U19088 (N_19088,N_18680,N_18453);
nand U19089 (N_19089,N_18513,N_18700);
xnor U19090 (N_19090,N_18633,N_18492);
nor U19091 (N_19091,N_18546,N_18520);
nand U19092 (N_19092,N_18412,N_18763);
or U19093 (N_19093,N_18650,N_18678);
or U19094 (N_19094,N_18582,N_18645);
or U19095 (N_19095,N_18440,N_18748);
or U19096 (N_19096,N_18499,N_18400);
nand U19097 (N_19097,N_18657,N_18559);
xor U19098 (N_19098,N_18415,N_18571);
xor U19099 (N_19099,N_18528,N_18591);
nand U19100 (N_19100,N_18652,N_18439);
and U19101 (N_19101,N_18536,N_18403);
and U19102 (N_19102,N_18779,N_18485);
nand U19103 (N_19103,N_18763,N_18509);
nor U19104 (N_19104,N_18619,N_18482);
nand U19105 (N_19105,N_18428,N_18459);
or U19106 (N_19106,N_18467,N_18502);
xnor U19107 (N_19107,N_18419,N_18601);
and U19108 (N_19108,N_18608,N_18554);
nand U19109 (N_19109,N_18573,N_18420);
nor U19110 (N_19110,N_18590,N_18410);
nand U19111 (N_19111,N_18404,N_18611);
xnor U19112 (N_19112,N_18633,N_18724);
nor U19113 (N_19113,N_18687,N_18636);
nor U19114 (N_19114,N_18451,N_18442);
xor U19115 (N_19115,N_18564,N_18659);
or U19116 (N_19116,N_18543,N_18795);
xor U19117 (N_19117,N_18606,N_18781);
nand U19118 (N_19118,N_18507,N_18717);
nor U19119 (N_19119,N_18636,N_18620);
and U19120 (N_19120,N_18781,N_18436);
or U19121 (N_19121,N_18767,N_18635);
nor U19122 (N_19122,N_18677,N_18497);
xor U19123 (N_19123,N_18471,N_18659);
nor U19124 (N_19124,N_18402,N_18529);
xor U19125 (N_19125,N_18586,N_18613);
or U19126 (N_19126,N_18472,N_18770);
nor U19127 (N_19127,N_18436,N_18730);
and U19128 (N_19128,N_18645,N_18792);
or U19129 (N_19129,N_18587,N_18711);
nor U19130 (N_19130,N_18788,N_18699);
nor U19131 (N_19131,N_18655,N_18714);
nor U19132 (N_19132,N_18755,N_18571);
xnor U19133 (N_19133,N_18597,N_18460);
xnor U19134 (N_19134,N_18670,N_18726);
or U19135 (N_19135,N_18540,N_18515);
xor U19136 (N_19136,N_18789,N_18402);
nand U19137 (N_19137,N_18560,N_18788);
xnor U19138 (N_19138,N_18527,N_18540);
xnor U19139 (N_19139,N_18698,N_18704);
and U19140 (N_19140,N_18510,N_18593);
xnor U19141 (N_19141,N_18483,N_18430);
and U19142 (N_19142,N_18443,N_18403);
xnor U19143 (N_19143,N_18426,N_18666);
nand U19144 (N_19144,N_18592,N_18407);
nand U19145 (N_19145,N_18453,N_18458);
nand U19146 (N_19146,N_18777,N_18701);
xor U19147 (N_19147,N_18407,N_18441);
and U19148 (N_19148,N_18497,N_18500);
xnor U19149 (N_19149,N_18735,N_18554);
and U19150 (N_19150,N_18740,N_18646);
or U19151 (N_19151,N_18699,N_18516);
or U19152 (N_19152,N_18637,N_18666);
nor U19153 (N_19153,N_18743,N_18685);
nor U19154 (N_19154,N_18504,N_18476);
nor U19155 (N_19155,N_18630,N_18772);
nand U19156 (N_19156,N_18623,N_18747);
xnor U19157 (N_19157,N_18425,N_18678);
nand U19158 (N_19158,N_18761,N_18655);
nor U19159 (N_19159,N_18759,N_18740);
nand U19160 (N_19160,N_18598,N_18553);
xor U19161 (N_19161,N_18683,N_18720);
nor U19162 (N_19162,N_18411,N_18562);
and U19163 (N_19163,N_18650,N_18586);
nand U19164 (N_19164,N_18763,N_18494);
nand U19165 (N_19165,N_18592,N_18687);
or U19166 (N_19166,N_18562,N_18727);
nand U19167 (N_19167,N_18413,N_18505);
and U19168 (N_19168,N_18576,N_18521);
xnor U19169 (N_19169,N_18412,N_18627);
and U19170 (N_19170,N_18407,N_18731);
xnor U19171 (N_19171,N_18464,N_18777);
and U19172 (N_19172,N_18701,N_18499);
and U19173 (N_19173,N_18794,N_18498);
and U19174 (N_19174,N_18607,N_18528);
nand U19175 (N_19175,N_18698,N_18534);
or U19176 (N_19176,N_18584,N_18718);
nor U19177 (N_19177,N_18767,N_18415);
nor U19178 (N_19178,N_18424,N_18585);
nor U19179 (N_19179,N_18711,N_18404);
nand U19180 (N_19180,N_18781,N_18723);
nor U19181 (N_19181,N_18461,N_18651);
nor U19182 (N_19182,N_18777,N_18501);
xor U19183 (N_19183,N_18567,N_18532);
and U19184 (N_19184,N_18773,N_18559);
and U19185 (N_19185,N_18568,N_18631);
xor U19186 (N_19186,N_18414,N_18611);
xnor U19187 (N_19187,N_18551,N_18734);
xnor U19188 (N_19188,N_18547,N_18560);
and U19189 (N_19189,N_18423,N_18468);
nor U19190 (N_19190,N_18486,N_18474);
and U19191 (N_19191,N_18436,N_18539);
nand U19192 (N_19192,N_18455,N_18661);
xor U19193 (N_19193,N_18522,N_18460);
and U19194 (N_19194,N_18584,N_18775);
xnor U19195 (N_19195,N_18505,N_18427);
nand U19196 (N_19196,N_18613,N_18469);
nand U19197 (N_19197,N_18457,N_18676);
and U19198 (N_19198,N_18402,N_18581);
or U19199 (N_19199,N_18543,N_18704);
and U19200 (N_19200,N_18901,N_19158);
and U19201 (N_19201,N_19169,N_18819);
nand U19202 (N_19202,N_19061,N_19025);
nand U19203 (N_19203,N_18868,N_18908);
xnor U19204 (N_19204,N_18900,N_18934);
nor U19205 (N_19205,N_18814,N_19083);
nor U19206 (N_19206,N_19167,N_18966);
or U19207 (N_19207,N_19133,N_18969);
nor U19208 (N_19208,N_19106,N_18957);
or U19209 (N_19209,N_18986,N_19073);
and U19210 (N_19210,N_18983,N_19148);
nand U19211 (N_19211,N_19130,N_18919);
xnor U19212 (N_19212,N_18939,N_19132);
xor U19213 (N_19213,N_18841,N_19194);
nor U19214 (N_19214,N_19165,N_18977);
or U19215 (N_19215,N_18857,N_19175);
nor U19216 (N_19216,N_19003,N_18816);
and U19217 (N_19217,N_18802,N_18932);
nand U19218 (N_19218,N_19191,N_19096);
xnor U19219 (N_19219,N_18850,N_19118);
nand U19220 (N_19220,N_19173,N_18898);
nor U19221 (N_19221,N_19015,N_19182);
nor U19222 (N_19222,N_18876,N_18935);
or U19223 (N_19223,N_19028,N_18884);
or U19224 (N_19224,N_19070,N_18829);
nand U19225 (N_19225,N_19052,N_18834);
nor U19226 (N_19226,N_19026,N_19049);
nand U19227 (N_19227,N_18922,N_18897);
nor U19228 (N_19228,N_19050,N_18989);
nor U19229 (N_19229,N_18862,N_18980);
nand U19230 (N_19230,N_19105,N_19045);
xor U19231 (N_19231,N_18863,N_18998);
or U19232 (N_19232,N_19195,N_18886);
xnor U19233 (N_19233,N_19150,N_18889);
nor U19234 (N_19234,N_19102,N_19024);
xor U19235 (N_19235,N_18993,N_18811);
nor U19236 (N_19236,N_18856,N_19019);
nand U19237 (N_19237,N_19198,N_19099);
and U19238 (N_19238,N_19186,N_18975);
nor U19239 (N_19239,N_19031,N_18847);
or U19240 (N_19240,N_18895,N_19101);
nor U19241 (N_19241,N_18818,N_18849);
xor U19242 (N_19242,N_18842,N_19016);
nor U19243 (N_19243,N_18823,N_19170);
or U19244 (N_19244,N_19190,N_19141);
nor U19245 (N_19245,N_18858,N_18833);
xnor U19246 (N_19246,N_18815,N_18910);
nand U19247 (N_19247,N_18881,N_19153);
or U19248 (N_19248,N_19059,N_18888);
xor U19249 (N_19249,N_19154,N_18978);
nand U19250 (N_19250,N_18896,N_18882);
and U19251 (N_19251,N_19104,N_19172);
xnor U19252 (N_19252,N_19076,N_19152);
and U19253 (N_19253,N_19164,N_18880);
nand U19254 (N_19254,N_18912,N_18808);
nor U19255 (N_19255,N_18955,N_19111);
nand U19256 (N_19256,N_19184,N_19072);
nor U19257 (N_19257,N_19007,N_18916);
or U19258 (N_19258,N_19174,N_19149);
and U19259 (N_19259,N_19185,N_19146);
or U19260 (N_19260,N_19008,N_19095);
and U19261 (N_19261,N_18931,N_19183);
nor U19262 (N_19262,N_19004,N_18801);
and U19263 (N_19263,N_19188,N_19121);
xnor U19264 (N_19264,N_18893,N_18873);
nor U19265 (N_19265,N_19078,N_18942);
nor U19266 (N_19266,N_19035,N_18928);
xor U19267 (N_19267,N_19068,N_19001);
or U19268 (N_19268,N_18949,N_18970);
nand U19269 (N_19269,N_19138,N_18920);
and U19270 (N_19270,N_18930,N_19017);
xor U19271 (N_19271,N_18953,N_18813);
or U19272 (N_19272,N_18902,N_18956);
xor U19273 (N_19273,N_19089,N_18810);
nor U19274 (N_19274,N_18804,N_19043);
nand U19275 (N_19275,N_19145,N_18954);
nor U19276 (N_19276,N_18806,N_18911);
nor U19277 (N_19277,N_18883,N_19077);
xor U19278 (N_19278,N_18965,N_19088);
xnor U19279 (N_19279,N_19042,N_18860);
nor U19280 (N_19280,N_18952,N_18994);
nor U19281 (N_19281,N_18803,N_19038);
nor U19282 (N_19282,N_19115,N_19181);
and U19283 (N_19283,N_18821,N_19196);
nand U19284 (N_19284,N_18878,N_18976);
xnor U19285 (N_19285,N_18947,N_18997);
and U19286 (N_19286,N_18971,N_19166);
nand U19287 (N_19287,N_19087,N_19143);
nand U19288 (N_19288,N_19081,N_19147);
xor U19289 (N_19289,N_18865,N_19039);
nor U19290 (N_19290,N_18830,N_18864);
or U19291 (N_19291,N_19009,N_18915);
nor U19292 (N_19292,N_19180,N_18996);
nand U19293 (N_19293,N_18959,N_19041);
or U19294 (N_19294,N_18924,N_19063);
nor U19295 (N_19295,N_19018,N_18923);
nand U19296 (N_19296,N_18807,N_18872);
xor U19297 (N_19297,N_18972,N_19137);
nand U19298 (N_19298,N_19090,N_18974);
xor U19299 (N_19299,N_19192,N_19048);
or U19300 (N_19300,N_18995,N_18874);
nor U19301 (N_19301,N_19162,N_19054);
xor U19302 (N_19302,N_19020,N_18824);
nor U19303 (N_19303,N_18867,N_18914);
nand U19304 (N_19304,N_19051,N_19062);
xnor U19305 (N_19305,N_19125,N_19069);
and U19306 (N_19306,N_18979,N_19010);
xnor U19307 (N_19307,N_18960,N_19021);
nor U19308 (N_19308,N_19123,N_18946);
or U19309 (N_19309,N_19189,N_18866);
or U19310 (N_19310,N_19122,N_18987);
nor U19311 (N_19311,N_19114,N_18812);
nor U19312 (N_19312,N_18875,N_18940);
and U19313 (N_19313,N_19056,N_18909);
xnor U19314 (N_19314,N_19168,N_19040);
nor U19315 (N_19315,N_19079,N_19187);
or U19316 (N_19316,N_19064,N_18904);
or U19317 (N_19317,N_18926,N_18870);
or U19318 (N_19318,N_18905,N_18852);
and U19319 (N_19319,N_19134,N_18846);
nor U19320 (N_19320,N_18948,N_19053);
xnor U19321 (N_19321,N_18853,N_19109);
or U19322 (N_19322,N_18973,N_18885);
xor U19323 (N_19323,N_19177,N_19080);
or U19324 (N_19324,N_18961,N_18929);
nor U19325 (N_19325,N_18871,N_18851);
or U19326 (N_19326,N_19058,N_18907);
nand U19327 (N_19327,N_18837,N_18950);
or U19328 (N_19328,N_19107,N_18985);
nor U19329 (N_19329,N_19176,N_19171);
nor U19330 (N_19330,N_18887,N_19030);
or U19331 (N_19331,N_19097,N_18982);
nand U19332 (N_19332,N_18831,N_19000);
or U19333 (N_19333,N_19098,N_19159);
xnor U19334 (N_19334,N_19012,N_18861);
nor U19335 (N_19335,N_18917,N_19011);
and U19336 (N_19336,N_19140,N_18877);
and U19337 (N_19337,N_18828,N_19112);
or U19338 (N_19338,N_18951,N_19074);
nand U19339 (N_19339,N_18990,N_19108);
nor U19340 (N_19340,N_19093,N_19091);
nor U19341 (N_19341,N_18927,N_18820);
xnor U19342 (N_19342,N_19193,N_19065);
nor U19343 (N_19343,N_18817,N_18967);
nand U19344 (N_19344,N_19144,N_19199);
nand U19345 (N_19345,N_19027,N_19047);
and U19346 (N_19346,N_19155,N_19117);
nand U19347 (N_19347,N_18991,N_19151);
nor U19348 (N_19348,N_18822,N_18906);
or U19349 (N_19349,N_18968,N_18869);
nor U19350 (N_19350,N_19094,N_18809);
nor U19351 (N_19351,N_18944,N_19135);
nor U19352 (N_19352,N_19055,N_19002);
and U19353 (N_19353,N_18843,N_19163);
nand U19354 (N_19354,N_19005,N_18839);
nor U19355 (N_19355,N_18826,N_18936);
nor U19356 (N_19356,N_19128,N_18992);
or U19357 (N_19357,N_18962,N_19029);
or U19358 (N_19358,N_19179,N_19082);
or U19359 (N_19359,N_18892,N_18943);
xnor U19360 (N_19360,N_19100,N_18918);
xor U19361 (N_19361,N_18999,N_18899);
or U19362 (N_19362,N_18925,N_19129);
nor U19363 (N_19363,N_19127,N_19131);
nand U19364 (N_19364,N_18945,N_18981);
nor U19365 (N_19365,N_19075,N_19119);
or U19366 (N_19366,N_19142,N_19197);
and U19367 (N_19367,N_19103,N_18984);
or U19368 (N_19368,N_18921,N_18835);
nand U19369 (N_19369,N_18879,N_19067);
and U19370 (N_19370,N_19034,N_19092);
nand U19371 (N_19371,N_19046,N_19178);
and U19372 (N_19372,N_18913,N_19116);
and U19373 (N_19373,N_19057,N_19037);
and U19374 (N_19374,N_19156,N_18933);
nor U19375 (N_19375,N_18832,N_18891);
and U19376 (N_19376,N_18838,N_18825);
and U19377 (N_19377,N_18827,N_19084);
nor U19378 (N_19378,N_19124,N_18941);
xnor U19379 (N_19379,N_18845,N_18848);
and U19380 (N_19380,N_19161,N_18938);
xor U19381 (N_19381,N_19036,N_19120);
nand U19382 (N_19382,N_19113,N_18800);
or U19383 (N_19383,N_18894,N_18958);
and U19384 (N_19384,N_19014,N_19157);
or U19385 (N_19385,N_19086,N_19033);
nand U19386 (N_19386,N_19023,N_18855);
nand U19387 (N_19387,N_18854,N_18859);
nand U19388 (N_19388,N_18840,N_18890);
or U19389 (N_19389,N_18836,N_19160);
nor U19390 (N_19390,N_18844,N_19032);
and U19391 (N_19391,N_19022,N_19066);
nor U19392 (N_19392,N_19071,N_19013);
xnor U19393 (N_19393,N_18988,N_18805);
and U19394 (N_19394,N_19110,N_18937);
nand U19395 (N_19395,N_19126,N_19044);
xor U19396 (N_19396,N_19060,N_19139);
nor U19397 (N_19397,N_19006,N_18964);
nand U19398 (N_19398,N_18963,N_19085);
and U19399 (N_19399,N_18903,N_19136);
or U19400 (N_19400,N_18926,N_19146);
and U19401 (N_19401,N_19079,N_18930);
nor U19402 (N_19402,N_18931,N_19078);
xnor U19403 (N_19403,N_19147,N_18992);
xnor U19404 (N_19404,N_18914,N_18988);
and U19405 (N_19405,N_19081,N_18846);
nor U19406 (N_19406,N_19136,N_18889);
nand U19407 (N_19407,N_18834,N_18967);
and U19408 (N_19408,N_18982,N_18937);
or U19409 (N_19409,N_18966,N_19076);
xor U19410 (N_19410,N_18957,N_19012);
nand U19411 (N_19411,N_19168,N_19098);
xnor U19412 (N_19412,N_19066,N_18960);
xor U19413 (N_19413,N_19104,N_19194);
or U19414 (N_19414,N_19179,N_18891);
nor U19415 (N_19415,N_19031,N_18917);
and U19416 (N_19416,N_18904,N_18888);
and U19417 (N_19417,N_19084,N_19171);
nand U19418 (N_19418,N_19186,N_18907);
xnor U19419 (N_19419,N_19060,N_19064);
nand U19420 (N_19420,N_19073,N_18908);
or U19421 (N_19421,N_18944,N_19027);
xor U19422 (N_19422,N_18912,N_18862);
xor U19423 (N_19423,N_19190,N_18954);
xnor U19424 (N_19424,N_19079,N_19114);
nor U19425 (N_19425,N_19061,N_18871);
nand U19426 (N_19426,N_19046,N_19154);
xor U19427 (N_19427,N_19005,N_18942);
or U19428 (N_19428,N_19066,N_18984);
nor U19429 (N_19429,N_19058,N_19096);
and U19430 (N_19430,N_19026,N_18849);
xnor U19431 (N_19431,N_18887,N_18916);
nor U19432 (N_19432,N_19171,N_19024);
and U19433 (N_19433,N_19088,N_19078);
or U19434 (N_19434,N_19140,N_19099);
and U19435 (N_19435,N_19134,N_19055);
nand U19436 (N_19436,N_18955,N_18884);
nand U19437 (N_19437,N_18812,N_18924);
or U19438 (N_19438,N_19024,N_18815);
and U19439 (N_19439,N_18885,N_18803);
and U19440 (N_19440,N_19166,N_18957);
xor U19441 (N_19441,N_18853,N_18945);
or U19442 (N_19442,N_19074,N_19057);
xnor U19443 (N_19443,N_19016,N_19186);
nand U19444 (N_19444,N_18889,N_18965);
xnor U19445 (N_19445,N_19138,N_18815);
or U19446 (N_19446,N_18825,N_18868);
and U19447 (N_19447,N_18990,N_19099);
nand U19448 (N_19448,N_18990,N_18971);
or U19449 (N_19449,N_18871,N_19133);
and U19450 (N_19450,N_19164,N_19014);
or U19451 (N_19451,N_19097,N_19148);
xor U19452 (N_19452,N_18945,N_18801);
xnor U19453 (N_19453,N_19028,N_19019);
nor U19454 (N_19454,N_19158,N_19113);
and U19455 (N_19455,N_18823,N_18848);
xor U19456 (N_19456,N_19184,N_18815);
or U19457 (N_19457,N_19001,N_18995);
nand U19458 (N_19458,N_19008,N_19190);
and U19459 (N_19459,N_18953,N_19111);
or U19460 (N_19460,N_19065,N_18809);
nand U19461 (N_19461,N_19172,N_19131);
xor U19462 (N_19462,N_19162,N_18935);
nand U19463 (N_19463,N_18912,N_18876);
or U19464 (N_19464,N_19058,N_18978);
nor U19465 (N_19465,N_19055,N_19121);
and U19466 (N_19466,N_19067,N_18884);
or U19467 (N_19467,N_18915,N_19162);
or U19468 (N_19468,N_19162,N_18936);
or U19469 (N_19469,N_18801,N_18948);
xnor U19470 (N_19470,N_19193,N_18852);
and U19471 (N_19471,N_19049,N_19004);
xnor U19472 (N_19472,N_19007,N_18847);
nor U19473 (N_19473,N_18863,N_18876);
xor U19474 (N_19474,N_18976,N_19116);
nor U19475 (N_19475,N_18848,N_19139);
and U19476 (N_19476,N_19110,N_18845);
nor U19477 (N_19477,N_18914,N_19152);
or U19478 (N_19478,N_19021,N_19153);
or U19479 (N_19479,N_18987,N_19158);
nand U19480 (N_19480,N_18987,N_18942);
nor U19481 (N_19481,N_18955,N_18886);
or U19482 (N_19482,N_18843,N_18872);
or U19483 (N_19483,N_18820,N_19092);
and U19484 (N_19484,N_19068,N_18892);
nand U19485 (N_19485,N_18854,N_19108);
or U19486 (N_19486,N_18811,N_18918);
nor U19487 (N_19487,N_19029,N_18849);
nor U19488 (N_19488,N_18946,N_19118);
xnor U19489 (N_19489,N_19048,N_19050);
xor U19490 (N_19490,N_19146,N_19138);
and U19491 (N_19491,N_18975,N_18965);
and U19492 (N_19492,N_18885,N_18999);
xnor U19493 (N_19493,N_18900,N_19052);
xor U19494 (N_19494,N_18996,N_18852);
and U19495 (N_19495,N_18963,N_19093);
nand U19496 (N_19496,N_18860,N_19059);
nand U19497 (N_19497,N_19134,N_18961);
nand U19498 (N_19498,N_19072,N_18904);
xnor U19499 (N_19499,N_18948,N_19025);
and U19500 (N_19500,N_19063,N_19177);
xor U19501 (N_19501,N_18941,N_18931);
and U19502 (N_19502,N_18881,N_18996);
nor U19503 (N_19503,N_19119,N_19104);
and U19504 (N_19504,N_18864,N_19094);
or U19505 (N_19505,N_18883,N_18976);
nand U19506 (N_19506,N_18837,N_18851);
and U19507 (N_19507,N_19046,N_18978);
and U19508 (N_19508,N_18934,N_19023);
nand U19509 (N_19509,N_19045,N_18805);
nor U19510 (N_19510,N_18823,N_19062);
or U19511 (N_19511,N_19069,N_19126);
or U19512 (N_19512,N_18968,N_18949);
nor U19513 (N_19513,N_18929,N_18974);
nor U19514 (N_19514,N_18969,N_19129);
nor U19515 (N_19515,N_18935,N_18879);
nor U19516 (N_19516,N_19140,N_18937);
and U19517 (N_19517,N_18952,N_18893);
or U19518 (N_19518,N_18877,N_18862);
and U19519 (N_19519,N_19088,N_19017);
or U19520 (N_19520,N_19137,N_18865);
or U19521 (N_19521,N_18827,N_19188);
nor U19522 (N_19522,N_19050,N_18912);
xnor U19523 (N_19523,N_18817,N_19032);
or U19524 (N_19524,N_19064,N_18895);
or U19525 (N_19525,N_18995,N_19162);
and U19526 (N_19526,N_18991,N_19045);
and U19527 (N_19527,N_19106,N_18966);
nor U19528 (N_19528,N_18811,N_19176);
xnor U19529 (N_19529,N_19099,N_19155);
xnor U19530 (N_19530,N_19035,N_19027);
nand U19531 (N_19531,N_18944,N_19138);
nand U19532 (N_19532,N_19112,N_18993);
nor U19533 (N_19533,N_18964,N_19048);
nand U19534 (N_19534,N_19064,N_18884);
xnor U19535 (N_19535,N_18966,N_18837);
nor U19536 (N_19536,N_18972,N_18958);
xnor U19537 (N_19537,N_18942,N_19140);
nor U19538 (N_19538,N_19177,N_18873);
or U19539 (N_19539,N_18841,N_18927);
or U19540 (N_19540,N_18832,N_18997);
nor U19541 (N_19541,N_19048,N_18900);
nor U19542 (N_19542,N_19019,N_19157);
or U19543 (N_19543,N_18922,N_18953);
and U19544 (N_19544,N_19004,N_19147);
or U19545 (N_19545,N_18875,N_19030);
nor U19546 (N_19546,N_19036,N_18888);
xnor U19547 (N_19547,N_18932,N_19115);
and U19548 (N_19548,N_19044,N_19124);
nand U19549 (N_19549,N_19128,N_18870);
xnor U19550 (N_19550,N_18885,N_18958);
xor U19551 (N_19551,N_18956,N_18801);
nor U19552 (N_19552,N_19110,N_19033);
nand U19553 (N_19553,N_19161,N_18918);
nor U19554 (N_19554,N_19177,N_19123);
nand U19555 (N_19555,N_18928,N_19121);
nand U19556 (N_19556,N_19050,N_18988);
and U19557 (N_19557,N_18804,N_19136);
xnor U19558 (N_19558,N_19143,N_18892);
nand U19559 (N_19559,N_19009,N_18920);
nand U19560 (N_19560,N_18962,N_18948);
nand U19561 (N_19561,N_19179,N_19135);
xnor U19562 (N_19562,N_18958,N_18819);
or U19563 (N_19563,N_18810,N_19184);
xnor U19564 (N_19564,N_19155,N_19184);
and U19565 (N_19565,N_19056,N_18904);
xor U19566 (N_19566,N_19181,N_19065);
xor U19567 (N_19567,N_19113,N_19124);
and U19568 (N_19568,N_18846,N_18952);
nor U19569 (N_19569,N_18982,N_18975);
and U19570 (N_19570,N_19103,N_19044);
and U19571 (N_19571,N_19074,N_19160);
nor U19572 (N_19572,N_18907,N_19056);
or U19573 (N_19573,N_18864,N_19086);
nand U19574 (N_19574,N_19031,N_19109);
or U19575 (N_19575,N_18913,N_18827);
xnor U19576 (N_19576,N_18818,N_18899);
and U19577 (N_19577,N_18805,N_18836);
nand U19578 (N_19578,N_19184,N_18992);
xnor U19579 (N_19579,N_19160,N_19064);
and U19580 (N_19580,N_19129,N_18997);
or U19581 (N_19581,N_18987,N_18823);
xnor U19582 (N_19582,N_19022,N_19000);
nand U19583 (N_19583,N_19061,N_18890);
nor U19584 (N_19584,N_19119,N_19089);
nor U19585 (N_19585,N_19128,N_18985);
nand U19586 (N_19586,N_19150,N_19056);
and U19587 (N_19587,N_18856,N_19137);
and U19588 (N_19588,N_18974,N_19136);
nand U19589 (N_19589,N_18903,N_18909);
or U19590 (N_19590,N_18911,N_19010);
xor U19591 (N_19591,N_19025,N_19185);
nand U19592 (N_19592,N_19169,N_19122);
nand U19593 (N_19593,N_19121,N_18946);
and U19594 (N_19594,N_18839,N_19015);
xor U19595 (N_19595,N_18846,N_18843);
nand U19596 (N_19596,N_18960,N_19045);
or U19597 (N_19597,N_19022,N_19097);
and U19598 (N_19598,N_19067,N_19138);
nor U19599 (N_19599,N_19051,N_18929);
nor U19600 (N_19600,N_19207,N_19303);
or U19601 (N_19601,N_19427,N_19435);
xor U19602 (N_19602,N_19379,N_19281);
nand U19603 (N_19603,N_19422,N_19497);
xor U19604 (N_19604,N_19211,N_19239);
and U19605 (N_19605,N_19584,N_19486);
nand U19606 (N_19606,N_19515,N_19592);
xnor U19607 (N_19607,N_19595,N_19276);
nand U19608 (N_19608,N_19439,N_19569);
nand U19609 (N_19609,N_19254,N_19394);
nor U19610 (N_19610,N_19321,N_19540);
xnor U19611 (N_19611,N_19307,N_19457);
nand U19612 (N_19612,N_19443,N_19252);
nand U19613 (N_19613,N_19258,N_19598);
and U19614 (N_19614,N_19524,N_19314);
or U19615 (N_19615,N_19347,N_19375);
xor U19616 (N_19616,N_19361,N_19348);
nor U19617 (N_19617,N_19465,N_19277);
nor U19618 (N_19618,N_19514,N_19417);
nand U19619 (N_19619,N_19248,N_19449);
nor U19620 (N_19620,N_19519,N_19520);
xor U19621 (N_19621,N_19311,N_19237);
or U19622 (N_19622,N_19392,N_19505);
or U19623 (N_19623,N_19345,N_19201);
nand U19624 (N_19624,N_19489,N_19358);
xnor U19625 (N_19625,N_19401,N_19460);
nor U19626 (N_19626,N_19441,N_19330);
nor U19627 (N_19627,N_19442,N_19426);
xor U19628 (N_19628,N_19255,N_19571);
xnor U19629 (N_19629,N_19354,N_19395);
or U19630 (N_19630,N_19472,N_19455);
nor U19631 (N_19631,N_19333,N_19283);
and U19632 (N_19632,N_19591,N_19549);
xnor U19633 (N_19633,N_19499,N_19225);
nor U19634 (N_19634,N_19240,N_19493);
nand U19635 (N_19635,N_19300,N_19544);
or U19636 (N_19636,N_19272,N_19495);
nand U19637 (N_19637,N_19336,N_19326);
or U19638 (N_19638,N_19398,N_19387);
nand U19639 (N_19639,N_19425,N_19205);
nand U19640 (N_19640,N_19257,N_19391);
nand U19641 (N_19641,N_19535,N_19492);
nand U19642 (N_19642,N_19464,N_19301);
or U19643 (N_19643,N_19586,N_19378);
or U19644 (N_19644,N_19561,N_19341);
xor U19645 (N_19645,N_19230,N_19485);
or U19646 (N_19646,N_19452,N_19528);
or U19647 (N_19647,N_19318,N_19253);
or U19648 (N_19648,N_19367,N_19434);
and U19649 (N_19649,N_19344,N_19288);
nor U19650 (N_19650,N_19545,N_19218);
and U19651 (N_19651,N_19558,N_19384);
or U19652 (N_19652,N_19407,N_19305);
nand U19653 (N_19653,N_19403,N_19278);
and U19654 (N_19654,N_19555,N_19510);
and U19655 (N_19655,N_19374,N_19414);
and U19656 (N_19656,N_19372,N_19292);
and U19657 (N_19657,N_19491,N_19597);
nand U19658 (N_19658,N_19547,N_19376);
and U19659 (N_19659,N_19355,N_19212);
xor U19660 (N_19660,N_19568,N_19327);
nand U19661 (N_19661,N_19266,N_19263);
or U19662 (N_19662,N_19578,N_19506);
and U19663 (N_19663,N_19533,N_19313);
and U19664 (N_19664,N_19260,N_19550);
nand U19665 (N_19665,N_19328,N_19484);
nor U19666 (N_19666,N_19477,N_19593);
or U19667 (N_19667,N_19294,N_19329);
and U19668 (N_19668,N_19397,N_19575);
nand U19669 (N_19669,N_19279,N_19476);
nor U19670 (N_19670,N_19388,N_19436);
xnor U19671 (N_19671,N_19390,N_19302);
or U19672 (N_19672,N_19286,N_19536);
nand U19673 (N_19673,N_19501,N_19356);
nand U19674 (N_19674,N_19352,N_19461);
or U19675 (N_19675,N_19487,N_19264);
xor U19676 (N_19676,N_19368,N_19440);
nor U19677 (N_19677,N_19382,N_19249);
xor U19678 (N_19678,N_19469,N_19265);
nor U19679 (N_19679,N_19463,N_19430);
nand U19680 (N_19680,N_19518,N_19413);
xnor U19681 (N_19681,N_19418,N_19468);
nand U19682 (N_19682,N_19583,N_19581);
and U19683 (N_19683,N_19498,N_19538);
xor U19684 (N_19684,N_19360,N_19325);
nand U19685 (N_19685,N_19516,N_19227);
nand U19686 (N_19686,N_19529,N_19589);
and U19687 (N_19687,N_19339,N_19428);
nor U19688 (N_19688,N_19511,N_19206);
nor U19689 (N_19689,N_19539,N_19331);
and U19690 (N_19690,N_19251,N_19503);
nand U19691 (N_19691,N_19373,N_19215);
nand U19692 (N_19692,N_19433,N_19412);
or U19693 (N_19693,N_19396,N_19399);
or U19694 (N_19694,N_19351,N_19259);
nor U19695 (N_19695,N_19445,N_19210);
nor U19696 (N_19696,N_19308,N_19274);
nor U19697 (N_19697,N_19480,N_19243);
nor U19698 (N_19698,N_19228,N_19590);
nand U19699 (N_19699,N_19411,N_19381);
or U19700 (N_19700,N_19234,N_19543);
or U19701 (N_19701,N_19562,N_19365);
xor U19702 (N_19702,N_19599,N_19342);
nor U19703 (N_19703,N_19517,N_19319);
xnor U19704 (N_19704,N_19291,N_19221);
nand U19705 (N_19705,N_19542,N_19566);
xnor U19706 (N_19706,N_19316,N_19389);
xnor U19707 (N_19707,N_19541,N_19500);
xor U19708 (N_19708,N_19438,N_19408);
nand U19709 (N_19709,N_19548,N_19502);
nor U19710 (N_19710,N_19304,N_19450);
nor U19711 (N_19711,N_19467,N_19369);
nor U19712 (N_19712,N_19315,N_19245);
nor U19713 (N_19713,N_19534,N_19377);
nor U19714 (N_19714,N_19559,N_19474);
or U19715 (N_19715,N_19431,N_19312);
nand U19716 (N_19716,N_19479,N_19322);
nand U19717 (N_19717,N_19563,N_19262);
nand U19718 (N_19718,N_19564,N_19223);
and U19719 (N_19719,N_19466,N_19522);
xnor U19720 (N_19720,N_19587,N_19523);
or U19721 (N_19721,N_19437,N_19432);
or U19722 (N_19722,N_19456,N_19579);
and U19723 (N_19723,N_19483,N_19448);
xnor U19724 (N_19724,N_19573,N_19481);
nor U19725 (N_19725,N_19216,N_19268);
nor U19726 (N_19726,N_19309,N_19349);
nand U19727 (N_19727,N_19400,N_19530);
and U19728 (N_19728,N_19409,N_19335);
and U19729 (N_19729,N_19200,N_19370);
nand U19730 (N_19730,N_19393,N_19214);
nor U19731 (N_19731,N_19423,N_19494);
or U19732 (N_19732,N_19273,N_19531);
or U19733 (N_19733,N_19299,N_19509);
or U19734 (N_19734,N_19596,N_19585);
or U19735 (N_19735,N_19306,N_19235);
nor U19736 (N_19736,N_19203,N_19453);
and U19737 (N_19737,N_19363,N_19204);
and U19738 (N_19738,N_19537,N_19527);
xor U19739 (N_19739,N_19482,N_19250);
nand U19740 (N_19740,N_19582,N_19220);
nor U19741 (N_19741,N_19416,N_19462);
nand U19742 (N_19742,N_19324,N_19310);
and U19743 (N_19743,N_19280,N_19219);
or U19744 (N_19744,N_19429,N_19421);
xor U19745 (N_19745,N_19317,N_19554);
xnor U19746 (N_19746,N_19565,N_19267);
and U19747 (N_19747,N_19553,N_19246);
and U19748 (N_19748,N_19525,N_19405);
nand U19749 (N_19749,N_19385,N_19357);
nor U19750 (N_19750,N_19337,N_19512);
or U19751 (N_19751,N_19383,N_19298);
and U19752 (N_19752,N_19572,N_19570);
and U19753 (N_19753,N_19295,N_19580);
or U19754 (N_19754,N_19446,N_19334);
nand U19755 (N_19755,N_19320,N_19366);
and U19756 (N_19756,N_19289,N_19232);
nor U19757 (N_19757,N_19475,N_19271);
xor U19758 (N_19758,N_19594,N_19415);
xnor U19759 (N_19759,N_19242,N_19222);
xnor U19760 (N_19760,N_19419,N_19386);
xnor U19761 (N_19761,N_19567,N_19241);
or U19762 (N_19762,N_19444,N_19451);
and U19763 (N_19763,N_19380,N_19224);
or U19764 (N_19764,N_19209,N_19346);
nor U19765 (N_19765,N_19261,N_19454);
nand U19766 (N_19766,N_19217,N_19546);
nor U19767 (N_19767,N_19473,N_19532);
nor U19768 (N_19768,N_19496,N_19447);
or U19769 (N_19769,N_19371,N_19213);
nor U19770 (N_19770,N_19247,N_19290);
nor U19771 (N_19771,N_19362,N_19275);
and U19772 (N_19772,N_19424,N_19420);
nor U19773 (N_19773,N_19574,N_19208);
nor U19774 (N_19774,N_19282,N_19285);
nor U19775 (N_19775,N_19233,N_19521);
and U19776 (N_19776,N_19478,N_19338);
or U19777 (N_19777,N_19340,N_19552);
and U19778 (N_19778,N_19490,N_19560);
and U19779 (N_19779,N_19470,N_19364);
xnor U19780 (N_19780,N_19332,N_19577);
nand U19781 (N_19781,N_19556,N_19526);
or U19782 (N_19782,N_19269,N_19353);
xnor U19783 (N_19783,N_19244,N_19323);
nor U19784 (N_19784,N_19588,N_19350);
xnor U19785 (N_19785,N_19229,N_19270);
and U19786 (N_19786,N_19557,N_19202);
or U19787 (N_19787,N_19284,N_19404);
nand U19788 (N_19788,N_19504,N_19236);
and U19789 (N_19789,N_19459,N_19513);
nor U19790 (N_19790,N_19402,N_19458);
or U19791 (N_19791,N_19359,N_19410);
or U19792 (N_19792,N_19508,N_19296);
or U19793 (N_19793,N_19256,N_19551);
xor U19794 (N_19794,N_19406,N_19488);
nor U19795 (N_19795,N_19238,N_19226);
or U19796 (N_19796,N_19507,N_19297);
xor U19797 (N_19797,N_19231,N_19293);
nor U19798 (N_19798,N_19287,N_19576);
xor U19799 (N_19799,N_19343,N_19471);
or U19800 (N_19800,N_19469,N_19331);
xor U19801 (N_19801,N_19308,N_19520);
xnor U19802 (N_19802,N_19436,N_19367);
or U19803 (N_19803,N_19452,N_19394);
nor U19804 (N_19804,N_19428,N_19511);
nand U19805 (N_19805,N_19431,N_19570);
and U19806 (N_19806,N_19289,N_19488);
xnor U19807 (N_19807,N_19226,N_19547);
nor U19808 (N_19808,N_19551,N_19426);
nor U19809 (N_19809,N_19412,N_19532);
or U19810 (N_19810,N_19400,N_19376);
nor U19811 (N_19811,N_19449,N_19316);
and U19812 (N_19812,N_19474,N_19380);
and U19813 (N_19813,N_19218,N_19537);
nor U19814 (N_19814,N_19210,N_19443);
xnor U19815 (N_19815,N_19563,N_19550);
or U19816 (N_19816,N_19252,N_19380);
xnor U19817 (N_19817,N_19507,N_19482);
xnor U19818 (N_19818,N_19303,N_19355);
or U19819 (N_19819,N_19481,N_19291);
or U19820 (N_19820,N_19483,N_19336);
or U19821 (N_19821,N_19528,N_19467);
nand U19822 (N_19822,N_19231,N_19322);
or U19823 (N_19823,N_19445,N_19515);
and U19824 (N_19824,N_19357,N_19380);
xor U19825 (N_19825,N_19217,N_19240);
xnor U19826 (N_19826,N_19418,N_19236);
or U19827 (N_19827,N_19456,N_19446);
xor U19828 (N_19828,N_19578,N_19270);
and U19829 (N_19829,N_19347,N_19200);
and U19830 (N_19830,N_19526,N_19243);
nand U19831 (N_19831,N_19281,N_19365);
and U19832 (N_19832,N_19528,N_19317);
and U19833 (N_19833,N_19287,N_19414);
xor U19834 (N_19834,N_19573,N_19544);
nor U19835 (N_19835,N_19217,N_19504);
nand U19836 (N_19836,N_19458,N_19366);
or U19837 (N_19837,N_19231,N_19387);
nand U19838 (N_19838,N_19289,N_19357);
nand U19839 (N_19839,N_19306,N_19342);
nor U19840 (N_19840,N_19591,N_19203);
and U19841 (N_19841,N_19597,N_19527);
nor U19842 (N_19842,N_19542,N_19444);
xnor U19843 (N_19843,N_19285,N_19224);
xnor U19844 (N_19844,N_19244,N_19379);
nor U19845 (N_19845,N_19288,N_19442);
nand U19846 (N_19846,N_19393,N_19286);
nand U19847 (N_19847,N_19340,N_19208);
xnor U19848 (N_19848,N_19451,N_19265);
nand U19849 (N_19849,N_19543,N_19279);
and U19850 (N_19850,N_19582,N_19288);
nor U19851 (N_19851,N_19201,N_19327);
or U19852 (N_19852,N_19468,N_19337);
nor U19853 (N_19853,N_19266,N_19236);
and U19854 (N_19854,N_19412,N_19408);
and U19855 (N_19855,N_19285,N_19502);
nor U19856 (N_19856,N_19236,N_19496);
or U19857 (N_19857,N_19378,N_19232);
or U19858 (N_19858,N_19210,N_19474);
nand U19859 (N_19859,N_19404,N_19206);
nand U19860 (N_19860,N_19306,N_19478);
xnor U19861 (N_19861,N_19577,N_19518);
nand U19862 (N_19862,N_19473,N_19336);
nand U19863 (N_19863,N_19288,N_19468);
nand U19864 (N_19864,N_19503,N_19435);
nand U19865 (N_19865,N_19585,N_19506);
xnor U19866 (N_19866,N_19433,N_19554);
nor U19867 (N_19867,N_19306,N_19459);
nor U19868 (N_19868,N_19236,N_19262);
xor U19869 (N_19869,N_19281,N_19566);
nor U19870 (N_19870,N_19551,N_19472);
or U19871 (N_19871,N_19580,N_19395);
and U19872 (N_19872,N_19208,N_19300);
nand U19873 (N_19873,N_19333,N_19404);
xnor U19874 (N_19874,N_19512,N_19475);
or U19875 (N_19875,N_19545,N_19328);
nor U19876 (N_19876,N_19482,N_19406);
and U19877 (N_19877,N_19384,N_19529);
and U19878 (N_19878,N_19482,N_19481);
xor U19879 (N_19879,N_19511,N_19346);
nor U19880 (N_19880,N_19226,N_19391);
or U19881 (N_19881,N_19433,N_19246);
or U19882 (N_19882,N_19409,N_19206);
or U19883 (N_19883,N_19383,N_19504);
nand U19884 (N_19884,N_19232,N_19478);
nor U19885 (N_19885,N_19314,N_19276);
nor U19886 (N_19886,N_19342,N_19412);
nand U19887 (N_19887,N_19365,N_19269);
nor U19888 (N_19888,N_19216,N_19528);
and U19889 (N_19889,N_19579,N_19566);
nor U19890 (N_19890,N_19266,N_19447);
nor U19891 (N_19891,N_19479,N_19436);
and U19892 (N_19892,N_19276,N_19299);
xnor U19893 (N_19893,N_19262,N_19374);
xor U19894 (N_19894,N_19529,N_19292);
nor U19895 (N_19895,N_19518,N_19260);
nor U19896 (N_19896,N_19589,N_19404);
nand U19897 (N_19897,N_19577,N_19246);
nand U19898 (N_19898,N_19349,N_19297);
nor U19899 (N_19899,N_19361,N_19401);
or U19900 (N_19900,N_19322,N_19313);
nand U19901 (N_19901,N_19577,N_19230);
or U19902 (N_19902,N_19419,N_19467);
nand U19903 (N_19903,N_19567,N_19496);
nor U19904 (N_19904,N_19513,N_19304);
nand U19905 (N_19905,N_19587,N_19467);
nor U19906 (N_19906,N_19366,N_19446);
nand U19907 (N_19907,N_19556,N_19365);
nand U19908 (N_19908,N_19542,N_19350);
and U19909 (N_19909,N_19489,N_19319);
nand U19910 (N_19910,N_19512,N_19218);
or U19911 (N_19911,N_19428,N_19458);
xnor U19912 (N_19912,N_19374,N_19443);
xnor U19913 (N_19913,N_19500,N_19588);
nand U19914 (N_19914,N_19577,N_19361);
or U19915 (N_19915,N_19224,N_19243);
and U19916 (N_19916,N_19348,N_19449);
and U19917 (N_19917,N_19563,N_19496);
nand U19918 (N_19918,N_19467,N_19344);
xnor U19919 (N_19919,N_19329,N_19533);
and U19920 (N_19920,N_19483,N_19278);
nand U19921 (N_19921,N_19486,N_19430);
xor U19922 (N_19922,N_19293,N_19306);
nor U19923 (N_19923,N_19219,N_19541);
nor U19924 (N_19924,N_19521,N_19268);
nand U19925 (N_19925,N_19256,N_19320);
nor U19926 (N_19926,N_19270,N_19561);
and U19927 (N_19927,N_19458,N_19374);
nand U19928 (N_19928,N_19376,N_19391);
or U19929 (N_19929,N_19263,N_19400);
nand U19930 (N_19930,N_19333,N_19366);
nor U19931 (N_19931,N_19435,N_19321);
nor U19932 (N_19932,N_19470,N_19518);
or U19933 (N_19933,N_19583,N_19366);
and U19934 (N_19934,N_19249,N_19512);
nand U19935 (N_19935,N_19489,N_19477);
nand U19936 (N_19936,N_19399,N_19446);
or U19937 (N_19937,N_19294,N_19240);
nand U19938 (N_19938,N_19452,N_19210);
nor U19939 (N_19939,N_19269,N_19375);
or U19940 (N_19940,N_19456,N_19410);
or U19941 (N_19941,N_19223,N_19295);
xor U19942 (N_19942,N_19209,N_19385);
nor U19943 (N_19943,N_19504,N_19211);
and U19944 (N_19944,N_19404,N_19493);
nor U19945 (N_19945,N_19289,N_19361);
nor U19946 (N_19946,N_19476,N_19596);
nand U19947 (N_19947,N_19481,N_19415);
xnor U19948 (N_19948,N_19352,N_19293);
and U19949 (N_19949,N_19417,N_19304);
nor U19950 (N_19950,N_19275,N_19239);
nor U19951 (N_19951,N_19533,N_19410);
nor U19952 (N_19952,N_19367,N_19331);
nand U19953 (N_19953,N_19205,N_19440);
xnor U19954 (N_19954,N_19392,N_19289);
and U19955 (N_19955,N_19292,N_19293);
or U19956 (N_19956,N_19349,N_19243);
nor U19957 (N_19957,N_19384,N_19565);
nand U19958 (N_19958,N_19249,N_19398);
nor U19959 (N_19959,N_19498,N_19460);
and U19960 (N_19960,N_19265,N_19206);
nor U19961 (N_19961,N_19367,N_19534);
or U19962 (N_19962,N_19596,N_19599);
or U19963 (N_19963,N_19338,N_19441);
or U19964 (N_19964,N_19590,N_19215);
nand U19965 (N_19965,N_19561,N_19583);
nand U19966 (N_19966,N_19539,N_19354);
nor U19967 (N_19967,N_19409,N_19492);
nor U19968 (N_19968,N_19588,N_19585);
nor U19969 (N_19969,N_19500,N_19312);
and U19970 (N_19970,N_19242,N_19408);
xor U19971 (N_19971,N_19509,N_19540);
nor U19972 (N_19972,N_19310,N_19234);
nand U19973 (N_19973,N_19484,N_19488);
nand U19974 (N_19974,N_19350,N_19473);
or U19975 (N_19975,N_19483,N_19527);
nand U19976 (N_19976,N_19538,N_19319);
nor U19977 (N_19977,N_19547,N_19225);
nand U19978 (N_19978,N_19375,N_19533);
nand U19979 (N_19979,N_19511,N_19463);
xnor U19980 (N_19980,N_19474,N_19311);
and U19981 (N_19981,N_19203,N_19248);
xnor U19982 (N_19982,N_19579,N_19266);
and U19983 (N_19983,N_19263,N_19315);
and U19984 (N_19984,N_19549,N_19302);
and U19985 (N_19985,N_19363,N_19504);
and U19986 (N_19986,N_19440,N_19306);
or U19987 (N_19987,N_19541,N_19354);
and U19988 (N_19988,N_19223,N_19257);
nand U19989 (N_19989,N_19530,N_19271);
nor U19990 (N_19990,N_19481,N_19450);
nor U19991 (N_19991,N_19418,N_19353);
xor U19992 (N_19992,N_19424,N_19555);
xnor U19993 (N_19993,N_19388,N_19459);
and U19994 (N_19994,N_19453,N_19304);
nor U19995 (N_19995,N_19550,N_19493);
nor U19996 (N_19996,N_19558,N_19504);
and U19997 (N_19997,N_19580,N_19313);
and U19998 (N_19998,N_19200,N_19395);
and U19999 (N_19999,N_19200,N_19401);
and UO_0 (O_0,N_19914,N_19671);
or UO_1 (O_1,N_19611,N_19768);
or UO_2 (O_2,N_19635,N_19825);
nor UO_3 (O_3,N_19636,N_19723);
nor UO_4 (O_4,N_19837,N_19986);
nor UO_5 (O_5,N_19661,N_19776);
nand UO_6 (O_6,N_19948,N_19988);
nand UO_7 (O_7,N_19769,N_19619);
nor UO_8 (O_8,N_19958,N_19873);
and UO_9 (O_9,N_19838,N_19628);
and UO_10 (O_10,N_19775,N_19884);
or UO_11 (O_11,N_19657,N_19889);
xnor UO_12 (O_12,N_19650,N_19814);
or UO_13 (O_13,N_19966,N_19708);
nor UO_14 (O_14,N_19920,N_19836);
xnor UO_15 (O_15,N_19679,N_19941);
or UO_16 (O_16,N_19917,N_19688);
or UO_17 (O_17,N_19716,N_19706);
nand UO_18 (O_18,N_19753,N_19692);
and UO_19 (O_19,N_19784,N_19990);
and UO_20 (O_20,N_19796,N_19739);
and UO_21 (O_21,N_19842,N_19911);
nand UO_22 (O_22,N_19809,N_19841);
and UO_23 (O_23,N_19861,N_19789);
nand UO_24 (O_24,N_19823,N_19655);
or UO_25 (O_25,N_19924,N_19746);
nand UO_26 (O_26,N_19699,N_19890);
xnor UO_27 (O_27,N_19742,N_19811);
and UO_28 (O_28,N_19799,N_19980);
nor UO_29 (O_29,N_19759,N_19881);
nand UO_30 (O_30,N_19639,N_19664);
and UO_31 (O_31,N_19645,N_19749);
nor UO_32 (O_32,N_19646,N_19850);
xor UO_33 (O_33,N_19955,N_19909);
and UO_34 (O_34,N_19745,N_19950);
xor UO_35 (O_35,N_19731,N_19854);
xor UO_36 (O_36,N_19694,N_19963);
and UO_37 (O_37,N_19906,N_19703);
and UO_38 (O_38,N_19886,N_19615);
nand UO_39 (O_39,N_19621,N_19818);
or UO_40 (O_40,N_19905,N_19761);
xnor UO_41 (O_41,N_19620,N_19701);
and UO_42 (O_42,N_19808,N_19943);
nand UO_43 (O_43,N_19868,N_19665);
or UO_44 (O_44,N_19855,N_19649);
and UO_45 (O_45,N_19623,N_19616);
nor UO_46 (O_46,N_19942,N_19627);
nand UO_47 (O_47,N_19816,N_19912);
or UO_48 (O_48,N_19953,N_19826);
nor UO_49 (O_49,N_19751,N_19788);
xor UO_50 (O_50,N_19651,N_19896);
nor UO_51 (O_51,N_19954,N_19964);
or UO_52 (O_52,N_19669,N_19951);
nor UO_53 (O_53,N_19853,N_19702);
or UO_54 (O_54,N_19726,N_19780);
nand UO_55 (O_55,N_19656,N_19767);
or UO_56 (O_56,N_19613,N_19936);
or UO_57 (O_57,N_19972,N_19847);
or UO_58 (O_58,N_19949,N_19893);
xor UO_59 (O_59,N_19633,N_19778);
and UO_60 (O_60,N_19935,N_19790);
nor UO_61 (O_61,N_19845,N_19987);
nor UO_62 (O_62,N_19762,N_19965);
nor UO_63 (O_63,N_19741,N_19857);
xor UO_64 (O_64,N_19604,N_19737);
and UO_65 (O_65,N_19607,N_19773);
nand UO_66 (O_66,N_19766,N_19887);
or UO_67 (O_67,N_19642,N_19791);
nand UO_68 (O_68,N_19760,N_19974);
nand UO_69 (O_69,N_19998,N_19698);
nor UO_70 (O_70,N_19872,N_19653);
or UO_71 (O_71,N_19786,N_19680);
and UO_72 (O_72,N_19637,N_19844);
xor UO_73 (O_73,N_19795,N_19687);
nor UO_74 (O_74,N_19644,N_19812);
and UO_75 (O_75,N_19971,N_19970);
or UO_76 (O_76,N_19967,N_19711);
nor UO_77 (O_77,N_19713,N_19659);
and UO_78 (O_78,N_19922,N_19710);
and UO_79 (O_79,N_19982,N_19682);
nor UO_80 (O_80,N_19923,N_19876);
nor UO_81 (O_81,N_19629,N_19793);
and UO_82 (O_82,N_19928,N_19654);
nand UO_83 (O_83,N_19984,N_19678);
nand UO_84 (O_84,N_19758,N_19681);
nor UO_85 (O_85,N_19901,N_19744);
nand UO_86 (O_86,N_19973,N_19631);
nand UO_87 (O_87,N_19763,N_19968);
nand UO_88 (O_88,N_19648,N_19719);
nand UO_89 (O_89,N_19771,N_19748);
or UO_90 (O_90,N_19691,N_19938);
or UO_91 (O_91,N_19632,N_19675);
nand UO_92 (O_92,N_19772,N_19902);
or UO_93 (O_93,N_19714,N_19672);
and UO_94 (O_94,N_19625,N_19765);
nand UO_95 (O_95,N_19940,N_19848);
nor UO_96 (O_96,N_19819,N_19601);
xnor UO_97 (O_97,N_19874,N_19722);
nor UO_98 (O_98,N_19695,N_19666);
nor UO_99 (O_99,N_19618,N_19652);
xor UO_100 (O_100,N_19870,N_19820);
nand UO_101 (O_101,N_19730,N_19851);
nor UO_102 (O_102,N_19658,N_19801);
and UO_103 (O_103,N_19718,N_19932);
or UO_104 (O_104,N_19693,N_19794);
xor UO_105 (O_105,N_19704,N_19662);
nor UO_106 (O_106,N_19724,N_19921);
nor UO_107 (O_107,N_19946,N_19858);
or UO_108 (O_108,N_19833,N_19999);
and UO_109 (O_109,N_19898,N_19700);
or UO_110 (O_110,N_19805,N_19840);
nand UO_111 (O_111,N_19899,N_19734);
or UO_112 (O_112,N_19736,N_19959);
or UO_113 (O_113,N_19600,N_19830);
or UO_114 (O_114,N_19919,N_19609);
or UO_115 (O_115,N_19685,N_19931);
xnor UO_116 (O_116,N_19952,N_19978);
or UO_117 (O_117,N_19747,N_19683);
or UO_118 (O_118,N_19866,N_19994);
and UO_119 (O_119,N_19864,N_19879);
xnor UO_120 (O_120,N_19624,N_19933);
or UO_121 (O_121,N_19908,N_19783);
or UO_122 (O_122,N_19750,N_19832);
nor UO_123 (O_123,N_19829,N_19641);
xor UO_124 (O_124,N_19843,N_19960);
xor UO_125 (O_125,N_19839,N_19690);
xor UO_126 (O_126,N_19725,N_19862);
or UO_127 (O_127,N_19782,N_19663);
or UO_128 (O_128,N_19673,N_19989);
nor UO_129 (O_129,N_19860,N_19732);
nand UO_130 (O_130,N_19991,N_19622);
or UO_131 (O_131,N_19797,N_19715);
or UO_132 (O_132,N_19810,N_19913);
nor UO_133 (O_133,N_19821,N_19916);
xor UO_134 (O_134,N_19617,N_19976);
nor UO_135 (O_135,N_19944,N_19712);
nand UO_136 (O_136,N_19785,N_19939);
xor UO_137 (O_137,N_19630,N_19640);
and UO_138 (O_138,N_19817,N_19777);
xnor UO_139 (O_139,N_19754,N_19962);
xnor UO_140 (O_140,N_19910,N_19930);
xnor UO_141 (O_141,N_19674,N_19867);
or UO_142 (O_142,N_19667,N_19875);
nand UO_143 (O_143,N_19869,N_19729);
and UO_144 (O_144,N_19945,N_19883);
nor UO_145 (O_145,N_19787,N_19852);
nand UO_146 (O_146,N_19983,N_19720);
xnor UO_147 (O_147,N_19888,N_19903);
nand UO_148 (O_148,N_19638,N_19705);
and UO_149 (O_149,N_19670,N_19877);
or UO_150 (O_150,N_19668,N_19897);
nor UO_151 (O_151,N_19689,N_19800);
xnor UO_152 (O_152,N_19880,N_19728);
xnor UO_153 (O_153,N_19806,N_19802);
nand UO_154 (O_154,N_19686,N_19781);
or UO_155 (O_155,N_19827,N_19803);
nand UO_156 (O_156,N_19849,N_19756);
nor UO_157 (O_157,N_19798,N_19740);
or UO_158 (O_158,N_19878,N_19774);
nand UO_159 (O_159,N_19915,N_19975);
nor UO_160 (O_160,N_19807,N_19981);
and UO_161 (O_161,N_19634,N_19610);
and UO_162 (O_162,N_19614,N_19996);
nor UO_163 (O_163,N_19907,N_19770);
or UO_164 (O_164,N_19871,N_19643);
nand UO_165 (O_165,N_19697,N_19961);
nand UO_166 (O_166,N_19929,N_19602);
nand UO_167 (O_167,N_19743,N_19997);
or UO_168 (O_168,N_19894,N_19608);
xor UO_169 (O_169,N_19934,N_19733);
and UO_170 (O_170,N_19927,N_19926);
or UO_171 (O_171,N_19605,N_19738);
and UO_172 (O_172,N_19822,N_19835);
nor UO_173 (O_173,N_19992,N_19717);
and UO_174 (O_174,N_19856,N_19885);
or UO_175 (O_175,N_19985,N_19612);
nand UO_176 (O_176,N_19676,N_19834);
or UO_177 (O_177,N_19813,N_19969);
xnor UO_178 (O_178,N_19709,N_19993);
nand UO_179 (O_179,N_19757,N_19831);
nor UO_180 (O_180,N_19696,N_19863);
or UO_181 (O_181,N_19752,N_19995);
nor UO_182 (O_182,N_19937,N_19815);
and UO_183 (O_183,N_19707,N_19824);
and UO_184 (O_184,N_19904,N_19977);
or UO_185 (O_185,N_19684,N_19956);
and UO_186 (O_186,N_19677,N_19647);
xor UO_187 (O_187,N_19882,N_19626);
nand UO_188 (O_188,N_19603,N_19865);
nor UO_189 (O_189,N_19925,N_19900);
xnor UO_190 (O_190,N_19660,N_19957);
xor UO_191 (O_191,N_19892,N_19755);
nor UO_192 (O_192,N_19606,N_19947);
nand UO_193 (O_193,N_19727,N_19828);
nor UO_194 (O_194,N_19804,N_19891);
nor UO_195 (O_195,N_19859,N_19846);
or UO_196 (O_196,N_19721,N_19764);
xnor UO_197 (O_197,N_19979,N_19918);
xor UO_198 (O_198,N_19792,N_19895);
nand UO_199 (O_199,N_19779,N_19735);
xnor UO_200 (O_200,N_19887,N_19600);
nand UO_201 (O_201,N_19672,N_19670);
and UO_202 (O_202,N_19669,N_19619);
or UO_203 (O_203,N_19751,N_19642);
or UO_204 (O_204,N_19733,N_19779);
nand UO_205 (O_205,N_19860,N_19985);
nand UO_206 (O_206,N_19815,N_19953);
nor UO_207 (O_207,N_19950,N_19871);
nand UO_208 (O_208,N_19636,N_19820);
xnor UO_209 (O_209,N_19665,N_19719);
xnor UO_210 (O_210,N_19716,N_19679);
nand UO_211 (O_211,N_19995,N_19608);
and UO_212 (O_212,N_19651,N_19794);
nor UO_213 (O_213,N_19904,N_19818);
xnor UO_214 (O_214,N_19752,N_19743);
xnor UO_215 (O_215,N_19697,N_19767);
nand UO_216 (O_216,N_19667,N_19891);
nand UO_217 (O_217,N_19640,N_19634);
or UO_218 (O_218,N_19745,N_19769);
nor UO_219 (O_219,N_19834,N_19757);
xor UO_220 (O_220,N_19876,N_19976);
xor UO_221 (O_221,N_19933,N_19616);
and UO_222 (O_222,N_19878,N_19885);
or UO_223 (O_223,N_19709,N_19734);
and UO_224 (O_224,N_19899,N_19770);
or UO_225 (O_225,N_19937,N_19881);
and UO_226 (O_226,N_19819,N_19643);
nand UO_227 (O_227,N_19897,N_19855);
nand UO_228 (O_228,N_19972,N_19747);
nand UO_229 (O_229,N_19834,N_19656);
xnor UO_230 (O_230,N_19691,N_19642);
or UO_231 (O_231,N_19699,N_19682);
and UO_232 (O_232,N_19693,N_19849);
nand UO_233 (O_233,N_19775,N_19864);
nor UO_234 (O_234,N_19631,N_19734);
nor UO_235 (O_235,N_19623,N_19948);
nor UO_236 (O_236,N_19724,N_19606);
or UO_237 (O_237,N_19918,N_19631);
nor UO_238 (O_238,N_19924,N_19728);
xnor UO_239 (O_239,N_19805,N_19632);
xnor UO_240 (O_240,N_19913,N_19966);
and UO_241 (O_241,N_19692,N_19918);
xnor UO_242 (O_242,N_19854,N_19786);
and UO_243 (O_243,N_19917,N_19613);
xnor UO_244 (O_244,N_19972,N_19613);
and UO_245 (O_245,N_19857,N_19665);
xnor UO_246 (O_246,N_19718,N_19633);
nand UO_247 (O_247,N_19676,N_19600);
or UO_248 (O_248,N_19832,N_19992);
or UO_249 (O_249,N_19620,N_19771);
nor UO_250 (O_250,N_19938,N_19673);
or UO_251 (O_251,N_19688,N_19979);
nor UO_252 (O_252,N_19733,N_19780);
nor UO_253 (O_253,N_19679,N_19851);
or UO_254 (O_254,N_19959,N_19830);
nand UO_255 (O_255,N_19797,N_19981);
and UO_256 (O_256,N_19930,N_19921);
or UO_257 (O_257,N_19729,N_19932);
and UO_258 (O_258,N_19650,N_19919);
nand UO_259 (O_259,N_19971,N_19796);
or UO_260 (O_260,N_19639,N_19814);
nor UO_261 (O_261,N_19713,N_19707);
or UO_262 (O_262,N_19718,N_19616);
nor UO_263 (O_263,N_19968,N_19704);
xnor UO_264 (O_264,N_19909,N_19918);
xnor UO_265 (O_265,N_19646,N_19729);
and UO_266 (O_266,N_19600,N_19855);
or UO_267 (O_267,N_19799,N_19691);
or UO_268 (O_268,N_19901,N_19829);
or UO_269 (O_269,N_19614,N_19817);
nand UO_270 (O_270,N_19807,N_19888);
and UO_271 (O_271,N_19619,N_19855);
and UO_272 (O_272,N_19862,N_19866);
nor UO_273 (O_273,N_19695,N_19788);
and UO_274 (O_274,N_19884,N_19600);
nor UO_275 (O_275,N_19695,N_19759);
and UO_276 (O_276,N_19738,N_19647);
and UO_277 (O_277,N_19742,N_19785);
xnor UO_278 (O_278,N_19665,N_19729);
or UO_279 (O_279,N_19651,N_19825);
and UO_280 (O_280,N_19964,N_19782);
nor UO_281 (O_281,N_19646,N_19723);
nand UO_282 (O_282,N_19789,N_19691);
or UO_283 (O_283,N_19671,N_19847);
and UO_284 (O_284,N_19883,N_19706);
nor UO_285 (O_285,N_19968,N_19646);
nand UO_286 (O_286,N_19807,N_19731);
nor UO_287 (O_287,N_19622,N_19668);
nor UO_288 (O_288,N_19867,N_19606);
nand UO_289 (O_289,N_19739,N_19681);
or UO_290 (O_290,N_19604,N_19879);
nor UO_291 (O_291,N_19823,N_19905);
nand UO_292 (O_292,N_19890,N_19785);
nor UO_293 (O_293,N_19625,N_19680);
or UO_294 (O_294,N_19659,N_19908);
nand UO_295 (O_295,N_19654,N_19775);
nor UO_296 (O_296,N_19704,N_19806);
nand UO_297 (O_297,N_19720,N_19898);
xnor UO_298 (O_298,N_19747,N_19898);
nand UO_299 (O_299,N_19897,N_19871);
and UO_300 (O_300,N_19839,N_19955);
xor UO_301 (O_301,N_19811,N_19781);
nor UO_302 (O_302,N_19808,N_19942);
xnor UO_303 (O_303,N_19949,N_19931);
nor UO_304 (O_304,N_19985,N_19716);
nand UO_305 (O_305,N_19824,N_19763);
nand UO_306 (O_306,N_19650,N_19810);
nor UO_307 (O_307,N_19996,N_19775);
or UO_308 (O_308,N_19707,N_19884);
and UO_309 (O_309,N_19806,N_19610);
xnor UO_310 (O_310,N_19963,N_19660);
xor UO_311 (O_311,N_19914,N_19651);
and UO_312 (O_312,N_19623,N_19969);
nor UO_313 (O_313,N_19939,N_19622);
and UO_314 (O_314,N_19829,N_19697);
xor UO_315 (O_315,N_19933,N_19975);
nand UO_316 (O_316,N_19708,N_19904);
xnor UO_317 (O_317,N_19665,N_19815);
nand UO_318 (O_318,N_19981,N_19618);
nand UO_319 (O_319,N_19697,N_19652);
or UO_320 (O_320,N_19770,N_19648);
nor UO_321 (O_321,N_19656,N_19940);
xor UO_322 (O_322,N_19867,N_19807);
and UO_323 (O_323,N_19936,N_19809);
nand UO_324 (O_324,N_19653,N_19919);
or UO_325 (O_325,N_19978,N_19690);
nor UO_326 (O_326,N_19988,N_19704);
and UO_327 (O_327,N_19671,N_19748);
nand UO_328 (O_328,N_19860,N_19657);
xnor UO_329 (O_329,N_19845,N_19606);
and UO_330 (O_330,N_19708,N_19897);
and UO_331 (O_331,N_19928,N_19774);
nor UO_332 (O_332,N_19749,N_19795);
or UO_333 (O_333,N_19629,N_19912);
nand UO_334 (O_334,N_19703,N_19892);
nand UO_335 (O_335,N_19755,N_19712);
or UO_336 (O_336,N_19967,N_19746);
and UO_337 (O_337,N_19698,N_19841);
or UO_338 (O_338,N_19810,N_19891);
nand UO_339 (O_339,N_19851,N_19810);
and UO_340 (O_340,N_19864,N_19981);
xor UO_341 (O_341,N_19800,N_19828);
xnor UO_342 (O_342,N_19754,N_19941);
nand UO_343 (O_343,N_19630,N_19712);
nand UO_344 (O_344,N_19986,N_19795);
nor UO_345 (O_345,N_19992,N_19658);
and UO_346 (O_346,N_19687,N_19625);
xor UO_347 (O_347,N_19705,N_19757);
and UO_348 (O_348,N_19671,N_19855);
xnor UO_349 (O_349,N_19963,N_19869);
nor UO_350 (O_350,N_19990,N_19694);
or UO_351 (O_351,N_19945,N_19775);
nor UO_352 (O_352,N_19658,N_19924);
nand UO_353 (O_353,N_19947,N_19814);
and UO_354 (O_354,N_19887,N_19732);
and UO_355 (O_355,N_19662,N_19679);
and UO_356 (O_356,N_19827,N_19764);
nand UO_357 (O_357,N_19856,N_19764);
and UO_358 (O_358,N_19962,N_19615);
nand UO_359 (O_359,N_19995,N_19690);
or UO_360 (O_360,N_19760,N_19710);
nand UO_361 (O_361,N_19828,N_19689);
nor UO_362 (O_362,N_19854,N_19777);
nor UO_363 (O_363,N_19982,N_19968);
nand UO_364 (O_364,N_19881,N_19871);
or UO_365 (O_365,N_19768,N_19686);
and UO_366 (O_366,N_19981,N_19983);
nor UO_367 (O_367,N_19859,N_19936);
nand UO_368 (O_368,N_19757,N_19928);
nor UO_369 (O_369,N_19955,N_19731);
nor UO_370 (O_370,N_19919,N_19811);
xor UO_371 (O_371,N_19991,N_19792);
nor UO_372 (O_372,N_19895,N_19994);
nor UO_373 (O_373,N_19913,N_19910);
nor UO_374 (O_374,N_19725,N_19773);
nand UO_375 (O_375,N_19920,N_19805);
xnor UO_376 (O_376,N_19610,N_19850);
xor UO_377 (O_377,N_19990,N_19896);
nand UO_378 (O_378,N_19696,N_19630);
xnor UO_379 (O_379,N_19821,N_19658);
and UO_380 (O_380,N_19661,N_19872);
or UO_381 (O_381,N_19698,N_19769);
and UO_382 (O_382,N_19615,N_19829);
and UO_383 (O_383,N_19810,N_19653);
or UO_384 (O_384,N_19749,N_19951);
and UO_385 (O_385,N_19697,N_19724);
xnor UO_386 (O_386,N_19652,N_19696);
nand UO_387 (O_387,N_19619,N_19622);
xnor UO_388 (O_388,N_19673,N_19867);
nand UO_389 (O_389,N_19630,N_19816);
nand UO_390 (O_390,N_19957,N_19889);
xnor UO_391 (O_391,N_19826,N_19866);
and UO_392 (O_392,N_19917,N_19777);
and UO_393 (O_393,N_19644,N_19780);
or UO_394 (O_394,N_19902,N_19769);
or UO_395 (O_395,N_19935,N_19926);
xnor UO_396 (O_396,N_19618,N_19794);
and UO_397 (O_397,N_19658,N_19962);
nand UO_398 (O_398,N_19704,N_19631);
xnor UO_399 (O_399,N_19604,N_19697);
and UO_400 (O_400,N_19947,N_19637);
nand UO_401 (O_401,N_19674,N_19851);
and UO_402 (O_402,N_19991,N_19731);
xor UO_403 (O_403,N_19709,N_19977);
nor UO_404 (O_404,N_19946,N_19925);
and UO_405 (O_405,N_19647,N_19695);
and UO_406 (O_406,N_19856,N_19931);
and UO_407 (O_407,N_19924,N_19731);
nand UO_408 (O_408,N_19640,N_19636);
and UO_409 (O_409,N_19679,N_19974);
and UO_410 (O_410,N_19636,N_19713);
and UO_411 (O_411,N_19773,N_19861);
xor UO_412 (O_412,N_19803,N_19974);
and UO_413 (O_413,N_19862,N_19819);
and UO_414 (O_414,N_19993,N_19884);
or UO_415 (O_415,N_19750,N_19679);
xnor UO_416 (O_416,N_19804,N_19643);
and UO_417 (O_417,N_19858,N_19940);
or UO_418 (O_418,N_19901,N_19802);
and UO_419 (O_419,N_19727,N_19897);
or UO_420 (O_420,N_19600,N_19900);
nand UO_421 (O_421,N_19678,N_19831);
and UO_422 (O_422,N_19688,N_19900);
nor UO_423 (O_423,N_19747,N_19823);
and UO_424 (O_424,N_19715,N_19823);
and UO_425 (O_425,N_19639,N_19633);
nand UO_426 (O_426,N_19930,N_19627);
and UO_427 (O_427,N_19828,N_19928);
nor UO_428 (O_428,N_19683,N_19911);
nand UO_429 (O_429,N_19701,N_19826);
xnor UO_430 (O_430,N_19637,N_19806);
nand UO_431 (O_431,N_19765,N_19827);
and UO_432 (O_432,N_19646,N_19654);
nor UO_433 (O_433,N_19815,N_19983);
nand UO_434 (O_434,N_19618,N_19666);
nor UO_435 (O_435,N_19950,N_19729);
nand UO_436 (O_436,N_19673,N_19873);
or UO_437 (O_437,N_19969,N_19684);
nor UO_438 (O_438,N_19741,N_19854);
xor UO_439 (O_439,N_19873,N_19878);
and UO_440 (O_440,N_19767,N_19894);
xor UO_441 (O_441,N_19682,N_19994);
or UO_442 (O_442,N_19877,N_19917);
nor UO_443 (O_443,N_19708,N_19611);
or UO_444 (O_444,N_19991,N_19763);
and UO_445 (O_445,N_19811,N_19821);
nor UO_446 (O_446,N_19864,N_19661);
xor UO_447 (O_447,N_19707,N_19918);
nor UO_448 (O_448,N_19868,N_19869);
or UO_449 (O_449,N_19902,N_19778);
and UO_450 (O_450,N_19947,N_19611);
or UO_451 (O_451,N_19648,N_19980);
xnor UO_452 (O_452,N_19844,N_19859);
and UO_453 (O_453,N_19885,N_19615);
nand UO_454 (O_454,N_19660,N_19867);
nand UO_455 (O_455,N_19868,N_19721);
xnor UO_456 (O_456,N_19738,N_19603);
nor UO_457 (O_457,N_19810,N_19973);
nand UO_458 (O_458,N_19690,N_19744);
nand UO_459 (O_459,N_19772,N_19603);
and UO_460 (O_460,N_19843,N_19833);
nor UO_461 (O_461,N_19787,N_19767);
xnor UO_462 (O_462,N_19682,N_19833);
nor UO_463 (O_463,N_19951,N_19883);
or UO_464 (O_464,N_19658,N_19965);
xnor UO_465 (O_465,N_19856,N_19714);
and UO_466 (O_466,N_19928,N_19740);
nor UO_467 (O_467,N_19959,N_19895);
xnor UO_468 (O_468,N_19702,N_19641);
and UO_469 (O_469,N_19641,N_19989);
and UO_470 (O_470,N_19932,N_19724);
and UO_471 (O_471,N_19722,N_19962);
nand UO_472 (O_472,N_19945,N_19634);
nor UO_473 (O_473,N_19633,N_19807);
nor UO_474 (O_474,N_19628,N_19742);
nand UO_475 (O_475,N_19971,N_19892);
nor UO_476 (O_476,N_19679,N_19821);
xor UO_477 (O_477,N_19791,N_19994);
or UO_478 (O_478,N_19977,N_19874);
nor UO_479 (O_479,N_19844,N_19797);
nor UO_480 (O_480,N_19626,N_19718);
nand UO_481 (O_481,N_19683,N_19969);
or UO_482 (O_482,N_19651,N_19964);
nor UO_483 (O_483,N_19914,N_19769);
or UO_484 (O_484,N_19601,N_19637);
xnor UO_485 (O_485,N_19803,N_19854);
nand UO_486 (O_486,N_19824,N_19612);
nand UO_487 (O_487,N_19686,N_19982);
and UO_488 (O_488,N_19651,N_19968);
nor UO_489 (O_489,N_19604,N_19646);
xor UO_490 (O_490,N_19819,N_19901);
xor UO_491 (O_491,N_19824,N_19942);
or UO_492 (O_492,N_19675,N_19789);
or UO_493 (O_493,N_19866,N_19886);
nand UO_494 (O_494,N_19846,N_19681);
and UO_495 (O_495,N_19698,N_19669);
xnor UO_496 (O_496,N_19996,N_19768);
and UO_497 (O_497,N_19833,N_19625);
nand UO_498 (O_498,N_19935,N_19818);
or UO_499 (O_499,N_19969,N_19999);
and UO_500 (O_500,N_19654,N_19681);
and UO_501 (O_501,N_19609,N_19657);
and UO_502 (O_502,N_19615,N_19673);
xor UO_503 (O_503,N_19671,N_19689);
or UO_504 (O_504,N_19700,N_19920);
and UO_505 (O_505,N_19945,N_19968);
or UO_506 (O_506,N_19977,N_19656);
nand UO_507 (O_507,N_19652,N_19722);
and UO_508 (O_508,N_19898,N_19851);
nor UO_509 (O_509,N_19865,N_19721);
and UO_510 (O_510,N_19792,N_19617);
nand UO_511 (O_511,N_19611,N_19660);
and UO_512 (O_512,N_19730,N_19971);
nand UO_513 (O_513,N_19766,N_19828);
or UO_514 (O_514,N_19822,N_19745);
nand UO_515 (O_515,N_19791,N_19630);
and UO_516 (O_516,N_19723,N_19866);
and UO_517 (O_517,N_19649,N_19788);
nor UO_518 (O_518,N_19714,N_19802);
or UO_519 (O_519,N_19886,N_19671);
xor UO_520 (O_520,N_19703,N_19990);
xnor UO_521 (O_521,N_19614,N_19929);
and UO_522 (O_522,N_19751,N_19738);
and UO_523 (O_523,N_19949,N_19790);
or UO_524 (O_524,N_19670,N_19826);
nor UO_525 (O_525,N_19870,N_19805);
and UO_526 (O_526,N_19769,N_19689);
xor UO_527 (O_527,N_19686,N_19627);
or UO_528 (O_528,N_19811,N_19884);
xor UO_529 (O_529,N_19736,N_19965);
nor UO_530 (O_530,N_19655,N_19867);
xor UO_531 (O_531,N_19940,N_19939);
nand UO_532 (O_532,N_19938,N_19908);
xor UO_533 (O_533,N_19948,N_19740);
xnor UO_534 (O_534,N_19982,N_19612);
nand UO_535 (O_535,N_19930,N_19787);
nor UO_536 (O_536,N_19805,N_19828);
nand UO_537 (O_537,N_19625,N_19630);
and UO_538 (O_538,N_19770,N_19857);
or UO_539 (O_539,N_19797,N_19850);
xnor UO_540 (O_540,N_19756,N_19843);
or UO_541 (O_541,N_19704,N_19789);
nand UO_542 (O_542,N_19862,N_19680);
xnor UO_543 (O_543,N_19802,N_19602);
and UO_544 (O_544,N_19698,N_19688);
nor UO_545 (O_545,N_19686,N_19747);
nand UO_546 (O_546,N_19783,N_19645);
or UO_547 (O_547,N_19953,N_19944);
xor UO_548 (O_548,N_19926,N_19756);
and UO_549 (O_549,N_19710,N_19891);
nor UO_550 (O_550,N_19719,N_19623);
and UO_551 (O_551,N_19951,N_19907);
and UO_552 (O_552,N_19973,N_19951);
nor UO_553 (O_553,N_19734,N_19811);
xor UO_554 (O_554,N_19738,N_19846);
and UO_555 (O_555,N_19833,N_19732);
nand UO_556 (O_556,N_19671,N_19754);
and UO_557 (O_557,N_19732,N_19675);
nand UO_558 (O_558,N_19748,N_19741);
nand UO_559 (O_559,N_19965,N_19613);
nor UO_560 (O_560,N_19652,N_19690);
nor UO_561 (O_561,N_19806,N_19811);
nand UO_562 (O_562,N_19859,N_19832);
nor UO_563 (O_563,N_19699,N_19737);
or UO_564 (O_564,N_19852,N_19716);
xor UO_565 (O_565,N_19874,N_19800);
nand UO_566 (O_566,N_19663,N_19893);
and UO_567 (O_567,N_19685,N_19759);
nor UO_568 (O_568,N_19996,N_19860);
nand UO_569 (O_569,N_19923,N_19899);
nand UO_570 (O_570,N_19915,N_19679);
or UO_571 (O_571,N_19772,N_19878);
nand UO_572 (O_572,N_19642,N_19832);
nand UO_573 (O_573,N_19909,N_19688);
xnor UO_574 (O_574,N_19724,N_19774);
xnor UO_575 (O_575,N_19867,N_19648);
xnor UO_576 (O_576,N_19898,N_19975);
or UO_577 (O_577,N_19956,N_19937);
nor UO_578 (O_578,N_19843,N_19941);
or UO_579 (O_579,N_19852,N_19913);
nand UO_580 (O_580,N_19994,N_19673);
nor UO_581 (O_581,N_19688,N_19866);
nand UO_582 (O_582,N_19825,N_19804);
nor UO_583 (O_583,N_19673,N_19761);
xor UO_584 (O_584,N_19755,N_19763);
nand UO_585 (O_585,N_19634,N_19832);
or UO_586 (O_586,N_19955,N_19993);
or UO_587 (O_587,N_19811,N_19676);
and UO_588 (O_588,N_19811,N_19715);
nor UO_589 (O_589,N_19839,N_19628);
or UO_590 (O_590,N_19729,N_19990);
and UO_591 (O_591,N_19890,N_19805);
nand UO_592 (O_592,N_19688,N_19862);
or UO_593 (O_593,N_19688,N_19804);
nor UO_594 (O_594,N_19665,N_19943);
xnor UO_595 (O_595,N_19755,N_19727);
or UO_596 (O_596,N_19914,N_19606);
or UO_597 (O_597,N_19961,N_19672);
nor UO_598 (O_598,N_19875,N_19701);
nor UO_599 (O_599,N_19987,N_19894);
nor UO_600 (O_600,N_19830,N_19929);
nand UO_601 (O_601,N_19879,N_19836);
or UO_602 (O_602,N_19602,N_19644);
nor UO_603 (O_603,N_19874,N_19952);
and UO_604 (O_604,N_19799,N_19908);
nand UO_605 (O_605,N_19880,N_19976);
or UO_606 (O_606,N_19658,N_19949);
nand UO_607 (O_607,N_19691,N_19958);
and UO_608 (O_608,N_19991,N_19931);
xor UO_609 (O_609,N_19722,N_19800);
nand UO_610 (O_610,N_19770,N_19822);
and UO_611 (O_611,N_19972,N_19986);
or UO_612 (O_612,N_19914,N_19742);
xnor UO_613 (O_613,N_19762,N_19854);
or UO_614 (O_614,N_19641,N_19861);
or UO_615 (O_615,N_19810,N_19637);
and UO_616 (O_616,N_19917,N_19837);
or UO_617 (O_617,N_19802,N_19722);
nand UO_618 (O_618,N_19895,N_19637);
nor UO_619 (O_619,N_19621,N_19976);
nand UO_620 (O_620,N_19929,N_19794);
xnor UO_621 (O_621,N_19968,N_19724);
and UO_622 (O_622,N_19732,N_19662);
nor UO_623 (O_623,N_19825,N_19727);
or UO_624 (O_624,N_19881,N_19884);
nand UO_625 (O_625,N_19664,N_19923);
nor UO_626 (O_626,N_19632,N_19871);
and UO_627 (O_627,N_19888,N_19701);
nand UO_628 (O_628,N_19878,N_19679);
or UO_629 (O_629,N_19924,N_19985);
nor UO_630 (O_630,N_19746,N_19688);
or UO_631 (O_631,N_19664,N_19872);
xor UO_632 (O_632,N_19725,N_19795);
and UO_633 (O_633,N_19602,N_19781);
nor UO_634 (O_634,N_19888,N_19926);
xnor UO_635 (O_635,N_19780,N_19878);
xnor UO_636 (O_636,N_19709,N_19908);
and UO_637 (O_637,N_19831,N_19871);
nor UO_638 (O_638,N_19886,N_19938);
and UO_639 (O_639,N_19955,N_19615);
nor UO_640 (O_640,N_19676,N_19757);
or UO_641 (O_641,N_19822,N_19786);
nand UO_642 (O_642,N_19745,N_19735);
nand UO_643 (O_643,N_19629,N_19861);
nand UO_644 (O_644,N_19847,N_19664);
nand UO_645 (O_645,N_19741,N_19790);
xnor UO_646 (O_646,N_19966,N_19816);
nand UO_647 (O_647,N_19996,N_19731);
nor UO_648 (O_648,N_19735,N_19738);
or UO_649 (O_649,N_19909,N_19846);
or UO_650 (O_650,N_19675,N_19676);
and UO_651 (O_651,N_19752,N_19701);
nand UO_652 (O_652,N_19957,N_19728);
and UO_653 (O_653,N_19883,N_19785);
and UO_654 (O_654,N_19979,N_19770);
or UO_655 (O_655,N_19702,N_19686);
nor UO_656 (O_656,N_19970,N_19698);
nor UO_657 (O_657,N_19701,N_19764);
nand UO_658 (O_658,N_19908,N_19662);
xor UO_659 (O_659,N_19818,N_19996);
and UO_660 (O_660,N_19913,N_19973);
nor UO_661 (O_661,N_19897,N_19910);
nor UO_662 (O_662,N_19853,N_19865);
nand UO_663 (O_663,N_19975,N_19688);
xor UO_664 (O_664,N_19931,N_19601);
and UO_665 (O_665,N_19718,N_19780);
or UO_666 (O_666,N_19964,N_19889);
xor UO_667 (O_667,N_19793,N_19951);
nand UO_668 (O_668,N_19715,N_19710);
xor UO_669 (O_669,N_19937,N_19990);
and UO_670 (O_670,N_19801,N_19680);
or UO_671 (O_671,N_19989,N_19948);
nor UO_672 (O_672,N_19931,N_19701);
and UO_673 (O_673,N_19707,N_19801);
xor UO_674 (O_674,N_19803,N_19713);
nor UO_675 (O_675,N_19769,N_19906);
nor UO_676 (O_676,N_19684,N_19850);
and UO_677 (O_677,N_19754,N_19966);
nor UO_678 (O_678,N_19993,N_19806);
nand UO_679 (O_679,N_19670,N_19928);
xor UO_680 (O_680,N_19613,N_19746);
nor UO_681 (O_681,N_19638,N_19802);
nand UO_682 (O_682,N_19770,N_19643);
or UO_683 (O_683,N_19624,N_19910);
or UO_684 (O_684,N_19946,N_19715);
xor UO_685 (O_685,N_19684,N_19897);
nor UO_686 (O_686,N_19700,N_19858);
nand UO_687 (O_687,N_19747,N_19937);
and UO_688 (O_688,N_19929,N_19825);
xor UO_689 (O_689,N_19726,N_19656);
and UO_690 (O_690,N_19859,N_19927);
nand UO_691 (O_691,N_19976,N_19721);
nand UO_692 (O_692,N_19669,N_19933);
nor UO_693 (O_693,N_19955,N_19626);
xor UO_694 (O_694,N_19610,N_19768);
nand UO_695 (O_695,N_19666,N_19935);
and UO_696 (O_696,N_19810,N_19930);
xnor UO_697 (O_697,N_19795,N_19662);
and UO_698 (O_698,N_19688,N_19719);
xnor UO_699 (O_699,N_19742,N_19796);
and UO_700 (O_700,N_19851,N_19971);
xnor UO_701 (O_701,N_19741,N_19783);
and UO_702 (O_702,N_19664,N_19996);
and UO_703 (O_703,N_19822,N_19821);
and UO_704 (O_704,N_19948,N_19806);
nand UO_705 (O_705,N_19917,N_19671);
or UO_706 (O_706,N_19752,N_19943);
xor UO_707 (O_707,N_19652,N_19942);
xnor UO_708 (O_708,N_19614,N_19928);
xor UO_709 (O_709,N_19683,N_19919);
or UO_710 (O_710,N_19640,N_19744);
xor UO_711 (O_711,N_19690,N_19698);
nor UO_712 (O_712,N_19659,N_19816);
nand UO_713 (O_713,N_19682,N_19708);
nor UO_714 (O_714,N_19816,N_19662);
and UO_715 (O_715,N_19739,N_19794);
xor UO_716 (O_716,N_19635,N_19713);
or UO_717 (O_717,N_19944,N_19637);
nand UO_718 (O_718,N_19827,N_19938);
or UO_719 (O_719,N_19681,N_19772);
and UO_720 (O_720,N_19695,N_19963);
or UO_721 (O_721,N_19609,N_19689);
nand UO_722 (O_722,N_19997,N_19760);
and UO_723 (O_723,N_19601,N_19789);
nand UO_724 (O_724,N_19961,N_19943);
nand UO_725 (O_725,N_19828,N_19723);
nand UO_726 (O_726,N_19652,N_19713);
or UO_727 (O_727,N_19791,N_19917);
nor UO_728 (O_728,N_19727,N_19965);
xnor UO_729 (O_729,N_19653,N_19903);
nand UO_730 (O_730,N_19776,N_19720);
xnor UO_731 (O_731,N_19799,N_19795);
and UO_732 (O_732,N_19674,N_19850);
xnor UO_733 (O_733,N_19907,N_19698);
nand UO_734 (O_734,N_19853,N_19971);
and UO_735 (O_735,N_19798,N_19618);
xnor UO_736 (O_736,N_19805,N_19716);
nor UO_737 (O_737,N_19716,N_19980);
nor UO_738 (O_738,N_19701,N_19841);
xor UO_739 (O_739,N_19856,N_19727);
or UO_740 (O_740,N_19719,N_19820);
nor UO_741 (O_741,N_19608,N_19781);
and UO_742 (O_742,N_19706,N_19887);
nor UO_743 (O_743,N_19654,N_19786);
and UO_744 (O_744,N_19972,N_19748);
nand UO_745 (O_745,N_19980,N_19618);
nor UO_746 (O_746,N_19839,N_19852);
nor UO_747 (O_747,N_19764,N_19684);
nor UO_748 (O_748,N_19973,N_19845);
nor UO_749 (O_749,N_19920,N_19927);
and UO_750 (O_750,N_19854,N_19780);
or UO_751 (O_751,N_19663,N_19985);
nand UO_752 (O_752,N_19897,N_19677);
and UO_753 (O_753,N_19718,N_19723);
nor UO_754 (O_754,N_19784,N_19846);
and UO_755 (O_755,N_19786,N_19892);
or UO_756 (O_756,N_19753,N_19789);
xor UO_757 (O_757,N_19767,N_19794);
xor UO_758 (O_758,N_19871,N_19885);
nand UO_759 (O_759,N_19683,N_19705);
nor UO_760 (O_760,N_19742,N_19679);
nand UO_761 (O_761,N_19977,N_19843);
nor UO_762 (O_762,N_19820,N_19603);
nor UO_763 (O_763,N_19845,N_19800);
or UO_764 (O_764,N_19631,N_19699);
and UO_765 (O_765,N_19725,N_19927);
or UO_766 (O_766,N_19868,N_19886);
xnor UO_767 (O_767,N_19804,N_19675);
or UO_768 (O_768,N_19943,N_19761);
nand UO_769 (O_769,N_19720,N_19843);
nor UO_770 (O_770,N_19659,N_19656);
and UO_771 (O_771,N_19631,N_19895);
xnor UO_772 (O_772,N_19770,N_19953);
or UO_773 (O_773,N_19755,N_19956);
nor UO_774 (O_774,N_19967,N_19946);
nand UO_775 (O_775,N_19634,N_19970);
or UO_776 (O_776,N_19827,N_19825);
nor UO_777 (O_777,N_19983,N_19766);
xnor UO_778 (O_778,N_19921,N_19761);
xor UO_779 (O_779,N_19953,N_19661);
xor UO_780 (O_780,N_19785,N_19637);
nand UO_781 (O_781,N_19607,N_19651);
nor UO_782 (O_782,N_19937,N_19846);
nand UO_783 (O_783,N_19680,N_19730);
nor UO_784 (O_784,N_19774,N_19768);
and UO_785 (O_785,N_19728,N_19650);
nor UO_786 (O_786,N_19653,N_19915);
nand UO_787 (O_787,N_19805,N_19901);
nor UO_788 (O_788,N_19603,N_19678);
nor UO_789 (O_789,N_19999,N_19921);
or UO_790 (O_790,N_19622,N_19723);
or UO_791 (O_791,N_19908,N_19926);
and UO_792 (O_792,N_19989,N_19695);
or UO_793 (O_793,N_19920,N_19951);
nand UO_794 (O_794,N_19702,N_19766);
nor UO_795 (O_795,N_19688,N_19950);
nor UO_796 (O_796,N_19667,N_19944);
and UO_797 (O_797,N_19916,N_19681);
and UO_798 (O_798,N_19866,N_19647);
or UO_799 (O_799,N_19976,N_19902);
nor UO_800 (O_800,N_19696,N_19972);
or UO_801 (O_801,N_19711,N_19962);
xnor UO_802 (O_802,N_19643,N_19857);
and UO_803 (O_803,N_19946,N_19981);
xnor UO_804 (O_804,N_19921,N_19695);
nand UO_805 (O_805,N_19678,N_19781);
and UO_806 (O_806,N_19615,N_19947);
and UO_807 (O_807,N_19884,N_19949);
and UO_808 (O_808,N_19652,N_19833);
and UO_809 (O_809,N_19714,N_19844);
nand UO_810 (O_810,N_19811,N_19907);
and UO_811 (O_811,N_19939,N_19917);
nand UO_812 (O_812,N_19968,N_19655);
xnor UO_813 (O_813,N_19661,N_19770);
or UO_814 (O_814,N_19850,N_19612);
and UO_815 (O_815,N_19977,N_19996);
or UO_816 (O_816,N_19720,N_19626);
xnor UO_817 (O_817,N_19952,N_19937);
or UO_818 (O_818,N_19754,N_19619);
xnor UO_819 (O_819,N_19686,N_19834);
nor UO_820 (O_820,N_19673,N_19808);
or UO_821 (O_821,N_19917,N_19620);
nor UO_822 (O_822,N_19709,N_19724);
nor UO_823 (O_823,N_19671,N_19845);
nor UO_824 (O_824,N_19927,N_19751);
nor UO_825 (O_825,N_19716,N_19625);
xor UO_826 (O_826,N_19822,N_19974);
nand UO_827 (O_827,N_19811,N_19942);
nand UO_828 (O_828,N_19661,N_19602);
nor UO_829 (O_829,N_19694,N_19657);
nand UO_830 (O_830,N_19688,N_19944);
and UO_831 (O_831,N_19981,N_19732);
or UO_832 (O_832,N_19696,N_19893);
nand UO_833 (O_833,N_19658,N_19614);
nand UO_834 (O_834,N_19719,N_19787);
nand UO_835 (O_835,N_19747,N_19834);
xor UO_836 (O_836,N_19977,N_19776);
and UO_837 (O_837,N_19995,N_19857);
nor UO_838 (O_838,N_19837,N_19805);
and UO_839 (O_839,N_19928,N_19761);
nand UO_840 (O_840,N_19686,N_19800);
xor UO_841 (O_841,N_19890,N_19674);
or UO_842 (O_842,N_19899,N_19879);
or UO_843 (O_843,N_19953,N_19918);
or UO_844 (O_844,N_19812,N_19786);
nor UO_845 (O_845,N_19820,N_19944);
or UO_846 (O_846,N_19651,N_19922);
nor UO_847 (O_847,N_19854,N_19938);
nand UO_848 (O_848,N_19918,N_19626);
xor UO_849 (O_849,N_19772,N_19975);
and UO_850 (O_850,N_19792,N_19663);
nand UO_851 (O_851,N_19922,N_19954);
nand UO_852 (O_852,N_19990,N_19768);
and UO_853 (O_853,N_19729,N_19907);
xor UO_854 (O_854,N_19771,N_19619);
and UO_855 (O_855,N_19774,N_19682);
and UO_856 (O_856,N_19853,N_19667);
nor UO_857 (O_857,N_19801,N_19620);
or UO_858 (O_858,N_19876,N_19608);
xnor UO_859 (O_859,N_19846,N_19621);
nor UO_860 (O_860,N_19776,N_19785);
and UO_861 (O_861,N_19897,N_19908);
and UO_862 (O_862,N_19969,N_19699);
or UO_863 (O_863,N_19836,N_19858);
or UO_864 (O_864,N_19902,N_19800);
nand UO_865 (O_865,N_19778,N_19855);
or UO_866 (O_866,N_19869,N_19937);
nand UO_867 (O_867,N_19914,N_19836);
nand UO_868 (O_868,N_19600,N_19629);
xnor UO_869 (O_869,N_19682,N_19946);
nor UO_870 (O_870,N_19699,N_19961);
xnor UO_871 (O_871,N_19805,N_19951);
nor UO_872 (O_872,N_19975,N_19905);
nor UO_873 (O_873,N_19885,N_19666);
or UO_874 (O_874,N_19892,N_19778);
or UO_875 (O_875,N_19694,N_19849);
and UO_876 (O_876,N_19614,N_19924);
nor UO_877 (O_877,N_19787,N_19793);
and UO_878 (O_878,N_19867,N_19824);
nand UO_879 (O_879,N_19627,N_19951);
xor UO_880 (O_880,N_19971,N_19702);
or UO_881 (O_881,N_19911,N_19788);
xnor UO_882 (O_882,N_19789,N_19671);
nor UO_883 (O_883,N_19839,N_19735);
and UO_884 (O_884,N_19714,N_19848);
xor UO_885 (O_885,N_19792,N_19729);
xnor UO_886 (O_886,N_19665,N_19836);
nand UO_887 (O_887,N_19806,N_19645);
nand UO_888 (O_888,N_19852,N_19624);
xor UO_889 (O_889,N_19800,N_19974);
nand UO_890 (O_890,N_19810,N_19833);
and UO_891 (O_891,N_19835,N_19743);
nor UO_892 (O_892,N_19926,N_19910);
and UO_893 (O_893,N_19618,N_19784);
xor UO_894 (O_894,N_19735,N_19845);
or UO_895 (O_895,N_19988,N_19878);
or UO_896 (O_896,N_19659,N_19934);
xnor UO_897 (O_897,N_19705,N_19633);
or UO_898 (O_898,N_19896,N_19637);
xnor UO_899 (O_899,N_19753,N_19847);
xnor UO_900 (O_900,N_19745,N_19664);
and UO_901 (O_901,N_19673,N_19871);
or UO_902 (O_902,N_19695,N_19747);
nand UO_903 (O_903,N_19915,N_19868);
nand UO_904 (O_904,N_19761,N_19936);
or UO_905 (O_905,N_19780,N_19934);
xor UO_906 (O_906,N_19751,N_19628);
xor UO_907 (O_907,N_19601,N_19749);
nor UO_908 (O_908,N_19602,N_19653);
nand UO_909 (O_909,N_19863,N_19625);
nor UO_910 (O_910,N_19686,N_19670);
and UO_911 (O_911,N_19723,N_19838);
or UO_912 (O_912,N_19967,N_19776);
nor UO_913 (O_913,N_19743,N_19758);
nand UO_914 (O_914,N_19893,N_19954);
nand UO_915 (O_915,N_19883,N_19694);
nor UO_916 (O_916,N_19757,N_19752);
or UO_917 (O_917,N_19906,N_19899);
xnor UO_918 (O_918,N_19770,N_19880);
nand UO_919 (O_919,N_19608,N_19990);
xnor UO_920 (O_920,N_19642,N_19975);
nand UO_921 (O_921,N_19698,N_19692);
xnor UO_922 (O_922,N_19667,N_19636);
nand UO_923 (O_923,N_19739,N_19990);
nor UO_924 (O_924,N_19790,N_19762);
xnor UO_925 (O_925,N_19780,N_19603);
xnor UO_926 (O_926,N_19691,N_19656);
or UO_927 (O_927,N_19819,N_19733);
nand UO_928 (O_928,N_19942,N_19847);
and UO_929 (O_929,N_19815,N_19934);
nand UO_930 (O_930,N_19690,N_19948);
xnor UO_931 (O_931,N_19672,N_19988);
xor UO_932 (O_932,N_19803,N_19607);
xor UO_933 (O_933,N_19707,N_19851);
nand UO_934 (O_934,N_19632,N_19641);
or UO_935 (O_935,N_19760,N_19826);
nor UO_936 (O_936,N_19704,N_19938);
or UO_937 (O_937,N_19815,N_19615);
nor UO_938 (O_938,N_19901,N_19854);
or UO_939 (O_939,N_19742,N_19858);
and UO_940 (O_940,N_19739,N_19840);
nand UO_941 (O_941,N_19776,N_19829);
xor UO_942 (O_942,N_19668,N_19858);
nand UO_943 (O_943,N_19853,N_19997);
nand UO_944 (O_944,N_19839,N_19695);
nand UO_945 (O_945,N_19651,N_19876);
or UO_946 (O_946,N_19690,N_19893);
xor UO_947 (O_947,N_19783,N_19765);
and UO_948 (O_948,N_19656,N_19820);
and UO_949 (O_949,N_19739,N_19979);
or UO_950 (O_950,N_19875,N_19873);
or UO_951 (O_951,N_19938,N_19682);
xnor UO_952 (O_952,N_19618,N_19732);
nor UO_953 (O_953,N_19642,N_19879);
and UO_954 (O_954,N_19834,N_19890);
nand UO_955 (O_955,N_19902,N_19919);
or UO_956 (O_956,N_19654,N_19843);
or UO_957 (O_957,N_19907,N_19938);
nand UO_958 (O_958,N_19992,N_19804);
nand UO_959 (O_959,N_19671,N_19932);
xnor UO_960 (O_960,N_19900,N_19947);
nand UO_961 (O_961,N_19698,N_19854);
nor UO_962 (O_962,N_19791,N_19645);
nand UO_963 (O_963,N_19773,N_19908);
nand UO_964 (O_964,N_19619,N_19869);
nor UO_965 (O_965,N_19923,N_19788);
or UO_966 (O_966,N_19659,N_19694);
nor UO_967 (O_967,N_19658,N_19736);
xnor UO_968 (O_968,N_19869,N_19670);
or UO_969 (O_969,N_19870,N_19762);
xnor UO_970 (O_970,N_19638,N_19953);
and UO_971 (O_971,N_19737,N_19793);
and UO_972 (O_972,N_19925,N_19731);
nand UO_973 (O_973,N_19913,N_19664);
and UO_974 (O_974,N_19808,N_19867);
xnor UO_975 (O_975,N_19782,N_19718);
or UO_976 (O_976,N_19905,N_19908);
xnor UO_977 (O_977,N_19955,N_19629);
nand UO_978 (O_978,N_19751,N_19727);
and UO_979 (O_979,N_19868,N_19631);
nand UO_980 (O_980,N_19807,N_19858);
nor UO_981 (O_981,N_19778,N_19761);
nand UO_982 (O_982,N_19667,N_19624);
xor UO_983 (O_983,N_19727,N_19919);
nor UO_984 (O_984,N_19899,N_19635);
xnor UO_985 (O_985,N_19608,N_19782);
and UO_986 (O_986,N_19740,N_19996);
xnor UO_987 (O_987,N_19720,N_19947);
and UO_988 (O_988,N_19841,N_19894);
xnor UO_989 (O_989,N_19996,N_19864);
nand UO_990 (O_990,N_19654,N_19987);
and UO_991 (O_991,N_19601,N_19706);
or UO_992 (O_992,N_19828,N_19858);
nand UO_993 (O_993,N_19783,N_19971);
nand UO_994 (O_994,N_19730,N_19693);
nor UO_995 (O_995,N_19994,N_19765);
nand UO_996 (O_996,N_19607,N_19836);
nand UO_997 (O_997,N_19700,N_19831);
nor UO_998 (O_998,N_19923,N_19970);
or UO_999 (O_999,N_19813,N_19650);
and UO_1000 (O_1000,N_19801,N_19894);
nand UO_1001 (O_1001,N_19897,N_19689);
xnor UO_1002 (O_1002,N_19946,N_19634);
and UO_1003 (O_1003,N_19974,N_19868);
nand UO_1004 (O_1004,N_19790,N_19725);
nor UO_1005 (O_1005,N_19602,N_19829);
and UO_1006 (O_1006,N_19929,N_19666);
nand UO_1007 (O_1007,N_19700,N_19646);
and UO_1008 (O_1008,N_19994,N_19784);
xnor UO_1009 (O_1009,N_19692,N_19850);
and UO_1010 (O_1010,N_19724,N_19890);
nand UO_1011 (O_1011,N_19918,N_19656);
nand UO_1012 (O_1012,N_19891,N_19862);
and UO_1013 (O_1013,N_19605,N_19659);
nor UO_1014 (O_1014,N_19639,N_19723);
and UO_1015 (O_1015,N_19800,N_19759);
xnor UO_1016 (O_1016,N_19948,N_19869);
nor UO_1017 (O_1017,N_19612,N_19807);
xnor UO_1018 (O_1018,N_19770,N_19832);
nor UO_1019 (O_1019,N_19895,N_19725);
nand UO_1020 (O_1020,N_19720,N_19941);
and UO_1021 (O_1021,N_19687,N_19834);
and UO_1022 (O_1022,N_19918,N_19781);
nor UO_1023 (O_1023,N_19759,N_19676);
or UO_1024 (O_1024,N_19928,N_19813);
or UO_1025 (O_1025,N_19722,N_19854);
or UO_1026 (O_1026,N_19826,N_19885);
or UO_1027 (O_1027,N_19968,N_19741);
and UO_1028 (O_1028,N_19989,N_19683);
xor UO_1029 (O_1029,N_19847,N_19636);
nor UO_1030 (O_1030,N_19937,N_19630);
nor UO_1031 (O_1031,N_19971,N_19795);
or UO_1032 (O_1032,N_19837,N_19655);
xor UO_1033 (O_1033,N_19658,N_19957);
xnor UO_1034 (O_1034,N_19915,N_19883);
or UO_1035 (O_1035,N_19993,N_19799);
xor UO_1036 (O_1036,N_19883,N_19790);
nand UO_1037 (O_1037,N_19858,N_19884);
nor UO_1038 (O_1038,N_19616,N_19608);
nor UO_1039 (O_1039,N_19697,N_19779);
nand UO_1040 (O_1040,N_19872,N_19781);
nor UO_1041 (O_1041,N_19906,N_19704);
nor UO_1042 (O_1042,N_19984,N_19704);
or UO_1043 (O_1043,N_19888,N_19912);
nor UO_1044 (O_1044,N_19867,N_19619);
or UO_1045 (O_1045,N_19790,N_19673);
and UO_1046 (O_1046,N_19781,N_19859);
and UO_1047 (O_1047,N_19620,N_19722);
or UO_1048 (O_1048,N_19951,N_19863);
and UO_1049 (O_1049,N_19994,N_19940);
xor UO_1050 (O_1050,N_19873,N_19779);
xor UO_1051 (O_1051,N_19989,N_19783);
xor UO_1052 (O_1052,N_19982,N_19868);
and UO_1053 (O_1053,N_19911,N_19645);
nand UO_1054 (O_1054,N_19726,N_19762);
xor UO_1055 (O_1055,N_19964,N_19751);
or UO_1056 (O_1056,N_19928,N_19626);
nand UO_1057 (O_1057,N_19803,N_19616);
nand UO_1058 (O_1058,N_19701,N_19937);
and UO_1059 (O_1059,N_19748,N_19695);
and UO_1060 (O_1060,N_19980,N_19708);
xnor UO_1061 (O_1061,N_19902,N_19679);
xor UO_1062 (O_1062,N_19661,N_19998);
nor UO_1063 (O_1063,N_19696,N_19771);
nor UO_1064 (O_1064,N_19905,N_19866);
nor UO_1065 (O_1065,N_19634,N_19684);
or UO_1066 (O_1066,N_19726,N_19805);
or UO_1067 (O_1067,N_19953,N_19697);
nand UO_1068 (O_1068,N_19642,N_19724);
and UO_1069 (O_1069,N_19865,N_19726);
nor UO_1070 (O_1070,N_19920,N_19651);
or UO_1071 (O_1071,N_19801,N_19939);
nor UO_1072 (O_1072,N_19872,N_19971);
or UO_1073 (O_1073,N_19952,N_19887);
and UO_1074 (O_1074,N_19703,N_19956);
nor UO_1075 (O_1075,N_19861,N_19842);
or UO_1076 (O_1076,N_19986,N_19640);
or UO_1077 (O_1077,N_19763,N_19634);
nor UO_1078 (O_1078,N_19841,N_19653);
xnor UO_1079 (O_1079,N_19766,N_19948);
and UO_1080 (O_1080,N_19800,N_19822);
and UO_1081 (O_1081,N_19876,N_19657);
nand UO_1082 (O_1082,N_19885,N_19731);
or UO_1083 (O_1083,N_19661,N_19813);
nand UO_1084 (O_1084,N_19646,N_19849);
nor UO_1085 (O_1085,N_19842,N_19728);
nand UO_1086 (O_1086,N_19725,N_19655);
nor UO_1087 (O_1087,N_19935,N_19774);
nand UO_1088 (O_1088,N_19633,N_19928);
nor UO_1089 (O_1089,N_19819,N_19956);
and UO_1090 (O_1090,N_19664,N_19794);
xnor UO_1091 (O_1091,N_19891,N_19842);
nand UO_1092 (O_1092,N_19965,N_19608);
nand UO_1093 (O_1093,N_19670,N_19757);
xor UO_1094 (O_1094,N_19884,N_19642);
nand UO_1095 (O_1095,N_19892,N_19875);
nand UO_1096 (O_1096,N_19955,N_19920);
nor UO_1097 (O_1097,N_19997,N_19626);
nor UO_1098 (O_1098,N_19780,N_19869);
xnor UO_1099 (O_1099,N_19685,N_19972);
nand UO_1100 (O_1100,N_19817,N_19850);
nand UO_1101 (O_1101,N_19783,N_19748);
xnor UO_1102 (O_1102,N_19614,N_19998);
xnor UO_1103 (O_1103,N_19847,N_19836);
xor UO_1104 (O_1104,N_19882,N_19970);
or UO_1105 (O_1105,N_19647,N_19942);
nor UO_1106 (O_1106,N_19915,N_19958);
xnor UO_1107 (O_1107,N_19883,N_19627);
and UO_1108 (O_1108,N_19983,N_19653);
or UO_1109 (O_1109,N_19697,N_19784);
nor UO_1110 (O_1110,N_19929,N_19990);
nor UO_1111 (O_1111,N_19760,N_19612);
or UO_1112 (O_1112,N_19815,N_19869);
or UO_1113 (O_1113,N_19737,N_19963);
and UO_1114 (O_1114,N_19613,N_19876);
and UO_1115 (O_1115,N_19811,N_19859);
nor UO_1116 (O_1116,N_19869,N_19944);
xor UO_1117 (O_1117,N_19993,N_19808);
nand UO_1118 (O_1118,N_19858,N_19876);
nand UO_1119 (O_1119,N_19831,N_19952);
or UO_1120 (O_1120,N_19753,N_19948);
xnor UO_1121 (O_1121,N_19799,N_19921);
nand UO_1122 (O_1122,N_19846,N_19988);
nand UO_1123 (O_1123,N_19832,N_19820);
or UO_1124 (O_1124,N_19998,N_19662);
nand UO_1125 (O_1125,N_19779,N_19606);
or UO_1126 (O_1126,N_19756,N_19835);
nand UO_1127 (O_1127,N_19830,N_19623);
or UO_1128 (O_1128,N_19732,N_19615);
nor UO_1129 (O_1129,N_19981,N_19661);
xor UO_1130 (O_1130,N_19672,N_19667);
and UO_1131 (O_1131,N_19640,N_19639);
or UO_1132 (O_1132,N_19660,N_19651);
xor UO_1133 (O_1133,N_19783,N_19897);
nand UO_1134 (O_1134,N_19824,N_19683);
or UO_1135 (O_1135,N_19643,N_19690);
nand UO_1136 (O_1136,N_19865,N_19963);
xnor UO_1137 (O_1137,N_19954,N_19754);
and UO_1138 (O_1138,N_19689,N_19688);
or UO_1139 (O_1139,N_19908,N_19958);
xnor UO_1140 (O_1140,N_19954,N_19762);
and UO_1141 (O_1141,N_19814,N_19604);
nand UO_1142 (O_1142,N_19744,N_19740);
nand UO_1143 (O_1143,N_19623,N_19915);
nand UO_1144 (O_1144,N_19679,N_19925);
nor UO_1145 (O_1145,N_19730,N_19662);
nand UO_1146 (O_1146,N_19604,N_19956);
xor UO_1147 (O_1147,N_19602,N_19959);
or UO_1148 (O_1148,N_19784,N_19657);
or UO_1149 (O_1149,N_19802,N_19821);
nor UO_1150 (O_1150,N_19655,N_19668);
nand UO_1151 (O_1151,N_19895,N_19714);
nor UO_1152 (O_1152,N_19897,N_19768);
xnor UO_1153 (O_1153,N_19603,N_19846);
nor UO_1154 (O_1154,N_19630,N_19962);
nand UO_1155 (O_1155,N_19715,N_19602);
xnor UO_1156 (O_1156,N_19888,N_19995);
nor UO_1157 (O_1157,N_19655,N_19673);
xor UO_1158 (O_1158,N_19616,N_19909);
nand UO_1159 (O_1159,N_19710,N_19765);
nor UO_1160 (O_1160,N_19745,N_19844);
nor UO_1161 (O_1161,N_19821,N_19969);
or UO_1162 (O_1162,N_19630,N_19677);
nor UO_1163 (O_1163,N_19869,N_19966);
or UO_1164 (O_1164,N_19788,N_19719);
xnor UO_1165 (O_1165,N_19896,N_19648);
and UO_1166 (O_1166,N_19782,N_19821);
and UO_1167 (O_1167,N_19806,N_19924);
nand UO_1168 (O_1168,N_19698,N_19646);
and UO_1169 (O_1169,N_19965,N_19913);
nor UO_1170 (O_1170,N_19745,N_19833);
nand UO_1171 (O_1171,N_19765,N_19971);
nand UO_1172 (O_1172,N_19626,N_19897);
nand UO_1173 (O_1173,N_19656,N_19697);
nand UO_1174 (O_1174,N_19737,N_19935);
or UO_1175 (O_1175,N_19638,N_19698);
and UO_1176 (O_1176,N_19841,N_19737);
and UO_1177 (O_1177,N_19838,N_19624);
or UO_1178 (O_1178,N_19771,N_19889);
nand UO_1179 (O_1179,N_19973,N_19881);
and UO_1180 (O_1180,N_19874,N_19998);
nand UO_1181 (O_1181,N_19837,N_19735);
nand UO_1182 (O_1182,N_19907,N_19783);
nor UO_1183 (O_1183,N_19655,N_19715);
and UO_1184 (O_1184,N_19922,N_19837);
nor UO_1185 (O_1185,N_19755,N_19765);
and UO_1186 (O_1186,N_19846,N_19804);
nand UO_1187 (O_1187,N_19765,N_19995);
or UO_1188 (O_1188,N_19664,N_19644);
xnor UO_1189 (O_1189,N_19807,N_19958);
and UO_1190 (O_1190,N_19684,N_19781);
xor UO_1191 (O_1191,N_19785,N_19955);
or UO_1192 (O_1192,N_19728,N_19716);
or UO_1193 (O_1193,N_19644,N_19726);
nor UO_1194 (O_1194,N_19657,N_19847);
and UO_1195 (O_1195,N_19951,N_19922);
or UO_1196 (O_1196,N_19745,N_19605);
nand UO_1197 (O_1197,N_19658,N_19817);
or UO_1198 (O_1198,N_19853,N_19693);
or UO_1199 (O_1199,N_19752,N_19731);
nand UO_1200 (O_1200,N_19745,N_19754);
or UO_1201 (O_1201,N_19790,N_19826);
or UO_1202 (O_1202,N_19880,N_19762);
nor UO_1203 (O_1203,N_19779,N_19604);
nand UO_1204 (O_1204,N_19949,N_19778);
xnor UO_1205 (O_1205,N_19853,N_19819);
or UO_1206 (O_1206,N_19690,N_19655);
nor UO_1207 (O_1207,N_19865,N_19931);
or UO_1208 (O_1208,N_19923,N_19622);
nor UO_1209 (O_1209,N_19752,N_19605);
nor UO_1210 (O_1210,N_19892,N_19728);
and UO_1211 (O_1211,N_19657,N_19963);
xnor UO_1212 (O_1212,N_19773,N_19712);
or UO_1213 (O_1213,N_19730,N_19792);
nor UO_1214 (O_1214,N_19761,N_19852);
nand UO_1215 (O_1215,N_19672,N_19974);
nand UO_1216 (O_1216,N_19925,N_19885);
nand UO_1217 (O_1217,N_19700,N_19770);
or UO_1218 (O_1218,N_19799,N_19867);
nor UO_1219 (O_1219,N_19680,N_19702);
and UO_1220 (O_1220,N_19739,N_19803);
or UO_1221 (O_1221,N_19940,N_19616);
xor UO_1222 (O_1222,N_19751,N_19712);
nor UO_1223 (O_1223,N_19601,N_19855);
xnor UO_1224 (O_1224,N_19980,N_19706);
nand UO_1225 (O_1225,N_19915,N_19992);
or UO_1226 (O_1226,N_19724,N_19911);
and UO_1227 (O_1227,N_19744,N_19629);
or UO_1228 (O_1228,N_19938,N_19803);
and UO_1229 (O_1229,N_19770,N_19788);
xor UO_1230 (O_1230,N_19668,N_19663);
and UO_1231 (O_1231,N_19991,N_19871);
xnor UO_1232 (O_1232,N_19879,N_19602);
xor UO_1233 (O_1233,N_19927,N_19866);
and UO_1234 (O_1234,N_19701,N_19816);
nor UO_1235 (O_1235,N_19706,N_19996);
or UO_1236 (O_1236,N_19672,N_19718);
xor UO_1237 (O_1237,N_19776,N_19687);
xnor UO_1238 (O_1238,N_19989,N_19996);
nand UO_1239 (O_1239,N_19649,N_19833);
or UO_1240 (O_1240,N_19633,N_19803);
or UO_1241 (O_1241,N_19924,N_19670);
or UO_1242 (O_1242,N_19655,N_19884);
or UO_1243 (O_1243,N_19891,N_19985);
and UO_1244 (O_1244,N_19874,N_19675);
and UO_1245 (O_1245,N_19868,N_19739);
and UO_1246 (O_1246,N_19796,N_19618);
nand UO_1247 (O_1247,N_19899,N_19709);
nor UO_1248 (O_1248,N_19788,N_19811);
nand UO_1249 (O_1249,N_19946,N_19887);
nand UO_1250 (O_1250,N_19682,N_19918);
and UO_1251 (O_1251,N_19612,N_19835);
xor UO_1252 (O_1252,N_19635,N_19781);
xnor UO_1253 (O_1253,N_19644,N_19830);
xor UO_1254 (O_1254,N_19725,N_19628);
nor UO_1255 (O_1255,N_19844,N_19783);
nor UO_1256 (O_1256,N_19804,N_19745);
nand UO_1257 (O_1257,N_19857,N_19605);
nor UO_1258 (O_1258,N_19802,N_19745);
or UO_1259 (O_1259,N_19975,N_19765);
nor UO_1260 (O_1260,N_19771,N_19870);
and UO_1261 (O_1261,N_19758,N_19825);
nor UO_1262 (O_1262,N_19967,N_19684);
nand UO_1263 (O_1263,N_19757,N_19867);
nor UO_1264 (O_1264,N_19633,N_19670);
xnor UO_1265 (O_1265,N_19853,N_19957);
nor UO_1266 (O_1266,N_19701,N_19821);
and UO_1267 (O_1267,N_19849,N_19850);
or UO_1268 (O_1268,N_19732,N_19946);
or UO_1269 (O_1269,N_19746,N_19863);
and UO_1270 (O_1270,N_19718,N_19964);
xnor UO_1271 (O_1271,N_19815,N_19814);
nor UO_1272 (O_1272,N_19631,N_19831);
xor UO_1273 (O_1273,N_19639,N_19662);
and UO_1274 (O_1274,N_19736,N_19669);
or UO_1275 (O_1275,N_19837,N_19702);
or UO_1276 (O_1276,N_19939,N_19863);
or UO_1277 (O_1277,N_19943,N_19676);
and UO_1278 (O_1278,N_19837,N_19900);
and UO_1279 (O_1279,N_19867,N_19775);
xor UO_1280 (O_1280,N_19728,N_19813);
nand UO_1281 (O_1281,N_19661,N_19686);
or UO_1282 (O_1282,N_19928,N_19784);
nand UO_1283 (O_1283,N_19896,N_19829);
xnor UO_1284 (O_1284,N_19763,N_19764);
nand UO_1285 (O_1285,N_19750,N_19614);
nor UO_1286 (O_1286,N_19788,N_19715);
nor UO_1287 (O_1287,N_19898,N_19665);
nor UO_1288 (O_1288,N_19809,N_19955);
or UO_1289 (O_1289,N_19676,N_19840);
nor UO_1290 (O_1290,N_19657,N_19660);
or UO_1291 (O_1291,N_19749,N_19628);
nor UO_1292 (O_1292,N_19719,N_19798);
nand UO_1293 (O_1293,N_19837,N_19842);
nor UO_1294 (O_1294,N_19659,N_19849);
or UO_1295 (O_1295,N_19664,N_19981);
nor UO_1296 (O_1296,N_19910,N_19770);
nor UO_1297 (O_1297,N_19968,N_19782);
nor UO_1298 (O_1298,N_19932,N_19662);
xnor UO_1299 (O_1299,N_19884,N_19611);
and UO_1300 (O_1300,N_19845,N_19981);
nor UO_1301 (O_1301,N_19859,N_19753);
xnor UO_1302 (O_1302,N_19769,N_19725);
and UO_1303 (O_1303,N_19629,N_19944);
nor UO_1304 (O_1304,N_19612,N_19752);
or UO_1305 (O_1305,N_19624,N_19847);
xnor UO_1306 (O_1306,N_19946,N_19997);
xor UO_1307 (O_1307,N_19938,N_19708);
nand UO_1308 (O_1308,N_19766,N_19659);
nand UO_1309 (O_1309,N_19624,N_19698);
nand UO_1310 (O_1310,N_19855,N_19816);
xor UO_1311 (O_1311,N_19972,N_19882);
and UO_1312 (O_1312,N_19881,N_19848);
nand UO_1313 (O_1313,N_19834,N_19695);
and UO_1314 (O_1314,N_19651,N_19937);
nor UO_1315 (O_1315,N_19973,N_19868);
nand UO_1316 (O_1316,N_19661,N_19869);
or UO_1317 (O_1317,N_19740,N_19855);
xnor UO_1318 (O_1318,N_19869,N_19651);
xnor UO_1319 (O_1319,N_19985,N_19620);
xor UO_1320 (O_1320,N_19732,N_19704);
nor UO_1321 (O_1321,N_19643,N_19985);
xor UO_1322 (O_1322,N_19798,N_19859);
nand UO_1323 (O_1323,N_19851,N_19688);
nand UO_1324 (O_1324,N_19603,N_19639);
or UO_1325 (O_1325,N_19782,N_19774);
nand UO_1326 (O_1326,N_19914,N_19786);
nand UO_1327 (O_1327,N_19640,N_19784);
and UO_1328 (O_1328,N_19643,N_19738);
nor UO_1329 (O_1329,N_19801,N_19642);
or UO_1330 (O_1330,N_19903,N_19741);
xnor UO_1331 (O_1331,N_19699,N_19609);
or UO_1332 (O_1332,N_19619,N_19904);
nor UO_1333 (O_1333,N_19649,N_19677);
and UO_1334 (O_1334,N_19800,N_19798);
nor UO_1335 (O_1335,N_19992,N_19965);
and UO_1336 (O_1336,N_19759,N_19861);
nand UO_1337 (O_1337,N_19673,N_19647);
nor UO_1338 (O_1338,N_19668,N_19841);
xnor UO_1339 (O_1339,N_19898,N_19760);
or UO_1340 (O_1340,N_19908,N_19970);
or UO_1341 (O_1341,N_19753,N_19959);
nand UO_1342 (O_1342,N_19733,N_19670);
nand UO_1343 (O_1343,N_19911,N_19776);
nand UO_1344 (O_1344,N_19672,N_19923);
and UO_1345 (O_1345,N_19643,N_19822);
nor UO_1346 (O_1346,N_19976,N_19792);
and UO_1347 (O_1347,N_19766,N_19886);
nor UO_1348 (O_1348,N_19947,N_19878);
xor UO_1349 (O_1349,N_19752,N_19667);
nand UO_1350 (O_1350,N_19784,N_19868);
xnor UO_1351 (O_1351,N_19817,N_19840);
and UO_1352 (O_1352,N_19616,N_19821);
nand UO_1353 (O_1353,N_19736,N_19828);
nand UO_1354 (O_1354,N_19847,N_19826);
nand UO_1355 (O_1355,N_19988,N_19777);
and UO_1356 (O_1356,N_19654,N_19912);
xor UO_1357 (O_1357,N_19678,N_19676);
xor UO_1358 (O_1358,N_19880,N_19833);
and UO_1359 (O_1359,N_19718,N_19948);
and UO_1360 (O_1360,N_19806,N_19640);
nor UO_1361 (O_1361,N_19779,N_19857);
and UO_1362 (O_1362,N_19755,N_19930);
and UO_1363 (O_1363,N_19658,N_19907);
and UO_1364 (O_1364,N_19956,N_19905);
or UO_1365 (O_1365,N_19870,N_19786);
or UO_1366 (O_1366,N_19915,N_19816);
or UO_1367 (O_1367,N_19883,N_19874);
or UO_1368 (O_1368,N_19922,N_19748);
nor UO_1369 (O_1369,N_19822,N_19889);
or UO_1370 (O_1370,N_19936,N_19625);
xor UO_1371 (O_1371,N_19902,N_19666);
and UO_1372 (O_1372,N_19620,N_19705);
or UO_1373 (O_1373,N_19860,N_19891);
nand UO_1374 (O_1374,N_19771,N_19615);
and UO_1375 (O_1375,N_19876,N_19778);
or UO_1376 (O_1376,N_19933,N_19888);
nor UO_1377 (O_1377,N_19705,N_19892);
nor UO_1378 (O_1378,N_19623,N_19859);
nor UO_1379 (O_1379,N_19881,N_19846);
or UO_1380 (O_1380,N_19967,N_19674);
and UO_1381 (O_1381,N_19869,N_19779);
or UO_1382 (O_1382,N_19977,N_19851);
nor UO_1383 (O_1383,N_19667,N_19613);
or UO_1384 (O_1384,N_19868,N_19857);
xor UO_1385 (O_1385,N_19910,N_19701);
xnor UO_1386 (O_1386,N_19670,N_19850);
and UO_1387 (O_1387,N_19811,N_19762);
and UO_1388 (O_1388,N_19686,N_19789);
and UO_1389 (O_1389,N_19630,N_19886);
nor UO_1390 (O_1390,N_19975,N_19977);
nor UO_1391 (O_1391,N_19771,N_19610);
xnor UO_1392 (O_1392,N_19814,N_19621);
or UO_1393 (O_1393,N_19763,N_19814);
nor UO_1394 (O_1394,N_19748,N_19909);
xor UO_1395 (O_1395,N_19601,N_19969);
nor UO_1396 (O_1396,N_19829,N_19714);
or UO_1397 (O_1397,N_19680,N_19954);
nand UO_1398 (O_1398,N_19781,N_19905);
nor UO_1399 (O_1399,N_19668,N_19988);
xnor UO_1400 (O_1400,N_19905,N_19639);
nand UO_1401 (O_1401,N_19718,N_19800);
nand UO_1402 (O_1402,N_19996,N_19738);
nand UO_1403 (O_1403,N_19635,N_19797);
or UO_1404 (O_1404,N_19842,N_19973);
nand UO_1405 (O_1405,N_19802,N_19699);
nor UO_1406 (O_1406,N_19604,N_19615);
and UO_1407 (O_1407,N_19664,N_19755);
and UO_1408 (O_1408,N_19820,N_19679);
xor UO_1409 (O_1409,N_19848,N_19678);
and UO_1410 (O_1410,N_19737,N_19826);
and UO_1411 (O_1411,N_19914,N_19630);
xor UO_1412 (O_1412,N_19958,N_19600);
nor UO_1413 (O_1413,N_19681,N_19799);
nor UO_1414 (O_1414,N_19765,N_19651);
xor UO_1415 (O_1415,N_19606,N_19967);
nand UO_1416 (O_1416,N_19823,N_19874);
or UO_1417 (O_1417,N_19618,N_19822);
or UO_1418 (O_1418,N_19930,N_19788);
or UO_1419 (O_1419,N_19949,N_19612);
or UO_1420 (O_1420,N_19876,N_19768);
and UO_1421 (O_1421,N_19789,N_19933);
and UO_1422 (O_1422,N_19820,N_19633);
or UO_1423 (O_1423,N_19773,N_19621);
nand UO_1424 (O_1424,N_19960,N_19614);
xor UO_1425 (O_1425,N_19818,N_19741);
or UO_1426 (O_1426,N_19640,N_19613);
or UO_1427 (O_1427,N_19653,N_19631);
and UO_1428 (O_1428,N_19662,N_19894);
xor UO_1429 (O_1429,N_19916,N_19975);
nand UO_1430 (O_1430,N_19721,N_19818);
nor UO_1431 (O_1431,N_19710,N_19631);
or UO_1432 (O_1432,N_19942,N_19628);
xor UO_1433 (O_1433,N_19928,N_19659);
or UO_1434 (O_1434,N_19950,N_19643);
nand UO_1435 (O_1435,N_19954,N_19848);
or UO_1436 (O_1436,N_19815,N_19708);
or UO_1437 (O_1437,N_19831,N_19626);
xnor UO_1438 (O_1438,N_19952,N_19716);
nor UO_1439 (O_1439,N_19801,N_19717);
nand UO_1440 (O_1440,N_19718,N_19797);
xnor UO_1441 (O_1441,N_19938,N_19884);
nor UO_1442 (O_1442,N_19719,N_19956);
or UO_1443 (O_1443,N_19922,N_19771);
xnor UO_1444 (O_1444,N_19970,N_19998);
nand UO_1445 (O_1445,N_19741,N_19891);
nand UO_1446 (O_1446,N_19857,N_19908);
nor UO_1447 (O_1447,N_19942,N_19613);
nor UO_1448 (O_1448,N_19719,N_19712);
nor UO_1449 (O_1449,N_19846,N_19658);
and UO_1450 (O_1450,N_19974,N_19854);
or UO_1451 (O_1451,N_19626,N_19746);
or UO_1452 (O_1452,N_19769,N_19904);
nor UO_1453 (O_1453,N_19711,N_19783);
and UO_1454 (O_1454,N_19924,N_19779);
nand UO_1455 (O_1455,N_19714,N_19737);
xor UO_1456 (O_1456,N_19608,N_19871);
nand UO_1457 (O_1457,N_19771,N_19670);
nor UO_1458 (O_1458,N_19987,N_19692);
and UO_1459 (O_1459,N_19828,N_19721);
xor UO_1460 (O_1460,N_19779,N_19992);
nor UO_1461 (O_1461,N_19666,N_19681);
nor UO_1462 (O_1462,N_19861,N_19876);
nor UO_1463 (O_1463,N_19770,N_19652);
nand UO_1464 (O_1464,N_19894,N_19869);
nor UO_1465 (O_1465,N_19968,N_19947);
nor UO_1466 (O_1466,N_19915,N_19865);
nor UO_1467 (O_1467,N_19671,N_19799);
or UO_1468 (O_1468,N_19825,N_19795);
nor UO_1469 (O_1469,N_19651,N_19983);
and UO_1470 (O_1470,N_19842,N_19945);
nand UO_1471 (O_1471,N_19857,N_19925);
and UO_1472 (O_1472,N_19782,N_19984);
or UO_1473 (O_1473,N_19658,N_19986);
nand UO_1474 (O_1474,N_19731,N_19649);
or UO_1475 (O_1475,N_19921,N_19830);
nand UO_1476 (O_1476,N_19952,N_19917);
nor UO_1477 (O_1477,N_19811,N_19886);
and UO_1478 (O_1478,N_19636,N_19941);
xnor UO_1479 (O_1479,N_19956,N_19976);
nand UO_1480 (O_1480,N_19718,N_19973);
nand UO_1481 (O_1481,N_19717,N_19803);
nor UO_1482 (O_1482,N_19780,N_19651);
and UO_1483 (O_1483,N_19852,N_19642);
and UO_1484 (O_1484,N_19711,N_19734);
and UO_1485 (O_1485,N_19899,N_19896);
xnor UO_1486 (O_1486,N_19965,N_19787);
nand UO_1487 (O_1487,N_19711,N_19947);
xor UO_1488 (O_1488,N_19787,N_19875);
xnor UO_1489 (O_1489,N_19768,N_19879);
nor UO_1490 (O_1490,N_19814,N_19656);
or UO_1491 (O_1491,N_19754,N_19850);
or UO_1492 (O_1492,N_19954,N_19979);
nor UO_1493 (O_1493,N_19718,N_19708);
nor UO_1494 (O_1494,N_19783,N_19637);
nor UO_1495 (O_1495,N_19680,N_19970);
nor UO_1496 (O_1496,N_19992,N_19929);
nor UO_1497 (O_1497,N_19798,N_19860);
and UO_1498 (O_1498,N_19811,N_19783);
nor UO_1499 (O_1499,N_19951,N_19810);
xor UO_1500 (O_1500,N_19897,N_19928);
nor UO_1501 (O_1501,N_19816,N_19787);
and UO_1502 (O_1502,N_19693,N_19869);
xor UO_1503 (O_1503,N_19774,N_19800);
nand UO_1504 (O_1504,N_19788,N_19795);
and UO_1505 (O_1505,N_19986,N_19875);
nor UO_1506 (O_1506,N_19955,N_19952);
and UO_1507 (O_1507,N_19606,N_19900);
nor UO_1508 (O_1508,N_19871,N_19955);
xor UO_1509 (O_1509,N_19711,N_19718);
and UO_1510 (O_1510,N_19825,N_19791);
and UO_1511 (O_1511,N_19653,N_19771);
nor UO_1512 (O_1512,N_19825,N_19761);
nand UO_1513 (O_1513,N_19721,N_19636);
or UO_1514 (O_1514,N_19904,N_19633);
nor UO_1515 (O_1515,N_19611,N_19885);
nor UO_1516 (O_1516,N_19860,N_19855);
nor UO_1517 (O_1517,N_19868,N_19883);
nor UO_1518 (O_1518,N_19888,N_19991);
xor UO_1519 (O_1519,N_19918,N_19934);
xor UO_1520 (O_1520,N_19732,N_19805);
nor UO_1521 (O_1521,N_19703,N_19733);
and UO_1522 (O_1522,N_19687,N_19702);
nor UO_1523 (O_1523,N_19600,N_19832);
xor UO_1524 (O_1524,N_19847,N_19893);
and UO_1525 (O_1525,N_19866,N_19738);
nor UO_1526 (O_1526,N_19664,N_19774);
and UO_1527 (O_1527,N_19719,N_19630);
or UO_1528 (O_1528,N_19787,N_19666);
and UO_1529 (O_1529,N_19612,N_19991);
and UO_1530 (O_1530,N_19630,N_19798);
nand UO_1531 (O_1531,N_19707,N_19722);
xnor UO_1532 (O_1532,N_19759,N_19628);
nand UO_1533 (O_1533,N_19659,N_19875);
xor UO_1534 (O_1534,N_19770,N_19747);
nor UO_1535 (O_1535,N_19664,N_19935);
xnor UO_1536 (O_1536,N_19720,N_19739);
nor UO_1537 (O_1537,N_19800,N_19835);
nor UO_1538 (O_1538,N_19624,N_19883);
nand UO_1539 (O_1539,N_19887,N_19747);
or UO_1540 (O_1540,N_19661,N_19916);
or UO_1541 (O_1541,N_19656,N_19891);
xor UO_1542 (O_1542,N_19835,N_19975);
xor UO_1543 (O_1543,N_19779,N_19968);
nand UO_1544 (O_1544,N_19742,N_19790);
or UO_1545 (O_1545,N_19880,N_19970);
xor UO_1546 (O_1546,N_19701,N_19674);
nor UO_1547 (O_1547,N_19755,N_19767);
or UO_1548 (O_1548,N_19967,N_19770);
xor UO_1549 (O_1549,N_19867,N_19657);
and UO_1550 (O_1550,N_19610,N_19649);
or UO_1551 (O_1551,N_19915,N_19646);
nand UO_1552 (O_1552,N_19812,N_19982);
xnor UO_1553 (O_1553,N_19924,N_19755);
nand UO_1554 (O_1554,N_19600,N_19829);
or UO_1555 (O_1555,N_19664,N_19830);
nand UO_1556 (O_1556,N_19828,N_19777);
or UO_1557 (O_1557,N_19875,N_19632);
xnor UO_1558 (O_1558,N_19940,N_19729);
nor UO_1559 (O_1559,N_19647,N_19820);
nand UO_1560 (O_1560,N_19934,N_19993);
xnor UO_1561 (O_1561,N_19689,N_19717);
xnor UO_1562 (O_1562,N_19975,N_19717);
xnor UO_1563 (O_1563,N_19729,N_19843);
nor UO_1564 (O_1564,N_19955,N_19861);
xor UO_1565 (O_1565,N_19858,N_19967);
and UO_1566 (O_1566,N_19933,N_19630);
xnor UO_1567 (O_1567,N_19913,N_19703);
nand UO_1568 (O_1568,N_19801,N_19880);
and UO_1569 (O_1569,N_19778,N_19981);
nor UO_1570 (O_1570,N_19817,N_19686);
nand UO_1571 (O_1571,N_19923,N_19663);
xnor UO_1572 (O_1572,N_19939,N_19988);
xnor UO_1573 (O_1573,N_19967,N_19773);
nand UO_1574 (O_1574,N_19974,N_19864);
nor UO_1575 (O_1575,N_19786,N_19719);
nand UO_1576 (O_1576,N_19860,N_19871);
nand UO_1577 (O_1577,N_19899,N_19807);
nor UO_1578 (O_1578,N_19849,N_19600);
xor UO_1579 (O_1579,N_19912,N_19929);
nor UO_1580 (O_1580,N_19825,N_19691);
nor UO_1581 (O_1581,N_19966,N_19935);
nand UO_1582 (O_1582,N_19771,N_19760);
xor UO_1583 (O_1583,N_19998,N_19864);
nor UO_1584 (O_1584,N_19882,N_19736);
nand UO_1585 (O_1585,N_19904,N_19713);
nand UO_1586 (O_1586,N_19631,N_19927);
nand UO_1587 (O_1587,N_19830,N_19680);
xor UO_1588 (O_1588,N_19793,N_19715);
nand UO_1589 (O_1589,N_19951,N_19924);
and UO_1590 (O_1590,N_19953,N_19758);
xnor UO_1591 (O_1591,N_19688,N_19645);
and UO_1592 (O_1592,N_19673,N_19661);
nand UO_1593 (O_1593,N_19934,N_19859);
nand UO_1594 (O_1594,N_19954,N_19952);
nand UO_1595 (O_1595,N_19856,N_19726);
or UO_1596 (O_1596,N_19749,N_19755);
or UO_1597 (O_1597,N_19725,N_19767);
or UO_1598 (O_1598,N_19953,N_19858);
nand UO_1599 (O_1599,N_19857,N_19998);
or UO_1600 (O_1600,N_19752,N_19727);
xnor UO_1601 (O_1601,N_19869,N_19650);
or UO_1602 (O_1602,N_19866,N_19771);
nand UO_1603 (O_1603,N_19776,N_19624);
or UO_1604 (O_1604,N_19633,N_19618);
xnor UO_1605 (O_1605,N_19830,N_19790);
nand UO_1606 (O_1606,N_19667,N_19621);
nand UO_1607 (O_1607,N_19807,N_19914);
and UO_1608 (O_1608,N_19899,N_19620);
nor UO_1609 (O_1609,N_19994,N_19806);
xor UO_1610 (O_1610,N_19648,N_19977);
or UO_1611 (O_1611,N_19610,N_19965);
nor UO_1612 (O_1612,N_19703,N_19741);
nor UO_1613 (O_1613,N_19981,N_19738);
xnor UO_1614 (O_1614,N_19613,N_19826);
nor UO_1615 (O_1615,N_19852,N_19879);
nor UO_1616 (O_1616,N_19871,N_19798);
nand UO_1617 (O_1617,N_19604,N_19902);
or UO_1618 (O_1618,N_19846,N_19925);
nand UO_1619 (O_1619,N_19780,N_19997);
nand UO_1620 (O_1620,N_19993,N_19687);
xnor UO_1621 (O_1621,N_19834,N_19831);
xor UO_1622 (O_1622,N_19672,N_19663);
xnor UO_1623 (O_1623,N_19798,N_19975);
nor UO_1624 (O_1624,N_19937,N_19954);
xnor UO_1625 (O_1625,N_19652,N_19926);
xor UO_1626 (O_1626,N_19831,N_19974);
xnor UO_1627 (O_1627,N_19781,N_19651);
nor UO_1628 (O_1628,N_19729,N_19734);
and UO_1629 (O_1629,N_19715,N_19902);
and UO_1630 (O_1630,N_19815,N_19759);
or UO_1631 (O_1631,N_19928,N_19719);
nor UO_1632 (O_1632,N_19934,N_19945);
nor UO_1633 (O_1633,N_19645,N_19845);
nand UO_1634 (O_1634,N_19813,N_19617);
nand UO_1635 (O_1635,N_19873,N_19847);
nand UO_1636 (O_1636,N_19855,N_19615);
nand UO_1637 (O_1637,N_19712,N_19977);
xnor UO_1638 (O_1638,N_19922,N_19888);
xnor UO_1639 (O_1639,N_19748,N_19699);
or UO_1640 (O_1640,N_19997,N_19963);
xor UO_1641 (O_1641,N_19740,N_19977);
nand UO_1642 (O_1642,N_19979,N_19764);
or UO_1643 (O_1643,N_19989,N_19701);
or UO_1644 (O_1644,N_19616,N_19848);
nor UO_1645 (O_1645,N_19727,N_19665);
or UO_1646 (O_1646,N_19944,N_19646);
and UO_1647 (O_1647,N_19685,N_19891);
xor UO_1648 (O_1648,N_19635,N_19848);
and UO_1649 (O_1649,N_19996,N_19771);
and UO_1650 (O_1650,N_19620,N_19878);
and UO_1651 (O_1651,N_19637,N_19826);
or UO_1652 (O_1652,N_19666,N_19898);
xnor UO_1653 (O_1653,N_19627,N_19740);
or UO_1654 (O_1654,N_19624,N_19810);
nor UO_1655 (O_1655,N_19662,N_19764);
xnor UO_1656 (O_1656,N_19629,N_19933);
nor UO_1657 (O_1657,N_19693,N_19976);
nor UO_1658 (O_1658,N_19987,N_19630);
or UO_1659 (O_1659,N_19921,N_19822);
and UO_1660 (O_1660,N_19675,N_19765);
and UO_1661 (O_1661,N_19752,N_19788);
nand UO_1662 (O_1662,N_19664,N_19920);
xnor UO_1663 (O_1663,N_19889,N_19950);
nand UO_1664 (O_1664,N_19839,N_19877);
or UO_1665 (O_1665,N_19630,N_19658);
nand UO_1666 (O_1666,N_19899,N_19851);
nor UO_1667 (O_1667,N_19718,N_19924);
nand UO_1668 (O_1668,N_19866,N_19706);
or UO_1669 (O_1669,N_19908,N_19916);
and UO_1670 (O_1670,N_19651,N_19662);
or UO_1671 (O_1671,N_19898,N_19621);
or UO_1672 (O_1672,N_19939,N_19758);
nor UO_1673 (O_1673,N_19650,N_19607);
or UO_1674 (O_1674,N_19882,N_19674);
and UO_1675 (O_1675,N_19686,N_19930);
nand UO_1676 (O_1676,N_19762,N_19791);
or UO_1677 (O_1677,N_19814,N_19965);
or UO_1678 (O_1678,N_19686,N_19843);
or UO_1679 (O_1679,N_19794,N_19854);
xor UO_1680 (O_1680,N_19662,N_19957);
and UO_1681 (O_1681,N_19893,N_19850);
nand UO_1682 (O_1682,N_19896,N_19663);
nand UO_1683 (O_1683,N_19995,N_19800);
xor UO_1684 (O_1684,N_19981,N_19813);
nand UO_1685 (O_1685,N_19972,N_19663);
or UO_1686 (O_1686,N_19741,N_19853);
or UO_1687 (O_1687,N_19917,N_19886);
or UO_1688 (O_1688,N_19672,N_19699);
xor UO_1689 (O_1689,N_19653,N_19615);
or UO_1690 (O_1690,N_19682,N_19984);
and UO_1691 (O_1691,N_19708,N_19628);
nand UO_1692 (O_1692,N_19770,N_19940);
and UO_1693 (O_1693,N_19724,N_19974);
nor UO_1694 (O_1694,N_19820,N_19824);
or UO_1695 (O_1695,N_19890,N_19663);
nor UO_1696 (O_1696,N_19614,N_19823);
xnor UO_1697 (O_1697,N_19890,N_19764);
or UO_1698 (O_1698,N_19660,N_19974);
nor UO_1699 (O_1699,N_19973,N_19694);
nor UO_1700 (O_1700,N_19660,N_19871);
nor UO_1701 (O_1701,N_19746,N_19745);
and UO_1702 (O_1702,N_19973,N_19628);
and UO_1703 (O_1703,N_19600,N_19631);
nand UO_1704 (O_1704,N_19743,N_19801);
and UO_1705 (O_1705,N_19672,N_19627);
and UO_1706 (O_1706,N_19977,N_19938);
and UO_1707 (O_1707,N_19686,N_19765);
and UO_1708 (O_1708,N_19789,N_19892);
or UO_1709 (O_1709,N_19941,N_19907);
nand UO_1710 (O_1710,N_19686,N_19757);
and UO_1711 (O_1711,N_19677,N_19803);
nor UO_1712 (O_1712,N_19820,N_19995);
nand UO_1713 (O_1713,N_19736,N_19843);
nand UO_1714 (O_1714,N_19835,N_19784);
nor UO_1715 (O_1715,N_19997,N_19884);
and UO_1716 (O_1716,N_19978,N_19876);
xor UO_1717 (O_1717,N_19955,N_19753);
nand UO_1718 (O_1718,N_19914,N_19779);
and UO_1719 (O_1719,N_19668,N_19875);
nor UO_1720 (O_1720,N_19697,N_19893);
or UO_1721 (O_1721,N_19853,N_19691);
xor UO_1722 (O_1722,N_19721,N_19772);
and UO_1723 (O_1723,N_19982,N_19727);
nand UO_1724 (O_1724,N_19811,N_19922);
or UO_1725 (O_1725,N_19670,N_19856);
nor UO_1726 (O_1726,N_19924,N_19774);
nand UO_1727 (O_1727,N_19992,N_19731);
nand UO_1728 (O_1728,N_19917,N_19677);
nand UO_1729 (O_1729,N_19987,N_19603);
or UO_1730 (O_1730,N_19871,N_19970);
nor UO_1731 (O_1731,N_19726,N_19699);
and UO_1732 (O_1732,N_19800,N_19659);
and UO_1733 (O_1733,N_19987,N_19993);
nand UO_1734 (O_1734,N_19932,N_19909);
or UO_1735 (O_1735,N_19626,N_19810);
nor UO_1736 (O_1736,N_19844,N_19979);
xnor UO_1737 (O_1737,N_19879,N_19862);
nor UO_1738 (O_1738,N_19654,N_19937);
and UO_1739 (O_1739,N_19872,N_19780);
nand UO_1740 (O_1740,N_19772,N_19844);
xor UO_1741 (O_1741,N_19821,N_19991);
or UO_1742 (O_1742,N_19872,N_19626);
nor UO_1743 (O_1743,N_19630,N_19988);
nand UO_1744 (O_1744,N_19855,N_19910);
xor UO_1745 (O_1745,N_19917,N_19975);
or UO_1746 (O_1746,N_19826,N_19652);
xor UO_1747 (O_1747,N_19753,N_19757);
and UO_1748 (O_1748,N_19692,N_19619);
nor UO_1749 (O_1749,N_19780,N_19768);
and UO_1750 (O_1750,N_19956,N_19842);
nand UO_1751 (O_1751,N_19622,N_19760);
nor UO_1752 (O_1752,N_19942,N_19630);
xnor UO_1753 (O_1753,N_19715,N_19964);
and UO_1754 (O_1754,N_19644,N_19743);
nor UO_1755 (O_1755,N_19811,N_19818);
xor UO_1756 (O_1756,N_19943,N_19873);
and UO_1757 (O_1757,N_19879,N_19994);
or UO_1758 (O_1758,N_19905,N_19845);
xnor UO_1759 (O_1759,N_19886,N_19861);
nor UO_1760 (O_1760,N_19920,N_19994);
nand UO_1761 (O_1761,N_19707,N_19699);
nor UO_1762 (O_1762,N_19996,N_19901);
nand UO_1763 (O_1763,N_19745,N_19920);
nand UO_1764 (O_1764,N_19612,N_19644);
xnor UO_1765 (O_1765,N_19948,N_19736);
or UO_1766 (O_1766,N_19605,N_19662);
nor UO_1767 (O_1767,N_19731,N_19747);
or UO_1768 (O_1768,N_19736,N_19710);
or UO_1769 (O_1769,N_19764,N_19974);
xnor UO_1770 (O_1770,N_19870,N_19809);
or UO_1771 (O_1771,N_19965,N_19858);
and UO_1772 (O_1772,N_19913,N_19782);
nor UO_1773 (O_1773,N_19833,N_19605);
and UO_1774 (O_1774,N_19668,N_19821);
xnor UO_1775 (O_1775,N_19845,N_19777);
nand UO_1776 (O_1776,N_19902,N_19831);
nor UO_1777 (O_1777,N_19642,N_19726);
nand UO_1778 (O_1778,N_19899,N_19835);
or UO_1779 (O_1779,N_19727,N_19659);
nand UO_1780 (O_1780,N_19662,N_19711);
nor UO_1781 (O_1781,N_19889,N_19888);
or UO_1782 (O_1782,N_19765,N_19667);
xnor UO_1783 (O_1783,N_19984,N_19735);
or UO_1784 (O_1784,N_19617,N_19807);
and UO_1785 (O_1785,N_19841,N_19657);
nor UO_1786 (O_1786,N_19642,N_19794);
nand UO_1787 (O_1787,N_19744,N_19651);
xnor UO_1788 (O_1788,N_19889,N_19856);
nand UO_1789 (O_1789,N_19693,N_19711);
or UO_1790 (O_1790,N_19700,N_19935);
nor UO_1791 (O_1791,N_19780,N_19714);
xor UO_1792 (O_1792,N_19676,N_19719);
and UO_1793 (O_1793,N_19606,N_19966);
nor UO_1794 (O_1794,N_19787,N_19696);
xnor UO_1795 (O_1795,N_19672,N_19883);
nor UO_1796 (O_1796,N_19634,N_19681);
or UO_1797 (O_1797,N_19791,N_19981);
or UO_1798 (O_1798,N_19646,N_19616);
xnor UO_1799 (O_1799,N_19871,N_19934);
and UO_1800 (O_1800,N_19756,N_19656);
xnor UO_1801 (O_1801,N_19833,N_19757);
nand UO_1802 (O_1802,N_19851,N_19903);
xnor UO_1803 (O_1803,N_19636,N_19607);
or UO_1804 (O_1804,N_19705,N_19666);
xor UO_1805 (O_1805,N_19794,N_19779);
xor UO_1806 (O_1806,N_19982,N_19616);
or UO_1807 (O_1807,N_19674,N_19997);
xor UO_1808 (O_1808,N_19735,N_19833);
nand UO_1809 (O_1809,N_19673,N_19911);
nand UO_1810 (O_1810,N_19636,N_19834);
xnor UO_1811 (O_1811,N_19660,N_19604);
xor UO_1812 (O_1812,N_19659,N_19807);
or UO_1813 (O_1813,N_19820,N_19963);
or UO_1814 (O_1814,N_19684,N_19921);
xnor UO_1815 (O_1815,N_19626,N_19908);
or UO_1816 (O_1816,N_19653,N_19849);
nor UO_1817 (O_1817,N_19617,N_19675);
xor UO_1818 (O_1818,N_19867,N_19822);
or UO_1819 (O_1819,N_19961,N_19964);
or UO_1820 (O_1820,N_19973,N_19734);
nor UO_1821 (O_1821,N_19763,N_19792);
and UO_1822 (O_1822,N_19895,N_19829);
and UO_1823 (O_1823,N_19877,N_19868);
nor UO_1824 (O_1824,N_19706,N_19685);
and UO_1825 (O_1825,N_19781,N_19842);
or UO_1826 (O_1826,N_19930,N_19747);
or UO_1827 (O_1827,N_19921,N_19612);
nor UO_1828 (O_1828,N_19820,N_19745);
or UO_1829 (O_1829,N_19735,N_19810);
and UO_1830 (O_1830,N_19654,N_19661);
or UO_1831 (O_1831,N_19731,N_19827);
or UO_1832 (O_1832,N_19920,N_19876);
and UO_1833 (O_1833,N_19665,N_19872);
or UO_1834 (O_1834,N_19816,N_19651);
nand UO_1835 (O_1835,N_19955,N_19604);
and UO_1836 (O_1836,N_19792,N_19645);
and UO_1837 (O_1837,N_19853,N_19626);
or UO_1838 (O_1838,N_19824,N_19983);
or UO_1839 (O_1839,N_19917,N_19948);
nor UO_1840 (O_1840,N_19619,N_19789);
and UO_1841 (O_1841,N_19754,N_19664);
xnor UO_1842 (O_1842,N_19900,N_19905);
xor UO_1843 (O_1843,N_19675,N_19754);
nand UO_1844 (O_1844,N_19838,N_19759);
and UO_1845 (O_1845,N_19879,N_19989);
nor UO_1846 (O_1846,N_19904,N_19679);
and UO_1847 (O_1847,N_19858,N_19998);
xnor UO_1848 (O_1848,N_19874,N_19730);
xnor UO_1849 (O_1849,N_19720,N_19836);
or UO_1850 (O_1850,N_19716,N_19801);
nor UO_1851 (O_1851,N_19822,N_19855);
and UO_1852 (O_1852,N_19748,N_19724);
nor UO_1853 (O_1853,N_19892,N_19669);
nand UO_1854 (O_1854,N_19660,N_19763);
nor UO_1855 (O_1855,N_19663,N_19722);
xor UO_1856 (O_1856,N_19806,N_19873);
xnor UO_1857 (O_1857,N_19980,N_19686);
or UO_1858 (O_1858,N_19854,N_19611);
and UO_1859 (O_1859,N_19729,N_19991);
nand UO_1860 (O_1860,N_19851,N_19668);
nor UO_1861 (O_1861,N_19891,N_19765);
xnor UO_1862 (O_1862,N_19636,N_19643);
and UO_1863 (O_1863,N_19631,N_19984);
and UO_1864 (O_1864,N_19800,N_19738);
or UO_1865 (O_1865,N_19902,N_19771);
nor UO_1866 (O_1866,N_19757,N_19891);
and UO_1867 (O_1867,N_19866,N_19742);
nor UO_1868 (O_1868,N_19814,N_19730);
nand UO_1869 (O_1869,N_19880,N_19924);
nand UO_1870 (O_1870,N_19824,N_19779);
and UO_1871 (O_1871,N_19961,N_19862);
xor UO_1872 (O_1872,N_19768,N_19809);
nand UO_1873 (O_1873,N_19980,N_19663);
and UO_1874 (O_1874,N_19985,N_19798);
nor UO_1875 (O_1875,N_19749,N_19920);
xor UO_1876 (O_1876,N_19638,N_19722);
nor UO_1877 (O_1877,N_19983,N_19800);
nor UO_1878 (O_1878,N_19712,N_19949);
and UO_1879 (O_1879,N_19772,N_19641);
or UO_1880 (O_1880,N_19682,N_19746);
nor UO_1881 (O_1881,N_19775,N_19949);
or UO_1882 (O_1882,N_19613,N_19880);
xor UO_1883 (O_1883,N_19986,N_19958);
or UO_1884 (O_1884,N_19712,N_19614);
nor UO_1885 (O_1885,N_19642,N_19859);
nor UO_1886 (O_1886,N_19650,N_19647);
and UO_1887 (O_1887,N_19930,N_19829);
nor UO_1888 (O_1888,N_19878,N_19650);
or UO_1889 (O_1889,N_19628,N_19739);
nand UO_1890 (O_1890,N_19724,N_19807);
or UO_1891 (O_1891,N_19767,N_19623);
nor UO_1892 (O_1892,N_19794,N_19652);
or UO_1893 (O_1893,N_19661,N_19636);
and UO_1894 (O_1894,N_19985,N_19780);
nor UO_1895 (O_1895,N_19856,N_19616);
nand UO_1896 (O_1896,N_19900,N_19736);
xnor UO_1897 (O_1897,N_19991,N_19704);
nor UO_1898 (O_1898,N_19881,N_19877);
xnor UO_1899 (O_1899,N_19947,N_19710);
and UO_1900 (O_1900,N_19748,N_19816);
nand UO_1901 (O_1901,N_19878,N_19890);
nand UO_1902 (O_1902,N_19630,N_19832);
nand UO_1903 (O_1903,N_19637,N_19845);
xnor UO_1904 (O_1904,N_19640,N_19759);
nand UO_1905 (O_1905,N_19779,N_19755);
nand UO_1906 (O_1906,N_19782,N_19752);
and UO_1907 (O_1907,N_19733,N_19671);
or UO_1908 (O_1908,N_19867,N_19821);
nor UO_1909 (O_1909,N_19817,N_19884);
and UO_1910 (O_1910,N_19703,N_19977);
nand UO_1911 (O_1911,N_19780,N_19914);
or UO_1912 (O_1912,N_19756,N_19824);
nor UO_1913 (O_1913,N_19978,N_19602);
nand UO_1914 (O_1914,N_19799,N_19760);
nor UO_1915 (O_1915,N_19961,N_19711);
or UO_1916 (O_1916,N_19775,N_19625);
nor UO_1917 (O_1917,N_19738,N_19820);
or UO_1918 (O_1918,N_19713,N_19792);
nand UO_1919 (O_1919,N_19925,N_19975);
or UO_1920 (O_1920,N_19990,N_19855);
or UO_1921 (O_1921,N_19957,N_19852);
nand UO_1922 (O_1922,N_19778,N_19788);
nor UO_1923 (O_1923,N_19778,N_19957);
or UO_1924 (O_1924,N_19674,N_19646);
nand UO_1925 (O_1925,N_19875,N_19674);
xnor UO_1926 (O_1926,N_19904,N_19678);
or UO_1927 (O_1927,N_19781,N_19946);
nand UO_1928 (O_1928,N_19622,N_19856);
and UO_1929 (O_1929,N_19605,N_19992);
or UO_1930 (O_1930,N_19765,N_19662);
or UO_1931 (O_1931,N_19921,N_19776);
or UO_1932 (O_1932,N_19785,N_19812);
nor UO_1933 (O_1933,N_19966,N_19998);
nand UO_1934 (O_1934,N_19947,N_19616);
nor UO_1935 (O_1935,N_19673,N_19894);
or UO_1936 (O_1936,N_19991,N_19982);
nor UO_1937 (O_1937,N_19931,N_19925);
nor UO_1938 (O_1938,N_19665,N_19627);
nand UO_1939 (O_1939,N_19814,N_19741);
or UO_1940 (O_1940,N_19983,N_19968);
nand UO_1941 (O_1941,N_19707,N_19921);
xor UO_1942 (O_1942,N_19689,N_19776);
and UO_1943 (O_1943,N_19826,N_19649);
nand UO_1944 (O_1944,N_19626,N_19865);
or UO_1945 (O_1945,N_19940,N_19787);
nand UO_1946 (O_1946,N_19862,N_19818);
xnor UO_1947 (O_1947,N_19777,N_19832);
nor UO_1948 (O_1948,N_19706,N_19695);
or UO_1949 (O_1949,N_19990,N_19833);
and UO_1950 (O_1950,N_19736,N_19938);
nor UO_1951 (O_1951,N_19826,N_19743);
or UO_1952 (O_1952,N_19607,N_19863);
nor UO_1953 (O_1953,N_19971,N_19964);
nor UO_1954 (O_1954,N_19702,N_19620);
and UO_1955 (O_1955,N_19810,N_19920);
or UO_1956 (O_1956,N_19979,N_19672);
or UO_1957 (O_1957,N_19978,N_19868);
xnor UO_1958 (O_1958,N_19778,N_19650);
nor UO_1959 (O_1959,N_19920,N_19677);
and UO_1960 (O_1960,N_19821,N_19755);
xor UO_1961 (O_1961,N_19714,N_19719);
nand UO_1962 (O_1962,N_19617,N_19627);
nand UO_1963 (O_1963,N_19922,N_19804);
nor UO_1964 (O_1964,N_19955,N_19812);
and UO_1965 (O_1965,N_19853,N_19808);
or UO_1966 (O_1966,N_19860,N_19791);
nor UO_1967 (O_1967,N_19808,N_19969);
nand UO_1968 (O_1968,N_19667,N_19970);
and UO_1969 (O_1969,N_19978,N_19794);
nor UO_1970 (O_1970,N_19978,N_19628);
xor UO_1971 (O_1971,N_19764,N_19766);
nor UO_1972 (O_1972,N_19809,N_19948);
and UO_1973 (O_1973,N_19725,N_19722);
or UO_1974 (O_1974,N_19867,N_19930);
xor UO_1975 (O_1975,N_19992,N_19981);
nand UO_1976 (O_1976,N_19705,N_19728);
and UO_1977 (O_1977,N_19843,N_19600);
xnor UO_1978 (O_1978,N_19734,N_19702);
nor UO_1979 (O_1979,N_19846,N_19948);
nand UO_1980 (O_1980,N_19988,N_19813);
xor UO_1981 (O_1981,N_19877,N_19748);
and UO_1982 (O_1982,N_19965,N_19859);
nand UO_1983 (O_1983,N_19981,N_19798);
or UO_1984 (O_1984,N_19873,N_19637);
nand UO_1985 (O_1985,N_19886,N_19764);
nand UO_1986 (O_1986,N_19787,N_19859);
xnor UO_1987 (O_1987,N_19784,N_19912);
xor UO_1988 (O_1988,N_19612,N_19898);
nor UO_1989 (O_1989,N_19624,N_19948);
and UO_1990 (O_1990,N_19950,N_19945);
or UO_1991 (O_1991,N_19605,N_19636);
nand UO_1992 (O_1992,N_19630,N_19796);
and UO_1993 (O_1993,N_19964,N_19903);
and UO_1994 (O_1994,N_19980,N_19956);
xnor UO_1995 (O_1995,N_19852,N_19759);
nand UO_1996 (O_1996,N_19720,N_19728);
nor UO_1997 (O_1997,N_19875,N_19738);
xor UO_1998 (O_1998,N_19716,N_19923);
nand UO_1999 (O_1999,N_19871,N_19638);
nand UO_2000 (O_2000,N_19986,N_19762);
nor UO_2001 (O_2001,N_19682,N_19666);
nand UO_2002 (O_2002,N_19753,N_19765);
xor UO_2003 (O_2003,N_19714,N_19977);
nand UO_2004 (O_2004,N_19656,N_19770);
or UO_2005 (O_2005,N_19804,N_19723);
or UO_2006 (O_2006,N_19821,N_19756);
nand UO_2007 (O_2007,N_19921,N_19920);
or UO_2008 (O_2008,N_19840,N_19921);
and UO_2009 (O_2009,N_19988,N_19934);
nand UO_2010 (O_2010,N_19626,N_19920);
nor UO_2011 (O_2011,N_19634,N_19897);
and UO_2012 (O_2012,N_19626,N_19695);
and UO_2013 (O_2013,N_19761,N_19600);
or UO_2014 (O_2014,N_19910,N_19807);
and UO_2015 (O_2015,N_19602,N_19636);
and UO_2016 (O_2016,N_19676,N_19718);
and UO_2017 (O_2017,N_19821,N_19982);
nor UO_2018 (O_2018,N_19675,N_19851);
nor UO_2019 (O_2019,N_19604,N_19883);
xor UO_2020 (O_2020,N_19732,N_19821);
xnor UO_2021 (O_2021,N_19922,N_19788);
and UO_2022 (O_2022,N_19808,N_19690);
nand UO_2023 (O_2023,N_19767,N_19846);
nor UO_2024 (O_2024,N_19737,N_19700);
or UO_2025 (O_2025,N_19967,N_19627);
or UO_2026 (O_2026,N_19780,N_19679);
and UO_2027 (O_2027,N_19682,N_19901);
or UO_2028 (O_2028,N_19743,N_19792);
nand UO_2029 (O_2029,N_19626,N_19705);
nand UO_2030 (O_2030,N_19802,N_19785);
nor UO_2031 (O_2031,N_19712,N_19757);
xnor UO_2032 (O_2032,N_19640,N_19770);
and UO_2033 (O_2033,N_19939,N_19630);
nand UO_2034 (O_2034,N_19936,N_19863);
xor UO_2035 (O_2035,N_19735,N_19807);
nand UO_2036 (O_2036,N_19969,N_19616);
and UO_2037 (O_2037,N_19984,N_19976);
nor UO_2038 (O_2038,N_19978,N_19882);
xnor UO_2039 (O_2039,N_19886,N_19825);
or UO_2040 (O_2040,N_19727,N_19688);
nand UO_2041 (O_2041,N_19629,N_19879);
and UO_2042 (O_2042,N_19678,N_19966);
and UO_2043 (O_2043,N_19700,N_19664);
nand UO_2044 (O_2044,N_19756,N_19638);
nor UO_2045 (O_2045,N_19658,N_19752);
and UO_2046 (O_2046,N_19726,N_19603);
and UO_2047 (O_2047,N_19612,N_19876);
xnor UO_2048 (O_2048,N_19758,N_19920);
nand UO_2049 (O_2049,N_19811,N_19659);
or UO_2050 (O_2050,N_19638,N_19954);
or UO_2051 (O_2051,N_19862,N_19805);
nor UO_2052 (O_2052,N_19948,N_19819);
and UO_2053 (O_2053,N_19933,N_19847);
nor UO_2054 (O_2054,N_19889,N_19693);
xnor UO_2055 (O_2055,N_19665,N_19676);
or UO_2056 (O_2056,N_19621,N_19816);
xnor UO_2057 (O_2057,N_19775,N_19749);
or UO_2058 (O_2058,N_19968,N_19645);
nor UO_2059 (O_2059,N_19731,N_19781);
nand UO_2060 (O_2060,N_19991,N_19748);
and UO_2061 (O_2061,N_19650,N_19602);
nor UO_2062 (O_2062,N_19744,N_19962);
nor UO_2063 (O_2063,N_19654,N_19694);
and UO_2064 (O_2064,N_19701,N_19654);
nor UO_2065 (O_2065,N_19804,N_19724);
xnor UO_2066 (O_2066,N_19854,N_19993);
or UO_2067 (O_2067,N_19878,N_19851);
or UO_2068 (O_2068,N_19959,N_19919);
or UO_2069 (O_2069,N_19883,N_19954);
or UO_2070 (O_2070,N_19873,N_19991);
xor UO_2071 (O_2071,N_19966,N_19628);
and UO_2072 (O_2072,N_19747,N_19994);
and UO_2073 (O_2073,N_19724,N_19658);
nand UO_2074 (O_2074,N_19607,N_19687);
nor UO_2075 (O_2075,N_19928,N_19829);
or UO_2076 (O_2076,N_19929,N_19997);
xnor UO_2077 (O_2077,N_19736,N_19789);
and UO_2078 (O_2078,N_19795,N_19816);
xnor UO_2079 (O_2079,N_19775,N_19991);
and UO_2080 (O_2080,N_19652,N_19739);
nor UO_2081 (O_2081,N_19602,N_19709);
and UO_2082 (O_2082,N_19991,N_19689);
and UO_2083 (O_2083,N_19622,N_19728);
and UO_2084 (O_2084,N_19785,N_19913);
or UO_2085 (O_2085,N_19752,N_19991);
nor UO_2086 (O_2086,N_19973,N_19982);
nor UO_2087 (O_2087,N_19645,N_19966);
nand UO_2088 (O_2088,N_19607,N_19816);
nor UO_2089 (O_2089,N_19771,N_19960);
xnor UO_2090 (O_2090,N_19741,N_19894);
nor UO_2091 (O_2091,N_19962,N_19614);
nor UO_2092 (O_2092,N_19671,N_19627);
or UO_2093 (O_2093,N_19778,N_19733);
or UO_2094 (O_2094,N_19959,N_19617);
xnor UO_2095 (O_2095,N_19715,N_19709);
or UO_2096 (O_2096,N_19941,N_19746);
nand UO_2097 (O_2097,N_19978,N_19739);
nor UO_2098 (O_2098,N_19856,N_19894);
nor UO_2099 (O_2099,N_19783,N_19819);
nand UO_2100 (O_2100,N_19681,N_19814);
and UO_2101 (O_2101,N_19797,N_19772);
nor UO_2102 (O_2102,N_19945,N_19830);
nor UO_2103 (O_2103,N_19981,N_19746);
xor UO_2104 (O_2104,N_19771,N_19664);
nand UO_2105 (O_2105,N_19849,N_19927);
nand UO_2106 (O_2106,N_19801,N_19721);
xor UO_2107 (O_2107,N_19687,N_19630);
nor UO_2108 (O_2108,N_19896,N_19856);
xor UO_2109 (O_2109,N_19666,N_19655);
xnor UO_2110 (O_2110,N_19827,N_19695);
or UO_2111 (O_2111,N_19743,N_19976);
and UO_2112 (O_2112,N_19921,N_19654);
xor UO_2113 (O_2113,N_19983,N_19716);
nand UO_2114 (O_2114,N_19709,N_19802);
nand UO_2115 (O_2115,N_19602,N_19779);
xnor UO_2116 (O_2116,N_19622,N_19645);
nor UO_2117 (O_2117,N_19978,N_19983);
or UO_2118 (O_2118,N_19725,N_19642);
and UO_2119 (O_2119,N_19794,N_19721);
xnor UO_2120 (O_2120,N_19724,N_19751);
nor UO_2121 (O_2121,N_19727,N_19915);
nand UO_2122 (O_2122,N_19648,N_19984);
or UO_2123 (O_2123,N_19912,N_19899);
or UO_2124 (O_2124,N_19923,N_19681);
and UO_2125 (O_2125,N_19709,N_19945);
nor UO_2126 (O_2126,N_19871,N_19891);
or UO_2127 (O_2127,N_19997,N_19673);
or UO_2128 (O_2128,N_19652,N_19648);
and UO_2129 (O_2129,N_19675,N_19630);
xnor UO_2130 (O_2130,N_19710,N_19664);
and UO_2131 (O_2131,N_19775,N_19646);
and UO_2132 (O_2132,N_19733,N_19692);
nor UO_2133 (O_2133,N_19928,N_19780);
nand UO_2134 (O_2134,N_19654,N_19834);
nor UO_2135 (O_2135,N_19852,N_19800);
or UO_2136 (O_2136,N_19623,N_19747);
or UO_2137 (O_2137,N_19905,N_19766);
nor UO_2138 (O_2138,N_19628,N_19941);
nor UO_2139 (O_2139,N_19946,N_19707);
xor UO_2140 (O_2140,N_19620,N_19710);
nand UO_2141 (O_2141,N_19665,N_19733);
xor UO_2142 (O_2142,N_19850,N_19698);
or UO_2143 (O_2143,N_19780,N_19748);
nor UO_2144 (O_2144,N_19775,N_19744);
or UO_2145 (O_2145,N_19660,N_19991);
xnor UO_2146 (O_2146,N_19853,N_19734);
and UO_2147 (O_2147,N_19886,N_19941);
or UO_2148 (O_2148,N_19891,N_19797);
xor UO_2149 (O_2149,N_19618,N_19833);
xor UO_2150 (O_2150,N_19848,N_19769);
and UO_2151 (O_2151,N_19963,N_19975);
nor UO_2152 (O_2152,N_19614,N_19871);
and UO_2153 (O_2153,N_19804,N_19614);
nand UO_2154 (O_2154,N_19676,N_19646);
nand UO_2155 (O_2155,N_19758,N_19654);
xor UO_2156 (O_2156,N_19759,N_19870);
xnor UO_2157 (O_2157,N_19769,N_19913);
xnor UO_2158 (O_2158,N_19917,N_19964);
nand UO_2159 (O_2159,N_19714,N_19816);
nand UO_2160 (O_2160,N_19822,N_19674);
or UO_2161 (O_2161,N_19967,N_19616);
or UO_2162 (O_2162,N_19967,N_19762);
nand UO_2163 (O_2163,N_19815,N_19915);
xnor UO_2164 (O_2164,N_19992,N_19925);
or UO_2165 (O_2165,N_19605,N_19747);
or UO_2166 (O_2166,N_19963,N_19978);
nor UO_2167 (O_2167,N_19863,N_19999);
and UO_2168 (O_2168,N_19936,N_19860);
or UO_2169 (O_2169,N_19874,N_19818);
nand UO_2170 (O_2170,N_19670,N_19875);
xor UO_2171 (O_2171,N_19689,N_19945);
nor UO_2172 (O_2172,N_19883,N_19964);
or UO_2173 (O_2173,N_19636,N_19816);
nor UO_2174 (O_2174,N_19709,N_19796);
or UO_2175 (O_2175,N_19775,N_19717);
nand UO_2176 (O_2176,N_19750,N_19918);
xnor UO_2177 (O_2177,N_19890,N_19871);
and UO_2178 (O_2178,N_19765,N_19794);
nor UO_2179 (O_2179,N_19984,N_19914);
nor UO_2180 (O_2180,N_19856,N_19799);
and UO_2181 (O_2181,N_19631,N_19993);
nor UO_2182 (O_2182,N_19676,N_19673);
and UO_2183 (O_2183,N_19994,N_19653);
nor UO_2184 (O_2184,N_19720,N_19609);
xor UO_2185 (O_2185,N_19779,N_19846);
and UO_2186 (O_2186,N_19632,N_19619);
nor UO_2187 (O_2187,N_19982,N_19863);
or UO_2188 (O_2188,N_19772,N_19932);
or UO_2189 (O_2189,N_19804,N_19727);
or UO_2190 (O_2190,N_19822,N_19914);
and UO_2191 (O_2191,N_19938,N_19940);
or UO_2192 (O_2192,N_19681,N_19691);
xnor UO_2193 (O_2193,N_19941,N_19737);
nand UO_2194 (O_2194,N_19957,N_19763);
xnor UO_2195 (O_2195,N_19705,N_19641);
or UO_2196 (O_2196,N_19789,N_19841);
and UO_2197 (O_2197,N_19697,N_19958);
or UO_2198 (O_2198,N_19867,N_19620);
or UO_2199 (O_2199,N_19656,N_19808);
and UO_2200 (O_2200,N_19832,N_19618);
xor UO_2201 (O_2201,N_19904,N_19890);
xnor UO_2202 (O_2202,N_19970,N_19609);
or UO_2203 (O_2203,N_19893,N_19790);
xnor UO_2204 (O_2204,N_19618,N_19663);
xor UO_2205 (O_2205,N_19711,N_19950);
nand UO_2206 (O_2206,N_19824,N_19646);
xnor UO_2207 (O_2207,N_19962,N_19806);
xor UO_2208 (O_2208,N_19982,N_19795);
or UO_2209 (O_2209,N_19714,N_19843);
xor UO_2210 (O_2210,N_19863,N_19738);
xor UO_2211 (O_2211,N_19605,N_19606);
xnor UO_2212 (O_2212,N_19866,N_19871);
nand UO_2213 (O_2213,N_19629,N_19970);
xor UO_2214 (O_2214,N_19899,N_19947);
nor UO_2215 (O_2215,N_19763,N_19876);
nor UO_2216 (O_2216,N_19936,N_19646);
xor UO_2217 (O_2217,N_19669,N_19695);
nand UO_2218 (O_2218,N_19874,N_19779);
and UO_2219 (O_2219,N_19861,N_19619);
or UO_2220 (O_2220,N_19793,N_19891);
or UO_2221 (O_2221,N_19856,N_19658);
nand UO_2222 (O_2222,N_19772,N_19894);
nand UO_2223 (O_2223,N_19987,N_19612);
nor UO_2224 (O_2224,N_19742,N_19680);
or UO_2225 (O_2225,N_19629,N_19623);
nand UO_2226 (O_2226,N_19740,N_19775);
and UO_2227 (O_2227,N_19914,N_19916);
nor UO_2228 (O_2228,N_19648,N_19798);
nand UO_2229 (O_2229,N_19996,N_19890);
nand UO_2230 (O_2230,N_19853,N_19828);
nor UO_2231 (O_2231,N_19668,N_19833);
and UO_2232 (O_2232,N_19615,N_19738);
xnor UO_2233 (O_2233,N_19745,N_19868);
nor UO_2234 (O_2234,N_19684,N_19971);
and UO_2235 (O_2235,N_19783,N_19972);
xnor UO_2236 (O_2236,N_19845,N_19761);
nand UO_2237 (O_2237,N_19619,N_19808);
or UO_2238 (O_2238,N_19905,N_19755);
or UO_2239 (O_2239,N_19979,N_19927);
nand UO_2240 (O_2240,N_19600,N_19821);
or UO_2241 (O_2241,N_19679,N_19961);
nor UO_2242 (O_2242,N_19806,N_19760);
xnor UO_2243 (O_2243,N_19870,N_19995);
or UO_2244 (O_2244,N_19717,N_19822);
and UO_2245 (O_2245,N_19900,N_19797);
and UO_2246 (O_2246,N_19646,N_19990);
and UO_2247 (O_2247,N_19665,N_19949);
or UO_2248 (O_2248,N_19731,N_19997);
nor UO_2249 (O_2249,N_19696,N_19666);
and UO_2250 (O_2250,N_19895,N_19722);
nor UO_2251 (O_2251,N_19860,N_19849);
or UO_2252 (O_2252,N_19611,N_19765);
or UO_2253 (O_2253,N_19765,N_19824);
and UO_2254 (O_2254,N_19655,N_19844);
nand UO_2255 (O_2255,N_19804,N_19986);
nand UO_2256 (O_2256,N_19755,N_19681);
xor UO_2257 (O_2257,N_19613,N_19762);
nor UO_2258 (O_2258,N_19630,N_19766);
and UO_2259 (O_2259,N_19646,N_19955);
or UO_2260 (O_2260,N_19854,N_19982);
nor UO_2261 (O_2261,N_19729,N_19801);
and UO_2262 (O_2262,N_19813,N_19676);
nand UO_2263 (O_2263,N_19923,N_19974);
or UO_2264 (O_2264,N_19943,N_19882);
nand UO_2265 (O_2265,N_19906,N_19824);
nand UO_2266 (O_2266,N_19961,N_19920);
or UO_2267 (O_2267,N_19707,N_19822);
nand UO_2268 (O_2268,N_19609,N_19674);
nand UO_2269 (O_2269,N_19974,N_19899);
nor UO_2270 (O_2270,N_19789,N_19630);
or UO_2271 (O_2271,N_19910,N_19806);
xnor UO_2272 (O_2272,N_19790,N_19827);
xnor UO_2273 (O_2273,N_19975,N_19848);
nand UO_2274 (O_2274,N_19708,N_19730);
nor UO_2275 (O_2275,N_19832,N_19648);
nor UO_2276 (O_2276,N_19961,N_19919);
and UO_2277 (O_2277,N_19672,N_19978);
nand UO_2278 (O_2278,N_19962,N_19761);
or UO_2279 (O_2279,N_19813,N_19956);
xnor UO_2280 (O_2280,N_19902,N_19710);
and UO_2281 (O_2281,N_19875,N_19914);
nor UO_2282 (O_2282,N_19743,N_19786);
nor UO_2283 (O_2283,N_19872,N_19770);
or UO_2284 (O_2284,N_19611,N_19621);
or UO_2285 (O_2285,N_19660,N_19821);
or UO_2286 (O_2286,N_19727,N_19760);
nand UO_2287 (O_2287,N_19982,N_19654);
nand UO_2288 (O_2288,N_19776,N_19769);
xor UO_2289 (O_2289,N_19744,N_19710);
and UO_2290 (O_2290,N_19661,N_19674);
nand UO_2291 (O_2291,N_19636,N_19889);
nand UO_2292 (O_2292,N_19968,N_19927);
or UO_2293 (O_2293,N_19927,N_19730);
and UO_2294 (O_2294,N_19872,N_19903);
nand UO_2295 (O_2295,N_19849,N_19733);
xor UO_2296 (O_2296,N_19720,N_19635);
or UO_2297 (O_2297,N_19989,N_19874);
nand UO_2298 (O_2298,N_19642,N_19782);
xor UO_2299 (O_2299,N_19834,N_19907);
nor UO_2300 (O_2300,N_19659,N_19775);
or UO_2301 (O_2301,N_19624,N_19630);
nand UO_2302 (O_2302,N_19956,N_19992);
nand UO_2303 (O_2303,N_19746,N_19687);
xnor UO_2304 (O_2304,N_19878,N_19930);
nand UO_2305 (O_2305,N_19711,N_19649);
or UO_2306 (O_2306,N_19772,N_19753);
and UO_2307 (O_2307,N_19775,N_19791);
or UO_2308 (O_2308,N_19618,N_19672);
or UO_2309 (O_2309,N_19991,N_19618);
and UO_2310 (O_2310,N_19720,N_19956);
or UO_2311 (O_2311,N_19638,N_19961);
nand UO_2312 (O_2312,N_19742,N_19806);
and UO_2313 (O_2313,N_19789,N_19636);
or UO_2314 (O_2314,N_19936,N_19752);
nor UO_2315 (O_2315,N_19895,N_19724);
xor UO_2316 (O_2316,N_19923,N_19744);
xor UO_2317 (O_2317,N_19944,N_19828);
or UO_2318 (O_2318,N_19948,N_19654);
xnor UO_2319 (O_2319,N_19967,N_19769);
xor UO_2320 (O_2320,N_19826,N_19874);
nand UO_2321 (O_2321,N_19912,N_19862);
or UO_2322 (O_2322,N_19820,N_19819);
nor UO_2323 (O_2323,N_19739,N_19738);
nand UO_2324 (O_2324,N_19665,N_19734);
nor UO_2325 (O_2325,N_19740,N_19665);
or UO_2326 (O_2326,N_19640,N_19807);
nor UO_2327 (O_2327,N_19705,N_19762);
nor UO_2328 (O_2328,N_19703,N_19604);
xor UO_2329 (O_2329,N_19691,N_19731);
nor UO_2330 (O_2330,N_19804,N_19656);
or UO_2331 (O_2331,N_19963,N_19934);
and UO_2332 (O_2332,N_19809,N_19618);
xor UO_2333 (O_2333,N_19871,N_19692);
xor UO_2334 (O_2334,N_19713,N_19722);
nor UO_2335 (O_2335,N_19654,N_19988);
nand UO_2336 (O_2336,N_19670,N_19899);
xor UO_2337 (O_2337,N_19990,N_19963);
xnor UO_2338 (O_2338,N_19988,N_19853);
and UO_2339 (O_2339,N_19738,N_19935);
nand UO_2340 (O_2340,N_19896,N_19870);
nand UO_2341 (O_2341,N_19779,N_19796);
nor UO_2342 (O_2342,N_19753,N_19844);
nor UO_2343 (O_2343,N_19795,N_19955);
nor UO_2344 (O_2344,N_19849,N_19631);
and UO_2345 (O_2345,N_19687,N_19875);
nor UO_2346 (O_2346,N_19985,N_19692);
nor UO_2347 (O_2347,N_19719,N_19973);
or UO_2348 (O_2348,N_19694,N_19843);
or UO_2349 (O_2349,N_19626,N_19815);
or UO_2350 (O_2350,N_19675,N_19662);
nor UO_2351 (O_2351,N_19604,N_19634);
nor UO_2352 (O_2352,N_19824,N_19697);
xor UO_2353 (O_2353,N_19819,N_19851);
or UO_2354 (O_2354,N_19820,N_19780);
or UO_2355 (O_2355,N_19721,N_19672);
nor UO_2356 (O_2356,N_19628,N_19710);
nor UO_2357 (O_2357,N_19671,N_19679);
xor UO_2358 (O_2358,N_19967,N_19685);
and UO_2359 (O_2359,N_19692,N_19939);
and UO_2360 (O_2360,N_19915,N_19788);
nor UO_2361 (O_2361,N_19853,N_19955);
and UO_2362 (O_2362,N_19990,N_19725);
nor UO_2363 (O_2363,N_19903,N_19812);
and UO_2364 (O_2364,N_19734,N_19842);
xor UO_2365 (O_2365,N_19776,N_19984);
nand UO_2366 (O_2366,N_19828,N_19707);
or UO_2367 (O_2367,N_19946,N_19860);
nor UO_2368 (O_2368,N_19600,N_19647);
or UO_2369 (O_2369,N_19846,N_19642);
nand UO_2370 (O_2370,N_19721,N_19919);
and UO_2371 (O_2371,N_19709,N_19654);
xor UO_2372 (O_2372,N_19840,N_19848);
and UO_2373 (O_2373,N_19895,N_19745);
nand UO_2374 (O_2374,N_19951,N_19648);
and UO_2375 (O_2375,N_19996,N_19988);
nand UO_2376 (O_2376,N_19645,N_19794);
xor UO_2377 (O_2377,N_19794,N_19938);
nor UO_2378 (O_2378,N_19770,N_19746);
or UO_2379 (O_2379,N_19659,N_19828);
nand UO_2380 (O_2380,N_19899,N_19940);
nor UO_2381 (O_2381,N_19795,N_19637);
xor UO_2382 (O_2382,N_19988,N_19752);
and UO_2383 (O_2383,N_19714,N_19753);
nand UO_2384 (O_2384,N_19766,N_19719);
nor UO_2385 (O_2385,N_19880,N_19948);
and UO_2386 (O_2386,N_19728,N_19608);
nand UO_2387 (O_2387,N_19859,N_19973);
nor UO_2388 (O_2388,N_19774,N_19720);
xnor UO_2389 (O_2389,N_19735,N_19947);
nor UO_2390 (O_2390,N_19934,N_19961);
or UO_2391 (O_2391,N_19911,N_19651);
and UO_2392 (O_2392,N_19810,N_19966);
and UO_2393 (O_2393,N_19624,N_19641);
xor UO_2394 (O_2394,N_19788,N_19899);
xor UO_2395 (O_2395,N_19784,N_19670);
xor UO_2396 (O_2396,N_19702,N_19862);
and UO_2397 (O_2397,N_19696,N_19872);
nand UO_2398 (O_2398,N_19826,N_19619);
or UO_2399 (O_2399,N_19893,N_19678);
and UO_2400 (O_2400,N_19922,N_19797);
nor UO_2401 (O_2401,N_19626,N_19866);
or UO_2402 (O_2402,N_19829,N_19606);
nand UO_2403 (O_2403,N_19878,N_19843);
nand UO_2404 (O_2404,N_19816,N_19969);
xor UO_2405 (O_2405,N_19692,N_19937);
nor UO_2406 (O_2406,N_19943,N_19960);
or UO_2407 (O_2407,N_19638,N_19949);
nor UO_2408 (O_2408,N_19897,N_19989);
or UO_2409 (O_2409,N_19925,N_19829);
or UO_2410 (O_2410,N_19855,N_19983);
or UO_2411 (O_2411,N_19642,N_19790);
nand UO_2412 (O_2412,N_19906,N_19903);
nand UO_2413 (O_2413,N_19880,N_19681);
xnor UO_2414 (O_2414,N_19778,N_19972);
xor UO_2415 (O_2415,N_19983,N_19645);
and UO_2416 (O_2416,N_19716,N_19610);
xor UO_2417 (O_2417,N_19863,N_19906);
or UO_2418 (O_2418,N_19843,N_19876);
nand UO_2419 (O_2419,N_19848,N_19721);
and UO_2420 (O_2420,N_19749,N_19984);
or UO_2421 (O_2421,N_19886,N_19687);
nor UO_2422 (O_2422,N_19735,N_19647);
nor UO_2423 (O_2423,N_19985,N_19921);
xnor UO_2424 (O_2424,N_19811,N_19935);
xnor UO_2425 (O_2425,N_19860,N_19719);
and UO_2426 (O_2426,N_19784,N_19736);
or UO_2427 (O_2427,N_19702,N_19653);
or UO_2428 (O_2428,N_19645,N_19804);
and UO_2429 (O_2429,N_19669,N_19900);
nor UO_2430 (O_2430,N_19856,N_19665);
nor UO_2431 (O_2431,N_19905,N_19811);
xor UO_2432 (O_2432,N_19994,N_19799);
nor UO_2433 (O_2433,N_19845,N_19693);
or UO_2434 (O_2434,N_19885,N_19671);
and UO_2435 (O_2435,N_19974,N_19609);
nor UO_2436 (O_2436,N_19948,N_19812);
or UO_2437 (O_2437,N_19653,N_19820);
and UO_2438 (O_2438,N_19708,N_19637);
nand UO_2439 (O_2439,N_19811,N_19680);
nor UO_2440 (O_2440,N_19653,N_19833);
nor UO_2441 (O_2441,N_19794,N_19740);
xnor UO_2442 (O_2442,N_19626,N_19842);
and UO_2443 (O_2443,N_19669,N_19707);
or UO_2444 (O_2444,N_19953,N_19884);
xor UO_2445 (O_2445,N_19842,N_19624);
nor UO_2446 (O_2446,N_19761,N_19769);
xnor UO_2447 (O_2447,N_19923,N_19728);
nor UO_2448 (O_2448,N_19815,N_19877);
nand UO_2449 (O_2449,N_19958,N_19671);
xnor UO_2450 (O_2450,N_19859,N_19884);
and UO_2451 (O_2451,N_19724,N_19967);
nand UO_2452 (O_2452,N_19847,N_19980);
and UO_2453 (O_2453,N_19909,N_19929);
or UO_2454 (O_2454,N_19975,N_19970);
or UO_2455 (O_2455,N_19863,N_19840);
or UO_2456 (O_2456,N_19674,N_19956);
nor UO_2457 (O_2457,N_19686,N_19609);
nand UO_2458 (O_2458,N_19996,N_19984);
nor UO_2459 (O_2459,N_19611,N_19771);
nor UO_2460 (O_2460,N_19829,N_19624);
xor UO_2461 (O_2461,N_19769,N_19772);
nand UO_2462 (O_2462,N_19614,N_19820);
or UO_2463 (O_2463,N_19798,N_19601);
nor UO_2464 (O_2464,N_19604,N_19610);
nand UO_2465 (O_2465,N_19905,N_19846);
and UO_2466 (O_2466,N_19987,N_19613);
xnor UO_2467 (O_2467,N_19879,N_19669);
xor UO_2468 (O_2468,N_19825,N_19685);
or UO_2469 (O_2469,N_19629,N_19853);
or UO_2470 (O_2470,N_19689,N_19858);
nor UO_2471 (O_2471,N_19664,N_19802);
or UO_2472 (O_2472,N_19963,N_19762);
or UO_2473 (O_2473,N_19964,N_19829);
xnor UO_2474 (O_2474,N_19675,N_19928);
and UO_2475 (O_2475,N_19948,N_19799);
or UO_2476 (O_2476,N_19766,N_19725);
nor UO_2477 (O_2477,N_19625,N_19759);
nor UO_2478 (O_2478,N_19775,N_19757);
nor UO_2479 (O_2479,N_19915,N_19734);
or UO_2480 (O_2480,N_19786,N_19807);
or UO_2481 (O_2481,N_19742,N_19687);
or UO_2482 (O_2482,N_19784,N_19898);
nand UO_2483 (O_2483,N_19996,N_19891);
or UO_2484 (O_2484,N_19752,N_19984);
xor UO_2485 (O_2485,N_19808,N_19783);
and UO_2486 (O_2486,N_19857,N_19685);
xor UO_2487 (O_2487,N_19601,N_19829);
xor UO_2488 (O_2488,N_19785,N_19765);
nand UO_2489 (O_2489,N_19775,N_19990);
or UO_2490 (O_2490,N_19605,N_19975);
xnor UO_2491 (O_2491,N_19625,N_19962);
and UO_2492 (O_2492,N_19605,N_19980);
and UO_2493 (O_2493,N_19999,N_19877);
xnor UO_2494 (O_2494,N_19696,N_19615);
xor UO_2495 (O_2495,N_19885,N_19724);
nand UO_2496 (O_2496,N_19861,N_19734);
nor UO_2497 (O_2497,N_19762,N_19782);
nor UO_2498 (O_2498,N_19896,N_19836);
nor UO_2499 (O_2499,N_19744,N_19931);
endmodule