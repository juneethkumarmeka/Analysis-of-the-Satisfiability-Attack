module basic_500_3000_500_6_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_214,In_196);
and U1 (N_1,In_493,In_10);
nand U2 (N_2,In_295,In_387);
nand U3 (N_3,In_421,In_277);
and U4 (N_4,In_301,In_153);
nand U5 (N_5,In_152,In_81);
nor U6 (N_6,In_477,In_429);
nand U7 (N_7,In_275,In_341);
and U8 (N_8,In_417,In_130);
nand U9 (N_9,In_18,In_405);
nand U10 (N_10,In_229,In_476);
or U11 (N_11,In_172,In_423);
or U12 (N_12,In_7,In_372);
nor U13 (N_13,In_98,In_350);
nand U14 (N_14,In_95,In_159);
nor U15 (N_15,In_227,In_288);
nor U16 (N_16,In_323,In_237);
and U17 (N_17,In_435,In_15);
nor U18 (N_18,In_106,In_117);
nor U19 (N_19,In_382,In_182);
and U20 (N_20,In_384,In_321);
nand U21 (N_21,In_120,In_238);
nor U22 (N_22,In_254,In_151);
nand U23 (N_23,In_181,In_201);
and U24 (N_24,In_378,In_426);
nand U25 (N_25,In_99,In_162);
and U26 (N_26,In_441,In_428);
nor U27 (N_27,In_290,In_313);
nand U28 (N_28,In_243,In_217);
or U29 (N_29,In_444,In_221);
nand U30 (N_30,In_498,In_17);
and U31 (N_31,In_209,In_205);
and U32 (N_32,In_414,In_434);
xnor U33 (N_33,In_128,In_266);
nor U34 (N_34,In_80,In_94);
and U35 (N_35,In_83,In_215);
and U36 (N_36,In_459,In_482);
nand U37 (N_37,In_442,In_241);
xor U38 (N_38,In_346,In_437);
nand U39 (N_39,In_456,In_294);
xor U40 (N_40,In_85,In_291);
or U41 (N_41,In_9,In_416);
nor U42 (N_42,In_267,In_143);
nand U43 (N_43,In_96,In_269);
xor U44 (N_44,In_110,In_61);
and U45 (N_45,In_486,In_474);
or U46 (N_46,In_169,In_413);
and U47 (N_47,In_150,In_121);
xor U48 (N_48,In_166,In_114);
and U49 (N_49,In_395,In_379);
nand U50 (N_50,In_145,In_282);
nand U51 (N_51,In_1,In_411);
xor U52 (N_52,In_90,In_102);
and U53 (N_53,In_67,In_357);
and U54 (N_54,In_356,In_156);
and U55 (N_55,In_298,In_133);
or U56 (N_56,In_163,In_213);
xnor U57 (N_57,In_125,In_144);
or U58 (N_58,In_33,In_281);
or U59 (N_59,In_412,In_19);
nor U60 (N_60,In_306,In_367);
nor U61 (N_61,In_257,In_70);
or U62 (N_62,In_154,In_253);
and U63 (N_63,In_390,In_72);
nand U64 (N_64,In_119,In_101);
and U65 (N_65,In_135,In_465);
nor U66 (N_66,In_364,In_28);
nand U67 (N_67,In_250,In_158);
nor U68 (N_68,In_147,In_419);
nor U69 (N_69,In_6,In_11);
nand U70 (N_70,In_82,In_433);
nand U71 (N_71,In_199,In_293);
nand U72 (N_72,In_25,In_249);
or U73 (N_73,In_161,In_454);
nand U74 (N_74,In_193,In_400);
or U75 (N_75,In_328,In_363);
nor U76 (N_76,In_60,In_348);
or U77 (N_77,In_463,In_78);
nor U78 (N_78,In_491,In_483);
or U79 (N_79,In_409,In_452);
and U80 (N_80,In_109,In_113);
nor U81 (N_81,In_351,In_494);
and U82 (N_82,In_183,In_418);
nor U83 (N_83,In_475,In_338);
nand U84 (N_84,In_189,In_402);
or U85 (N_85,In_398,In_297);
nor U86 (N_86,In_174,In_289);
or U87 (N_87,In_79,In_30);
and U88 (N_88,In_165,In_440);
nor U89 (N_89,In_232,In_93);
or U90 (N_90,In_479,In_29);
nor U91 (N_91,In_252,In_100);
nor U92 (N_92,In_342,In_256);
xnor U93 (N_93,In_26,In_74);
nand U94 (N_94,In_54,In_103);
or U95 (N_95,In_233,In_311);
and U96 (N_96,In_484,In_447);
xor U97 (N_97,In_322,In_24);
nand U98 (N_98,In_432,In_271);
or U99 (N_99,In_450,In_198);
nand U100 (N_100,In_222,In_326);
and U101 (N_101,In_68,In_31);
or U102 (N_102,In_499,In_284);
nand U103 (N_103,In_137,In_138);
and U104 (N_104,In_122,In_404);
xor U105 (N_105,In_263,In_470);
or U106 (N_106,In_292,In_131);
nand U107 (N_107,In_49,In_126);
nand U108 (N_108,In_425,In_64);
nor U109 (N_109,In_139,In_449);
nor U110 (N_110,In_420,In_365);
or U111 (N_111,In_343,In_300);
or U112 (N_112,In_280,In_206);
and U113 (N_113,In_200,In_88);
nor U114 (N_114,In_468,In_220);
nand U115 (N_115,In_488,In_248);
and U116 (N_116,In_388,In_191);
nand U117 (N_117,In_71,In_337);
nor U118 (N_118,In_273,In_391);
nand U119 (N_119,In_264,In_230);
and U120 (N_120,In_132,In_448);
or U121 (N_121,In_473,In_308);
xor U122 (N_122,In_329,In_140);
or U123 (N_123,In_204,In_335);
nand U124 (N_124,In_92,In_492);
nand U125 (N_125,In_176,In_251);
or U126 (N_126,In_0,In_164);
nand U127 (N_127,In_286,In_385);
nand U128 (N_128,In_146,In_353);
nand U129 (N_129,In_123,In_23);
nor U130 (N_130,In_345,In_389);
nand U131 (N_131,In_44,In_401);
nand U132 (N_132,In_369,In_236);
nor U133 (N_133,In_407,In_12);
xnor U134 (N_134,In_481,In_272);
nand U135 (N_135,In_39,In_157);
nor U136 (N_136,In_36,In_246);
nand U137 (N_137,In_55,In_320);
nand U138 (N_138,In_324,In_490);
or U139 (N_139,In_279,In_394);
and U140 (N_140,In_406,In_50);
or U141 (N_141,In_155,In_489);
and U142 (N_142,In_334,In_14);
or U143 (N_143,In_265,In_259);
xnor U144 (N_144,In_118,In_467);
nor U145 (N_145,In_2,In_455);
nor U146 (N_146,In_453,In_462);
and U147 (N_147,In_330,In_360);
and U148 (N_148,In_315,In_192);
or U149 (N_149,In_410,In_276);
or U150 (N_150,In_312,In_469);
and U151 (N_151,In_53,In_149);
and U152 (N_152,In_278,In_376);
or U153 (N_153,In_141,In_45);
and U154 (N_154,In_299,In_66);
or U155 (N_155,In_124,In_202);
and U156 (N_156,In_208,In_16);
xor U157 (N_157,In_451,In_42);
and U158 (N_158,In_347,In_244);
nor U159 (N_159,In_325,In_5);
nor U160 (N_160,In_47,In_160);
or U161 (N_161,In_51,In_107);
nor U162 (N_162,In_458,In_35);
nand U163 (N_163,In_445,In_438);
and U164 (N_164,In_104,In_485);
nand U165 (N_165,In_355,In_3);
nor U166 (N_166,In_58,In_22);
and U167 (N_167,In_317,In_431);
and U168 (N_168,In_415,In_75);
and U169 (N_169,In_207,In_436);
nand U170 (N_170,In_142,In_168);
nand U171 (N_171,In_59,In_274);
and U172 (N_172,In_197,In_359);
and U173 (N_173,In_296,In_173);
and U174 (N_174,In_20,In_304);
nand U175 (N_175,In_129,In_76);
or U176 (N_176,In_305,In_302);
and U177 (N_177,In_87,In_316);
nand U178 (N_178,In_86,In_349);
or U179 (N_179,In_399,In_134);
or U180 (N_180,In_472,In_108);
and U181 (N_181,In_224,In_333);
or U182 (N_182,In_8,In_339);
xor U183 (N_183,In_480,In_430);
nor U184 (N_184,In_190,In_371);
and U185 (N_185,In_188,In_186);
or U186 (N_186,In_307,In_37);
or U187 (N_187,In_443,In_57);
and U188 (N_188,In_211,In_32);
and U189 (N_189,In_65,In_177);
nor U190 (N_190,In_56,In_424);
and U191 (N_191,In_336,In_392);
nor U192 (N_192,In_344,In_318);
nand U193 (N_193,In_352,In_368);
or U194 (N_194,In_487,In_239);
and U195 (N_195,In_216,In_13);
and U196 (N_196,In_234,In_84);
or U197 (N_197,In_40,In_219);
or U198 (N_198,In_258,In_77);
or U199 (N_199,In_427,In_466);
and U200 (N_200,In_373,In_340);
or U201 (N_201,In_116,In_268);
nand U202 (N_202,In_184,In_261);
nand U203 (N_203,In_73,In_247);
nor U204 (N_204,In_89,In_226);
nor U205 (N_205,In_4,In_21);
and U206 (N_206,In_112,In_136);
xnor U207 (N_207,In_218,In_185);
nand U208 (N_208,In_52,In_408);
nand U209 (N_209,In_370,In_380);
nand U210 (N_210,In_194,In_223);
or U211 (N_211,In_175,In_439);
and U212 (N_212,In_115,In_255);
and U213 (N_213,In_178,In_203);
nand U214 (N_214,In_422,In_231);
nor U215 (N_215,In_262,In_366);
nor U216 (N_216,In_383,In_332);
or U217 (N_217,In_381,In_358);
nor U218 (N_218,In_170,In_270);
nor U219 (N_219,In_69,In_127);
nand U220 (N_220,In_283,In_235);
and U221 (N_221,In_497,In_41);
nor U222 (N_222,In_496,In_287);
xor U223 (N_223,In_319,In_471);
and U224 (N_224,In_393,In_180);
nand U225 (N_225,In_97,In_187);
and U226 (N_226,In_195,In_285);
and U227 (N_227,In_43,In_354);
nor U228 (N_228,In_309,In_396);
xor U229 (N_229,In_105,In_245);
and U230 (N_230,In_375,In_38);
and U231 (N_231,In_457,In_331);
nor U232 (N_232,In_374,In_495);
nor U233 (N_233,In_212,In_464);
or U234 (N_234,In_446,In_242);
or U235 (N_235,In_327,In_303);
and U236 (N_236,In_478,In_310);
nand U237 (N_237,In_111,In_225);
or U238 (N_238,In_461,In_46);
or U239 (N_239,In_260,In_62);
xnor U240 (N_240,In_403,In_48);
and U241 (N_241,In_34,In_397);
nor U242 (N_242,In_240,In_361);
or U243 (N_243,In_148,In_460);
nor U244 (N_244,In_171,In_27);
xnor U245 (N_245,In_228,In_91);
nor U246 (N_246,In_314,In_210);
or U247 (N_247,In_167,In_386);
xnor U248 (N_248,In_362,In_377);
nand U249 (N_249,In_179,In_63);
xor U250 (N_250,In_242,In_147);
nand U251 (N_251,In_172,In_387);
nor U252 (N_252,In_457,In_468);
xor U253 (N_253,In_420,In_314);
xnor U254 (N_254,In_426,In_292);
nand U255 (N_255,In_194,In_408);
or U256 (N_256,In_167,In_0);
or U257 (N_257,In_244,In_325);
nor U258 (N_258,In_84,In_82);
and U259 (N_259,In_350,In_31);
and U260 (N_260,In_435,In_194);
nand U261 (N_261,In_467,In_226);
nand U262 (N_262,In_491,In_304);
and U263 (N_263,In_434,In_464);
nor U264 (N_264,In_248,In_387);
nand U265 (N_265,In_456,In_81);
or U266 (N_266,In_282,In_351);
xnor U267 (N_267,In_208,In_179);
or U268 (N_268,In_303,In_407);
nand U269 (N_269,In_86,In_60);
or U270 (N_270,In_176,In_149);
and U271 (N_271,In_355,In_374);
nor U272 (N_272,In_161,In_140);
and U273 (N_273,In_276,In_34);
or U274 (N_274,In_139,In_8);
nor U275 (N_275,In_44,In_444);
xnor U276 (N_276,In_289,In_57);
xor U277 (N_277,In_185,In_478);
or U278 (N_278,In_119,In_388);
nand U279 (N_279,In_2,In_450);
and U280 (N_280,In_148,In_18);
or U281 (N_281,In_77,In_61);
nor U282 (N_282,In_154,In_50);
xor U283 (N_283,In_429,In_171);
and U284 (N_284,In_342,In_355);
nor U285 (N_285,In_304,In_471);
nor U286 (N_286,In_33,In_147);
or U287 (N_287,In_232,In_360);
nand U288 (N_288,In_102,In_106);
nand U289 (N_289,In_370,In_15);
nand U290 (N_290,In_108,In_241);
nor U291 (N_291,In_195,In_249);
nand U292 (N_292,In_61,In_419);
nor U293 (N_293,In_331,In_214);
and U294 (N_294,In_432,In_409);
nor U295 (N_295,In_124,In_344);
nor U296 (N_296,In_473,In_207);
nor U297 (N_297,In_139,In_216);
nand U298 (N_298,In_282,In_85);
nor U299 (N_299,In_106,In_225);
xnor U300 (N_300,In_87,In_453);
and U301 (N_301,In_292,In_73);
nand U302 (N_302,In_161,In_481);
or U303 (N_303,In_339,In_372);
nor U304 (N_304,In_280,In_184);
xnor U305 (N_305,In_169,In_64);
xor U306 (N_306,In_489,In_55);
or U307 (N_307,In_126,In_187);
nand U308 (N_308,In_2,In_479);
nand U309 (N_309,In_47,In_323);
or U310 (N_310,In_375,In_31);
and U311 (N_311,In_48,In_36);
and U312 (N_312,In_227,In_191);
and U313 (N_313,In_335,In_343);
nand U314 (N_314,In_201,In_364);
nor U315 (N_315,In_278,In_257);
nand U316 (N_316,In_351,In_460);
nand U317 (N_317,In_29,In_116);
and U318 (N_318,In_290,In_48);
nor U319 (N_319,In_3,In_141);
or U320 (N_320,In_397,In_453);
xor U321 (N_321,In_45,In_179);
nand U322 (N_322,In_474,In_96);
and U323 (N_323,In_141,In_454);
nand U324 (N_324,In_389,In_33);
or U325 (N_325,In_27,In_394);
xor U326 (N_326,In_359,In_130);
and U327 (N_327,In_146,In_325);
or U328 (N_328,In_297,In_25);
nor U329 (N_329,In_376,In_235);
nand U330 (N_330,In_98,In_187);
nor U331 (N_331,In_342,In_379);
and U332 (N_332,In_164,In_248);
and U333 (N_333,In_78,In_192);
nor U334 (N_334,In_271,In_80);
or U335 (N_335,In_229,In_0);
and U336 (N_336,In_175,In_133);
nor U337 (N_337,In_35,In_273);
and U338 (N_338,In_274,In_71);
xnor U339 (N_339,In_284,In_66);
or U340 (N_340,In_238,In_253);
nor U341 (N_341,In_317,In_90);
or U342 (N_342,In_161,In_203);
xnor U343 (N_343,In_192,In_209);
nand U344 (N_344,In_358,In_64);
and U345 (N_345,In_235,In_17);
xnor U346 (N_346,In_293,In_280);
or U347 (N_347,In_398,In_179);
or U348 (N_348,In_143,In_458);
nand U349 (N_349,In_54,In_267);
and U350 (N_350,In_303,In_253);
nand U351 (N_351,In_103,In_275);
nor U352 (N_352,In_23,In_292);
and U353 (N_353,In_22,In_186);
nor U354 (N_354,In_286,In_81);
nor U355 (N_355,In_443,In_90);
and U356 (N_356,In_239,In_328);
nand U357 (N_357,In_469,In_87);
nor U358 (N_358,In_303,In_138);
nor U359 (N_359,In_377,In_40);
xor U360 (N_360,In_449,In_408);
or U361 (N_361,In_438,In_286);
xor U362 (N_362,In_29,In_133);
nor U363 (N_363,In_283,In_0);
nand U364 (N_364,In_449,In_265);
nand U365 (N_365,In_247,In_128);
nor U366 (N_366,In_96,In_455);
xor U367 (N_367,In_298,In_435);
and U368 (N_368,In_148,In_319);
nand U369 (N_369,In_39,In_122);
nand U370 (N_370,In_7,In_155);
and U371 (N_371,In_494,In_226);
nand U372 (N_372,In_24,In_213);
nand U373 (N_373,In_123,In_441);
or U374 (N_374,In_475,In_499);
and U375 (N_375,In_230,In_10);
or U376 (N_376,In_372,In_454);
or U377 (N_377,In_250,In_349);
and U378 (N_378,In_268,In_186);
or U379 (N_379,In_268,In_99);
nor U380 (N_380,In_227,In_499);
and U381 (N_381,In_158,In_15);
nor U382 (N_382,In_242,In_442);
and U383 (N_383,In_67,In_337);
or U384 (N_384,In_337,In_377);
and U385 (N_385,In_265,In_142);
or U386 (N_386,In_365,In_85);
and U387 (N_387,In_407,In_296);
nor U388 (N_388,In_452,In_307);
or U389 (N_389,In_88,In_4);
or U390 (N_390,In_129,In_224);
or U391 (N_391,In_434,In_373);
and U392 (N_392,In_365,In_82);
nand U393 (N_393,In_77,In_33);
nand U394 (N_394,In_333,In_221);
or U395 (N_395,In_9,In_272);
nor U396 (N_396,In_125,In_97);
nor U397 (N_397,In_118,In_421);
and U398 (N_398,In_247,In_235);
and U399 (N_399,In_55,In_385);
nand U400 (N_400,In_243,In_332);
and U401 (N_401,In_378,In_231);
and U402 (N_402,In_334,In_204);
nand U403 (N_403,In_259,In_429);
xor U404 (N_404,In_440,In_338);
nor U405 (N_405,In_292,In_191);
nand U406 (N_406,In_259,In_403);
xnor U407 (N_407,In_191,In_472);
or U408 (N_408,In_75,In_209);
nor U409 (N_409,In_81,In_472);
and U410 (N_410,In_414,In_189);
and U411 (N_411,In_103,In_464);
nor U412 (N_412,In_365,In_368);
and U413 (N_413,In_299,In_124);
or U414 (N_414,In_129,In_174);
nand U415 (N_415,In_405,In_139);
nand U416 (N_416,In_468,In_103);
and U417 (N_417,In_219,In_127);
nand U418 (N_418,In_174,In_197);
and U419 (N_419,In_197,In_441);
and U420 (N_420,In_211,In_158);
or U421 (N_421,In_286,In_423);
or U422 (N_422,In_361,In_192);
or U423 (N_423,In_269,In_299);
and U424 (N_424,In_412,In_494);
or U425 (N_425,In_118,In_194);
nand U426 (N_426,In_446,In_161);
nor U427 (N_427,In_144,In_351);
nand U428 (N_428,In_366,In_329);
nor U429 (N_429,In_443,In_330);
and U430 (N_430,In_359,In_261);
or U431 (N_431,In_24,In_124);
nand U432 (N_432,In_176,In_419);
xnor U433 (N_433,In_338,In_41);
nand U434 (N_434,In_237,In_225);
nor U435 (N_435,In_238,In_442);
nor U436 (N_436,In_172,In_65);
nor U437 (N_437,In_242,In_218);
nor U438 (N_438,In_290,In_221);
nand U439 (N_439,In_97,In_336);
or U440 (N_440,In_29,In_432);
xor U441 (N_441,In_47,In_372);
nand U442 (N_442,In_97,In_5);
nor U443 (N_443,In_279,In_104);
and U444 (N_444,In_167,In_102);
or U445 (N_445,In_45,In_173);
nand U446 (N_446,In_427,In_149);
or U447 (N_447,In_179,In_204);
or U448 (N_448,In_153,In_131);
nor U449 (N_449,In_315,In_79);
nor U450 (N_450,In_399,In_33);
nor U451 (N_451,In_236,In_244);
nand U452 (N_452,In_232,In_363);
and U453 (N_453,In_298,In_470);
and U454 (N_454,In_178,In_372);
and U455 (N_455,In_279,In_466);
and U456 (N_456,In_361,In_52);
and U457 (N_457,In_32,In_93);
xor U458 (N_458,In_138,In_186);
nand U459 (N_459,In_225,In_468);
nor U460 (N_460,In_166,In_241);
or U461 (N_461,In_56,In_111);
and U462 (N_462,In_359,In_26);
nand U463 (N_463,In_489,In_140);
nor U464 (N_464,In_354,In_246);
xnor U465 (N_465,In_495,In_175);
nor U466 (N_466,In_449,In_16);
nor U467 (N_467,In_398,In_118);
nor U468 (N_468,In_112,In_407);
or U469 (N_469,In_241,In_438);
nand U470 (N_470,In_45,In_459);
nor U471 (N_471,In_264,In_307);
or U472 (N_472,In_248,In_299);
nand U473 (N_473,In_195,In_409);
nor U474 (N_474,In_370,In_240);
nand U475 (N_475,In_53,In_410);
nor U476 (N_476,In_227,In_307);
xor U477 (N_477,In_263,In_267);
and U478 (N_478,In_144,In_97);
nor U479 (N_479,In_241,In_332);
or U480 (N_480,In_323,In_409);
or U481 (N_481,In_471,In_386);
nand U482 (N_482,In_404,In_44);
or U483 (N_483,In_77,In_215);
nand U484 (N_484,In_41,In_408);
and U485 (N_485,In_443,In_388);
or U486 (N_486,In_107,In_156);
and U487 (N_487,In_495,In_286);
nand U488 (N_488,In_253,In_342);
and U489 (N_489,In_425,In_462);
nor U490 (N_490,In_345,In_361);
or U491 (N_491,In_121,In_327);
and U492 (N_492,In_17,In_122);
nor U493 (N_493,In_371,In_0);
nor U494 (N_494,In_82,In_208);
nor U495 (N_495,In_31,In_50);
xor U496 (N_496,In_303,In_100);
nor U497 (N_497,In_111,In_459);
and U498 (N_498,In_387,In_30);
nand U499 (N_499,In_465,In_171);
and U500 (N_500,N_481,N_193);
and U501 (N_501,N_216,N_188);
or U502 (N_502,N_292,N_486);
or U503 (N_503,N_124,N_43);
or U504 (N_504,N_280,N_147);
or U505 (N_505,N_51,N_376);
or U506 (N_506,N_152,N_319);
or U507 (N_507,N_108,N_338);
xnor U508 (N_508,N_359,N_125);
and U509 (N_509,N_207,N_453);
or U510 (N_510,N_466,N_160);
nand U511 (N_511,N_121,N_276);
or U512 (N_512,N_383,N_80);
or U513 (N_513,N_149,N_7);
nand U514 (N_514,N_205,N_26);
and U515 (N_515,N_213,N_409);
and U516 (N_516,N_123,N_284);
and U517 (N_517,N_454,N_435);
and U518 (N_518,N_267,N_187);
and U519 (N_519,N_106,N_170);
and U520 (N_520,N_459,N_233);
nor U521 (N_521,N_257,N_477);
or U522 (N_522,N_374,N_394);
or U523 (N_523,N_371,N_138);
or U524 (N_524,N_350,N_455);
nor U525 (N_525,N_315,N_365);
and U526 (N_526,N_9,N_151);
nand U527 (N_527,N_402,N_73);
or U528 (N_528,N_8,N_64);
and U529 (N_529,N_404,N_272);
xnor U530 (N_530,N_490,N_169);
or U531 (N_531,N_268,N_426);
xor U532 (N_532,N_97,N_388);
nand U533 (N_533,N_443,N_334);
or U534 (N_534,N_136,N_153);
and U535 (N_535,N_59,N_61);
nand U536 (N_536,N_133,N_57);
nand U537 (N_537,N_415,N_56);
or U538 (N_538,N_194,N_69);
nand U539 (N_539,N_163,N_174);
or U540 (N_540,N_273,N_444);
nor U541 (N_541,N_183,N_295);
nand U542 (N_542,N_68,N_297);
nand U543 (N_543,N_15,N_29);
and U544 (N_544,N_399,N_261);
nand U545 (N_545,N_231,N_202);
and U546 (N_546,N_175,N_158);
nor U547 (N_547,N_236,N_333);
nor U548 (N_548,N_422,N_178);
nor U549 (N_549,N_11,N_200);
nand U550 (N_550,N_498,N_52);
or U551 (N_551,N_14,N_358);
nand U552 (N_552,N_439,N_421);
xor U553 (N_553,N_162,N_309);
or U554 (N_554,N_21,N_89);
nand U555 (N_555,N_234,N_214);
nor U556 (N_556,N_90,N_131);
nor U557 (N_557,N_62,N_127);
or U558 (N_558,N_237,N_351);
and U559 (N_559,N_128,N_396);
nand U560 (N_560,N_217,N_122);
or U561 (N_561,N_173,N_400);
or U562 (N_562,N_203,N_497);
and U563 (N_563,N_141,N_375);
or U564 (N_564,N_253,N_289);
nand U565 (N_565,N_5,N_177);
nor U566 (N_566,N_274,N_419);
nand U567 (N_567,N_196,N_380);
nand U568 (N_568,N_204,N_304);
and U569 (N_569,N_485,N_215);
or U570 (N_570,N_85,N_356);
xor U571 (N_571,N_135,N_168);
or U572 (N_572,N_101,N_457);
nand U573 (N_573,N_437,N_346);
and U574 (N_574,N_30,N_58);
nor U575 (N_575,N_171,N_357);
or U576 (N_576,N_305,N_251);
xnor U577 (N_577,N_16,N_464);
or U578 (N_578,N_260,N_201);
nand U579 (N_579,N_82,N_499);
or U580 (N_580,N_329,N_195);
or U581 (N_581,N_244,N_35);
or U582 (N_582,N_287,N_102);
or U583 (N_583,N_142,N_219);
nor U584 (N_584,N_489,N_316);
or U585 (N_585,N_28,N_386);
and U586 (N_586,N_473,N_296);
nand U587 (N_587,N_487,N_472);
xnor U588 (N_588,N_463,N_208);
or U589 (N_589,N_34,N_46);
or U590 (N_590,N_243,N_345);
nand U591 (N_591,N_0,N_112);
nor U592 (N_592,N_335,N_32);
or U593 (N_593,N_339,N_103);
and U594 (N_594,N_199,N_181);
and U595 (N_595,N_120,N_172);
xnor U596 (N_596,N_155,N_495);
nand U597 (N_597,N_38,N_478);
and U598 (N_598,N_407,N_191);
nor U599 (N_599,N_84,N_33);
and U600 (N_600,N_352,N_382);
nand U601 (N_601,N_332,N_161);
nand U602 (N_602,N_54,N_156);
nand U603 (N_603,N_37,N_465);
xnor U604 (N_604,N_265,N_442);
xnor U605 (N_605,N_456,N_27);
nor U606 (N_606,N_362,N_418);
nor U607 (N_607,N_104,N_23);
and U608 (N_608,N_119,N_398);
nor U609 (N_609,N_303,N_293);
xnor U610 (N_610,N_431,N_475);
nand U611 (N_611,N_238,N_269);
and U612 (N_612,N_159,N_72);
xnor U613 (N_613,N_401,N_474);
nor U614 (N_614,N_348,N_414);
and U615 (N_615,N_307,N_197);
or U616 (N_616,N_99,N_228);
and U617 (N_617,N_255,N_258);
nand U618 (N_618,N_143,N_450);
nand U619 (N_619,N_259,N_392);
or U620 (N_620,N_283,N_310);
nand U621 (N_621,N_93,N_134);
xnor U622 (N_622,N_91,N_471);
nor U623 (N_623,N_210,N_406);
or U624 (N_624,N_446,N_167);
or U625 (N_625,N_55,N_118);
nor U626 (N_626,N_291,N_330);
and U627 (N_627,N_311,N_229);
xnor U628 (N_628,N_343,N_360);
or U629 (N_629,N_427,N_189);
nor U630 (N_630,N_412,N_440);
and U631 (N_631,N_278,N_98);
nor U632 (N_632,N_479,N_71);
and U633 (N_633,N_100,N_462);
nand U634 (N_634,N_45,N_209);
or U635 (N_635,N_340,N_96);
nor U636 (N_636,N_239,N_468);
or U637 (N_637,N_266,N_429);
nor U638 (N_638,N_282,N_331);
and U639 (N_639,N_230,N_77);
nand U640 (N_640,N_290,N_405);
or U641 (N_641,N_366,N_279);
nand U642 (N_642,N_18,N_250);
or U643 (N_643,N_460,N_328);
and U644 (N_644,N_241,N_146);
nand U645 (N_645,N_19,N_86);
nand U646 (N_646,N_354,N_300);
xor U647 (N_647,N_67,N_433);
nor U648 (N_648,N_342,N_49);
and U649 (N_649,N_185,N_313);
or U650 (N_650,N_70,N_115);
nor U651 (N_651,N_299,N_370);
nand U652 (N_652,N_94,N_325);
and U653 (N_653,N_111,N_379);
and U654 (N_654,N_397,N_150);
nor U655 (N_655,N_186,N_470);
and U656 (N_656,N_347,N_182);
nand U657 (N_657,N_166,N_434);
nand U658 (N_658,N_324,N_116);
nand U659 (N_659,N_137,N_17);
xnor U660 (N_660,N_192,N_249);
and U661 (N_661,N_294,N_107);
and U662 (N_662,N_66,N_323);
xor U663 (N_663,N_242,N_246);
or U664 (N_664,N_417,N_109);
nand U665 (N_665,N_469,N_372);
xnor U666 (N_666,N_132,N_312);
and U667 (N_667,N_441,N_391);
and U668 (N_668,N_78,N_224);
nor U669 (N_669,N_20,N_467);
or U670 (N_670,N_378,N_320);
and U671 (N_671,N_218,N_165);
xnor U672 (N_672,N_13,N_321);
nand U673 (N_673,N_390,N_318);
or U674 (N_674,N_263,N_286);
and U675 (N_675,N_48,N_252);
nand U676 (N_676,N_484,N_423);
nor U677 (N_677,N_75,N_126);
nand U678 (N_678,N_113,N_3);
nor U679 (N_679,N_271,N_39);
nor U680 (N_680,N_413,N_377);
or U681 (N_681,N_449,N_416);
nor U682 (N_682,N_164,N_395);
and U683 (N_683,N_81,N_226);
nor U684 (N_684,N_47,N_428);
or U685 (N_685,N_410,N_384);
nand U686 (N_686,N_227,N_448);
nor U687 (N_687,N_387,N_1);
and U688 (N_688,N_31,N_425);
or U689 (N_689,N_198,N_496);
and U690 (N_690,N_190,N_306);
and U691 (N_691,N_301,N_245);
nor U692 (N_692,N_24,N_341);
nor U693 (N_693,N_285,N_317);
and U694 (N_694,N_447,N_211);
and U695 (N_695,N_420,N_83);
or U696 (N_696,N_248,N_50);
nor U697 (N_697,N_275,N_40);
and U698 (N_698,N_270,N_247);
or U699 (N_699,N_88,N_436);
and U700 (N_700,N_117,N_353);
or U701 (N_701,N_488,N_432);
or U702 (N_702,N_87,N_438);
or U703 (N_703,N_95,N_368);
xnor U704 (N_704,N_389,N_74);
and U705 (N_705,N_298,N_483);
nor U706 (N_706,N_129,N_491);
nor U707 (N_707,N_349,N_385);
or U708 (N_708,N_277,N_308);
or U709 (N_709,N_336,N_355);
and U710 (N_710,N_10,N_110);
nand U711 (N_711,N_105,N_184);
nor U712 (N_712,N_452,N_139);
or U713 (N_713,N_369,N_256);
nor U714 (N_714,N_140,N_367);
nand U715 (N_715,N_322,N_212);
or U716 (N_716,N_65,N_53);
or U717 (N_717,N_25,N_424);
and U718 (N_718,N_36,N_206);
nand U719 (N_719,N_364,N_180);
nor U720 (N_720,N_6,N_492);
and U721 (N_721,N_326,N_281);
nor U722 (N_722,N_222,N_344);
nor U723 (N_723,N_148,N_114);
or U724 (N_724,N_176,N_411);
and U725 (N_725,N_327,N_408);
or U726 (N_726,N_363,N_157);
nand U727 (N_727,N_76,N_144);
or U728 (N_728,N_4,N_240);
nor U729 (N_729,N_92,N_232);
nor U730 (N_730,N_373,N_288);
nand U731 (N_731,N_381,N_337);
or U732 (N_732,N_41,N_476);
or U733 (N_733,N_42,N_430);
nand U734 (N_734,N_393,N_179);
and U735 (N_735,N_145,N_79);
and U736 (N_736,N_254,N_154);
and U737 (N_737,N_223,N_130);
and U738 (N_738,N_2,N_314);
nand U739 (N_739,N_451,N_480);
nand U740 (N_740,N_44,N_445);
nor U741 (N_741,N_302,N_225);
or U742 (N_742,N_22,N_60);
nor U743 (N_743,N_63,N_220);
or U744 (N_744,N_235,N_403);
xnor U745 (N_745,N_221,N_461);
xor U746 (N_746,N_12,N_493);
or U747 (N_747,N_361,N_494);
or U748 (N_748,N_482,N_458);
nand U749 (N_749,N_262,N_264);
or U750 (N_750,N_144,N_116);
xor U751 (N_751,N_120,N_371);
nor U752 (N_752,N_208,N_333);
or U753 (N_753,N_235,N_379);
or U754 (N_754,N_395,N_148);
and U755 (N_755,N_60,N_95);
or U756 (N_756,N_160,N_388);
nand U757 (N_757,N_86,N_187);
or U758 (N_758,N_148,N_152);
nor U759 (N_759,N_328,N_172);
nor U760 (N_760,N_4,N_214);
or U761 (N_761,N_98,N_86);
and U762 (N_762,N_148,N_105);
nand U763 (N_763,N_85,N_163);
nand U764 (N_764,N_179,N_18);
nor U765 (N_765,N_156,N_439);
xnor U766 (N_766,N_247,N_314);
or U767 (N_767,N_435,N_407);
or U768 (N_768,N_74,N_123);
xnor U769 (N_769,N_214,N_199);
or U770 (N_770,N_368,N_231);
nand U771 (N_771,N_92,N_58);
nor U772 (N_772,N_367,N_283);
or U773 (N_773,N_352,N_239);
nor U774 (N_774,N_60,N_308);
nand U775 (N_775,N_368,N_136);
and U776 (N_776,N_422,N_433);
nor U777 (N_777,N_221,N_38);
nand U778 (N_778,N_210,N_9);
nand U779 (N_779,N_259,N_174);
and U780 (N_780,N_397,N_342);
and U781 (N_781,N_333,N_101);
nor U782 (N_782,N_222,N_346);
or U783 (N_783,N_211,N_289);
nand U784 (N_784,N_348,N_89);
and U785 (N_785,N_255,N_123);
xor U786 (N_786,N_352,N_363);
nand U787 (N_787,N_447,N_344);
xor U788 (N_788,N_219,N_20);
and U789 (N_789,N_39,N_399);
nor U790 (N_790,N_147,N_168);
nand U791 (N_791,N_372,N_347);
nand U792 (N_792,N_316,N_71);
nor U793 (N_793,N_181,N_50);
xor U794 (N_794,N_373,N_63);
xnor U795 (N_795,N_317,N_406);
or U796 (N_796,N_44,N_38);
nor U797 (N_797,N_100,N_27);
nand U798 (N_798,N_426,N_208);
xor U799 (N_799,N_234,N_223);
and U800 (N_800,N_497,N_242);
and U801 (N_801,N_203,N_335);
and U802 (N_802,N_165,N_243);
and U803 (N_803,N_80,N_329);
and U804 (N_804,N_100,N_225);
and U805 (N_805,N_279,N_344);
nor U806 (N_806,N_216,N_25);
or U807 (N_807,N_400,N_221);
and U808 (N_808,N_69,N_13);
nor U809 (N_809,N_146,N_374);
nand U810 (N_810,N_312,N_196);
nor U811 (N_811,N_164,N_329);
nor U812 (N_812,N_180,N_281);
nor U813 (N_813,N_352,N_2);
nand U814 (N_814,N_47,N_349);
and U815 (N_815,N_15,N_167);
or U816 (N_816,N_2,N_471);
nor U817 (N_817,N_338,N_254);
or U818 (N_818,N_126,N_434);
nand U819 (N_819,N_454,N_448);
nand U820 (N_820,N_79,N_443);
or U821 (N_821,N_145,N_326);
nor U822 (N_822,N_153,N_11);
nand U823 (N_823,N_164,N_435);
or U824 (N_824,N_233,N_169);
and U825 (N_825,N_240,N_117);
and U826 (N_826,N_440,N_365);
nand U827 (N_827,N_416,N_46);
nand U828 (N_828,N_8,N_348);
nand U829 (N_829,N_230,N_487);
xnor U830 (N_830,N_229,N_437);
and U831 (N_831,N_423,N_264);
and U832 (N_832,N_320,N_245);
and U833 (N_833,N_388,N_61);
nor U834 (N_834,N_205,N_487);
or U835 (N_835,N_263,N_465);
and U836 (N_836,N_135,N_419);
nand U837 (N_837,N_345,N_408);
nand U838 (N_838,N_416,N_209);
nand U839 (N_839,N_480,N_210);
and U840 (N_840,N_378,N_51);
nor U841 (N_841,N_159,N_100);
or U842 (N_842,N_114,N_431);
and U843 (N_843,N_130,N_261);
or U844 (N_844,N_421,N_176);
nand U845 (N_845,N_97,N_233);
or U846 (N_846,N_122,N_328);
nor U847 (N_847,N_105,N_114);
nor U848 (N_848,N_273,N_457);
or U849 (N_849,N_140,N_416);
and U850 (N_850,N_409,N_336);
xnor U851 (N_851,N_172,N_460);
nand U852 (N_852,N_94,N_480);
nand U853 (N_853,N_321,N_252);
nand U854 (N_854,N_330,N_108);
nand U855 (N_855,N_17,N_124);
nand U856 (N_856,N_288,N_446);
or U857 (N_857,N_14,N_220);
nor U858 (N_858,N_146,N_292);
or U859 (N_859,N_47,N_294);
nand U860 (N_860,N_471,N_71);
nor U861 (N_861,N_104,N_20);
and U862 (N_862,N_327,N_145);
and U863 (N_863,N_447,N_147);
or U864 (N_864,N_289,N_305);
nor U865 (N_865,N_342,N_439);
or U866 (N_866,N_60,N_418);
or U867 (N_867,N_461,N_7);
and U868 (N_868,N_340,N_493);
or U869 (N_869,N_58,N_36);
and U870 (N_870,N_454,N_201);
nor U871 (N_871,N_349,N_343);
and U872 (N_872,N_263,N_225);
nor U873 (N_873,N_296,N_90);
nand U874 (N_874,N_140,N_214);
or U875 (N_875,N_310,N_301);
or U876 (N_876,N_428,N_491);
nand U877 (N_877,N_92,N_469);
or U878 (N_878,N_355,N_431);
or U879 (N_879,N_137,N_479);
nand U880 (N_880,N_192,N_402);
nor U881 (N_881,N_184,N_160);
or U882 (N_882,N_151,N_95);
and U883 (N_883,N_494,N_245);
or U884 (N_884,N_2,N_419);
or U885 (N_885,N_137,N_101);
nor U886 (N_886,N_173,N_42);
nand U887 (N_887,N_257,N_130);
and U888 (N_888,N_90,N_8);
or U889 (N_889,N_278,N_211);
nor U890 (N_890,N_457,N_94);
or U891 (N_891,N_188,N_198);
or U892 (N_892,N_411,N_31);
and U893 (N_893,N_304,N_360);
and U894 (N_894,N_11,N_174);
nor U895 (N_895,N_187,N_274);
nor U896 (N_896,N_220,N_387);
and U897 (N_897,N_133,N_69);
and U898 (N_898,N_117,N_415);
and U899 (N_899,N_262,N_495);
and U900 (N_900,N_369,N_462);
and U901 (N_901,N_436,N_146);
nand U902 (N_902,N_391,N_236);
or U903 (N_903,N_89,N_6);
xnor U904 (N_904,N_307,N_444);
nor U905 (N_905,N_178,N_158);
nand U906 (N_906,N_259,N_40);
or U907 (N_907,N_292,N_192);
or U908 (N_908,N_200,N_417);
nor U909 (N_909,N_498,N_25);
or U910 (N_910,N_361,N_76);
or U911 (N_911,N_496,N_86);
or U912 (N_912,N_163,N_186);
and U913 (N_913,N_292,N_356);
or U914 (N_914,N_238,N_198);
or U915 (N_915,N_341,N_485);
nor U916 (N_916,N_134,N_2);
and U917 (N_917,N_47,N_434);
and U918 (N_918,N_203,N_337);
or U919 (N_919,N_68,N_186);
nand U920 (N_920,N_388,N_253);
or U921 (N_921,N_228,N_283);
and U922 (N_922,N_97,N_121);
or U923 (N_923,N_43,N_442);
nand U924 (N_924,N_0,N_2);
nor U925 (N_925,N_41,N_356);
and U926 (N_926,N_112,N_422);
and U927 (N_927,N_206,N_228);
and U928 (N_928,N_109,N_384);
xor U929 (N_929,N_7,N_470);
nand U930 (N_930,N_425,N_201);
xor U931 (N_931,N_76,N_64);
xnor U932 (N_932,N_282,N_426);
nand U933 (N_933,N_303,N_208);
or U934 (N_934,N_100,N_24);
nor U935 (N_935,N_242,N_12);
and U936 (N_936,N_42,N_119);
nor U937 (N_937,N_22,N_375);
xor U938 (N_938,N_96,N_138);
and U939 (N_939,N_96,N_487);
nor U940 (N_940,N_381,N_435);
nor U941 (N_941,N_41,N_71);
nor U942 (N_942,N_153,N_276);
nor U943 (N_943,N_462,N_85);
nand U944 (N_944,N_244,N_395);
nand U945 (N_945,N_124,N_116);
and U946 (N_946,N_368,N_477);
nor U947 (N_947,N_363,N_268);
nor U948 (N_948,N_331,N_475);
or U949 (N_949,N_314,N_21);
xnor U950 (N_950,N_179,N_306);
and U951 (N_951,N_111,N_76);
nand U952 (N_952,N_337,N_407);
nor U953 (N_953,N_373,N_377);
nand U954 (N_954,N_1,N_435);
xnor U955 (N_955,N_337,N_453);
or U956 (N_956,N_28,N_282);
nand U957 (N_957,N_34,N_63);
nor U958 (N_958,N_225,N_156);
or U959 (N_959,N_120,N_464);
nand U960 (N_960,N_375,N_63);
and U961 (N_961,N_384,N_22);
and U962 (N_962,N_287,N_406);
or U963 (N_963,N_273,N_140);
nor U964 (N_964,N_168,N_21);
and U965 (N_965,N_409,N_291);
nand U966 (N_966,N_37,N_395);
xor U967 (N_967,N_321,N_134);
nor U968 (N_968,N_401,N_181);
nor U969 (N_969,N_29,N_459);
or U970 (N_970,N_11,N_344);
nor U971 (N_971,N_137,N_455);
nor U972 (N_972,N_458,N_470);
nor U973 (N_973,N_115,N_89);
or U974 (N_974,N_460,N_482);
nand U975 (N_975,N_263,N_145);
or U976 (N_976,N_64,N_73);
nand U977 (N_977,N_344,N_388);
nor U978 (N_978,N_89,N_192);
and U979 (N_979,N_200,N_415);
and U980 (N_980,N_106,N_30);
or U981 (N_981,N_433,N_112);
nand U982 (N_982,N_196,N_348);
nor U983 (N_983,N_281,N_450);
nand U984 (N_984,N_213,N_128);
nand U985 (N_985,N_394,N_275);
nand U986 (N_986,N_260,N_29);
or U987 (N_987,N_99,N_420);
nand U988 (N_988,N_485,N_34);
and U989 (N_989,N_497,N_491);
and U990 (N_990,N_41,N_9);
nor U991 (N_991,N_329,N_78);
and U992 (N_992,N_447,N_74);
nor U993 (N_993,N_166,N_488);
or U994 (N_994,N_415,N_261);
nand U995 (N_995,N_15,N_225);
or U996 (N_996,N_65,N_187);
and U997 (N_997,N_25,N_436);
or U998 (N_998,N_349,N_369);
xnor U999 (N_999,N_104,N_446);
nor U1000 (N_1000,N_531,N_884);
nand U1001 (N_1001,N_858,N_551);
xnor U1002 (N_1002,N_801,N_800);
nor U1003 (N_1003,N_512,N_698);
or U1004 (N_1004,N_802,N_608);
nand U1005 (N_1005,N_534,N_899);
xor U1006 (N_1006,N_723,N_612);
xnor U1007 (N_1007,N_553,N_909);
nand U1008 (N_1008,N_713,N_677);
and U1009 (N_1009,N_572,N_836);
or U1010 (N_1010,N_936,N_826);
xnor U1011 (N_1011,N_813,N_564);
or U1012 (N_1012,N_992,N_834);
nand U1013 (N_1013,N_778,N_971);
and U1014 (N_1014,N_558,N_573);
xor U1015 (N_1015,N_975,N_959);
and U1016 (N_1016,N_565,N_591);
nand U1017 (N_1017,N_883,N_650);
nor U1018 (N_1018,N_900,N_871);
and U1019 (N_1019,N_961,N_576);
and U1020 (N_1020,N_599,N_841);
nor U1021 (N_1021,N_995,N_970);
or U1022 (N_1022,N_745,N_821);
and U1023 (N_1023,N_810,N_803);
or U1024 (N_1024,N_860,N_822);
nor U1025 (N_1025,N_525,N_504);
nor U1026 (N_1026,N_919,N_736);
and U1027 (N_1027,N_503,N_615);
xor U1028 (N_1028,N_830,N_845);
xnor U1029 (N_1029,N_928,N_777);
xor U1030 (N_1030,N_976,N_655);
or U1031 (N_1031,N_501,N_543);
xnor U1032 (N_1032,N_942,N_738);
nor U1033 (N_1033,N_637,N_704);
nand U1034 (N_1034,N_596,N_526);
and U1035 (N_1035,N_540,N_852);
nand U1036 (N_1036,N_545,N_740);
or U1037 (N_1037,N_958,N_869);
and U1038 (N_1038,N_706,N_683);
nor U1039 (N_1039,N_644,N_763);
or U1040 (N_1040,N_873,N_952);
xnor U1041 (N_1041,N_996,N_586);
and U1042 (N_1042,N_623,N_921);
nor U1043 (N_1043,N_661,N_533);
and U1044 (N_1044,N_855,N_787);
nor U1045 (N_1045,N_933,N_818);
nand U1046 (N_1046,N_729,N_686);
nor U1047 (N_1047,N_577,N_805);
xor U1048 (N_1048,N_658,N_929);
and U1049 (N_1049,N_710,N_681);
nand U1050 (N_1050,N_627,N_832);
xnor U1051 (N_1051,N_878,N_897);
nand U1052 (N_1052,N_766,N_735);
and U1053 (N_1053,N_542,N_775);
nand U1054 (N_1054,N_946,N_838);
or U1055 (N_1055,N_638,N_752);
nand U1056 (N_1056,N_554,N_879);
and U1057 (N_1057,N_980,N_550);
and U1058 (N_1058,N_772,N_833);
nand U1059 (N_1059,N_786,N_672);
and U1060 (N_1060,N_981,N_730);
nor U1061 (N_1061,N_908,N_569);
nand U1062 (N_1062,N_774,N_593);
or U1063 (N_1063,N_506,N_732);
nand U1064 (N_1064,N_597,N_825);
or U1065 (N_1065,N_788,N_937);
nor U1066 (N_1066,N_758,N_560);
nor U1067 (N_1067,N_820,N_588);
or U1068 (N_1068,N_541,N_768);
and U1069 (N_1069,N_977,N_982);
nand U1070 (N_1070,N_633,N_598);
nor U1071 (N_1071,N_514,N_868);
or U1072 (N_1072,N_848,N_515);
nor U1073 (N_1073,N_875,N_892);
or U1074 (N_1074,N_876,N_762);
or U1075 (N_1075,N_656,N_857);
or U1076 (N_1076,N_864,N_549);
nor U1077 (N_1077,N_502,N_718);
nand U1078 (N_1078,N_679,N_648);
nor U1079 (N_1079,N_993,N_764);
and U1080 (N_1080,N_931,N_642);
and U1081 (N_1081,N_643,N_898);
or U1082 (N_1082,N_944,N_707);
or U1083 (N_1083,N_853,N_951);
nor U1084 (N_1084,N_570,N_746);
nand U1085 (N_1085,N_782,N_687);
or U1086 (N_1086,N_722,N_695);
nor U1087 (N_1087,N_585,N_603);
nor U1088 (N_1088,N_584,N_537);
and U1089 (N_1089,N_694,N_624);
and U1090 (N_1090,N_755,N_626);
or U1091 (N_1091,N_602,N_907);
xor U1092 (N_1092,N_817,N_799);
nor U1093 (N_1093,N_893,N_609);
nor U1094 (N_1094,N_916,N_751);
nand U1095 (N_1095,N_945,N_999);
xnor U1096 (N_1096,N_923,N_610);
nor U1097 (N_1097,N_911,N_712);
nor U1098 (N_1098,N_770,N_957);
nand U1099 (N_1099,N_927,N_819);
nor U1100 (N_1100,N_891,N_966);
and U1101 (N_1101,N_562,N_646);
and U1102 (N_1102,N_932,N_566);
and U1103 (N_1103,N_508,N_987);
and U1104 (N_1104,N_631,N_831);
nor U1105 (N_1105,N_641,N_634);
xnor U1106 (N_1106,N_716,N_605);
and U1107 (N_1107,N_872,N_500);
nor U1108 (N_1108,N_827,N_618);
nand U1109 (N_1109,N_964,N_797);
or U1110 (N_1110,N_913,N_988);
nand U1111 (N_1111,N_779,N_524);
xnor U1112 (N_1112,N_865,N_749);
nand U1113 (N_1113,N_689,N_973);
and U1114 (N_1114,N_846,N_954);
or U1115 (N_1115,N_684,N_934);
and U1116 (N_1116,N_614,N_555);
nor U1117 (N_1117,N_556,N_939);
xor U1118 (N_1118,N_914,N_956);
nand U1119 (N_1119,N_582,N_874);
and U1120 (N_1120,N_776,N_986);
nand U1121 (N_1121,N_839,N_847);
nand U1122 (N_1122,N_673,N_544);
nor U1123 (N_1123,N_998,N_619);
and U1124 (N_1124,N_769,N_635);
nand U1125 (N_1125,N_589,N_651);
nor U1126 (N_1126,N_997,N_784);
or U1127 (N_1127,N_750,N_580);
nor U1128 (N_1128,N_968,N_794);
xor U1129 (N_1129,N_528,N_906);
or U1130 (N_1130,N_639,N_559);
nand U1131 (N_1131,N_791,N_807);
nand U1132 (N_1132,N_924,N_666);
nand U1133 (N_1133,N_756,N_620);
and U1134 (N_1134,N_519,N_604);
or U1135 (N_1135,N_509,N_521);
and U1136 (N_1136,N_719,N_856);
and U1137 (N_1137,N_652,N_809);
or U1138 (N_1138,N_910,N_765);
or U1139 (N_1139,N_835,N_926);
and U1140 (N_1140,N_709,N_674);
or U1141 (N_1141,N_811,N_849);
xnor U1142 (N_1142,N_726,N_816);
xor U1143 (N_1143,N_955,N_571);
nand U1144 (N_1144,N_815,N_983);
nand U1145 (N_1145,N_930,N_915);
or U1146 (N_1146,N_690,N_715);
and U1147 (N_1147,N_994,N_522);
and U1148 (N_1148,N_861,N_731);
nand U1149 (N_1149,N_792,N_617);
nand U1150 (N_1150,N_851,N_796);
nor U1151 (N_1151,N_814,N_904);
xnor U1152 (N_1152,N_882,N_532);
nand U1153 (N_1153,N_567,N_721);
or U1154 (N_1154,N_510,N_536);
or U1155 (N_1155,N_889,N_943);
or U1156 (N_1156,N_863,N_960);
xnor U1157 (N_1157,N_967,N_840);
nor U1158 (N_1158,N_940,N_705);
and U1159 (N_1159,N_702,N_630);
nor U1160 (N_1160,N_828,N_592);
xnor U1161 (N_1161,N_979,N_901);
nand U1162 (N_1162,N_862,N_963);
nor U1163 (N_1163,N_767,N_965);
or U1164 (N_1164,N_663,N_887);
nand U1165 (N_1165,N_972,N_737);
nor U1166 (N_1166,N_747,N_785);
or U1167 (N_1167,N_824,N_516);
or U1168 (N_1168,N_742,N_783);
nand U1169 (N_1169,N_653,N_859);
nand U1170 (N_1170,N_692,N_985);
and U1171 (N_1171,N_728,N_511);
nor U1172 (N_1172,N_579,N_594);
xor U1173 (N_1173,N_659,N_953);
nand U1174 (N_1174,N_905,N_903);
nand U1175 (N_1175,N_613,N_804);
and U1176 (N_1176,N_669,N_668);
nand U1177 (N_1177,N_760,N_561);
or U1178 (N_1178,N_890,N_505);
nor U1179 (N_1179,N_667,N_708);
nor U1180 (N_1180,N_563,N_685);
xnor U1181 (N_1181,N_557,N_538);
and U1182 (N_1182,N_535,N_654);
xor U1183 (N_1183,N_991,N_739);
or U1184 (N_1184,N_670,N_518);
nor U1185 (N_1185,N_632,N_867);
nand U1186 (N_1186,N_741,N_866);
xor U1187 (N_1187,N_880,N_912);
or U1188 (N_1188,N_529,N_665);
nor U1189 (N_1189,N_717,N_829);
nand U1190 (N_1190,N_989,N_808);
or U1191 (N_1191,N_574,N_854);
and U1192 (N_1192,N_688,N_812);
and U1193 (N_1193,N_675,N_720);
nor U1194 (N_1194,N_877,N_917);
and U1195 (N_1195,N_693,N_714);
nand U1196 (N_1196,N_881,N_568);
nand U1197 (N_1197,N_795,N_941);
nand U1198 (N_1198,N_798,N_699);
or U1199 (N_1199,N_724,N_616);
nand U1200 (N_1200,N_948,N_649);
and U1201 (N_1201,N_743,N_628);
and U1202 (N_1202,N_950,N_581);
nand U1203 (N_1203,N_520,N_711);
xor U1204 (N_1204,N_920,N_680);
nand U1205 (N_1205,N_984,N_691);
xnor U1206 (N_1206,N_662,N_748);
xnor U1207 (N_1207,N_513,N_587);
or U1208 (N_1208,N_725,N_601);
and U1209 (N_1209,N_625,N_575);
nor U1210 (N_1210,N_761,N_607);
nand U1211 (N_1211,N_676,N_922);
and U1212 (N_1212,N_870,N_793);
nand U1213 (N_1213,N_629,N_744);
nand U1214 (N_1214,N_823,N_781);
nor U1215 (N_1215,N_647,N_547);
nand U1216 (N_1216,N_590,N_896);
nor U1217 (N_1217,N_843,N_844);
nand U1218 (N_1218,N_727,N_888);
nor U1219 (N_1219,N_578,N_894);
xor U1220 (N_1220,N_771,N_523);
nand U1221 (N_1221,N_949,N_935);
or U1222 (N_1222,N_697,N_700);
nor U1223 (N_1223,N_507,N_759);
or U1224 (N_1224,N_611,N_583);
and U1225 (N_1225,N_548,N_606);
nor U1226 (N_1226,N_842,N_546);
xor U1227 (N_1227,N_978,N_754);
or U1228 (N_1228,N_806,N_780);
and U1229 (N_1229,N_789,N_895);
or U1230 (N_1230,N_595,N_837);
xor U1231 (N_1231,N_678,N_539);
nor U1232 (N_1232,N_753,N_757);
and U1233 (N_1233,N_969,N_850);
nand U1234 (N_1234,N_703,N_885);
or U1235 (N_1235,N_527,N_990);
or U1236 (N_1236,N_660,N_517);
and U1237 (N_1237,N_773,N_918);
nor U1238 (N_1238,N_733,N_636);
or U1239 (N_1239,N_657,N_696);
and U1240 (N_1240,N_925,N_886);
or U1241 (N_1241,N_600,N_640);
nand U1242 (N_1242,N_645,N_974);
and U1243 (N_1243,N_902,N_664);
nand U1244 (N_1244,N_962,N_947);
nand U1245 (N_1245,N_938,N_530);
and U1246 (N_1246,N_622,N_790);
or U1247 (N_1247,N_671,N_701);
and U1248 (N_1248,N_682,N_621);
and U1249 (N_1249,N_552,N_734);
and U1250 (N_1250,N_675,N_970);
and U1251 (N_1251,N_796,N_844);
or U1252 (N_1252,N_886,N_542);
xnor U1253 (N_1253,N_623,N_583);
and U1254 (N_1254,N_832,N_752);
nand U1255 (N_1255,N_552,N_536);
nor U1256 (N_1256,N_769,N_784);
nand U1257 (N_1257,N_965,N_998);
nand U1258 (N_1258,N_729,N_769);
and U1259 (N_1259,N_740,N_730);
xor U1260 (N_1260,N_614,N_810);
nor U1261 (N_1261,N_680,N_903);
nor U1262 (N_1262,N_830,N_761);
and U1263 (N_1263,N_675,N_773);
xor U1264 (N_1264,N_789,N_827);
xor U1265 (N_1265,N_555,N_787);
nor U1266 (N_1266,N_783,N_815);
or U1267 (N_1267,N_604,N_807);
nand U1268 (N_1268,N_666,N_769);
nand U1269 (N_1269,N_619,N_632);
or U1270 (N_1270,N_641,N_636);
xor U1271 (N_1271,N_648,N_801);
xnor U1272 (N_1272,N_893,N_557);
nor U1273 (N_1273,N_725,N_724);
nand U1274 (N_1274,N_879,N_832);
nor U1275 (N_1275,N_911,N_638);
or U1276 (N_1276,N_664,N_811);
and U1277 (N_1277,N_993,N_896);
or U1278 (N_1278,N_681,N_903);
nand U1279 (N_1279,N_965,N_845);
nand U1280 (N_1280,N_888,N_754);
nor U1281 (N_1281,N_848,N_708);
and U1282 (N_1282,N_911,N_881);
nand U1283 (N_1283,N_941,N_753);
and U1284 (N_1284,N_532,N_898);
nor U1285 (N_1285,N_561,N_680);
or U1286 (N_1286,N_609,N_573);
and U1287 (N_1287,N_924,N_706);
or U1288 (N_1288,N_556,N_954);
nand U1289 (N_1289,N_818,N_901);
nor U1290 (N_1290,N_585,N_715);
and U1291 (N_1291,N_797,N_552);
nand U1292 (N_1292,N_899,N_861);
or U1293 (N_1293,N_564,N_914);
or U1294 (N_1294,N_784,N_776);
or U1295 (N_1295,N_943,N_867);
nand U1296 (N_1296,N_816,N_932);
nor U1297 (N_1297,N_599,N_667);
nor U1298 (N_1298,N_933,N_535);
nor U1299 (N_1299,N_823,N_937);
and U1300 (N_1300,N_939,N_592);
and U1301 (N_1301,N_509,N_593);
and U1302 (N_1302,N_754,N_554);
nor U1303 (N_1303,N_997,N_759);
or U1304 (N_1304,N_525,N_528);
or U1305 (N_1305,N_866,N_913);
nor U1306 (N_1306,N_587,N_676);
and U1307 (N_1307,N_949,N_895);
and U1308 (N_1308,N_553,N_867);
nor U1309 (N_1309,N_986,N_840);
and U1310 (N_1310,N_998,N_562);
and U1311 (N_1311,N_590,N_685);
nor U1312 (N_1312,N_658,N_834);
nand U1313 (N_1313,N_915,N_743);
nand U1314 (N_1314,N_925,N_616);
nor U1315 (N_1315,N_919,N_908);
nor U1316 (N_1316,N_695,N_553);
or U1317 (N_1317,N_930,N_980);
and U1318 (N_1318,N_663,N_876);
or U1319 (N_1319,N_697,N_565);
or U1320 (N_1320,N_899,N_916);
nor U1321 (N_1321,N_853,N_840);
nand U1322 (N_1322,N_984,N_513);
nand U1323 (N_1323,N_540,N_753);
or U1324 (N_1324,N_836,N_951);
and U1325 (N_1325,N_835,N_674);
nand U1326 (N_1326,N_734,N_614);
or U1327 (N_1327,N_980,N_936);
xnor U1328 (N_1328,N_862,N_519);
nor U1329 (N_1329,N_713,N_863);
nor U1330 (N_1330,N_983,N_884);
nand U1331 (N_1331,N_931,N_751);
or U1332 (N_1332,N_859,N_936);
nor U1333 (N_1333,N_763,N_600);
or U1334 (N_1334,N_750,N_528);
nor U1335 (N_1335,N_933,N_542);
or U1336 (N_1336,N_812,N_510);
nand U1337 (N_1337,N_915,N_689);
or U1338 (N_1338,N_661,N_560);
nand U1339 (N_1339,N_890,N_885);
xnor U1340 (N_1340,N_732,N_657);
nand U1341 (N_1341,N_821,N_951);
nor U1342 (N_1342,N_650,N_689);
nand U1343 (N_1343,N_538,N_704);
nor U1344 (N_1344,N_598,N_853);
or U1345 (N_1345,N_628,N_765);
or U1346 (N_1346,N_613,N_769);
nor U1347 (N_1347,N_952,N_912);
nor U1348 (N_1348,N_765,N_987);
and U1349 (N_1349,N_878,N_754);
and U1350 (N_1350,N_546,N_517);
xnor U1351 (N_1351,N_910,N_588);
nand U1352 (N_1352,N_867,N_713);
nor U1353 (N_1353,N_794,N_604);
nor U1354 (N_1354,N_947,N_525);
and U1355 (N_1355,N_597,N_509);
and U1356 (N_1356,N_859,N_528);
nor U1357 (N_1357,N_674,N_777);
xnor U1358 (N_1358,N_889,N_718);
nand U1359 (N_1359,N_909,N_878);
and U1360 (N_1360,N_935,N_818);
and U1361 (N_1361,N_513,N_614);
and U1362 (N_1362,N_622,N_960);
nand U1363 (N_1363,N_794,N_504);
nand U1364 (N_1364,N_691,N_739);
nand U1365 (N_1365,N_968,N_691);
and U1366 (N_1366,N_907,N_758);
nor U1367 (N_1367,N_609,N_877);
nor U1368 (N_1368,N_548,N_993);
and U1369 (N_1369,N_612,N_587);
or U1370 (N_1370,N_807,N_614);
nand U1371 (N_1371,N_715,N_890);
nor U1372 (N_1372,N_933,N_696);
and U1373 (N_1373,N_954,N_537);
nor U1374 (N_1374,N_612,N_624);
and U1375 (N_1375,N_804,N_870);
and U1376 (N_1376,N_993,N_734);
nor U1377 (N_1377,N_554,N_646);
or U1378 (N_1378,N_751,N_528);
or U1379 (N_1379,N_567,N_802);
and U1380 (N_1380,N_988,N_789);
xor U1381 (N_1381,N_923,N_842);
and U1382 (N_1382,N_822,N_899);
nor U1383 (N_1383,N_668,N_878);
or U1384 (N_1384,N_832,N_754);
and U1385 (N_1385,N_989,N_860);
nand U1386 (N_1386,N_873,N_801);
or U1387 (N_1387,N_557,N_550);
and U1388 (N_1388,N_660,N_897);
nand U1389 (N_1389,N_784,N_958);
and U1390 (N_1390,N_806,N_937);
nand U1391 (N_1391,N_676,N_847);
xor U1392 (N_1392,N_877,N_786);
xnor U1393 (N_1393,N_693,N_525);
and U1394 (N_1394,N_678,N_715);
and U1395 (N_1395,N_785,N_863);
nand U1396 (N_1396,N_780,N_773);
nand U1397 (N_1397,N_892,N_736);
nor U1398 (N_1398,N_858,N_552);
nand U1399 (N_1399,N_544,N_888);
and U1400 (N_1400,N_586,N_908);
or U1401 (N_1401,N_705,N_901);
nand U1402 (N_1402,N_906,N_779);
nand U1403 (N_1403,N_731,N_749);
nor U1404 (N_1404,N_950,N_860);
nor U1405 (N_1405,N_545,N_883);
nand U1406 (N_1406,N_804,N_650);
and U1407 (N_1407,N_621,N_970);
and U1408 (N_1408,N_922,N_672);
or U1409 (N_1409,N_981,N_637);
or U1410 (N_1410,N_504,N_818);
nor U1411 (N_1411,N_635,N_552);
nor U1412 (N_1412,N_683,N_864);
nand U1413 (N_1413,N_721,N_931);
or U1414 (N_1414,N_613,N_839);
or U1415 (N_1415,N_672,N_928);
or U1416 (N_1416,N_737,N_902);
nand U1417 (N_1417,N_624,N_951);
and U1418 (N_1418,N_581,N_812);
nand U1419 (N_1419,N_771,N_650);
or U1420 (N_1420,N_548,N_639);
or U1421 (N_1421,N_737,N_798);
nor U1422 (N_1422,N_754,N_616);
and U1423 (N_1423,N_947,N_724);
and U1424 (N_1424,N_645,N_857);
nor U1425 (N_1425,N_869,N_674);
and U1426 (N_1426,N_950,N_738);
nand U1427 (N_1427,N_626,N_832);
nor U1428 (N_1428,N_815,N_966);
or U1429 (N_1429,N_597,N_962);
nand U1430 (N_1430,N_717,N_611);
nor U1431 (N_1431,N_582,N_990);
nor U1432 (N_1432,N_765,N_554);
and U1433 (N_1433,N_598,N_726);
nand U1434 (N_1434,N_983,N_685);
xor U1435 (N_1435,N_747,N_959);
and U1436 (N_1436,N_500,N_734);
or U1437 (N_1437,N_868,N_607);
nor U1438 (N_1438,N_876,N_991);
nor U1439 (N_1439,N_588,N_508);
and U1440 (N_1440,N_994,N_828);
nand U1441 (N_1441,N_739,N_561);
xnor U1442 (N_1442,N_628,N_749);
or U1443 (N_1443,N_605,N_743);
or U1444 (N_1444,N_991,N_518);
nor U1445 (N_1445,N_547,N_875);
nor U1446 (N_1446,N_629,N_905);
nand U1447 (N_1447,N_525,N_909);
nor U1448 (N_1448,N_964,N_971);
and U1449 (N_1449,N_905,N_680);
or U1450 (N_1450,N_734,N_653);
nand U1451 (N_1451,N_827,N_933);
nor U1452 (N_1452,N_740,N_874);
xnor U1453 (N_1453,N_716,N_577);
nor U1454 (N_1454,N_504,N_754);
nand U1455 (N_1455,N_713,N_551);
or U1456 (N_1456,N_954,N_851);
and U1457 (N_1457,N_764,N_782);
nor U1458 (N_1458,N_788,N_722);
nand U1459 (N_1459,N_563,N_939);
nor U1460 (N_1460,N_985,N_674);
nand U1461 (N_1461,N_986,N_506);
and U1462 (N_1462,N_745,N_985);
or U1463 (N_1463,N_563,N_524);
and U1464 (N_1464,N_973,N_893);
and U1465 (N_1465,N_955,N_811);
or U1466 (N_1466,N_796,N_515);
and U1467 (N_1467,N_868,N_961);
and U1468 (N_1468,N_634,N_965);
and U1469 (N_1469,N_748,N_721);
and U1470 (N_1470,N_994,N_526);
or U1471 (N_1471,N_837,N_620);
nor U1472 (N_1472,N_775,N_847);
nor U1473 (N_1473,N_790,N_644);
nor U1474 (N_1474,N_725,N_915);
or U1475 (N_1475,N_789,N_901);
and U1476 (N_1476,N_665,N_730);
and U1477 (N_1477,N_584,N_789);
nor U1478 (N_1478,N_876,N_799);
nand U1479 (N_1479,N_955,N_694);
and U1480 (N_1480,N_658,N_905);
or U1481 (N_1481,N_864,N_816);
or U1482 (N_1482,N_508,N_874);
nor U1483 (N_1483,N_724,N_738);
nand U1484 (N_1484,N_979,N_546);
and U1485 (N_1485,N_964,N_835);
and U1486 (N_1486,N_789,N_875);
nand U1487 (N_1487,N_887,N_530);
or U1488 (N_1488,N_599,N_863);
nor U1489 (N_1489,N_603,N_613);
or U1490 (N_1490,N_670,N_645);
xor U1491 (N_1491,N_994,N_942);
nand U1492 (N_1492,N_573,N_738);
and U1493 (N_1493,N_540,N_882);
or U1494 (N_1494,N_531,N_897);
nor U1495 (N_1495,N_824,N_771);
xor U1496 (N_1496,N_988,N_876);
and U1497 (N_1497,N_573,N_967);
or U1498 (N_1498,N_625,N_814);
nor U1499 (N_1499,N_872,N_806);
nand U1500 (N_1500,N_1014,N_1478);
or U1501 (N_1501,N_1005,N_1351);
nor U1502 (N_1502,N_1272,N_1196);
and U1503 (N_1503,N_1058,N_1019);
nand U1504 (N_1504,N_1316,N_1096);
nor U1505 (N_1505,N_1353,N_1022);
and U1506 (N_1506,N_1108,N_1294);
xnor U1507 (N_1507,N_1453,N_1232);
nor U1508 (N_1508,N_1178,N_1048);
nand U1509 (N_1509,N_1053,N_1166);
or U1510 (N_1510,N_1193,N_1254);
nor U1511 (N_1511,N_1070,N_1282);
nand U1512 (N_1512,N_1361,N_1073);
or U1513 (N_1513,N_1270,N_1265);
nand U1514 (N_1514,N_1101,N_1261);
and U1515 (N_1515,N_1032,N_1391);
or U1516 (N_1516,N_1063,N_1148);
nand U1517 (N_1517,N_1304,N_1362);
nor U1518 (N_1518,N_1025,N_1332);
xor U1519 (N_1519,N_1258,N_1429);
nor U1520 (N_1520,N_1045,N_1028);
nand U1521 (N_1521,N_1203,N_1385);
and U1522 (N_1522,N_1341,N_1420);
nor U1523 (N_1523,N_1015,N_1112);
nand U1524 (N_1524,N_1320,N_1078);
and U1525 (N_1525,N_1379,N_1447);
and U1526 (N_1526,N_1100,N_1207);
or U1527 (N_1527,N_1162,N_1291);
and U1528 (N_1528,N_1010,N_1360);
nor U1529 (N_1529,N_1071,N_1230);
or U1530 (N_1530,N_1284,N_1173);
or U1531 (N_1531,N_1404,N_1457);
nor U1532 (N_1532,N_1184,N_1325);
or U1533 (N_1533,N_1264,N_1387);
or U1534 (N_1534,N_1013,N_1080);
and U1535 (N_1535,N_1378,N_1458);
and U1536 (N_1536,N_1443,N_1476);
nand U1537 (N_1537,N_1105,N_1008);
nand U1538 (N_1538,N_1036,N_1314);
nand U1539 (N_1539,N_1052,N_1283);
or U1540 (N_1540,N_1201,N_1029);
nand U1541 (N_1541,N_1170,N_1038);
or U1542 (N_1542,N_1066,N_1221);
nand U1543 (N_1543,N_1222,N_1095);
and U1544 (N_1544,N_1084,N_1090);
or U1545 (N_1545,N_1020,N_1302);
nand U1546 (N_1546,N_1384,N_1396);
nand U1547 (N_1547,N_1278,N_1017);
or U1548 (N_1548,N_1004,N_1431);
and U1549 (N_1549,N_1436,N_1299);
and U1550 (N_1550,N_1160,N_1062);
and U1551 (N_1551,N_1144,N_1410);
and U1552 (N_1552,N_1474,N_1035);
and U1553 (N_1553,N_1297,N_1397);
nor U1554 (N_1554,N_1484,N_1192);
nor U1555 (N_1555,N_1043,N_1459);
nand U1556 (N_1556,N_1466,N_1422);
nor U1557 (N_1557,N_1081,N_1295);
nor U1558 (N_1558,N_1037,N_1381);
and U1559 (N_1559,N_1167,N_1271);
xnor U1560 (N_1560,N_1357,N_1375);
nand U1561 (N_1561,N_1369,N_1155);
or U1562 (N_1562,N_1206,N_1414);
xnor U1563 (N_1563,N_1123,N_1439);
nor U1564 (N_1564,N_1285,N_1204);
nand U1565 (N_1565,N_1398,N_1076);
or U1566 (N_1566,N_1475,N_1092);
and U1567 (N_1567,N_1156,N_1141);
xor U1568 (N_1568,N_1248,N_1001);
nand U1569 (N_1569,N_1292,N_1250);
nand U1570 (N_1570,N_1229,N_1116);
nor U1571 (N_1571,N_1340,N_1403);
xor U1572 (N_1572,N_1089,N_1212);
nor U1573 (N_1573,N_1169,N_1243);
or U1574 (N_1574,N_1055,N_1305);
and U1575 (N_1575,N_1049,N_1134);
or U1576 (N_1576,N_1237,N_1269);
nor U1577 (N_1577,N_1321,N_1335);
or U1578 (N_1578,N_1149,N_1392);
nor U1579 (N_1579,N_1202,N_1275);
nor U1580 (N_1580,N_1473,N_1256);
and U1581 (N_1581,N_1068,N_1454);
or U1582 (N_1582,N_1047,N_1034);
or U1583 (N_1583,N_1483,N_1465);
or U1584 (N_1584,N_1494,N_1121);
nand U1585 (N_1585,N_1296,N_1463);
nor U1586 (N_1586,N_1138,N_1240);
nand U1587 (N_1587,N_1133,N_1370);
and U1588 (N_1588,N_1328,N_1456);
and U1589 (N_1589,N_1236,N_1041);
or U1590 (N_1590,N_1194,N_1267);
or U1591 (N_1591,N_1417,N_1452);
and U1592 (N_1592,N_1446,N_1288);
and U1593 (N_1593,N_1315,N_1077);
and U1594 (N_1594,N_1132,N_1199);
and U1595 (N_1595,N_1190,N_1338);
and U1596 (N_1596,N_1142,N_1400);
nor U1597 (N_1597,N_1147,N_1130);
nand U1598 (N_1598,N_1430,N_1437);
nor U1599 (N_1599,N_1485,N_1313);
nor U1600 (N_1600,N_1342,N_1247);
and U1601 (N_1601,N_1424,N_1383);
or U1602 (N_1602,N_1006,N_1177);
or U1603 (N_1603,N_1356,N_1083);
or U1604 (N_1604,N_1421,N_1214);
or U1605 (N_1605,N_1218,N_1471);
nor U1606 (N_1606,N_1311,N_1345);
nor U1607 (N_1607,N_1115,N_1179);
nand U1608 (N_1608,N_1493,N_1412);
and U1609 (N_1609,N_1354,N_1161);
nor U1610 (N_1610,N_1491,N_1432);
and U1611 (N_1611,N_1492,N_1349);
nor U1612 (N_1612,N_1268,N_1205);
nor U1613 (N_1613,N_1317,N_1176);
nor U1614 (N_1614,N_1064,N_1119);
or U1615 (N_1615,N_1187,N_1303);
nand U1616 (N_1616,N_1098,N_1364);
and U1617 (N_1617,N_1486,N_1257);
and U1618 (N_1618,N_1408,N_1225);
and U1619 (N_1619,N_1213,N_1109);
xnor U1620 (N_1620,N_1208,N_1394);
xor U1621 (N_1621,N_1152,N_1151);
xnor U1622 (N_1622,N_1495,N_1227);
nand U1623 (N_1623,N_1343,N_1003);
nor U1624 (N_1624,N_1125,N_1241);
xor U1625 (N_1625,N_1352,N_1406);
or U1626 (N_1626,N_1235,N_1002);
nor U1627 (N_1627,N_1046,N_1106);
nor U1628 (N_1628,N_1211,N_1300);
nor U1629 (N_1629,N_1128,N_1368);
or U1630 (N_1630,N_1310,N_1118);
or U1631 (N_1631,N_1231,N_1198);
and U1632 (N_1632,N_1031,N_1154);
and U1633 (N_1633,N_1409,N_1434);
nand U1634 (N_1634,N_1312,N_1301);
nand U1635 (N_1635,N_1181,N_1326);
or U1636 (N_1636,N_1382,N_1067);
and U1637 (N_1637,N_1079,N_1386);
or U1638 (N_1638,N_1244,N_1146);
nor U1639 (N_1639,N_1479,N_1153);
nor U1640 (N_1640,N_1188,N_1127);
or U1641 (N_1641,N_1330,N_1481);
nor U1642 (N_1642,N_1497,N_1136);
and U1643 (N_1643,N_1122,N_1371);
or U1644 (N_1644,N_1468,N_1407);
or U1645 (N_1645,N_1433,N_1441);
xor U1646 (N_1646,N_1057,N_1344);
and U1647 (N_1647,N_1060,N_1168);
xor U1648 (N_1648,N_1329,N_1273);
nand U1649 (N_1649,N_1336,N_1489);
xor U1650 (N_1650,N_1039,N_1131);
nand U1651 (N_1651,N_1103,N_1016);
xor U1652 (N_1652,N_1044,N_1224);
and U1653 (N_1653,N_1307,N_1094);
or U1654 (N_1654,N_1054,N_1099);
nand U1655 (N_1655,N_1159,N_1395);
nand U1656 (N_1656,N_1197,N_1480);
nand U1657 (N_1657,N_1334,N_1255);
or U1658 (N_1658,N_1467,N_1377);
nand U1659 (N_1659,N_1117,N_1007);
nor U1660 (N_1660,N_1027,N_1435);
or U1661 (N_1661,N_1065,N_1346);
nor U1662 (N_1662,N_1263,N_1318);
and U1663 (N_1663,N_1000,N_1350);
or U1664 (N_1664,N_1373,N_1145);
and U1665 (N_1665,N_1365,N_1274);
nor U1666 (N_1666,N_1135,N_1220);
nor U1667 (N_1667,N_1245,N_1327);
and U1668 (N_1668,N_1171,N_1498);
nor U1669 (N_1669,N_1140,N_1215);
nand U1670 (N_1670,N_1180,N_1189);
nor U1671 (N_1671,N_1411,N_1359);
nand U1672 (N_1672,N_1246,N_1487);
xor U1673 (N_1673,N_1279,N_1195);
nand U1674 (N_1674,N_1238,N_1075);
nor U1675 (N_1675,N_1388,N_1413);
nand U1676 (N_1676,N_1488,N_1009);
and U1677 (N_1677,N_1438,N_1219);
or U1678 (N_1678,N_1448,N_1158);
or U1679 (N_1679,N_1042,N_1372);
nand U1680 (N_1680,N_1186,N_1234);
and U1681 (N_1681,N_1293,N_1499);
nor U1682 (N_1682,N_1376,N_1126);
xor U1683 (N_1683,N_1228,N_1209);
nor U1684 (N_1684,N_1088,N_1290);
or U1685 (N_1685,N_1223,N_1040);
or U1686 (N_1686,N_1110,N_1389);
nor U1687 (N_1687,N_1374,N_1324);
nand U1688 (N_1688,N_1012,N_1150);
nand U1689 (N_1689,N_1026,N_1276);
nand U1690 (N_1690,N_1440,N_1306);
or U1691 (N_1691,N_1451,N_1210);
or U1692 (N_1692,N_1124,N_1085);
nand U1693 (N_1693,N_1113,N_1086);
or U1694 (N_1694,N_1280,N_1470);
and U1695 (N_1695,N_1143,N_1464);
or U1696 (N_1696,N_1051,N_1174);
nor U1697 (N_1697,N_1427,N_1490);
nor U1698 (N_1698,N_1164,N_1418);
nor U1699 (N_1699,N_1426,N_1129);
or U1700 (N_1700,N_1337,N_1097);
and U1701 (N_1701,N_1091,N_1157);
nand U1702 (N_1702,N_1281,N_1242);
nor U1703 (N_1703,N_1074,N_1323);
or U1704 (N_1704,N_1226,N_1163);
nor U1705 (N_1705,N_1460,N_1200);
or U1706 (N_1706,N_1423,N_1030);
or U1707 (N_1707,N_1309,N_1107);
and U1708 (N_1708,N_1216,N_1355);
or U1709 (N_1709,N_1322,N_1056);
or U1710 (N_1710,N_1185,N_1380);
and U1711 (N_1711,N_1333,N_1191);
or U1712 (N_1712,N_1018,N_1183);
nor U1713 (N_1713,N_1445,N_1114);
or U1714 (N_1714,N_1358,N_1393);
nand U1715 (N_1715,N_1120,N_1239);
nand U1716 (N_1716,N_1286,N_1419);
and U1717 (N_1717,N_1455,N_1469);
nand U1718 (N_1718,N_1401,N_1172);
xor U1719 (N_1719,N_1348,N_1050);
and U1720 (N_1720,N_1450,N_1021);
nor U1721 (N_1721,N_1496,N_1182);
or U1722 (N_1722,N_1308,N_1259);
or U1723 (N_1723,N_1482,N_1425);
xor U1724 (N_1724,N_1069,N_1102);
and U1725 (N_1725,N_1462,N_1233);
or U1726 (N_1726,N_1087,N_1428);
nor U1727 (N_1727,N_1266,N_1472);
nor U1728 (N_1728,N_1024,N_1347);
nor U1729 (N_1729,N_1390,N_1175);
and U1730 (N_1730,N_1277,N_1477);
or U1731 (N_1731,N_1298,N_1367);
xor U1732 (N_1732,N_1319,N_1444);
nand U1733 (N_1733,N_1137,N_1251);
and U1734 (N_1734,N_1405,N_1072);
or U1735 (N_1735,N_1416,N_1442);
xnor U1736 (N_1736,N_1033,N_1363);
and U1737 (N_1737,N_1093,N_1287);
xnor U1738 (N_1738,N_1252,N_1111);
xnor U1739 (N_1739,N_1061,N_1260);
and U1740 (N_1740,N_1253,N_1461);
nand U1741 (N_1741,N_1402,N_1366);
nand U1742 (N_1742,N_1415,N_1217);
or U1743 (N_1743,N_1011,N_1249);
nor U1744 (N_1744,N_1331,N_1289);
nor U1745 (N_1745,N_1082,N_1059);
or U1746 (N_1746,N_1165,N_1449);
nor U1747 (N_1747,N_1339,N_1139);
nor U1748 (N_1748,N_1104,N_1023);
or U1749 (N_1749,N_1262,N_1399);
and U1750 (N_1750,N_1220,N_1363);
and U1751 (N_1751,N_1053,N_1464);
or U1752 (N_1752,N_1185,N_1088);
and U1753 (N_1753,N_1249,N_1371);
nor U1754 (N_1754,N_1037,N_1456);
xnor U1755 (N_1755,N_1317,N_1046);
nand U1756 (N_1756,N_1388,N_1338);
nor U1757 (N_1757,N_1382,N_1438);
xor U1758 (N_1758,N_1302,N_1265);
or U1759 (N_1759,N_1411,N_1099);
and U1760 (N_1760,N_1397,N_1204);
nor U1761 (N_1761,N_1162,N_1386);
nand U1762 (N_1762,N_1182,N_1000);
nand U1763 (N_1763,N_1199,N_1213);
nand U1764 (N_1764,N_1448,N_1036);
xor U1765 (N_1765,N_1140,N_1194);
and U1766 (N_1766,N_1199,N_1127);
nor U1767 (N_1767,N_1488,N_1089);
nor U1768 (N_1768,N_1239,N_1398);
or U1769 (N_1769,N_1425,N_1308);
and U1770 (N_1770,N_1225,N_1476);
xor U1771 (N_1771,N_1472,N_1101);
nand U1772 (N_1772,N_1450,N_1123);
xnor U1773 (N_1773,N_1442,N_1079);
nor U1774 (N_1774,N_1150,N_1352);
nand U1775 (N_1775,N_1038,N_1179);
or U1776 (N_1776,N_1136,N_1153);
xnor U1777 (N_1777,N_1192,N_1058);
or U1778 (N_1778,N_1194,N_1062);
and U1779 (N_1779,N_1357,N_1180);
nand U1780 (N_1780,N_1288,N_1363);
or U1781 (N_1781,N_1273,N_1258);
or U1782 (N_1782,N_1043,N_1423);
xnor U1783 (N_1783,N_1028,N_1141);
nor U1784 (N_1784,N_1146,N_1279);
nor U1785 (N_1785,N_1108,N_1135);
or U1786 (N_1786,N_1395,N_1002);
or U1787 (N_1787,N_1490,N_1338);
nand U1788 (N_1788,N_1472,N_1347);
or U1789 (N_1789,N_1296,N_1124);
nand U1790 (N_1790,N_1354,N_1366);
nor U1791 (N_1791,N_1169,N_1452);
or U1792 (N_1792,N_1214,N_1441);
nand U1793 (N_1793,N_1367,N_1277);
or U1794 (N_1794,N_1283,N_1279);
or U1795 (N_1795,N_1494,N_1492);
or U1796 (N_1796,N_1259,N_1388);
and U1797 (N_1797,N_1368,N_1490);
or U1798 (N_1798,N_1187,N_1181);
nor U1799 (N_1799,N_1462,N_1050);
and U1800 (N_1800,N_1462,N_1030);
nor U1801 (N_1801,N_1010,N_1262);
nand U1802 (N_1802,N_1079,N_1320);
nor U1803 (N_1803,N_1379,N_1258);
and U1804 (N_1804,N_1005,N_1245);
and U1805 (N_1805,N_1403,N_1456);
and U1806 (N_1806,N_1226,N_1385);
or U1807 (N_1807,N_1179,N_1336);
and U1808 (N_1808,N_1023,N_1498);
nand U1809 (N_1809,N_1106,N_1104);
nand U1810 (N_1810,N_1005,N_1481);
or U1811 (N_1811,N_1127,N_1443);
nand U1812 (N_1812,N_1473,N_1126);
or U1813 (N_1813,N_1417,N_1091);
nand U1814 (N_1814,N_1257,N_1105);
nand U1815 (N_1815,N_1041,N_1168);
and U1816 (N_1816,N_1382,N_1112);
or U1817 (N_1817,N_1252,N_1393);
or U1818 (N_1818,N_1407,N_1287);
and U1819 (N_1819,N_1122,N_1146);
nand U1820 (N_1820,N_1261,N_1426);
and U1821 (N_1821,N_1348,N_1062);
or U1822 (N_1822,N_1325,N_1373);
or U1823 (N_1823,N_1001,N_1014);
nor U1824 (N_1824,N_1262,N_1208);
nor U1825 (N_1825,N_1261,N_1349);
nand U1826 (N_1826,N_1115,N_1000);
or U1827 (N_1827,N_1054,N_1247);
xnor U1828 (N_1828,N_1296,N_1408);
and U1829 (N_1829,N_1240,N_1418);
or U1830 (N_1830,N_1326,N_1052);
or U1831 (N_1831,N_1314,N_1294);
and U1832 (N_1832,N_1400,N_1039);
nand U1833 (N_1833,N_1276,N_1037);
or U1834 (N_1834,N_1012,N_1395);
nor U1835 (N_1835,N_1132,N_1188);
or U1836 (N_1836,N_1086,N_1059);
xor U1837 (N_1837,N_1212,N_1088);
nor U1838 (N_1838,N_1205,N_1140);
or U1839 (N_1839,N_1405,N_1056);
nand U1840 (N_1840,N_1118,N_1176);
or U1841 (N_1841,N_1001,N_1116);
nand U1842 (N_1842,N_1024,N_1454);
xnor U1843 (N_1843,N_1439,N_1033);
and U1844 (N_1844,N_1261,N_1270);
nand U1845 (N_1845,N_1473,N_1378);
nand U1846 (N_1846,N_1209,N_1374);
and U1847 (N_1847,N_1484,N_1088);
and U1848 (N_1848,N_1308,N_1017);
or U1849 (N_1849,N_1030,N_1396);
and U1850 (N_1850,N_1214,N_1399);
nor U1851 (N_1851,N_1199,N_1277);
nand U1852 (N_1852,N_1240,N_1253);
and U1853 (N_1853,N_1496,N_1230);
nor U1854 (N_1854,N_1130,N_1311);
nand U1855 (N_1855,N_1093,N_1131);
and U1856 (N_1856,N_1211,N_1086);
and U1857 (N_1857,N_1029,N_1386);
and U1858 (N_1858,N_1372,N_1445);
and U1859 (N_1859,N_1469,N_1434);
nor U1860 (N_1860,N_1133,N_1251);
or U1861 (N_1861,N_1309,N_1094);
nor U1862 (N_1862,N_1247,N_1412);
xnor U1863 (N_1863,N_1437,N_1479);
nor U1864 (N_1864,N_1190,N_1085);
and U1865 (N_1865,N_1002,N_1195);
nand U1866 (N_1866,N_1487,N_1025);
xnor U1867 (N_1867,N_1209,N_1333);
and U1868 (N_1868,N_1039,N_1186);
or U1869 (N_1869,N_1061,N_1451);
nor U1870 (N_1870,N_1104,N_1011);
and U1871 (N_1871,N_1112,N_1050);
or U1872 (N_1872,N_1429,N_1326);
nor U1873 (N_1873,N_1033,N_1283);
and U1874 (N_1874,N_1237,N_1324);
nand U1875 (N_1875,N_1060,N_1204);
xor U1876 (N_1876,N_1276,N_1488);
and U1877 (N_1877,N_1389,N_1441);
nand U1878 (N_1878,N_1173,N_1407);
nor U1879 (N_1879,N_1185,N_1026);
xnor U1880 (N_1880,N_1171,N_1376);
and U1881 (N_1881,N_1388,N_1181);
or U1882 (N_1882,N_1418,N_1168);
nand U1883 (N_1883,N_1043,N_1230);
or U1884 (N_1884,N_1094,N_1440);
nor U1885 (N_1885,N_1077,N_1072);
nand U1886 (N_1886,N_1429,N_1254);
or U1887 (N_1887,N_1295,N_1226);
nor U1888 (N_1888,N_1309,N_1361);
and U1889 (N_1889,N_1439,N_1395);
and U1890 (N_1890,N_1004,N_1400);
nor U1891 (N_1891,N_1263,N_1218);
or U1892 (N_1892,N_1496,N_1195);
xor U1893 (N_1893,N_1023,N_1236);
nand U1894 (N_1894,N_1074,N_1070);
and U1895 (N_1895,N_1313,N_1339);
nand U1896 (N_1896,N_1043,N_1253);
nor U1897 (N_1897,N_1282,N_1495);
nor U1898 (N_1898,N_1068,N_1493);
nor U1899 (N_1899,N_1378,N_1282);
nor U1900 (N_1900,N_1074,N_1238);
and U1901 (N_1901,N_1403,N_1440);
and U1902 (N_1902,N_1394,N_1034);
or U1903 (N_1903,N_1404,N_1275);
nor U1904 (N_1904,N_1422,N_1102);
and U1905 (N_1905,N_1102,N_1356);
and U1906 (N_1906,N_1107,N_1180);
nand U1907 (N_1907,N_1401,N_1429);
nor U1908 (N_1908,N_1308,N_1054);
xnor U1909 (N_1909,N_1414,N_1427);
nand U1910 (N_1910,N_1467,N_1465);
nor U1911 (N_1911,N_1440,N_1350);
and U1912 (N_1912,N_1392,N_1222);
or U1913 (N_1913,N_1017,N_1166);
nor U1914 (N_1914,N_1034,N_1123);
or U1915 (N_1915,N_1024,N_1097);
nand U1916 (N_1916,N_1120,N_1375);
nand U1917 (N_1917,N_1190,N_1079);
and U1918 (N_1918,N_1360,N_1388);
nand U1919 (N_1919,N_1246,N_1195);
or U1920 (N_1920,N_1408,N_1279);
and U1921 (N_1921,N_1061,N_1257);
nand U1922 (N_1922,N_1454,N_1104);
nand U1923 (N_1923,N_1285,N_1321);
xor U1924 (N_1924,N_1430,N_1310);
nand U1925 (N_1925,N_1385,N_1341);
xnor U1926 (N_1926,N_1200,N_1333);
and U1927 (N_1927,N_1248,N_1302);
or U1928 (N_1928,N_1210,N_1303);
or U1929 (N_1929,N_1023,N_1000);
nor U1930 (N_1930,N_1255,N_1392);
and U1931 (N_1931,N_1241,N_1351);
or U1932 (N_1932,N_1339,N_1281);
nand U1933 (N_1933,N_1038,N_1027);
and U1934 (N_1934,N_1483,N_1210);
or U1935 (N_1935,N_1187,N_1006);
nand U1936 (N_1936,N_1380,N_1453);
nand U1937 (N_1937,N_1222,N_1132);
or U1938 (N_1938,N_1263,N_1378);
or U1939 (N_1939,N_1064,N_1367);
nor U1940 (N_1940,N_1220,N_1225);
or U1941 (N_1941,N_1275,N_1062);
xor U1942 (N_1942,N_1080,N_1380);
xor U1943 (N_1943,N_1337,N_1351);
and U1944 (N_1944,N_1423,N_1352);
or U1945 (N_1945,N_1426,N_1400);
and U1946 (N_1946,N_1325,N_1297);
nand U1947 (N_1947,N_1323,N_1231);
nor U1948 (N_1948,N_1279,N_1088);
nand U1949 (N_1949,N_1235,N_1478);
nor U1950 (N_1950,N_1086,N_1484);
xor U1951 (N_1951,N_1108,N_1304);
nand U1952 (N_1952,N_1384,N_1292);
nand U1953 (N_1953,N_1147,N_1004);
xor U1954 (N_1954,N_1031,N_1285);
nor U1955 (N_1955,N_1400,N_1293);
and U1956 (N_1956,N_1216,N_1335);
or U1957 (N_1957,N_1251,N_1288);
xnor U1958 (N_1958,N_1139,N_1314);
and U1959 (N_1959,N_1186,N_1076);
nor U1960 (N_1960,N_1100,N_1493);
nor U1961 (N_1961,N_1012,N_1110);
or U1962 (N_1962,N_1221,N_1262);
and U1963 (N_1963,N_1270,N_1263);
and U1964 (N_1964,N_1269,N_1105);
nand U1965 (N_1965,N_1426,N_1258);
nand U1966 (N_1966,N_1089,N_1329);
nand U1967 (N_1967,N_1017,N_1197);
and U1968 (N_1968,N_1298,N_1005);
and U1969 (N_1969,N_1387,N_1100);
nand U1970 (N_1970,N_1297,N_1271);
nor U1971 (N_1971,N_1037,N_1277);
nand U1972 (N_1972,N_1173,N_1297);
or U1973 (N_1973,N_1397,N_1084);
nor U1974 (N_1974,N_1418,N_1137);
nor U1975 (N_1975,N_1316,N_1180);
or U1976 (N_1976,N_1083,N_1328);
nand U1977 (N_1977,N_1189,N_1305);
nor U1978 (N_1978,N_1483,N_1395);
or U1979 (N_1979,N_1180,N_1346);
and U1980 (N_1980,N_1053,N_1387);
and U1981 (N_1981,N_1468,N_1159);
nor U1982 (N_1982,N_1073,N_1461);
nand U1983 (N_1983,N_1242,N_1023);
nor U1984 (N_1984,N_1037,N_1454);
nand U1985 (N_1985,N_1363,N_1058);
or U1986 (N_1986,N_1251,N_1257);
nand U1987 (N_1987,N_1159,N_1126);
nand U1988 (N_1988,N_1433,N_1338);
and U1989 (N_1989,N_1354,N_1097);
or U1990 (N_1990,N_1013,N_1148);
and U1991 (N_1991,N_1278,N_1267);
nor U1992 (N_1992,N_1156,N_1381);
nor U1993 (N_1993,N_1204,N_1376);
and U1994 (N_1994,N_1314,N_1250);
nand U1995 (N_1995,N_1074,N_1395);
nor U1996 (N_1996,N_1315,N_1314);
nand U1997 (N_1997,N_1411,N_1169);
nand U1998 (N_1998,N_1202,N_1177);
nor U1999 (N_1999,N_1189,N_1280);
nand U2000 (N_2000,N_1927,N_1807);
nand U2001 (N_2001,N_1622,N_1873);
nand U2002 (N_2002,N_1975,N_1752);
nor U2003 (N_2003,N_1683,N_1598);
xnor U2004 (N_2004,N_1884,N_1613);
nor U2005 (N_2005,N_1582,N_1788);
nor U2006 (N_2006,N_1737,N_1718);
nand U2007 (N_2007,N_1572,N_1559);
nand U2008 (N_2008,N_1770,N_1554);
nand U2009 (N_2009,N_1930,N_1716);
nand U2010 (N_2010,N_1519,N_1581);
and U2011 (N_2011,N_1684,N_1655);
nor U2012 (N_2012,N_1616,N_1506);
xor U2013 (N_2013,N_1798,N_1571);
nor U2014 (N_2014,N_1819,N_1955);
nor U2015 (N_2015,N_1913,N_1841);
and U2016 (N_2016,N_1688,N_1646);
and U2017 (N_2017,N_1544,N_1829);
or U2018 (N_2018,N_1886,N_1708);
and U2019 (N_2019,N_1721,N_1872);
and U2020 (N_2020,N_1689,N_1508);
xor U2021 (N_2021,N_1533,N_1522);
or U2022 (N_2022,N_1728,N_1738);
nand U2023 (N_2023,N_1957,N_1909);
and U2024 (N_2024,N_1833,N_1802);
xnor U2025 (N_2025,N_1670,N_1625);
or U2026 (N_2026,N_1686,N_1675);
and U2027 (N_2027,N_1780,N_1972);
or U2028 (N_2028,N_1871,N_1532);
nand U2029 (N_2029,N_1535,N_1576);
and U2030 (N_2030,N_1887,N_1612);
and U2031 (N_2031,N_1722,N_1929);
nor U2032 (N_2032,N_1593,N_1850);
nand U2033 (N_2033,N_1600,N_1945);
or U2034 (N_2034,N_1846,N_1771);
nor U2035 (N_2035,N_1792,N_1667);
and U2036 (N_2036,N_1836,N_1500);
nor U2037 (N_2037,N_1740,N_1720);
xnor U2038 (N_2038,N_1677,N_1697);
nor U2039 (N_2039,N_1703,N_1779);
or U2040 (N_2040,N_1628,N_1803);
and U2041 (N_2041,N_1526,N_1735);
nand U2042 (N_2042,N_1632,N_1690);
or U2043 (N_2043,N_1777,N_1503);
nand U2044 (N_2044,N_1907,N_1524);
nand U2045 (N_2045,N_1513,N_1620);
nor U2046 (N_2046,N_1789,N_1637);
or U2047 (N_2047,N_1996,N_1758);
nand U2048 (N_2048,N_1921,N_1812);
and U2049 (N_2049,N_1960,N_1521);
and U2050 (N_2050,N_1710,N_1530);
and U2051 (N_2051,N_1865,N_1711);
nand U2052 (N_2052,N_1810,N_1669);
nand U2053 (N_2053,N_1992,N_1561);
and U2054 (N_2054,N_1741,N_1531);
or U2055 (N_2055,N_1775,N_1785);
and U2056 (N_2056,N_1860,N_1980);
nand U2057 (N_2057,N_1952,N_1864);
nor U2058 (N_2058,N_1774,N_1617);
nor U2059 (N_2059,N_1642,N_1650);
or U2060 (N_2060,N_1555,N_1847);
and U2061 (N_2061,N_1589,N_1848);
nor U2062 (N_2062,N_1984,N_1811);
or U2063 (N_2063,N_1974,N_1851);
nand U2064 (N_2064,N_1587,N_1990);
or U2065 (N_2065,N_1967,N_1993);
xnor U2066 (N_2066,N_1528,N_1880);
nand U2067 (N_2067,N_1795,N_1977);
nand U2068 (N_2068,N_1680,N_1827);
nor U2069 (N_2069,N_1712,N_1797);
or U2070 (N_2070,N_1610,N_1601);
and U2071 (N_2071,N_1910,N_1895);
or U2072 (N_2072,N_1941,N_1515);
or U2073 (N_2073,N_1618,N_1825);
and U2074 (N_2074,N_1552,N_1736);
and U2075 (N_2075,N_1747,N_1653);
nor U2076 (N_2076,N_1707,N_1982);
nand U2077 (N_2077,N_1664,N_1994);
nand U2078 (N_2078,N_1558,N_1787);
or U2079 (N_2079,N_1963,N_1983);
nor U2080 (N_2080,N_1687,N_1536);
nor U2081 (N_2081,N_1824,N_1892);
nand U2082 (N_2082,N_1548,N_1856);
nor U2083 (N_2083,N_1916,N_1549);
nor U2084 (N_2084,N_1999,N_1845);
xor U2085 (N_2085,N_1938,N_1609);
and U2086 (N_2086,N_1654,N_1926);
or U2087 (N_2087,N_1764,N_1691);
nand U2088 (N_2088,N_1917,N_1937);
and U2089 (N_2089,N_1709,N_1849);
or U2090 (N_2090,N_1765,N_1804);
or U2091 (N_2091,N_1896,N_1665);
xor U2092 (N_2092,N_1885,N_1585);
or U2093 (N_2093,N_1959,N_1900);
nand U2094 (N_2094,N_1776,N_1726);
and U2095 (N_2095,N_1783,N_1744);
nand U2096 (N_2096,N_1782,N_1615);
or U2097 (N_2097,N_1767,N_1987);
nand U2098 (N_2098,N_1590,N_1922);
nand U2099 (N_2099,N_1640,N_1925);
and U2100 (N_2100,N_1878,N_1899);
and U2101 (N_2101,N_1979,N_1773);
or U2102 (N_2102,N_1826,N_1934);
or U2103 (N_2103,N_1954,N_1599);
or U2104 (N_2104,N_1951,N_1820);
and U2105 (N_2105,N_1969,N_1840);
or U2106 (N_2106,N_1717,N_1801);
and U2107 (N_2107,N_1540,N_1725);
and U2108 (N_2108,N_1762,N_1939);
or U2109 (N_2109,N_1908,N_1748);
or U2110 (N_2110,N_1897,N_1918);
nor U2111 (N_2111,N_1839,N_1766);
nand U2112 (N_2112,N_1817,N_1502);
nand U2113 (N_2113,N_1681,N_1893);
and U2114 (N_2114,N_1924,N_1568);
nor U2115 (N_2115,N_1719,N_1869);
xnor U2116 (N_2116,N_1518,N_1673);
nand U2117 (N_2117,N_1901,N_1631);
or U2118 (N_2118,N_1603,N_1875);
or U2119 (N_2119,N_1523,N_1757);
and U2120 (N_2120,N_1932,N_1547);
nor U2121 (N_2121,N_1731,N_1835);
nor U2122 (N_2122,N_1695,N_1877);
or U2123 (N_2123,N_1838,N_1739);
and U2124 (N_2124,N_1964,N_1574);
and U2125 (N_2125,N_1986,N_1541);
xor U2126 (N_2126,N_1715,N_1816);
xnor U2127 (N_2127,N_1511,N_1671);
nand U2128 (N_2128,N_1751,N_1753);
and U2129 (N_2129,N_1516,N_1727);
and U2130 (N_2130,N_1904,N_1696);
or U2131 (N_2131,N_1557,N_1543);
or U2132 (N_2132,N_1584,N_1633);
xnor U2133 (N_2133,N_1966,N_1867);
and U2134 (N_2134,N_1823,N_1855);
and U2135 (N_2135,N_1988,N_1588);
xnor U2136 (N_2136,N_1950,N_1520);
and U2137 (N_2137,N_1635,N_1958);
nand U2138 (N_2138,N_1575,N_1693);
and U2139 (N_2139,N_1942,N_1551);
or U2140 (N_2140,N_1949,N_1553);
xor U2141 (N_2141,N_1881,N_1989);
nor U2142 (N_2142,N_1874,N_1834);
nand U2143 (N_2143,N_1976,N_1517);
nand U2144 (N_2144,N_1702,N_1981);
nand U2145 (N_2145,N_1911,N_1538);
nand U2146 (N_2146,N_1843,N_1882);
or U2147 (N_2147,N_1563,N_1594);
nor U2148 (N_2148,N_1651,N_1808);
nor U2149 (N_2149,N_1906,N_1923);
or U2150 (N_2150,N_1743,N_1894);
nor U2151 (N_2151,N_1933,N_1602);
or U2152 (N_2152,N_1556,N_1772);
or U2153 (N_2153,N_1668,N_1946);
nor U2154 (N_2154,N_1970,N_1573);
xnor U2155 (N_2155,N_1888,N_1705);
or U2156 (N_2156,N_1944,N_1604);
xor U2157 (N_2157,N_1562,N_1962);
nand U2158 (N_2158,N_1914,N_1968);
or U2159 (N_2159,N_1978,N_1624);
and U2160 (N_2160,N_1746,N_1868);
or U2161 (N_2161,N_1997,N_1936);
or U2162 (N_2162,N_1956,N_1569);
and U2163 (N_2163,N_1991,N_1611);
nor U2164 (N_2164,N_1733,N_1920);
and U2165 (N_2165,N_1662,N_1545);
nor U2166 (N_2166,N_1828,N_1876);
nand U2167 (N_2167,N_1948,N_1786);
nor U2168 (N_2168,N_1866,N_1619);
and U2169 (N_2169,N_1799,N_1639);
or U2170 (N_2170,N_1723,N_1935);
or U2171 (N_2171,N_1755,N_1698);
nand U2172 (N_2172,N_1605,N_1529);
or U2173 (N_2173,N_1706,N_1586);
and U2174 (N_2174,N_1760,N_1621);
nand U2175 (N_2175,N_1915,N_1761);
nand U2176 (N_2176,N_1636,N_1870);
and U2177 (N_2177,N_1537,N_1634);
nor U2178 (N_2178,N_1890,N_1995);
nand U2179 (N_2179,N_1729,N_1863);
and U2180 (N_2180,N_1608,N_1854);
or U2181 (N_2181,N_1732,N_1793);
and U2182 (N_2182,N_1592,N_1791);
nor U2183 (N_2183,N_1660,N_1769);
xor U2184 (N_2184,N_1831,N_1796);
nor U2185 (N_2185,N_1629,N_1837);
and U2186 (N_2186,N_1853,N_1965);
and U2187 (N_2187,N_1504,N_1596);
and U2188 (N_2188,N_1985,N_1560);
nand U2189 (N_2189,N_1694,N_1679);
or U2190 (N_2190,N_1861,N_1658);
and U2191 (N_2191,N_1657,N_1510);
nor U2192 (N_2192,N_1685,N_1832);
or U2193 (N_2193,N_1507,N_1701);
xor U2194 (N_2194,N_1889,N_1822);
xnor U2195 (N_2195,N_1809,N_1614);
or U2196 (N_2196,N_1534,N_1713);
xnor U2197 (N_2197,N_1704,N_1644);
or U2198 (N_2198,N_1891,N_1659);
xor U2199 (N_2199,N_1842,N_1857);
nor U2200 (N_2200,N_1768,N_1566);
nor U2201 (N_2201,N_1943,N_1591);
nor U2202 (N_2202,N_1649,N_1645);
nor U2203 (N_2203,N_1953,N_1903);
nand U2204 (N_2204,N_1501,N_1666);
and U2205 (N_2205,N_1577,N_1879);
or U2206 (N_2206,N_1940,N_1902);
nand U2207 (N_2207,N_1626,N_1778);
nor U2208 (N_2208,N_1759,N_1998);
or U2209 (N_2209,N_1539,N_1597);
or U2210 (N_2210,N_1700,N_1971);
xnor U2211 (N_2211,N_1674,N_1742);
or U2212 (N_2212,N_1606,N_1805);
or U2213 (N_2213,N_1542,N_1578);
nor U2214 (N_2214,N_1734,N_1567);
and U2215 (N_2215,N_1905,N_1595);
nand U2216 (N_2216,N_1790,N_1883);
nor U2217 (N_2217,N_1564,N_1678);
or U2218 (N_2218,N_1749,N_1763);
or U2219 (N_2219,N_1583,N_1699);
nand U2220 (N_2220,N_1745,N_1730);
nand U2221 (N_2221,N_1919,N_1565);
and U2222 (N_2222,N_1676,N_1579);
nand U2223 (N_2223,N_1830,N_1928);
nor U2224 (N_2224,N_1821,N_1648);
or U2225 (N_2225,N_1931,N_1794);
and U2226 (N_2226,N_1750,N_1754);
or U2227 (N_2227,N_1550,N_1814);
or U2228 (N_2228,N_1858,N_1844);
or U2229 (N_2229,N_1512,N_1813);
or U2230 (N_2230,N_1912,N_1509);
nor U2231 (N_2231,N_1692,N_1527);
or U2232 (N_2232,N_1661,N_1514);
xor U2233 (N_2233,N_1862,N_1630);
nor U2234 (N_2234,N_1570,N_1898);
nand U2235 (N_2235,N_1973,N_1818);
nor U2236 (N_2236,N_1672,N_1724);
and U2237 (N_2237,N_1800,N_1961);
and U2238 (N_2238,N_1546,N_1852);
or U2239 (N_2239,N_1781,N_1638);
or U2240 (N_2240,N_1505,N_1682);
or U2241 (N_2241,N_1647,N_1652);
nand U2242 (N_2242,N_1643,N_1756);
and U2243 (N_2243,N_1714,N_1806);
nor U2244 (N_2244,N_1627,N_1656);
and U2245 (N_2245,N_1580,N_1623);
or U2246 (N_2246,N_1663,N_1641);
or U2247 (N_2247,N_1525,N_1607);
and U2248 (N_2248,N_1784,N_1815);
or U2249 (N_2249,N_1859,N_1947);
xnor U2250 (N_2250,N_1806,N_1778);
nor U2251 (N_2251,N_1837,N_1901);
xnor U2252 (N_2252,N_1880,N_1819);
nand U2253 (N_2253,N_1557,N_1975);
nand U2254 (N_2254,N_1877,N_1518);
and U2255 (N_2255,N_1879,N_1976);
and U2256 (N_2256,N_1570,N_1740);
and U2257 (N_2257,N_1725,N_1526);
nor U2258 (N_2258,N_1759,N_1878);
or U2259 (N_2259,N_1978,N_1988);
nor U2260 (N_2260,N_1851,N_1757);
nor U2261 (N_2261,N_1875,N_1857);
or U2262 (N_2262,N_1958,N_1746);
nor U2263 (N_2263,N_1976,N_1571);
nor U2264 (N_2264,N_1984,N_1708);
nand U2265 (N_2265,N_1849,N_1937);
and U2266 (N_2266,N_1685,N_1628);
or U2267 (N_2267,N_1546,N_1597);
or U2268 (N_2268,N_1607,N_1614);
or U2269 (N_2269,N_1611,N_1803);
or U2270 (N_2270,N_1614,N_1658);
and U2271 (N_2271,N_1629,N_1875);
nor U2272 (N_2272,N_1680,N_1966);
nor U2273 (N_2273,N_1997,N_1829);
nand U2274 (N_2274,N_1873,N_1633);
or U2275 (N_2275,N_1912,N_1636);
xnor U2276 (N_2276,N_1736,N_1731);
nor U2277 (N_2277,N_1895,N_1977);
nor U2278 (N_2278,N_1967,N_1880);
nor U2279 (N_2279,N_1603,N_1662);
and U2280 (N_2280,N_1727,N_1697);
nand U2281 (N_2281,N_1926,N_1973);
nand U2282 (N_2282,N_1880,N_1841);
nand U2283 (N_2283,N_1948,N_1732);
and U2284 (N_2284,N_1949,N_1933);
nand U2285 (N_2285,N_1952,N_1715);
nand U2286 (N_2286,N_1558,N_1745);
nand U2287 (N_2287,N_1807,N_1680);
xnor U2288 (N_2288,N_1614,N_1582);
nand U2289 (N_2289,N_1820,N_1840);
and U2290 (N_2290,N_1520,N_1911);
and U2291 (N_2291,N_1919,N_1507);
nor U2292 (N_2292,N_1649,N_1790);
nor U2293 (N_2293,N_1782,N_1724);
nand U2294 (N_2294,N_1507,N_1869);
or U2295 (N_2295,N_1529,N_1687);
and U2296 (N_2296,N_1725,N_1935);
nand U2297 (N_2297,N_1736,N_1576);
and U2298 (N_2298,N_1678,N_1865);
or U2299 (N_2299,N_1517,N_1658);
and U2300 (N_2300,N_1608,N_1579);
and U2301 (N_2301,N_1962,N_1704);
nand U2302 (N_2302,N_1777,N_1670);
or U2303 (N_2303,N_1557,N_1965);
xnor U2304 (N_2304,N_1644,N_1637);
xor U2305 (N_2305,N_1593,N_1953);
and U2306 (N_2306,N_1714,N_1963);
nor U2307 (N_2307,N_1969,N_1712);
xnor U2308 (N_2308,N_1726,N_1589);
and U2309 (N_2309,N_1690,N_1744);
xnor U2310 (N_2310,N_1695,N_1984);
nor U2311 (N_2311,N_1997,N_1962);
nor U2312 (N_2312,N_1679,N_1999);
and U2313 (N_2313,N_1696,N_1882);
and U2314 (N_2314,N_1819,N_1830);
nand U2315 (N_2315,N_1934,N_1618);
nor U2316 (N_2316,N_1739,N_1528);
or U2317 (N_2317,N_1841,N_1968);
and U2318 (N_2318,N_1614,N_1870);
or U2319 (N_2319,N_1878,N_1580);
nand U2320 (N_2320,N_1546,N_1746);
or U2321 (N_2321,N_1546,N_1667);
nor U2322 (N_2322,N_1718,N_1595);
or U2323 (N_2323,N_1998,N_1938);
nor U2324 (N_2324,N_1570,N_1566);
nand U2325 (N_2325,N_1706,N_1997);
nand U2326 (N_2326,N_1554,N_1958);
or U2327 (N_2327,N_1682,N_1942);
nand U2328 (N_2328,N_1832,N_1997);
nand U2329 (N_2329,N_1671,N_1669);
nand U2330 (N_2330,N_1883,N_1541);
and U2331 (N_2331,N_1863,N_1717);
or U2332 (N_2332,N_1541,N_1855);
and U2333 (N_2333,N_1751,N_1852);
xor U2334 (N_2334,N_1683,N_1956);
nand U2335 (N_2335,N_1844,N_1646);
nor U2336 (N_2336,N_1561,N_1713);
nand U2337 (N_2337,N_1827,N_1524);
nand U2338 (N_2338,N_1731,N_1523);
xor U2339 (N_2339,N_1699,N_1537);
nor U2340 (N_2340,N_1782,N_1703);
nand U2341 (N_2341,N_1687,N_1889);
or U2342 (N_2342,N_1713,N_1788);
nand U2343 (N_2343,N_1537,N_1866);
nand U2344 (N_2344,N_1903,N_1766);
nand U2345 (N_2345,N_1665,N_1688);
or U2346 (N_2346,N_1907,N_1564);
xor U2347 (N_2347,N_1727,N_1710);
and U2348 (N_2348,N_1928,N_1734);
nor U2349 (N_2349,N_1526,N_1876);
or U2350 (N_2350,N_1975,N_1874);
xor U2351 (N_2351,N_1763,N_1982);
or U2352 (N_2352,N_1560,N_1510);
nand U2353 (N_2353,N_1787,N_1686);
or U2354 (N_2354,N_1755,N_1996);
xor U2355 (N_2355,N_1824,N_1582);
nor U2356 (N_2356,N_1584,N_1882);
and U2357 (N_2357,N_1888,N_1516);
nand U2358 (N_2358,N_1551,N_1790);
and U2359 (N_2359,N_1741,N_1533);
or U2360 (N_2360,N_1903,N_1512);
xnor U2361 (N_2361,N_1876,N_1566);
and U2362 (N_2362,N_1616,N_1564);
and U2363 (N_2363,N_1596,N_1795);
or U2364 (N_2364,N_1546,N_1914);
or U2365 (N_2365,N_1554,N_1568);
and U2366 (N_2366,N_1912,N_1910);
and U2367 (N_2367,N_1859,N_1555);
or U2368 (N_2368,N_1700,N_1881);
xnor U2369 (N_2369,N_1843,N_1990);
nand U2370 (N_2370,N_1712,N_1610);
nor U2371 (N_2371,N_1823,N_1576);
nor U2372 (N_2372,N_1809,N_1576);
xor U2373 (N_2373,N_1696,N_1642);
or U2374 (N_2374,N_1545,N_1888);
and U2375 (N_2375,N_1842,N_1759);
or U2376 (N_2376,N_1851,N_1728);
nor U2377 (N_2377,N_1550,N_1990);
nand U2378 (N_2378,N_1638,N_1650);
xor U2379 (N_2379,N_1960,N_1620);
or U2380 (N_2380,N_1892,N_1762);
nor U2381 (N_2381,N_1617,N_1904);
nand U2382 (N_2382,N_1756,N_1940);
and U2383 (N_2383,N_1598,N_1701);
nand U2384 (N_2384,N_1839,N_1982);
nand U2385 (N_2385,N_1813,N_1565);
nor U2386 (N_2386,N_1724,N_1911);
or U2387 (N_2387,N_1701,N_1765);
and U2388 (N_2388,N_1683,N_1560);
or U2389 (N_2389,N_1687,N_1964);
or U2390 (N_2390,N_1999,N_1839);
nor U2391 (N_2391,N_1777,N_1844);
and U2392 (N_2392,N_1623,N_1964);
or U2393 (N_2393,N_1639,N_1860);
xnor U2394 (N_2394,N_1988,N_1834);
nor U2395 (N_2395,N_1717,N_1803);
and U2396 (N_2396,N_1913,N_1606);
nand U2397 (N_2397,N_1647,N_1507);
nor U2398 (N_2398,N_1681,N_1838);
xor U2399 (N_2399,N_1813,N_1946);
nor U2400 (N_2400,N_1605,N_1718);
or U2401 (N_2401,N_1678,N_1749);
or U2402 (N_2402,N_1950,N_1856);
or U2403 (N_2403,N_1703,N_1610);
nand U2404 (N_2404,N_1536,N_1582);
and U2405 (N_2405,N_1981,N_1562);
nand U2406 (N_2406,N_1575,N_1774);
and U2407 (N_2407,N_1911,N_1780);
and U2408 (N_2408,N_1658,N_1582);
nor U2409 (N_2409,N_1966,N_1910);
or U2410 (N_2410,N_1719,N_1902);
or U2411 (N_2411,N_1525,N_1950);
nor U2412 (N_2412,N_1912,N_1652);
nor U2413 (N_2413,N_1778,N_1688);
or U2414 (N_2414,N_1882,N_1689);
nand U2415 (N_2415,N_1760,N_1938);
nand U2416 (N_2416,N_1668,N_1550);
and U2417 (N_2417,N_1916,N_1564);
or U2418 (N_2418,N_1635,N_1664);
or U2419 (N_2419,N_1822,N_1774);
and U2420 (N_2420,N_1840,N_1809);
and U2421 (N_2421,N_1678,N_1577);
nand U2422 (N_2422,N_1706,N_1919);
nor U2423 (N_2423,N_1755,N_1915);
nor U2424 (N_2424,N_1651,N_1585);
or U2425 (N_2425,N_1917,N_1977);
and U2426 (N_2426,N_1828,N_1749);
nand U2427 (N_2427,N_1986,N_1547);
and U2428 (N_2428,N_1598,N_1506);
nor U2429 (N_2429,N_1890,N_1972);
nor U2430 (N_2430,N_1823,N_1904);
or U2431 (N_2431,N_1811,N_1713);
or U2432 (N_2432,N_1640,N_1564);
and U2433 (N_2433,N_1979,N_1846);
nand U2434 (N_2434,N_1920,N_1701);
xor U2435 (N_2435,N_1631,N_1859);
or U2436 (N_2436,N_1558,N_1999);
and U2437 (N_2437,N_1776,N_1841);
nor U2438 (N_2438,N_1519,N_1961);
nor U2439 (N_2439,N_1602,N_1749);
xor U2440 (N_2440,N_1609,N_1954);
or U2441 (N_2441,N_1826,N_1967);
xnor U2442 (N_2442,N_1630,N_1985);
nand U2443 (N_2443,N_1544,N_1659);
nor U2444 (N_2444,N_1808,N_1757);
nand U2445 (N_2445,N_1742,N_1760);
xor U2446 (N_2446,N_1615,N_1663);
and U2447 (N_2447,N_1862,N_1914);
nor U2448 (N_2448,N_1598,N_1758);
nand U2449 (N_2449,N_1726,N_1851);
or U2450 (N_2450,N_1703,N_1768);
xor U2451 (N_2451,N_1955,N_1796);
or U2452 (N_2452,N_1734,N_1729);
nand U2453 (N_2453,N_1510,N_1620);
nor U2454 (N_2454,N_1663,N_1803);
and U2455 (N_2455,N_1661,N_1993);
or U2456 (N_2456,N_1677,N_1896);
nand U2457 (N_2457,N_1606,N_1620);
nor U2458 (N_2458,N_1692,N_1848);
xor U2459 (N_2459,N_1686,N_1699);
nand U2460 (N_2460,N_1957,N_1950);
and U2461 (N_2461,N_1892,N_1534);
and U2462 (N_2462,N_1950,N_1887);
nand U2463 (N_2463,N_1906,N_1546);
xnor U2464 (N_2464,N_1879,N_1646);
nor U2465 (N_2465,N_1663,N_1716);
or U2466 (N_2466,N_1972,N_1792);
or U2467 (N_2467,N_1656,N_1886);
nand U2468 (N_2468,N_1912,N_1518);
or U2469 (N_2469,N_1709,N_1774);
nand U2470 (N_2470,N_1939,N_1640);
nor U2471 (N_2471,N_1998,N_1571);
xor U2472 (N_2472,N_1755,N_1939);
and U2473 (N_2473,N_1612,N_1717);
or U2474 (N_2474,N_1814,N_1908);
nor U2475 (N_2475,N_1719,N_1908);
nand U2476 (N_2476,N_1665,N_1941);
nor U2477 (N_2477,N_1818,N_1806);
or U2478 (N_2478,N_1842,N_1735);
or U2479 (N_2479,N_1585,N_1822);
and U2480 (N_2480,N_1855,N_1522);
or U2481 (N_2481,N_1695,N_1533);
or U2482 (N_2482,N_1823,N_1637);
nor U2483 (N_2483,N_1662,N_1591);
and U2484 (N_2484,N_1880,N_1641);
nand U2485 (N_2485,N_1746,N_1889);
nor U2486 (N_2486,N_1620,N_1987);
or U2487 (N_2487,N_1626,N_1845);
nand U2488 (N_2488,N_1778,N_1630);
and U2489 (N_2489,N_1970,N_1853);
nor U2490 (N_2490,N_1754,N_1588);
nand U2491 (N_2491,N_1522,N_1566);
or U2492 (N_2492,N_1624,N_1914);
nor U2493 (N_2493,N_1884,N_1825);
or U2494 (N_2494,N_1584,N_1906);
or U2495 (N_2495,N_1916,N_1947);
and U2496 (N_2496,N_1753,N_1850);
nor U2497 (N_2497,N_1681,N_1816);
and U2498 (N_2498,N_1590,N_1533);
nand U2499 (N_2499,N_1737,N_1526);
nor U2500 (N_2500,N_2056,N_2266);
nor U2501 (N_2501,N_2111,N_2413);
nand U2502 (N_2502,N_2408,N_2343);
nor U2503 (N_2503,N_2020,N_2189);
nor U2504 (N_2504,N_2326,N_2317);
nand U2505 (N_2505,N_2180,N_2361);
and U2506 (N_2506,N_2208,N_2392);
and U2507 (N_2507,N_2109,N_2076);
or U2508 (N_2508,N_2384,N_2337);
nand U2509 (N_2509,N_2154,N_2456);
nand U2510 (N_2510,N_2077,N_2254);
nor U2511 (N_2511,N_2146,N_2350);
or U2512 (N_2512,N_2386,N_2393);
nor U2513 (N_2513,N_2289,N_2410);
and U2514 (N_2514,N_2140,N_2046);
nand U2515 (N_2515,N_2333,N_2259);
or U2516 (N_2516,N_2043,N_2421);
nor U2517 (N_2517,N_2198,N_2472);
or U2518 (N_2518,N_2000,N_2011);
nor U2519 (N_2519,N_2003,N_2340);
xnor U2520 (N_2520,N_2390,N_2196);
nand U2521 (N_2521,N_2192,N_2462);
nand U2522 (N_2522,N_2325,N_2296);
nand U2523 (N_2523,N_2488,N_2074);
nor U2524 (N_2524,N_2226,N_2403);
nand U2525 (N_2525,N_2485,N_2396);
nand U2526 (N_2526,N_2080,N_2092);
or U2527 (N_2527,N_2032,N_2318);
nor U2528 (N_2528,N_2104,N_2084);
nand U2529 (N_2529,N_2257,N_2021);
nor U2530 (N_2530,N_2299,N_2121);
nand U2531 (N_2531,N_2187,N_2212);
and U2532 (N_2532,N_2055,N_2108);
nor U2533 (N_2533,N_2057,N_2453);
nand U2534 (N_2534,N_2238,N_2063);
xor U2535 (N_2535,N_2124,N_2490);
nand U2536 (N_2536,N_2136,N_2079);
or U2537 (N_2537,N_2006,N_2487);
nand U2538 (N_2538,N_2151,N_2245);
or U2539 (N_2539,N_2068,N_2400);
nand U2540 (N_2540,N_2036,N_2088);
or U2541 (N_2541,N_2090,N_2031);
or U2542 (N_2542,N_2148,N_2481);
nor U2543 (N_2543,N_2066,N_2041);
or U2544 (N_2544,N_2191,N_2203);
and U2545 (N_2545,N_2402,N_2370);
or U2546 (N_2546,N_2336,N_2139);
nand U2547 (N_2547,N_2160,N_2356);
nor U2548 (N_2548,N_2280,N_2156);
nor U2549 (N_2549,N_2119,N_2070);
xnor U2550 (N_2550,N_2310,N_2166);
nor U2551 (N_2551,N_2051,N_2422);
nor U2552 (N_2552,N_2125,N_2425);
nor U2553 (N_2553,N_2012,N_2093);
nor U2554 (N_2554,N_2072,N_2123);
nand U2555 (N_2555,N_2405,N_2428);
nand U2556 (N_2556,N_2364,N_2232);
nand U2557 (N_2557,N_2231,N_2237);
nand U2558 (N_2558,N_2253,N_2323);
xnor U2559 (N_2559,N_2330,N_2352);
nor U2560 (N_2560,N_2186,N_2368);
nand U2561 (N_2561,N_2258,N_2168);
or U2562 (N_2562,N_2223,N_2439);
nand U2563 (N_2563,N_2301,N_2214);
nand U2564 (N_2564,N_2058,N_2346);
and U2565 (N_2565,N_2242,N_2349);
nor U2566 (N_2566,N_2217,N_2022);
nand U2567 (N_2567,N_2159,N_2277);
nor U2568 (N_2568,N_2427,N_2061);
nor U2569 (N_2569,N_2401,N_2300);
nor U2570 (N_2570,N_2222,N_2050);
and U2571 (N_2571,N_2177,N_2086);
or U2572 (N_2572,N_2447,N_2412);
xor U2573 (N_2573,N_2024,N_2312);
nand U2574 (N_2574,N_2335,N_2047);
and U2575 (N_2575,N_2465,N_2145);
or U2576 (N_2576,N_2004,N_2176);
nor U2577 (N_2577,N_2175,N_2045);
nor U2578 (N_2578,N_2389,N_2482);
or U2579 (N_2579,N_2426,N_2397);
xnor U2580 (N_2580,N_2193,N_2302);
nor U2581 (N_2581,N_2309,N_2010);
nor U2582 (N_2582,N_2044,N_2415);
xor U2583 (N_2583,N_2001,N_2244);
or U2584 (N_2584,N_2452,N_2054);
or U2585 (N_2585,N_2429,N_2339);
nor U2586 (N_2586,N_2144,N_2475);
and U2587 (N_2587,N_2264,N_2195);
or U2588 (N_2588,N_2181,N_2105);
and U2589 (N_2589,N_2272,N_2229);
and U2590 (N_2590,N_2313,N_2486);
nor U2591 (N_2591,N_2423,N_2081);
or U2592 (N_2592,N_2286,N_2157);
and U2593 (N_2593,N_2455,N_2027);
nand U2594 (N_2594,N_2069,N_2362);
and U2595 (N_2595,N_2469,N_2457);
nand U2596 (N_2596,N_2210,N_2284);
and U2597 (N_2597,N_2150,N_2329);
or U2598 (N_2598,N_2221,N_2274);
and U2599 (N_2599,N_2129,N_2184);
nand U2600 (N_2600,N_2252,N_2363);
xor U2601 (N_2601,N_2378,N_2407);
nand U2602 (N_2602,N_2211,N_2065);
or U2603 (N_2603,N_2225,N_2170);
and U2604 (N_2604,N_2357,N_2243);
nand U2605 (N_2605,N_2134,N_2255);
or U2606 (N_2606,N_2265,N_2479);
nor U2607 (N_2607,N_2048,N_2089);
or U2608 (N_2608,N_2260,N_2230);
nand U2609 (N_2609,N_2461,N_2030);
or U2610 (N_2610,N_2449,N_2083);
nand U2611 (N_2611,N_2498,N_2248);
nand U2612 (N_2612,N_2307,N_2158);
nor U2613 (N_2613,N_2443,N_2279);
and U2614 (N_2614,N_2276,N_2122);
nand U2615 (N_2615,N_2322,N_2354);
nand U2616 (N_2616,N_2269,N_2023);
and U2617 (N_2617,N_2082,N_2328);
and U2618 (N_2618,N_2493,N_2239);
nor U2619 (N_2619,N_2434,N_2314);
nor U2620 (N_2620,N_2064,N_2446);
nand U2621 (N_2621,N_2102,N_2440);
nand U2622 (N_2622,N_2360,N_2009);
or U2623 (N_2623,N_2233,N_2353);
or U2624 (N_2624,N_2411,N_2261);
nand U2625 (N_2625,N_2141,N_2182);
and U2626 (N_2626,N_2463,N_2101);
or U2627 (N_2627,N_2120,N_2473);
nor U2628 (N_2628,N_2404,N_2297);
nor U2629 (N_2629,N_2178,N_2110);
and U2630 (N_2630,N_2251,N_2497);
nor U2631 (N_2631,N_2075,N_2127);
nor U2632 (N_2632,N_2394,N_2118);
nor U2633 (N_2633,N_2294,N_2137);
and U2634 (N_2634,N_2435,N_2438);
or U2635 (N_2635,N_2149,N_2372);
xnor U2636 (N_2636,N_2142,N_2477);
nand U2637 (N_2637,N_2355,N_2320);
or U2638 (N_2638,N_2291,N_2365);
nand U2639 (N_2639,N_2098,N_2096);
and U2640 (N_2640,N_2053,N_2085);
nand U2641 (N_2641,N_2029,N_2037);
xnor U2642 (N_2642,N_2433,N_2062);
and U2643 (N_2643,N_2117,N_2132);
and U2644 (N_2644,N_2256,N_2067);
or U2645 (N_2645,N_2460,N_2419);
xnor U2646 (N_2646,N_2420,N_2334);
nor U2647 (N_2647,N_2155,N_2444);
nor U2648 (N_2648,N_2327,N_2113);
nand U2649 (N_2649,N_2162,N_2483);
xor U2650 (N_2650,N_2344,N_2321);
nor U2651 (N_2651,N_2234,N_2342);
nor U2652 (N_2652,N_2017,N_2052);
nor U2653 (N_2653,N_2116,N_2227);
nor U2654 (N_2654,N_2106,N_2441);
and U2655 (N_2655,N_2138,N_2263);
nor U2656 (N_2656,N_2199,N_2437);
nand U2657 (N_2657,N_2188,N_2078);
or U2658 (N_2658,N_2247,N_2167);
and U2659 (N_2659,N_2095,N_2375);
or U2660 (N_2660,N_2163,N_2060);
and U2661 (N_2661,N_2492,N_2406);
or U2662 (N_2662,N_2305,N_2262);
and U2663 (N_2663,N_2015,N_2218);
or U2664 (N_2664,N_2224,N_2351);
or U2665 (N_2665,N_2107,N_2450);
xnor U2666 (N_2666,N_2275,N_2039);
and U2667 (N_2667,N_2002,N_2374);
xnor U2668 (N_2668,N_2376,N_2358);
xnor U2669 (N_2669,N_2097,N_2236);
xor U2670 (N_2670,N_2290,N_2209);
xnor U2671 (N_2671,N_2112,N_2018);
or U2672 (N_2672,N_2100,N_2197);
xor U2673 (N_2673,N_2311,N_2319);
nand U2674 (N_2674,N_2282,N_2431);
or U2675 (N_2675,N_2215,N_2071);
nor U2676 (N_2676,N_2174,N_2474);
or U2677 (N_2677,N_2202,N_2073);
or U2678 (N_2678,N_2103,N_2040);
or U2679 (N_2679,N_2331,N_2359);
and U2680 (N_2680,N_2172,N_2033);
nor U2681 (N_2681,N_2216,N_2267);
nand U2682 (N_2682,N_2417,N_2458);
xor U2683 (N_2683,N_2087,N_2049);
nor U2684 (N_2684,N_2194,N_2005);
nand U2685 (N_2685,N_2304,N_2213);
nand U2686 (N_2686,N_2464,N_2173);
nor U2687 (N_2687,N_2026,N_2204);
nand U2688 (N_2688,N_2185,N_2496);
or U2689 (N_2689,N_2383,N_2271);
nor U2690 (N_2690,N_2367,N_2007);
nand U2691 (N_2691,N_2377,N_2008);
xor U2692 (N_2692,N_2130,N_2016);
xnor U2693 (N_2693,N_2347,N_2099);
or U2694 (N_2694,N_2494,N_2432);
nand U2695 (N_2695,N_2179,N_2468);
xor U2696 (N_2696,N_2143,N_2228);
or U2697 (N_2697,N_2476,N_2345);
xor U2698 (N_2698,N_2380,N_2306);
or U2699 (N_2699,N_2038,N_2391);
nand U2700 (N_2700,N_2281,N_2385);
nand U2701 (N_2701,N_2341,N_2489);
nand U2702 (N_2702,N_2287,N_2424);
or U2703 (N_2703,N_2094,N_2398);
xor U2704 (N_2704,N_2324,N_2495);
nand U2705 (N_2705,N_2366,N_2442);
nor U2706 (N_2706,N_2133,N_2241);
xor U2707 (N_2707,N_2152,N_2268);
or U2708 (N_2708,N_2164,N_2219);
and U2709 (N_2709,N_2035,N_2308);
and U2710 (N_2710,N_2165,N_2387);
xnor U2711 (N_2711,N_2348,N_2315);
xnor U2712 (N_2712,N_2207,N_2491);
nor U2713 (N_2713,N_2201,N_2034);
xnor U2714 (N_2714,N_2459,N_2478);
nand U2715 (N_2715,N_2028,N_2014);
and U2716 (N_2716,N_2042,N_2338);
or U2717 (N_2717,N_2013,N_2153);
nor U2718 (N_2718,N_2295,N_2471);
or U2719 (N_2719,N_2270,N_2115);
nor U2720 (N_2720,N_2249,N_2169);
nand U2721 (N_2721,N_2273,N_2147);
nand U2722 (N_2722,N_2126,N_2235);
xor U2723 (N_2723,N_2220,N_2131);
nand U2724 (N_2724,N_2332,N_2409);
nand U2725 (N_2725,N_2448,N_2399);
nor U2726 (N_2726,N_2288,N_2388);
xnor U2727 (N_2727,N_2484,N_2128);
and U2728 (N_2728,N_2206,N_2395);
nand U2729 (N_2729,N_2454,N_2298);
xnor U2730 (N_2730,N_2416,N_2293);
and U2731 (N_2731,N_2161,N_2467);
nand U2732 (N_2732,N_2240,N_2499);
or U2733 (N_2733,N_2025,N_2285);
nor U2734 (N_2734,N_2114,N_2445);
nand U2735 (N_2735,N_2414,N_2059);
or U2736 (N_2736,N_2470,N_2278);
xor U2737 (N_2737,N_2373,N_2381);
nor U2738 (N_2738,N_2466,N_2418);
nand U2739 (N_2739,N_2379,N_2250);
nand U2740 (N_2740,N_2200,N_2430);
or U2741 (N_2741,N_2190,N_2436);
and U2742 (N_2742,N_2246,N_2135);
or U2743 (N_2743,N_2480,N_2183);
nor U2744 (N_2744,N_2292,N_2371);
or U2745 (N_2745,N_2091,N_2451);
nand U2746 (N_2746,N_2382,N_2369);
nor U2747 (N_2747,N_2205,N_2303);
xnor U2748 (N_2748,N_2019,N_2171);
nand U2749 (N_2749,N_2283,N_2316);
and U2750 (N_2750,N_2112,N_2331);
nand U2751 (N_2751,N_2368,N_2374);
and U2752 (N_2752,N_2075,N_2141);
and U2753 (N_2753,N_2091,N_2015);
nor U2754 (N_2754,N_2354,N_2038);
nand U2755 (N_2755,N_2274,N_2231);
xor U2756 (N_2756,N_2116,N_2124);
and U2757 (N_2757,N_2017,N_2152);
nor U2758 (N_2758,N_2330,N_2423);
nand U2759 (N_2759,N_2333,N_2343);
nor U2760 (N_2760,N_2341,N_2176);
or U2761 (N_2761,N_2082,N_2150);
nor U2762 (N_2762,N_2320,N_2297);
nor U2763 (N_2763,N_2439,N_2084);
or U2764 (N_2764,N_2413,N_2361);
nand U2765 (N_2765,N_2490,N_2323);
and U2766 (N_2766,N_2125,N_2097);
nand U2767 (N_2767,N_2002,N_2193);
or U2768 (N_2768,N_2159,N_2424);
nand U2769 (N_2769,N_2380,N_2126);
nor U2770 (N_2770,N_2398,N_2081);
and U2771 (N_2771,N_2325,N_2059);
xor U2772 (N_2772,N_2367,N_2362);
xor U2773 (N_2773,N_2127,N_2407);
nor U2774 (N_2774,N_2476,N_2479);
xnor U2775 (N_2775,N_2005,N_2140);
nor U2776 (N_2776,N_2055,N_2017);
or U2777 (N_2777,N_2426,N_2095);
nand U2778 (N_2778,N_2120,N_2470);
nor U2779 (N_2779,N_2280,N_2057);
nand U2780 (N_2780,N_2369,N_2373);
and U2781 (N_2781,N_2221,N_2289);
nand U2782 (N_2782,N_2020,N_2110);
and U2783 (N_2783,N_2298,N_2198);
xor U2784 (N_2784,N_2115,N_2148);
nor U2785 (N_2785,N_2415,N_2358);
or U2786 (N_2786,N_2171,N_2120);
nand U2787 (N_2787,N_2251,N_2105);
nor U2788 (N_2788,N_2141,N_2274);
or U2789 (N_2789,N_2141,N_2203);
and U2790 (N_2790,N_2408,N_2411);
xnor U2791 (N_2791,N_2330,N_2191);
and U2792 (N_2792,N_2280,N_2240);
xnor U2793 (N_2793,N_2354,N_2193);
and U2794 (N_2794,N_2208,N_2431);
or U2795 (N_2795,N_2171,N_2352);
and U2796 (N_2796,N_2360,N_2474);
nor U2797 (N_2797,N_2231,N_2497);
or U2798 (N_2798,N_2219,N_2276);
nor U2799 (N_2799,N_2408,N_2382);
nor U2800 (N_2800,N_2406,N_2307);
nor U2801 (N_2801,N_2183,N_2485);
and U2802 (N_2802,N_2294,N_2014);
or U2803 (N_2803,N_2192,N_2342);
or U2804 (N_2804,N_2374,N_2460);
nand U2805 (N_2805,N_2163,N_2082);
and U2806 (N_2806,N_2094,N_2401);
nand U2807 (N_2807,N_2074,N_2146);
nand U2808 (N_2808,N_2184,N_2183);
nor U2809 (N_2809,N_2129,N_2422);
and U2810 (N_2810,N_2339,N_2127);
or U2811 (N_2811,N_2191,N_2178);
nand U2812 (N_2812,N_2096,N_2361);
or U2813 (N_2813,N_2297,N_2499);
or U2814 (N_2814,N_2433,N_2124);
xor U2815 (N_2815,N_2326,N_2168);
nor U2816 (N_2816,N_2301,N_2485);
or U2817 (N_2817,N_2062,N_2415);
or U2818 (N_2818,N_2330,N_2136);
nand U2819 (N_2819,N_2436,N_2475);
and U2820 (N_2820,N_2266,N_2474);
and U2821 (N_2821,N_2066,N_2391);
or U2822 (N_2822,N_2033,N_2495);
nor U2823 (N_2823,N_2416,N_2486);
nand U2824 (N_2824,N_2443,N_2465);
nand U2825 (N_2825,N_2315,N_2377);
or U2826 (N_2826,N_2404,N_2335);
or U2827 (N_2827,N_2126,N_2433);
and U2828 (N_2828,N_2396,N_2112);
nor U2829 (N_2829,N_2336,N_2064);
and U2830 (N_2830,N_2134,N_2403);
nor U2831 (N_2831,N_2209,N_2258);
nand U2832 (N_2832,N_2069,N_2434);
and U2833 (N_2833,N_2295,N_2204);
nor U2834 (N_2834,N_2068,N_2115);
xor U2835 (N_2835,N_2231,N_2005);
and U2836 (N_2836,N_2487,N_2079);
xnor U2837 (N_2837,N_2388,N_2465);
nand U2838 (N_2838,N_2063,N_2415);
and U2839 (N_2839,N_2389,N_2291);
and U2840 (N_2840,N_2481,N_2156);
or U2841 (N_2841,N_2010,N_2234);
nor U2842 (N_2842,N_2307,N_2290);
and U2843 (N_2843,N_2325,N_2493);
nand U2844 (N_2844,N_2272,N_2176);
or U2845 (N_2845,N_2333,N_2065);
or U2846 (N_2846,N_2139,N_2340);
nor U2847 (N_2847,N_2293,N_2410);
nor U2848 (N_2848,N_2401,N_2354);
nor U2849 (N_2849,N_2111,N_2225);
and U2850 (N_2850,N_2165,N_2404);
nand U2851 (N_2851,N_2130,N_2070);
and U2852 (N_2852,N_2305,N_2302);
nand U2853 (N_2853,N_2091,N_2089);
and U2854 (N_2854,N_2312,N_2125);
or U2855 (N_2855,N_2016,N_2304);
or U2856 (N_2856,N_2431,N_2097);
and U2857 (N_2857,N_2388,N_2190);
or U2858 (N_2858,N_2311,N_2483);
nor U2859 (N_2859,N_2042,N_2452);
xor U2860 (N_2860,N_2041,N_2274);
or U2861 (N_2861,N_2081,N_2126);
nor U2862 (N_2862,N_2361,N_2166);
and U2863 (N_2863,N_2499,N_2123);
nand U2864 (N_2864,N_2273,N_2170);
or U2865 (N_2865,N_2219,N_2455);
nor U2866 (N_2866,N_2059,N_2301);
nand U2867 (N_2867,N_2172,N_2472);
or U2868 (N_2868,N_2273,N_2470);
nand U2869 (N_2869,N_2387,N_2442);
and U2870 (N_2870,N_2346,N_2052);
and U2871 (N_2871,N_2335,N_2393);
and U2872 (N_2872,N_2360,N_2250);
or U2873 (N_2873,N_2410,N_2489);
nor U2874 (N_2874,N_2195,N_2394);
nor U2875 (N_2875,N_2146,N_2452);
and U2876 (N_2876,N_2084,N_2494);
or U2877 (N_2877,N_2432,N_2447);
or U2878 (N_2878,N_2283,N_2308);
nand U2879 (N_2879,N_2335,N_2100);
nand U2880 (N_2880,N_2256,N_2473);
nor U2881 (N_2881,N_2403,N_2384);
nand U2882 (N_2882,N_2406,N_2236);
xnor U2883 (N_2883,N_2271,N_2209);
and U2884 (N_2884,N_2405,N_2231);
nand U2885 (N_2885,N_2144,N_2087);
and U2886 (N_2886,N_2303,N_2083);
nor U2887 (N_2887,N_2135,N_2305);
and U2888 (N_2888,N_2016,N_2385);
or U2889 (N_2889,N_2451,N_2316);
and U2890 (N_2890,N_2465,N_2304);
nor U2891 (N_2891,N_2296,N_2499);
nor U2892 (N_2892,N_2253,N_2057);
or U2893 (N_2893,N_2416,N_2362);
nand U2894 (N_2894,N_2388,N_2137);
nand U2895 (N_2895,N_2440,N_2088);
and U2896 (N_2896,N_2490,N_2368);
xnor U2897 (N_2897,N_2498,N_2466);
and U2898 (N_2898,N_2476,N_2414);
nand U2899 (N_2899,N_2178,N_2183);
nor U2900 (N_2900,N_2324,N_2052);
or U2901 (N_2901,N_2232,N_2152);
or U2902 (N_2902,N_2185,N_2429);
nor U2903 (N_2903,N_2194,N_2088);
nor U2904 (N_2904,N_2256,N_2046);
nor U2905 (N_2905,N_2324,N_2155);
and U2906 (N_2906,N_2445,N_2058);
or U2907 (N_2907,N_2376,N_2244);
xnor U2908 (N_2908,N_2154,N_2314);
xor U2909 (N_2909,N_2289,N_2048);
or U2910 (N_2910,N_2104,N_2463);
nand U2911 (N_2911,N_2081,N_2025);
nor U2912 (N_2912,N_2108,N_2021);
and U2913 (N_2913,N_2177,N_2435);
nor U2914 (N_2914,N_2477,N_2331);
and U2915 (N_2915,N_2434,N_2494);
xor U2916 (N_2916,N_2476,N_2122);
nor U2917 (N_2917,N_2365,N_2438);
and U2918 (N_2918,N_2162,N_2206);
and U2919 (N_2919,N_2069,N_2302);
and U2920 (N_2920,N_2029,N_2441);
nand U2921 (N_2921,N_2379,N_2322);
and U2922 (N_2922,N_2225,N_2231);
nand U2923 (N_2923,N_2444,N_2325);
nand U2924 (N_2924,N_2003,N_2392);
or U2925 (N_2925,N_2068,N_2138);
nand U2926 (N_2926,N_2205,N_2329);
and U2927 (N_2927,N_2221,N_2426);
nor U2928 (N_2928,N_2489,N_2085);
and U2929 (N_2929,N_2322,N_2232);
nor U2930 (N_2930,N_2161,N_2445);
and U2931 (N_2931,N_2242,N_2475);
xor U2932 (N_2932,N_2003,N_2261);
nor U2933 (N_2933,N_2422,N_2181);
nor U2934 (N_2934,N_2135,N_2459);
or U2935 (N_2935,N_2067,N_2071);
and U2936 (N_2936,N_2381,N_2403);
and U2937 (N_2937,N_2312,N_2009);
nor U2938 (N_2938,N_2012,N_2257);
and U2939 (N_2939,N_2370,N_2457);
or U2940 (N_2940,N_2182,N_2078);
nor U2941 (N_2941,N_2363,N_2303);
xnor U2942 (N_2942,N_2024,N_2244);
and U2943 (N_2943,N_2320,N_2123);
or U2944 (N_2944,N_2305,N_2006);
or U2945 (N_2945,N_2047,N_2212);
nand U2946 (N_2946,N_2425,N_2377);
nor U2947 (N_2947,N_2173,N_2136);
or U2948 (N_2948,N_2161,N_2237);
and U2949 (N_2949,N_2412,N_2391);
nor U2950 (N_2950,N_2098,N_2058);
nand U2951 (N_2951,N_2323,N_2462);
nand U2952 (N_2952,N_2237,N_2305);
or U2953 (N_2953,N_2068,N_2495);
or U2954 (N_2954,N_2279,N_2257);
and U2955 (N_2955,N_2481,N_2033);
nand U2956 (N_2956,N_2434,N_2473);
and U2957 (N_2957,N_2407,N_2006);
nand U2958 (N_2958,N_2232,N_2154);
xor U2959 (N_2959,N_2185,N_2107);
nor U2960 (N_2960,N_2093,N_2240);
nor U2961 (N_2961,N_2237,N_2306);
or U2962 (N_2962,N_2159,N_2019);
and U2963 (N_2963,N_2239,N_2171);
and U2964 (N_2964,N_2194,N_2198);
xnor U2965 (N_2965,N_2273,N_2220);
nand U2966 (N_2966,N_2299,N_2066);
or U2967 (N_2967,N_2141,N_2052);
or U2968 (N_2968,N_2358,N_2163);
and U2969 (N_2969,N_2181,N_2433);
nand U2970 (N_2970,N_2161,N_2129);
nand U2971 (N_2971,N_2243,N_2285);
and U2972 (N_2972,N_2175,N_2386);
xor U2973 (N_2973,N_2413,N_2141);
or U2974 (N_2974,N_2370,N_2036);
nor U2975 (N_2975,N_2051,N_2328);
nor U2976 (N_2976,N_2077,N_2159);
nand U2977 (N_2977,N_2102,N_2407);
nor U2978 (N_2978,N_2383,N_2267);
nand U2979 (N_2979,N_2423,N_2055);
and U2980 (N_2980,N_2233,N_2122);
nor U2981 (N_2981,N_2374,N_2324);
xor U2982 (N_2982,N_2011,N_2027);
and U2983 (N_2983,N_2034,N_2204);
nand U2984 (N_2984,N_2278,N_2039);
or U2985 (N_2985,N_2102,N_2141);
nor U2986 (N_2986,N_2054,N_2438);
nor U2987 (N_2987,N_2162,N_2419);
and U2988 (N_2988,N_2112,N_2229);
or U2989 (N_2989,N_2198,N_2457);
and U2990 (N_2990,N_2226,N_2395);
and U2991 (N_2991,N_2163,N_2365);
or U2992 (N_2992,N_2236,N_2317);
nand U2993 (N_2993,N_2453,N_2132);
xor U2994 (N_2994,N_2323,N_2027);
nand U2995 (N_2995,N_2465,N_2180);
or U2996 (N_2996,N_2190,N_2290);
nor U2997 (N_2997,N_2333,N_2384);
xnor U2998 (N_2998,N_2282,N_2353);
and U2999 (N_2999,N_2062,N_2191);
xnor UO_0 (O_0,N_2535,N_2935);
nand UO_1 (O_1,N_2528,N_2986);
or UO_2 (O_2,N_2878,N_2712);
nor UO_3 (O_3,N_2888,N_2625);
nand UO_4 (O_4,N_2823,N_2575);
and UO_5 (O_5,N_2720,N_2862);
and UO_6 (O_6,N_2793,N_2969);
xnor UO_7 (O_7,N_2604,N_2874);
and UO_8 (O_8,N_2883,N_2928);
or UO_9 (O_9,N_2696,N_2879);
or UO_10 (O_10,N_2939,N_2880);
and UO_11 (O_11,N_2779,N_2988);
xnor UO_12 (O_12,N_2852,N_2724);
or UO_13 (O_13,N_2542,N_2867);
nor UO_14 (O_14,N_2964,N_2804);
or UO_15 (O_15,N_2552,N_2849);
and UO_16 (O_16,N_2923,N_2802);
and UO_17 (O_17,N_2978,N_2596);
xor UO_18 (O_18,N_2768,N_2548);
xnor UO_19 (O_19,N_2872,N_2967);
xor UO_20 (O_20,N_2798,N_2581);
xnor UO_21 (O_21,N_2844,N_2841);
xor UO_22 (O_22,N_2739,N_2685);
nor UO_23 (O_23,N_2819,N_2508);
or UO_24 (O_24,N_2714,N_2626);
xor UO_25 (O_25,N_2505,N_2646);
nor UO_26 (O_26,N_2837,N_2910);
or UO_27 (O_27,N_2507,N_2737);
nand UO_28 (O_28,N_2790,N_2827);
and UO_29 (O_29,N_2560,N_2527);
or UO_30 (O_30,N_2949,N_2977);
nand UO_31 (O_31,N_2567,N_2989);
and UO_32 (O_32,N_2759,N_2900);
and UO_33 (O_33,N_2886,N_2729);
or UO_34 (O_34,N_2840,N_2921);
nand UO_35 (O_35,N_2635,N_2856);
nor UO_36 (O_36,N_2601,N_2975);
nor UO_37 (O_37,N_2769,N_2589);
or UO_38 (O_38,N_2943,N_2621);
nand UO_39 (O_39,N_2632,N_2814);
nand UO_40 (O_40,N_2728,N_2937);
or UO_41 (O_41,N_2771,N_2733);
nor UO_42 (O_42,N_2584,N_2904);
nand UO_43 (O_43,N_2531,N_2898);
nor UO_44 (O_44,N_2922,N_2981);
and UO_45 (O_45,N_2812,N_2833);
and UO_46 (O_46,N_2640,N_2639);
nor UO_47 (O_47,N_2780,N_2829);
or UO_48 (O_48,N_2583,N_2607);
nor UO_49 (O_49,N_2866,N_2875);
nor UO_50 (O_50,N_2671,N_2645);
xor UO_51 (O_51,N_2563,N_2914);
nand UO_52 (O_52,N_2760,N_2927);
xor UO_53 (O_53,N_2553,N_2913);
or UO_54 (O_54,N_2711,N_2805);
nor UO_55 (O_55,N_2803,N_2847);
nand UO_56 (O_56,N_2579,N_2690);
and UO_57 (O_57,N_2620,N_2501);
and UO_58 (O_58,N_2722,N_2948);
nor UO_59 (O_59,N_2970,N_2545);
nor UO_60 (O_60,N_2952,N_2870);
and UO_61 (O_61,N_2695,N_2958);
or UO_62 (O_62,N_2945,N_2756);
or UO_63 (O_63,N_2821,N_2820);
and UO_64 (O_64,N_2515,N_2736);
and UO_65 (O_65,N_2555,N_2777);
or UO_66 (O_66,N_2594,N_2735);
nand UO_67 (O_67,N_2502,N_2938);
xnor UO_68 (O_68,N_2857,N_2854);
nand UO_69 (O_69,N_2745,N_2889);
and UO_70 (O_70,N_2773,N_2983);
nand UO_71 (O_71,N_2936,N_2905);
nor UO_72 (O_72,N_2623,N_2734);
and UO_73 (O_73,N_2959,N_2511);
nand UO_74 (O_74,N_2518,N_2656);
xnor UO_75 (O_75,N_2707,N_2687);
nand UO_76 (O_76,N_2573,N_2578);
nor UO_77 (O_77,N_2896,N_2658);
and UO_78 (O_78,N_2593,N_2895);
and UO_79 (O_79,N_2873,N_2860);
xnor UO_80 (O_80,N_2636,N_2950);
or UO_81 (O_81,N_2766,N_2911);
nand UO_82 (O_82,N_2562,N_2655);
xor UO_83 (O_83,N_2513,N_2679);
or UO_84 (O_84,N_2674,N_2569);
or UO_85 (O_85,N_2672,N_2686);
and UO_86 (O_86,N_2550,N_2549);
and UO_87 (O_87,N_2710,N_2525);
nor UO_88 (O_88,N_2908,N_2976);
xnor UO_89 (O_89,N_2912,N_2617);
nand UO_90 (O_90,N_2629,N_2524);
nand UO_91 (O_91,N_2526,N_2903);
nand UO_92 (O_92,N_2586,N_2846);
nor UO_93 (O_93,N_2761,N_2770);
and UO_94 (O_94,N_2561,N_2746);
and UO_95 (O_95,N_2916,N_2719);
nor UO_96 (O_96,N_2654,N_2996);
xnor UO_97 (O_97,N_2678,N_2708);
nor UO_98 (O_98,N_2638,N_2726);
nor UO_99 (O_99,N_2642,N_2539);
nor UO_100 (O_100,N_2801,N_2861);
nand UO_101 (O_101,N_2954,N_2644);
nor UO_102 (O_102,N_2884,N_2605);
or UO_103 (O_103,N_2772,N_2946);
xor UO_104 (O_104,N_2909,N_2570);
xor UO_105 (O_105,N_2876,N_2985);
and UO_106 (O_106,N_2919,N_2512);
xnor UO_107 (O_107,N_2509,N_2877);
nand UO_108 (O_108,N_2666,N_2659);
and UO_109 (O_109,N_2701,N_2557);
and UO_110 (O_110,N_2980,N_2715);
or UO_111 (O_111,N_2647,N_2891);
and UO_112 (O_112,N_2998,N_2500);
nor UO_113 (O_113,N_2706,N_2649);
nor UO_114 (O_114,N_2681,N_2554);
or UO_115 (O_115,N_2807,N_2982);
and UO_116 (O_116,N_2997,N_2758);
nor UO_117 (O_117,N_2546,N_2665);
nand UO_118 (O_118,N_2740,N_2999);
and UO_119 (O_119,N_2630,N_2944);
or UO_120 (O_120,N_2973,N_2587);
and UO_121 (O_121,N_2885,N_2754);
or UO_122 (O_122,N_2915,N_2755);
or UO_123 (O_123,N_2799,N_2520);
nand UO_124 (O_124,N_2816,N_2931);
or UO_125 (O_125,N_2574,N_2782);
or UO_126 (O_126,N_2848,N_2648);
or UO_127 (O_127,N_2951,N_2813);
xnor UO_128 (O_128,N_2956,N_2599);
nand UO_129 (O_129,N_2651,N_2942);
and UO_130 (O_130,N_2743,N_2811);
nor UO_131 (O_131,N_2634,N_2536);
nand UO_132 (O_132,N_2698,N_2716);
xor UO_133 (O_133,N_2519,N_2689);
nor UO_134 (O_134,N_2667,N_2993);
or UO_135 (O_135,N_2530,N_2602);
nand UO_136 (O_136,N_2955,N_2660);
nor UO_137 (O_137,N_2868,N_2537);
or UO_138 (O_138,N_2785,N_2987);
or UO_139 (O_139,N_2850,N_2697);
xor UO_140 (O_140,N_2556,N_2824);
nand UO_141 (O_141,N_2568,N_2723);
nor UO_142 (O_142,N_2920,N_2677);
nand UO_143 (O_143,N_2517,N_2595);
and UO_144 (O_144,N_2566,N_2953);
xor UO_145 (O_145,N_2683,N_2929);
xor UO_146 (O_146,N_2616,N_2699);
nor UO_147 (O_147,N_2932,N_2830);
nor UO_148 (O_148,N_2882,N_2506);
nand UO_149 (O_149,N_2972,N_2522);
nor UO_150 (O_150,N_2907,N_2751);
and UO_151 (O_151,N_2700,N_2748);
and UO_152 (O_152,N_2789,N_2890);
nor UO_153 (O_153,N_2673,N_2828);
or UO_154 (O_154,N_2992,N_2631);
nor UO_155 (O_155,N_2806,N_2995);
nand UO_156 (O_156,N_2984,N_2957);
xor UO_157 (O_157,N_2692,N_2628);
and UO_158 (O_158,N_2826,N_2676);
xor UO_159 (O_159,N_2808,N_2622);
or UO_160 (O_160,N_2611,N_2514);
nand UO_161 (O_161,N_2540,N_2994);
and UO_162 (O_162,N_2899,N_2688);
and UO_163 (O_163,N_2893,N_2504);
or UO_164 (O_164,N_2691,N_2979);
xnor UO_165 (O_165,N_2834,N_2637);
and UO_166 (O_166,N_2917,N_2767);
and UO_167 (O_167,N_2965,N_2796);
nor UO_168 (O_168,N_2551,N_2831);
nand UO_169 (O_169,N_2534,N_2741);
and UO_170 (O_170,N_2791,N_2906);
or UO_171 (O_171,N_2933,N_2529);
and UO_172 (O_172,N_2962,N_2835);
xor UO_173 (O_173,N_2612,N_2762);
or UO_174 (O_174,N_2727,N_2843);
nor UO_175 (O_175,N_2925,N_2547);
and UO_176 (O_176,N_2705,N_2597);
nor UO_177 (O_177,N_2624,N_2657);
nand UO_178 (O_178,N_2558,N_2794);
nor UO_179 (O_179,N_2960,N_2591);
nand UO_180 (O_180,N_2764,N_2732);
nor UO_181 (O_181,N_2797,N_2718);
nor UO_182 (O_182,N_2851,N_2694);
nor UO_183 (O_183,N_2703,N_2863);
or UO_184 (O_184,N_2717,N_2516);
nand UO_185 (O_185,N_2778,N_2565);
nor UO_186 (O_186,N_2930,N_2775);
and UO_187 (O_187,N_2572,N_2842);
xnor UO_188 (O_188,N_2838,N_2961);
nor UO_189 (O_189,N_2947,N_2788);
nor UO_190 (O_190,N_2892,N_2822);
nor UO_191 (O_191,N_2742,N_2704);
or UO_192 (O_192,N_2974,N_2503);
or UO_193 (O_193,N_2680,N_2564);
or UO_194 (O_194,N_2653,N_2859);
nand UO_195 (O_195,N_2776,N_2963);
xor UO_196 (O_196,N_2940,N_2571);
nand UO_197 (O_197,N_2684,N_2924);
nor UO_198 (O_198,N_2783,N_2747);
nor UO_199 (O_199,N_2702,N_2968);
nand UO_200 (O_200,N_2817,N_2598);
nand UO_201 (O_201,N_2971,N_2721);
nand UO_202 (O_202,N_2609,N_2661);
and UO_203 (O_203,N_2619,N_2869);
and UO_204 (O_204,N_2669,N_2588);
or UO_205 (O_205,N_2836,N_2784);
xor UO_206 (O_206,N_2865,N_2795);
and UO_207 (O_207,N_2966,N_2615);
or UO_208 (O_208,N_2901,N_2815);
nand UO_209 (O_209,N_2902,N_2641);
or UO_210 (O_210,N_2990,N_2675);
nor UO_211 (O_211,N_2544,N_2725);
xor UO_212 (O_212,N_2765,N_2749);
nor UO_213 (O_213,N_2590,N_2610);
nand UO_214 (O_214,N_2744,N_2709);
and UO_215 (O_215,N_2991,N_2613);
or UO_216 (O_216,N_2786,N_2538);
xor UO_217 (O_217,N_2585,N_2523);
nand UO_218 (O_218,N_2713,N_2576);
and UO_219 (O_219,N_2652,N_2663);
nor UO_220 (O_220,N_2693,N_2926);
nand UO_221 (O_221,N_2533,N_2858);
nand UO_222 (O_222,N_2543,N_2810);
xnor UO_223 (O_223,N_2668,N_2662);
and UO_224 (O_224,N_2800,N_2832);
xor UO_225 (O_225,N_2627,N_2825);
nor UO_226 (O_226,N_2510,N_2845);
and UO_227 (O_227,N_2855,N_2792);
and UO_228 (O_228,N_2670,N_2614);
nor UO_229 (O_229,N_2580,N_2603);
xnor UO_230 (O_230,N_2774,N_2592);
nor UO_231 (O_231,N_2897,N_2934);
and UO_232 (O_232,N_2643,N_2818);
nand UO_233 (O_233,N_2894,N_2532);
and UO_234 (O_234,N_2731,N_2608);
xnor UO_235 (O_235,N_2738,N_2941);
nor UO_236 (O_236,N_2664,N_2521);
or UO_237 (O_237,N_2730,N_2559);
nand UO_238 (O_238,N_2787,N_2606);
nand UO_239 (O_239,N_2650,N_2752);
xnor UO_240 (O_240,N_2682,N_2864);
or UO_241 (O_241,N_2541,N_2633);
or UO_242 (O_242,N_2582,N_2753);
xor UO_243 (O_243,N_2918,N_2763);
xor UO_244 (O_244,N_2881,N_2853);
nor UO_245 (O_245,N_2809,N_2600);
nor UO_246 (O_246,N_2781,N_2750);
and UO_247 (O_247,N_2839,N_2887);
nand UO_248 (O_248,N_2618,N_2757);
nand UO_249 (O_249,N_2577,N_2871);
nand UO_250 (O_250,N_2572,N_2696);
nor UO_251 (O_251,N_2918,N_2773);
nor UO_252 (O_252,N_2878,N_2727);
and UO_253 (O_253,N_2967,N_2528);
nand UO_254 (O_254,N_2815,N_2854);
nand UO_255 (O_255,N_2781,N_2721);
and UO_256 (O_256,N_2670,N_2574);
nor UO_257 (O_257,N_2806,N_2981);
nand UO_258 (O_258,N_2673,N_2578);
and UO_259 (O_259,N_2668,N_2998);
nor UO_260 (O_260,N_2930,N_2516);
or UO_261 (O_261,N_2785,N_2666);
xnor UO_262 (O_262,N_2580,N_2794);
nor UO_263 (O_263,N_2863,N_2659);
nor UO_264 (O_264,N_2603,N_2982);
or UO_265 (O_265,N_2614,N_2530);
and UO_266 (O_266,N_2957,N_2672);
and UO_267 (O_267,N_2824,N_2852);
nand UO_268 (O_268,N_2558,N_2772);
or UO_269 (O_269,N_2924,N_2853);
and UO_270 (O_270,N_2508,N_2768);
xnor UO_271 (O_271,N_2757,N_2797);
and UO_272 (O_272,N_2651,N_2978);
nand UO_273 (O_273,N_2546,N_2809);
or UO_274 (O_274,N_2937,N_2884);
or UO_275 (O_275,N_2741,N_2767);
nand UO_276 (O_276,N_2781,N_2903);
or UO_277 (O_277,N_2976,N_2861);
nor UO_278 (O_278,N_2559,N_2829);
or UO_279 (O_279,N_2726,N_2999);
and UO_280 (O_280,N_2670,N_2543);
nor UO_281 (O_281,N_2856,N_2841);
nor UO_282 (O_282,N_2741,N_2765);
nor UO_283 (O_283,N_2819,N_2838);
or UO_284 (O_284,N_2999,N_2758);
nand UO_285 (O_285,N_2696,N_2982);
nor UO_286 (O_286,N_2979,N_2599);
and UO_287 (O_287,N_2930,N_2679);
or UO_288 (O_288,N_2723,N_2969);
nand UO_289 (O_289,N_2923,N_2644);
nor UO_290 (O_290,N_2558,N_2586);
nand UO_291 (O_291,N_2965,N_2657);
or UO_292 (O_292,N_2564,N_2807);
nand UO_293 (O_293,N_2979,N_2727);
nand UO_294 (O_294,N_2926,N_2565);
xnor UO_295 (O_295,N_2744,N_2671);
or UO_296 (O_296,N_2936,N_2665);
xor UO_297 (O_297,N_2829,N_2791);
or UO_298 (O_298,N_2665,N_2824);
or UO_299 (O_299,N_2900,N_2650);
and UO_300 (O_300,N_2563,N_2609);
nor UO_301 (O_301,N_2594,N_2989);
or UO_302 (O_302,N_2955,N_2629);
and UO_303 (O_303,N_2748,N_2690);
and UO_304 (O_304,N_2704,N_2999);
or UO_305 (O_305,N_2926,N_2848);
xor UO_306 (O_306,N_2550,N_2733);
nor UO_307 (O_307,N_2643,N_2935);
nor UO_308 (O_308,N_2679,N_2988);
or UO_309 (O_309,N_2751,N_2755);
nand UO_310 (O_310,N_2856,N_2878);
and UO_311 (O_311,N_2843,N_2695);
or UO_312 (O_312,N_2705,N_2817);
and UO_313 (O_313,N_2714,N_2734);
nand UO_314 (O_314,N_2932,N_2659);
nand UO_315 (O_315,N_2946,N_2618);
xor UO_316 (O_316,N_2575,N_2558);
and UO_317 (O_317,N_2787,N_2978);
and UO_318 (O_318,N_2821,N_2740);
or UO_319 (O_319,N_2606,N_2741);
or UO_320 (O_320,N_2817,N_2656);
and UO_321 (O_321,N_2736,N_2791);
nand UO_322 (O_322,N_2796,N_2926);
and UO_323 (O_323,N_2647,N_2857);
nor UO_324 (O_324,N_2779,N_2898);
nand UO_325 (O_325,N_2977,N_2687);
nand UO_326 (O_326,N_2805,N_2938);
or UO_327 (O_327,N_2804,N_2988);
nor UO_328 (O_328,N_2719,N_2821);
nand UO_329 (O_329,N_2916,N_2583);
or UO_330 (O_330,N_2707,N_2886);
and UO_331 (O_331,N_2670,N_2905);
nand UO_332 (O_332,N_2690,N_2563);
or UO_333 (O_333,N_2865,N_2773);
nor UO_334 (O_334,N_2537,N_2999);
nand UO_335 (O_335,N_2804,N_2773);
nand UO_336 (O_336,N_2502,N_2874);
nand UO_337 (O_337,N_2691,N_2606);
or UO_338 (O_338,N_2791,N_2986);
and UO_339 (O_339,N_2873,N_2831);
xnor UO_340 (O_340,N_2726,N_2740);
or UO_341 (O_341,N_2522,N_2623);
or UO_342 (O_342,N_2685,N_2824);
and UO_343 (O_343,N_2819,N_2897);
or UO_344 (O_344,N_2978,N_2549);
nand UO_345 (O_345,N_2986,N_2605);
nand UO_346 (O_346,N_2765,N_2692);
xor UO_347 (O_347,N_2573,N_2769);
nand UO_348 (O_348,N_2546,N_2860);
nand UO_349 (O_349,N_2944,N_2608);
nand UO_350 (O_350,N_2813,N_2913);
and UO_351 (O_351,N_2549,N_2617);
or UO_352 (O_352,N_2539,N_2884);
nand UO_353 (O_353,N_2792,N_2537);
nand UO_354 (O_354,N_2602,N_2639);
or UO_355 (O_355,N_2776,N_2968);
or UO_356 (O_356,N_2715,N_2908);
nor UO_357 (O_357,N_2502,N_2682);
or UO_358 (O_358,N_2639,N_2900);
or UO_359 (O_359,N_2781,N_2562);
nand UO_360 (O_360,N_2644,N_2882);
xor UO_361 (O_361,N_2806,N_2512);
xnor UO_362 (O_362,N_2632,N_2707);
xnor UO_363 (O_363,N_2708,N_2685);
or UO_364 (O_364,N_2962,N_2848);
and UO_365 (O_365,N_2791,N_2618);
or UO_366 (O_366,N_2726,N_2596);
xor UO_367 (O_367,N_2650,N_2515);
xnor UO_368 (O_368,N_2809,N_2898);
and UO_369 (O_369,N_2601,N_2899);
nor UO_370 (O_370,N_2518,N_2933);
or UO_371 (O_371,N_2543,N_2786);
xor UO_372 (O_372,N_2522,N_2585);
nor UO_373 (O_373,N_2848,N_2684);
nor UO_374 (O_374,N_2628,N_2560);
and UO_375 (O_375,N_2669,N_2696);
and UO_376 (O_376,N_2997,N_2934);
and UO_377 (O_377,N_2991,N_2587);
nand UO_378 (O_378,N_2518,N_2706);
or UO_379 (O_379,N_2612,N_2936);
nand UO_380 (O_380,N_2810,N_2502);
or UO_381 (O_381,N_2719,N_2500);
nand UO_382 (O_382,N_2696,N_2658);
and UO_383 (O_383,N_2945,N_2874);
nor UO_384 (O_384,N_2786,N_2711);
and UO_385 (O_385,N_2774,N_2743);
and UO_386 (O_386,N_2840,N_2912);
nor UO_387 (O_387,N_2539,N_2752);
nor UO_388 (O_388,N_2854,N_2539);
nor UO_389 (O_389,N_2947,N_2887);
nand UO_390 (O_390,N_2810,N_2586);
and UO_391 (O_391,N_2523,N_2868);
nand UO_392 (O_392,N_2654,N_2692);
nor UO_393 (O_393,N_2556,N_2575);
nand UO_394 (O_394,N_2697,N_2615);
or UO_395 (O_395,N_2830,N_2666);
and UO_396 (O_396,N_2667,N_2771);
or UO_397 (O_397,N_2597,N_2975);
nand UO_398 (O_398,N_2925,N_2565);
nor UO_399 (O_399,N_2888,N_2922);
and UO_400 (O_400,N_2595,N_2695);
or UO_401 (O_401,N_2883,N_2959);
or UO_402 (O_402,N_2633,N_2625);
or UO_403 (O_403,N_2826,N_2627);
nor UO_404 (O_404,N_2814,N_2989);
and UO_405 (O_405,N_2748,N_2660);
nor UO_406 (O_406,N_2736,N_2720);
nand UO_407 (O_407,N_2893,N_2630);
or UO_408 (O_408,N_2631,N_2556);
or UO_409 (O_409,N_2553,N_2648);
nand UO_410 (O_410,N_2704,N_2956);
or UO_411 (O_411,N_2825,N_2719);
and UO_412 (O_412,N_2520,N_2978);
nand UO_413 (O_413,N_2702,N_2590);
or UO_414 (O_414,N_2600,N_2531);
nand UO_415 (O_415,N_2577,N_2575);
nor UO_416 (O_416,N_2791,N_2916);
nand UO_417 (O_417,N_2675,N_2836);
and UO_418 (O_418,N_2857,N_2990);
or UO_419 (O_419,N_2790,N_2676);
and UO_420 (O_420,N_2575,N_2798);
or UO_421 (O_421,N_2520,N_2934);
nor UO_422 (O_422,N_2715,N_2690);
nand UO_423 (O_423,N_2556,N_2517);
nand UO_424 (O_424,N_2961,N_2618);
or UO_425 (O_425,N_2642,N_2503);
nand UO_426 (O_426,N_2978,N_2760);
xnor UO_427 (O_427,N_2726,N_2709);
or UO_428 (O_428,N_2507,N_2759);
or UO_429 (O_429,N_2776,N_2680);
and UO_430 (O_430,N_2894,N_2957);
or UO_431 (O_431,N_2666,N_2585);
or UO_432 (O_432,N_2651,N_2997);
and UO_433 (O_433,N_2591,N_2909);
or UO_434 (O_434,N_2716,N_2542);
nor UO_435 (O_435,N_2710,N_2848);
nor UO_436 (O_436,N_2787,N_2835);
nor UO_437 (O_437,N_2764,N_2748);
nand UO_438 (O_438,N_2877,N_2641);
nor UO_439 (O_439,N_2781,N_2532);
nor UO_440 (O_440,N_2927,N_2630);
or UO_441 (O_441,N_2738,N_2887);
nand UO_442 (O_442,N_2903,N_2732);
nor UO_443 (O_443,N_2764,N_2876);
and UO_444 (O_444,N_2808,N_2783);
nor UO_445 (O_445,N_2722,N_2729);
xnor UO_446 (O_446,N_2954,N_2501);
nor UO_447 (O_447,N_2810,N_2518);
nand UO_448 (O_448,N_2931,N_2559);
nor UO_449 (O_449,N_2538,N_2940);
xnor UO_450 (O_450,N_2703,N_2837);
or UO_451 (O_451,N_2723,N_2569);
xnor UO_452 (O_452,N_2852,N_2768);
or UO_453 (O_453,N_2670,N_2591);
xnor UO_454 (O_454,N_2744,N_2994);
nand UO_455 (O_455,N_2696,N_2500);
xnor UO_456 (O_456,N_2993,N_2661);
nand UO_457 (O_457,N_2626,N_2760);
xnor UO_458 (O_458,N_2922,N_2925);
nor UO_459 (O_459,N_2811,N_2530);
nand UO_460 (O_460,N_2925,N_2966);
nand UO_461 (O_461,N_2643,N_2707);
and UO_462 (O_462,N_2890,N_2808);
xnor UO_463 (O_463,N_2744,N_2714);
nand UO_464 (O_464,N_2833,N_2937);
and UO_465 (O_465,N_2634,N_2730);
and UO_466 (O_466,N_2508,N_2561);
or UO_467 (O_467,N_2567,N_2662);
or UO_468 (O_468,N_2926,N_2853);
or UO_469 (O_469,N_2633,N_2568);
nand UO_470 (O_470,N_2607,N_2653);
or UO_471 (O_471,N_2501,N_2808);
or UO_472 (O_472,N_2738,N_2728);
nor UO_473 (O_473,N_2755,N_2639);
or UO_474 (O_474,N_2671,N_2777);
nand UO_475 (O_475,N_2680,N_2992);
nand UO_476 (O_476,N_2543,N_2947);
nor UO_477 (O_477,N_2931,N_2515);
nand UO_478 (O_478,N_2611,N_2600);
nand UO_479 (O_479,N_2555,N_2898);
or UO_480 (O_480,N_2820,N_2597);
nand UO_481 (O_481,N_2855,N_2563);
xnor UO_482 (O_482,N_2575,N_2672);
nor UO_483 (O_483,N_2635,N_2755);
nor UO_484 (O_484,N_2906,N_2526);
and UO_485 (O_485,N_2850,N_2535);
or UO_486 (O_486,N_2691,N_2811);
or UO_487 (O_487,N_2835,N_2502);
nor UO_488 (O_488,N_2526,N_2633);
nand UO_489 (O_489,N_2791,N_2548);
or UO_490 (O_490,N_2814,N_2996);
nor UO_491 (O_491,N_2941,N_2807);
nor UO_492 (O_492,N_2922,N_2524);
and UO_493 (O_493,N_2986,N_2792);
nor UO_494 (O_494,N_2558,N_2731);
nand UO_495 (O_495,N_2508,N_2872);
nand UO_496 (O_496,N_2932,N_2539);
nor UO_497 (O_497,N_2929,N_2713);
and UO_498 (O_498,N_2837,N_2678);
or UO_499 (O_499,N_2623,N_2529);
endmodule