module basic_500_3000_500_40_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_167,In_322);
nand U1 (N_1,In_395,In_188);
or U2 (N_2,In_238,In_106);
nor U3 (N_3,In_251,In_38);
nor U4 (N_4,In_494,In_276);
or U5 (N_5,In_182,In_163);
and U6 (N_6,In_399,In_194);
xor U7 (N_7,In_176,In_434);
or U8 (N_8,In_409,In_398);
or U9 (N_9,In_135,In_459);
nand U10 (N_10,In_295,In_408);
nor U11 (N_11,In_103,In_485);
and U12 (N_12,In_283,In_444);
or U13 (N_13,In_420,In_7);
and U14 (N_14,In_56,In_456);
and U15 (N_15,In_370,In_275);
and U16 (N_16,In_385,In_457);
or U17 (N_17,In_102,In_467);
and U18 (N_18,In_120,In_104);
or U19 (N_19,In_392,In_29);
and U20 (N_20,In_393,In_209);
and U21 (N_21,In_156,In_458);
or U22 (N_22,In_235,In_247);
or U23 (N_23,In_481,In_292);
nor U24 (N_24,In_415,In_166);
nand U25 (N_25,In_119,In_112);
and U26 (N_26,In_476,In_412);
or U27 (N_27,In_67,In_495);
nor U28 (N_28,In_35,In_315);
nor U29 (N_29,In_333,In_452);
nor U30 (N_30,In_498,In_88);
and U31 (N_31,In_34,In_468);
and U32 (N_32,In_100,In_221);
and U33 (N_33,In_255,In_319);
or U34 (N_34,In_219,In_285);
nor U35 (N_35,In_271,In_410);
or U36 (N_36,In_310,In_232);
or U37 (N_37,In_157,In_348);
nor U38 (N_38,In_63,In_391);
nand U39 (N_39,In_294,In_215);
nor U40 (N_40,In_321,In_225);
or U41 (N_41,In_186,In_107);
nor U42 (N_42,In_33,In_201);
or U43 (N_43,In_281,In_93);
nor U44 (N_44,In_496,In_358);
nor U45 (N_45,In_82,In_473);
nand U46 (N_46,In_447,In_413);
or U47 (N_47,In_65,In_31);
nor U48 (N_48,In_70,In_486);
nor U49 (N_49,In_224,In_222);
or U50 (N_50,In_170,In_461);
nand U51 (N_51,In_228,In_161);
and U52 (N_52,In_90,In_363);
nor U53 (N_53,In_328,In_58);
and U54 (N_54,In_8,In_20);
or U55 (N_55,In_84,In_68);
nor U56 (N_56,In_350,In_14);
and U57 (N_57,In_424,In_37);
nor U58 (N_58,In_440,In_105);
nand U59 (N_59,In_454,In_180);
nor U60 (N_60,In_139,In_52);
nor U61 (N_61,In_24,In_10);
nand U62 (N_62,In_162,In_448);
nand U63 (N_63,In_158,In_325);
nand U64 (N_64,In_89,In_150);
nand U65 (N_65,In_282,In_378);
nand U66 (N_66,In_323,In_324);
or U67 (N_67,In_168,In_347);
nor U68 (N_68,In_472,In_195);
nand U69 (N_69,In_76,In_335);
nor U70 (N_70,In_55,In_446);
nor U71 (N_71,In_435,In_354);
nand U72 (N_72,In_18,In_305);
and U73 (N_73,In_451,In_164);
or U74 (N_74,In_236,In_192);
nor U75 (N_75,In_425,In_353);
or U76 (N_76,In_183,In_470);
nand U77 (N_77,In_369,In_288);
or U78 (N_78,In_109,In_124);
and U79 (N_79,N_2,N_43);
nand U80 (N_80,In_75,In_404);
and U81 (N_81,In_60,In_240);
or U82 (N_82,In_421,In_289);
nor U83 (N_83,In_118,In_433);
and U84 (N_84,N_8,In_401);
and U85 (N_85,In_359,N_3);
xor U86 (N_86,In_250,In_185);
nor U87 (N_87,In_334,In_389);
or U88 (N_88,In_122,In_26);
nand U89 (N_89,In_491,In_422);
nor U90 (N_90,In_368,In_50);
and U91 (N_91,In_87,In_173);
or U92 (N_92,In_307,In_216);
or U93 (N_93,In_145,In_212);
nand U94 (N_94,In_474,In_407);
and U95 (N_95,In_441,In_9);
nor U96 (N_96,N_35,N_32);
and U97 (N_97,In_121,In_267);
nand U98 (N_98,In_460,In_92);
or U99 (N_99,In_297,In_95);
or U100 (N_100,In_260,In_390);
and U101 (N_101,N_67,In_367);
and U102 (N_102,In_462,In_202);
and U103 (N_103,In_246,In_445);
nor U104 (N_104,In_141,In_364);
nor U105 (N_105,In_40,In_428);
nand U106 (N_106,In_177,In_419);
nand U107 (N_107,In_205,In_365);
and U108 (N_108,In_306,N_31);
nor U109 (N_109,In_361,In_355);
and U110 (N_110,In_326,N_23);
or U111 (N_111,N_28,In_455);
and U112 (N_112,In_349,In_85);
nor U113 (N_113,In_77,In_142);
and U114 (N_114,N_4,N_70);
nand U115 (N_115,N_49,In_4);
or U116 (N_116,In_264,In_175);
nor U117 (N_117,In_160,In_430);
nand U118 (N_118,In_406,N_33);
or U119 (N_119,N_19,N_24);
nand U120 (N_120,In_108,In_482);
nor U121 (N_121,In_366,In_165);
or U122 (N_122,In_133,In_19);
or U123 (N_123,In_449,In_475);
and U124 (N_124,In_479,In_181);
or U125 (N_125,In_6,In_290);
nor U126 (N_126,N_15,In_371);
nor U127 (N_127,In_218,In_72);
and U128 (N_128,In_465,In_230);
and U129 (N_129,In_45,N_27);
nor U130 (N_130,In_394,In_111);
and U131 (N_131,In_253,In_477);
nand U132 (N_132,In_471,In_488);
nor U133 (N_133,In_98,N_39);
and U134 (N_134,In_15,In_2);
and U135 (N_135,N_69,In_234);
and U136 (N_136,In_416,In_48);
nand U137 (N_137,N_63,In_134);
nand U138 (N_138,In_155,N_16);
or U139 (N_139,N_20,N_44);
nor U140 (N_140,In_317,In_376);
or U141 (N_141,In_483,N_64);
nand U142 (N_142,N_1,N_37);
or U143 (N_143,In_61,In_5);
nand U144 (N_144,In_339,In_402);
and U145 (N_145,In_388,In_360);
and U146 (N_146,In_336,In_492);
nand U147 (N_147,N_11,In_439);
and U148 (N_148,In_136,N_66);
and U149 (N_149,In_280,N_52);
nor U150 (N_150,N_13,N_55);
and U151 (N_151,In_258,In_387);
nor U152 (N_152,In_153,N_149);
or U153 (N_153,In_229,N_6);
and U154 (N_154,In_32,N_90);
nor U155 (N_155,In_41,In_73);
nor U156 (N_156,In_78,N_61);
nand U157 (N_157,N_78,In_97);
nor U158 (N_158,N_41,In_128);
or U159 (N_159,In_331,In_478);
nand U160 (N_160,N_46,N_100);
and U161 (N_161,N_112,In_96);
nand U162 (N_162,In_261,In_127);
and U163 (N_163,In_223,N_18);
or U164 (N_164,In_397,N_29);
or U165 (N_165,In_342,In_79);
or U166 (N_166,N_57,In_208);
and U167 (N_167,In_263,In_42);
nand U168 (N_168,In_21,N_54);
and U169 (N_169,N_118,In_129);
nor U170 (N_170,In_345,N_105);
nor U171 (N_171,In_43,In_47);
xnor U172 (N_172,In_278,In_254);
nand U173 (N_173,In_28,In_356);
nand U174 (N_174,N_113,In_381);
and U175 (N_175,N_101,N_141);
nor U176 (N_176,N_30,N_21);
nor U177 (N_177,In_154,N_98);
nor U178 (N_178,In_302,In_436);
nand U179 (N_179,In_231,In_343);
nor U180 (N_180,N_53,In_206);
nand U181 (N_181,In_341,N_131);
and U182 (N_182,N_50,In_309);
and U183 (N_183,In_137,N_82);
or U184 (N_184,In_316,N_74);
nor U185 (N_185,In_0,In_346);
and U186 (N_186,N_106,N_95);
and U187 (N_187,In_184,N_120);
nand U188 (N_188,In_116,In_62);
nor U189 (N_189,In_405,N_26);
or U190 (N_190,N_79,In_362);
nand U191 (N_191,N_68,N_126);
nor U192 (N_192,In_17,In_36);
nor U193 (N_193,In_99,In_12);
or U194 (N_194,In_450,In_132);
nor U195 (N_195,In_148,In_330);
and U196 (N_196,In_373,In_466);
and U197 (N_197,N_134,In_344);
and U198 (N_198,In_384,In_418);
or U199 (N_199,In_114,In_16);
or U200 (N_200,N_147,In_277);
or U201 (N_201,N_92,N_97);
nand U202 (N_202,In_338,In_71);
or U203 (N_203,N_60,N_115);
or U204 (N_204,N_122,In_140);
nand U205 (N_205,In_248,In_25);
and U206 (N_206,In_259,In_241);
and U207 (N_207,N_148,N_22);
and U208 (N_208,In_199,N_132);
nor U209 (N_209,N_38,In_337);
nor U210 (N_210,N_47,In_423);
nor U211 (N_211,N_107,In_357);
and U212 (N_212,In_81,In_211);
and U213 (N_213,N_81,In_442);
and U214 (N_214,In_300,N_83);
or U215 (N_215,In_200,N_34);
or U216 (N_216,N_77,In_286);
or U217 (N_217,N_121,In_101);
nor U218 (N_218,In_327,In_308);
nand U219 (N_219,In_203,In_414);
nor U220 (N_220,In_190,N_143);
nor U221 (N_221,In_427,In_91);
nor U222 (N_222,In_113,N_62);
and U223 (N_223,In_379,In_411);
and U224 (N_224,In_198,In_123);
nor U225 (N_225,N_5,In_332);
and U226 (N_226,N_179,In_152);
xnor U227 (N_227,N_36,N_117);
nor U228 (N_228,In_493,N_59);
or U229 (N_229,N_166,N_174);
nand U230 (N_230,N_172,N_116);
and U231 (N_231,N_99,N_9);
nand U232 (N_232,In_54,In_386);
and U233 (N_233,In_227,N_216);
nor U234 (N_234,N_133,N_175);
nand U235 (N_235,N_164,N_127);
nor U236 (N_236,In_179,In_64);
nor U237 (N_237,In_274,In_53);
and U238 (N_238,N_176,In_239);
and U239 (N_239,In_245,In_320);
nor U240 (N_240,N_14,In_147);
nand U241 (N_241,N_86,In_453);
and U242 (N_242,N_209,In_318);
and U243 (N_243,In_27,N_185);
nand U244 (N_244,N_171,In_11);
nand U245 (N_245,In_464,N_48);
nor U246 (N_246,In_143,N_220);
or U247 (N_247,In_144,In_30);
or U248 (N_248,N_222,N_168);
and U249 (N_249,In_375,In_189);
or U250 (N_250,In_438,N_205);
and U251 (N_251,N_42,In_57);
nand U252 (N_252,N_110,In_220);
nand U253 (N_253,N_200,In_149);
nand U254 (N_254,N_125,In_51);
nor U255 (N_255,In_44,N_84);
nand U256 (N_256,In_396,In_39);
nand U257 (N_257,In_86,In_174);
nor U258 (N_258,N_192,N_96);
nor U259 (N_259,N_211,In_311);
or U260 (N_260,N_218,N_189);
nor U261 (N_261,N_158,In_299);
nand U262 (N_262,N_102,N_130);
and U263 (N_263,In_279,In_298);
or U264 (N_264,N_123,N_163);
or U265 (N_265,N_224,N_207);
or U266 (N_266,N_201,In_138);
nor U267 (N_267,N_199,In_80);
or U268 (N_268,N_187,In_146);
and U269 (N_269,N_111,In_329);
nor U270 (N_270,In_207,In_352);
nand U271 (N_271,In_266,N_88);
nand U272 (N_272,N_144,In_287);
nor U273 (N_273,In_351,N_193);
or U274 (N_274,N_161,N_157);
and U275 (N_275,In_380,N_214);
nand U276 (N_276,N_169,In_273);
or U277 (N_277,N_197,N_124);
xnor U278 (N_278,In_265,In_463);
or U279 (N_279,In_270,N_146);
xnor U280 (N_280,In_469,N_93);
and U281 (N_281,N_103,N_195);
or U282 (N_282,In_1,N_137);
and U283 (N_283,In_169,N_180);
and U284 (N_284,N_51,N_188);
nor U285 (N_285,N_203,In_193);
nand U286 (N_286,N_76,In_303);
and U287 (N_287,In_242,N_71);
and U288 (N_288,In_497,N_72);
or U289 (N_289,N_85,In_499);
nand U290 (N_290,In_210,In_151);
and U291 (N_291,In_204,In_237);
or U292 (N_292,In_426,N_212);
nand U293 (N_293,N_223,In_196);
nor U294 (N_294,N_75,N_136);
nor U295 (N_295,N_150,In_59);
nand U296 (N_296,In_304,In_244);
or U297 (N_297,N_160,N_56);
nor U298 (N_298,In_197,In_443);
or U299 (N_299,N_215,In_214);
nand U300 (N_300,In_432,N_273);
and U301 (N_301,N_270,N_231);
nor U302 (N_302,In_178,N_65);
nand U303 (N_303,In_284,In_49);
nor U304 (N_304,N_248,In_226);
and U305 (N_305,N_221,N_204);
or U306 (N_306,N_249,In_130);
and U307 (N_307,N_153,N_217);
nand U308 (N_308,N_232,N_236);
or U309 (N_309,N_155,N_94);
and U310 (N_310,In_66,N_229);
and U311 (N_311,N_138,In_13);
and U312 (N_312,N_292,N_73);
nand U313 (N_313,N_165,N_173);
or U314 (N_314,N_279,N_109);
nand U315 (N_315,In_256,N_288);
nand U316 (N_316,In_489,N_282);
nand U317 (N_317,N_80,N_264);
or U318 (N_318,In_400,In_23);
nand U319 (N_319,N_259,N_108);
and U320 (N_320,N_267,N_276);
nand U321 (N_321,In_125,N_234);
nand U322 (N_322,In_252,In_74);
nand U323 (N_323,In_484,In_480);
and U324 (N_324,N_119,N_285);
nand U325 (N_325,N_265,N_152);
nand U326 (N_326,In_171,N_89);
or U327 (N_327,N_281,N_17);
nand U328 (N_328,N_258,In_213);
nor U329 (N_329,In_372,In_403);
nand U330 (N_330,In_115,In_3);
nor U331 (N_331,N_206,N_295);
nand U332 (N_332,N_114,N_289);
nor U333 (N_333,N_280,N_241);
or U334 (N_334,N_278,N_40);
nor U335 (N_335,N_170,N_210);
and U336 (N_336,In_340,In_131);
nor U337 (N_337,N_182,N_291);
or U338 (N_338,N_202,In_126);
and U339 (N_339,In_262,N_151);
or U340 (N_340,N_247,In_110);
nand U341 (N_341,In_383,N_253);
and U342 (N_342,N_191,N_178);
and U343 (N_343,N_240,N_0);
or U344 (N_344,N_244,N_45);
nand U345 (N_345,In_377,N_239);
and U346 (N_346,N_58,N_237);
and U347 (N_347,N_266,N_286);
and U348 (N_348,N_225,N_140);
and U349 (N_349,N_228,In_382);
or U350 (N_350,N_233,N_261);
and U351 (N_351,N_219,N_159);
nand U352 (N_352,N_260,N_181);
and U353 (N_353,In_296,In_22);
and U354 (N_354,In_293,N_298);
and U355 (N_355,N_167,In_159);
or U356 (N_356,N_277,N_245);
and U357 (N_357,N_91,In_272);
nand U358 (N_358,In_429,N_274);
and U359 (N_359,N_284,N_196);
nor U360 (N_360,N_128,N_104);
or U361 (N_361,N_296,In_46);
nor U362 (N_362,In_291,N_263);
and U363 (N_363,N_251,N_272);
nor U364 (N_364,N_87,N_268);
and U365 (N_365,In_217,In_490);
nand U366 (N_366,In_94,N_275);
and U367 (N_367,In_257,N_213);
nor U368 (N_368,N_145,N_271);
or U369 (N_369,N_162,N_194);
nor U370 (N_370,In_374,In_301);
or U371 (N_371,N_156,N_262);
and U372 (N_372,N_294,N_226);
nor U373 (N_373,N_252,N_12);
nor U374 (N_374,N_154,In_417);
xor U375 (N_375,N_316,In_243);
or U376 (N_376,N_356,N_307);
xor U377 (N_377,In_187,N_366);
nor U378 (N_378,N_255,N_319);
or U379 (N_379,N_311,N_332);
and U380 (N_380,N_326,N_177);
nand U381 (N_381,N_365,N_334);
or U382 (N_382,N_313,N_341);
nor U383 (N_383,N_359,N_355);
nand U384 (N_384,N_230,N_374);
nor U385 (N_385,N_246,N_338);
or U386 (N_386,N_329,N_333);
or U387 (N_387,N_10,N_310);
or U388 (N_388,N_320,N_142);
or U389 (N_389,N_372,N_331);
xor U390 (N_390,N_293,In_313);
nand U391 (N_391,N_243,In_83);
xnor U392 (N_392,N_340,In_312);
or U393 (N_393,N_328,N_301);
nand U394 (N_394,N_350,N_290);
nand U395 (N_395,N_327,N_312);
nor U396 (N_396,In_117,N_25);
and U397 (N_397,N_371,N_325);
nor U398 (N_398,N_324,N_357);
or U399 (N_399,N_297,N_306);
nor U400 (N_400,N_322,N_238);
nand U401 (N_401,N_323,N_364);
and U402 (N_402,N_309,N_250);
and U403 (N_403,N_361,N_363);
xor U404 (N_404,N_369,N_342);
nor U405 (N_405,N_308,N_184);
or U406 (N_406,In_191,N_337);
and U407 (N_407,In_69,In_249);
nor U408 (N_408,N_336,N_139);
nor U409 (N_409,N_190,N_254);
or U410 (N_410,N_135,N_367);
or U411 (N_411,N_287,In_431);
and U412 (N_412,N_299,N_362);
and U413 (N_413,N_339,N_283);
nor U414 (N_414,N_227,N_208);
nor U415 (N_415,N_235,N_370);
nor U416 (N_416,N_198,In_487);
nor U417 (N_417,In_268,N_256);
nand U418 (N_418,N_315,In_269);
or U419 (N_419,N_353,N_343);
or U420 (N_420,N_129,In_233);
nand U421 (N_421,N_346,N_300);
nor U422 (N_422,N_257,N_348);
and U423 (N_423,N_304,N_358);
and U424 (N_424,N_303,N_360);
or U425 (N_425,N_368,N_335);
and U426 (N_426,N_345,N_373);
nand U427 (N_427,In_314,N_330);
nor U428 (N_428,N_347,N_305);
or U429 (N_429,N_269,In_172);
nor U430 (N_430,N_318,In_437);
nor U431 (N_431,N_183,N_344);
nand U432 (N_432,N_321,N_242);
or U433 (N_433,N_352,N_354);
nand U434 (N_434,N_186,N_317);
or U435 (N_435,N_7,N_302);
or U436 (N_436,N_314,N_351);
nor U437 (N_437,N_349,N_364);
or U438 (N_438,N_250,N_340);
nor U439 (N_439,N_337,In_437);
and U440 (N_440,N_374,N_357);
nor U441 (N_441,N_330,N_302);
nand U442 (N_442,N_313,N_364);
nand U443 (N_443,N_227,N_360);
and U444 (N_444,In_313,N_341);
nand U445 (N_445,N_354,N_363);
or U446 (N_446,N_301,N_329);
nand U447 (N_447,N_368,N_309);
or U448 (N_448,N_186,N_363);
nor U449 (N_449,N_350,In_117);
nand U450 (N_450,N_448,N_424);
and U451 (N_451,N_431,N_392);
nor U452 (N_452,N_449,N_417);
or U453 (N_453,N_444,N_399);
nand U454 (N_454,N_402,N_391);
and U455 (N_455,N_405,N_435);
or U456 (N_456,N_383,N_390);
nor U457 (N_457,N_422,N_419);
and U458 (N_458,N_426,N_420);
nand U459 (N_459,N_400,N_427);
or U460 (N_460,N_428,N_441);
nor U461 (N_461,N_416,N_437);
or U462 (N_462,N_388,N_410);
or U463 (N_463,N_376,N_386);
and U464 (N_464,N_415,N_398);
or U465 (N_465,N_443,N_396);
nand U466 (N_466,N_377,N_442);
or U467 (N_467,N_379,N_434);
nand U468 (N_468,N_447,N_446);
nor U469 (N_469,N_412,N_421);
nand U470 (N_470,N_433,N_432);
or U471 (N_471,N_384,N_378);
nand U472 (N_472,N_394,N_401);
and U473 (N_473,N_381,N_380);
or U474 (N_474,N_429,N_404);
and U475 (N_475,N_406,N_413);
and U476 (N_476,N_418,N_414);
nand U477 (N_477,N_385,N_389);
or U478 (N_478,N_440,N_439);
nand U479 (N_479,N_425,N_375);
or U480 (N_480,N_430,N_438);
or U481 (N_481,N_411,N_397);
and U482 (N_482,N_393,N_387);
or U483 (N_483,N_436,N_409);
nand U484 (N_484,N_382,N_403);
nand U485 (N_485,N_423,N_408);
nor U486 (N_486,N_445,N_407);
or U487 (N_487,N_395,N_415);
nand U488 (N_488,N_433,N_408);
nor U489 (N_489,N_416,N_447);
or U490 (N_490,N_389,N_424);
nand U491 (N_491,N_387,N_406);
or U492 (N_492,N_422,N_406);
or U493 (N_493,N_413,N_388);
or U494 (N_494,N_447,N_439);
and U495 (N_495,N_382,N_407);
or U496 (N_496,N_404,N_423);
and U497 (N_497,N_375,N_410);
and U498 (N_498,N_439,N_376);
and U499 (N_499,N_414,N_429);
or U500 (N_500,N_430,N_402);
nor U501 (N_501,N_430,N_446);
and U502 (N_502,N_440,N_393);
and U503 (N_503,N_400,N_387);
nand U504 (N_504,N_394,N_441);
nor U505 (N_505,N_381,N_377);
and U506 (N_506,N_417,N_391);
and U507 (N_507,N_404,N_398);
or U508 (N_508,N_433,N_401);
nor U509 (N_509,N_418,N_407);
or U510 (N_510,N_391,N_432);
nor U511 (N_511,N_448,N_386);
or U512 (N_512,N_395,N_428);
nand U513 (N_513,N_436,N_379);
and U514 (N_514,N_422,N_441);
and U515 (N_515,N_405,N_411);
nor U516 (N_516,N_427,N_388);
nand U517 (N_517,N_446,N_395);
and U518 (N_518,N_399,N_376);
or U519 (N_519,N_415,N_424);
nand U520 (N_520,N_420,N_412);
and U521 (N_521,N_398,N_387);
nand U522 (N_522,N_425,N_376);
nand U523 (N_523,N_390,N_399);
nand U524 (N_524,N_419,N_391);
nor U525 (N_525,N_518,N_502);
nor U526 (N_526,N_463,N_513);
or U527 (N_527,N_454,N_494);
and U528 (N_528,N_508,N_484);
or U529 (N_529,N_524,N_512);
nand U530 (N_530,N_523,N_517);
and U531 (N_531,N_453,N_455);
nor U532 (N_532,N_481,N_495);
nor U533 (N_533,N_476,N_488);
nor U534 (N_534,N_489,N_470);
or U535 (N_535,N_464,N_472);
nand U536 (N_536,N_451,N_515);
nand U537 (N_537,N_521,N_474);
and U538 (N_538,N_466,N_467);
and U539 (N_539,N_485,N_458);
and U540 (N_540,N_461,N_496);
or U541 (N_541,N_511,N_473);
nand U542 (N_542,N_469,N_457);
and U543 (N_543,N_465,N_482);
nor U544 (N_544,N_462,N_509);
or U545 (N_545,N_487,N_516);
or U546 (N_546,N_493,N_504);
and U547 (N_547,N_483,N_506);
nand U548 (N_548,N_490,N_503);
or U549 (N_549,N_491,N_450);
and U550 (N_550,N_486,N_507);
nor U551 (N_551,N_468,N_460);
nor U552 (N_552,N_501,N_522);
xnor U553 (N_553,N_497,N_519);
and U554 (N_554,N_456,N_471);
nand U555 (N_555,N_514,N_520);
nand U556 (N_556,N_499,N_498);
nor U557 (N_557,N_492,N_510);
and U558 (N_558,N_500,N_479);
and U559 (N_559,N_475,N_477);
nand U560 (N_560,N_505,N_452);
nor U561 (N_561,N_478,N_480);
nor U562 (N_562,N_459,N_461);
and U563 (N_563,N_500,N_456);
nand U564 (N_564,N_502,N_457);
or U565 (N_565,N_500,N_482);
or U566 (N_566,N_489,N_493);
and U567 (N_567,N_464,N_475);
nand U568 (N_568,N_460,N_472);
or U569 (N_569,N_483,N_488);
nor U570 (N_570,N_518,N_461);
or U571 (N_571,N_512,N_522);
or U572 (N_572,N_477,N_458);
and U573 (N_573,N_450,N_497);
or U574 (N_574,N_523,N_511);
or U575 (N_575,N_523,N_483);
or U576 (N_576,N_474,N_454);
or U577 (N_577,N_462,N_471);
nand U578 (N_578,N_467,N_512);
or U579 (N_579,N_511,N_477);
and U580 (N_580,N_524,N_513);
or U581 (N_581,N_508,N_461);
nor U582 (N_582,N_476,N_486);
and U583 (N_583,N_494,N_517);
nor U584 (N_584,N_488,N_458);
nor U585 (N_585,N_458,N_516);
nand U586 (N_586,N_490,N_488);
or U587 (N_587,N_492,N_465);
or U588 (N_588,N_466,N_490);
nor U589 (N_589,N_501,N_453);
xnor U590 (N_590,N_461,N_488);
and U591 (N_591,N_474,N_450);
and U592 (N_592,N_515,N_480);
and U593 (N_593,N_513,N_523);
and U594 (N_594,N_487,N_455);
or U595 (N_595,N_456,N_460);
nor U596 (N_596,N_451,N_480);
nor U597 (N_597,N_451,N_460);
nor U598 (N_598,N_505,N_461);
nor U599 (N_599,N_452,N_493);
and U600 (N_600,N_575,N_574);
or U601 (N_601,N_536,N_532);
nor U602 (N_602,N_525,N_587);
nand U603 (N_603,N_565,N_544);
nand U604 (N_604,N_555,N_535);
or U605 (N_605,N_589,N_583);
and U606 (N_606,N_599,N_567);
and U607 (N_607,N_527,N_569);
and U608 (N_608,N_551,N_579);
nand U609 (N_609,N_597,N_542);
nor U610 (N_610,N_592,N_546);
and U611 (N_611,N_553,N_563);
nand U612 (N_612,N_571,N_550);
or U613 (N_613,N_529,N_533);
and U614 (N_614,N_576,N_573);
and U615 (N_615,N_584,N_552);
or U616 (N_616,N_526,N_598);
nor U617 (N_617,N_547,N_570);
nand U618 (N_618,N_568,N_591);
nand U619 (N_619,N_578,N_585);
nor U620 (N_620,N_566,N_586);
nand U621 (N_621,N_590,N_572);
and U622 (N_622,N_549,N_561);
and U623 (N_623,N_548,N_593);
nor U624 (N_624,N_540,N_538);
or U625 (N_625,N_595,N_558);
or U626 (N_626,N_556,N_562);
nand U627 (N_627,N_581,N_588);
nor U628 (N_628,N_531,N_564);
and U629 (N_629,N_537,N_557);
or U630 (N_630,N_594,N_530);
or U631 (N_631,N_541,N_560);
nand U632 (N_632,N_539,N_577);
and U633 (N_633,N_596,N_543);
or U634 (N_634,N_528,N_545);
nor U635 (N_635,N_534,N_582);
and U636 (N_636,N_580,N_554);
or U637 (N_637,N_559,N_595);
nand U638 (N_638,N_592,N_530);
and U639 (N_639,N_566,N_576);
and U640 (N_640,N_593,N_562);
xnor U641 (N_641,N_548,N_557);
nand U642 (N_642,N_564,N_525);
nor U643 (N_643,N_534,N_525);
nand U644 (N_644,N_569,N_572);
nor U645 (N_645,N_588,N_551);
and U646 (N_646,N_531,N_554);
nor U647 (N_647,N_595,N_564);
and U648 (N_648,N_588,N_531);
nor U649 (N_649,N_572,N_593);
nand U650 (N_650,N_543,N_552);
nand U651 (N_651,N_585,N_551);
and U652 (N_652,N_539,N_593);
or U653 (N_653,N_541,N_583);
nor U654 (N_654,N_555,N_590);
nand U655 (N_655,N_550,N_551);
and U656 (N_656,N_564,N_570);
nand U657 (N_657,N_560,N_556);
nand U658 (N_658,N_534,N_538);
nand U659 (N_659,N_562,N_594);
or U660 (N_660,N_537,N_565);
nand U661 (N_661,N_562,N_537);
nor U662 (N_662,N_545,N_532);
or U663 (N_663,N_577,N_535);
nor U664 (N_664,N_592,N_587);
nand U665 (N_665,N_572,N_548);
or U666 (N_666,N_576,N_575);
nand U667 (N_667,N_558,N_582);
nor U668 (N_668,N_555,N_546);
or U669 (N_669,N_595,N_542);
or U670 (N_670,N_580,N_576);
or U671 (N_671,N_569,N_549);
nor U672 (N_672,N_587,N_583);
nand U673 (N_673,N_598,N_559);
nor U674 (N_674,N_531,N_593);
and U675 (N_675,N_674,N_641);
nand U676 (N_676,N_623,N_630);
and U677 (N_677,N_661,N_655);
and U678 (N_678,N_657,N_658);
nor U679 (N_679,N_669,N_637);
or U680 (N_680,N_666,N_645);
nor U681 (N_681,N_607,N_644);
nand U682 (N_682,N_602,N_673);
or U683 (N_683,N_609,N_651);
nor U684 (N_684,N_634,N_670);
and U685 (N_685,N_653,N_610);
and U686 (N_686,N_652,N_663);
nand U687 (N_687,N_659,N_668);
nand U688 (N_688,N_646,N_631);
or U689 (N_689,N_617,N_672);
or U690 (N_690,N_662,N_648);
nor U691 (N_691,N_611,N_643);
nand U692 (N_692,N_627,N_603);
nand U693 (N_693,N_650,N_660);
nand U694 (N_694,N_638,N_640);
or U695 (N_695,N_622,N_635);
or U696 (N_696,N_605,N_601);
nor U697 (N_697,N_616,N_619);
nor U698 (N_698,N_612,N_649);
nor U699 (N_699,N_633,N_642);
nor U700 (N_700,N_656,N_632);
nor U701 (N_701,N_606,N_620);
nand U702 (N_702,N_608,N_665);
nand U703 (N_703,N_671,N_621);
nand U704 (N_704,N_628,N_639);
and U705 (N_705,N_654,N_647);
nor U706 (N_706,N_664,N_667);
or U707 (N_707,N_629,N_626);
and U708 (N_708,N_614,N_625);
nor U709 (N_709,N_615,N_618);
or U710 (N_710,N_600,N_624);
or U711 (N_711,N_604,N_636);
and U712 (N_712,N_613,N_620);
nand U713 (N_713,N_639,N_640);
nand U714 (N_714,N_665,N_663);
nand U715 (N_715,N_633,N_649);
and U716 (N_716,N_612,N_607);
nor U717 (N_717,N_662,N_605);
or U718 (N_718,N_603,N_623);
nor U719 (N_719,N_635,N_655);
or U720 (N_720,N_610,N_658);
and U721 (N_721,N_659,N_635);
nor U722 (N_722,N_642,N_660);
and U723 (N_723,N_632,N_634);
or U724 (N_724,N_629,N_612);
nor U725 (N_725,N_608,N_672);
nand U726 (N_726,N_656,N_635);
nor U727 (N_727,N_625,N_646);
or U728 (N_728,N_632,N_624);
and U729 (N_729,N_660,N_674);
or U730 (N_730,N_648,N_604);
nor U731 (N_731,N_651,N_670);
or U732 (N_732,N_636,N_613);
nor U733 (N_733,N_606,N_624);
nand U734 (N_734,N_635,N_633);
nor U735 (N_735,N_661,N_667);
or U736 (N_736,N_658,N_642);
or U737 (N_737,N_621,N_650);
nor U738 (N_738,N_672,N_612);
nand U739 (N_739,N_637,N_602);
nand U740 (N_740,N_633,N_660);
nor U741 (N_741,N_609,N_605);
nand U742 (N_742,N_603,N_638);
xor U743 (N_743,N_632,N_665);
nor U744 (N_744,N_621,N_641);
and U745 (N_745,N_668,N_633);
and U746 (N_746,N_672,N_671);
nand U747 (N_747,N_645,N_642);
nand U748 (N_748,N_648,N_664);
nand U749 (N_749,N_650,N_600);
or U750 (N_750,N_693,N_699);
or U751 (N_751,N_726,N_747);
and U752 (N_752,N_714,N_695);
nand U753 (N_753,N_731,N_701);
nand U754 (N_754,N_703,N_724);
nand U755 (N_755,N_677,N_690);
or U756 (N_756,N_702,N_738);
or U757 (N_757,N_676,N_709);
and U758 (N_758,N_733,N_692);
nand U759 (N_759,N_749,N_687);
nor U760 (N_760,N_694,N_711);
nor U761 (N_761,N_725,N_739);
or U762 (N_762,N_715,N_685);
and U763 (N_763,N_740,N_743);
or U764 (N_764,N_741,N_704);
and U765 (N_765,N_727,N_688);
nand U766 (N_766,N_697,N_730);
nand U767 (N_767,N_718,N_728);
or U768 (N_768,N_732,N_720);
nor U769 (N_769,N_700,N_713);
nor U770 (N_770,N_746,N_680);
nor U771 (N_771,N_722,N_708);
nor U772 (N_772,N_742,N_748);
or U773 (N_773,N_675,N_723);
and U774 (N_774,N_716,N_705);
or U775 (N_775,N_734,N_736);
and U776 (N_776,N_737,N_744);
nand U777 (N_777,N_691,N_735);
and U778 (N_778,N_707,N_717);
nor U779 (N_779,N_721,N_689);
nor U780 (N_780,N_682,N_683);
nand U781 (N_781,N_706,N_678);
nand U782 (N_782,N_719,N_710);
nor U783 (N_783,N_698,N_679);
nor U784 (N_784,N_745,N_681);
and U785 (N_785,N_712,N_686);
nor U786 (N_786,N_729,N_696);
and U787 (N_787,N_684,N_715);
or U788 (N_788,N_704,N_707);
and U789 (N_789,N_694,N_678);
nor U790 (N_790,N_682,N_734);
nor U791 (N_791,N_739,N_740);
or U792 (N_792,N_744,N_691);
or U793 (N_793,N_706,N_698);
nor U794 (N_794,N_706,N_701);
or U795 (N_795,N_741,N_720);
and U796 (N_796,N_695,N_725);
or U797 (N_797,N_743,N_701);
nand U798 (N_798,N_727,N_746);
and U799 (N_799,N_680,N_723);
nand U800 (N_800,N_739,N_688);
and U801 (N_801,N_687,N_726);
nand U802 (N_802,N_720,N_701);
and U803 (N_803,N_696,N_740);
and U804 (N_804,N_742,N_712);
nand U805 (N_805,N_731,N_748);
nand U806 (N_806,N_690,N_679);
or U807 (N_807,N_675,N_722);
or U808 (N_808,N_720,N_736);
nor U809 (N_809,N_692,N_736);
nand U810 (N_810,N_703,N_739);
nand U811 (N_811,N_691,N_697);
and U812 (N_812,N_678,N_734);
or U813 (N_813,N_677,N_717);
or U814 (N_814,N_737,N_678);
or U815 (N_815,N_693,N_718);
or U816 (N_816,N_725,N_696);
or U817 (N_817,N_721,N_691);
nand U818 (N_818,N_717,N_748);
nor U819 (N_819,N_744,N_701);
nor U820 (N_820,N_685,N_704);
nor U821 (N_821,N_698,N_719);
nor U822 (N_822,N_733,N_747);
nor U823 (N_823,N_747,N_713);
nor U824 (N_824,N_711,N_697);
or U825 (N_825,N_776,N_794);
nor U826 (N_826,N_767,N_792);
or U827 (N_827,N_779,N_785);
and U828 (N_828,N_803,N_778);
or U829 (N_829,N_798,N_789);
and U830 (N_830,N_805,N_791);
or U831 (N_831,N_796,N_770);
nor U832 (N_832,N_799,N_758);
nand U833 (N_833,N_808,N_815);
nor U834 (N_834,N_802,N_809);
nand U835 (N_835,N_800,N_810);
nor U836 (N_836,N_823,N_786);
nor U837 (N_837,N_817,N_795);
or U838 (N_838,N_766,N_821);
or U839 (N_839,N_757,N_813);
or U840 (N_840,N_750,N_793);
or U841 (N_841,N_752,N_782);
nor U842 (N_842,N_819,N_764);
nand U843 (N_843,N_822,N_788);
and U844 (N_844,N_760,N_751);
nand U845 (N_845,N_806,N_787);
and U846 (N_846,N_765,N_804);
and U847 (N_847,N_820,N_816);
or U848 (N_848,N_761,N_768);
nand U849 (N_849,N_783,N_773);
and U850 (N_850,N_762,N_771);
and U851 (N_851,N_801,N_807);
nor U852 (N_852,N_814,N_769);
nand U853 (N_853,N_781,N_811);
nand U854 (N_854,N_784,N_759);
nand U855 (N_855,N_790,N_775);
nand U856 (N_856,N_763,N_754);
or U857 (N_857,N_774,N_755);
or U858 (N_858,N_812,N_780);
and U859 (N_859,N_824,N_772);
and U860 (N_860,N_753,N_777);
or U861 (N_861,N_756,N_818);
and U862 (N_862,N_797,N_766);
or U863 (N_863,N_761,N_812);
or U864 (N_864,N_815,N_792);
or U865 (N_865,N_816,N_813);
and U866 (N_866,N_811,N_809);
or U867 (N_867,N_821,N_815);
nand U868 (N_868,N_794,N_758);
nor U869 (N_869,N_759,N_755);
nor U870 (N_870,N_780,N_757);
nor U871 (N_871,N_773,N_758);
nor U872 (N_872,N_766,N_779);
nand U873 (N_873,N_791,N_778);
nand U874 (N_874,N_788,N_753);
nand U875 (N_875,N_787,N_778);
nand U876 (N_876,N_799,N_818);
or U877 (N_877,N_769,N_792);
and U878 (N_878,N_756,N_809);
or U879 (N_879,N_780,N_753);
and U880 (N_880,N_817,N_768);
and U881 (N_881,N_762,N_822);
nand U882 (N_882,N_807,N_809);
and U883 (N_883,N_781,N_753);
nand U884 (N_884,N_815,N_779);
nand U885 (N_885,N_778,N_764);
nor U886 (N_886,N_765,N_758);
nand U887 (N_887,N_759,N_758);
nor U888 (N_888,N_797,N_820);
nand U889 (N_889,N_783,N_764);
nand U890 (N_890,N_799,N_812);
nor U891 (N_891,N_764,N_801);
or U892 (N_892,N_808,N_797);
nand U893 (N_893,N_814,N_815);
nand U894 (N_894,N_794,N_766);
or U895 (N_895,N_807,N_768);
nand U896 (N_896,N_757,N_788);
xnor U897 (N_897,N_808,N_803);
nor U898 (N_898,N_770,N_793);
nor U899 (N_899,N_768,N_765);
nor U900 (N_900,N_869,N_889);
and U901 (N_901,N_856,N_881);
nand U902 (N_902,N_836,N_842);
nor U903 (N_903,N_826,N_868);
nand U904 (N_904,N_897,N_832);
or U905 (N_905,N_892,N_859);
and U906 (N_906,N_893,N_866);
nand U907 (N_907,N_840,N_885);
nor U908 (N_908,N_841,N_849);
nor U909 (N_909,N_828,N_872);
or U910 (N_910,N_888,N_862);
nand U911 (N_911,N_830,N_879);
and U912 (N_912,N_878,N_837);
nand U913 (N_913,N_898,N_851);
and U914 (N_914,N_899,N_839);
or U915 (N_915,N_876,N_834);
nor U916 (N_916,N_867,N_844);
and U917 (N_917,N_863,N_861);
nor U918 (N_918,N_838,N_835);
and U919 (N_919,N_843,N_890);
or U920 (N_920,N_895,N_860);
nand U921 (N_921,N_825,N_833);
or U922 (N_922,N_871,N_854);
nor U923 (N_923,N_829,N_846);
or U924 (N_924,N_847,N_874);
xnor U925 (N_925,N_886,N_896);
and U926 (N_926,N_848,N_865);
nand U927 (N_927,N_852,N_883);
nor U928 (N_928,N_894,N_870);
and U929 (N_929,N_875,N_853);
or U930 (N_930,N_850,N_884);
nor U931 (N_931,N_831,N_877);
and U932 (N_932,N_858,N_855);
and U933 (N_933,N_887,N_857);
nand U934 (N_934,N_827,N_880);
and U935 (N_935,N_882,N_845);
and U936 (N_936,N_891,N_873);
and U937 (N_937,N_864,N_826);
nor U938 (N_938,N_837,N_845);
nand U939 (N_939,N_889,N_858);
nand U940 (N_940,N_835,N_832);
nand U941 (N_941,N_845,N_835);
nor U942 (N_942,N_830,N_827);
nor U943 (N_943,N_832,N_869);
nand U944 (N_944,N_865,N_847);
and U945 (N_945,N_829,N_888);
nor U946 (N_946,N_879,N_825);
nand U947 (N_947,N_835,N_834);
nor U948 (N_948,N_896,N_861);
nor U949 (N_949,N_889,N_841);
nand U950 (N_950,N_888,N_851);
nor U951 (N_951,N_892,N_862);
nor U952 (N_952,N_842,N_862);
and U953 (N_953,N_885,N_842);
nor U954 (N_954,N_882,N_877);
nor U955 (N_955,N_836,N_872);
nor U956 (N_956,N_841,N_851);
nand U957 (N_957,N_832,N_834);
or U958 (N_958,N_827,N_856);
nor U959 (N_959,N_894,N_832);
nor U960 (N_960,N_868,N_878);
or U961 (N_961,N_888,N_866);
or U962 (N_962,N_895,N_868);
nor U963 (N_963,N_848,N_857);
nand U964 (N_964,N_874,N_890);
and U965 (N_965,N_868,N_850);
nor U966 (N_966,N_829,N_884);
nand U967 (N_967,N_834,N_846);
and U968 (N_968,N_860,N_865);
or U969 (N_969,N_887,N_843);
and U970 (N_970,N_831,N_845);
and U971 (N_971,N_890,N_832);
or U972 (N_972,N_826,N_892);
nand U973 (N_973,N_870,N_885);
nand U974 (N_974,N_831,N_826);
or U975 (N_975,N_927,N_952);
or U976 (N_976,N_957,N_972);
nand U977 (N_977,N_919,N_963);
or U978 (N_978,N_907,N_964);
and U979 (N_979,N_910,N_956);
nand U980 (N_980,N_913,N_949);
and U981 (N_981,N_925,N_928);
nand U982 (N_982,N_936,N_933);
nand U983 (N_983,N_905,N_923);
and U984 (N_984,N_948,N_940);
and U985 (N_985,N_945,N_903);
nor U986 (N_986,N_924,N_902);
or U987 (N_987,N_962,N_951);
or U988 (N_988,N_926,N_904);
and U989 (N_989,N_973,N_953);
nor U990 (N_990,N_942,N_974);
or U991 (N_991,N_922,N_970);
nor U992 (N_992,N_965,N_938);
nand U993 (N_993,N_920,N_954);
and U994 (N_994,N_930,N_932);
or U995 (N_995,N_929,N_947);
or U996 (N_996,N_916,N_935);
and U997 (N_997,N_909,N_914);
nor U998 (N_998,N_950,N_968);
or U999 (N_999,N_934,N_921);
nor U1000 (N_1000,N_955,N_967);
or U1001 (N_1001,N_900,N_946);
and U1002 (N_1002,N_918,N_959);
nor U1003 (N_1003,N_906,N_915);
nor U1004 (N_1004,N_971,N_944);
nand U1005 (N_1005,N_911,N_943);
or U1006 (N_1006,N_908,N_939);
nand U1007 (N_1007,N_969,N_931);
nand U1008 (N_1008,N_960,N_912);
or U1009 (N_1009,N_901,N_961);
nor U1010 (N_1010,N_917,N_966);
nor U1011 (N_1011,N_937,N_941);
nand U1012 (N_1012,N_958,N_954);
or U1013 (N_1013,N_942,N_907);
and U1014 (N_1014,N_903,N_941);
nand U1015 (N_1015,N_916,N_948);
nor U1016 (N_1016,N_943,N_970);
nor U1017 (N_1017,N_931,N_901);
and U1018 (N_1018,N_943,N_923);
or U1019 (N_1019,N_938,N_957);
or U1020 (N_1020,N_907,N_952);
or U1021 (N_1021,N_953,N_933);
nor U1022 (N_1022,N_957,N_908);
and U1023 (N_1023,N_958,N_929);
nor U1024 (N_1024,N_970,N_927);
nor U1025 (N_1025,N_952,N_974);
or U1026 (N_1026,N_968,N_913);
nor U1027 (N_1027,N_973,N_935);
or U1028 (N_1028,N_915,N_944);
and U1029 (N_1029,N_954,N_950);
or U1030 (N_1030,N_966,N_920);
nor U1031 (N_1031,N_932,N_921);
and U1032 (N_1032,N_970,N_957);
and U1033 (N_1033,N_940,N_906);
nand U1034 (N_1034,N_962,N_939);
or U1035 (N_1035,N_938,N_942);
nor U1036 (N_1036,N_943,N_909);
nor U1037 (N_1037,N_914,N_940);
and U1038 (N_1038,N_948,N_902);
and U1039 (N_1039,N_933,N_955);
nor U1040 (N_1040,N_966,N_954);
and U1041 (N_1041,N_971,N_973);
and U1042 (N_1042,N_901,N_922);
or U1043 (N_1043,N_947,N_907);
and U1044 (N_1044,N_958,N_904);
or U1045 (N_1045,N_930,N_973);
xor U1046 (N_1046,N_931,N_913);
nor U1047 (N_1047,N_971,N_918);
nand U1048 (N_1048,N_921,N_947);
nand U1049 (N_1049,N_966,N_928);
nand U1050 (N_1050,N_985,N_981);
nand U1051 (N_1051,N_1007,N_1013);
nor U1052 (N_1052,N_1029,N_1024);
or U1053 (N_1053,N_1048,N_1044);
or U1054 (N_1054,N_1021,N_1036);
and U1055 (N_1055,N_986,N_1003);
or U1056 (N_1056,N_1010,N_1006);
or U1057 (N_1057,N_983,N_978);
nor U1058 (N_1058,N_977,N_1042);
and U1059 (N_1059,N_1041,N_1046);
nand U1060 (N_1060,N_1014,N_1035);
or U1061 (N_1061,N_1017,N_1025);
or U1062 (N_1062,N_1004,N_979);
and U1063 (N_1063,N_980,N_1000);
nor U1064 (N_1064,N_1039,N_1027);
or U1065 (N_1065,N_999,N_1028);
and U1066 (N_1066,N_1032,N_997);
nand U1067 (N_1067,N_992,N_1008);
nor U1068 (N_1068,N_976,N_1020);
nand U1069 (N_1069,N_1043,N_1030);
and U1070 (N_1070,N_1040,N_1018);
or U1071 (N_1071,N_1019,N_998);
and U1072 (N_1072,N_1012,N_975);
or U1073 (N_1073,N_996,N_1011);
nand U1074 (N_1074,N_1002,N_1009);
and U1075 (N_1075,N_993,N_1005);
nor U1076 (N_1076,N_995,N_994);
nor U1077 (N_1077,N_1049,N_1001);
or U1078 (N_1078,N_1038,N_990);
nor U1079 (N_1079,N_1023,N_1047);
or U1080 (N_1080,N_987,N_1022);
nor U1081 (N_1081,N_989,N_982);
or U1082 (N_1082,N_1026,N_1045);
or U1083 (N_1083,N_1016,N_988);
and U1084 (N_1084,N_1034,N_1033);
nand U1085 (N_1085,N_1031,N_984);
and U1086 (N_1086,N_991,N_1037);
and U1087 (N_1087,N_1015,N_1044);
nor U1088 (N_1088,N_1040,N_1029);
nand U1089 (N_1089,N_993,N_1049);
nor U1090 (N_1090,N_1015,N_980);
nand U1091 (N_1091,N_997,N_986);
nand U1092 (N_1092,N_1028,N_1022);
nand U1093 (N_1093,N_998,N_991);
or U1094 (N_1094,N_1041,N_977);
nand U1095 (N_1095,N_996,N_982);
or U1096 (N_1096,N_1018,N_1042);
and U1097 (N_1097,N_1029,N_1018);
nand U1098 (N_1098,N_1029,N_1026);
and U1099 (N_1099,N_1018,N_978);
or U1100 (N_1100,N_1008,N_983);
or U1101 (N_1101,N_998,N_1029);
nand U1102 (N_1102,N_1030,N_1012);
nor U1103 (N_1103,N_1019,N_1023);
and U1104 (N_1104,N_1006,N_1024);
nand U1105 (N_1105,N_990,N_1007);
nand U1106 (N_1106,N_978,N_1048);
or U1107 (N_1107,N_1013,N_981);
and U1108 (N_1108,N_1037,N_983);
nor U1109 (N_1109,N_1044,N_993);
or U1110 (N_1110,N_988,N_990);
nand U1111 (N_1111,N_980,N_1009);
nor U1112 (N_1112,N_1019,N_1005);
nor U1113 (N_1113,N_1034,N_1035);
and U1114 (N_1114,N_983,N_1026);
nor U1115 (N_1115,N_1037,N_980);
nor U1116 (N_1116,N_989,N_1013);
or U1117 (N_1117,N_1010,N_978);
and U1118 (N_1118,N_1035,N_997);
nand U1119 (N_1119,N_1005,N_1032);
and U1120 (N_1120,N_1042,N_1002);
or U1121 (N_1121,N_982,N_1033);
and U1122 (N_1122,N_995,N_993);
nor U1123 (N_1123,N_1019,N_1027);
and U1124 (N_1124,N_1015,N_979);
and U1125 (N_1125,N_1088,N_1121);
nor U1126 (N_1126,N_1076,N_1073);
and U1127 (N_1127,N_1052,N_1075);
nor U1128 (N_1128,N_1069,N_1085);
nand U1129 (N_1129,N_1117,N_1053);
and U1130 (N_1130,N_1093,N_1072);
nor U1131 (N_1131,N_1054,N_1098);
nand U1132 (N_1132,N_1087,N_1084);
and U1133 (N_1133,N_1086,N_1094);
and U1134 (N_1134,N_1119,N_1120);
or U1135 (N_1135,N_1077,N_1092);
or U1136 (N_1136,N_1065,N_1109);
nand U1137 (N_1137,N_1070,N_1114);
nand U1138 (N_1138,N_1071,N_1057);
and U1139 (N_1139,N_1083,N_1108);
nand U1140 (N_1140,N_1097,N_1079);
nor U1141 (N_1141,N_1103,N_1116);
nand U1142 (N_1142,N_1105,N_1111);
or U1143 (N_1143,N_1110,N_1062);
or U1144 (N_1144,N_1078,N_1080);
or U1145 (N_1145,N_1064,N_1100);
or U1146 (N_1146,N_1060,N_1115);
or U1147 (N_1147,N_1056,N_1113);
nand U1148 (N_1148,N_1099,N_1082);
nor U1149 (N_1149,N_1051,N_1104);
or U1150 (N_1150,N_1081,N_1095);
nor U1151 (N_1151,N_1063,N_1096);
nand U1152 (N_1152,N_1068,N_1123);
nor U1153 (N_1153,N_1118,N_1107);
nand U1154 (N_1154,N_1122,N_1055);
or U1155 (N_1155,N_1050,N_1102);
nand U1156 (N_1156,N_1112,N_1124);
and U1157 (N_1157,N_1074,N_1066);
nor U1158 (N_1158,N_1106,N_1067);
or U1159 (N_1159,N_1059,N_1089);
and U1160 (N_1160,N_1101,N_1090);
nand U1161 (N_1161,N_1091,N_1061);
or U1162 (N_1162,N_1058,N_1069);
nand U1163 (N_1163,N_1105,N_1091);
or U1164 (N_1164,N_1079,N_1084);
and U1165 (N_1165,N_1059,N_1072);
nand U1166 (N_1166,N_1064,N_1071);
and U1167 (N_1167,N_1086,N_1123);
nor U1168 (N_1168,N_1057,N_1062);
and U1169 (N_1169,N_1071,N_1062);
nor U1170 (N_1170,N_1090,N_1096);
nor U1171 (N_1171,N_1071,N_1086);
nand U1172 (N_1172,N_1108,N_1050);
nand U1173 (N_1173,N_1087,N_1109);
nand U1174 (N_1174,N_1082,N_1074);
nor U1175 (N_1175,N_1055,N_1097);
nor U1176 (N_1176,N_1104,N_1115);
nand U1177 (N_1177,N_1089,N_1095);
nand U1178 (N_1178,N_1116,N_1053);
or U1179 (N_1179,N_1121,N_1055);
xor U1180 (N_1180,N_1063,N_1111);
nor U1181 (N_1181,N_1056,N_1072);
and U1182 (N_1182,N_1075,N_1072);
nor U1183 (N_1183,N_1077,N_1087);
nand U1184 (N_1184,N_1096,N_1080);
nor U1185 (N_1185,N_1078,N_1079);
nand U1186 (N_1186,N_1064,N_1106);
or U1187 (N_1187,N_1064,N_1092);
and U1188 (N_1188,N_1072,N_1070);
nor U1189 (N_1189,N_1093,N_1095);
nand U1190 (N_1190,N_1115,N_1112);
or U1191 (N_1191,N_1067,N_1069);
or U1192 (N_1192,N_1095,N_1078);
nor U1193 (N_1193,N_1121,N_1066);
and U1194 (N_1194,N_1070,N_1058);
nand U1195 (N_1195,N_1091,N_1080);
or U1196 (N_1196,N_1072,N_1103);
or U1197 (N_1197,N_1061,N_1058);
nor U1198 (N_1198,N_1070,N_1122);
or U1199 (N_1199,N_1117,N_1076);
nand U1200 (N_1200,N_1183,N_1137);
and U1201 (N_1201,N_1188,N_1155);
and U1202 (N_1202,N_1184,N_1161);
nand U1203 (N_1203,N_1152,N_1169);
nand U1204 (N_1204,N_1174,N_1164);
and U1205 (N_1205,N_1172,N_1159);
or U1206 (N_1206,N_1129,N_1194);
nand U1207 (N_1207,N_1135,N_1178);
nor U1208 (N_1208,N_1181,N_1142);
or U1209 (N_1209,N_1197,N_1154);
and U1210 (N_1210,N_1145,N_1146);
and U1211 (N_1211,N_1198,N_1147);
nand U1212 (N_1212,N_1156,N_1132);
and U1213 (N_1213,N_1173,N_1162);
or U1214 (N_1214,N_1150,N_1157);
or U1215 (N_1215,N_1141,N_1185);
nand U1216 (N_1216,N_1138,N_1191);
and U1217 (N_1217,N_1175,N_1126);
nor U1218 (N_1218,N_1167,N_1131);
xor U1219 (N_1219,N_1176,N_1158);
or U1220 (N_1220,N_1151,N_1140);
or U1221 (N_1221,N_1195,N_1179);
and U1222 (N_1222,N_1163,N_1166);
nor U1223 (N_1223,N_1144,N_1165);
or U1224 (N_1224,N_1186,N_1125);
nand U1225 (N_1225,N_1170,N_1192);
or U1226 (N_1226,N_1128,N_1182);
or U1227 (N_1227,N_1133,N_1153);
nand U1228 (N_1228,N_1130,N_1149);
nand U1229 (N_1229,N_1168,N_1171);
and U1230 (N_1230,N_1143,N_1134);
nand U1231 (N_1231,N_1127,N_1148);
and U1232 (N_1232,N_1190,N_1160);
and U1233 (N_1233,N_1177,N_1136);
and U1234 (N_1234,N_1189,N_1199);
nand U1235 (N_1235,N_1193,N_1139);
and U1236 (N_1236,N_1196,N_1187);
nor U1237 (N_1237,N_1180,N_1156);
or U1238 (N_1238,N_1184,N_1198);
nand U1239 (N_1239,N_1192,N_1171);
and U1240 (N_1240,N_1189,N_1157);
nor U1241 (N_1241,N_1156,N_1198);
or U1242 (N_1242,N_1191,N_1190);
or U1243 (N_1243,N_1125,N_1197);
or U1244 (N_1244,N_1142,N_1136);
nand U1245 (N_1245,N_1158,N_1152);
nor U1246 (N_1246,N_1193,N_1164);
or U1247 (N_1247,N_1164,N_1173);
or U1248 (N_1248,N_1139,N_1127);
nor U1249 (N_1249,N_1149,N_1181);
and U1250 (N_1250,N_1179,N_1166);
and U1251 (N_1251,N_1172,N_1158);
nand U1252 (N_1252,N_1136,N_1176);
nand U1253 (N_1253,N_1175,N_1180);
xor U1254 (N_1254,N_1183,N_1143);
nor U1255 (N_1255,N_1126,N_1164);
or U1256 (N_1256,N_1142,N_1126);
or U1257 (N_1257,N_1168,N_1144);
or U1258 (N_1258,N_1169,N_1179);
nand U1259 (N_1259,N_1129,N_1199);
and U1260 (N_1260,N_1184,N_1199);
and U1261 (N_1261,N_1166,N_1149);
nor U1262 (N_1262,N_1194,N_1142);
nand U1263 (N_1263,N_1159,N_1170);
and U1264 (N_1264,N_1159,N_1175);
nor U1265 (N_1265,N_1181,N_1130);
nand U1266 (N_1266,N_1169,N_1142);
nand U1267 (N_1267,N_1165,N_1170);
or U1268 (N_1268,N_1173,N_1148);
and U1269 (N_1269,N_1181,N_1131);
nor U1270 (N_1270,N_1185,N_1178);
nor U1271 (N_1271,N_1141,N_1192);
nor U1272 (N_1272,N_1197,N_1186);
nor U1273 (N_1273,N_1153,N_1196);
nor U1274 (N_1274,N_1153,N_1184);
and U1275 (N_1275,N_1206,N_1243);
or U1276 (N_1276,N_1266,N_1257);
nand U1277 (N_1277,N_1250,N_1268);
or U1278 (N_1278,N_1252,N_1225);
and U1279 (N_1279,N_1271,N_1203);
or U1280 (N_1280,N_1222,N_1246);
nor U1281 (N_1281,N_1213,N_1220);
nor U1282 (N_1282,N_1239,N_1260);
nand U1283 (N_1283,N_1200,N_1207);
or U1284 (N_1284,N_1241,N_1212);
xnor U1285 (N_1285,N_1272,N_1269);
or U1286 (N_1286,N_1228,N_1262);
nand U1287 (N_1287,N_1216,N_1255);
or U1288 (N_1288,N_1267,N_1215);
nand U1289 (N_1289,N_1232,N_1273);
nor U1290 (N_1290,N_1259,N_1251);
nor U1291 (N_1291,N_1261,N_1234);
nor U1292 (N_1292,N_1211,N_1221);
nor U1293 (N_1293,N_1202,N_1235);
and U1294 (N_1294,N_1238,N_1227);
nand U1295 (N_1295,N_1253,N_1242);
and U1296 (N_1296,N_1245,N_1204);
nor U1297 (N_1297,N_1258,N_1264);
and U1298 (N_1298,N_1263,N_1201);
or U1299 (N_1299,N_1240,N_1237);
or U1300 (N_1300,N_1248,N_1270);
nand U1301 (N_1301,N_1229,N_1224);
nor U1302 (N_1302,N_1209,N_1254);
nand U1303 (N_1303,N_1233,N_1244);
nand U1304 (N_1304,N_1217,N_1214);
and U1305 (N_1305,N_1256,N_1274);
and U1306 (N_1306,N_1205,N_1223);
or U1307 (N_1307,N_1219,N_1208);
or U1308 (N_1308,N_1249,N_1236);
nor U1309 (N_1309,N_1265,N_1226);
and U1310 (N_1310,N_1230,N_1218);
nand U1311 (N_1311,N_1247,N_1210);
and U1312 (N_1312,N_1231,N_1230);
nor U1313 (N_1313,N_1258,N_1224);
and U1314 (N_1314,N_1271,N_1243);
xnor U1315 (N_1315,N_1211,N_1237);
or U1316 (N_1316,N_1238,N_1249);
and U1317 (N_1317,N_1215,N_1212);
nor U1318 (N_1318,N_1262,N_1252);
nand U1319 (N_1319,N_1251,N_1270);
nand U1320 (N_1320,N_1262,N_1226);
or U1321 (N_1321,N_1264,N_1251);
and U1322 (N_1322,N_1251,N_1239);
nor U1323 (N_1323,N_1219,N_1238);
and U1324 (N_1324,N_1251,N_1241);
nor U1325 (N_1325,N_1265,N_1215);
and U1326 (N_1326,N_1214,N_1235);
nor U1327 (N_1327,N_1234,N_1211);
nor U1328 (N_1328,N_1268,N_1222);
or U1329 (N_1329,N_1221,N_1235);
nand U1330 (N_1330,N_1264,N_1212);
nand U1331 (N_1331,N_1245,N_1270);
or U1332 (N_1332,N_1264,N_1225);
nor U1333 (N_1333,N_1230,N_1245);
nor U1334 (N_1334,N_1213,N_1274);
nor U1335 (N_1335,N_1257,N_1270);
and U1336 (N_1336,N_1259,N_1230);
nand U1337 (N_1337,N_1265,N_1232);
or U1338 (N_1338,N_1225,N_1202);
xor U1339 (N_1339,N_1221,N_1238);
and U1340 (N_1340,N_1252,N_1224);
or U1341 (N_1341,N_1241,N_1257);
and U1342 (N_1342,N_1257,N_1212);
nand U1343 (N_1343,N_1216,N_1205);
or U1344 (N_1344,N_1204,N_1254);
nand U1345 (N_1345,N_1210,N_1274);
or U1346 (N_1346,N_1264,N_1270);
nor U1347 (N_1347,N_1256,N_1217);
nand U1348 (N_1348,N_1239,N_1225);
and U1349 (N_1349,N_1213,N_1202);
nor U1350 (N_1350,N_1291,N_1275);
nor U1351 (N_1351,N_1337,N_1300);
or U1352 (N_1352,N_1289,N_1285);
nand U1353 (N_1353,N_1284,N_1320);
nor U1354 (N_1354,N_1345,N_1328);
xor U1355 (N_1355,N_1304,N_1347);
nand U1356 (N_1356,N_1343,N_1287);
nand U1357 (N_1357,N_1313,N_1305);
and U1358 (N_1358,N_1292,N_1293);
and U1359 (N_1359,N_1340,N_1331);
or U1360 (N_1360,N_1312,N_1295);
nand U1361 (N_1361,N_1298,N_1333);
and U1362 (N_1362,N_1286,N_1318);
nor U1363 (N_1363,N_1299,N_1311);
nand U1364 (N_1364,N_1277,N_1308);
nor U1365 (N_1365,N_1338,N_1322);
nand U1366 (N_1366,N_1321,N_1294);
nand U1367 (N_1367,N_1342,N_1329);
or U1368 (N_1368,N_1335,N_1302);
and U1369 (N_1369,N_1290,N_1319);
and U1370 (N_1370,N_1309,N_1327);
or U1371 (N_1371,N_1326,N_1334);
or U1372 (N_1372,N_1301,N_1324);
or U1373 (N_1373,N_1288,N_1303);
and U1374 (N_1374,N_1283,N_1296);
nor U1375 (N_1375,N_1307,N_1348);
and U1376 (N_1376,N_1317,N_1276);
nand U1377 (N_1377,N_1344,N_1323);
nand U1378 (N_1378,N_1315,N_1330);
nor U1379 (N_1379,N_1306,N_1281);
nor U1380 (N_1380,N_1341,N_1282);
and U1381 (N_1381,N_1325,N_1314);
nor U1382 (N_1382,N_1346,N_1332);
nand U1383 (N_1383,N_1310,N_1349);
nor U1384 (N_1384,N_1339,N_1316);
and U1385 (N_1385,N_1297,N_1278);
or U1386 (N_1386,N_1280,N_1279);
nor U1387 (N_1387,N_1336,N_1290);
nor U1388 (N_1388,N_1319,N_1286);
nand U1389 (N_1389,N_1338,N_1325);
nand U1390 (N_1390,N_1346,N_1293);
or U1391 (N_1391,N_1331,N_1283);
and U1392 (N_1392,N_1348,N_1280);
nor U1393 (N_1393,N_1314,N_1280);
nand U1394 (N_1394,N_1318,N_1289);
or U1395 (N_1395,N_1292,N_1334);
or U1396 (N_1396,N_1334,N_1316);
nand U1397 (N_1397,N_1294,N_1340);
or U1398 (N_1398,N_1323,N_1341);
nor U1399 (N_1399,N_1337,N_1348);
and U1400 (N_1400,N_1275,N_1330);
or U1401 (N_1401,N_1308,N_1347);
or U1402 (N_1402,N_1346,N_1311);
nand U1403 (N_1403,N_1291,N_1313);
nand U1404 (N_1404,N_1338,N_1290);
or U1405 (N_1405,N_1349,N_1312);
nor U1406 (N_1406,N_1285,N_1311);
and U1407 (N_1407,N_1324,N_1314);
and U1408 (N_1408,N_1302,N_1311);
and U1409 (N_1409,N_1342,N_1333);
or U1410 (N_1410,N_1303,N_1330);
nor U1411 (N_1411,N_1336,N_1323);
or U1412 (N_1412,N_1343,N_1298);
or U1413 (N_1413,N_1317,N_1280);
or U1414 (N_1414,N_1287,N_1300);
nand U1415 (N_1415,N_1317,N_1275);
nand U1416 (N_1416,N_1278,N_1308);
nor U1417 (N_1417,N_1280,N_1328);
and U1418 (N_1418,N_1313,N_1323);
or U1419 (N_1419,N_1323,N_1349);
and U1420 (N_1420,N_1280,N_1313);
nor U1421 (N_1421,N_1307,N_1290);
nand U1422 (N_1422,N_1295,N_1332);
nand U1423 (N_1423,N_1275,N_1340);
or U1424 (N_1424,N_1321,N_1318);
nand U1425 (N_1425,N_1378,N_1407);
nor U1426 (N_1426,N_1395,N_1385);
nor U1427 (N_1427,N_1360,N_1383);
nor U1428 (N_1428,N_1406,N_1398);
nand U1429 (N_1429,N_1411,N_1413);
nor U1430 (N_1430,N_1373,N_1379);
and U1431 (N_1431,N_1358,N_1388);
and U1432 (N_1432,N_1387,N_1376);
and U1433 (N_1433,N_1408,N_1423);
xor U1434 (N_1434,N_1389,N_1396);
and U1435 (N_1435,N_1369,N_1390);
or U1436 (N_1436,N_1399,N_1393);
nand U1437 (N_1437,N_1362,N_1424);
or U1438 (N_1438,N_1400,N_1380);
nor U1439 (N_1439,N_1391,N_1386);
and U1440 (N_1440,N_1355,N_1415);
or U1441 (N_1441,N_1374,N_1404);
nor U1442 (N_1442,N_1409,N_1417);
nand U1443 (N_1443,N_1359,N_1416);
nor U1444 (N_1444,N_1392,N_1403);
and U1445 (N_1445,N_1357,N_1377);
nand U1446 (N_1446,N_1382,N_1397);
or U1447 (N_1447,N_1418,N_1366);
nand U1448 (N_1448,N_1410,N_1363);
nand U1449 (N_1449,N_1370,N_1350);
nand U1450 (N_1450,N_1351,N_1401);
nand U1451 (N_1451,N_1394,N_1368);
nand U1452 (N_1452,N_1352,N_1414);
or U1453 (N_1453,N_1375,N_1421);
nand U1454 (N_1454,N_1356,N_1367);
or U1455 (N_1455,N_1420,N_1381);
nor U1456 (N_1456,N_1419,N_1384);
nand U1457 (N_1457,N_1422,N_1371);
nand U1458 (N_1458,N_1402,N_1372);
or U1459 (N_1459,N_1405,N_1353);
and U1460 (N_1460,N_1364,N_1365);
or U1461 (N_1461,N_1354,N_1412);
nand U1462 (N_1462,N_1361,N_1356);
nor U1463 (N_1463,N_1367,N_1399);
nor U1464 (N_1464,N_1424,N_1386);
and U1465 (N_1465,N_1374,N_1414);
or U1466 (N_1466,N_1403,N_1385);
nor U1467 (N_1467,N_1385,N_1363);
nor U1468 (N_1468,N_1389,N_1375);
or U1469 (N_1469,N_1398,N_1409);
or U1470 (N_1470,N_1352,N_1391);
or U1471 (N_1471,N_1374,N_1351);
and U1472 (N_1472,N_1418,N_1356);
or U1473 (N_1473,N_1372,N_1387);
and U1474 (N_1474,N_1355,N_1392);
and U1475 (N_1475,N_1384,N_1407);
nor U1476 (N_1476,N_1382,N_1369);
and U1477 (N_1477,N_1399,N_1385);
or U1478 (N_1478,N_1365,N_1386);
nand U1479 (N_1479,N_1366,N_1362);
xor U1480 (N_1480,N_1350,N_1400);
and U1481 (N_1481,N_1378,N_1397);
nand U1482 (N_1482,N_1394,N_1414);
or U1483 (N_1483,N_1406,N_1360);
or U1484 (N_1484,N_1351,N_1406);
and U1485 (N_1485,N_1410,N_1369);
or U1486 (N_1486,N_1388,N_1411);
and U1487 (N_1487,N_1384,N_1394);
and U1488 (N_1488,N_1387,N_1406);
or U1489 (N_1489,N_1383,N_1390);
and U1490 (N_1490,N_1353,N_1396);
nand U1491 (N_1491,N_1361,N_1351);
nand U1492 (N_1492,N_1409,N_1389);
or U1493 (N_1493,N_1424,N_1374);
nand U1494 (N_1494,N_1406,N_1373);
and U1495 (N_1495,N_1399,N_1392);
nand U1496 (N_1496,N_1411,N_1383);
nor U1497 (N_1497,N_1391,N_1361);
nor U1498 (N_1498,N_1369,N_1381);
nand U1499 (N_1499,N_1379,N_1378);
and U1500 (N_1500,N_1469,N_1455);
or U1501 (N_1501,N_1450,N_1438);
and U1502 (N_1502,N_1464,N_1454);
and U1503 (N_1503,N_1493,N_1427);
nand U1504 (N_1504,N_1472,N_1482);
and U1505 (N_1505,N_1446,N_1485);
nor U1506 (N_1506,N_1480,N_1468);
or U1507 (N_1507,N_1476,N_1494);
and U1508 (N_1508,N_1444,N_1434);
and U1509 (N_1509,N_1498,N_1462);
or U1510 (N_1510,N_1437,N_1445);
nand U1511 (N_1511,N_1457,N_1443);
nand U1512 (N_1512,N_1491,N_1449);
nor U1513 (N_1513,N_1436,N_1432);
nor U1514 (N_1514,N_1435,N_1456);
and U1515 (N_1515,N_1459,N_1448);
or U1516 (N_1516,N_1429,N_1467);
nor U1517 (N_1517,N_1471,N_1473);
nor U1518 (N_1518,N_1496,N_1497);
or U1519 (N_1519,N_1486,N_1484);
and U1520 (N_1520,N_1483,N_1490);
or U1521 (N_1521,N_1458,N_1465);
nor U1522 (N_1522,N_1489,N_1428);
nand U1523 (N_1523,N_1442,N_1431);
nor U1524 (N_1524,N_1433,N_1481);
or U1525 (N_1525,N_1441,N_1477);
or U1526 (N_1526,N_1430,N_1425);
nor U1527 (N_1527,N_1466,N_1487);
nand U1528 (N_1528,N_1426,N_1440);
and U1529 (N_1529,N_1475,N_1461);
and U1530 (N_1530,N_1474,N_1453);
nor U1531 (N_1531,N_1463,N_1460);
and U1532 (N_1532,N_1451,N_1495);
or U1533 (N_1533,N_1478,N_1492);
and U1534 (N_1534,N_1470,N_1452);
nand U1535 (N_1535,N_1499,N_1479);
or U1536 (N_1536,N_1488,N_1439);
or U1537 (N_1537,N_1447,N_1479);
and U1538 (N_1538,N_1482,N_1431);
and U1539 (N_1539,N_1477,N_1426);
or U1540 (N_1540,N_1446,N_1453);
nand U1541 (N_1541,N_1460,N_1497);
and U1542 (N_1542,N_1442,N_1459);
nand U1543 (N_1543,N_1490,N_1494);
or U1544 (N_1544,N_1484,N_1495);
and U1545 (N_1545,N_1493,N_1435);
or U1546 (N_1546,N_1468,N_1488);
nor U1547 (N_1547,N_1473,N_1459);
or U1548 (N_1548,N_1481,N_1429);
nor U1549 (N_1549,N_1498,N_1430);
nor U1550 (N_1550,N_1431,N_1428);
and U1551 (N_1551,N_1449,N_1460);
nand U1552 (N_1552,N_1434,N_1463);
and U1553 (N_1553,N_1466,N_1431);
or U1554 (N_1554,N_1435,N_1438);
and U1555 (N_1555,N_1452,N_1454);
nor U1556 (N_1556,N_1427,N_1435);
nor U1557 (N_1557,N_1467,N_1458);
and U1558 (N_1558,N_1478,N_1447);
nor U1559 (N_1559,N_1499,N_1430);
xor U1560 (N_1560,N_1435,N_1484);
or U1561 (N_1561,N_1456,N_1465);
and U1562 (N_1562,N_1433,N_1434);
nand U1563 (N_1563,N_1452,N_1437);
or U1564 (N_1564,N_1456,N_1496);
and U1565 (N_1565,N_1482,N_1469);
or U1566 (N_1566,N_1485,N_1440);
nand U1567 (N_1567,N_1484,N_1445);
and U1568 (N_1568,N_1443,N_1447);
or U1569 (N_1569,N_1479,N_1489);
nand U1570 (N_1570,N_1432,N_1471);
nor U1571 (N_1571,N_1433,N_1490);
or U1572 (N_1572,N_1444,N_1446);
nand U1573 (N_1573,N_1493,N_1460);
nand U1574 (N_1574,N_1465,N_1478);
and U1575 (N_1575,N_1551,N_1571);
nand U1576 (N_1576,N_1526,N_1547);
nand U1577 (N_1577,N_1554,N_1565);
or U1578 (N_1578,N_1503,N_1518);
nor U1579 (N_1579,N_1573,N_1550);
and U1580 (N_1580,N_1540,N_1556);
nor U1581 (N_1581,N_1562,N_1519);
and U1582 (N_1582,N_1521,N_1515);
nand U1583 (N_1583,N_1555,N_1512);
and U1584 (N_1584,N_1528,N_1536);
and U1585 (N_1585,N_1560,N_1549);
and U1586 (N_1586,N_1531,N_1569);
or U1587 (N_1587,N_1523,N_1516);
or U1588 (N_1588,N_1566,N_1541);
or U1589 (N_1589,N_1552,N_1525);
and U1590 (N_1590,N_1539,N_1535);
or U1591 (N_1591,N_1538,N_1563);
and U1592 (N_1592,N_1530,N_1542);
nand U1593 (N_1593,N_1557,N_1506);
nor U1594 (N_1594,N_1533,N_1534);
nand U1595 (N_1595,N_1559,N_1553);
nand U1596 (N_1596,N_1500,N_1504);
nand U1597 (N_1597,N_1505,N_1510);
nand U1598 (N_1598,N_1514,N_1513);
nor U1599 (N_1599,N_1524,N_1561);
nand U1600 (N_1600,N_1501,N_1532);
or U1601 (N_1601,N_1517,N_1545);
and U1602 (N_1602,N_1570,N_1546);
nor U1603 (N_1603,N_1574,N_1543);
and U1604 (N_1604,N_1572,N_1509);
nor U1605 (N_1605,N_1508,N_1507);
or U1606 (N_1606,N_1502,N_1558);
or U1607 (N_1607,N_1564,N_1537);
nand U1608 (N_1608,N_1522,N_1527);
nor U1609 (N_1609,N_1548,N_1529);
and U1610 (N_1610,N_1544,N_1567);
or U1611 (N_1611,N_1511,N_1568);
or U1612 (N_1612,N_1520,N_1509);
nor U1613 (N_1613,N_1520,N_1561);
xnor U1614 (N_1614,N_1526,N_1507);
nand U1615 (N_1615,N_1508,N_1547);
and U1616 (N_1616,N_1502,N_1568);
nand U1617 (N_1617,N_1562,N_1545);
nor U1618 (N_1618,N_1527,N_1554);
or U1619 (N_1619,N_1507,N_1513);
nor U1620 (N_1620,N_1519,N_1565);
nor U1621 (N_1621,N_1517,N_1566);
or U1622 (N_1622,N_1536,N_1558);
or U1623 (N_1623,N_1517,N_1572);
nor U1624 (N_1624,N_1540,N_1552);
and U1625 (N_1625,N_1515,N_1522);
nor U1626 (N_1626,N_1544,N_1554);
nand U1627 (N_1627,N_1555,N_1519);
xnor U1628 (N_1628,N_1532,N_1536);
nand U1629 (N_1629,N_1567,N_1531);
or U1630 (N_1630,N_1572,N_1522);
nand U1631 (N_1631,N_1503,N_1543);
and U1632 (N_1632,N_1540,N_1514);
and U1633 (N_1633,N_1501,N_1504);
and U1634 (N_1634,N_1567,N_1570);
or U1635 (N_1635,N_1522,N_1521);
and U1636 (N_1636,N_1564,N_1548);
and U1637 (N_1637,N_1523,N_1524);
or U1638 (N_1638,N_1565,N_1569);
or U1639 (N_1639,N_1518,N_1570);
or U1640 (N_1640,N_1542,N_1515);
nand U1641 (N_1641,N_1533,N_1564);
and U1642 (N_1642,N_1523,N_1508);
nor U1643 (N_1643,N_1563,N_1559);
nor U1644 (N_1644,N_1542,N_1564);
nor U1645 (N_1645,N_1523,N_1536);
or U1646 (N_1646,N_1538,N_1526);
nand U1647 (N_1647,N_1548,N_1536);
nand U1648 (N_1648,N_1514,N_1556);
nor U1649 (N_1649,N_1520,N_1558);
and U1650 (N_1650,N_1639,N_1601);
or U1651 (N_1651,N_1597,N_1578);
and U1652 (N_1652,N_1622,N_1629);
and U1653 (N_1653,N_1640,N_1646);
nor U1654 (N_1654,N_1630,N_1645);
nor U1655 (N_1655,N_1592,N_1624);
nor U1656 (N_1656,N_1598,N_1605);
or U1657 (N_1657,N_1631,N_1596);
and U1658 (N_1658,N_1633,N_1583);
nor U1659 (N_1659,N_1620,N_1638);
or U1660 (N_1660,N_1619,N_1577);
nand U1661 (N_1661,N_1628,N_1627);
or U1662 (N_1662,N_1641,N_1575);
nand U1663 (N_1663,N_1582,N_1586);
nand U1664 (N_1664,N_1635,N_1637);
nor U1665 (N_1665,N_1616,N_1587);
and U1666 (N_1666,N_1595,N_1590);
xnor U1667 (N_1667,N_1623,N_1618);
or U1668 (N_1668,N_1621,N_1584);
nand U1669 (N_1669,N_1581,N_1602);
nand U1670 (N_1670,N_1606,N_1612);
nand U1671 (N_1671,N_1588,N_1649);
and U1672 (N_1672,N_1610,N_1647);
and U1673 (N_1673,N_1604,N_1603);
or U1674 (N_1674,N_1591,N_1615);
and U1675 (N_1675,N_1599,N_1585);
nand U1676 (N_1676,N_1611,N_1625);
or U1677 (N_1677,N_1644,N_1608);
and U1678 (N_1678,N_1614,N_1643);
and U1679 (N_1679,N_1607,N_1579);
nand U1680 (N_1680,N_1648,N_1589);
nand U1681 (N_1681,N_1609,N_1594);
nand U1682 (N_1682,N_1626,N_1576);
or U1683 (N_1683,N_1634,N_1593);
or U1684 (N_1684,N_1580,N_1642);
nor U1685 (N_1685,N_1613,N_1632);
nor U1686 (N_1686,N_1636,N_1600);
or U1687 (N_1687,N_1617,N_1639);
and U1688 (N_1688,N_1605,N_1631);
and U1689 (N_1689,N_1633,N_1646);
or U1690 (N_1690,N_1607,N_1637);
nor U1691 (N_1691,N_1616,N_1589);
and U1692 (N_1692,N_1607,N_1636);
and U1693 (N_1693,N_1575,N_1601);
nand U1694 (N_1694,N_1643,N_1618);
nor U1695 (N_1695,N_1602,N_1637);
nor U1696 (N_1696,N_1635,N_1585);
xnor U1697 (N_1697,N_1614,N_1584);
and U1698 (N_1698,N_1625,N_1639);
nor U1699 (N_1699,N_1593,N_1625);
and U1700 (N_1700,N_1642,N_1595);
nand U1701 (N_1701,N_1620,N_1621);
nor U1702 (N_1702,N_1630,N_1576);
nor U1703 (N_1703,N_1619,N_1646);
and U1704 (N_1704,N_1605,N_1638);
or U1705 (N_1705,N_1593,N_1595);
and U1706 (N_1706,N_1634,N_1601);
and U1707 (N_1707,N_1626,N_1648);
nor U1708 (N_1708,N_1645,N_1589);
nand U1709 (N_1709,N_1599,N_1649);
and U1710 (N_1710,N_1589,N_1634);
or U1711 (N_1711,N_1632,N_1631);
and U1712 (N_1712,N_1615,N_1605);
nand U1713 (N_1713,N_1633,N_1629);
nor U1714 (N_1714,N_1636,N_1619);
xnor U1715 (N_1715,N_1633,N_1619);
nor U1716 (N_1716,N_1632,N_1603);
or U1717 (N_1717,N_1633,N_1593);
and U1718 (N_1718,N_1599,N_1648);
and U1719 (N_1719,N_1613,N_1584);
and U1720 (N_1720,N_1642,N_1636);
and U1721 (N_1721,N_1614,N_1617);
and U1722 (N_1722,N_1578,N_1613);
and U1723 (N_1723,N_1632,N_1602);
nand U1724 (N_1724,N_1632,N_1583);
nor U1725 (N_1725,N_1670,N_1718);
or U1726 (N_1726,N_1689,N_1708);
or U1727 (N_1727,N_1676,N_1691);
nand U1728 (N_1728,N_1700,N_1664);
nor U1729 (N_1729,N_1680,N_1688);
nand U1730 (N_1730,N_1720,N_1724);
and U1731 (N_1731,N_1692,N_1697);
and U1732 (N_1732,N_1661,N_1681);
xnor U1733 (N_1733,N_1683,N_1712);
and U1734 (N_1734,N_1709,N_1687);
nor U1735 (N_1735,N_1650,N_1694);
and U1736 (N_1736,N_1722,N_1677);
nand U1737 (N_1737,N_1721,N_1665);
nand U1738 (N_1738,N_1707,N_1673);
nor U1739 (N_1739,N_1686,N_1705);
nor U1740 (N_1740,N_1653,N_1666);
nand U1741 (N_1741,N_1685,N_1668);
or U1742 (N_1742,N_1716,N_1696);
or U1743 (N_1743,N_1671,N_1657);
xnor U1744 (N_1744,N_1672,N_1706);
nor U1745 (N_1745,N_1723,N_1698);
nor U1746 (N_1746,N_1651,N_1662);
nand U1747 (N_1747,N_1659,N_1703);
nor U1748 (N_1748,N_1717,N_1656);
nor U1749 (N_1749,N_1711,N_1715);
and U1750 (N_1750,N_1679,N_1682);
nand U1751 (N_1751,N_1684,N_1675);
or U1752 (N_1752,N_1710,N_1667);
nand U1753 (N_1753,N_1704,N_1719);
and U1754 (N_1754,N_1652,N_1663);
nand U1755 (N_1755,N_1695,N_1654);
or U1756 (N_1756,N_1714,N_1701);
nor U1757 (N_1757,N_1669,N_1702);
or U1758 (N_1758,N_1678,N_1693);
nor U1759 (N_1759,N_1690,N_1655);
nand U1760 (N_1760,N_1674,N_1660);
nand U1761 (N_1761,N_1713,N_1658);
nand U1762 (N_1762,N_1699,N_1658);
nor U1763 (N_1763,N_1687,N_1710);
nor U1764 (N_1764,N_1658,N_1687);
nand U1765 (N_1765,N_1711,N_1671);
and U1766 (N_1766,N_1710,N_1689);
nor U1767 (N_1767,N_1699,N_1676);
or U1768 (N_1768,N_1665,N_1661);
nand U1769 (N_1769,N_1714,N_1724);
or U1770 (N_1770,N_1704,N_1652);
or U1771 (N_1771,N_1690,N_1686);
or U1772 (N_1772,N_1693,N_1690);
or U1773 (N_1773,N_1685,N_1699);
or U1774 (N_1774,N_1659,N_1713);
or U1775 (N_1775,N_1701,N_1702);
and U1776 (N_1776,N_1713,N_1685);
nand U1777 (N_1777,N_1698,N_1661);
nor U1778 (N_1778,N_1678,N_1694);
nor U1779 (N_1779,N_1713,N_1721);
or U1780 (N_1780,N_1665,N_1680);
or U1781 (N_1781,N_1713,N_1723);
nand U1782 (N_1782,N_1706,N_1687);
and U1783 (N_1783,N_1714,N_1662);
nor U1784 (N_1784,N_1656,N_1716);
nor U1785 (N_1785,N_1653,N_1665);
nor U1786 (N_1786,N_1684,N_1718);
or U1787 (N_1787,N_1705,N_1671);
nand U1788 (N_1788,N_1717,N_1660);
nor U1789 (N_1789,N_1689,N_1704);
or U1790 (N_1790,N_1663,N_1702);
and U1791 (N_1791,N_1663,N_1669);
or U1792 (N_1792,N_1660,N_1715);
and U1793 (N_1793,N_1722,N_1697);
nor U1794 (N_1794,N_1711,N_1713);
nor U1795 (N_1795,N_1685,N_1653);
nand U1796 (N_1796,N_1710,N_1704);
and U1797 (N_1797,N_1684,N_1693);
or U1798 (N_1798,N_1666,N_1665);
nand U1799 (N_1799,N_1667,N_1664);
nand U1800 (N_1800,N_1744,N_1746);
or U1801 (N_1801,N_1736,N_1741);
or U1802 (N_1802,N_1737,N_1764);
or U1803 (N_1803,N_1785,N_1748);
nand U1804 (N_1804,N_1765,N_1732);
and U1805 (N_1805,N_1799,N_1756);
and U1806 (N_1806,N_1782,N_1772);
or U1807 (N_1807,N_1747,N_1754);
and U1808 (N_1808,N_1725,N_1729);
or U1809 (N_1809,N_1774,N_1770);
or U1810 (N_1810,N_1792,N_1735);
nand U1811 (N_1811,N_1797,N_1791);
or U1812 (N_1812,N_1787,N_1749);
or U1813 (N_1813,N_1763,N_1734);
or U1814 (N_1814,N_1780,N_1727);
or U1815 (N_1815,N_1739,N_1793);
and U1816 (N_1816,N_1776,N_1728);
and U1817 (N_1817,N_1771,N_1726);
nand U1818 (N_1818,N_1745,N_1798);
nand U1819 (N_1819,N_1794,N_1761);
nand U1820 (N_1820,N_1759,N_1796);
nand U1821 (N_1821,N_1740,N_1773);
nor U1822 (N_1822,N_1767,N_1742);
nor U1823 (N_1823,N_1777,N_1784);
and U1824 (N_1824,N_1790,N_1786);
nand U1825 (N_1825,N_1755,N_1731);
nand U1826 (N_1826,N_1769,N_1750);
nand U1827 (N_1827,N_1779,N_1752);
and U1828 (N_1828,N_1775,N_1753);
and U1829 (N_1829,N_1743,N_1788);
and U1830 (N_1830,N_1758,N_1760);
and U1831 (N_1831,N_1789,N_1751);
nand U1832 (N_1832,N_1795,N_1778);
nand U1833 (N_1833,N_1768,N_1781);
or U1834 (N_1834,N_1766,N_1738);
nor U1835 (N_1835,N_1733,N_1783);
and U1836 (N_1836,N_1762,N_1757);
and U1837 (N_1837,N_1730,N_1752);
and U1838 (N_1838,N_1777,N_1767);
nor U1839 (N_1839,N_1745,N_1776);
or U1840 (N_1840,N_1794,N_1796);
and U1841 (N_1841,N_1764,N_1766);
and U1842 (N_1842,N_1738,N_1765);
nand U1843 (N_1843,N_1792,N_1783);
and U1844 (N_1844,N_1752,N_1784);
nand U1845 (N_1845,N_1786,N_1738);
or U1846 (N_1846,N_1749,N_1795);
or U1847 (N_1847,N_1725,N_1766);
and U1848 (N_1848,N_1786,N_1736);
or U1849 (N_1849,N_1759,N_1756);
and U1850 (N_1850,N_1774,N_1740);
and U1851 (N_1851,N_1758,N_1749);
or U1852 (N_1852,N_1775,N_1764);
or U1853 (N_1853,N_1793,N_1785);
and U1854 (N_1854,N_1745,N_1746);
xor U1855 (N_1855,N_1794,N_1769);
nor U1856 (N_1856,N_1763,N_1796);
nand U1857 (N_1857,N_1771,N_1780);
or U1858 (N_1858,N_1753,N_1782);
nor U1859 (N_1859,N_1786,N_1789);
xor U1860 (N_1860,N_1797,N_1762);
nand U1861 (N_1861,N_1730,N_1737);
nand U1862 (N_1862,N_1794,N_1741);
or U1863 (N_1863,N_1787,N_1778);
and U1864 (N_1864,N_1741,N_1761);
nand U1865 (N_1865,N_1737,N_1776);
nor U1866 (N_1866,N_1730,N_1770);
or U1867 (N_1867,N_1750,N_1782);
nor U1868 (N_1868,N_1787,N_1774);
or U1869 (N_1869,N_1740,N_1795);
or U1870 (N_1870,N_1737,N_1735);
and U1871 (N_1871,N_1735,N_1746);
nand U1872 (N_1872,N_1740,N_1768);
nor U1873 (N_1873,N_1793,N_1736);
and U1874 (N_1874,N_1759,N_1781);
xnor U1875 (N_1875,N_1874,N_1842);
nand U1876 (N_1876,N_1828,N_1854);
and U1877 (N_1877,N_1840,N_1860);
nor U1878 (N_1878,N_1831,N_1872);
and U1879 (N_1879,N_1849,N_1853);
nand U1880 (N_1880,N_1843,N_1812);
nand U1881 (N_1881,N_1858,N_1855);
and U1882 (N_1882,N_1862,N_1807);
or U1883 (N_1883,N_1845,N_1869);
and U1884 (N_1884,N_1815,N_1844);
and U1885 (N_1885,N_1867,N_1816);
or U1886 (N_1886,N_1825,N_1804);
or U1887 (N_1887,N_1859,N_1838);
or U1888 (N_1888,N_1852,N_1801);
nand U1889 (N_1889,N_1835,N_1822);
or U1890 (N_1890,N_1805,N_1871);
or U1891 (N_1891,N_1810,N_1802);
nor U1892 (N_1892,N_1847,N_1836);
and U1893 (N_1893,N_1865,N_1813);
nand U1894 (N_1894,N_1806,N_1823);
nand U1895 (N_1895,N_1864,N_1821);
or U1896 (N_1896,N_1826,N_1870);
nand U1897 (N_1897,N_1841,N_1808);
nand U1898 (N_1898,N_1833,N_1827);
nand U1899 (N_1899,N_1819,N_1866);
or U1900 (N_1900,N_1814,N_1848);
or U1901 (N_1901,N_1857,N_1818);
or U1902 (N_1902,N_1803,N_1834);
or U1903 (N_1903,N_1817,N_1824);
nand U1904 (N_1904,N_1832,N_1830);
nor U1905 (N_1905,N_1800,N_1868);
nand U1906 (N_1906,N_1873,N_1846);
nor U1907 (N_1907,N_1839,N_1861);
and U1908 (N_1908,N_1837,N_1850);
and U1909 (N_1909,N_1820,N_1856);
nor U1910 (N_1910,N_1809,N_1851);
or U1911 (N_1911,N_1829,N_1863);
or U1912 (N_1912,N_1811,N_1803);
nor U1913 (N_1913,N_1864,N_1812);
and U1914 (N_1914,N_1819,N_1856);
nand U1915 (N_1915,N_1845,N_1870);
and U1916 (N_1916,N_1831,N_1855);
or U1917 (N_1917,N_1848,N_1866);
nor U1918 (N_1918,N_1847,N_1857);
or U1919 (N_1919,N_1845,N_1854);
and U1920 (N_1920,N_1867,N_1870);
nand U1921 (N_1921,N_1841,N_1827);
nor U1922 (N_1922,N_1824,N_1861);
and U1923 (N_1923,N_1836,N_1869);
nor U1924 (N_1924,N_1818,N_1865);
or U1925 (N_1925,N_1874,N_1862);
nor U1926 (N_1926,N_1815,N_1813);
nor U1927 (N_1927,N_1865,N_1812);
nand U1928 (N_1928,N_1843,N_1811);
or U1929 (N_1929,N_1836,N_1800);
or U1930 (N_1930,N_1800,N_1860);
or U1931 (N_1931,N_1852,N_1825);
or U1932 (N_1932,N_1848,N_1811);
nand U1933 (N_1933,N_1840,N_1865);
nor U1934 (N_1934,N_1821,N_1812);
nor U1935 (N_1935,N_1849,N_1803);
nor U1936 (N_1936,N_1833,N_1865);
nor U1937 (N_1937,N_1804,N_1855);
nor U1938 (N_1938,N_1857,N_1853);
or U1939 (N_1939,N_1832,N_1842);
xnor U1940 (N_1940,N_1819,N_1862);
and U1941 (N_1941,N_1829,N_1813);
or U1942 (N_1942,N_1842,N_1840);
and U1943 (N_1943,N_1809,N_1835);
nor U1944 (N_1944,N_1849,N_1839);
nand U1945 (N_1945,N_1810,N_1823);
or U1946 (N_1946,N_1817,N_1838);
nand U1947 (N_1947,N_1868,N_1858);
nand U1948 (N_1948,N_1809,N_1832);
or U1949 (N_1949,N_1863,N_1836);
nand U1950 (N_1950,N_1912,N_1900);
and U1951 (N_1951,N_1884,N_1937);
or U1952 (N_1952,N_1939,N_1885);
nor U1953 (N_1953,N_1922,N_1936);
and U1954 (N_1954,N_1904,N_1919);
or U1955 (N_1955,N_1903,N_1901);
nand U1956 (N_1956,N_1926,N_1932);
or U1957 (N_1957,N_1890,N_1945);
nand U1958 (N_1958,N_1879,N_1946);
nor U1959 (N_1959,N_1940,N_1877);
or U1960 (N_1960,N_1938,N_1893);
and U1961 (N_1961,N_1910,N_1899);
or U1962 (N_1962,N_1941,N_1875);
and U1963 (N_1963,N_1949,N_1913);
nor U1964 (N_1964,N_1933,N_1942);
nor U1965 (N_1965,N_1886,N_1924);
nor U1966 (N_1966,N_1916,N_1881);
or U1967 (N_1967,N_1928,N_1898);
nand U1968 (N_1968,N_1920,N_1947);
nand U1969 (N_1969,N_1915,N_1891);
nor U1970 (N_1970,N_1896,N_1902);
nor U1971 (N_1971,N_1908,N_1880);
and U1972 (N_1972,N_1907,N_1925);
nand U1973 (N_1973,N_1929,N_1930);
or U1974 (N_1974,N_1897,N_1921);
nand U1975 (N_1975,N_1917,N_1894);
and U1976 (N_1976,N_1889,N_1895);
and U1977 (N_1977,N_1887,N_1892);
and U1978 (N_1978,N_1935,N_1905);
nand U1979 (N_1979,N_1934,N_1948);
nand U1980 (N_1980,N_1914,N_1927);
or U1981 (N_1981,N_1883,N_1882);
or U1982 (N_1982,N_1906,N_1931);
nand U1983 (N_1983,N_1911,N_1918);
or U1984 (N_1984,N_1878,N_1944);
or U1985 (N_1985,N_1923,N_1876);
and U1986 (N_1986,N_1888,N_1943);
or U1987 (N_1987,N_1909,N_1907);
and U1988 (N_1988,N_1906,N_1908);
or U1989 (N_1989,N_1932,N_1916);
or U1990 (N_1990,N_1923,N_1930);
and U1991 (N_1991,N_1911,N_1907);
and U1992 (N_1992,N_1949,N_1925);
or U1993 (N_1993,N_1890,N_1946);
nand U1994 (N_1994,N_1937,N_1897);
and U1995 (N_1995,N_1885,N_1889);
or U1996 (N_1996,N_1913,N_1882);
and U1997 (N_1997,N_1901,N_1937);
nand U1998 (N_1998,N_1937,N_1912);
nor U1999 (N_1999,N_1883,N_1910);
nand U2000 (N_2000,N_1904,N_1883);
or U2001 (N_2001,N_1887,N_1942);
nor U2002 (N_2002,N_1901,N_1949);
nor U2003 (N_2003,N_1895,N_1891);
or U2004 (N_2004,N_1919,N_1911);
nor U2005 (N_2005,N_1936,N_1885);
and U2006 (N_2006,N_1882,N_1910);
nand U2007 (N_2007,N_1905,N_1918);
nor U2008 (N_2008,N_1927,N_1885);
nor U2009 (N_2009,N_1936,N_1929);
nand U2010 (N_2010,N_1942,N_1897);
and U2011 (N_2011,N_1908,N_1942);
nor U2012 (N_2012,N_1883,N_1945);
or U2013 (N_2013,N_1943,N_1909);
nor U2014 (N_2014,N_1885,N_1921);
nand U2015 (N_2015,N_1919,N_1898);
or U2016 (N_2016,N_1899,N_1942);
xnor U2017 (N_2017,N_1944,N_1889);
or U2018 (N_2018,N_1888,N_1881);
nor U2019 (N_2019,N_1921,N_1884);
and U2020 (N_2020,N_1924,N_1942);
and U2021 (N_2021,N_1887,N_1896);
and U2022 (N_2022,N_1917,N_1933);
nor U2023 (N_2023,N_1894,N_1876);
and U2024 (N_2024,N_1888,N_1949);
nor U2025 (N_2025,N_1980,N_1971);
and U2026 (N_2026,N_1951,N_2010);
nand U2027 (N_2027,N_1956,N_1970);
and U2028 (N_2028,N_1992,N_2012);
nand U2029 (N_2029,N_1967,N_2023);
or U2030 (N_2030,N_1972,N_1952);
and U2031 (N_2031,N_1983,N_1994);
nor U2032 (N_2032,N_1965,N_1950);
nand U2033 (N_2033,N_1966,N_1988);
and U2034 (N_2034,N_2018,N_1999);
xnor U2035 (N_2035,N_1973,N_1987);
nor U2036 (N_2036,N_2011,N_1993);
or U2037 (N_2037,N_2001,N_1996);
nand U2038 (N_2038,N_1986,N_2003);
or U2039 (N_2039,N_1954,N_1997);
nand U2040 (N_2040,N_2006,N_1998);
nor U2041 (N_2041,N_1982,N_2007);
nand U2042 (N_2042,N_2004,N_1974);
nand U2043 (N_2043,N_1963,N_1958);
nor U2044 (N_2044,N_1959,N_1969);
nand U2045 (N_2045,N_2005,N_1962);
or U2046 (N_2046,N_2000,N_1985);
or U2047 (N_2047,N_1976,N_2009);
and U2048 (N_2048,N_1991,N_2016);
nand U2049 (N_2049,N_2021,N_1995);
nand U2050 (N_2050,N_2015,N_1968);
nor U2051 (N_2051,N_2020,N_2014);
nor U2052 (N_2052,N_1989,N_1990);
xnor U2053 (N_2053,N_1960,N_2024);
and U2054 (N_2054,N_1981,N_2002);
or U2055 (N_2055,N_2008,N_1984);
or U2056 (N_2056,N_2017,N_1977);
or U2057 (N_2057,N_1955,N_2022);
or U2058 (N_2058,N_1957,N_1975);
or U2059 (N_2059,N_2013,N_1964);
and U2060 (N_2060,N_1953,N_1978);
and U2061 (N_2061,N_1979,N_2019);
nor U2062 (N_2062,N_1961,N_2014);
and U2063 (N_2063,N_2007,N_2005);
xor U2064 (N_2064,N_2005,N_2001);
nand U2065 (N_2065,N_1965,N_2014);
nand U2066 (N_2066,N_1971,N_1986);
nand U2067 (N_2067,N_1976,N_2004);
nor U2068 (N_2068,N_2018,N_1952);
nor U2069 (N_2069,N_1980,N_1979);
or U2070 (N_2070,N_1959,N_1979);
nand U2071 (N_2071,N_2006,N_1997);
and U2072 (N_2072,N_2006,N_1952);
and U2073 (N_2073,N_1952,N_1974);
and U2074 (N_2074,N_1950,N_2006);
or U2075 (N_2075,N_1989,N_1959);
nor U2076 (N_2076,N_1954,N_2007);
and U2077 (N_2077,N_1952,N_1987);
nor U2078 (N_2078,N_1950,N_2005);
nand U2079 (N_2079,N_1974,N_1950);
and U2080 (N_2080,N_1975,N_2023);
nand U2081 (N_2081,N_1967,N_1981);
nand U2082 (N_2082,N_1964,N_2001);
or U2083 (N_2083,N_1972,N_1957);
nand U2084 (N_2084,N_1974,N_1977);
nand U2085 (N_2085,N_1954,N_1989);
nand U2086 (N_2086,N_1965,N_1953);
nor U2087 (N_2087,N_1964,N_1960);
and U2088 (N_2088,N_1984,N_1982);
and U2089 (N_2089,N_1983,N_1991);
nor U2090 (N_2090,N_1997,N_2018);
or U2091 (N_2091,N_1973,N_2022);
nor U2092 (N_2092,N_1950,N_2017);
or U2093 (N_2093,N_2018,N_2023);
nor U2094 (N_2094,N_1990,N_1988);
or U2095 (N_2095,N_1997,N_1992);
or U2096 (N_2096,N_1979,N_1995);
nor U2097 (N_2097,N_2010,N_1969);
nand U2098 (N_2098,N_1985,N_1991);
nand U2099 (N_2099,N_2023,N_2003);
nand U2100 (N_2100,N_2064,N_2098);
nor U2101 (N_2101,N_2031,N_2045);
or U2102 (N_2102,N_2062,N_2082);
xnor U2103 (N_2103,N_2095,N_2077);
or U2104 (N_2104,N_2089,N_2058);
or U2105 (N_2105,N_2041,N_2099);
or U2106 (N_2106,N_2043,N_2063);
and U2107 (N_2107,N_2050,N_2026);
nor U2108 (N_2108,N_2085,N_2061);
or U2109 (N_2109,N_2066,N_2097);
or U2110 (N_2110,N_2025,N_2088);
and U2111 (N_2111,N_2084,N_2081);
nor U2112 (N_2112,N_2076,N_2091);
and U2113 (N_2113,N_2078,N_2072);
nor U2114 (N_2114,N_2055,N_2047);
nor U2115 (N_2115,N_2034,N_2054);
xor U2116 (N_2116,N_2068,N_2059);
or U2117 (N_2117,N_2074,N_2090);
and U2118 (N_2118,N_2037,N_2093);
or U2119 (N_2119,N_2060,N_2042);
nor U2120 (N_2120,N_2071,N_2065);
or U2121 (N_2121,N_2028,N_2044);
nor U2122 (N_2122,N_2067,N_2094);
nor U2123 (N_2123,N_2052,N_2030);
nand U2124 (N_2124,N_2073,N_2036);
nor U2125 (N_2125,N_2038,N_2080);
and U2126 (N_2126,N_2053,N_2039);
nand U2127 (N_2127,N_2032,N_2069);
nor U2128 (N_2128,N_2033,N_2048);
and U2129 (N_2129,N_2086,N_2040);
nand U2130 (N_2130,N_2035,N_2096);
nand U2131 (N_2131,N_2092,N_2049);
and U2132 (N_2132,N_2046,N_2079);
and U2133 (N_2133,N_2057,N_2056);
nor U2134 (N_2134,N_2070,N_2075);
and U2135 (N_2135,N_2029,N_2027);
and U2136 (N_2136,N_2083,N_2051);
and U2137 (N_2137,N_2087,N_2039);
or U2138 (N_2138,N_2093,N_2044);
nor U2139 (N_2139,N_2095,N_2035);
nand U2140 (N_2140,N_2025,N_2085);
nand U2141 (N_2141,N_2028,N_2070);
nor U2142 (N_2142,N_2051,N_2028);
nor U2143 (N_2143,N_2030,N_2082);
xnor U2144 (N_2144,N_2087,N_2042);
or U2145 (N_2145,N_2081,N_2037);
and U2146 (N_2146,N_2039,N_2078);
and U2147 (N_2147,N_2065,N_2067);
nand U2148 (N_2148,N_2057,N_2031);
nand U2149 (N_2149,N_2036,N_2046);
and U2150 (N_2150,N_2089,N_2035);
or U2151 (N_2151,N_2063,N_2083);
and U2152 (N_2152,N_2041,N_2080);
nor U2153 (N_2153,N_2045,N_2033);
nor U2154 (N_2154,N_2045,N_2037);
and U2155 (N_2155,N_2084,N_2039);
nor U2156 (N_2156,N_2032,N_2067);
and U2157 (N_2157,N_2059,N_2043);
and U2158 (N_2158,N_2066,N_2077);
or U2159 (N_2159,N_2027,N_2076);
nor U2160 (N_2160,N_2030,N_2034);
nor U2161 (N_2161,N_2029,N_2065);
and U2162 (N_2162,N_2092,N_2029);
and U2163 (N_2163,N_2029,N_2082);
or U2164 (N_2164,N_2089,N_2049);
nand U2165 (N_2165,N_2066,N_2095);
nor U2166 (N_2166,N_2041,N_2088);
or U2167 (N_2167,N_2049,N_2035);
or U2168 (N_2168,N_2076,N_2070);
nand U2169 (N_2169,N_2031,N_2073);
nor U2170 (N_2170,N_2096,N_2085);
nor U2171 (N_2171,N_2079,N_2078);
nor U2172 (N_2172,N_2036,N_2082);
nand U2173 (N_2173,N_2065,N_2082);
or U2174 (N_2174,N_2034,N_2048);
nor U2175 (N_2175,N_2106,N_2151);
or U2176 (N_2176,N_2162,N_2110);
or U2177 (N_2177,N_2131,N_2174);
and U2178 (N_2178,N_2113,N_2173);
and U2179 (N_2179,N_2140,N_2124);
nand U2180 (N_2180,N_2115,N_2130);
and U2181 (N_2181,N_2147,N_2121);
or U2182 (N_2182,N_2132,N_2150);
nor U2183 (N_2183,N_2123,N_2139);
nand U2184 (N_2184,N_2102,N_2105);
and U2185 (N_2185,N_2136,N_2142);
nand U2186 (N_2186,N_2170,N_2167);
or U2187 (N_2187,N_2122,N_2117);
and U2188 (N_2188,N_2171,N_2146);
or U2189 (N_2189,N_2137,N_2125);
or U2190 (N_2190,N_2127,N_2152);
nor U2191 (N_2191,N_2120,N_2119);
nor U2192 (N_2192,N_2163,N_2135);
nor U2193 (N_2193,N_2168,N_2145);
nor U2194 (N_2194,N_2118,N_2101);
nor U2195 (N_2195,N_2169,N_2148);
nand U2196 (N_2196,N_2109,N_2141);
and U2197 (N_2197,N_2157,N_2112);
nor U2198 (N_2198,N_2108,N_2160);
nor U2199 (N_2199,N_2166,N_2153);
and U2200 (N_2200,N_2159,N_2172);
nand U2201 (N_2201,N_2155,N_2158);
nand U2202 (N_2202,N_2134,N_2100);
nor U2203 (N_2203,N_2111,N_2126);
nand U2204 (N_2204,N_2116,N_2103);
nor U2205 (N_2205,N_2161,N_2128);
nor U2206 (N_2206,N_2107,N_2133);
nor U2207 (N_2207,N_2114,N_2165);
or U2208 (N_2208,N_2138,N_2164);
and U2209 (N_2209,N_2129,N_2104);
and U2210 (N_2210,N_2149,N_2143);
nand U2211 (N_2211,N_2156,N_2144);
and U2212 (N_2212,N_2154,N_2169);
or U2213 (N_2213,N_2174,N_2162);
or U2214 (N_2214,N_2105,N_2132);
nand U2215 (N_2215,N_2148,N_2158);
nand U2216 (N_2216,N_2106,N_2161);
nand U2217 (N_2217,N_2163,N_2166);
nor U2218 (N_2218,N_2119,N_2155);
xnor U2219 (N_2219,N_2103,N_2125);
nor U2220 (N_2220,N_2172,N_2135);
or U2221 (N_2221,N_2114,N_2148);
nor U2222 (N_2222,N_2168,N_2106);
and U2223 (N_2223,N_2124,N_2160);
or U2224 (N_2224,N_2173,N_2174);
and U2225 (N_2225,N_2119,N_2102);
or U2226 (N_2226,N_2135,N_2141);
nor U2227 (N_2227,N_2158,N_2125);
or U2228 (N_2228,N_2133,N_2116);
nand U2229 (N_2229,N_2157,N_2129);
xnor U2230 (N_2230,N_2122,N_2173);
nand U2231 (N_2231,N_2111,N_2165);
and U2232 (N_2232,N_2169,N_2104);
and U2233 (N_2233,N_2169,N_2170);
nor U2234 (N_2234,N_2149,N_2133);
nand U2235 (N_2235,N_2127,N_2171);
nand U2236 (N_2236,N_2124,N_2114);
or U2237 (N_2237,N_2153,N_2160);
or U2238 (N_2238,N_2101,N_2151);
nand U2239 (N_2239,N_2172,N_2104);
and U2240 (N_2240,N_2145,N_2159);
nor U2241 (N_2241,N_2172,N_2164);
nand U2242 (N_2242,N_2108,N_2149);
nor U2243 (N_2243,N_2137,N_2114);
nor U2244 (N_2244,N_2129,N_2127);
or U2245 (N_2245,N_2172,N_2124);
xnor U2246 (N_2246,N_2153,N_2130);
or U2247 (N_2247,N_2151,N_2129);
nand U2248 (N_2248,N_2139,N_2143);
or U2249 (N_2249,N_2117,N_2152);
and U2250 (N_2250,N_2227,N_2196);
and U2251 (N_2251,N_2236,N_2183);
or U2252 (N_2252,N_2179,N_2238);
nand U2253 (N_2253,N_2243,N_2247);
xnor U2254 (N_2254,N_2189,N_2195);
or U2255 (N_2255,N_2233,N_2180);
or U2256 (N_2256,N_2178,N_2232);
nor U2257 (N_2257,N_2200,N_2210);
and U2258 (N_2258,N_2234,N_2192);
and U2259 (N_2259,N_2220,N_2224);
or U2260 (N_2260,N_2175,N_2201);
nand U2261 (N_2261,N_2219,N_2222);
and U2262 (N_2262,N_2241,N_2181);
nand U2263 (N_2263,N_2223,N_2240);
nand U2264 (N_2264,N_2217,N_2177);
nor U2265 (N_2265,N_2245,N_2215);
or U2266 (N_2266,N_2199,N_2186);
nor U2267 (N_2267,N_2185,N_2229);
nand U2268 (N_2268,N_2194,N_2197);
nor U2269 (N_2269,N_2190,N_2225);
or U2270 (N_2270,N_2202,N_2198);
or U2271 (N_2271,N_2184,N_2212);
or U2272 (N_2272,N_2203,N_2221);
and U2273 (N_2273,N_2208,N_2218);
xor U2274 (N_2274,N_2214,N_2204);
nand U2275 (N_2275,N_2188,N_2244);
nand U2276 (N_2276,N_2235,N_2211);
nand U2277 (N_2277,N_2246,N_2193);
nor U2278 (N_2278,N_2205,N_2176);
nor U2279 (N_2279,N_2231,N_2207);
nor U2280 (N_2280,N_2216,N_2239);
or U2281 (N_2281,N_2228,N_2209);
and U2282 (N_2282,N_2248,N_2213);
and U2283 (N_2283,N_2182,N_2226);
nor U2284 (N_2284,N_2237,N_2249);
nand U2285 (N_2285,N_2187,N_2206);
or U2286 (N_2286,N_2191,N_2230);
nor U2287 (N_2287,N_2242,N_2240);
nand U2288 (N_2288,N_2206,N_2241);
nand U2289 (N_2289,N_2210,N_2233);
nor U2290 (N_2290,N_2192,N_2194);
nand U2291 (N_2291,N_2179,N_2222);
nand U2292 (N_2292,N_2222,N_2194);
nor U2293 (N_2293,N_2206,N_2244);
or U2294 (N_2294,N_2179,N_2233);
nand U2295 (N_2295,N_2184,N_2244);
xor U2296 (N_2296,N_2234,N_2187);
or U2297 (N_2297,N_2188,N_2246);
nor U2298 (N_2298,N_2180,N_2177);
nor U2299 (N_2299,N_2244,N_2243);
nand U2300 (N_2300,N_2206,N_2208);
and U2301 (N_2301,N_2207,N_2182);
nand U2302 (N_2302,N_2198,N_2175);
and U2303 (N_2303,N_2217,N_2224);
or U2304 (N_2304,N_2193,N_2191);
nor U2305 (N_2305,N_2196,N_2245);
nor U2306 (N_2306,N_2188,N_2219);
nand U2307 (N_2307,N_2176,N_2220);
nor U2308 (N_2308,N_2178,N_2231);
and U2309 (N_2309,N_2224,N_2229);
or U2310 (N_2310,N_2211,N_2183);
nor U2311 (N_2311,N_2237,N_2198);
and U2312 (N_2312,N_2196,N_2238);
nand U2313 (N_2313,N_2244,N_2215);
and U2314 (N_2314,N_2186,N_2218);
nor U2315 (N_2315,N_2182,N_2249);
or U2316 (N_2316,N_2248,N_2247);
and U2317 (N_2317,N_2209,N_2183);
nand U2318 (N_2318,N_2193,N_2215);
or U2319 (N_2319,N_2219,N_2225);
and U2320 (N_2320,N_2207,N_2192);
nor U2321 (N_2321,N_2201,N_2237);
nand U2322 (N_2322,N_2186,N_2225);
or U2323 (N_2323,N_2175,N_2235);
nor U2324 (N_2324,N_2219,N_2235);
or U2325 (N_2325,N_2311,N_2270);
nand U2326 (N_2326,N_2284,N_2285);
or U2327 (N_2327,N_2263,N_2282);
or U2328 (N_2328,N_2324,N_2286);
nor U2329 (N_2329,N_2250,N_2255);
nor U2330 (N_2330,N_2264,N_2271);
and U2331 (N_2331,N_2275,N_2261);
xnor U2332 (N_2332,N_2302,N_2276);
nor U2333 (N_2333,N_2309,N_2296);
nor U2334 (N_2334,N_2319,N_2259);
and U2335 (N_2335,N_2318,N_2283);
nor U2336 (N_2336,N_2252,N_2322);
nand U2337 (N_2337,N_2274,N_2305);
nand U2338 (N_2338,N_2320,N_2306);
nand U2339 (N_2339,N_2269,N_2298);
nand U2340 (N_2340,N_2303,N_2289);
or U2341 (N_2341,N_2315,N_2257);
nand U2342 (N_2342,N_2297,N_2317);
nor U2343 (N_2343,N_2266,N_2278);
and U2344 (N_2344,N_2299,N_2251);
nand U2345 (N_2345,N_2288,N_2295);
or U2346 (N_2346,N_2300,N_2272);
or U2347 (N_2347,N_2304,N_2277);
nand U2348 (N_2348,N_2312,N_2253);
nand U2349 (N_2349,N_2291,N_2258);
and U2350 (N_2350,N_2265,N_2268);
nand U2351 (N_2351,N_2321,N_2308);
and U2352 (N_2352,N_2294,N_2310);
and U2353 (N_2353,N_2313,N_2287);
and U2354 (N_2354,N_2290,N_2256);
or U2355 (N_2355,N_2301,N_2307);
nand U2356 (N_2356,N_2292,N_2280);
nor U2357 (N_2357,N_2314,N_2262);
and U2358 (N_2358,N_2316,N_2260);
or U2359 (N_2359,N_2293,N_2254);
and U2360 (N_2360,N_2273,N_2323);
nor U2361 (N_2361,N_2279,N_2267);
nor U2362 (N_2362,N_2281,N_2261);
nor U2363 (N_2363,N_2313,N_2281);
nor U2364 (N_2364,N_2295,N_2283);
nand U2365 (N_2365,N_2261,N_2299);
nor U2366 (N_2366,N_2280,N_2324);
or U2367 (N_2367,N_2303,N_2267);
or U2368 (N_2368,N_2267,N_2315);
and U2369 (N_2369,N_2263,N_2320);
nand U2370 (N_2370,N_2296,N_2310);
and U2371 (N_2371,N_2289,N_2310);
nand U2372 (N_2372,N_2294,N_2323);
and U2373 (N_2373,N_2303,N_2257);
or U2374 (N_2374,N_2299,N_2279);
nand U2375 (N_2375,N_2305,N_2262);
or U2376 (N_2376,N_2293,N_2292);
nand U2377 (N_2377,N_2308,N_2302);
and U2378 (N_2378,N_2282,N_2277);
and U2379 (N_2379,N_2304,N_2284);
nor U2380 (N_2380,N_2291,N_2302);
or U2381 (N_2381,N_2280,N_2317);
nand U2382 (N_2382,N_2254,N_2316);
nor U2383 (N_2383,N_2292,N_2323);
and U2384 (N_2384,N_2291,N_2267);
or U2385 (N_2385,N_2288,N_2256);
nand U2386 (N_2386,N_2273,N_2251);
nand U2387 (N_2387,N_2318,N_2263);
or U2388 (N_2388,N_2276,N_2268);
nor U2389 (N_2389,N_2322,N_2289);
nand U2390 (N_2390,N_2302,N_2311);
or U2391 (N_2391,N_2290,N_2282);
nor U2392 (N_2392,N_2281,N_2272);
and U2393 (N_2393,N_2290,N_2280);
or U2394 (N_2394,N_2267,N_2270);
and U2395 (N_2395,N_2309,N_2257);
or U2396 (N_2396,N_2251,N_2269);
nand U2397 (N_2397,N_2298,N_2294);
nand U2398 (N_2398,N_2281,N_2296);
nand U2399 (N_2399,N_2302,N_2280);
nand U2400 (N_2400,N_2363,N_2362);
and U2401 (N_2401,N_2372,N_2374);
or U2402 (N_2402,N_2341,N_2384);
and U2403 (N_2403,N_2385,N_2387);
nor U2404 (N_2404,N_2397,N_2349);
nor U2405 (N_2405,N_2382,N_2381);
or U2406 (N_2406,N_2366,N_2361);
nand U2407 (N_2407,N_2336,N_2376);
and U2408 (N_2408,N_2367,N_2375);
and U2409 (N_2409,N_2391,N_2328);
and U2410 (N_2410,N_2357,N_2371);
nor U2411 (N_2411,N_2343,N_2398);
or U2412 (N_2412,N_2327,N_2390);
and U2413 (N_2413,N_2364,N_2331);
or U2414 (N_2414,N_2380,N_2353);
nor U2415 (N_2415,N_2338,N_2347);
or U2416 (N_2416,N_2365,N_2370);
nor U2417 (N_2417,N_2326,N_2339);
or U2418 (N_2418,N_2344,N_2356);
and U2419 (N_2419,N_2389,N_2392);
and U2420 (N_2420,N_2334,N_2393);
nand U2421 (N_2421,N_2379,N_2369);
and U2422 (N_2422,N_2340,N_2329);
or U2423 (N_2423,N_2333,N_2350);
and U2424 (N_2424,N_2394,N_2359);
nor U2425 (N_2425,N_2325,N_2396);
or U2426 (N_2426,N_2352,N_2335);
and U2427 (N_2427,N_2358,N_2342);
nor U2428 (N_2428,N_2386,N_2399);
or U2429 (N_2429,N_2377,N_2368);
nor U2430 (N_2430,N_2332,N_2346);
nand U2431 (N_2431,N_2383,N_2373);
nand U2432 (N_2432,N_2378,N_2351);
nor U2433 (N_2433,N_2345,N_2348);
and U2434 (N_2434,N_2330,N_2355);
or U2435 (N_2435,N_2388,N_2337);
nor U2436 (N_2436,N_2360,N_2395);
or U2437 (N_2437,N_2354,N_2395);
nor U2438 (N_2438,N_2392,N_2359);
nor U2439 (N_2439,N_2363,N_2345);
or U2440 (N_2440,N_2358,N_2339);
nor U2441 (N_2441,N_2368,N_2359);
or U2442 (N_2442,N_2328,N_2363);
nor U2443 (N_2443,N_2351,N_2388);
nand U2444 (N_2444,N_2342,N_2340);
xnor U2445 (N_2445,N_2344,N_2361);
or U2446 (N_2446,N_2397,N_2338);
and U2447 (N_2447,N_2380,N_2325);
or U2448 (N_2448,N_2387,N_2329);
or U2449 (N_2449,N_2332,N_2341);
nor U2450 (N_2450,N_2388,N_2371);
or U2451 (N_2451,N_2389,N_2382);
nand U2452 (N_2452,N_2380,N_2352);
or U2453 (N_2453,N_2373,N_2389);
nand U2454 (N_2454,N_2355,N_2386);
nor U2455 (N_2455,N_2356,N_2366);
nor U2456 (N_2456,N_2366,N_2386);
or U2457 (N_2457,N_2370,N_2327);
and U2458 (N_2458,N_2395,N_2332);
and U2459 (N_2459,N_2325,N_2365);
nor U2460 (N_2460,N_2363,N_2327);
or U2461 (N_2461,N_2389,N_2398);
nor U2462 (N_2462,N_2365,N_2333);
and U2463 (N_2463,N_2388,N_2355);
nor U2464 (N_2464,N_2367,N_2360);
or U2465 (N_2465,N_2380,N_2393);
and U2466 (N_2466,N_2347,N_2348);
and U2467 (N_2467,N_2378,N_2331);
nand U2468 (N_2468,N_2375,N_2357);
nand U2469 (N_2469,N_2347,N_2354);
or U2470 (N_2470,N_2343,N_2390);
nor U2471 (N_2471,N_2364,N_2379);
nand U2472 (N_2472,N_2345,N_2332);
xnor U2473 (N_2473,N_2397,N_2395);
nand U2474 (N_2474,N_2377,N_2394);
nand U2475 (N_2475,N_2447,N_2423);
nor U2476 (N_2476,N_2430,N_2422);
nor U2477 (N_2477,N_2411,N_2457);
nand U2478 (N_2478,N_2408,N_2431);
and U2479 (N_2479,N_2460,N_2453);
nand U2480 (N_2480,N_2458,N_2469);
nor U2481 (N_2481,N_2419,N_2444);
nor U2482 (N_2482,N_2424,N_2445);
or U2483 (N_2483,N_2450,N_2425);
nand U2484 (N_2484,N_2401,N_2432);
or U2485 (N_2485,N_2446,N_2433);
and U2486 (N_2486,N_2402,N_2407);
and U2487 (N_2487,N_2451,N_2442);
nand U2488 (N_2488,N_2437,N_2435);
nor U2489 (N_2489,N_2473,N_2455);
and U2490 (N_2490,N_2434,N_2454);
nor U2491 (N_2491,N_2404,N_2436);
or U2492 (N_2492,N_2406,N_2418);
or U2493 (N_2493,N_2461,N_2405);
and U2494 (N_2494,N_2420,N_2466);
nand U2495 (N_2495,N_2449,N_2462);
and U2496 (N_2496,N_2463,N_2440);
and U2497 (N_2497,N_2467,N_2413);
or U2498 (N_2498,N_2412,N_2414);
nor U2499 (N_2499,N_2443,N_2456);
nor U2500 (N_2500,N_2468,N_2464);
nand U2501 (N_2501,N_2410,N_2459);
or U2502 (N_2502,N_2415,N_2403);
nor U2503 (N_2503,N_2429,N_2426);
nor U2504 (N_2504,N_2470,N_2439);
nand U2505 (N_2505,N_2428,N_2465);
nor U2506 (N_2506,N_2438,N_2452);
and U2507 (N_2507,N_2474,N_2416);
nand U2508 (N_2508,N_2421,N_2417);
and U2509 (N_2509,N_2400,N_2441);
nand U2510 (N_2510,N_2448,N_2472);
nand U2511 (N_2511,N_2471,N_2409);
nand U2512 (N_2512,N_2427,N_2443);
or U2513 (N_2513,N_2453,N_2474);
and U2514 (N_2514,N_2442,N_2406);
nand U2515 (N_2515,N_2421,N_2462);
nand U2516 (N_2516,N_2463,N_2438);
nor U2517 (N_2517,N_2441,N_2462);
or U2518 (N_2518,N_2422,N_2458);
xnor U2519 (N_2519,N_2447,N_2422);
nor U2520 (N_2520,N_2431,N_2465);
and U2521 (N_2521,N_2429,N_2418);
nor U2522 (N_2522,N_2442,N_2415);
nor U2523 (N_2523,N_2412,N_2461);
nand U2524 (N_2524,N_2423,N_2456);
or U2525 (N_2525,N_2400,N_2402);
nor U2526 (N_2526,N_2459,N_2467);
and U2527 (N_2527,N_2401,N_2409);
or U2528 (N_2528,N_2400,N_2431);
nor U2529 (N_2529,N_2455,N_2418);
and U2530 (N_2530,N_2467,N_2408);
nand U2531 (N_2531,N_2457,N_2465);
nand U2532 (N_2532,N_2425,N_2401);
and U2533 (N_2533,N_2427,N_2422);
or U2534 (N_2534,N_2450,N_2412);
nand U2535 (N_2535,N_2412,N_2429);
nor U2536 (N_2536,N_2468,N_2409);
and U2537 (N_2537,N_2467,N_2430);
nor U2538 (N_2538,N_2435,N_2400);
and U2539 (N_2539,N_2404,N_2427);
xor U2540 (N_2540,N_2453,N_2466);
nand U2541 (N_2541,N_2403,N_2401);
and U2542 (N_2542,N_2437,N_2434);
nand U2543 (N_2543,N_2404,N_2429);
or U2544 (N_2544,N_2408,N_2462);
nand U2545 (N_2545,N_2417,N_2437);
nand U2546 (N_2546,N_2433,N_2452);
nand U2547 (N_2547,N_2412,N_2442);
nand U2548 (N_2548,N_2423,N_2465);
nand U2549 (N_2549,N_2435,N_2414);
or U2550 (N_2550,N_2531,N_2523);
or U2551 (N_2551,N_2510,N_2537);
nand U2552 (N_2552,N_2539,N_2543);
nor U2553 (N_2553,N_2522,N_2506);
or U2554 (N_2554,N_2535,N_2492);
and U2555 (N_2555,N_2482,N_2478);
nor U2556 (N_2556,N_2538,N_2509);
nand U2557 (N_2557,N_2485,N_2475);
or U2558 (N_2558,N_2484,N_2507);
nand U2559 (N_2559,N_2513,N_2521);
and U2560 (N_2560,N_2483,N_2514);
and U2561 (N_2561,N_2545,N_2501);
nand U2562 (N_2562,N_2527,N_2549);
or U2563 (N_2563,N_2520,N_2479);
or U2564 (N_2564,N_2536,N_2491);
nand U2565 (N_2565,N_2493,N_2533);
nor U2566 (N_2566,N_2502,N_2548);
nand U2567 (N_2567,N_2498,N_2499);
nand U2568 (N_2568,N_2525,N_2541);
or U2569 (N_2569,N_2490,N_2497);
and U2570 (N_2570,N_2504,N_2517);
nand U2571 (N_2571,N_2519,N_2528);
and U2572 (N_2572,N_2547,N_2532);
nor U2573 (N_2573,N_2489,N_2546);
nand U2574 (N_2574,N_2544,N_2496);
or U2575 (N_2575,N_2516,N_2542);
nand U2576 (N_2576,N_2534,N_2511);
and U2577 (N_2577,N_2526,N_2524);
or U2578 (N_2578,N_2503,N_2481);
or U2579 (N_2579,N_2495,N_2515);
nand U2580 (N_2580,N_2530,N_2500);
nor U2581 (N_2581,N_2480,N_2486);
and U2582 (N_2582,N_2512,N_2477);
or U2583 (N_2583,N_2487,N_2508);
or U2584 (N_2584,N_2518,N_2540);
or U2585 (N_2585,N_2494,N_2505);
or U2586 (N_2586,N_2476,N_2529);
and U2587 (N_2587,N_2488,N_2502);
nor U2588 (N_2588,N_2549,N_2476);
and U2589 (N_2589,N_2509,N_2486);
nor U2590 (N_2590,N_2541,N_2478);
or U2591 (N_2591,N_2548,N_2512);
and U2592 (N_2592,N_2491,N_2508);
nand U2593 (N_2593,N_2481,N_2509);
nor U2594 (N_2594,N_2506,N_2538);
nand U2595 (N_2595,N_2490,N_2499);
nor U2596 (N_2596,N_2535,N_2523);
xnor U2597 (N_2597,N_2513,N_2516);
nand U2598 (N_2598,N_2544,N_2543);
nor U2599 (N_2599,N_2533,N_2511);
and U2600 (N_2600,N_2548,N_2533);
or U2601 (N_2601,N_2493,N_2507);
and U2602 (N_2602,N_2531,N_2518);
and U2603 (N_2603,N_2523,N_2526);
and U2604 (N_2604,N_2535,N_2493);
nor U2605 (N_2605,N_2480,N_2542);
nand U2606 (N_2606,N_2531,N_2477);
nor U2607 (N_2607,N_2515,N_2503);
or U2608 (N_2608,N_2501,N_2482);
nor U2609 (N_2609,N_2524,N_2496);
and U2610 (N_2610,N_2487,N_2493);
and U2611 (N_2611,N_2540,N_2500);
nand U2612 (N_2612,N_2545,N_2528);
xnor U2613 (N_2613,N_2512,N_2491);
and U2614 (N_2614,N_2521,N_2524);
or U2615 (N_2615,N_2529,N_2531);
nand U2616 (N_2616,N_2516,N_2487);
or U2617 (N_2617,N_2532,N_2519);
and U2618 (N_2618,N_2545,N_2494);
and U2619 (N_2619,N_2537,N_2496);
nand U2620 (N_2620,N_2538,N_2514);
nor U2621 (N_2621,N_2505,N_2487);
and U2622 (N_2622,N_2502,N_2519);
or U2623 (N_2623,N_2505,N_2519);
or U2624 (N_2624,N_2539,N_2487);
or U2625 (N_2625,N_2584,N_2607);
nor U2626 (N_2626,N_2615,N_2595);
and U2627 (N_2627,N_2573,N_2561);
and U2628 (N_2628,N_2623,N_2599);
and U2629 (N_2629,N_2596,N_2578);
nand U2630 (N_2630,N_2594,N_2581);
or U2631 (N_2631,N_2583,N_2574);
and U2632 (N_2632,N_2557,N_2559);
or U2633 (N_2633,N_2603,N_2586);
or U2634 (N_2634,N_2554,N_2562);
nand U2635 (N_2635,N_2566,N_2568);
nor U2636 (N_2636,N_2567,N_2553);
and U2637 (N_2637,N_2597,N_2592);
nor U2638 (N_2638,N_2616,N_2598);
nor U2639 (N_2639,N_2564,N_2591);
or U2640 (N_2640,N_2622,N_2612);
nor U2641 (N_2641,N_2570,N_2608);
nor U2642 (N_2642,N_2618,N_2609);
nand U2643 (N_2643,N_2606,N_2600);
or U2644 (N_2644,N_2556,N_2621);
and U2645 (N_2645,N_2613,N_2582);
nor U2646 (N_2646,N_2602,N_2577);
nor U2647 (N_2647,N_2575,N_2558);
nand U2648 (N_2648,N_2551,N_2614);
and U2649 (N_2649,N_2589,N_2605);
nor U2650 (N_2650,N_2619,N_2611);
or U2651 (N_2651,N_2601,N_2587);
nand U2652 (N_2652,N_2565,N_2590);
nand U2653 (N_2653,N_2604,N_2572);
nor U2654 (N_2654,N_2563,N_2555);
and U2655 (N_2655,N_2593,N_2560);
nor U2656 (N_2656,N_2580,N_2624);
and U2657 (N_2657,N_2552,N_2617);
nor U2658 (N_2658,N_2571,N_2585);
nand U2659 (N_2659,N_2588,N_2576);
nor U2660 (N_2660,N_2610,N_2569);
nand U2661 (N_2661,N_2620,N_2579);
nand U2662 (N_2662,N_2550,N_2603);
nor U2663 (N_2663,N_2617,N_2577);
or U2664 (N_2664,N_2597,N_2563);
nand U2665 (N_2665,N_2617,N_2572);
nor U2666 (N_2666,N_2559,N_2558);
nor U2667 (N_2667,N_2579,N_2557);
nand U2668 (N_2668,N_2614,N_2608);
nand U2669 (N_2669,N_2605,N_2614);
or U2670 (N_2670,N_2615,N_2611);
nand U2671 (N_2671,N_2567,N_2615);
or U2672 (N_2672,N_2581,N_2585);
or U2673 (N_2673,N_2619,N_2601);
and U2674 (N_2674,N_2592,N_2599);
nor U2675 (N_2675,N_2613,N_2554);
or U2676 (N_2676,N_2606,N_2611);
or U2677 (N_2677,N_2579,N_2601);
and U2678 (N_2678,N_2605,N_2555);
and U2679 (N_2679,N_2619,N_2607);
or U2680 (N_2680,N_2586,N_2612);
or U2681 (N_2681,N_2621,N_2596);
nand U2682 (N_2682,N_2556,N_2551);
nand U2683 (N_2683,N_2587,N_2583);
nand U2684 (N_2684,N_2597,N_2584);
and U2685 (N_2685,N_2550,N_2601);
nor U2686 (N_2686,N_2604,N_2621);
nor U2687 (N_2687,N_2605,N_2574);
and U2688 (N_2688,N_2579,N_2589);
and U2689 (N_2689,N_2567,N_2601);
and U2690 (N_2690,N_2607,N_2564);
nor U2691 (N_2691,N_2574,N_2593);
nand U2692 (N_2692,N_2559,N_2554);
or U2693 (N_2693,N_2616,N_2554);
and U2694 (N_2694,N_2588,N_2559);
nor U2695 (N_2695,N_2593,N_2569);
nand U2696 (N_2696,N_2615,N_2554);
and U2697 (N_2697,N_2552,N_2604);
nand U2698 (N_2698,N_2562,N_2556);
or U2699 (N_2699,N_2604,N_2582);
nor U2700 (N_2700,N_2647,N_2643);
or U2701 (N_2701,N_2652,N_2675);
nand U2702 (N_2702,N_2674,N_2698);
or U2703 (N_2703,N_2661,N_2654);
nor U2704 (N_2704,N_2628,N_2683);
or U2705 (N_2705,N_2638,N_2676);
or U2706 (N_2706,N_2670,N_2692);
nand U2707 (N_2707,N_2679,N_2663);
and U2708 (N_2708,N_2671,N_2686);
nand U2709 (N_2709,N_2688,N_2699);
or U2710 (N_2710,N_2627,N_2687);
nand U2711 (N_2711,N_2629,N_2660);
nor U2712 (N_2712,N_2649,N_2639);
nand U2713 (N_2713,N_2693,N_2642);
nand U2714 (N_2714,N_2681,N_2672);
nand U2715 (N_2715,N_2678,N_2684);
nor U2716 (N_2716,N_2685,N_2697);
or U2717 (N_2717,N_2631,N_2650);
or U2718 (N_2718,N_2656,N_2634);
nand U2719 (N_2719,N_2648,N_2651);
nand U2720 (N_2720,N_2696,N_2667);
nor U2721 (N_2721,N_2680,N_2633);
nand U2722 (N_2722,N_2662,N_2626);
or U2723 (N_2723,N_2635,N_2636);
xnor U2724 (N_2724,N_2646,N_2694);
or U2725 (N_2725,N_2640,N_2695);
nor U2726 (N_2726,N_2666,N_2658);
nor U2727 (N_2727,N_2655,N_2659);
nor U2728 (N_2728,N_2641,N_2689);
nand U2729 (N_2729,N_2625,N_2632);
and U2730 (N_2730,N_2677,N_2669);
and U2731 (N_2731,N_2665,N_2637);
nor U2732 (N_2732,N_2653,N_2690);
nand U2733 (N_2733,N_2691,N_2645);
nor U2734 (N_2734,N_2657,N_2668);
and U2735 (N_2735,N_2664,N_2673);
and U2736 (N_2736,N_2682,N_2644);
nand U2737 (N_2737,N_2630,N_2699);
or U2738 (N_2738,N_2647,N_2652);
nor U2739 (N_2739,N_2667,N_2646);
or U2740 (N_2740,N_2651,N_2696);
nand U2741 (N_2741,N_2634,N_2689);
nor U2742 (N_2742,N_2646,N_2661);
nand U2743 (N_2743,N_2632,N_2627);
and U2744 (N_2744,N_2695,N_2672);
nor U2745 (N_2745,N_2684,N_2625);
and U2746 (N_2746,N_2641,N_2630);
nand U2747 (N_2747,N_2678,N_2655);
nor U2748 (N_2748,N_2646,N_2665);
nor U2749 (N_2749,N_2694,N_2674);
nor U2750 (N_2750,N_2696,N_2689);
nor U2751 (N_2751,N_2626,N_2648);
nor U2752 (N_2752,N_2642,N_2640);
nand U2753 (N_2753,N_2660,N_2678);
and U2754 (N_2754,N_2651,N_2634);
nor U2755 (N_2755,N_2694,N_2670);
nor U2756 (N_2756,N_2658,N_2636);
nand U2757 (N_2757,N_2687,N_2670);
and U2758 (N_2758,N_2631,N_2698);
and U2759 (N_2759,N_2697,N_2654);
nor U2760 (N_2760,N_2654,N_2663);
nor U2761 (N_2761,N_2675,N_2637);
nor U2762 (N_2762,N_2632,N_2694);
and U2763 (N_2763,N_2669,N_2652);
nor U2764 (N_2764,N_2664,N_2625);
nand U2765 (N_2765,N_2671,N_2682);
nand U2766 (N_2766,N_2674,N_2627);
or U2767 (N_2767,N_2686,N_2646);
and U2768 (N_2768,N_2646,N_2627);
or U2769 (N_2769,N_2674,N_2653);
or U2770 (N_2770,N_2637,N_2679);
nor U2771 (N_2771,N_2647,N_2630);
nand U2772 (N_2772,N_2646,N_2631);
nor U2773 (N_2773,N_2677,N_2650);
and U2774 (N_2774,N_2658,N_2682);
or U2775 (N_2775,N_2726,N_2729);
nand U2776 (N_2776,N_2745,N_2723);
or U2777 (N_2777,N_2754,N_2734);
nand U2778 (N_2778,N_2764,N_2717);
or U2779 (N_2779,N_2701,N_2759);
and U2780 (N_2780,N_2702,N_2756);
nand U2781 (N_2781,N_2733,N_2735);
nor U2782 (N_2782,N_2766,N_2769);
nor U2783 (N_2783,N_2748,N_2763);
nor U2784 (N_2784,N_2770,N_2721);
nand U2785 (N_2785,N_2711,N_2713);
nor U2786 (N_2786,N_2738,N_2750);
nand U2787 (N_2787,N_2737,N_2742);
and U2788 (N_2788,N_2714,N_2749);
or U2789 (N_2789,N_2715,N_2725);
or U2790 (N_2790,N_2761,N_2716);
nand U2791 (N_2791,N_2762,N_2774);
nor U2792 (N_2792,N_2718,N_2719);
nand U2793 (N_2793,N_2758,N_2730);
nand U2794 (N_2794,N_2746,N_2705);
or U2795 (N_2795,N_2771,N_2751);
and U2796 (N_2796,N_2732,N_2743);
nand U2797 (N_2797,N_2740,N_2747);
or U2798 (N_2798,N_2760,N_2720);
and U2799 (N_2799,N_2700,N_2707);
nor U2800 (N_2800,N_2772,N_2724);
nor U2801 (N_2801,N_2706,N_2703);
and U2802 (N_2802,N_2727,N_2709);
and U2803 (N_2803,N_2712,N_2708);
nand U2804 (N_2804,N_2757,N_2767);
nand U2805 (N_2805,N_2722,N_2736);
xnor U2806 (N_2806,N_2753,N_2728);
nor U2807 (N_2807,N_2765,N_2755);
and U2808 (N_2808,N_2710,N_2744);
or U2809 (N_2809,N_2741,N_2768);
nand U2810 (N_2810,N_2731,N_2752);
nand U2811 (N_2811,N_2704,N_2739);
nand U2812 (N_2812,N_2773,N_2759);
or U2813 (N_2813,N_2744,N_2733);
and U2814 (N_2814,N_2751,N_2708);
and U2815 (N_2815,N_2747,N_2756);
or U2816 (N_2816,N_2761,N_2746);
and U2817 (N_2817,N_2765,N_2727);
and U2818 (N_2818,N_2771,N_2713);
nor U2819 (N_2819,N_2730,N_2729);
or U2820 (N_2820,N_2707,N_2726);
nor U2821 (N_2821,N_2745,N_2724);
nand U2822 (N_2822,N_2703,N_2716);
or U2823 (N_2823,N_2724,N_2714);
nand U2824 (N_2824,N_2707,N_2756);
nand U2825 (N_2825,N_2758,N_2743);
and U2826 (N_2826,N_2769,N_2756);
or U2827 (N_2827,N_2761,N_2751);
nor U2828 (N_2828,N_2714,N_2726);
or U2829 (N_2829,N_2726,N_2759);
nor U2830 (N_2830,N_2730,N_2749);
and U2831 (N_2831,N_2762,N_2729);
and U2832 (N_2832,N_2724,N_2721);
and U2833 (N_2833,N_2719,N_2713);
and U2834 (N_2834,N_2715,N_2703);
or U2835 (N_2835,N_2758,N_2709);
and U2836 (N_2836,N_2738,N_2749);
or U2837 (N_2837,N_2764,N_2733);
and U2838 (N_2838,N_2722,N_2707);
nor U2839 (N_2839,N_2770,N_2753);
or U2840 (N_2840,N_2771,N_2702);
nor U2841 (N_2841,N_2729,N_2738);
nand U2842 (N_2842,N_2770,N_2712);
nand U2843 (N_2843,N_2707,N_2760);
and U2844 (N_2844,N_2770,N_2711);
nor U2845 (N_2845,N_2762,N_2770);
and U2846 (N_2846,N_2757,N_2748);
or U2847 (N_2847,N_2752,N_2709);
or U2848 (N_2848,N_2711,N_2724);
nor U2849 (N_2849,N_2734,N_2762);
nor U2850 (N_2850,N_2777,N_2792);
nand U2851 (N_2851,N_2807,N_2784);
and U2852 (N_2852,N_2811,N_2814);
nor U2853 (N_2853,N_2823,N_2796);
nand U2854 (N_2854,N_2810,N_2795);
nor U2855 (N_2855,N_2776,N_2826);
nor U2856 (N_2856,N_2786,N_2835);
or U2857 (N_2857,N_2779,N_2843);
nand U2858 (N_2858,N_2824,N_2829);
or U2859 (N_2859,N_2831,N_2830);
and U2860 (N_2860,N_2803,N_2788);
nand U2861 (N_2861,N_2790,N_2794);
nand U2862 (N_2862,N_2842,N_2801);
nor U2863 (N_2863,N_2775,N_2781);
nand U2864 (N_2864,N_2839,N_2833);
or U2865 (N_2865,N_2804,N_2845);
nor U2866 (N_2866,N_2782,N_2819);
or U2867 (N_2867,N_2780,N_2806);
or U2868 (N_2868,N_2805,N_2822);
and U2869 (N_2869,N_2820,N_2847);
nand U2870 (N_2870,N_2838,N_2808);
and U2871 (N_2871,N_2837,N_2849);
nand U2872 (N_2872,N_2813,N_2799);
and U2873 (N_2873,N_2840,N_2798);
nor U2874 (N_2874,N_2778,N_2791);
nand U2875 (N_2875,N_2821,N_2817);
nand U2876 (N_2876,N_2834,N_2802);
nor U2877 (N_2877,N_2793,N_2841);
xnor U2878 (N_2878,N_2844,N_2848);
nor U2879 (N_2879,N_2785,N_2836);
or U2880 (N_2880,N_2816,N_2789);
and U2881 (N_2881,N_2832,N_2825);
or U2882 (N_2882,N_2783,N_2787);
nand U2883 (N_2883,N_2818,N_2809);
or U2884 (N_2884,N_2828,N_2815);
nand U2885 (N_2885,N_2800,N_2827);
or U2886 (N_2886,N_2812,N_2846);
and U2887 (N_2887,N_2797,N_2813);
nand U2888 (N_2888,N_2846,N_2810);
nor U2889 (N_2889,N_2811,N_2846);
or U2890 (N_2890,N_2776,N_2791);
and U2891 (N_2891,N_2829,N_2788);
and U2892 (N_2892,N_2843,N_2800);
nor U2893 (N_2893,N_2833,N_2815);
nor U2894 (N_2894,N_2826,N_2844);
or U2895 (N_2895,N_2835,N_2842);
nand U2896 (N_2896,N_2787,N_2807);
nor U2897 (N_2897,N_2827,N_2825);
nor U2898 (N_2898,N_2809,N_2837);
nand U2899 (N_2899,N_2822,N_2831);
or U2900 (N_2900,N_2786,N_2843);
or U2901 (N_2901,N_2803,N_2839);
or U2902 (N_2902,N_2847,N_2804);
or U2903 (N_2903,N_2797,N_2824);
or U2904 (N_2904,N_2839,N_2829);
nor U2905 (N_2905,N_2819,N_2821);
nor U2906 (N_2906,N_2840,N_2830);
nor U2907 (N_2907,N_2819,N_2789);
nor U2908 (N_2908,N_2815,N_2844);
nor U2909 (N_2909,N_2788,N_2833);
and U2910 (N_2910,N_2827,N_2790);
nor U2911 (N_2911,N_2822,N_2799);
or U2912 (N_2912,N_2819,N_2820);
and U2913 (N_2913,N_2781,N_2831);
nor U2914 (N_2914,N_2810,N_2847);
nor U2915 (N_2915,N_2835,N_2803);
or U2916 (N_2916,N_2775,N_2809);
or U2917 (N_2917,N_2832,N_2829);
nand U2918 (N_2918,N_2845,N_2808);
and U2919 (N_2919,N_2785,N_2823);
nor U2920 (N_2920,N_2789,N_2837);
and U2921 (N_2921,N_2791,N_2843);
nor U2922 (N_2922,N_2841,N_2831);
or U2923 (N_2923,N_2827,N_2793);
and U2924 (N_2924,N_2776,N_2843);
nor U2925 (N_2925,N_2890,N_2856);
nor U2926 (N_2926,N_2923,N_2893);
nand U2927 (N_2927,N_2883,N_2892);
nor U2928 (N_2928,N_2870,N_2910);
nor U2929 (N_2929,N_2908,N_2859);
and U2930 (N_2930,N_2898,N_2888);
nor U2931 (N_2931,N_2924,N_2904);
or U2932 (N_2932,N_2884,N_2863);
and U2933 (N_2933,N_2868,N_2912);
nor U2934 (N_2934,N_2920,N_2918);
nor U2935 (N_2935,N_2894,N_2913);
and U2936 (N_2936,N_2907,N_2903);
or U2937 (N_2937,N_2876,N_2861);
or U2938 (N_2938,N_2916,N_2895);
nor U2939 (N_2939,N_2864,N_2886);
or U2940 (N_2940,N_2889,N_2911);
and U2941 (N_2941,N_2882,N_2867);
nor U2942 (N_2942,N_2854,N_2857);
nand U2943 (N_2943,N_2852,N_2906);
nor U2944 (N_2944,N_2875,N_2891);
or U2945 (N_2945,N_2860,N_2914);
or U2946 (N_2946,N_2905,N_2879);
nand U2947 (N_2947,N_2872,N_2851);
and U2948 (N_2948,N_2922,N_2871);
or U2949 (N_2949,N_2865,N_2917);
nor U2950 (N_2950,N_2885,N_2869);
nor U2951 (N_2951,N_2881,N_2866);
and U2952 (N_2952,N_2873,N_2850);
nand U2953 (N_2953,N_2862,N_2878);
nand U2954 (N_2954,N_2921,N_2899);
nand U2955 (N_2955,N_2915,N_2902);
or U2956 (N_2956,N_2901,N_2877);
and U2957 (N_2957,N_2900,N_2909);
or U2958 (N_2958,N_2919,N_2896);
nand U2959 (N_2959,N_2874,N_2897);
and U2960 (N_2960,N_2853,N_2880);
or U2961 (N_2961,N_2855,N_2887);
nand U2962 (N_2962,N_2858,N_2901);
nand U2963 (N_2963,N_2910,N_2893);
nor U2964 (N_2964,N_2919,N_2911);
nor U2965 (N_2965,N_2877,N_2887);
nand U2966 (N_2966,N_2857,N_2882);
nor U2967 (N_2967,N_2867,N_2909);
nor U2968 (N_2968,N_2905,N_2866);
and U2969 (N_2969,N_2857,N_2893);
and U2970 (N_2970,N_2853,N_2881);
and U2971 (N_2971,N_2901,N_2892);
nand U2972 (N_2972,N_2871,N_2921);
nor U2973 (N_2973,N_2922,N_2892);
and U2974 (N_2974,N_2857,N_2894);
and U2975 (N_2975,N_2890,N_2915);
nand U2976 (N_2976,N_2871,N_2884);
nand U2977 (N_2977,N_2916,N_2855);
nor U2978 (N_2978,N_2893,N_2874);
or U2979 (N_2979,N_2886,N_2905);
and U2980 (N_2980,N_2885,N_2874);
nor U2981 (N_2981,N_2923,N_2880);
and U2982 (N_2982,N_2869,N_2871);
or U2983 (N_2983,N_2856,N_2909);
nor U2984 (N_2984,N_2890,N_2865);
or U2985 (N_2985,N_2854,N_2880);
and U2986 (N_2986,N_2856,N_2879);
nor U2987 (N_2987,N_2883,N_2919);
or U2988 (N_2988,N_2875,N_2908);
or U2989 (N_2989,N_2912,N_2876);
or U2990 (N_2990,N_2898,N_2882);
and U2991 (N_2991,N_2851,N_2907);
and U2992 (N_2992,N_2916,N_2877);
or U2993 (N_2993,N_2884,N_2917);
nor U2994 (N_2994,N_2852,N_2888);
or U2995 (N_2995,N_2907,N_2853);
nor U2996 (N_2996,N_2903,N_2852);
or U2997 (N_2997,N_2917,N_2895);
nor U2998 (N_2998,N_2900,N_2855);
nor U2999 (N_2999,N_2901,N_2887);
nand UO_0 (O_0,N_2983,N_2979);
nor UO_1 (O_1,N_2931,N_2992);
nand UO_2 (O_2,N_2968,N_2941);
xor UO_3 (O_3,N_2993,N_2974);
nand UO_4 (O_4,N_2995,N_2972);
and UO_5 (O_5,N_2945,N_2960);
or UO_6 (O_6,N_2997,N_2929);
nand UO_7 (O_7,N_2950,N_2999);
and UO_8 (O_8,N_2935,N_2985);
nor UO_9 (O_9,N_2963,N_2980);
or UO_10 (O_10,N_2933,N_2961);
nand UO_11 (O_11,N_2973,N_2952);
nor UO_12 (O_12,N_2943,N_2932);
nor UO_13 (O_13,N_2956,N_2962);
and UO_14 (O_14,N_2965,N_2936);
or UO_15 (O_15,N_2994,N_2971);
nand UO_16 (O_16,N_2955,N_2990);
nand UO_17 (O_17,N_2926,N_2967);
or UO_18 (O_18,N_2937,N_2951);
or UO_19 (O_19,N_2940,N_2976);
and UO_20 (O_20,N_2977,N_2925);
and UO_21 (O_21,N_2942,N_2930);
nor UO_22 (O_22,N_2988,N_2986);
nand UO_23 (O_23,N_2970,N_2927);
or UO_24 (O_24,N_2928,N_2998);
nand UO_25 (O_25,N_2948,N_2953);
or UO_26 (O_26,N_2944,N_2969);
nor UO_27 (O_27,N_2975,N_2982);
nor UO_28 (O_28,N_2958,N_2938);
or UO_29 (O_29,N_2939,N_2959);
nand UO_30 (O_30,N_2966,N_2989);
or UO_31 (O_31,N_2949,N_2947);
nor UO_32 (O_32,N_2954,N_2964);
and UO_33 (O_33,N_2978,N_2957);
and UO_34 (O_34,N_2996,N_2984);
nor UO_35 (O_35,N_2987,N_2934);
or UO_36 (O_36,N_2946,N_2981);
or UO_37 (O_37,N_2991,N_2990);
and UO_38 (O_38,N_2939,N_2965);
nand UO_39 (O_39,N_2977,N_2941);
nor UO_40 (O_40,N_2938,N_2954);
nand UO_41 (O_41,N_2936,N_2967);
and UO_42 (O_42,N_2957,N_2964);
nand UO_43 (O_43,N_2956,N_2976);
or UO_44 (O_44,N_2987,N_2989);
or UO_45 (O_45,N_2940,N_2934);
nor UO_46 (O_46,N_2925,N_2975);
or UO_47 (O_47,N_2976,N_2930);
nand UO_48 (O_48,N_2957,N_2970);
nand UO_49 (O_49,N_2998,N_2992);
nor UO_50 (O_50,N_2971,N_2977);
nor UO_51 (O_51,N_2980,N_2930);
and UO_52 (O_52,N_2972,N_2928);
nor UO_53 (O_53,N_2938,N_2955);
or UO_54 (O_54,N_2946,N_2948);
nor UO_55 (O_55,N_2989,N_2957);
and UO_56 (O_56,N_2930,N_2970);
and UO_57 (O_57,N_2993,N_2965);
nor UO_58 (O_58,N_2928,N_2965);
nand UO_59 (O_59,N_2986,N_2997);
and UO_60 (O_60,N_2938,N_2932);
and UO_61 (O_61,N_2973,N_2956);
nand UO_62 (O_62,N_2950,N_2968);
or UO_63 (O_63,N_2930,N_2953);
nand UO_64 (O_64,N_2957,N_2951);
and UO_65 (O_65,N_2976,N_2989);
xor UO_66 (O_66,N_2933,N_2926);
nor UO_67 (O_67,N_2927,N_2997);
nand UO_68 (O_68,N_2962,N_2981);
and UO_69 (O_69,N_2931,N_2993);
and UO_70 (O_70,N_2998,N_2953);
nand UO_71 (O_71,N_2959,N_2956);
nand UO_72 (O_72,N_2995,N_2954);
nor UO_73 (O_73,N_2963,N_2998);
and UO_74 (O_74,N_2936,N_2944);
nor UO_75 (O_75,N_2998,N_2966);
or UO_76 (O_76,N_2979,N_2935);
and UO_77 (O_77,N_2963,N_2975);
nor UO_78 (O_78,N_2970,N_2972);
nand UO_79 (O_79,N_2954,N_2989);
or UO_80 (O_80,N_2970,N_2953);
xnor UO_81 (O_81,N_2983,N_2942);
or UO_82 (O_82,N_2976,N_2960);
or UO_83 (O_83,N_2926,N_2965);
or UO_84 (O_84,N_2952,N_2930);
or UO_85 (O_85,N_2978,N_2976);
and UO_86 (O_86,N_2936,N_2996);
or UO_87 (O_87,N_2938,N_2940);
nor UO_88 (O_88,N_2933,N_2977);
nand UO_89 (O_89,N_2944,N_2988);
nor UO_90 (O_90,N_2929,N_2954);
nand UO_91 (O_91,N_2927,N_2962);
or UO_92 (O_92,N_2996,N_2999);
or UO_93 (O_93,N_2999,N_2989);
nand UO_94 (O_94,N_2976,N_2955);
or UO_95 (O_95,N_2943,N_2962);
or UO_96 (O_96,N_2969,N_2931);
or UO_97 (O_97,N_2952,N_2995);
nand UO_98 (O_98,N_2947,N_2957);
or UO_99 (O_99,N_2932,N_2973);
nand UO_100 (O_100,N_2950,N_2957);
and UO_101 (O_101,N_2982,N_2967);
or UO_102 (O_102,N_2970,N_2977);
and UO_103 (O_103,N_2988,N_2991);
or UO_104 (O_104,N_2969,N_2940);
nor UO_105 (O_105,N_2950,N_2973);
or UO_106 (O_106,N_2979,N_2928);
nand UO_107 (O_107,N_2944,N_2946);
or UO_108 (O_108,N_2948,N_2991);
nor UO_109 (O_109,N_2958,N_2966);
or UO_110 (O_110,N_2961,N_2934);
nor UO_111 (O_111,N_2998,N_2949);
nand UO_112 (O_112,N_2955,N_2985);
nor UO_113 (O_113,N_2970,N_2967);
nand UO_114 (O_114,N_2995,N_2944);
nor UO_115 (O_115,N_2972,N_2990);
nand UO_116 (O_116,N_2939,N_2952);
nand UO_117 (O_117,N_2977,N_2927);
and UO_118 (O_118,N_2987,N_2971);
or UO_119 (O_119,N_2947,N_2926);
nor UO_120 (O_120,N_2925,N_2991);
and UO_121 (O_121,N_2994,N_2977);
and UO_122 (O_122,N_2935,N_2999);
and UO_123 (O_123,N_2931,N_2958);
nor UO_124 (O_124,N_2926,N_2943);
nor UO_125 (O_125,N_2948,N_2965);
and UO_126 (O_126,N_2980,N_2971);
nand UO_127 (O_127,N_2994,N_2947);
and UO_128 (O_128,N_2978,N_2963);
nor UO_129 (O_129,N_2934,N_2980);
or UO_130 (O_130,N_2987,N_2955);
and UO_131 (O_131,N_2950,N_2955);
xor UO_132 (O_132,N_2945,N_2975);
nand UO_133 (O_133,N_2942,N_2952);
or UO_134 (O_134,N_2979,N_2977);
nand UO_135 (O_135,N_2976,N_2953);
nor UO_136 (O_136,N_2985,N_2961);
or UO_137 (O_137,N_2967,N_2974);
nor UO_138 (O_138,N_2967,N_2935);
or UO_139 (O_139,N_2967,N_2938);
nor UO_140 (O_140,N_2995,N_2931);
or UO_141 (O_141,N_2942,N_2951);
nor UO_142 (O_142,N_2952,N_2949);
nand UO_143 (O_143,N_2974,N_2942);
or UO_144 (O_144,N_2935,N_2974);
or UO_145 (O_145,N_2932,N_2949);
nand UO_146 (O_146,N_2954,N_2957);
or UO_147 (O_147,N_2972,N_2932);
and UO_148 (O_148,N_2969,N_2942);
and UO_149 (O_149,N_2966,N_2936);
and UO_150 (O_150,N_2935,N_2972);
nand UO_151 (O_151,N_2977,N_2964);
and UO_152 (O_152,N_2991,N_2938);
nor UO_153 (O_153,N_2958,N_2988);
nor UO_154 (O_154,N_2953,N_2991);
or UO_155 (O_155,N_2967,N_2957);
nor UO_156 (O_156,N_2950,N_2982);
or UO_157 (O_157,N_2986,N_2972);
and UO_158 (O_158,N_2936,N_2986);
and UO_159 (O_159,N_2964,N_2969);
nand UO_160 (O_160,N_2958,N_2974);
or UO_161 (O_161,N_2956,N_2989);
or UO_162 (O_162,N_2928,N_2999);
nand UO_163 (O_163,N_2936,N_2981);
or UO_164 (O_164,N_2945,N_2993);
and UO_165 (O_165,N_2992,N_2984);
nor UO_166 (O_166,N_2930,N_2929);
nor UO_167 (O_167,N_2929,N_2934);
and UO_168 (O_168,N_2978,N_2992);
nor UO_169 (O_169,N_2948,N_2935);
nand UO_170 (O_170,N_2997,N_2935);
nand UO_171 (O_171,N_2929,N_2953);
nor UO_172 (O_172,N_2935,N_2960);
and UO_173 (O_173,N_2960,N_2975);
nand UO_174 (O_174,N_2968,N_2972);
nor UO_175 (O_175,N_2984,N_2994);
or UO_176 (O_176,N_2938,N_2973);
or UO_177 (O_177,N_2975,N_2930);
nand UO_178 (O_178,N_2967,N_2937);
nand UO_179 (O_179,N_2953,N_2966);
or UO_180 (O_180,N_2996,N_2928);
nand UO_181 (O_181,N_2949,N_2991);
or UO_182 (O_182,N_2993,N_2953);
nand UO_183 (O_183,N_2927,N_2985);
nand UO_184 (O_184,N_2993,N_2989);
or UO_185 (O_185,N_2957,N_2938);
xnor UO_186 (O_186,N_2928,N_2925);
and UO_187 (O_187,N_2987,N_2996);
nand UO_188 (O_188,N_2932,N_2955);
or UO_189 (O_189,N_2984,N_2926);
nor UO_190 (O_190,N_2940,N_2961);
nand UO_191 (O_191,N_2939,N_2937);
or UO_192 (O_192,N_2943,N_2959);
xor UO_193 (O_193,N_2931,N_2932);
and UO_194 (O_194,N_2935,N_2944);
and UO_195 (O_195,N_2954,N_2960);
nor UO_196 (O_196,N_2935,N_2958);
nor UO_197 (O_197,N_2979,N_2991);
nor UO_198 (O_198,N_2946,N_2943);
and UO_199 (O_199,N_2953,N_2935);
or UO_200 (O_200,N_2955,N_2999);
nor UO_201 (O_201,N_2940,N_2975);
and UO_202 (O_202,N_2980,N_2972);
nand UO_203 (O_203,N_2953,N_2986);
or UO_204 (O_204,N_2968,N_2929);
nor UO_205 (O_205,N_2945,N_2991);
nand UO_206 (O_206,N_2930,N_2936);
nor UO_207 (O_207,N_2952,N_2951);
nand UO_208 (O_208,N_2978,N_2953);
or UO_209 (O_209,N_2953,N_2983);
or UO_210 (O_210,N_2980,N_2966);
nand UO_211 (O_211,N_2929,N_2946);
and UO_212 (O_212,N_2930,N_2947);
or UO_213 (O_213,N_2943,N_2983);
nor UO_214 (O_214,N_2936,N_2994);
or UO_215 (O_215,N_2973,N_2986);
and UO_216 (O_216,N_2988,N_2953);
or UO_217 (O_217,N_2926,N_2987);
and UO_218 (O_218,N_2974,N_2980);
nand UO_219 (O_219,N_2927,N_2936);
nand UO_220 (O_220,N_2958,N_2937);
and UO_221 (O_221,N_2929,N_2994);
or UO_222 (O_222,N_2955,N_2935);
nor UO_223 (O_223,N_2936,N_2937);
and UO_224 (O_224,N_2977,N_2959);
and UO_225 (O_225,N_2943,N_2987);
nand UO_226 (O_226,N_2930,N_2926);
nor UO_227 (O_227,N_2984,N_2969);
nor UO_228 (O_228,N_2996,N_2970);
or UO_229 (O_229,N_2970,N_2971);
nand UO_230 (O_230,N_2968,N_2926);
nor UO_231 (O_231,N_2975,N_2934);
and UO_232 (O_232,N_2941,N_2957);
and UO_233 (O_233,N_2955,N_2978);
nor UO_234 (O_234,N_2940,N_2957);
nand UO_235 (O_235,N_2941,N_2940);
or UO_236 (O_236,N_2965,N_2961);
nand UO_237 (O_237,N_2938,N_2949);
nand UO_238 (O_238,N_2928,N_2991);
and UO_239 (O_239,N_2933,N_2940);
or UO_240 (O_240,N_2995,N_2962);
nand UO_241 (O_241,N_2978,N_2986);
and UO_242 (O_242,N_2983,N_2944);
nor UO_243 (O_243,N_2973,N_2936);
and UO_244 (O_244,N_2957,N_2930);
nor UO_245 (O_245,N_2955,N_2927);
nor UO_246 (O_246,N_2978,N_2936);
nor UO_247 (O_247,N_2976,N_2946);
and UO_248 (O_248,N_2943,N_2940);
nor UO_249 (O_249,N_2951,N_2950);
nor UO_250 (O_250,N_2943,N_2947);
nand UO_251 (O_251,N_2956,N_2952);
nor UO_252 (O_252,N_2932,N_2958);
nand UO_253 (O_253,N_2977,N_2972);
or UO_254 (O_254,N_2976,N_2948);
nor UO_255 (O_255,N_2968,N_2988);
and UO_256 (O_256,N_2993,N_2956);
or UO_257 (O_257,N_2999,N_2933);
nand UO_258 (O_258,N_2925,N_2943);
nor UO_259 (O_259,N_2949,N_2956);
and UO_260 (O_260,N_2935,N_2970);
nand UO_261 (O_261,N_2997,N_2988);
or UO_262 (O_262,N_2925,N_2995);
or UO_263 (O_263,N_2947,N_2973);
xnor UO_264 (O_264,N_2993,N_2979);
and UO_265 (O_265,N_2986,N_2935);
nor UO_266 (O_266,N_2926,N_2954);
nand UO_267 (O_267,N_2927,N_2965);
or UO_268 (O_268,N_2935,N_2941);
nand UO_269 (O_269,N_2982,N_2936);
nand UO_270 (O_270,N_2933,N_2959);
or UO_271 (O_271,N_2975,N_2962);
nor UO_272 (O_272,N_2946,N_2931);
nor UO_273 (O_273,N_2946,N_2952);
and UO_274 (O_274,N_2926,N_2950);
and UO_275 (O_275,N_2953,N_2925);
nor UO_276 (O_276,N_2985,N_2970);
or UO_277 (O_277,N_2995,N_2987);
nor UO_278 (O_278,N_2972,N_2951);
nor UO_279 (O_279,N_2963,N_2948);
nor UO_280 (O_280,N_2955,N_2960);
and UO_281 (O_281,N_2940,N_2996);
nor UO_282 (O_282,N_2969,N_2925);
xnor UO_283 (O_283,N_2933,N_2936);
or UO_284 (O_284,N_2939,N_2927);
and UO_285 (O_285,N_2973,N_2982);
nor UO_286 (O_286,N_2982,N_2998);
and UO_287 (O_287,N_2929,N_2937);
and UO_288 (O_288,N_2972,N_2979);
or UO_289 (O_289,N_2935,N_2930);
nor UO_290 (O_290,N_2927,N_2999);
or UO_291 (O_291,N_2942,N_2933);
nor UO_292 (O_292,N_2963,N_2961);
nand UO_293 (O_293,N_2952,N_2937);
nor UO_294 (O_294,N_2985,N_2931);
nand UO_295 (O_295,N_2995,N_2936);
or UO_296 (O_296,N_2955,N_2966);
nand UO_297 (O_297,N_2939,N_2934);
nor UO_298 (O_298,N_2975,N_2953);
or UO_299 (O_299,N_2955,N_2984);
nand UO_300 (O_300,N_2949,N_2936);
and UO_301 (O_301,N_2962,N_2997);
or UO_302 (O_302,N_2957,N_2965);
nand UO_303 (O_303,N_2946,N_2938);
nand UO_304 (O_304,N_2952,N_2983);
nor UO_305 (O_305,N_2948,N_2980);
or UO_306 (O_306,N_2941,N_2976);
and UO_307 (O_307,N_2976,N_2987);
and UO_308 (O_308,N_2991,N_2946);
or UO_309 (O_309,N_2952,N_2927);
nor UO_310 (O_310,N_2941,N_2972);
nor UO_311 (O_311,N_2952,N_2996);
nor UO_312 (O_312,N_2967,N_2998);
or UO_313 (O_313,N_2997,N_2994);
nand UO_314 (O_314,N_2978,N_2946);
and UO_315 (O_315,N_2927,N_2934);
and UO_316 (O_316,N_2960,N_2989);
nor UO_317 (O_317,N_2969,N_2937);
nor UO_318 (O_318,N_2980,N_2993);
and UO_319 (O_319,N_2999,N_2962);
or UO_320 (O_320,N_2975,N_2947);
and UO_321 (O_321,N_2971,N_2964);
nor UO_322 (O_322,N_2972,N_2996);
nor UO_323 (O_323,N_2990,N_2978);
nand UO_324 (O_324,N_2971,N_2972);
and UO_325 (O_325,N_2967,N_2977);
nand UO_326 (O_326,N_2953,N_2990);
nand UO_327 (O_327,N_2964,N_2976);
and UO_328 (O_328,N_2980,N_2954);
nand UO_329 (O_329,N_2989,N_2990);
and UO_330 (O_330,N_2970,N_2976);
nand UO_331 (O_331,N_2995,N_2933);
nand UO_332 (O_332,N_2962,N_2955);
nor UO_333 (O_333,N_2999,N_2954);
and UO_334 (O_334,N_2994,N_2941);
or UO_335 (O_335,N_2961,N_2980);
or UO_336 (O_336,N_2966,N_2947);
nor UO_337 (O_337,N_2997,N_2976);
nand UO_338 (O_338,N_2938,N_2988);
nand UO_339 (O_339,N_2993,N_2947);
nor UO_340 (O_340,N_2945,N_2974);
or UO_341 (O_341,N_2947,N_2998);
or UO_342 (O_342,N_2929,N_2982);
or UO_343 (O_343,N_2955,N_2941);
nand UO_344 (O_344,N_2969,N_2939);
nor UO_345 (O_345,N_2987,N_2931);
or UO_346 (O_346,N_2958,N_2980);
nor UO_347 (O_347,N_2942,N_2949);
xnor UO_348 (O_348,N_2927,N_2996);
and UO_349 (O_349,N_2936,N_2984);
nor UO_350 (O_350,N_2996,N_2983);
nor UO_351 (O_351,N_2925,N_2947);
nand UO_352 (O_352,N_2979,N_2937);
nor UO_353 (O_353,N_2983,N_2960);
and UO_354 (O_354,N_2929,N_2991);
or UO_355 (O_355,N_2964,N_2974);
nor UO_356 (O_356,N_2980,N_2964);
nor UO_357 (O_357,N_2958,N_2998);
nand UO_358 (O_358,N_2991,N_2963);
and UO_359 (O_359,N_2948,N_2990);
nand UO_360 (O_360,N_2968,N_2999);
nand UO_361 (O_361,N_2949,N_2978);
or UO_362 (O_362,N_2930,N_2939);
and UO_363 (O_363,N_2976,N_2927);
and UO_364 (O_364,N_2937,N_2970);
or UO_365 (O_365,N_2946,N_2935);
xor UO_366 (O_366,N_2927,N_2953);
nand UO_367 (O_367,N_2980,N_2928);
or UO_368 (O_368,N_2972,N_2926);
xor UO_369 (O_369,N_2935,N_2925);
or UO_370 (O_370,N_2928,N_2977);
or UO_371 (O_371,N_2994,N_2992);
and UO_372 (O_372,N_2946,N_2992);
or UO_373 (O_373,N_2962,N_2952);
and UO_374 (O_374,N_2957,N_2946);
nor UO_375 (O_375,N_2948,N_2973);
nor UO_376 (O_376,N_2974,N_2996);
or UO_377 (O_377,N_2987,N_2949);
or UO_378 (O_378,N_2999,N_2943);
and UO_379 (O_379,N_2954,N_2982);
nand UO_380 (O_380,N_2951,N_2930);
nand UO_381 (O_381,N_2999,N_2930);
nand UO_382 (O_382,N_2963,N_2938);
and UO_383 (O_383,N_2943,N_2981);
nor UO_384 (O_384,N_2933,N_2925);
and UO_385 (O_385,N_2996,N_2925);
nand UO_386 (O_386,N_2961,N_2975);
and UO_387 (O_387,N_2933,N_2951);
nor UO_388 (O_388,N_2960,N_2965);
nor UO_389 (O_389,N_2972,N_2967);
nor UO_390 (O_390,N_2933,N_2957);
and UO_391 (O_391,N_2934,N_2937);
nor UO_392 (O_392,N_2943,N_2944);
nand UO_393 (O_393,N_2940,N_2931);
or UO_394 (O_394,N_2983,N_2963);
nor UO_395 (O_395,N_2952,N_2991);
or UO_396 (O_396,N_2966,N_2949);
nor UO_397 (O_397,N_2933,N_2992);
nor UO_398 (O_398,N_2967,N_2965);
and UO_399 (O_399,N_2970,N_2941);
xor UO_400 (O_400,N_2940,N_2926);
nor UO_401 (O_401,N_2975,N_2936);
nand UO_402 (O_402,N_2938,N_2997);
or UO_403 (O_403,N_2965,N_2985);
nor UO_404 (O_404,N_2988,N_2981);
nand UO_405 (O_405,N_2928,N_2988);
and UO_406 (O_406,N_2940,N_2987);
and UO_407 (O_407,N_2933,N_2958);
nand UO_408 (O_408,N_2951,N_2975);
and UO_409 (O_409,N_2937,N_2956);
or UO_410 (O_410,N_2989,N_2984);
nand UO_411 (O_411,N_2943,N_2982);
nor UO_412 (O_412,N_2936,N_2997);
nand UO_413 (O_413,N_2954,N_2952);
or UO_414 (O_414,N_2997,N_2949);
or UO_415 (O_415,N_2959,N_2966);
and UO_416 (O_416,N_2939,N_2989);
nor UO_417 (O_417,N_2945,N_2967);
or UO_418 (O_418,N_2940,N_2979);
nand UO_419 (O_419,N_2994,N_2939);
or UO_420 (O_420,N_2927,N_2995);
or UO_421 (O_421,N_2991,N_2934);
nor UO_422 (O_422,N_2975,N_2968);
nand UO_423 (O_423,N_2992,N_2982);
or UO_424 (O_424,N_2948,N_2931);
or UO_425 (O_425,N_2970,N_2973);
nand UO_426 (O_426,N_2964,N_2970);
nor UO_427 (O_427,N_2965,N_2931);
or UO_428 (O_428,N_2970,N_2966);
or UO_429 (O_429,N_2958,N_2960);
nand UO_430 (O_430,N_2964,N_2995);
nand UO_431 (O_431,N_2949,N_2981);
nor UO_432 (O_432,N_2933,N_2970);
nand UO_433 (O_433,N_2987,N_2948);
and UO_434 (O_434,N_2967,N_2989);
or UO_435 (O_435,N_2947,N_2955);
nor UO_436 (O_436,N_2972,N_2944);
and UO_437 (O_437,N_2948,N_2940);
nand UO_438 (O_438,N_2969,N_2932);
and UO_439 (O_439,N_2976,N_2963);
nor UO_440 (O_440,N_2928,N_2976);
nand UO_441 (O_441,N_2946,N_2993);
and UO_442 (O_442,N_2982,N_2953);
nand UO_443 (O_443,N_2941,N_2998);
nand UO_444 (O_444,N_2947,N_2969);
nor UO_445 (O_445,N_2952,N_2950);
and UO_446 (O_446,N_2991,N_2956);
and UO_447 (O_447,N_2972,N_2960);
and UO_448 (O_448,N_2969,N_2970);
or UO_449 (O_449,N_2991,N_2971);
nand UO_450 (O_450,N_2993,N_2960);
nand UO_451 (O_451,N_2934,N_2953);
xnor UO_452 (O_452,N_2965,N_2978);
nor UO_453 (O_453,N_2926,N_2974);
nor UO_454 (O_454,N_2964,N_2943);
nand UO_455 (O_455,N_2937,N_2950);
and UO_456 (O_456,N_2960,N_2987);
or UO_457 (O_457,N_2961,N_2977);
nor UO_458 (O_458,N_2944,N_2960);
nor UO_459 (O_459,N_2967,N_2944);
nor UO_460 (O_460,N_2937,N_2974);
nand UO_461 (O_461,N_2977,N_2995);
and UO_462 (O_462,N_2997,N_2968);
and UO_463 (O_463,N_2994,N_2978);
and UO_464 (O_464,N_2930,N_2994);
nand UO_465 (O_465,N_2946,N_2977);
or UO_466 (O_466,N_2948,N_2926);
nor UO_467 (O_467,N_2926,N_2935);
nand UO_468 (O_468,N_2962,N_2998);
nand UO_469 (O_469,N_2933,N_2962);
nand UO_470 (O_470,N_2936,N_2951);
nand UO_471 (O_471,N_2986,N_2964);
nand UO_472 (O_472,N_2953,N_2951);
and UO_473 (O_473,N_2954,N_2997);
and UO_474 (O_474,N_2969,N_2962);
and UO_475 (O_475,N_2947,N_2941);
and UO_476 (O_476,N_2975,N_2944);
nor UO_477 (O_477,N_2963,N_2959);
nand UO_478 (O_478,N_2985,N_2979);
or UO_479 (O_479,N_2944,N_2985);
nor UO_480 (O_480,N_2946,N_2982);
or UO_481 (O_481,N_2941,N_2962);
or UO_482 (O_482,N_2993,N_2988);
or UO_483 (O_483,N_2984,N_2985);
nand UO_484 (O_484,N_2984,N_2946);
and UO_485 (O_485,N_2964,N_2994);
nand UO_486 (O_486,N_2982,N_2958);
and UO_487 (O_487,N_2979,N_2946);
or UO_488 (O_488,N_2953,N_2950);
and UO_489 (O_489,N_2964,N_2967);
and UO_490 (O_490,N_2978,N_2934);
nand UO_491 (O_491,N_2968,N_2958);
nor UO_492 (O_492,N_2955,N_2989);
nor UO_493 (O_493,N_2962,N_2979);
nor UO_494 (O_494,N_2977,N_2942);
and UO_495 (O_495,N_2993,N_2998);
nor UO_496 (O_496,N_2945,N_2966);
nor UO_497 (O_497,N_2997,N_2944);
and UO_498 (O_498,N_2935,N_2933);
or UO_499 (O_499,N_2996,N_2942);
endmodule