module basic_2500_25000_3000_125_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_564,In_1798);
and U1 (N_1,In_695,In_1081);
nand U2 (N_2,In_2013,In_878);
or U3 (N_3,In_1186,In_773);
and U4 (N_4,In_1549,In_120);
or U5 (N_5,In_1028,In_1618);
nor U6 (N_6,In_156,In_2475);
nand U7 (N_7,In_916,In_568);
or U8 (N_8,In_930,In_913);
nor U9 (N_9,In_1574,In_2189);
or U10 (N_10,In_914,In_1035);
nor U11 (N_11,In_789,In_2210);
nor U12 (N_12,In_2197,In_1361);
and U13 (N_13,In_1251,In_111);
xor U14 (N_14,In_881,In_260);
and U15 (N_15,In_418,In_809);
or U16 (N_16,In_787,In_1247);
or U17 (N_17,In_977,In_1522);
nor U18 (N_18,In_2206,In_35);
xnor U19 (N_19,In_1814,In_2236);
nand U20 (N_20,In_915,In_968);
and U21 (N_21,In_1052,In_850);
or U22 (N_22,In_305,In_1875);
nand U23 (N_23,In_1387,In_1780);
or U24 (N_24,In_1929,In_1625);
nand U25 (N_25,In_1627,In_1486);
and U26 (N_26,In_2134,In_2286);
and U27 (N_27,In_551,In_59);
and U28 (N_28,In_1356,In_338);
nor U29 (N_29,In_1435,In_2415);
nor U30 (N_30,In_99,In_836);
nor U31 (N_31,In_2014,In_872);
and U32 (N_32,In_1739,In_941);
nor U33 (N_33,In_1912,In_1523);
and U34 (N_34,In_2117,In_750);
nand U35 (N_35,In_609,In_2338);
nand U36 (N_36,In_664,In_1734);
nor U37 (N_37,In_2141,In_166);
nor U38 (N_38,In_1143,In_229);
nor U39 (N_39,In_2179,In_553);
nor U40 (N_40,In_1520,In_1181);
and U41 (N_41,In_535,In_1413);
nor U42 (N_42,In_1153,In_848);
and U43 (N_43,In_2455,In_962);
nand U44 (N_44,In_756,In_586);
or U45 (N_45,In_826,In_2221);
nand U46 (N_46,In_2322,In_1973);
nand U47 (N_47,In_782,In_1423);
nand U48 (N_48,In_1350,In_455);
or U49 (N_49,In_1114,In_1958);
nor U50 (N_50,In_323,In_693);
nor U51 (N_51,In_1258,In_33);
nor U52 (N_52,In_1490,In_170);
xor U53 (N_53,In_735,In_1284);
nand U54 (N_54,In_581,In_1243);
xor U55 (N_55,In_1190,In_28);
and U56 (N_56,In_2068,In_1675);
nand U57 (N_57,In_2484,In_2156);
nor U58 (N_58,In_784,In_1868);
nand U59 (N_59,In_255,In_67);
and U60 (N_60,In_998,In_2409);
and U61 (N_61,In_1926,In_433);
or U62 (N_62,In_722,In_2490);
or U63 (N_63,In_833,In_1833);
nor U64 (N_64,In_747,In_20);
or U65 (N_65,In_1691,In_1891);
and U66 (N_66,In_2103,In_272);
nand U67 (N_67,In_819,In_421);
and U68 (N_68,In_2074,In_791);
nor U69 (N_69,In_311,In_1678);
nand U70 (N_70,In_1959,In_282);
and U71 (N_71,In_2102,In_2171);
nor U72 (N_72,In_736,In_905);
and U73 (N_73,In_52,In_2241);
or U74 (N_74,In_2356,In_1381);
and U75 (N_75,In_1561,In_1591);
nor U76 (N_76,In_1744,In_65);
and U77 (N_77,In_2298,In_1826);
or U78 (N_78,In_1098,In_1882);
nand U79 (N_79,In_44,In_801);
and U80 (N_80,In_1424,In_2281);
nor U81 (N_81,In_2265,In_241);
or U82 (N_82,In_2367,In_292);
nor U83 (N_83,In_1097,In_2317);
or U84 (N_84,In_101,In_1550);
nor U85 (N_85,In_1472,In_1519);
nand U86 (N_86,In_712,In_741);
nand U87 (N_87,In_1645,In_1278);
nand U88 (N_88,In_774,In_2418);
nand U89 (N_89,In_2294,In_273);
nor U90 (N_90,In_1048,In_1215);
nand U91 (N_91,In_2349,In_749);
nand U92 (N_92,In_96,In_1341);
or U93 (N_93,In_2406,In_1211);
and U94 (N_94,In_638,In_1418);
or U95 (N_95,In_2440,In_1007);
xor U96 (N_96,In_249,In_1398);
or U97 (N_97,In_512,In_2231);
xnor U98 (N_98,In_2174,In_838);
or U99 (N_99,In_1493,In_1183);
and U100 (N_100,In_871,In_1610);
xnor U101 (N_101,In_2465,In_1126);
or U102 (N_102,In_1693,In_757);
and U103 (N_103,In_1012,In_810);
or U104 (N_104,In_1534,In_1303);
nor U105 (N_105,In_428,In_907);
nor U106 (N_106,In_1036,In_1282);
xnor U107 (N_107,In_1803,In_135);
or U108 (N_108,In_1664,In_999);
or U109 (N_109,In_1317,In_1174);
or U110 (N_110,In_640,In_1207);
or U111 (N_111,In_492,In_2434);
and U112 (N_112,In_371,In_1927);
and U113 (N_113,In_381,In_1784);
nor U114 (N_114,In_87,In_1400);
nor U115 (N_115,In_394,In_2421);
and U116 (N_116,In_714,In_1680);
nand U117 (N_117,In_1677,In_1853);
or U118 (N_118,In_1804,In_2203);
nor U119 (N_119,In_2385,In_958);
or U120 (N_120,In_1852,In_2373);
nor U121 (N_121,In_146,In_694);
xnor U122 (N_122,In_2289,In_1899);
and U123 (N_123,In_1898,In_2035);
nand U124 (N_124,In_1871,In_2175);
nand U125 (N_125,In_1507,In_676);
and U126 (N_126,In_100,In_1313);
nor U127 (N_127,In_301,In_1351);
nand U128 (N_128,In_1330,In_1306);
and U129 (N_129,In_2497,In_1681);
nor U130 (N_130,In_488,In_672);
and U131 (N_131,In_1011,In_1223);
or U132 (N_132,In_713,In_729);
or U133 (N_133,In_1893,In_1735);
nor U134 (N_134,In_115,In_1033);
or U135 (N_135,In_312,In_364);
and U136 (N_136,In_2127,In_274);
xnor U137 (N_137,In_1944,In_1983);
nand U138 (N_138,In_2052,In_2444);
nor U139 (N_139,In_2138,In_554);
or U140 (N_140,In_2381,In_1514);
or U141 (N_141,In_895,In_1483);
and U142 (N_142,In_2323,In_119);
nand U143 (N_143,In_45,In_608);
nand U144 (N_144,In_1428,In_1935);
and U145 (N_145,In_1373,In_327);
nand U146 (N_146,In_2291,In_1121);
and U147 (N_147,In_1308,In_2296);
and U148 (N_148,In_1980,In_781);
or U149 (N_149,In_330,In_767);
nand U150 (N_150,In_2047,In_1179);
and U151 (N_151,In_875,In_1296);
nand U152 (N_152,In_877,In_469);
nor U153 (N_153,In_588,In_725);
nand U154 (N_154,In_1042,In_2345);
nand U155 (N_155,In_2084,In_324);
or U156 (N_156,In_1000,In_1032);
and U157 (N_157,In_1575,In_1106);
xnor U158 (N_158,In_2195,In_1198);
or U159 (N_159,In_2049,In_1619);
nand U160 (N_160,In_1799,In_1951);
nor U161 (N_161,In_1995,In_1056);
and U162 (N_162,In_1392,In_2330);
xnor U163 (N_163,In_2372,In_1182);
and U164 (N_164,In_370,In_1405);
and U165 (N_165,In_2387,In_1706);
and U166 (N_166,In_75,In_755);
nor U167 (N_167,In_1123,In_1641);
and U168 (N_168,In_46,In_1782);
nor U169 (N_169,In_1811,In_1116);
nor U170 (N_170,In_1792,In_1046);
nand U171 (N_171,In_2267,In_1682);
and U172 (N_172,In_1332,In_963);
or U173 (N_173,In_2321,In_365);
nand U174 (N_174,In_1425,In_1727);
and U175 (N_175,In_546,In_443);
or U176 (N_176,In_1616,In_812);
xor U177 (N_177,In_1414,In_1378);
nand U178 (N_178,In_2213,In_2314);
nand U179 (N_179,In_2392,In_1656);
or U180 (N_180,In_1185,In_448);
and U181 (N_181,In_949,In_1805);
nor U182 (N_182,In_254,In_1749);
xnor U183 (N_183,In_172,In_1438);
or U184 (N_184,In_199,In_299);
nor U185 (N_185,In_577,In_1458);
or U186 (N_186,In_29,In_2097);
or U187 (N_187,In_2253,In_2266);
nor U188 (N_188,In_211,In_979);
xor U189 (N_189,In_110,In_2250);
nor U190 (N_190,In_1325,In_1745);
nand U191 (N_191,In_1846,In_1991);
or U192 (N_192,In_1269,In_390);
and U193 (N_193,In_2159,In_1346);
nor U194 (N_194,In_181,In_1091);
and U195 (N_195,In_1817,In_2028);
nand U196 (N_196,In_1216,In_527);
nand U197 (N_197,In_2079,In_2319);
and U198 (N_198,In_66,In_2350);
nor U199 (N_199,In_574,In_2009);
and U200 (N_200,In_495,In_2464);
and U201 (N_201,N_38,In_355);
or U202 (N_202,In_372,In_815);
nand U203 (N_203,In_206,In_1037);
or U204 (N_204,In_298,In_2332);
or U205 (N_205,In_710,In_912);
nand U206 (N_206,In_1924,In_345);
or U207 (N_207,In_195,In_2478);
or U208 (N_208,N_17,N_109);
and U209 (N_209,In_1698,In_1642);
nand U210 (N_210,In_1823,In_1213);
nand U211 (N_211,In_1460,In_131);
nand U212 (N_212,In_1650,In_674);
nor U213 (N_213,In_858,In_707);
or U214 (N_214,In_408,In_558);
and U215 (N_215,In_662,In_1430);
and U216 (N_216,In_653,In_1020);
and U217 (N_217,N_48,In_1595);
or U218 (N_218,In_1915,In_1570);
xnor U219 (N_219,N_89,In_16);
or U220 (N_220,N_44,In_547);
nor U221 (N_221,In_1477,In_2207);
xnor U222 (N_222,In_1933,In_700);
nor U223 (N_223,In_1071,In_2278);
or U224 (N_224,In_1367,In_532);
nand U225 (N_225,In_1402,In_2149);
or U226 (N_226,In_2087,In_1674);
nor U227 (N_227,In_171,N_148);
xor U228 (N_228,N_40,In_2311);
xor U229 (N_229,In_2243,In_366);
xnor U230 (N_230,In_1250,In_1286);
nor U231 (N_231,In_920,In_83);
xor U232 (N_232,In_552,In_2441);
and U233 (N_233,In_13,In_891);
or U234 (N_234,In_412,In_149);
nor U235 (N_235,In_2034,In_168);
nor U236 (N_236,In_490,In_2493);
nor U237 (N_237,In_9,In_1118);
and U238 (N_238,In_1231,In_927);
or U239 (N_239,In_541,In_1928);
and U240 (N_240,In_788,In_1562);
nor U241 (N_241,In_1975,In_884);
nor U242 (N_242,In_615,In_944);
nand U243 (N_243,In_1343,In_1352);
nand U244 (N_244,In_2402,In_2026);
nand U245 (N_245,In_1119,In_427);
xor U246 (N_246,In_1253,In_1128);
nor U247 (N_247,In_1669,N_167);
xor U248 (N_248,In_1446,N_19);
and U249 (N_249,In_1305,In_1019);
nor U250 (N_250,In_491,In_1781);
nor U251 (N_251,In_2164,In_2438);
nor U252 (N_252,In_2058,In_1828);
nor U253 (N_253,In_486,In_1512);
nand U254 (N_254,In_2252,In_2196);
or U255 (N_255,In_1726,In_2461);
nand U256 (N_256,In_1827,In_1429);
and U257 (N_257,In_106,N_74);
and U258 (N_258,In_1327,In_514);
nor U259 (N_259,In_2310,In_1531);
nand U260 (N_260,In_150,In_2437);
or U261 (N_261,In_2398,In_1360);
or U262 (N_262,In_477,N_165);
nand U263 (N_263,In_441,In_1696);
nor U264 (N_264,In_1450,In_1757);
nor U265 (N_265,In_1968,In_1785);
nor U266 (N_266,In_1015,In_824);
nor U267 (N_267,In_1221,In_1416);
nand U268 (N_268,In_2326,In_1358);
nor U269 (N_269,In_606,In_887);
or U270 (N_270,In_972,In_31);
and U271 (N_271,In_1851,In_1647);
or U272 (N_272,In_1344,In_1203);
and U273 (N_273,In_1265,In_1812);
xor U274 (N_274,In_2116,In_1025);
and U275 (N_275,In_198,In_1601);
or U276 (N_276,In_2090,In_2325);
and U277 (N_277,In_737,In_721);
or U278 (N_278,In_854,In_1314);
nand U279 (N_279,In_2128,In_2276);
nor U280 (N_280,In_1887,In_221);
and U281 (N_281,N_114,In_2254);
nor U282 (N_282,In_1234,In_1171);
nor U283 (N_283,In_2124,N_59);
and U284 (N_284,In_1932,In_2366);
xnor U285 (N_285,In_480,In_656);
and U286 (N_286,In_2401,In_616);
or U287 (N_287,N_95,N_9);
xnor U288 (N_288,In_169,In_2318);
or U289 (N_289,N_105,N_55);
nand U290 (N_290,In_349,In_2268);
nor U291 (N_291,In_1136,N_129);
and U292 (N_292,In_496,In_1431);
or U293 (N_293,In_2163,In_2428);
nor U294 (N_294,In_417,In_988);
nor U295 (N_295,In_2045,In_1130);
nand U296 (N_296,N_18,In_1956);
nor U297 (N_297,In_2077,N_1);
nor U298 (N_298,In_1504,N_132);
nand U299 (N_299,In_1553,In_752);
nor U300 (N_300,In_560,N_140);
nand U301 (N_301,In_405,In_1248);
or U302 (N_302,In_1612,In_2186);
or U303 (N_303,In_2146,In_2063);
or U304 (N_304,In_2153,In_2172);
or U305 (N_305,N_36,In_1333);
or U306 (N_306,In_1878,In_250);
nand U307 (N_307,In_2292,In_2282);
nor U308 (N_308,In_127,In_1637);
nor U309 (N_309,In_51,N_96);
nor U310 (N_310,In_23,In_689);
nand U311 (N_311,In_1235,In_1661);
and U312 (N_312,In_458,In_2046);
nor U313 (N_313,In_1527,In_1233);
nand U314 (N_314,In_2379,In_2155);
and U315 (N_315,In_1320,In_1560);
nand U316 (N_316,In_2358,N_158);
xor U317 (N_317,N_107,In_2498);
nor U318 (N_318,In_359,In_1873);
and U319 (N_319,In_1178,In_1173);
and U320 (N_320,In_1487,In_699);
xor U321 (N_321,In_2051,In_219);
nand U322 (N_322,In_1892,In_1663);
xor U323 (N_323,In_898,In_439);
or U324 (N_324,In_1009,In_476);
xor U325 (N_325,In_649,In_1708);
and U326 (N_326,In_524,N_72);
or U327 (N_327,In_504,In_526);
nor U328 (N_328,In_2093,In_1082);
nor U329 (N_329,In_2202,In_1822);
nand U330 (N_330,N_3,In_284);
nor U331 (N_331,In_683,In_1273);
nand U332 (N_332,In_573,In_2088);
or U333 (N_333,In_122,In_2222);
xor U334 (N_334,In_430,In_484);
and U335 (N_335,In_1068,In_1261);
or U336 (N_336,In_1966,N_197);
nor U337 (N_337,In_1748,In_503);
and U338 (N_338,In_77,In_1196);
or U339 (N_339,In_982,In_1163);
and U340 (N_340,N_71,In_2450);
nor U341 (N_341,In_230,In_317);
and U342 (N_342,In_378,In_1908);
nor U343 (N_343,In_460,In_1703);
and U344 (N_344,In_399,In_698);
nand U345 (N_345,In_1339,In_2369);
and U346 (N_346,In_465,In_2473);
nand U347 (N_347,In_2126,In_2426);
or U348 (N_348,In_1232,In_57);
and U349 (N_349,In_1224,In_436);
and U350 (N_350,In_933,In_187);
xnor U351 (N_351,In_1676,In_1403);
nor U352 (N_352,In_684,In_2239);
or U353 (N_353,In_572,In_522);
xor U354 (N_354,N_182,In_2148);
nor U355 (N_355,N_113,In_1724);
nor U356 (N_356,In_2200,In_776);
or U357 (N_357,In_207,In_2157);
and U358 (N_358,In_1302,In_1768);
nor U359 (N_359,In_2335,N_161);
nor U360 (N_360,In_2468,In_2371);
nor U361 (N_361,In_1571,In_598);
and U362 (N_362,In_1087,In_1750);
and U363 (N_363,In_1260,In_1517);
nand U364 (N_364,In_1292,In_2447);
nor U365 (N_365,In_2111,In_2359);
nor U366 (N_366,In_2181,In_1086);
nand U367 (N_367,In_61,In_911);
nor U368 (N_368,In_1689,In_1088);
and U369 (N_369,In_706,In_1996);
nor U370 (N_370,In_1964,In_2225);
or U371 (N_371,In_1095,In_1484);
or U372 (N_372,In_1267,In_1443);
nor U373 (N_373,In_2023,N_145);
or U374 (N_374,In_540,In_63);
or U375 (N_375,In_438,In_1532);
or U376 (N_376,In_1509,In_668);
or U377 (N_377,In_873,In_594);
nand U378 (N_378,N_97,In_2333);
nand U379 (N_379,In_582,In_1903);
nand U380 (N_380,In_825,N_42);
nand U381 (N_381,In_191,In_852);
and U382 (N_382,In_2050,In_1600);
xnor U383 (N_383,In_1976,In_406);
or U384 (N_384,In_1860,In_401);
or U385 (N_385,In_136,In_1329);
or U386 (N_386,In_1242,In_533);
or U387 (N_387,In_2378,In_2405);
or U388 (N_388,In_2086,In_2137);
or U389 (N_389,In_2062,In_2214);
xnor U390 (N_390,In_158,In_1658);
and U391 (N_391,In_1971,In_629);
nor U392 (N_392,In_2144,In_1201);
nand U393 (N_393,In_143,In_965);
and U394 (N_394,In_1038,In_74);
and U395 (N_395,In_233,In_992);
or U396 (N_396,In_1335,N_88);
nand U397 (N_397,In_1047,In_682);
nor U398 (N_398,In_658,In_280);
and U399 (N_399,In_753,In_1856);
nand U400 (N_400,In_2001,In_217);
and U401 (N_401,In_325,In_1107);
and U402 (N_402,In_1907,In_1217);
nand U403 (N_403,In_2451,In_1140);
and U404 (N_404,In_380,In_2389);
or U405 (N_405,In_1918,In_426);
nand U406 (N_406,In_623,In_2482);
and U407 (N_407,In_2071,In_543);
xnor U408 (N_408,In_917,In_1752);
and U409 (N_409,N_275,In_1569);
nand U410 (N_410,In_637,In_1440);
nor U411 (N_411,In_1919,N_386);
nand U412 (N_412,N_366,In_1659);
or U413 (N_413,In_1690,In_1717);
nor U414 (N_414,In_1800,In_925);
or U415 (N_415,In_1219,In_1420);
or U416 (N_416,In_1455,In_415);
nor U417 (N_417,In_373,In_1169);
nor U418 (N_418,In_626,In_1065);
and U419 (N_419,In_1679,In_2257);
and U420 (N_420,In_986,In_634);
nand U421 (N_421,In_2070,In_1589);
and U422 (N_422,In_2168,In_1218);
nand U423 (N_423,In_657,In_377);
xnor U424 (N_424,In_1204,In_152);
nor U425 (N_425,In_614,In_2040);
nor U426 (N_426,In_579,In_1779);
nor U427 (N_427,In_2057,In_353);
xor U428 (N_428,N_163,In_1010);
or U429 (N_429,In_1461,In_876);
nand U430 (N_430,In_1124,N_350);
nand U431 (N_431,In_2106,In_1939);
nand U432 (N_432,In_1567,In_1528);
nor U433 (N_433,In_2205,In_315);
and U434 (N_434,In_2476,In_1085);
xnor U435 (N_435,In_271,In_245);
nand U436 (N_436,N_0,In_341);
nor U437 (N_437,In_1579,In_1810);
nand U438 (N_438,In_2274,In_2204);
nand U439 (N_439,In_49,N_184);
nand U440 (N_440,In_1175,In_563);
or U441 (N_441,N_229,In_2185);
and U442 (N_442,In_402,In_2365);
nand U443 (N_443,In_73,In_1241);
nand U444 (N_444,In_2386,In_1298);
nand U445 (N_445,In_1023,In_334);
nor U446 (N_446,In_1945,In_1386);
and U447 (N_447,In_1767,N_273);
or U448 (N_448,In_1747,In_1322);
nand U449 (N_449,In_818,In_1214);
xnor U450 (N_450,N_378,In_516);
or U451 (N_451,In_2279,In_942);
nor U452 (N_452,In_599,In_310);
nand U453 (N_453,In_497,In_1411);
and U454 (N_454,N_336,In_2199);
or U455 (N_455,N_178,N_4);
nor U456 (N_456,In_314,N_360);
nand U457 (N_457,In_1969,In_845);
or U458 (N_458,In_1195,N_106);
nor U459 (N_459,In_1093,In_1603);
xor U460 (N_460,In_601,In_523);
or U461 (N_461,In_1067,In_981);
nand U462 (N_462,In_456,In_1276);
nor U463 (N_463,In_1469,In_2232);
nand U464 (N_464,In_1901,N_198);
nor U465 (N_465,In_995,In_1790);
nor U466 (N_466,In_1938,In_2457);
nor U467 (N_467,In_762,In_587);
and U468 (N_468,In_2011,In_1287);
nor U469 (N_469,In_388,In_1772);
and U470 (N_470,In_1736,N_238);
and U471 (N_471,In_1245,In_2076);
nor U472 (N_472,In_994,In_398);
nand U473 (N_473,In_1646,In_2099);
and U474 (N_474,In_155,N_194);
nand U475 (N_475,In_3,N_204);
nand U476 (N_476,In_795,N_177);
nor U477 (N_477,In_2108,N_31);
nor U478 (N_478,N_223,In_94);
nor U479 (N_479,In_566,In_1866);
xor U480 (N_480,In_660,In_1159);
and U481 (N_481,In_2165,In_639);
nor U482 (N_482,In_2041,In_1501);
nand U483 (N_483,N_252,N_85);
or U484 (N_484,In_2258,In_1883);
nand U485 (N_485,In_1089,In_1342);
or U486 (N_486,In_648,In_536);
nand U487 (N_487,In_1793,In_288);
nor U488 (N_488,In_95,In_244);
nand U489 (N_489,N_314,In_1725);
or U490 (N_490,In_1474,In_2091);
nand U491 (N_491,In_1709,In_98);
or U492 (N_492,N_24,In_1884);
nor U493 (N_493,In_655,In_337);
and U494 (N_494,In_368,In_403);
nand U495 (N_495,N_14,In_1756);
nand U496 (N_496,In_1092,In_1388);
or U497 (N_497,In_548,In_620);
xnor U498 (N_498,N_187,In_1791);
nand U499 (N_499,In_1459,In_759);
nor U500 (N_500,N_201,N_255);
and U501 (N_501,In_192,In_2064);
nand U502 (N_502,N_290,In_2242);
nor U503 (N_503,N_142,In_1340);
nand U504 (N_504,In_636,N_231);
or U505 (N_505,In_1577,In_996);
or U506 (N_506,In_1842,In_1626);
or U507 (N_507,N_311,In_2024);
and U508 (N_508,In_1802,N_69);
and U509 (N_509,In_1176,In_1321);
nand U510 (N_510,In_295,In_1497);
nand U511 (N_511,In_709,In_2218);
nand U512 (N_512,In_1862,In_1597);
or U513 (N_513,In_1004,In_190);
and U514 (N_514,In_1777,In_1002);
nand U515 (N_515,In_1746,In_1017);
nand U516 (N_516,In_724,In_1239);
nand U517 (N_517,In_1134,In_242);
or U518 (N_518,In_1132,In_1809);
nor U519 (N_519,In_2347,In_643);
nand U520 (N_520,In_1054,N_398);
xor U521 (N_521,In_1205,In_1513);
nor U522 (N_522,In_1156,In_2443);
or U523 (N_523,In_1835,In_137);
or U524 (N_524,In_2037,In_1816);
or U525 (N_525,In_517,In_356);
or U526 (N_526,In_437,In_903);
nor U527 (N_527,In_124,In_2439);
or U528 (N_528,In_866,In_163);
nor U529 (N_529,In_1877,N_175);
or U530 (N_530,In_1536,In_1266);
and U531 (N_531,In_1890,In_118);
nor U532 (N_532,In_1077,In_1640);
or U533 (N_533,N_137,In_926);
nand U534 (N_534,In_993,In_1848);
and U535 (N_535,In_772,In_1129);
or U536 (N_536,N_128,N_315);
nor U537 (N_537,In_1869,In_1967);
nor U538 (N_538,N_369,N_112);
nor U539 (N_539,In_2092,N_306);
nor U540 (N_540,In_126,N_349);
or U541 (N_541,In_1789,In_717);
nand U542 (N_542,In_1471,N_219);
nor U543 (N_543,In_2096,N_32);
and U544 (N_544,In_162,In_585);
and U545 (N_545,In_175,N_359);
and U546 (N_546,In_2491,N_218);
and U547 (N_547,In_2480,N_318);
nor U548 (N_548,In_1886,In_1328);
and U549 (N_549,In_2247,In_2104);
nor U550 (N_550,In_2417,N_217);
nand U551 (N_551,In_842,In_277);
or U552 (N_552,N_248,In_2269);
xnor U553 (N_553,In_1808,In_397);
and U554 (N_554,In_565,In_1863);
and U555 (N_555,In_204,N_171);
nor U556 (N_556,In_53,In_1565);
and U557 (N_557,In_68,In_1324);
nand U558 (N_558,In_1993,In_1593);
nand U559 (N_559,N_246,In_1421);
xnor U560 (N_560,In_2160,In_2320);
nand U561 (N_561,In_2255,In_893);
nor U562 (N_562,In_2223,In_470);
and U563 (N_563,In_2069,In_1319);
and U564 (N_564,In_2259,In_830);
nor U565 (N_565,In_287,In_76);
or U566 (N_566,N_141,In_602);
nand U567 (N_567,In_1475,N_381);
and U568 (N_568,In_343,In_1518);
nand U569 (N_569,In_2492,N_286);
nand U570 (N_570,In_1539,In_2256);
nand U571 (N_571,In_1547,In_1917);
nor U572 (N_572,In_2031,In_1788);
and U573 (N_573,In_921,In_1987);
nand U574 (N_574,In_596,In_1448);
or U575 (N_575,In_331,In_2394);
nor U576 (N_576,In_1075,In_975);
nand U577 (N_577,In_1662,In_2008);
nand U578 (N_578,In_748,In_1466);
or U579 (N_579,In_2288,In_159);
nand U580 (N_580,In_117,In_1230);
and U581 (N_581,In_1151,In_1096);
or U582 (N_582,In_1249,In_745);
and U583 (N_583,In_2382,In_870);
or U584 (N_584,N_155,In_1556);
nor U585 (N_585,In_1187,In_2328);
nand U586 (N_586,In_400,In_633);
or U587 (N_587,In_589,In_243);
or U588 (N_588,In_1997,In_419);
or U589 (N_589,In_2183,N_157);
nor U590 (N_590,In_1285,In_1657);
nor U591 (N_591,In_945,In_1079);
and U592 (N_592,In_2169,In_2147);
nand U593 (N_593,In_97,In_1592);
or U594 (N_594,In_1110,In_1016);
and U595 (N_595,In_860,In_807);
nor U596 (N_596,N_309,In_2101);
and U597 (N_597,In_1112,In_1741);
and U598 (N_598,In_1080,In_2234);
nand U599 (N_599,In_2121,In_1738);
or U600 (N_600,In_2229,In_392);
nand U601 (N_601,In_1061,In_1730);
nand U602 (N_602,In_2215,In_1439);
and U603 (N_603,N_70,In_2130);
and U604 (N_604,In_720,N_338);
or U605 (N_605,N_509,N_295);
or U606 (N_606,In_1410,N_445);
and U607 (N_607,N_83,In_2460);
nor U608 (N_608,In_1936,N_244);
nand U609 (N_609,In_1001,In_846);
or U610 (N_610,In_2361,N_450);
nand U611 (N_611,In_1632,In_1);
or U612 (N_612,N_63,N_25);
nand U613 (N_613,In_743,N_599);
nand U614 (N_614,In_2273,In_1353);
nand U615 (N_615,In_2302,In_2030);
nor U616 (N_616,In_584,In_145);
or U617 (N_617,In_1281,In_1422);
and U618 (N_618,N_515,In_2400);
and U619 (N_619,In_296,In_978);
nand U620 (N_620,In_1499,In_1700);
nand U621 (N_621,In_1986,In_2143);
and U622 (N_622,In_1395,In_1832);
and U623 (N_623,N_162,In_1259);
and U624 (N_624,In_141,N_412);
nand U625 (N_625,In_487,N_181);
nand U626 (N_626,In_1761,In_1737);
nor U627 (N_627,In_2033,In_294);
or U628 (N_628,In_519,In_1858);
and U629 (N_629,In_591,N_341);
or U630 (N_630,In_2238,In_1713);
and U631 (N_631,In_1583,N_335);
nor U632 (N_632,N_473,In_93);
or U633 (N_633,In_42,N_160);
or U634 (N_634,In_1844,N_514);
nor U635 (N_635,N_512,In_2495);
nand U636 (N_636,N_472,In_1865);
xnor U637 (N_637,In_1540,In_723);
or U638 (N_638,In_799,In_1376);
nor U639 (N_639,In_329,N_371);
and U640 (N_640,In_701,In_1120);
nand U641 (N_641,In_1309,N_356);
and U642 (N_642,In_113,In_1758);
and U643 (N_643,In_1293,In_733);
nor U644 (N_644,N_584,In_286);
and U645 (N_645,N_54,N_94);
nor U646 (N_646,N_153,In_622);
or U647 (N_647,N_591,In_1467);
and U648 (N_648,In_468,In_1371);
and U649 (N_649,In_928,In_2065);
nor U650 (N_650,In_531,In_1896);
xnor U651 (N_651,In_805,N_481);
nor U652 (N_652,In_2308,In_1359);
xnor U653 (N_653,In_708,In_410);
and U654 (N_654,N_556,In_2414);
nor U655 (N_655,In_798,In_1288);
nand U656 (N_656,N_419,In_220);
or U657 (N_657,In_1554,N_324);
nand U658 (N_658,In_950,In_974);
nor U659 (N_659,N_5,In_1576);
nand U660 (N_660,In_2227,N_496);
nand U661 (N_661,In_1906,In_461);
nor U662 (N_662,In_2006,In_1797);
nor U663 (N_663,In_1776,In_2140);
or U664 (N_664,N_285,N_365);
or U665 (N_665,In_1825,In_971);
nand U666 (N_666,N_457,In_562);
nor U667 (N_667,In_2125,In_2301);
or U668 (N_668,In_256,N_351);
and U669 (N_669,N_276,In_2413);
or U670 (N_670,N_299,N_483);
or U671 (N_671,In_2081,In_1541);
nor U672 (N_672,N_494,In_768);
nand U673 (N_673,In_1312,In_1733);
nor U674 (N_674,In_1974,N_189);
nand U675 (N_675,In_955,In_213);
or U676 (N_676,N_269,In_1502);
or U677 (N_677,In_1463,N_352);
and U678 (N_678,N_587,N_122);
xnor U679 (N_679,N_47,N_256);
and U680 (N_680,In_1003,In_1401);
or U681 (N_681,N_277,N_393);
and U682 (N_682,In_414,In_1948);
or U683 (N_683,In_2061,In_2262);
nand U684 (N_684,In_600,In_1099);
nor U685 (N_685,N_21,N_405);
nand U686 (N_686,In_1818,In_12);
nor U687 (N_687,In_1602,In_983);
nor U688 (N_688,In_1113,In_240);
nand U689 (N_689,In_2025,In_1783);
or U690 (N_690,In_1697,In_138);
nor U691 (N_691,In_2448,In_1962);
xnor U692 (N_692,In_922,N_588);
nand U693 (N_693,In_1586,In_530);
nand U694 (N_694,In_1949,In_1209);
or U695 (N_695,In_2383,In_1578);
or U696 (N_696,In_493,In_964);
nand U697 (N_697,In_2453,N_247);
nor U698 (N_698,In_1109,N_531);
xnor U699 (N_699,In_1755,In_1133);
nor U700 (N_700,N_569,In_246);
nand U701 (N_701,In_1914,In_1839);
or U702 (N_702,In_81,In_1615);
nor U703 (N_703,N_168,In_2340);
nand U704 (N_704,In_556,In_1830);
nand U705 (N_705,In_800,In_164);
or U706 (N_706,In_62,In_2483);
and U707 (N_707,In_114,In_1348);
or U708 (N_708,In_447,In_597);
nand U709 (N_709,In_1447,In_2284);
nand U710 (N_710,N_239,In_952);
or U711 (N_711,N_353,N_533);
and U712 (N_712,In_2407,In_1854);
xnor U713 (N_713,N_169,In_1950);
and U714 (N_714,In_1742,In_2173);
or U715 (N_715,In_2339,In_862);
or U716 (N_716,N_497,N_53);
or U717 (N_717,In_247,In_340);
and U718 (N_718,In_103,In_511);
or U719 (N_719,In_796,In_1686);
and U720 (N_720,In_104,In_885);
or U721 (N_721,In_2188,In_1062);
nor U722 (N_722,In_1670,In_1139);
or U723 (N_723,N_478,In_128);
nor U724 (N_724,In_1608,N_41);
or U725 (N_725,N_75,In_1694);
and U726 (N_726,In_1526,N_504);
nor U727 (N_727,In_901,In_37);
or U728 (N_728,In_1942,In_223);
or U729 (N_729,N_519,In_2219);
nor U730 (N_730,In_1323,In_1631);
nor U731 (N_731,In_2334,In_1363);
nor U732 (N_732,In_1409,In_1111);
nand U733 (N_733,N_125,N_343);
and U734 (N_734,In_420,In_931);
nor U735 (N_735,N_8,In_2010);
or U736 (N_736,In_1326,In_1551);
nand U737 (N_737,In_1444,In_1794);
or U738 (N_738,In_1045,In_1759);
nor U739 (N_739,N_489,In_322);
and U740 (N_740,N_133,In_675);
nor U741 (N_741,In_1672,N_300);
nand U742 (N_742,In_1984,In_386);
xnor U743 (N_743,In_1653,N_307);
nand U744 (N_744,In_627,In_278);
or U745 (N_745,In_70,N_374);
or U746 (N_746,In_2331,In_1829);
or U747 (N_747,In_186,In_1885);
nor U748 (N_748,In_1188,In_177);
nand U749 (N_749,In_1494,In_939);
and U750 (N_750,In_2246,In_940);
nand U751 (N_751,N_566,N_394);
nor U752 (N_752,In_2270,In_116);
and U753 (N_753,In_619,N_437);
or U754 (N_754,N_380,N_15);
nand U755 (N_755,N_424,In_650);
nand U756 (N_756,In_2363,In_1141);
or U757 (N_757,N_254,In_518);
or U758 (N_758,In_1102,N_60);
and U759 (N_759,N_399,N_232);
xor U760 (N_760,In_2235,N_573);
and U761 (N_761,In_459,In_671);
nor U762 (N_762,In_328,In_646);
or U763 (N_763,N_58,In_2139);
and U764 (N_764,In_984,N_313);
or U765 (N_765,In_2449,In_2353);
nand U766 (N_766,N_92,In_1345);
nand U767 (N_767,N_462,N_143);
nand U768 (N_768,In_1199,N_130);
or U769 (N_769,In_834,In_2022);
and U770 (N_770,In_2161,In_1030);
nor U771 (N_771,In_1338,In_218);
and U772 (N_772,In_1355,In_1607);
or U773 (N_773,In_2078,In_539);
and U774 (N_774,In_669,In_839);
or U775 (N_775,In_2194,In_841);
or U776 (N_776,N_339,In_2005);
nand U777 (N_777,N_267,In_463);
nand U778 (N_778,In_1720,In_308);
nand U779 (N_779,In_954,In_1990);
and U780 (N_780,N_527,In_959);
and U781 (N_781,In_2364,In_350);
nor U782 (N_782,In_432,In_1683);
nand U783 (N_783,In_1940,In_1389);
nand U784 (N_784,In_1718,In_79);
nand U785 (N_785,In_783,In_140);
nand U786 (N_786,N_51,N_347);
and U787 (N_787,In_583,In_2261);
or U788 (N_788,N_534,In_813);
or U789 (N_789,N_210,In_445);
and U790 (N_790,In_409,In_2154);
nand U791 (N_791,In_502,In_2425);
and U792 (N_792,In_2016,In_130);
xor U793 (N_793,In_1525,In_1390);
nand U794 (N_794,N_435,In_976);
nand U795 (N_795,In_1059,In_973);
nand U796 (N_796,In_2158,In_2211);
nor U797 (N_797,In_2240,N_195);
and U798 (N_798,In_567,N_530);
nor U799 (N_799,In_1406,In_2316);
nand U800 (N_800,In_25,In_261);
and U801 (N_801,In_1787,In_2120);
nor U802 (N_802,N_440,In_153);
and U803 (N_803,N_740,In_1500);
or U804 (N_804,N_752,In_1478);
nor U805 (N_805,In_411,In_139);
and U806 (N_806,In_1786,In_232);
and U807 (N_807,In_2263,In_2277);
and U808 (N_808,N_548,N_763);
and U809 (N_809,In_1872,In_840);
nor U810 (N_810,N_224,In_687);
or U811 (N_811,In_1297,In_2275);
nor U812 (N_812,In_936,N_718);
or U813 (N_813,In_515,In_1069);
nand U814 (N_814,N_305,In_2115);
xnor U815 (N_815,In_71,N_778);
xnor U816 (N_816,In_1889,In_1073);
nand U817 (N_817,In_811,N_52);
xnor U818 (N_818,In_1104,In_2228);
and U819 (N_819,N_700,N_340);
nand U820 (N_820,N_136,In_300);
and U821 (N_821,In_133,In_1044);
or U822 (N_822,In_252,N_80);
xor U823 (N_823,In_874,In_183);
nor U824 (N_824,In_2209,N_747);
nand U825 (N_825,In_1957,In_847);
or U826 (N_826,N_84,N_164);
nand U827 (N_827,In_335,In_422);
nor U828 (N_828,N_207,In_1841);
and U829 (N_829,N_425,In_228);
and U830 (N_830,N_423,In_1977);
nand U831 (N_831,In_879,In_2264);
or U832 (N_832,In_251,N_172);
nand U833 (N_833,N_687,N_570);
and U834 (N_834,N_723,In_2145);
nor U835 (N_835,N_701,N_671);
nand U836 (N_836,N_368,In_2245);
and U837 (N_837,In_1240,In_1555);
or U838 (N_838,N_441,N_783);
and U839 (N_839,In_1070,In_303);
nand U840 (N_840,In_890,In_1084);
xnor U841 (N_841,In_362,N_297);
xor U842 (N_842,In_1796,In_1246);
or U843 (N_843,In_1876,In_1628);
nor U844 (N_844,In_934,In_525);
nand U845 (N_845,In_2471,N_614);
nor U846 (N_846,In_2003,In_1336);
or U847 (N_847,N_131,In_1837);
xor U848 (N_848,N_216,In_1671);
xnor U849 (N_849,N_121,In_2374);
nor U850 (N_850,N_666,N_228);
nand U851 (N_851,N_692,N_235);
nor U852 (N_852,N_511,In_2454);
and U853 (N_853,In_2170,N_78);
and U854 (N_854,N_115,N_579);
nand U855 (N_855,In_2118,N_538);
or U856 (N_856,N_278,In_2136);
nor U857 (N_857,In_1530,N_541);
or U858 (N_858,In_1191,N_521);
nor U859 (N_859,N_750,N_432);
and U860 (N_860,In_344,In_58);
and U861 (N_861,N_501,In_1264);
xor U862 (N_862,N_91,In_1357);
and U863 (N_863,In_555,In_107);
and U864 (N_864,In_319,N_321);
nand U865 (N_865,In_857,In_744);
and U866 (N_866,N_657,N_203);
or U867 (N_867,In_215,In_2375);
and U868 (N_868,In_34,In_1573);
and U869 (N_869,In_2043,In_1369);
or U870 (N_870,N_22,N_719);
nand U871 (N_871,In_1417,In_1849);
nand U872 (N_872,In_142,In_1605);
nand U873 (N_873,In_454,In_779);
nand U874 (N_874,N_384,N_294);
xor U875 (N_875,In_446,N_586);
nand U876 (N_876,In_1277,In_888);
nand U877 (N_877,In_1456,N_337);
xor U878 (N_878,In_2481,N_429);
nor U879 (N_879,In_466,N_731);
nand U880 (N_880,In_644,In_2152);
nor U881 (N_881,In_1101,In_1925);
and U882 (N_882,In_1434,In_635);
nor U883 (N_883,N_377,In_1952);
nor U884 (N_884,In_1485,N_334);
nand U885 (N_885,N_392,N_649);
xor U886 (N_886,N_574,N_471);
and U887 (N_887,N_35,In_1621);
or U888 (N_888,In_2458,In_894);
nor U889 (N_889,In_716,In_262);
nand U890 (N_890,N_103,In_450);
and U891 (N_891,N_116,In_24);
xor U892 (N_892,N_698,In_184);
xnor U893 (N_893,In_1404,In_483);
or U894 (N_894,In_1117,In_1568);
nor U895 (N_895,In_1202,In_333);
nor U896 (N_896,N_688,In_1427);
xnor U897 (N_897,In_302,In_2477);
nor U898 (N_898,N_490,N_422);
nor U899 (N_899,In_861,In_1008);
or U900 (N_900,In_1147,In_1374);
and U901 (N_901,In_1972,In_808);
nor U902 (N_902,In_264,N_57);
nand U903 (N_903,N_522,N_427);
nand U904 (N_904,In_732,In_19);
nor U905 (N_905,In_844,In_2397);
nor U906 (N_906,N_590,In_1014);
and U907 (N_907,In_2072,In_510);
or U908 (N_908,N_225,In_2162);
nor U909 (N_909,In_151,In_147);
nand U910 (N_910,In_2119,In_1384);
and U911 (N_911,N_364,In_1257);
and U912 (N_912,N_99,In_222);
xor U913 (N_913,In_1751,N_785);
nand U914 (N_914,In_449,In_1652);
nor U915 (N_915,In_91,N_651);
or U916 (N_916,In_4,N_696);
or U917 (N_917,N_493,N_261);
nor U918 (N_918,N_765,N_608);
nand U919 (N_919,In_624,In_1208);
and U920 (N_920,In_416,N_746);
nor U921 (N_921,In_203,In_154);
or U922 (N_922,In_1180,N_571);
xnor U923 (N_923,In_1380,In_389);
nor U924 (N_924,In_180,In_534);
nand U925 (N_925,In_121,N_250);
xnor U926 (N_926,In_225,In_2393);
or U927 (N_927,In_804,N_332);
and U928 (N_928,In_667,In_2489);
and U929 (N_929,N_196,In_2337);
nor U930 (N_930,In_780,In_690);
xnor U931 (N_931,N_264,N_292);
nand U932 (N_932,In_1701,In_1283);
nand U933 (N_933,In_2346,In_821);
nand U934 (N_934,In_2190,N_491);
nor U935 (N_935,N_513,N_376);
and U936 (N_936,In_1006,N_611);
and U937 (N_937,In_1861,In_176);
or U938 (N_938,In_843,In_1765);
or U939 (N_939,N_798,In_1879);
nand U940 (N_940,N_220,N_199);
nand U941 (N_941,N_282,N_390);
nand U942 (N_942,In_823,N_470);
xor U943 (N_943,N_636,In_718);
nor U944 (N_944,In_234,In_2067);
nor U945 (N_945,In_47,In_1598);
and U946 (N_946,In_1639,In_1921);
or U947 (N_947,In_1888,In_346);
nand U948 (N_948,In_820,In_1963);
and U949 (N_949,N_382,N_754);
nand U950 (N_950,N_465,N_772);
nor U951 (N_951,N_606,In_938);
xor U952 (N_952,N_192,In_1074);
or U953 (N_953,In_1807,In_1587);
nor U954 (N_954,In_508,In_645);
nor U955 (N_955,In_1622,In_730);
nor U956 (N_956,In_923,N_756);
nand U957 (N_957,N_166,N_90);
nor U958 (N_958,N_134,In_613);
xor U959 (N_959,In_1588,In_2408);
or U960 (N_960,In_2429,In_889);
and U961 (N_961,In_48,N_385);
and U962 (N_962,N_344,In_966);
and U963 (N_963,N_535,N_355);
xnor U964 (N_964,In_1408,N_322);
nor U965 (N_965,N_316,N_346);
nor U966 (N_966,In_632,N_34);
and U967 (N_967,In_55,N_11);
xnor U968 (N_968,In_2342,N_650);
nor U969 (N_969,In_1815,N_630);
and U970 (N_970,N_648,N_755);
and U971 (N_971,N_793,In_766);
nand U972 (N_972,N_67,N_237);
nor U973 (N_973,In_1347,N_222);
or U974 (N_974,N_7,In_2036);
nor U975 (N_975,In_2248,In_961);
nand U976 (N_976,In_1855,In_306);
nor U977 (N_977,In_2351,N_737);
nor U978 (N_978,In_267,N_444);
or U979 (N_979,In_348,In_1192);
nand U980 (N_980,In_1563,In_1636);
or U981 (N_981,In_859,N_308);
or U982 (N_982,N_211,N_301);
nor U983 (N_983,In_1479,N_395);
nor U984 (N_984,N_565,In_2208);
nand U985 (N_985,N_708,In_1385);
nand U986 (N_986,In_361,In_2496);
and U987 (N_987,In_1161,In_2004);
nand U988 (N_988,In_178,In_1930);
and U989 (N_989,In_2431,In_1307);
xnor U990 (N_990,In_1961,In_1760);
and U991 (N_991,In_321,In_886);
nor U992 (N_992,In_1712,In_1978);
and U993 (N_993,N_387,N_634);
and U994 (N_994,In_1470,N_430);
nor U995 (N_995,In_60,In_865);
nor U996 (N_996,In_1262,N_738);
nor U997 (N_997,In_1913,In_32);
nand U998 (N_998,In_537,N_202);
or U999 (N_999,In_1022,N_516);
or U1000 (N_1000,In_1473,In_1704);
xor U1001 (N_1001,N_26,In_467);
nor U1002 (N_1002,In_10,In_144);
and U1003 (N_1003,In_1900,In_1634);
nand U1004 (N_1004,In_2306,N_302);
or U1005 (N_1005,In_631,N_669);
and U1006 (N_1006,N_876,N_751);
nand U1007 (N_1007,In_1454,N_652);
and U1008 (N_1008,N_660,In_1238);
and U1009 (N_1009,In_1992,N_77);
or U1010 (N_1010,N_950,N_104);
nand U1011 (N_1011,N_455,N_894);
and U1012 (N_1012,In_457,N_781);
and U1013 (N_1013,In_1904,In_2355);
and U1014 (N_1014,In_1144,N_486);
and U1015 (N_1015,In_1135,N_715);
nand U1016 (N_1016,In_1366,N_120);
nor U1017 (N_1017,In_1946,N_773);
xnor U1018 (N_1018,In_1167,N_933);
or U1019 (N_1019,In_1685,In_1985);
and U1020 (N_1020,In_1145,In_2094);
or U1021 (N_1021,In_1482,In_69);
or U1022 (N_1022,In_2470,In_1331);
and U1023 (N_1023,In_80,N_560);
or U1024 (N_1024,In_1692,In_1166);
nor U1025 (N_1025,In_1762,N_730);
nand U1026 (N_1026,N_801,N_987);
nand U1027 (N_1027,In_2048,In_1580);
and U1028 (N_1028,In_1290,N_190);
or U1029 (N_1029,In_2499,In_797);
nor U1030 (N_1030,In_413,In_2380);
or U1031 (N_1031,In_2403,N_812);
and U1032 (N_1032,In_790,N_279);
and U1033 (N_1033,N_873,In_727);
nor U1034 (N_1034,In_853,In_263);
nor U1035 (N_1035,N_787,In_1491);
nand U1036 (N_1036,N_838,N_354);
nor U1037 (N_1037,N_345,In_1437);
xnor U1038 (N_1038,N_833,In_1529);
and U1039 (N_1039,N_30,In_2467);
nor U1040 (N_1040,N_180,In_1609);
and U1041 (N_1041,N_461,In_7);
nor U1042 (N_1042,In_1256,In_1847);
nand U1043 (N_1043,In_980,In_2290);
and U1044 (N_1044,In_235,N_433);
or U1045 (N_1045,N_760,In_1629);
nor U1046 (N_1046,N_767,N_780);
and U1047 (N_1047,N_488,In_1498);
and U1048 (N_1048,N_73,N_668);
and U1049 (N_1049,In_1177,N_413);
and U1050 (N_1050,N_243,N_839);
nand U1051 (N_1051,In_2230,In_2412);
nor U1052 (N_1052,N_744,In_238);
and U1053 (N_1053,N_771,In_358);
nor U1054 (N_1054,In_612,N_317);
nand U1055 (N_1055,In_880,N_951);
nand U1056 (N_1056,N_921,N_994);
nand U1057 (N_1057,N_508,In_751);
xor U1058 (N_1058,In_2249,In_642);
and U1059 (N_1059,In_90,N_540);
nand U1060 (N_1060,N_379,In_2059);
or U1061 (N_1061,In_2184,In_0);
or U1062 (N_1062,N_712,N_583);
nand U1063 (N_1063,N_326,In_1165);
and U1064 (N_1064,In_731,In_326);
and U1065 (N_1065,N_790,N_811);
nand U1066 (N_1066,In_1859,N_460);
and U1067 (N_1067,In_2488,In_1684);
or U1068 (N_1068,N_803,N_485);
or U1069 (N_1069,In_2280,In_1620);
xnor U1070 (N_1070,N_39,In_1311);
or U1071 (N_1071,N_572,In_529);
or U1072 (N_1072,N_815,N_937);
and U1073 (N_1073,In_1289,N_866);
and U1074 (N_1074,In_792,In_1989);
and U1075 (N_1075,In_610,N_241);
or U1076 (N_1076,In_84,N_916);
nand U1077 (N_1077,In_194,N_10);
and U1078 (N_1078,In_1521,In_2391);
nor U1079 (N_1079,N_206,In_357);
nand U1080 (N_1080,In_1557,N_383);
and U1081 (N_1081,In_1778,In_1955);
or U1082 (N_1082,In_1538,N_962);
nand U1083 (N_1083,In_1769,N_555);
or U1084 (N_1084,In_2132,N_857);
nand U1085 (N_1085,In_2283,In_2416);
xor U1086 (N_1086,N_762,In_2336);
nor U1087 (N_1087,N_956,In_1222);
and U1088 (N_1088,N_550,In_89);
nor U1089 (N_1089,N_804,N_482);
nor U1090 (N_1090,In_1244,N_262);
or U1091 (N_1091,In_1916,In_2329);
xor U1092 (N_1092,In_507,N_678);
and U1093 (N_1093,In_2032,In_1433);
or U1094 (N_1094,N_179,In_946);
nor U1095 (N_1095,In_336,In_385);
nand U1096 (N_1096,N_372,In_1979);
and U1097 (N_1097,N_888,N_551);
nand U1098 (N_1098,In_1334,N_598);
and U1099 (N_1099,In_453,In_715);
nor U1100 (N_1100,N_363,In_1774);
or U1101 (N_1101,N_411,N_881);
or U1102 (N_1102,In_2089,N_582);
nor U1103 (N_1103,N_749,N_296);
nor U1104 (N_1104,N_632,N_761);
nor U1105 (N_1105,In_2110,In_1773);
or U1106 (N_1106,In_1655,In_1666);
and U1107 (N_1107,N_633,In_2177);
and U1108 (N_1108,In_1695,N_769);
or U1109 (N_1109,In_2419,N_500);
or U1110 (N_1110,N_638,In_1953);
nand U1111 (N_1111,In_36,N_799);
and U1112 (N_1112,N_82,In_603);
xor U1113 (N_1113,N_970,In_1599);
and U1114 (N_1114,N_110,In_1072);
and U1115 (N_1115,In_2327,N_330);
or U1116 (N_1116,In_1137,In_1349);
nor U1117 (N_1117,In_1146,In_1624);
or U1118 (N_1118,N_759,N_415);
nor U1119 (N_1119,N_362,N_446);
and U1120 (N_1120,N_561,N_917);
nand U1121 (N_1121,In_696,In_2054);
nor U1122 (N_1122,In_1488,In_21);
or U1123 (N_1123,In_1468,N_845);
nand U1124 (N_1124,In_630,In_1537);
or U1125 (N_1125,In_1154,In_2131);
and U1126 (N_1126,In_1510,N_626);
xor U1127 (N_1127,N_545,In_1943);
nor U1128 (N_1128,In_1824,N_265);
nor U1129 (N_1129,N_564,In_2324);
nand U1130 (N_1130,In_216,In_383);
nand U1131 (N_1131,In_1316,In_1960);
xor U1132 (N_1132,In_2411,In_1753);
nand U1133 (N_1133,In_442,N_943);
nor U1134 (N_1134,In_1766,In_770);
or U1135 (N_1135,In_2216,In_2388);
nor U1136 (N_1136,N_64,In_1026);
nor U1137 (N_1137,N_859,In_200);
or U1138 (N_1138,N_532,N_931);
or U1139 (N_1139,N_971,In_1543);
xnor U1140 (N_1140,N_623,N_138);
or U1141 (N_1141,In_227,In_2423);
and U1142 (N_1142,N_757,N_498);
nand U1143 (N_1143,N_961,N_724);
or U1144 (N_1144,In_702,N_594);
nand U1145 (N_1145,In_2176,N_526);
nand U1146 (N_1146,In_868,In_2487);
nand U1147 (N_1147,N_945,N_867);
nor U1148 (N_1148,N_442,In_647);
or U1149 (N_1149,In_1881,N_728);
nor U1150 (N_1150,In_462,N_567);
xor U1151 (N_1151,N_973,In_738);
or U1152 (N_1152,N_520,In_754);
nor U1153 (N_1153,N_159,N_23);
or U1154 (N_1154,In_1337,In_2456);
nor U1155 (N_1155,In_691,In_1981);
nand U1156 (N_1156,N_388,N_408);
and U1157 (N_1157,In_78,N_20);
nand U1158 (N_1158,In_1125,N_147);
or U1159 (N_1159,In_266,N_451);
nand U1160 (N_1160,In_1464,In_1923);
and U1161 (N_1161,In_2167,N_401);
or U1162 (N_1162,N_870,In_960);
and U1163 (N_1163,N_908,In_728);
and U1164 (N_1164,In_1638,In_665);
and U1165 (N_1165,N_645,In_785);
nor U1166 (N_1166,In_375,In_2135);
or U1167 (N_1167,N_589,In_125);
nand U1168 (N_1168,In_786,In_2445);
nor U1169 (N_1169,In_2344,In_1051);
nand U1170 (N_1170,In_182,N_969);
and U1171 (N_1171,N_802,In_1254);
nand U1172 (N_1172,In_482,In_1031);
nor U1173 (N_1173,N_438,In_1649);
nor U1174 (N_1174,In_703,In_1585);
nand U1175 (N_1175,N_274,In_369);
or U1176 (N_1176,In_1503,N_832);
nand U1177 (N_1177,N_310,N_2);
nand U1178 (N_1178,In_1127,In_1719);
nor U1179 (N_1179,N_826,N_808);
or U1180 (N_1180,In_1426,In_1728);
and U1181 (N_1181,In_1850,N_865);
and U1182 (N_1182,In_1197,In_1150);
nand U1183 (N_1183,In_673,In_2304);
nor U1184 (N_1184,N_847,In_2459);
and U1185 (N_1185,In_882,In_2224);
and U1186 (N_1186,N_436,In_1064);
or U1187 (N_1187,In_479,In_1843);
nor U1188 (N_1188,N_443,N_375);
or U1189 (N_1189,In_1368,In_2479);
nor U1190 (N_1190,N_953,In_902);
nand U1191 (N_1191,In_2377,N_889);
nor U1192 (N_1192,In_498,In_864);
nor U1193 (N_1193,In_26,In_313);
nand U1194 (N_1194,N_944,N_596);
nor U1195 (N_1195,In_2293,In_2271);
and U1196 (N_1196,In_2029,In_896);
or U1197 (N_1197,N_705,In_1902);
and U1198 (N_1198,In_475,N_896);
and U1199 (N_1199,N_260,N_431);
and U1200 (N_1200,N_1023,In_1393);
nand U1201 (N_1201,N_861,In_2396);
nor U1202 (N_1202,N_1060,N_1001);
nor U1203 (N_1203,In_832,In_165);
nor U1204 (N_1204,N_209,In_224);
and U1205 (N_1205,In_711,N_766);
nand U1206 (N_1206,N_1012,In_802);
nor U1207 (N_1207,In_618,N_1090);
xor U1208 (N_1208,N_985,In_680);
or U1209 (N_1209,In_291,N_1115);
or U1210 (N_1210,N_1169,In_2007);
or U1211 (N_1211,In_2220,N_995);
or U1212 (N_1212,In_1994,In_1415);
nand U1213 (N_1213,In_2309,N_544);
nand U1214 (N_1214,N_528,In_1722);
and U1215 (N_1215,In_803,N_578);
nand U1216 (N_1216,In_1673,N_681);
nand U1217 (N_1217,N_342,N_928);
and U1218 (N_1218,N_517,In_1383);
or U1219 (N_1219,In_932,In_434);
xnor U1220 (N_1220,In_1189,N_892);
nand U1221 (N_1221,N_854,N_1179);
and U1222 (N_1222,N_477,N_449);
xnor U1223 (N_1223,N_794,In_1379);
xor U1224 (N_1224,N_670,N_915);
nand U1225 (N_1225,N_93,N_1114);
nor U1226 (N_1226,In_1476,In_275);
nand U1227 (N_1227,In_1505,N_869);
and U1228 (N_1228,N_251,In_924);
nor U1229 (N_1229,In_189,N_1101);
and U1230 (N_1230,N_16,N_601);
nand U1231 (N_1231,N_1162,In_1304);
nor U1232 (N_1232,In_1078,N_941);
or U1233 (N_1233,In_989,N_577);
and U1234 (N_1234,N_146,In_943);
xnor U1235 (N_1235,N_562,N_536);
xnor U1236 (N_1236,In_265,In_2287);
nand U1237 (N_1237,N_453,In_41);
or U1238 (N_1238,N_842,N_697);
or U1239 (N_1239,In_2095,In_1138);
nand U1240 (N_1240,N_710,In_2212);
or U1241 (N_1241,N_117,In_2191);
nor U1242 (N_1242,N_242,In_1508);
and U1243 (N_1243,N_1098,N_1199);
xor U1244 (N_1244,In_1299,N_1033);
and U1245 (N_1245,In_2098,N_711);
and U1246 (N_1246,In_1999,N_102);
nor U1247 (N_1247,In_1489,In_763);
or U1248 (N_1248,N_537,N_725);
and U1249 (N_1249,N_1079,N_849);
and U1250 (N_1250,In_239,In_1432);
nor U1251 (N_1251,N_1111,In_1897);
xnor U1252 (N_1252,N_677,In_2430);
and U1253 (N_1253,N_79,N_418);
xor U1254 (N_1254,N_824,In_1465);
nand U1255 (N_1255,In_1905,N_927);
and U1256 (N_1256,N_1192,In_947);
nor U1257 (N_1257,In_544,In_304);
or U1258 (N_1258,N_581,In_1294);
nor U1259 (N_1259,In_909,In_226);
and U1260 (N_1260,In_1492,In_1419);
and U1261 (N_1261,In_1094,In_935);
nor U1262 (N_1262,In_967,In_2122);
nor U1263 (N_1263,In_1617,N_205);
or U1264 (N_1264,In_2436,In_2198);
xnor U1265 (N_1265,N_1155,In_670);
nor U1266 (N_1266,N_1164,In_339);
or U1267 (N_1267,N_1057,In_855);
nor U1268 (N_1268,N_850,In_948);
nand U1269 (N_1269,N_1131,N_370);
nor U1270 (N_1270,N_817,N_404);
nor U1271 (N_1271,In_212,N_880);
and U1272 (N_1272,In_1200,In_248);
and U1273 (N_1273,N_878,N_1040);
nor U1274 (N_1274,In_607,N_27);
and U1275 (N_1275,N_234,N_949);
and U1276 (N_1276,In_1083,In_1158);
and U1277 (N_1277,In_1845,N_739);
and U1278 (N_1278,N_922,N_736);
and U1279 (N_1279,In_2446,N_646);
nor U1280 (N_1280,N_946,N_914);
or U1281 (N_1281,N_291,In_1651);
nand U1282 (N_1282,In_2368,In_704);
nor U1283 (N_1283,N_1095,N_947);
nor U1284 (N_1284,In_1100,In_1274);
nand U1285 (N_1285,N_635,In_1668);
or U1286 (N_1286,In_2017,In_332);
nand U1287 (N_1287,N_200,N_1039);
xnor U1288 (N_1288,N_1092,N_1150);
or U1289 (N_1289,N_1055,N_689);
or U1290 (N_1290,N_475,N_333);
and U1291 (N_1291,N_403,In_1506);
nor U1292 (N_1292,In_1291,N_1146);
xnor U1293 (N_1293,N_714,In_1801);
nor U1294 (N_1294,N_554,In_2422);
or U1295 (N_1295,N_1087,In_545);
or U1296 (N_1296,N_396,N_1053);
or U1297 (N_1297,N_758,N_764);
nand U1298 (N_1298,In_50,In_374);
xor U1299 (N_1299,N_1173,In_39);
nand U1300 (N_1300,N_877,In_900);
and U1301 (N_1301,N_463,N_559);
or U1302 (N_1302,N_1028,N_348);
and U1303 (N_1303,N_549,N_1130);
or U1304 (N_1304,N_150,In_407);
and U1305 (N_1305,N_1045,In_1630);
or U1306 (N_1306,N_1097,In_1041);
nor U1307 (N_1307,N_1093,N_898);
and U1308 (N_1308,N_975,N_1134);
nand U1309 (N_1309,N_174,In_1066);
or U1310 (N_1310,N_1086,In_1564);
or U1311 (N_1311,N_855,In_425);
and U1312 (N_1312,N_312,N_1154);
or U1313 (N_1313,In_828,N_1081);
or U1314 (N_1314,N_797,N_329);
and U1315 (N_1315,In_677,In_1566);
xor U1316 (N_1316,In_112,In_1710);
and U1317 (N_1317,In_1937,N_402);
and U1318 (N_1318,In_205,N_524);
nand U1319 (N_1319,N_576,N_903);
nand U1320 (N_1320,N_875,In_237);
and U1321 (N_1321,In_899,In_1648);
xor U1322 (N_1322,In_1584,N_289);
nor U1323 (N_1323,In_14,In_1834);
and U1324 (N_1324,In_1813,N_929);
nand U1325 (N_1325,N_1151,N_690);
or U1326 (N_1326,N_863,In_2362);
nor U1327 (N_1327,N_819,N_86);
xor U1328 (N_1328,In_2312,In_1821);
nand U1329 (N_1329,In_2056,N_1084);
nand U1330 (N_1330,In_1838,N_835);
or U1331 (N_1331,In_969,N_1022);
or U1332 (N_1332,N_902,In_2018);
nand U1333 (N_1333,In_1535,N_523);
or U1334 (N_1334,N_1082,N_607);
nor U1335 (N_1335,N_964,N_726);
xor U1336 (N_1336,N_920,N_621);
xnor U1337 (N_1337,In_663,N_665);
or U1338 (N_1338,In_1988,In_1606);
and U1339 (N_1339,N_868,In_991);
nand U1340 (N_1340,N_745,N_1119);
nor U1341 (N_1341,In_1377,In_2109);
nand U1342 (N_1342,N_930,In_360);
xor U1343 (N_1343,In_231,In_2019);
nand U1344 (N_1344,N_788,N_603);
xor U1345 (N_1345,N_1068,In_513);
xor U1346 (N_1346,N_716,In_1397);
xnor U1347 (N_1347,In_173,In_557);
or U1348 (N_1348,N_940,In_1731);
or U1349 (N_1349,In_1210,In_910);
nand U1350 (N_1350,In_1372,In_827);
or U1351 (N_1351,In_1227,In_347);
or U1352 (N_1352,In_849,In_1160);
xor U1353 (N_1353,N_6,N_791);
or U1354 (N_1354,N_547,N_56);
and U1355 (N_1355,N_1159,In_652);
nand U1356 (N_1356,N_1144,In_258);
or U1357 (N_1357,In_1229,In_1633);
and U1358 (N_1358,N_1014,N_655);
or U1359 (N_1359,N_879,N_1011);
xor U1360 (N_1360,N_298,In_2150);
and U1361 (N_1361,N_1056,N_1189);
nor U1362 (N_1362,N_1015,N_734);
or U1363 (N_1363,In_1729,N_1175);
nor U1364 (N_1364,N_1153,In_2432);
or U1365 (N_1365,In_179,N_702);
nand U1366 (N_1366,In_1596,N_467);
xnor U1367 (N_1367,N_1049,N_183);
xnor U1368 (N_1368,N_679,N_389);
nand U1369 (N_1369,In_1280,In_1040);
and U1370 (N_1370,N_1075,N_152);
nand U1371 (N_1371,N_1197,In_1152);
nor U1372 (N_1372,In_892,In_1268);
or U1373 (N_1373,In_214,In_1831);
and U1374 (N_1374,N_287,N_883);
xor U1375 (N_1375,In_1820,N_1166);
or U1376 (N_1376,N_721,In_253);
and U1377 (N_1377,N_625,In_1164);
nand U1378 (N_1378,In_1714,In_318);
nand U1379 (N_1379,In_1764,N_807);
nand U1380 (N_1380,In_393,In_771);
and U1381 (N_1381,N_775,N_729);
and U1382 (N_1382,In_2201,In_2233);
and U1383 (N_1383,N_420,In_2390);
nand U1384 (N_1384,N_1193,N_1181);
and U1385 (N_1385,N_1138,N_695);
nor U1386 (N_1386,In_1157,N_620);
and U1387 (N_1387,N_1051,N_667);
nor U1388 (N_1388,N_12,In_109);
or U1389 (N_1389,N_934,N_476);
nor U1390 (N_1390,In_1604,In_2053);
nor U1391 (N_1391,In_2080,N_919);
and U1392 (N_1392,N_658,In_1053);
nor U1393 (N_1393,In_1715,In_1029);
nor U1394 (N_1394,N_1009,N_602);
or U1395 (N_1395,N_1152,In_1721);
or U1396 (N_1396,In_290,In_1723);
nand U1397 (N_1397,In_829,N_1145);
and U1398 (N_1398,In_1481,N_840);
and U1399 (N_1399,In_485,N_1182);
nand U1400 (N_1400,N_1121,In_1170);
or U1401 (N_1401,N_1042,N_1364);
or U1402 (N_1402,In_1194,N_795);
xor U1403 (N_1403,N_1135,N_257);
nand U1404 (N_1404,In_108,In_904);
nand U1405 (N_1405,In_1613,In_11);
nand U1406 (N_1406,In_538,In_1018);
nand U1407 (N_1407,N_1099,In_685);
nand U1408 (N_1408,In_2,N_963);
nand U1409 (N_1409,N_518,N_1207);
nor U1410 (N_1410,N_595,In_123);
nor U1411 (N_1411,N_1139,In_1453);
nor U1412 (N_1412,N_452,In_2466);
and U1413 (N_1413,N_1085,N_45);
or U1414 (N_1414,N_1279,N_662);
or U1415 (N_1415,N_1044,In_1546);
nor U1416 (N_1416,N_1373,In_1301);
xnor U1417 (N_1417,N_154,In_1910);
or U1418 (N_1418,N_81,N_1021);
xnor U1419 (N_1419,N_1335,In_8);
and U1420 (N_1420,N_327,In_210);
nor U1421 (N_1421,N_741,N_600);
or U1422 (N_1422,In_908,In_2021);
or U1423 (N_1423,In_734,N_918);
and U1424 (N_1424,In_611,In_1236);
nand U1425 (N_1425,In_1947,N_1186);
nand U1426 (N_1426,In_2244,N_1247);
and U1427 (N_1427,N_1100,In_1228);
nor U1428 (N_1428,N_1143,In_2151);
and U1429 (N_1429,N_111,In_27);
nand U1430 (N_1430,N_397,In_2133);
and U1431 (N_1431,N_1270,N_686);
xor U1432 (N_1432,N_1187,In_1688);
nor U1433 (N_1433,N_906,N_421);
nor U1434 (N_1434,In_1542,N_959);
xnor U1435 (N_1435,In_1445,In_1039);
nand U1436 (N_1436,In_2435,In_1819);
nand U1437 (N_1437,N_1030,N_887);
nor U1438 (N_1438,N_1102,In_2357);
or U1439 (N_1439,N_1122,In_1732);
or U1440 (N_1440,In_719,In_2075);
and U1441 (N_1441,In_88,N_805);
or U1442 (N_1442,N_1198,In_1552);
and U1443 (N_1443,N_557,In_1105);
nor U1444 (N_1444,N_1332,N_1225);
nor U1445 (N_1445,N_654,N_622);
nor U1446 (N_1446,N_605,N_61);
xnor U1447 (N_1447,N_996,N_1331);
or U1448 (N_1448,In_1771,N_1389);
nor U1449 (N_1449,N_454,In_956);
or U1450 (N_1450,In_1399,N_101);
nand U1451 (N_1451,In_1162,In_831);
nand U1452 (N_1452,N_249,N_1237);
nand U1453 (N_1453,N_978,In_764);
nor U1454 (N_1454,N_782,N_1167);
nor U1455 (N_1455,In_1122,In_1795);
and U1456 (N_1456,N_1007,N_1311);
or U1457 (N_1457,In_391,N_1211);
nand U1458 (N_1458,In_506,In_2472);
or U1459 (N_1459,In_236,N_1305);
and U1460 (N_1460,N_707,N_1374);
xor U1461 (N_1461,N_1377,N_221);
nor U1462 (N_1462,In_2485,N_1357);
nand U1463 (N_1463,In_1998,N_1204);
nand U1464 (N_1464,In_2060,N_882);
and U1465 (N_1465,N_1328,In_1667);
nand U1466 (N_1466,N_1020,N_1341);
nand U1467 (N_1467,In_1558,In_604);
or U1468 (N_1468,In_1909,In_2462);
and U1469 (N_1469,In_2297,N_1251);
or U1470 (N_1470,N_1083,In_1970);
nand U1471 (N_1471,In_22,In_1226);
nor U1472 (N_1472,N_1310,N_843);
xor U1473 (N_1473,N_1096,In_38);
nor U1474 (N_1474,N_50,In_816);
nor U1475 (N_1475,N_828,N_1327);
nand U1476 (N_1476,N_1107,In_569);
nand U1477 (N_1477,N_1160,N_428);
or U1478 (N_1478,In_777,In_1442);
nor U1479 (N_1479,N_170,In_697);
nand U1480 (N_1480,In_1024,In_2192);
or U1481 (N_1481,In_440,In_396);
and U1482 (N_1482,N_1047,In_2494);
nor U1483 (N_1483,N_968,N_809);
nand U1484 (N_1484,In_2341,N_1171);
and U1485 (N_1485,N_997,N_1337);
nor U1486 (N_1486,In_1743,N_1206);
or U1487 (N_1487,N_1219,In_2410);
and U1488 (N_1488,N_492,N_1036);
nor U1489 (N_1489,In_499,N_479);
xor U1490 (N_1490,N_1387,N_108);
or U1491 (N_1491,N_1080,In_56);
nor U1492 (N_1492,N_1017,In_814);
and U1493 (N_1493,N_1073,N_542);
or U1494 (N_1494,In_2015,N_506);
and U1495 (N_1495,N_1330,In_481);
or U1496 (N_1496,N_1067,N_1396);
nor U1497 (N_1497,N_87,N_76);
or U1498 (N_1498,N_722,N_1125);
nand U1499 (N_1499,N_1200,In_257);
xor U1500 (N_1500,In_2424,In_2193);
nand U1501 (N_1501,N_1046,N_932);
and U1502 (N_1502,N_1329,N_407);
or U1503 (N_1503,N_1343,N_552);
or U1504 (N_1504,N_821,N_784);
nand U1505 (N_1505,N_1334,N_320);
nor U1506 (N_1506,In_2178,N_1306);
or U1507 (N_1507,In_1049,N_439);
and U1508 (N_1508,N_1368,N_704);
nand U1509 (N_1509,In_1354,N_1297);
nor U1510 (N_1510,In_1705,In_1702);
nand U1511 (N_1511,In_1225,N_1392);
nand U1512 (N_1512,N_592,In_1168);
or U1513 (N_1513,In_575,In_1894);
nand U1514 (N_1514,In_134,In_1524);
nor U1515 (N_1515,N_1271,In_625);
nor U1516 (N_1516,N_1113,N_1163);
or U1517 (N_1517,N_268,N_706);
nor U1518 (N_1518,N_1127,In_739);
nor U1519 (N_1519,In_478,N_1295);
and U1520 (N_1520,N_814,In_2313);
nor U1521 (N_1521,N_226,N_1259);
nand U1522 (N_1522,N_1091,In_2433);
xnor U1523 (N_1523,N_525,N_862);
nor U1524 (N_1524,N_893,N_1293);
nor U1525 (N_1525,In_2107,N_1264);
xnor U1526 (N_1526,In_395,N_1054);
and U1527 (N_1527,N_1322,N_1356);
nand U1528 (N_1528,N_124,N_1191);
nor U1529 (N_1529,In_2237,N_972);
and U1530 (N_1530,N_1339,N_818);
nor U1531 (N_1531,N_1183,In_1711);
nand U1532 (N_1532,N_304,In_883);
or U1533 (N_1533,In_740,In_270);
and U1534 (N_1534,N_1016,N_816);
and U1535 (N_1535,In_1545,N_459);
nor U1536 (N_1536,In_897,N_43);
xor U1537 (N_1537,N_46,N_942);
nand U1538 (N_1538,In_1436,In_641);
nor U1539 (N_1539,N_1314,In_451);
or U1540 (N_1540,In_1480,In_1806);
nor U1541 (N_1541,In_2187,N_1383);
xor U1542 (N_1542,N_904,N_1378);
nor U1543 (N_1543,N_1027,N_1109);
and U1544 (N_1544,In_1315,N_999);
nand U1545 (N_1545,In_953,N_948);
and U1546 (N_1546,N_271,N_1375);
nand U1547 (N_1547,N_391,In_1412);
nand U1548 (N_1548,In_2066,N_361);
and U1549 (N_1549,In_1775,N_1064);
nand U1550 (N_1550,N_1124,N_1129);
and U1551 (N_1551,N_283,N_466);
and U1552 (N_1552,N_1117,N_864);
and U1553 (N_1553,N_675,In_2299);
nand U1554 (N_1554,N_1280,N_123);
xor U1555 (N_1555,In_404,In_1271);
xnor U1556 (N_1556,N_214,N_331);
or U1557 (N_1557,In_1611,In_1365);
or U1558 (N_1558,In_1255,N_1089);
nand U1559 (N_1559,In_758,In_293);
nor U1560 (N_1560,N_1205,In_351);
nor U1561 (N_1561,N_1019,N_1195);
nand U1562 (N_1562,N_647,In_1449);
and U1563 (N_1563,N_909,N_1319);
nor U1564 (N_1564,In_494,N_1398);
nand U1565 (N_1565,In_1548,N_939);
xor U1566 (N_1566,In_2100,N_998);
nand U1567 (N_1567,In_185,N_1240);
and U1568 (N_1568,In_471,In_593);
nand U1569 (N_1569,N_144,In_760);
and U1570 (N_1570,N_580,N_1312);
nor U1571 (N_1571,N_593,N_1287);
and U1572 (N_1572,N_967,N_456);
and U1573 (N_1573,N_1088,In_1515);
or U1574 (N_1574,N_1137,In_132);
and U1575 (N_1575,In_281,In_2073);
nor U1576 (N_1576,N_955,N_806);
nor U1577 (N_1577,In_429,N_673);
nand U1578 (N_1578,N_1333,N_1386);
nand U1579 (N_1579,N_618,In_2354);
nor U1580 (N_1580,In_2463,N_913);
and U1581 (N_1581,N_597,N_1303);
nor U1582 (N_1582,N_1229,N_29);
nand U1583 (N_1583,In_1496,N_503);
nand U1584 (N_1584,In_316,N_1394);
and U1585 (N_1585,N_487,In_1057);
nor U1586 (N_1586,In_957,N_966);
or U1587 (N_1587,N_990,N_1244);
xor U1588 (N_1588,N_1156,N_988);
nor U1589 (N_1589,N_1230,In_424);
and U1590 (N_1590,In_559,In_1279);
nor U1591 (N_1591,N_1037,In_85);
nand U1592 (N_1592,In_822,In_2055);
and U1593 (N_1593,N_1032,N_1243);
nor U1594 (N_1594,N_991,In_2251);
and U1595 (N_1595,In_387,N_126);
nand U1596 (N_1596,N_1013,N_1380);
nand U1597 (N_1597,In_1740,In_444);
xor U1598 (N_1598,In_997,N_1226);
xnor U1599 (N_1599,N_1382,N_974);
and U1600 (N_1600,N_1349,In_794);
xnor U1601 (N_1601,N_1004,In_987);
nand U1602 (N_1602,N_720,N_1212);
nand U1603 (N_1603,N_1252,In_1654);
and U1604 (N_1604,In_1699,In_1635);
nand U1605 (N_1605,N_510,In_82);
or U1606 (N_1606,In_1155,N_900);
nor U1607 (N_1607,N_1250,In_778);
nand U1608 (N_1608,N_1043,N_830);
nand U1609 (N_1609,N_1509,In_775);
and U1610 (N_1610,N_1320,N_1103);
nor U1611 (N_1611,In_201,In_937);
and U1612 (N_1612,N_1447,N_856);
nor U1613 (N_1613,N_1585,In_473);
and U1614 (N_1614,N_1575,In_161);
or U1615 (N_1615,N_98,In_1544);
or U1616 (N_1616,N_713,N_1561);
and U1617 (N_1617,N_293,In_1043);
and U1618 (N_1618,N_1568,N_1354);
and U1619 (N_1619,N_100,N_1170);
nor U1620 (N_1620,N_1262,In_464);
and U1621 (N_1621,In_1920,N_1110);
or U1622 (N_1622,N_1434,N_480);
and U1623 (N_1623,N_1094,N_409);
nor U1624 (N_1624,N_1344,N_1479);
or U1625 (N_1625,N_1524,N_191);
or U1626 (N_1626,N_507,N_558);
xnor U1627 (N_1627,N_410,N_1172);
xnor U1628 (N_1628,N_631,N_1555);
nand U1629 (N_1629,In_289,N_1307);
or U1630 (N_1630,N_1563,In_2180);
xnor U1631 (N_1631,In_1391,In_1252);
nor U1632 (N_1632,N_1041,In_590);
and U1633 (N_1633,N_328,N_1451);
or U1634 (N_1634,N_1457,N_682);
nand U1635 (N_1635,N_954,In_681);
nand U1636 (N_1636,In_521,In_307);
and U1637 (N_1637,N_1345,In_1394);
and U1638 (N_1638,N_1469,N_659);
nor U1639 (N_1639,N_848,N_236);
nor U1640 (N_1640,In_869,N_280);
or U1641 (N_1641,In_1149,N_1133);
nand U1642 (N_1642,N_1507,In_1594);
and U1643 (N_1643,In_2376,In_40);
nor U1644 (N_1644,N_1545,In_2399);
and U1645 (N_1645,N_1588,N_1541);
and U1646 (N_1646,N_499,In_1013);
nor U1647 (N_1647,N_543,N_1077);
and U1648 (N_1648,In_102,N_905);
nand U1649 (N_1649,N_624,N_1291);
xor U1650 (N_1650,In_1880,N_1358);
xor U1651 (N_1651,In_549,N_674);
nand U1652 (N_1652,N_1512,N_259);
nor U1653 (N_1653,N_1559,N_1063);
nand U1654 (N_1654,In_2042,N_895);
nand U1655 (N_1655,N_1257,N_1423);
or U1656 (N_1656,In_2044,N_1210);
nand U1657 (N_1657,N_1126,In_628);
or U1658 (N_1658,N_891,In_1582);
nor U1659 (N_1659,In_1050,N_1564);
nor U1660 (N_1660,N_1534,N_1294);
or U1661 (N_1661,N_884,In_765);
xnor U1662 (N_1662,In_1090,In_769);
nand U1663 (N_1663,N_1276,In_2020);
and U1664 (N_1664,In_856,N_1592);
nand U1665 (N_1665,N_1452,In_2343);
nand U1666 (N_1666,In_793,N_1203);
xor U1667 (N_1667,N_288,N_822);
and U1668 (N_1668,N_653,N_1518);
nand U1669 (N_1669,N_400,N_1454);
and U1670 (N_1670,In_15,N_1569);
nand U1671 (N_1671,In_2442,In_2300);
xor U1672 (N_1672,N_448,In_1840);
xnor U1673 (N_1673,In_1206,In_105);
and U1674 (N_1674,N_1490,In_1716);
and U1675 (N_1675,N_1442,N_1008);
xor U1676 (N_1676,N_1448,N_642);
nor U1677 (N_1677,N_796,In_951);
nand U1678 (N_1678,N_1265,In_528);
xor U1679 (N_1679,In_1559,N_1513);
nand U1680 (N_1680,N_820,N_661);
nor U1681 (N_1681,In_5,N_1256);
and U1682 (N_1682,In_30,N_604);
or U1683 (N_1683,In_1103,N_65);
nand U1684 (N_1684,In_2039,N_1432);
and U1685 (N_1685,N_1024,N_1520);
nor U1686 (N_1686,N_1116,N_230);
xnor U1687 (N_1687,In_160,N_546);
and U1688 (N_1688,In_1441,N_1213);
xnor U1689 (N_1689,N_1527,In_1895);
and U1690 (N_1690,N_1350,In_1911);
nor U1691 (N_1691,N_1006,N_1546);
nand U1692 (N_1692,In_1754,N_1149);
or U1693 (N_1693,N_357,N_1516);
nand U1694 (N_1694,N_1050,N_619);
or U1695 (N_1695,N_1363,N_1438);
nand U1696 (N_1696,N_1388,N_1369);
nand U1697 (N_1697,N_1360,In_817);
nor U1698 (N_1698,N_1220,N_1104);
nand U1699 (N_1699,N_1402,N_1583);
and U1700 (N_1700,N_1292,N_981);
nor U1701 (N_1701,N_1235,In_1643);
or U1702 (N_1702,In_382,N_1526);
or U1703 (N_1703,In_867,N_890);
and U1704 (N_1704,N_1494,In_474);
nor U1705 (N_1705,N_680,N_982);
nor U1706 (N_1706,N_609,N_1263);
or U1707 (N_1707,In_1462,In_550);
and U1708 (N_1708,N_1410,N_1260);
nor U1709 (N_1709,N_1466,N_1180);
and U1710 (N_1710,N_1370,N_834);
nor U1711 (N_1711,N_1362,In_1623);
and U1712 (N_1712,In_1763,N_1413);
or U1713 (N_1713,N_776,N_1161);
nand U1714 (N_1714,N_1463,N_1059);
or U1715 (N_1715,N_656,In_1836);
or U1716 (N_1716,N_1474,In_1457);
and U1717 (N_1717,N_1573,N_1565);
or U1718 (N_1718,In_1954,N_1478);
xnor U1719 (N_1719,N_1342,N_1218);
nor U1720 (N_1720,N_1052,N_1070);
nor U1721 (N_1721,N_529,N_1464);
nand U1722 (N_1722,N_1488,N_118);
or U1723 (N_1723,In_1270,N_1157);
nor U1724 (N_1724,In_2260,N_911);
nor U1725 (N_1725,N_925,In_2360);
and U1726 (N_1726,N_1562,N_1495);
or U1727 (N_1727,N_1486,In_1237);
or U1728 (N_1728,N_844,N_49);
nor U1729 (N_1729,In_651,N_1445);
xor U1730 (N_1730,In_2420,In_692);
or U1731 (N_1731,N_1458,N_1376);
nor U1732 (N_1732,N_1300,N_240);
and U1733 (N_1733,In_542,N_1551);
or U1734 (N_1734,In_2474,N_193);
nand U1735 (N_1735,N_831,N_1428);
nor U1736 (N_1736,In_1148,In_2295);
nor U1737 (N_1737,N_1168,N_774);
nand U1738 (N_1738,N_272,In_1660);
and U1739 (N_1739,N_800,N_188);
nor U1740 (N_1740,In_1452,N_860);
or U1741 (N_1741,In_580,N_709);
nand U1742 (N_1742,N_1018,In_2469);
xor U1743 (N_1743,N_1254,N_717);
nand U1744 (N_1744,N_699,N_135);
and U1745 (N_1745,In_678,N_852);
nand U1746 (N_1746,N_1366,N_1324);
xor U1747 (N_1747,N_640,In_1396);
or U1748 (N_1748,N_208,N_872);
nor U1749 (N_1749,N_641,In_1511);
nor U1750 (N_1750,In_726,N_1594);
nor U1751 (N_1751,N_1002,In_320);
xnor U1752 (N_1752,N_1106,N_37);
nor U1753 (N_1753,N_281,N_676);
nor U1754 (N_1754,N_1176,N_1470);
nor U1755 (N_1755,N_899,In_1864);
nor U1756 (N_1756,N_434,N_1399);
and U1757 (N_1757,N_1598,In_1867);
and U1758 (N_1758,N_897,In_2348);
or U1759 (N_1759,N_733,N_1078);
and U1760 (N_1760,In_571,N_1572);
and U1761 (N_1761,In_1027,N_1239);
or U1762 (N_1762,In_18,N_1108);
nor U1763 (N_1763,N_1026,N_1489);
or U1764 (N_1764,N_539,In_1965);
nand U1765 (N_1765,In_1034,N_1419);
and U1766 (N_1766,In_64,N_1236);
xnor U1767 (N_1767,In_2452,N_1417);
nand U1768 (N_1768,N_1554,In_1108);
nor U1769 (N_1769,In_520,In_6);
nor U1770 (N_1770,In_2307,N_732);
or U1771 (N_1771,N_1471,In_906);
nand U1772 (N_1772,N_1391,In_592);
or U1773 (N_1773,N_1424,N_639);
nand U1774 (N_1774,N_1285,N_1532);
or U1775 (N_1775,N_748,In_679);
nor U1776 (N_1776,In_285,In_501);
nor U1777 (N_1777,N_1313,N_858);
and U1778 (N_1778,N_1455,In_1058);
nor U1779 (N_1779,N_575,N_1499);
xnor U1780 (N_1780,N_979,In_2112);
and U1781 (N_1781,N_615,N_1487);
and U1782 (N_1782,N_1141,N_1482);
or U1783 (N_1783,N_1475,N_1558);
and U1784 (N_1784,N_1234,N_1476);
nor U1785 (N_1785,In_1941,In_43);
nand U1786 (N_1786,N_1112,N_1228);
and U1787 (N_1787,N_468,N_663);
xor U1788 (N_1788,N_1282,N_1496);
nor U1789 (N_1789,N_1446,In_384);
or U1790 (N_1790,In_2123,In_746);
nor U1791 (N_1791,N_874,N_1549);
nand U1792 (N_1792,N_1440,In_1055);
and U1793 (N_1793,N_1299,N_1530);
or U1794 (N_1794,N_62,N_986);
or U1795 (N_1795,N_373,N_1543);
nor U1796 (N_1796,N_1066,N_266);
or U1797 (N_1797,N_553,N_735);
nand U1798 (N_1798,N_1381,N_1427);
nor U1799 (N_1799,In_17,N_1472);
and U1800 (N_1800,In_309,In_2226);
nor U1801 (N_1801,N_1184,N_610);
and U1802 (N_1802,N_215,N_464);
xor U1803 (N_1803,N_1283,N_1048);
nor U1804 (N_1804,N_1485,In_970);
nand U1805 (N_1805,In_2114,N_1253);
and U1806 (N_1806,N_1582,N_1286);
or U1807 (N_1807,N_1760,N_1477);
and U1808 (N_1808,N_1723,N_1460);
and U1809 (N_1809,N_173,In_990);
or U1810 (N_1810,N_1619,N_1684);
or U1811 (N_1811,N_703,N_469);
or U1812 (N_1812,N_1224,N_1725);
xor U1813 (N_1813,In_666,N_1794);
nor U1814 (N_1814,N_1401,N_1693);
or U1815 (N_1815,N_1796,N_753);
nor U1816 (N_1816,N_1689,In_1263);
nor U1817 (N_1817,N_447,N_1700);
and U1818 (N_1818,N_1511,N_119);
or U1819 (N_1819,N_1790,N_1421);
or U1820 (N_1820,In_2012,N_1610);
and U1821 (N_1821,N_958,N_977);
xor U1822 (N_1822,N_1242,N_1694);
and U1823 (N_1823,In_1687,N_1570);
and U1824 (N_1824,N_1185,N_1744);
nand U1825 (N_1825,N_685,N_245);
or U1826 (N_1826,N_1679,N_1449);
or U1827 (N_1827,In_835,In_2395);
and U1828 (N_1828,N_1552,N_672);
xnor U1829 (N_1829,N_1290,N_1395);
nor U1830 (N_1830,N_976,N_983);
nor U1831 (N_1831,N_414,N_1778);
or U1832 (N_1832,N_1223,N_1074);
xnor U1833 (N_1833,N_1456,N_1346);
or U1834 (N_1834,N_1658,In_742);
xnor U1835 (N_1835,N_846,N_1425);
and U1836 (N_1836,In_472,N_1718);
and U1837 (N_1837,N_1418,N_1728);
and U1838 (N_1838,N_1606,N_416);
or U1839 (N_1839,N_1749,N_1351);
nand U1840 (N_1840,N_1667,N_1607);
or U1841 (N_1841,N_960,N_1574);
nor U1842 (N_1842,In_86,N_1730);
and U1843 (N_1843,N_1604,N_1289);
nand U1844 (N_1844,N_1795,N_1590);
nor U1845 (N_1845,N_1682,In_2000);
and U1846 (N_1846,N_1680,N_1523);
xor U1847 (N_1847,In_500,N_156);
and U1848 (N_1848,N_1576,N_1221);
or U1849 (N_1849,N_1517,N_1062);
nand U1850 (N_1850,N_957,In_1931);
nor U1851 (N_1851,N_1731,In_1665);
and U1852 (N_1852,N_1757,In_561);
or U1853 (N_1853,N_1497,N_1272);
nor U1854 (N_1854,N_1609,N_1635);
xor U1855 (N_1855,N_1058,N_1765);
nand U1856 (N_1856,N_1751,N_1702);
nor U1857 (N_1857,In_268,N_1510);
nand U1858 (N_1858,N_1636,N_1706);
nor U1859 (N_1859,N_1698,N_770);
nor U1860 (N_1860,N_1461,N_1709);
and U1861 (N_1861,In_1451,N_1762);
or U1862 (N_1862,N_1174,N_810);
or U1863 (N_1863,N_367,N_1766);
nor U1864 (N_1864,N_1249,N_1735);
nor U1865 (N_1865,N_1632,N_935);
nor U1866 (N_1866,N_1676,N_1281);
nor U1867 (N_1867,In_279,N_1400);
nor U1868 (N_1868,N_1429,In_2272);
nor U1869 (N_1869,N_151,N_1786);
nand U1870 (N_1870,N_406,N_1267);
and U1871 (N_1871,N_1713,In_1495);
nor U1872 (N_1872,N_1238,N_1061);
or U1873 (N_1873,In_761,N_1686);
nand U1874 (N_1874,N_1188,N_1318);
nor U1875 (N_1875,In_1076,N_1118);
nand U1876 (N_1876,N_1355,N_837);
nand U1877 (N_1877,In_1857,N_1750);
nor U1878 (N_1878,N_851,N_1232);
and U1879 (N_1879,N_186,N_1734);
and U1880 (N_1880,N_1727,N_1603);
nand U1881 (N_1881,N_1065,N_1508);
nor U1882 (N_1882,N_1165,N_1614);
and U1883 (N_1883,In_686,N_1653);
and U1884 (N_1884,N_1031,N_1278);
and U1885 (N_1885,N_936,N_1764);
and U1886 (N_1886,N_1404,In_376);
and U1887 (N_1887,In_1005,In_1131);
and U1888 (N_1888,N_1596,N_1678);
or U1889 (N_1889,N_1506,In_661);
nor U1890 (N_1890,N_1771,N_779);
nand U1891 (N_1891,N_1493,N_1784);
xor U1892 (N_1892,N_1540,In_269);
or U1893 (N_1893,N_1537,N_1365);
or U1894 (N_1894,N_1737,N_417);
or U1895 (N_1895,N_1261,N_1000);
and U1896 (N_1896,N_263,In_174);
nor U1897 (N_1897,N_1775,N_1384);
and U1898 (N_1898,N_694,N_1770);
and U1899 (N_1899,In_1021,N_1720);
nand U1900 (N_1900,In_367,N_924);
nand U1901 (N_1901,In_196,N_1255);
nand U1902 (N_1902,N_1755,N_1681);
and U1903 (N_1903,N_1772,N_1640);
nand U1904 (N_1904,N_253,N_1408);
and U1905 (N_1905,N_1674,In_2166);
and U1906 (N_1906,N_1444,N_1618);
nand U1907 (N_1907,In_2370,In_202);
or U1908 (N_1908,In_1590,N_1656);
or U1909 (N_1909,In_1572,In_2352);
and U1910 (N_1910,N_926,N_303);
and U1911 (N_1911,N_1641,N_1608);
nor U1912 (N_1912,In_1407,N_1616);
and U1913 (N_1913,N_637,N_1717);
nor U1914 (N_1914,N_1591,N_792);
nor U1915 (N_1915,N_325,N_1660);
or U1916 (N_1916,N_1481,N_1587);
and U1917 (N_1917,In_188,In_1063);
nand U1918 (N_1918,N_1414,N_1763);
nor U1919 (N_1919,N_1781,In_489);
and U1920 (N_1920,N_1502,In_2305);
nand U1921 (N_1921,N_1215,N_1620);
and U1922 (N_1922,N_1038,N_1633);
nand U1923 (N_1923,In_919,N_1148);
and U1924 (N_1924,N_1785,N_1441);
nor U1925 (N_1925,N_989,N_853);
nor U1926 (N_1926,N_1798,N_923);
nand U1927 (N_1927,In_1644,N_458);
and U1928 (N_1928,N_1359,N_1158);
nand U1929 (N_1929,N_1593,In_197);
and U1930 (N_1930,N_1675,In_54);
or U1931 (N_1931,In_2315,N_28);
xor U1932 (N_1932,N_1622,In_2083);
and U1933 (N_1933,N_1705,N_1274);
and U1934 (N_1934,N_1367,N_1567);
or U1935 (N_1935,N_127,N_1222);
nand U1936 (N_1936,N_13,N_1754);
xor U1937 (N_1937,In_1172,N_1774);
nand U1938 (N_1938,In_148,N_1379);
and U1939 (N_1939,N_1245,In_578);
or U1940 (N_1940,N_1566,N_1782);
nor U1941 (N_1941,N_1298,N_786);
or U1942 (N_1942,N_1637,In_2027);
or U1943 (N_1943,N_617,N_1069);
nand U1944 (N_1944,N_1792,N_1308);
nand U1945 (N_1945,N_1304,In_1770);
nand U1946 (N_1946,N_1538,N_1315);
or U1947 (N_1947,N_992,N_323);
or U1948 (N_1948,N_841,N_644);
nor U1949 (N_1949,N_213,N_1136);
or U1950 (N_1950,N_1246,In_2303);
xnor U1951 (N_1951,In_688,In_621);
nor U1952 (N_1952,N_1768,N_871);
or U1953 (N_1953,N_1268,N_952);
or U1954 (N_1954,N_1630,N_233);
nor U1955 (N_1955,N_1338,N_789);
and U1956 (N_1956,In_654,In_929);
and U1957 (N_1957,N_1703,N_1500);
and U1958 (N_1958,N_1664,N_1140);
and U1959 (N_1959,In_1142,N_1776);
or U1960 (N_1960,N_1787,N_1076);
nor U1961 (N_1961,In_705,N_1397);
nor U1962 (N_1962,N_1657,In_2142);
xor U1963 (N_1963,In_2285,N_1258);
or U1964 (N_1964,N_1696,N_1433);
nand U1965 (N_1965,N_1695,N_1571);
nor U1966 (N_1966,N_1670,N_1147);
nor U1967 (N_1967,N_1560,N_1227);
nor U1968 (N_1968,N_1348,In_2427);
nand U1969 (N_1969,N_1793,In_605);
nand U1970 (N_1970,In_1310,N_1557);
or U1971 (N_1971,In_576,In_193);
or U1972 (N_1972,N_1273,N_1586);
nor U1973 (N_1973,N_1627,N_1752);
nand U1974 (N_1974,N_1643,N_612);
nor U1975 (N_1975,N_139,In_129);
nor U1976 (N_1976,N_1688,N_1756);
and U1977 (N_1977,N_1712,N_1519);
nor U1978 (N_1978,N_1498,In_659);
xnor U1979 (N_1979,N_664,N_1648);
and U1980 (N_1980,N_683,In_2105);
nand U1981 (N_1981,N_1035,N_1409);
and U1982 (N_1982,In_1533,N_1321);
or U1983 (N_1983,N_1316,N_1601);
nand U1984 (N_1984,N_1128,N_1652);
and U1985 (N_1985,In_1614,N_1437);
or U1986 (N_1986,N_1721,N_1733);
nor U1987 (N_1987,N_1791,N_1483);
and U1988 (N_1988,N_1503,N_1767);
nor U1989 (N_1989,N_1634,N_176);
nand U1990 (N_1990,N_629,N_1196);
nand U1991 (N_1991,N_1783,N_1525);
and U1992 (N_1992,In_617,N_1639);
or U1993 (N_1993,N_1542,N_1430);
nand U1994 (N_1994,In_1193,N_1515);
xnor U1995 (N_1995,In_1874,N_628);
or U1996 (N_1996,N_1266,N_1645);
nor U1997 (N_1997,In_2384,In_431);
and U1998 (N_1998,N_1275,N_1480);
xor U1999 (N_1999,N_1553,N_1602);
nand U2000 (N_2000,N_1747,N_1952);
xor U2001 (N_2001,N_1840,N_1945);
or U2002 (N_2002,In_208,N_1915);
nor U2003 (N_2003,In_2038,In_1870);
nand U2004 (N_2004,N_1214,N_1863);
nor U2005 (N_2005,N_613,N_1025);
nor U2006 (N_2006,N_1352,In_863);
xnor U2007 (N_2007,N_1892,In_1707);
nor U2008 (N_2008,N_1820,N_1847);
or U2009 (N_2009,N_1903,N_1626);
nand U2010 (N_2010,N_1901,N_910);
or U2011 (N_2011,In_570,N_627);
nor U2012 (N_2012,In_509,In_2085);
xor U2013 (N_2013,In_1362,N_1966);
nor U2014 (N_2014,N_1909,N_1317);
and U2015 (N_2015,N_1836,N_319);
and U2016 (N_2016,N_1123,N_1842);
or U2017 (N_2017,N_1817,N_1937);
nor U2018 (N_2018,N_1999,N_1789);
nor U2019 (N_2019,N_1724,N_1371);
or U2020 (N_2020,N_1217,In_2113);
nand U2021 (N_2021,N_1822,N_1600);
and U2022 (N_2022,N_993,N_1514);
or U2023 (N_2023,N_1533,N_1529);
or U2024 (N_2024,N_912,N_1912);
xnor U2025 (N_2025,N_1969,N_1473);
and U2026 (N_2026,N_1827,In_851);
or U2027 (N_2027,In_1318,N_1621);
nand U2028 (N_2028,N_1647,N_1977);
and U2029 (N_2029,N_1411,N_227);
and U2030 (N_2030,N_1844,N_1872);
or U2031 (N_2031,N_901,In_1115);
xnor U2032 (N_2032,N_1759,N_1921);
nor U2033 (N_2033,N_1878,In_2002);
and U2034 (N_2034,In_595,N_1416);
and U2035 (N_2035,N_1450,N_1932);
and U2036 (N_2036,N_727,N_1659);
xor U2037 (N_2037,N_1501,N_1880);
nand U2038 (N_2038,N_1858,N_1807);
or U2039 (N_2039,N_1642,N_1231);
nor U2040 (N_2040,N_1005,N_1809);
nand U2041 (N_2041,N_1453,N_1738);
and U2042 (N_2042,N_1898,N_1815);
nor U2043 (N_2043,N_1142,In_1382);
or U2044 (N_2044,N_1935,N_1732);
nor U2045 (N_2045,N_1628,In_259);
xor U2046 (N_2046,In_2404,N_1985);
or U2047 (N_2047,N_1711,In_276);
nor U2048 (N_2048,N_1797,N_1917);
and U2049 (N_2049,N_1690,N_1710);
nand U2050 (N_2050,N_1924,N_938);
or U2051 (N_2051,N_1990,N_1974);
and U2052 (N_2052,N_212,N_813);
xor U2053 (N_2053,N_1665,In_806);
and U2054 (N_2054,N_1535,N_1920);
or U2055 (N_2055,N_1886,N_1739);
nand U2056 (N_2056,N_1323,N_1928);
nor U2057 (N_2057,N_185,N_1965);
nand U2058 (N_2058,In_423,N_1874);
or U2059 (N_2059,N_1629,N_1802);
or U2060 (N_2060,N_1876,N_1860);
nand U2061 (N_2061,N_829,N_1326);
xor U2062 (N_2062,N_1925,N_1962);
xnor U2063 (N_2063,N_827,N_1692);
and U2064 (N_2064,N_1799,N_1971);
nor U2065 (N_2065,N_1034,N_66);
nand U2066 (N_2066,N_1824,N_1811);
nand U2067 (N_2067,N_1816,N_1745);
nand U2068 (N_2068,N_1812,N_505);
and U2069 (N_2069,N_684,N_502);
and U2070 (N_2070,N_1989,N_1504);
and U2071 (N_2071,N_1927,N_1959);
nor U2072 (N_2072,N_1777,N_1010);
and U2073 (N_2073,In_1184,N_1407);
nor U2074 (N_2074,In_1220,In_1922);
nor U2075 (N_2075,N_1856,N_1105);
and U2076 (N_2076,N_1954,N_1578);
nor U2077 (N_2077,In_363,N_1677);
xnor U2078 (N_2078,N_1617,N_1406);
nor U2079 (N_2079,N_1631,N_1867);
nand U2080 (N_2080,N_1857,N_1743);
and U2081 (N_2081,In_167,N_1800);
nor U2082 (N_2082,In_1272,N_1707);
nor U2083 (N_2083,N_1947,N_568);
nor U2084 (N_2084,N_1589,N_1422);
nor U2085 (N_2085,N_1597,N_1851);
nor U2086 (N_2086,N_1548,In_837);
and U2087 (N_2087,N_836,N_1916);
and U2088 (N_2088,In_352,N_886);
nand U2089 (N_2089,N_1853,N_1340);
or U2090 (N_2090,In_1300,N_1655);
nor U2091 (N_2091,N_1850,N_1941);
xnor U2092 (N_2092,N_1813,N_1949);
and U2093 (N_2093,In_157,N_1780);
nand U2094 (N_2094,N_1788,N_1933);
xnor U2095 (N_2095,In_1060,N_1420);
or U2096 (N_2096,N_1580,N_1804);
and U2097 (N_2097,N_1996,N_1875);
nand U2098 (N_2098,N_1716,N_1269);
xnor U2099 (N_2099,N_474,N_1072);
and U2100 (N_2100,N_1987,N_1685);
nand U2101 (N_2101,N_1868,N_1216);
nand U2102 (N_2102,N_1669,N_1887);
xnor U2103 (N_2103,In_435,N_1885);
and U2104 (N_2104,N_1301,N_1870);
or U2105 (N_2105,N_1964,N_1861);
xnor U2106 (N_2106,N_1979,N_1922);
xnor U2107 (N_2107,N_1988,N_1336);
nor U2108 (N_2108,N_1746,N_1654);
or U2109 (N_2109,In_283,N_1761);
or U2110 (N_2110,N_1805,In_505);
or U2111 (N_2111,N_1889,N_1968);
nor U2112 (N_2112,N_1753,N_1855);
nand U2113 (N_2113,N_1910,N_1599);
nor U2114 (N_2114,N_1742,N_1859);
nor U2115 (N_2115,N_1913,N_984);
or U2116 (N_2116,N_1595,N_1862);
or U2117 (N_2117,N_743,N_1704);
nand U2118 (N_2118,N_1995,In_1370);
nand U2119 (N_2119,In_2217,N_1806);
xnor U2120 (N_2120,N_1939,N_1803);
and U2121 (N_2121,N_1845,N_1866);
or U2122 (N_2122,N_1940,N_1668);
and U2123 (N_2123,N_1907,N_1891);
and U2124 (N_2124,N_1646,N_1531);
and U2125 (N_2125,N_1825,In_72);
and U2126 (N_2126,N_1993,N_693);
and U2127 (N_2127,N_1661,N_1325);
nor U2128 (N_2128,In_1982,N_1521);
and U2129 (N_2129,N_1883,N_825);
nand U2130 (N_2130,N_1930,N_1881);
or U2131 (N_2131,N_1848,N_1484);
nor U2132 (N_2132,N_1919,N_1834);
xor U2133 (N_2133,In_1375,N_1843);
nand U2134 (N_2134,N_1492,N_1821);
nor U2135 (N_2135,In_2182,N_1201);
or U2136 (N_2136,N_1869,N_1177);
or U2137 (N_2137,N_1897,N_1906);
nor U2138 (N_2138,N_1405,N_1715);
nor U2139 (N_2139,N_1975,N_1651);
and U2140 (N_2140,N_1773,N_1431);
and U2141 (N_2141,N_1871,In_985);
and U2142 (N_2142,N_1963,In_379);
nand U2143 (N_2143,N_1814,N_1662);
nor U2144 (N_2144,N_768,N_691);
nand U2145 (N_2145,N_1997,N_1961);
nor U2146 (N_2146,N_1612,N_643);
and U2147 (N_2147,N_1003,N_1829);
nand U2148 (N_2148,N_1826,N_1972);
xnor U2149 (N_2149,N_68,N_1828);
and U2150 (N_2150,N_1838,N_1132);
nor U2151 (N_2151,N_495,N_1918);
nor U2152 (N_2152,N_1178,N_1624);
nor U2153 (N_2153,N_1931,N_1741);
nor U2154 (N_2154,In_1295,N_1819);
or U2155 (N_2155,N_1810,N_1719);
or U2156 (N_2156,N_1663,N_1528);
and U2157 (N_2157,N_1459,In_452);
nand U2158 (N_2158,In_1212,N_1967);
or U2159 (N_2159,N_1823,N_1714);
and U2160 (N_2160,N_1296,N_1650);
nor U2161 (N_2161,N_1958,N_1029);
and U2162 (N_2162,N_1412,N_1984);
nor U2163 (N_2163,N_1865,N_1839);
nor U2164 (N_2164,N_1190,N_1353);
and U2165 (N_2165,In_342,N_1248);
and U2166 (N_2166,N_1896,N_1904);
nand U2167 (N_2167,N_1467,In_918);
nand U2168 (N_2168,N_284,N_1944);
nand U2169 (N_2169,N_1726,N_1948);
nor U2170 (N_2170,N_358,N_1929);
or U2171 (N_2171,In_1364,N_1982);
and U2172 (N_2172,N_1701,N_1415);
or U2173 (N_2173,N_1505,N_1908);
or U2174 (N_2174,In_297,N_1539);
and U2175 (N_2175,N_1556,N_1623);
nor U2176 (N_2176,N_1544,N_1831);
nor U2177 (N_2177,N_1818,N_1841);
or U2178 (N_2178,N_1209,In_1275);
and U2179 (N_2179,N_1625,N_1864);
nand U2180 (N_2180,N_1550,N_1309);
or U2181 (N_2181,N_1649,N_484);
nand U2182 (N_2182,In_2082,N_1666);
and U2183 (N_2183,N_1914,N_1978);
and U2184 (N_2184,N_1846,N_563);
and U2185 (N_2185,N_1672,N_1071);
nor U2186 (N_2186,N_1938,N_777);
nand U2187 (N_2187,N_885,N_1436);
nand U2188 (N_2188,N_1983,N_1393);
xor U2189 (N_2189,N_1950,N_1208);
nand U2190 (N_2190,N_33,N_1808);
nor U2191 (N_2191,N_1960,N_1722);
nor U2192 (N_2192,N_1443,N_1740);
and U2193 (N_2193,N_270,N_1882);
and U2194 (N_2194,N_1832,N_1956);
and U2195 (N_2195,In_1934,N_1769);
or U2196 (N_2196,N_1347,N_1953);
or U2197 (N_2197,N_980,N_1638);
or U2198 (N_2198,N_1992,N_1202);
nor U2199 (N_2199,N_1491,N_1683);
nor U2200 (N_2200,N_2050,N_1536);
nor U2201 (N_2201,N_2069,N_2127);
or U2202 (N_2202,N_2077,N_2128);
nand U2203 (N_2203,N_2014,N_2130);
xor U2204 (N_2204,N_1426,N_2046);
and U2205 (N_2205,N_2089,N_2065);
xnor U2206 (N_2206,N_2041,N_2067);
xnor U2207 (N_2207,N_2189,N_2000);
or U2208 (N_2208,N_1233,N_2017);
nand U2209 (N_2209,N_1994,N_2031);
and U2210 (N_2210,N_2039,N_1852);
and U2211 (N_2211,N_1884,N_2152);
nand U2212 (N_2212,N_1615,N_1946);
nor U2213 (N_2213,N_2011,N_2148);
or U2214 (N_2214,N_2134,N_2122);
and U2215 (N_2215,N_1748,N_1911);
and U2216 (N_2216,N_2194,N_2157);
or U2217 (N_2217,N_2172,N_2083);
nand U2218 (N_2218,N_2044,N_1986);
or U2219 (N_2219,N_1691,N_1581);
or U2220 (N_2220,N_2097,N_1439);
nand U2221 (N_2221,N_2058,N_1973);
nand U2222 (N_2222,N_1957,N_2138);
nor U2223 (N_2223,N_1361,N_2188);
or U2224 (N_2224,N_2045,N_2190);
xor U2225 (N_2225,N_1893,N_2166);
nor U2226 (N_2226,N_2082,N_742);
or U2227 (N_2227,N_2020,N_2140);
and U2228 (N_2228,N_2175,N_2005);
nand U2229 (N_2229,N_1462,N_2197);
nand U2230 (N_2230,N_2023,N_1611);
and U2231 (N_2231,N_2125,N_2092);
nand U2232 (N_2232,N_2183,N_1194);
and U2233 (N_2233,N_2080,N_2158);
and U2234 (N_2234,N_2043,N_2033);
and U2235 (N_2235,N_1385,N_2117);
or U2236 (N_2236,N_2078,N_616);
or U2237 (N_2237,N_1801,N_1671);
and U2238 (N_2238,N_2191,N_2001);
nor U2239 (N_2239,N_2101,N_2156);
and U2240 (N_2240,N_1991,N_1970);
nand U2241 (N_2241,N_1936,N_2104);
nor U2242 (N_2242,N_2034,N_1926);
xnor U2243 (N_2243,N_1758,N_2195);
nand U2244 (N_2244,N_1943,N_2013);
xor U2245 (N_2245,N_2192,N_2162);
or U2246 (N_2246,N_2026,N_1673);
nor U2247 (N_2247,N_2179,N_1241);
and U2248 (N_2248,N_2198,In_209);
nand U2249 (N_2249,N_585,N_2151);
and U2250 (N_2250,N_2196,N_2135);
nor U2251 (N_2251,N_1390,N_2016);
and U2252 (N_2252,N_1277,N_2124);
nor U2253 (N_2253,N_2091,N_1854);
and U2254 (N_2254,N_2110,N_149);
nor U2255 (N_2255,N_2076,N_2012);
or U2256 (N_2256,N_1998,N_2113);
and U2257 (N_2257,N_2105,N_2003);
and U2258 (N_2258,N_2030,N_2123);
nor U2259 (N_2259,N_1547,N_2036);
and U2260 (N_2260,N_2167,N_907);
nand U2261 (N_2261,N_2047,N_1699);
and U2262 (N_2262,N_1833,N_2116);
xnor U2263 (N_2263,N_2006,N_1579);
or U2264 (N_2264,N_1522,N_2147);
nor U2265 (N_2265,N_1951,N_2090);
or U2266 (N_2266,N_1877,N_2131);
nor U2267 (N_2267,N_2181,N_1120);
nand U2268 (N_2268,N_2019,N_2093);
and U2269 (N_2269,N_2120,N_2165);
and U2270 (N_2270,N_2060,N_2027);
xnor U2271 (N_2271,N_2098,N_2129);
nand U2272 (N_2272,In_354,N_2074);
and U2273 (N_2273,N_2052,N_1584);
or U2274 (N_2274,N_2199,N_2141);
nand U2275 (N_2275,In_2129,N_2119);
nand U2276 (N_2276,N_2164,N_2009);
and U2277 (N_2277,N_1905,N_2004);
or U2278 (N_2278,N_2062,N_965);
xor U2279 (N_2279,N_2029,N_1613);
and U2280 (N_2280,N_1830,N_1873);
xnor U2281 (N_2281,N_2037,N_258);
nor U2282 (N_2282,N_2084,N_2021);
or U2283 (N_2283,In_1581,N_2168);
and U2284 (N_2284,N_2066,N_2018);
xor U2285 (N_2285,N_1687,N_2068);
or U2286 (N_2286,N_1890,N_2180);
nor U2287 (N_2287,N_2145,N_2112);
or U2288 (N_2288,N_2075,N_2055);
or U2289 (N_2289,N_2100,N_2024);
or U2290 (N_2290,N_2143,N_2184);
xor U2291 (N_2291,N_2010,N_2057);
nand U2292 (N_2292,N_1895,N_1894);
nor U2293 (N_2293,N_2187,N_2049);
nand U2294 (N_2294,N_1837,N_2109);
nor U2295 (N_2295,N_1605,N_2136);
and U2296 (N_2296,N_2154,N_1981);
or U2297 (N_2297,N_1923,N_1980);
nor U2298 (N_2298,N_2028,N_1468);
or U2299 (N_2299,N_2008,N_2161);
and U2300 (N_2300,N_1736,N_1955);
or U2301 (N_2301,N_2025,In_2486);
nand U2302 (N_2302,N_2106,N_2108);
nor U2303 (N_2303,N_1888,N_1729);
nor U2304 (N_2304,N_2153,N_1934);
nand U2305 (N_2305,N_823,N_2048);
nand U2306 (N_2306,N_2177,N_2111);
nor U2307 (N_2307,N_2146,N_2178);
nor U2308 (N_2308,N_1288,In_92);
nand U2309 (N_2309,N_2173,N_2085);
or U2310 (N_2310,N_2007,N_1372);
xor U2311 (N_2311,N_2061,N_1435);
nor U2312 (N_2312,N_1577,N_2176);
xor U2313 (N_2313,N_2149,N_1697);
nor U2314 (N_2314,N_2144,N_2186);
and U2315 (N_2315,N_2087,N_2171);
or U2316 (N_2316,N_1465,N_2079);
xnor U2317 (N_2317,N_2042,N_2053);
or U2318 (N_2318,N_2163,N_1779);
nor U2319 (N_2319,N_1849,N_2072);
nand U2320 (N_2320,N_2182,N_2185);
nand U2321 (N_2321,N_1879,N_2160);
nand U2322 (N_2322,N_1976,N_2137);
nor U2323 (N_2323,N_2054,N_2193);
nor U2324 (N_2324,N_2035,N_2032);
nor U2325 (N_2325,N_1899,N_2115);
nand U2326 (N_2326,N_2174,In_1516);
nand U2327 (N_2327,N_2169,N_2126);
and U2328 (N_2328,N_2139,N_2015);
or U2329 (N_2329,N_2103,N_2070);
nand U2330 (N_2330,N_2051,N_2159);
nor U2331 (N_2331,N_2088,N_1302);
nor U2332 (N_2332,N_2086,N_1708);
nand U2333 (N_2333,N_2155,N_2114);
or U2334 (N_2334,N_2002,N_2150);
nor U2335 (N_2335,N_1900,N_2099);
nor U2336 (N_2336,N_2071,N_1835);
nor U2337 (N_2337,N_2063,N_2073);
and U2338 (N_2338,N_426,N_2022);
and U2339 (N_2339,N_2142,N_2107);
and U2340 (N_2340,N_2038,N_2102);
nor U2341 (N_2341,N_2059,N_2132);
nor U2342 (N_2342,N_2040,N_2094);
nand U2343 (N_2343,N_1644,N_2095);
or U2344 (N_2344,N_2056,N_1403);
or U2345 (N_2345,N_2118,N_1902);
xnor U2346 (N_2346,N_2121,N_1942);
nor U2347 (N_2347,N_2133,N_1284);
nand U2348 (N_2348,N_2081,N_2170);
or U2349 (N_2349,N_2096,N_2064);
xor U2350 (N_2350,N_2071,N_2145);
nor U2351 (N_2351,N_1736,N_2046);
nor U2352 (N_2352,N_1644,N_1849);
xor U2353 (N_2353,N_2152,N_1361);
nand U2354 (N_2354,N_2178,N_2095);
nand U2355 (N_2355,N_2026,N_2042);
or U2356 (N_2356,N_2049,N_2046);
nand U2357 (N_2357,N_1943,N_1673);
nor U2358 (N_2358,N_2080,N_2186);
nand U2359 (N_2359,N_2198,N_2063);
nor U2360 (N_2360,N_2138,N_2124);
nand U2361 (N_2361,N_2006,N_2114);
nor U2362 (N_2362,N_2098,N_2077);
or U2363 (N_2363,N_2082,N_2056);
nand U2364 (N_2364,N_1888,N_2144);
xnor U2365 (N_2365,N_2012,N_1900);
nand U2366 (N_2366,N_1468,N_1801);
nor U2367 (N_2367,N_1893,N_2026);
nand U2368 (N_2368,N_1403,N_2019);
xnor U2369 (N_2369,N_1644,N_2064);
nor U2370 (N_2370,N_2017,N_1361);
nor U2371 (N_2371,N_1902,N_2133);
and U2372 (N_2372,N_2004,N_2175);
or U2373 (N_2373,N_823,N_1288);
xnor U2374 (N_2374,N_585,N_1435);
xor U2375 (N_2375,N_2163,N_2184);
nor U2376 (N_2376,N_2095,N_1708);
xnor U2377 (N_2377,N_1403,N_2119);
and U2378 (N_2378,N_2053,N_2017);
nand U2379 (N_2379,N_2140,N_2112);
nand U2380 (N_2380,N_1986,N_1849);
or U2381 (N_2381,N_2160,N_1611);
nand U2382 (N_2382,N_2001,N_2079);
or U2383 (N_2383,N_2038,N_2111);
or U2384 (N_2384,N_2052,N_2049);
nor U2385 (N_2385,N_1986,N_2061);
or U2386 (N_2386,In_92,N_2166);
nor U2387 (N_2387,N_2039,N_2021);
or U2388 (N_2388,N_1926,N_2130);
nand U2389 (N_2389,N_1951,N_1194);
or U2390 (N_2390,N_2154,N_2125);
and U2391 (N_2391,N_1936,N_2082);
and U2392 (N_2392,N_2105,In_209);
nand U2393 (N_2393,N_2095,N_1955);
nor U2394 (N_2394,N_2018,N_2041);
or U2395 (N_2395,N_2014,N_1893);
nand U2396 (N_2396,N_2119,N_2162);
nor U2397 (N_2397,N_1890,N_2111);
and U2398 (N_2398,N_2024,N_2118);
or U2399 (N_2399,N_2093,N_2056);
nor U2400 (N_2400,N_2348,N_2206);
or U2401 (N_2401,N_2388,N_2215);
or U2402 (N_2402,N_2383,N_2384);
and U2403 (N_2403,N_2373,N_2213);
and U2404 (N_2404,N_2211,N_2284);
and U2405 (N_2405,N_2238,N_2289);
and U2406 (N_2406,N_2262,N_2293);
or U2407 (N_2407,N_2325,N_2324);
nand U2408 (N_2408,N_2337,N_2263);
or U2409 (N_2409,N_2280,N_2239);
xor U2410 (N_2410,N_2236,N_2386);
and U2411 (N_2411,N_2226,N_2318);
nor U2412 (N_2412,N_2252,N_2269);
or U2413 (N_2413,N_2205,N_2359);
nor U2414 (N_2414,N_2278,N_2303);
or U2415 (N_2415,N_2378,N_2227);
or U2416 (N_2416,N_2264,N_2352);
and U2417 (N_2417,N_2322,N_2217);
nand U2418 (N_2418,N_2312,N_2207);
nor U2419 (N_2419,N_2241,N_2270);
nand U2420 (N_2420,N_2223,N_2328);
or U2421 (N_2421,N_2243,N_2363);
nor U2422 (N_2422,N_2333,N_2274);
nand U2423 (N_2423,N_2345,N_2275);
nand U2424 (N_2424,N_2225,N_2321);
nor U2425 (N_2425,N_2336,N_2355);
nor U2426 (N_2426,N_2240,N_2315);
or U2427 (N_2427,N_2347,N_2221);
nand U2428 (N_2428,N_2201,N_2272);
xor U2429 (N_2429,N_2385,N_2354);
and U2430 (N_2430,N_2212,N_2326);
nand U2431 (N_2431,N_2295,N_2249);
or U2432 (N_2432,N_2271,N_2398);
and U2433 (N_2433,N_2203,N_2380);
nor U2434 (N_2434,N_2297,N_2382);
nor U2435 (N_2435,N_2290,N_2260);
or U2436 (N_2436,N_2389,N_2330);
nor U2437 (N_2437,N_2287,N_2214);
or U2438 (N_2438,N_2381,N_2305);
nand U2439 (N_2439,N_2200,N_2282);
nor U2440 (N_2440,N_2332,N_2370);
and U2441 (N_2441,N_2235,N_2281);
xnor U2442 (N_2442,N_2371,N_2377);
and U2443 (N_2443,N_2334,N_2298);
nor U2444 (N_2444,N_2257,N_2313);
and U2445 (N_2445,N_2360,N_2277);
nor U2446 (N_2446,N_2259,N_2300);
nor U2447 (N_2447,N_2251,N_2361);
and U2448 (N_2448,N_2353,N_2311);
xnor U2449 (N_2449,N_2276,N_2246);
or U2450 (N_2450,N_2283,N_2341);
and U2451 (N_2451,N_2317,N_2390);
or U2452 (N_2452,N_2224,N_2357);
or U2453 (N_2453,N_2301,N_2242);
nor U2454 (N_2454,N_2218,N_2374);
nor U2455 (N_2455,N_2219,N_2306);
nor U2456 (N_2456,N_2208,N_2258);
nor U2457 (N_2457,N_2320,N_2366);
or U2458 (N_2458,N_2299,N_2209);
nand U2459 (N_2459,N_2216,N_2394);
nor U2460 (N_2460,N_2392,N_2395);
nand U2461 (N_2461,N_2229,N_2329);
and U2462 (N_2462,N_2393,N_2253);
nor U2463 (N_2463,N_2350,N_2286);
xor U2464 (N_2464,N_2204,N_2331);
or U2465 (N_2465,N_2247,N_2230);
or U2466 (N_2466,N_2372,N_2376);
and U2467 (N_2467,N_2302,N_2369);
or U2468 (N_2468,N_2340,N_2356);
or U2469 (N_2469,N_2296,N_2244);
or U2470 (N_2470,N_2256,N_2292);
xor U2471 (N_2471,N_2375,N_2358);
nor U2472 (N_2472,N_2291,N_2268);
or U2473 (N_2473,N_2327,N_2387);
nand U2474 (N_2474,N_2362,N_2288);
or U2475 (N_2475,N_2228,N_2265);
and U2476 (N_2476,N_2220,N_2365);
and U2477 (N_2477,N_2319,N_2279);
nand U2478 (N_2478,N_2349,N_2248);
nor U2479 (N_2479,N_2266,N_2346);
nor U2480 (N_2480,N_2367,N_2232);
and U2481 (N_2481,N_2237,N_2285);
xnor U2482 (N_2482,N_2339,N_2379);
and U2483 (N_2483,N_2323,N_2397);
nand U2484 (N_2484,N_2210,N_2308);
and U2485 (N_2485,N_2344,N_2343);
or U2486 (N_2486,N_2316,N_2307);
or U2487 (N_2487,N_2202,N_2255);
nor U2488 (N_2488,N_2233,N_2309);
and U2489 (N_2489,N_2254,N_2391);
nand U2490 (N_2490,N_2222,N_2294);
or U2491 (N_2491,N_2364,N_2335);
and U2492 (N_2492,N_2250,N_2351);
or U2493 (N_2493,N_2267,N_2261);
and U2494 (N_2494,N_2273,N_2245);
nor U2495 (N_2495,N_2310,N_2396);
and U2496 (N_2496,N_2368,N_2304);
and U2497 (N_2497,N_2399,N_2314);
or U2498 (N_2498,N_2338,N_2234);
nand U2499 (N_2499,N_2231,N_2342);
nor U2500 (N_2500,N_2289,N_2355);
or U2501 (N_2501,N_2212,N_2240);
nand U2502 (N_2502,N_2343,N_2328);
xor U2503 (N_2503,N_2228,N_2225);
and U2504 (N_2504,N_2251,N_2299);
and U2505 (N_2505,N_2388,N_2347);
nand U2506 (N_2506,N_2268,N_2318);
xnor U2507 (N_2507,N_2246,N_2216);
nand U2508 (N_2508,N_2256,N_2230);
nand U2509 (N_2509,N_2218,N_2260);
or U2510 (N_2510,N_2250,N_2301);
nor U2511 (N_2511,N_2321,N_2235);
xor U2512 (N_2512,N_2336,N_2283);
nand U2513 (N_2513,N_2258,N_2370);
nand U2514 (N_2514,N_2241,N_2378);
nor U2515 (N_2515,N_2272,N_2302);
and U2516 (N_2516,N_2360,N_2329);
nor U2517 (N_2517,N_2385,N_2222);
and U2518 (N_2518,N_2355,N_2207);
and U2519 (N_2519,N_2288,N_2256);
nand U2520 (N_2520,N_2241,N_2291);
nand U2521 (N_2521,N_2241,N_2342);
nand U2522 (N_2522,N_2373,N_2391);
nor U2523 (N_2523,N_2202,N_2372);
xnor U2524 (N_2524,N_2239,N_2261);
and U2525 (N_2525,N_2360,N_2236);
nand U2526 (N_2526,N_2236,N_2234);
nor U2527 (N_2527,N_2315,N_2228);
or U2528 (N_2528,N_2342,N_2254);
or U2529 (N_2529,N_2339,N_2240);
nand U2530 (N_2530,N_2329,N_2371);
xor U2531 (N_2531,N_2329,N_2298);
nand U2532 (N_2532,N_2325,N_2256);
or U2533 (N_2533,N_2349,N_2226);
nor U2534 (N_2534,N_2344,N_2275);
nand U2535 (N_2535,N_2325,N_2225);
and U2536 (N_2536,N_2314,N_2393);
nand U2537 (N_2537,N_2238,N_2302);
nor U2538 (N_2538,N_2243,N_2296);
nor U2539 (N_2539,N_2263,N_2340);
nor U2540 (N_2540,N_2261,N_2216);
nand U2541 (N_2541,N_2228,N_2226);
and U2542 (N_2542,N_2240,N_2344);
or U2543 (N_2543,N_2266,N_2290);
and U2544 (N_2544,N_2344,N_2390);
nor U2545 (N_2545,N_2376,N_2233);
or U2546 (N_2546,N_2232,N_2271);
nand U2547 (N_2547,N_2208,N_2375);
xor U2548 (N_2548,N_2219,N_2214);
nand U2549 (N_2549,N_2276,N_2368);
nor U2550 (N_2550,N_2330,N_2288);
or U2551 (N_2551,N_2251,N_2366);
or U2552 (N_2552,N_2324,N_2223);
nor U2553 (N_2553,N_2340,N_2280);
nand U2554 (N_2554,N_2295,N_2345);
and U2555 (N_2555,N_2337,N_2313);
and U2556 (N_2556,N_2371,N_2212);
nand U2557 (N_2557,N_2215,N_2327);
xor U2558 (N_2558,N_2278,N_2276);
or U2559 (N_2559,N_2303,N_2394);
xor U2560 (N_2560,N_2363,N_2317);
or U2561 (N_2561,N_2351,N_2356);
and U2562 (N_2562,N_2229,N_2246);
xor U2563 (N_2563,N_2224,N_2365);
or U2564 (N_2564,N_2238,N_2340);
and U2565 (N_2565,N_2212,N_2263);
and U2566 (N_2566,N_2356,N_2365);
and U2567 (N_2567,N_2232,N_2380);
or U2568 (N_2568,N_2230,N_2264);
nor U2569 (N_2569,N_2352,N_2260);
nand U2570 (N_2570,N_2386,N_2240);
or U2571 (N_2571,N_2239,N_2258);
or U2572 (N_2572,N_2320,N_2375);
xor U2573 (N_2573,N_2283,N_2214);
nor U2574 (N_2574,N_2244,N_2222);
or U2575 (N_2575,N_2246,N_2371);
or U2576 (N_2576,N_2289,N_2296);
nand U2577 (N_2577,N_2263,N_2230);
and U2578 (N_2578,N_2213,N_2296);
and U2579 (N_2579,N_2390,N_2293);
and U2580 (N_2580,N_2337,N_2323);
or U2581 (N_2581,N_2371,N_2247);
nand U2582 (N_2582,N_2286,N_2289);
and U2583 (N_2583,N_2269,N_2245);
nor U2584 (N_2584,N_2300,N_2307);
nand U2585 (N_2585,N_2296,N_2260);
and U2586 (N_2586,N_2273,N_2240);
xor U2587 (N_2587,N_2308,N_2200);
or U2588 (N_2588,N_2253,N_2205);
or U2589 (N_2589,N_2280,N_2375);
or U2590 (N_2590,N_2379,N_2216);
nand U2591 (N_2591,N_2372,N_2200);
nor U2592 (N_2592,N_2269,N_2393);
or U2593 (N_2593,N_2287,N_2203);
and U2594 (N_2594,N_2279,N_2259);
and U2595 (N_2595,N_2314,N_2305);
nand U2596 (N_2596,N_2239,N_2234);
nand U2597 (N_2597,N_2345,N_2318);
nor U2598 (N_2598,N_2259,N_2370);
nor U2599 (N_2599,N_2311,N_2369);
or U2600 (N_2600,N_2459,N_2509);
and U2601 (N_2601,N_2420,N_2506);
nor U2602 (N_2602,N_2480,N_2571);
nand U2603 (N_2603,N_2581,N_2537);
and U2604 (N_2604,N_2410,N_2515);
and U2605 (N_2605,N_2496,N_2475);
nand U2606 (N_2606,N_2556,N_2403);
nand U2607 (N_2607,N_2485,N_2598);
and U2608 (N_2608,N_2474,N_2540);
and U2609 (N_2609,N_2406,N_2401);
nor U2610 (N_2610,N_2414,N_2524);
and U2611 (N_2611,N_2586,N_2583);
nor U2612 (N_2612,N_2534,N_2546);
or U2613 (N_2613,N_2542,N_2590);
or U2614 (N_2614,N_2517,N_2466);
nand U2615 (N_2615,N_2487,N_2402);
xnor U2616 (N_2616,N_2400,N_2443);
and U2617 (N_2617,N_2527,N_2483);
xnor U2618 (N_2618,N_2467,N_2428);
nor U2619 (N_2619,N_2561,N_2539);
nand U2620 (N_2620,N_2503,N_2482);
or U2621 (N_2621,N_2407,N_2452);
nand U2622 (N_2622,N_2575,N_2526);
or U2623 (N_2623,N_2456,N_2536);
and U2624 (N_2624,N_2500,N_2419);
or U2625 (N_2625,N_2557,N_2425);
and U2626 (N_2626,N_2469,N_2530);
and U2627 (N_2627,N_2436,N_2566);
or U2628 (N_2628,N_2596,N_2578);
and U2629 (N_2629,N_2593,N_2434);
or U2630 (N_2630,N_2547,N_2535);
nor U2631 (N_2631,N_2440,N_2549);
and U2632 (N_2632,N_2550,N_2471);
nand U2633 (N_2633,N_2455,N_2424);
nand U2634 (N_2634,N_2544,N_2518);
nor U2635 (N_2635,N_2441,N_2555);
nor U2636 (N_2636,N_2577,N_2477);
nor U2637 (N_2637,N_2430,N_2404);
xnor U2638 (N_2638,N_2438,N_2574);
xor U2639 (N_2639,N_2573,N_2418);
or U2640 (N_2640,N_2444,N_2499);
or U2641 (N_2641,N_2568,N_2552);
nand U2642 (N_2642,N_2595,N_2551);
xnor U2643 (N_2643,N_2426,N_2461);
or U2644 (N_2644,N_2457,N_2435);
nor U2645 (N_2645,N_2416,N_2421);
nand U2646 (N_2646,N_2521,N_2522);
or U2647 (N_2647,N_2516,N_2447);
nor U2648 (N_2648,N_2429,N_2431);
and U2649 (N_2649,N_2585,N_2464);
nand U2650 (N_2650,N_2588,N_2560);
nand U2651 (N_2651,N_2520,N_2565);
nor U2652 (N_2652,N_2582,N_2533);
nand U2653 (N_2653,N_2584,N_2576);
or U2654 (N_2654,N_2538,N_2481);
nor U2655 (N_2655,N_2405,N_2514);
nand U2656 (N_2656,N_2413,N_2510);
or U2657 (N_2657,N_2417,N_2580);
nor U2658 (N_2658,N_2587,N_2427);
nor U2659 (N_2659,N_2458,N_2489);
and U2660 (N_2660,N_2529,N_2507);
nand U2661 (N_2661,N_2422,N_2570);
and U2662 (N_2662,N_2599,N_2470);
nor U2663 (N_2663,N_2488,N_2423);
nor U2664 (N_2664,N_2528,N_2553);
xnor U2665 (N_2665,N_2463,N_2572);
nand U2666 (N_2666,N_2504,N_2454);
or U2667 (N_2667,N_2589,N_2502);
or U2668 (N_2668,N_2476,N_2486);
or U2669 (N_2669,N_2493,N_2523);
or U2670 (N_2670,N_2433,N_2408);
and U2671 (N_2671,N_2498,N_2512);
nor U2672 (N_2672,N_2548,N_2472);
and U2673 (N_2673,N_2450,N_2451);
nor U2674 (N_2674,N_2591,N_2564);
and U2675 (N_2675,N_2569,N_2460);
or U2676 (N_2676,N_2409,N_2473);
and U2677 (N_2677,N_2567,N_2543);
nor U2678 (N_2678,N_2453,N_2479);
nand U2679 (N_2679,N_2491,N_2531);
nand U2680 (N_2680,N_2462,N_2592);
or U2681 (N_2681,N_2594,N_2446);
nor U2682 (N_2682,N_2559,N_2508);
and U2683 (N_2683,N_2497,N_2468);
and U2684 (N_2684,N_2545,N_2484);
nor U2685 (N_2685,N_2412,N_2439);
and U2686 (N_2686,N_2442,N_2541);
and U2687 (N_2687,N_2554,N_2445);
or U2688 (N_2688,N_2558,N_2511);
nor U2689 (N_2689,N_2448,N_2501);
and U2690 (N_2690,N_2432,N_2494);
nand U2691 (N_2691,N_2597,N_2579);
nand U2692 (N_2692,N_2415,N_2513);
nor U2693 (N_2693,N_2449,N_2490);
and U2694 (N_2694,N_2411,N_2519);
and U2695 (N_2695,N_2532,N_2492);
nor U2696 (N_2696,N_2505,N_2562);
and U2697 (N_2697,N_2437,N_2465);
or U2698 (N_2698,N_2563,N_2478);
nand U2699 (N_2699,N_2525,N_2495);
xor U2700 (N_2700,N_2498,N_2542);
or U2701 (N_2701,N_2410,N_2557);
nor U2702 (N_2702,N_2449,N_2511);
or U2703 (N_2703,N_2451,N_2556);
and U2704 (N_2704,N_2494,N_2503);
and U2705 (N_2705,N_2541,N_2502);
or U2706 (N_2706,N_2406,N_2435);
or U2707 (N_2707,N_2479,N_2412);
nor U2708 (N_2708,N_2406,N_2492);
and U2709 (N_2709,N_2450,N_2483);
and U2710 (N_2710,N_2556,N_2562);
or U2711 (N_2711,N_2518,N_2547);
and U2712 (N_2712,N_2494,N_2580);
or U2713 (N_2713,N_2472,N_2540);
and U2714 (N_2714,N_2585,N_2443);
nand U2715 (N_2715,N_2537,N_2499);
and U2716 (N_2716,N_2548,N_2560);
or U2717 (N_2717,N_2469,N_2453);
and U2718 (N_2718,N_2448,N_2464);
and U2719 (N_2719,N_2537,N_2543);
or U2720 (N_2720,N_2540,N_2432);
and U2721 (N_2721,N_2464,N_2444);
or U2722 (N_2722,N_2422,N_2504);
or U2723 (N_2723,N_2435,N_2550);
or U2724 (N_2724,N_2456,N_2500);
nor U2725 (N_2725,N_2489,N_2578);
nand U2726 (N_2726,N_2531,N_2562);
or U2727 (N_2727,N_2578,N_2577);
xor U2728 (N_2728,N_2460,N_2415);
nor U2729 (N_2729,N_2464,N_2452);
and U2730 (N_2730,N_2531,N_2417);
or U2731 (N_2731,N_2593,N_2455);
or U2732 (N_2732,N_2462,N_2568);
nor U2733 (N_2733,N_2433,N_2463);
nand U2734 (N_2734,N_2581,N_2450);
nand U2735 (N_2735,N_2549,N_2476);
and U2736 (N_2736,N_2585,N_2545);
nor U2737 (N_2737,N_2456,N_2426);
or U2738 (N_2738,N_2418,N_2441);
and U2739 (N_2739,N_2494,N_2452);
nor U2740 (N_2740,N_2415,N_2456);
nand U2741 (N_2741,N_2431,N_2421);
and U2742 (N_2742,N_2447,N_2540);
nor U2743 (N_2743,N_2439,N_2415);
nand U2744 (N_2744,N_2503,N_2421);
or U2745 (N_2745,N_2529,N_2453);
or U2746 (N_2746,N_2488,N_2592);
or U2747 (N_2747,N_2579,N_2560);
or U2748 (N_2748,N_2479,N_2428);
nor U2749 (N_2749,N_2459,N_2497);
nor U2750 (N_2750,N_2579,N_2575);
nand U2751 (N_2751,N_2587,N_2424);
xor U2752 (N_2752,N_2506,N_2498);
nand U2753 (N_2753,N_2516,N_2483);
and U2754 (N_2754,N_2596,N_2448);
or U2755 (N_2755,N_2448,N_2520);
or U2756 (N_2756,N_2561,N_2469);
nand U2757 (N_2757,N_2535,N_2514);
nand U2758 (N_2758,N_2414,N_2480);
nand U2759 (N_2759,N_2587,N_2543);
nor U2760 (N_2760,N_2566,N_2403);
and U2761 (N_2761,N_2578,N_2400);
nand U2762 (N_2762,N_2584,N_2513);
nor U2763 (N_2763,N_2401,N_2557);
or U2764 (N_2764,N_2564,N_2471);
or U2765 (N_2765,N_2572,N_2566);
nor U2766 (N_2766,N_2590,N_2440);
nor U2767 (N_2767,N_2512,N_2409);
nand U2768 (N_2768,N_2563,N_2476);
and U2769 (N_2769,N_2469,N_2433);
and U2770 (N_2770,N_2517,N_2484);
and U2771 (N_2771,N_2524,N_2540);
xor U2772 (N_2772,N_2485,N_2592);
or U2773 (N_2773,N_2453,N_2527);
xnor U2774 (N_2774,N_2475,N_2542);
nor U2775 (N_2775,N_2523,N_2490);
nand U2776 (N_2776,N_2406,N_2437);
xnor U2777 (N_2777,N_2431,N_2430);
and U2778 (N_2778,N_2437,N_2548);
xnor U2779 (N_2779,N_2415,N_2405);
nand U2780 (N_2780,N_2465,N_2523);
and U2781 (N_2781,N_2534,N_2526);
nand U2782 (N_2782,N_2410,N_2486);
nand U2783 (N_2783,N_2533,N_2545);
and U2784 (N_2784,N_2457,N_2505);
and U2785 (N_2785,N_2588,N_2525);
nand U2786 (N_2786,N_2509,N_2448);
or U2787 (N_2787,N_2478,N_2572);
and U2788 (N_2788,N_2455,N_2571);
nor U2789 (N_2789,N_2475,N_2546);
and U2790 (N_2790,N_2463,N_2413);
or U2791 (N_2791,N_2422,N_2574);
nor U2792 (N_2792,N_2460,N_2479);
and U2793 (N_2793,N_2468,N_2490);
and U2794 (N_2794,N_2466,N_2412);
and U2795 (N_2795,N_2433,N_2410);
or U2796 (N_2796,N_2471,N_2510);
or U2797 (N_2797,N_2413,N_2498);
nor U2798 (N_2798,N_2559,N_2495);
xor U2799 (N_2799,N_2423,N_2458);
nor U2800 (N_2800,N_2779,N_2649);
or U2801 (N_2801,N_2747,N_2703);
nand U2802 (N_2802,N_2627,N_2794);
nand U2803 (N_2803,N_2647,N_2764);
nand U2804 (N_2804,N_2695,N_2752);
nor U2805 (N_2805,N_2610,N_2772);
or U2806 (N_2806,N_2698,N_2663);
and U2807 (N_2807,N_2670,N_2688);
nor U2808 (N_2808,N_2659,N_2727);
and U2809 (N_2809,N_2740,N_2619);
xor U2810 (N_2810,N_2682,N_2611);
or U2811 (N_2811,N_2662,N_2768);
or U2812 (N_2812,N_2656,N_2783);
nand U2813 (N_2813,N_2701,N_2687);
or U2814 (N_2814,N_2660,N_2765);
and U2815 (N_2815,N_2689,N_2672);
nand U2816 (N_2816,N_2654,N_2648);
and U2817 (N_2817,N_2645,N_2677);
or U2818 (N_2818,N_2722,N_2616);
nand U2819 (N_2819,N_2710,N_2679);
nor U2820 (N_2820,N_2774,N_2756);
and U2821 (N_2821,N_2751,N_2725);
and U2822 (N_2822,N_2739,N_2726);
nor U2823 (N_2823,N_2719,N_2704);
nand U2824 (N_2824,N_2615,N_2644);
nand U2825 (N_2825,N_2736,N_2799);
nand U2826 (N_2826,N_2788,N_2620);
or U2827 (N_2827,N_2781,N_2797);
nor U2828 (N_2828,N_2762,N_2652);
and U2829 (N_2829,N_2641,N_2604);
nand U2830 (N_2830,N_2600,N_2785);
xor U2831 (N_2831,N_2617,N_2691);
and U2832 (N_2832,N_2778,N_2700);
nor U2833 (N_2833,N_2653,N_2712);
nand U2834 (N_2834,N_2786,N_2743);
and U2835 (N_2835,N_2667,N_2643);
nor U2836 (N_2836,N_2618,N_2798);
nand U2837 (N_2837,N_2613,N_2602);
or U2838 (N_2838,N_2761,N_2685);
xnor U2839 (N_2839,N_2792,N_2748);
nand U2840 (N_2840,N_2746,N_2637);
nor U2841 (N_2841,N_2657,N_2603);
nand U2842 (N_2842,N_2668,N_2721);
or U2843 (N_2843,N_2767,N_2763);
nor U2844 (N_2844,N_2623,N_2773);
nor U2845 (N_2845,N_2639,N_2735);
nor U2846 (N_2846,N_2650,N_2718);
or U2847 (N_2847,N_2661,N_2614);
and U2848 (N_2848,N_2741,N_2715);
and U2849 (N_2849,N_2694,N_2753);
or U2850 (N_2850,N_2629,N_2717);
xor U2851 (N_2851,N_2633,N_2699);
nor U2852 (N_2852,N_2665,N_2771);
nor U2853 (N_2853,N_2642,N_2666);
and U2854 (N_2854,N_2766,N_2730);
or U2855 (N_2855,N_2626,N_2608);
xnor U2856 (N_2856,N_2632,N_2723);
nand U2857 (N_2857,N_2795,N_2758);
nor U2858 (N_2858,N_2790,N_2733);
and U2859 (N_2859,N_2729,N_2707);
nand U2860 (N_2860,N_2775,N_2759);
or U2861 (N_2861,N_2731,N_2709);
or U2862 (N_2862,N_2681,N_2651);
nand U2863 (N_2863,N_2744,N_2606);
xnor U2864 (N_2864,N_2605,N_2636);
nor U2865 (N_2865,N_2655,N_2675);
or U2866 (N_2866,N_2769,N_2624);
nand U2867 (N_2867,N_2673,N_2686);
nor U2868 (N_2868,N_2658,N_2676);
or U2869 (N_2869,N_2671,N_2714);
and U2870 (N_2870,N_2776,N_2630);
nor U2871 (N_2871,N_2755,N_2702);
nor U2872 (N_2872,N_2749,N_2684);
xor U2873 (N_2873,N_2622,N_2669);
or U2874 (N_2874,N_2745,N_2780);
nor U2875 (N_2875,N_2734,N_2732);
and U2876 (N_2876,N_2696,N_2628);
xnor U2877 (N_2877,N_2697,N_2760);
nor U2878 (N_2878,N_2713,N_2612);
and U2879 (N_2879,N_2724,N_2625);
xnor U2880 (N_2880,N_2738,N_2787);
nand U2881 (N_2881,N_2757,N_2678);
and U2882 (N_2882,N_2601,N_2737);
or U2883 (N_2883,N_2607,N_2742);
or U2884 (N_2884,N_2664,N_2634);
and U2885 (N_2885,N_2711,N_2789);
nand U2886 (N_2886,N_2690,N_2692);
nor U2887 (N_2887,N_2706,N_2770);
and U2888 (N_2888,N_2683,N_2750);
and U2889 (N_2889,N_2708,N_2728);
and U2890 (N_2890,N_2784,N_2674);
and U2891 (N_2891,N_2777,N_2621);
or U2892 (N_2892,N_2680,N_2609);
or U2893 (N_2893,N_2791,N_2693);
and U2894 (N_2894,N_2796,N_2631);
xnor U2895 (N_2895,N_2638,N_2705);
and U2896 (N_2896,N_2646,N_2716);
nor U2897 (N_2897,N_2782,N_2793);
and U2898 (N_2898,N_2640,N_2754);
xor U2899 (N_2899,N_2720,N_2635);
nand U2900 (N_2900,N_2661,N_2655);
nand U2901 (N_2901,N_2640,N_2724);
or U2902 (N_2902,N_2675,N_2694);
or U2903 (N_2903,N_2710,N_2705);
and U2904 (N_2904,N_2769,N_2793);
nor U2905 (N_2905,N_2718,N_2625);
or U2906 (N_2906,N_2683,N_2688);
or U2907 (N_2907,N_2650,N_2708);
or U2908 (N_2908,N_2747,N_2632);
xor U2909 (N_2909,N_2746,N_2723);
and U2910 (N_2910,N_2670,N_2728);
nor U2911 (N_2911,N_2703,N_2687);
or U2912 (N_2912,N_2623,N_2657);
nor U2913 (N_2913,N_2718,N_2677);
and U2914 (N_2914,N_2698,N_2651);
nor U2915 (N_2915,N_2705,N_2733);
xnor U2916 (N_2916,N_2668,N_2687);
or U2917 (N_2917,N_2680,N_2706);
or U2918 (N_2918,N_2613,N_2745);
nor U2919 (N_2919,N_2624,N_2717);
nand U2920 (N_2920,N_2639,N_2734);
nand U2921 (N_2921,N_2750,N_2691);
or U2922 (N_2922,N_2637,N_2751);
or U2923 (N_2923,N_2690,N_2712);
nor U2924 (N_2924,N_2714,N_2794);
or U2925 (N_2925,N_2747,N_2668);
nand U2926 (N_2926,N_2603,N_2757);
nand U2927 (N_2927,N_2717,N_2647);
nor U2928 (N_2928,N_2633,N_2605);
nand U2929 (N_2929,N_2665,N_2680);
nor U2930 (N_2930,N_2717,N_2618);
nor U2931 (N_2931,N_2654,N_2667);
nand U2932 (N_2932,N_2661,N_2606);
nor U2933 (N_2933,N_2603,N_2742);
and U2934 (N_2934,N_2722,N_2739);
xnor U2935 (N_2935,N_2744,N_2675);
or U2936 (N_2936,N_2606,N_2698);
nor U2937 (N_2937,N_2618,N_2752);
xnor U2938 (N_2938,N_2636,N_2609);
or U2939 (N_2939,N_2644,N_2713);
nor U2940 (N_2940,N_2630,N_2704);
nand U2941 (N_2941,N_2738,N_2764);
nor U2942 (N_2942,N_2622,N_2659);
nand U2943 (N_2943,N_2744,N_2706);
nor U2944 (N_2944,N_2660,N_2795);
xnor U2945 (N_2945,N_2704,N_2603);
nor U2946 (N_2946,N_2606,N_2618);
nor U2947 (N_2947,N_2647,N_2631);
nor U2948 (N_2948,N_2771,N_2637);
nor U2949 (N_2949,N_2780,N_2663);
nor U2950 (N_2950,N_2766,N_2726);
and U2951 (N_2951,N_2612,N_2655);
and U2952 (N_2952,N_2718,N_2651);
nand U2953 (N_2953,N_2783,N_2613);
and U2954 (N_2954,N_2601,N_2703);
and U2955 (N_2955,N_2661,N_2680);
nand U2956 (N_2956,N_2681,N_2684);
nor U2957 (N_2957,N_2603,N_2666);
nand U2958 (N_2958,N_2700,N_2617);
and U2959 (N_2959,N_2681,N_2704);
nand U2960 (N_2960,N_2629,N_2723);
and U2961 (N_2961,N_2701,N_2648);
nor U2962 (N_2962,N_2711,N_2791);
or U2963 (N_2963,N_2746,N_2662);
and U2964 (N_2964,N_2715,N_2777);
and U2965 (N_2965,N_2747,N_2749);
and U2966 (N_2966,N_2657,N_2695);
and U2967 (N_2967,N_2748,N_2656);
nor U2968 (N_2968,N_2601,N_2794);
and U2969 (N_2969,N_2712,N_2604);
or U2970 (N_2970,N_2789,N_2716);
nor U2971 (N_2971,N_2664,N_2763);
xor U2972 (N_2972,N_2621,N_2760);
or U2973 (N_2973,N_2796,N_2688);
and U2974 (N_2974,N_2738,N_2697);
or U2975 (N_2975,N_2727,N_2769);
nand U2976 (N_2976,N_2705,N_2676);
nor U2977 (N_2977,N_2650,N_2660);
nor U2978 (N_2978,N_2601,N_2702);
nand U2979 (N_2979,N_2763,N_2607);
and U2980 (N_2980,N_2696,N_2782);
nand U2981 (N_2981,N_2626,N_2621);
and U2982 (N_2982,N_2698,N_2773);
nor U2983 (N_2983,N_2758,N_2751);
or U2984 (N_2984,N_2608,N_2767);
and U2985 (N_2985,N_2764,N_2662);
and U2986 (N_2986,N_2743,N_2775);
nand U2987 (N_2987,N_2739,N_2631);
or U2988 (N_2988,N_2773,N_2654);
xnor U2989 (N_2989,N_2631,N_2794);
and U2990 (N_2990,N_2746,N_2786);
or U2991 (N_2991,N_2719,N_2738);
or U2992 (N_2992,N_2671,N_2675);
xor U2993 (N_2993,N_2693,N_2612);
nand U2994 (N_2994,N_2719,N_2660);
nor U2995 (N_2995,N_2623,N_2751);
or U2996 (N_2996,N_2745,N_2712);
nand U2997 (N_2997,N_2747,N_2702);
nor U2998 (N_2998,N_2661,N_2659);
nand U2999 (N_2999,N_2612,N_2601);
and U3000 (N_3000,N_2888,N_2989);
and U3001 (N_3001,N_2961,N_2834);
and U3002 (N_3002,N_2860,N_2921);
nand U3003 (N_3003,N_2873,N_2844);
nor U3004 (N_3004,N_2970,N_2805);
nand U3005 (N_3005,N_2952,N_2818);
and U3006 (N_3006,N_2946,N_2942);
nand U3007 (N_3007,N_2838,N_2847);
nor U3008 (N_3008,N_2897,N_2924);
and U3009 (N_3009,N_2950,N_2922);
nor U3010 (N_3010,N_2831,N_2850);
nor U3011 (N_3011,N_2899,N_2857);
nor U3012 (N_3012,N_2965,N_2863);
and U3013 (N_3013,N_2839,N_2926);
nor U3014 (N_3014,N_2959,N_2992);
or U3015 (N_3015,N_2865,N_2994);
or U3016 (N_3016,N_2905,N_2813);
and U3017 (N_3017,N_2914,N_2830);
and U3018 (N_3018,N_2896,N_2918);
and U3019 (N_3019,N_2855,N_2967);
nand U3020 (N_3020,N_2803,N_2884);
or U3021 (N_3021,N_2953,N_2824);
nand U3022 (N_3022,N_2990,N_2912);
or U3023 (N_3023,N_2960,N_2939);
nor U3024 (N_3024,N_2971,N_2815);
nand U3025 (N_3025,N_2890,N_2816);
or U3026 (N_3026,N_2987,N_2991);
or U3027 (N_3027,N_2957,N_2973);
or U3028 (N_3028,N_2804,N_2846);
nand U3029 (N_3029,N_2995,N_2882);
or U3030 (N_3030,N_2972,N_2949);
nand U3031 (N_3031,N_2820,N_2903);
xnor U3032 (N_3032,N_2880,N_2917);
and U3033 (N_3033,N_2907,N_2968);
nand U3034 (N_3034,N_2821,N_2809);
nand U3035 (N_3035,N_2858,N_2974);
and U3036 (N_3036,N_2872,N_2893);
or U3037 (N_3037,N_2931,N_2900);
nor U3038 (N_3038,N_2866,N_2828);
nor U3039 (N_3039,N_2827,N_2996);
or U3040 (N_3040,N_2822,N_2867);
and U3041 (N_3041,N_2848,N_2840);
nor U3042 (N_3042,N_2930,N_2909);
nor U3043 (N_3043,N_2812,N_2997);
or U3044 (N_3044,N_2927,N_2800);
nor U3045 (N_3045,N_2913,N_2911);
or U3046 (N_3046,N_2883,N_2871);
or U3047 (N_3047,N_2856,N_2978);
nand U3048 (N_3048,N_2817,N_2843);
xnor U3049 (N_3049,N_2842,N_2869);
xor U3050 (N_3050,N_2947,N_2977);
nor U3051 (N_3051,N_2937,N_2979);
or U3052 (N_3052,N_2943,N_2825);
and U3053 (N_3053,N_2928,N_2886);
nand U3054 (N_3054,N_2932,N_2934);
and U3055 (N_3055,N_2808,N_2864);
nor U3056 (N_3056,N_2823,N_2810);
nor U3057 (N_3057,N_2845,N_2879);
nand U3058 (N_3058,N_2938,N_2983);
nor U3059 (N_3059,N_2854,N_2923);
and U3060 (N_3060,N_2876,N_2841);
nor U3061 (N_3061,N_2870,N_2852);
or U3062 (N_3062,N_2981,N_2906);
or U3063 (N_3063,N_2963,N_2925);
nand U3064 (N_3064,N_2941,N_2862);
or U3065 (N_3065,N_2853,N_2908);
and U3066 (N_3066,N_2984,N_2811);
nor U3067 (N_3067,N_2806,N_2975);
or U3068 (N_3068,N_2875,N_2935);
or U3069 (N_3069,N_2948,N_2904);
or U3070 (N_3070,N_2802,N_2920);
nor U3071 (N_3071,N_2887,N_2895);
nor U3072 (N_3072,N_2982,N_2929);
or U3073 (N_3073,N_2944,N_2998);
nand U3074 (N_3074,N_2851,N_2801);
nand U3075 (N_3075,N_2964,N_2829);
and U3076 (N_3076,N_2919,N_2892);
or U3077 (N_3077,N_2878,N_2894);
nand U3078 (N_3078,N_2962,N_2826);
nor U3079 (N_3079,N_2993,N_2915);
nor U3080 (N_3080,N_2901,N_2945);
nand U3081 (N_3081,N_2954,N_2966);
nor U3082 (N_3082,N_2837,N_2902);
nor U3083 (N_3083,N_2976,N_2849);
nand U3084 (N_3084,N_2885,N_2814);
and U3085 (N_3085,N_2940,N_2980);
or U3086 (N_3086,N_2936,N_2951);
nand U3087 (N_3087,N_2999,N_2889);
and U3088 (N_3088,N_2868,N_2988);
nand U3089 (N_3089,N_2859,N_2836);
and U3090 (N_3090,N_2874,N_2832);
xor U3091 (N_3091,N_2881,N_2916);
nor U3092 (N_3092,N_2956,N_2819);
xnor U3093 (N_3093,N_2986,N_2861);
xor U3094 (N_3094,N_2898,N_2891);
or U3095 (N_3095,N_2985,N_2877);
or U3096 (N_3096,N_2833,N_2910);
and U3097 (N_3097,N_2807,N_2958);
nand U3098 (N_3098,N_2969,N_2835);
nand U3099 (N_3099,N_2955,N_2933);
and U3100 (N_3100,N_2994,N_2947);
nand U3101 (N_3101,N_2820,N_2963);
nand U3102 (N_3102,N_2873,N_2935);
nor U3103 (N_3103,N_2845,N_2823);
or U3104 (N_3104,N_2920,N_2822);
nor U3105 (N_3105,N_2886,N_2984);
nor U3106 (N_3106,N_2851,N_2926);
nand U3107 (N_3107,N_2875,N_2821);
nor U3108 (N_3108,N_2943,N_2967);
or U3109 (N_3109,N_2913,N_2853);
nor U3110 (N_3110,N_2953,N_2863);
nor U3111 (N_3111,N_2819,N_2995);
nor U3112 (N_3112,N_2932,N_2945);
nand U3113 (N_3113,N_2955,N_2942);
nor U3114 (N_3114,N_2817,N_2969);
nand U3115 (N_3115,N_2885,N_2949);
and U3116 (N_3116,N_2807,N_2968);
nor U3117 (N_3117,N_2871,N_2844);
xnor U3118 (N_3118,N_2816,N_2995);
nand U3119 (N_3119,N_2921,N_2818);
and U3120 (N_3120,N_2854,N_2876);
or U3121 (N_3121,N_2802,N_2896);
nand U3122 (N_3122,N_2978,N_2984);
nand U3123 (N_3123,N_2806,N_2879);
xnor U3124 (N_3124,N_2872,N_2953);
or U3125 (N_3125,N_2818,N_2856);
nand U3126 (N_3126,N_2920,N_2927);
and U3127 (N_3127,N_2831,N_2878);
nand U3128 (N_3128,N_2937,N_2987);
nor U3129 (N_3129,N_2852,N_2807);
nand U3130 (N_3130,N_2837,N_2975);
xor U3131 (N_3131,N_2924,N_2808);
and U3132 (N_3132,N_2928,N_2973);
xor U3133 (N_3133,N_2893,N_2913);
xor U3134 (N_3134,N_2918,N_2825);
nor U3135 (N_3135,N_2956,N_2900);
nor U3136 (N_3136,N_2825,N_2957);
xor U3137 (N_3137,N_2950,N_2824);
nand U3138 (N_3138,N_2899,N_2846);
or U3139 (N_3139,N_2965,N_2918);
nor U3140 (N_3140,N_2910,N_2816);
nor U3141 (N_3141,N_2871,N_2979);
nand U3142 (N_3142,N_2994,N_2835);
nand U3143 (N_3143,N_2870,N_2835);
or U3144 (N_3144,N_2913,N_2816);
nor U3145 (N_3145,N_2813,N_2806);
nand U3146 (N_3146,N_2821,N_2876);
and U3147 (N_3147,N_2993,N_2821);
nor U3148 (N_3148,N_2866,N_2991);
nor U3149 (N_3149,N_2953,N_2986);
nor U3150 (N_3150,N_2850,N_2834);
and U3151 (N_3151,N_2914,N_2989);
or U3152 (N_3152,N_2878,N_2935);
nor U3153 (N_3153,N_2996,N_2994);
and U3154 (N_3154,N_2900,N_2842);
nor U3155 (N_3155,N_2846,N_2867);
nand U3156 (N_3156,N_2862,N_2828);
and U3157 (N_3157,N_2803,N_2988);
nor U3158 (N_3158,N_2958,N_2911);
nand U3159 (N_3159,N_2806,N_2905);
xor U3160 (N_3160,N_2878,N_2919);
nand U3161 (N_3161,N_2999,N_2925);
nor U3162 (N_3162,N_2821,N_2802);
nand U3163 (N_3163,N_2870,N_2972);
and U3164 (N_3164,N_2832,N_2916);
xnor U3165 (N_3165,N_2819,N_2887);
or U3166 (N_3166,N_2930,N_2883);
nor U3167 (N_3167,N_2950,N_2895);
xnor U3168 (N_3168,N_2924,N_2910);
xnor U3169 (N_3169,N_2992,N_2822);
and U3170 (N_3170,N_2915,N_2959);
nand U3171 (N_3171,N_2836,N_2861);
nor U3172 (N_3172,N_2999,N_2975);
or U3173 (N_3173,N_2868,N_2878);
xor U3174 (N_3174,N_2864,N_2944);
nand U3175 (N_3175,N_2861,N_2940);
nand U3176 (N_3176,N_2936,N_2836);
nand U3177 (N_3177,N_2998,N_2871);
xor U3178 (N_3178,N_2981,N_2949);
nor U3179 (N_3179,N_2847,N_2998);
nor U3180 (N_3180,N_2922,N_2989);
nand U3181 (N_3181,N_2929,N_2946);
and U3182 (N_3182,N_2850,N_2966);
nor U3183 (N_3183,N_2993,N_2989);
nor U3184 (N_3184,N_2990,N_2812);
xnor U3185 (N_3185,N_2852,N_2872);
xor U3186 (N_3186,N_2870,N_2906);
nor U3187 (N_3187,N_2997,N_2888);
or U3188 (N_3188,N_2983,N_2987);
or U3189 (N_3189,N_2915,N_2811);
and U3190 (N_3190,N_2918,N_2800);
and U3191 (N_3191,N_2842,N_2942);
or U3192 (N_3192,N_2812,N_2819);
nand U3193 (N_3193,N_2908,N_2803);
or U3194 (N_3194,N_2966,N_2880);
nand U3195 (N_3195,N_2979,N_2853);
nor U3196 (N_3196,N_2896,N_2813);
or U3197 (N_3197,N_2822,N_2811);
nor U3198 (N_3198,N_2977,N_2907);
nand U3199 (N_3199,N_2955,N_2801);
or U3200 (N_3200,N_3002,N_3004);
xor U3201 (N_3201,N_3006,N_3097);
nor U3202 (N_3202,N_3136,N_3089);
nor U3203 (N_3203,N_3079,N_3194);
or U3204 (N_3204,N_3174,N_3100);
and U3205 (N_3205,N_3177,N_3092);
nor U3206 (N_3206,N_3150,N_3042);
nand U3207 (N_3207,N_3055,N_3101);
nor U3208 (N_3208,N_3070,N_3170);
and U3209 (N_3209,N_3126,N_3140);
nand U3210 (N_3210,N_3062,N_3096);
nor U3211 (N_3211,N_3109,N_3088);
and U3212 (N_3212,N_3020,N_3027);
and U3213 (N_3213,N_3039,N_3017);
or U3214 (N_3214,N_3036,N_3037);
nand U3215 (N_3215,N_3035,N_3024);
xnor U3216 (N_3216,N_3044,N_3168);
nor U3217 (N_3217,N_3111,N_3154);
or U3218 (N_3218,N_3198,N_3139);
and U3219 (N_3219,N_3135,N_3009);
nand U3220 (N_3220,N_3078,N_3125);
nor U3221 (N_3221,N_3180,N_3143);
nand U3222 (N_3222,N_3137,N_3183);
or U3223 (N_3223,N_3115,N_3158);
and U3224 (N_3224,N_3189,N_3118);
nor U3225 (N_3225,N_3152,N_3195);
nand U3226 (N_3226,N_3072,N_3049);
nand U3227 (N_3227,N_3019,N_3094);
and U3228 (N_3228,N_3040,N_3102);
nand U3229 (N_3229,N_3075,N_3095);
and U3230 (N_3230,N_3169,N_3171);
and U3231 (N_3231,N_3054,N_3138);
nand U3232 (N_3232,N_3149,N_3110);
nor U3233 (N_3233,N_3005,N_3160);
nand U3234 (N_3234,N_3016,N_3184);
and U3235 (N_3235,N_3112,N_3058);
or U3236 (N_3236,N_3010,N_3098);
nor U3237 (N_3237,N_3012,N_3071);
or U3238 (N_3238,N_3166,N_3175);
or U3239 (N_3239,N_3033,N_3046);
and U3240 (N_3240,N_3060,N_3013);
nand U3241 (N_3241,N_3099,N_3031);
nand U3242 (N_3242,N_3133,N_3032);
nor U3243 (N_3243,N_3091,N_3197);
and U3244 (N_3244,N_3162,N_3146);
and U3245 (N_3245,N_3129,N_3053);
nor U3246 (N_3246,N_3068,N_3122);
and U3247 (N_3247,N_3090,N_3030);
nor U3248 (N_3248,N_3083,N_3085);
nand U3249 (N_3249,N_3043,N_3144);
xor U3250 (N_3250,N_3116,N_3008);
nand U3251 (N_3251,N_3186,N_3153);
nand U3252 (N_3252,N_3185,N_3131);
and U3253 (N_3253,N_3107,N_3081);
and U3254 (N_3254,N_3124,N_3157);
and U3255 (N_3255,N_3018,N_3014);
nand U3256 (N_3256,N_3034,N_3196);
and U3257 (N_3257,N_3045,N_3121);
nor U3258 (N_3258,N_3191,N_3038);
nand U3259 (N_3259,N_3134,N_3007);
nand U3260 (N_3260,N_3172,N_3155);
and U3261 (N_3261,N_3050,N_3128);
and U3262 (N_3262,N_3173,N_3114);
or U3263 (N_3263,N_3182,N_3056);
nand U3264 (N_3264,N_3059,N_3087);
and U3265 (N_3265,N_3145,N_3052);
nand U3266 (N_3266,N_3190,N_3080);
and U3267 (N_3267,N_3179,N_3086);
xor U3268 (N_3268,N_3077,N_3147);
and U3269 (N_3269,N_3067,N_3061);
xor U3270 (N_3270,N_3103,N_3064);
nor U3271 (N_3271,N_3015,N_3181);
nor U3272 (N_3272,N_3199,N_3066);
xnor U3273 (N_3273,N_3132,N_3151);
and U3274 (N_3274,N_3119,N_3193);
or U3275 (N_3275,N_3021,N_3120);
or U3276 (N_3276,N_3001,N_3141);
and U3277 (N_3277,N_3192,N_3084);
nand U3278 (N_3278,N_3106,N_3093);
and U3279 (N_3279,N_3029,N_3127);
or U3280 (N_3280,N_3022,N_3167);
or U3281 (N_3281,N_3113,N_3026);
and U3282 (N_3282,N_3117,N_3076);
and U3283 (N_3283,N_3011,N_3065);
or U3284 (N_3284,N_3047,N_3057);
xnor U3285 (N_3285,N_3074,N_3025);
nand U3286 (N_3286,N_3000,N_3130);
and U3287 (N_3287,N_3063,N_3163);
nor U3288 (N_3288,N_3073,N_3142);
nand U3289 (N_3289,N_3178,N_3108);
xnor U3290 (N_3290,N_3048,N_3159);
nand U3291 (N_3291,N_3069,N_3164);
and U3292 (N_3292,N_3104,N_3161);
nor U3293 (N_3293,N_3188,N_3187);
and U3294 (N_3294,N_3028,N_3148);
or U3295 (N_3295,N_3023,N_3051);
nor U3296 (N_3296,N_3105,N_3082);
nor U3297 (N_3297,N_3156,N_3003);
nor U3298 (N_3298,N_3176,N_3123);
and U3299 (N_3299,N_3041,N_3165);
nand U3300 (N_3300,N_3139,N_3096);
or U3301 (N_3301,N_3150,N_3114);
nor U3302 (N_3302,N_3056,N_3064);
nand U3303 (N_3303,N_3099,N_3135);
or U3304 (N_3304,N_3032,N_3017);
and U3305 (N_3305,N_3068,N_3075);
nor U3306 (N_3306,N_3011,N_3088);
nand U3307 (N_3307,N_3010,N_3115);
xnor U3308 (N_3308,N_3157,N_3135);
nand U3309 (N_3309,N_3073,N_3017);
nor U3310 (N_3310,N_3102,N_3184);
nor U3311 (N_3311,N_3081,N_3044);
xor U3312 (N_3312,N_3160,N_3190);
and U3313 (N_3313,N_3052,N_3014);
and U3314 (N_3314,N_3011,N_3155);
nor U3315 (N_3315,N_3163,N_3152);
and U3316 (N_3316,N_3095,N_3006);
or U3317 (N_3317,N_3030,N_3021);
nand U3318 (N_3318,N_3071,N_3101);
or U3319 (N_3319,N_3126,N_3037);
and U3320 (N_3320,N_3096,N_3074);
or U3321 (N_3321,N_3169,N_3181);
nand U3322 (N_3322,N_3054,N_3014);
or U3323 (N_3323,N_3142,N_3054);
or U3324 (N_3324,N_3122,N_3196);
and U3325 (N_3325,N_3114,N_3052);
or U3326 (N_3326,N_3178,N_3165);
or U3327 (N_3327,N_3028,N_3155);
nand U3328 (N_3328,N_3169,N_3113);
and U3329 (N_3329,N_3163,N_3118);
or U3330 (N_3330,N_3048,N_3035);
xnor U3331 (N_3331,N_3176,N_3106);
nor U3332 (N_3332,N_3156,N_3166);
and U3333 (N_3333,N_3104,N_3138);
or U3334 (N_3334,N_3142,N_3139);
nand U3335 (N_3335,N_3184,N_3124);
or U3336 (N_3336,N_3151,N_3180);
nand U3337 (N_3337,N_3165,N_3104);
nor U3338 (N_3338,N_3183,N_3003);
or U3339 (N_3339,N_3048,N_3156);
or U3340 (N_3340,N_3063,N_3198);
nor U3341 (N_3341,N_3169,N_3098);
nand U3342 (N_3342,N_3162,N_3001);
and U3343 (N_3343,N_3085,N_3136);
and U3344 (N_3344,N_3042,N_3065);
xor U3345 (N_3345,N_3055,N_3007);
and U3346 (N_3346,N_3111,N_3167);
nor U3347 (N_3347,N_3103,N_3131);
and U3348 (N_3348,N_3104,N_3136);
or U3349 (N_3349,N_3047,N_3115);
xnor U3350 (N_3350,N_3183,N_3063);
or U3351 (N_3351,N_3095,N_3109);
or U3352 (N_3352,N_3074,N_3173);
or U3353 (N_3353,N_3100,N_3017);
or U3354 (N_3354,N_3045,N_3122);
nand U3355 (N_3355,N_3057,N_3087);
or U3356 (N_3356,N_3165,N_3047);
and U3357 (N_3357,N_3171,N_3102);
nor U3358 (N_3358,N_3193,N_3157);
and U3359 (N_3359,N_3122,N_3156);
xnor U3360 (N_3360,N_3026,N_3040);
and U3361 (N_3361,N_3092,N_3032);
or U3362 (N_3362,N_3059,N_3136);
xnor U3363 (N_3363,N_3101,N_3198);
nor U3364 (N_3364,N_3100,N_3073);
and U3365 (N_3365,N_3068,N_3041);
xor U3366 (N_3366,N_3094,N_3122);
and U3367 (N_3367,N_3042,N_3075);
nor U3368 (N_3368,N_3133,N_3107);
nand U3369 (N_3369,N_3127,N_3188);
nand U3370 (N_3370,N_3037,N_3077);
nand U3371 (N_3371,N_3029,N_3105);
nor U3372 (N_3372,N_3003,N_3024);
or U3373 (N_3373,N_3121,N_3066);
and U3374 (N_3374,N_3111,N_3035);
nor U3375 (N_3375,N_3188,N_3013);
nor U3376 (N_3376,N_3004,N_3174);
and U3377 (N_3377,N_3085,N_3080);
nor U3378 (N_3378,N_3139,N_3065);
or U3379 (N_3379,N_3086,N_3164);
and U3380 (N_3380,N_3043,N_3191);
nand U3381 (N_3381,N_3147,N_3109);
nor U3382 (N_3382,N_3100,N_3163);
nand U3383 (N_3383,N_3196,N_3036);
and U3384 (N_3384,N_3101,N_3079);
and U3385 (N_3385,N_3018,N_3122);
and U3386 (N_3386,N_3100,N_3105);
xnor U3387 (N_3387,N_3006,N_3159);
nand U3388 (N_3388,N_3052,N_3151);
xor U3389 (N_3389,N_3143,N_3096);
xor U3390 (N_3390,N_3041,N_3043);
and U3391 (N_3391,N_3121,N_3044);
nor U3392 (N_3392,N_3194,N_3191);
or U3393 (N_3393,N_3062,N_3070);
nor U3394 (N_3394,N_3142,N_3098);
nand U3395 (N_3395,N_3112,N_3034);
nand U3396 (N_3396,N_3104,N_3158);
or U3397 (N_3397,N_3043,N_3121);
nor U3398 (N_3398,N_3125,N_3104);
or U3399 (N_3399,N_3002,N_3003);
and U3400 (N_3400,N_3251,N_3395);
nand U3401 (N_3401,N_3365,N_3333);
xor U3402 (N_3402,N_3260,N_3212);
and U3403 (N_3403,N_3254,N_3200);
or U3404 (N_3404,N_3296,N_3324);
nor U3405 (N_3405,N_3344,N_3343);
nand U3406 (N_3406,N_3244,N_3388);
and U3407 (N_3407,N_3261,N_3201);
and U3408 (N_3408,N_3317,N_3289);
or U3409 (N_3409,N_3308,N_3265);
nand U3410 (N_3410,N_3266,N_3275);
or U3411 (N_3411,N_3239,N_3358);
nor U3412 (N_3412,N_3224,N_3312);
nand U3413 (N_3413,N_3335,N_3277);
or U3414 (N_3414,N_3374,N_3379);
nand U3415 (N_3415,N_3382,N_3264);
or U3416 (N_3416,N_3357,N_3348);
and U3417 (N_3417,N_3286,N_3228);
nor U3418 (N_3418,N_3351,N_3233);
xnor U3419 (N_3419,N_3354,N_3257);
xnor U3420 (N_3420,N_3282,N_3340);
and U3421 (N_3421,N_3391,N_3226);
and U3422 (N_3422,N_3334,N_3283);
or U3423 (N_3423,N_3274,N_3370);
nand U3424 (N_3424,N_3246,N_3259);
xnor U3425 (N_3425,N_3380,N_3235);
and U3426 (N_3426,N_3318,N_3278);
nand U3427 (N_3427,N_3303,N_3225);
or U3428 (N_3428,N_3373,N_3216);
nand U3429 (N_3429,N_3315,N_3396);
nor U3430 (N_3430,N_3218,N_3258);
nand U3431 (N_3431,N_3346,N_3276);
or U3432 (N_3432,N_3353,N_3291);
xor U3433 (N_3433,N_3364,N_3309);
nand U3434 (N_3434,N_3304,N_3214);
and U3435 (N_3435,N_3394,N_3241);
nor U3436 (N_3436,N_3256,N_3386);
and U3437 (N_3437,N_3389,N_3284);
or U3438 (N_3438,N_3299,N_3230);
nand U3439 (N_3439,N_3295,N_3316);
nor U3440 (N_3440,N_3247,N_3285);
or U3441 (N_3441,N_3387,N_3223);
and U3442 (N_3442,N_3337,N_3271);
nand U3443 (N_3443,N_3281,N_3398);
and U3444 (N_3444,N_3345,N_3359);
or U3445 (N_3445,N_3210,N_3384);
or U3446 (N_3446,N_3305,N_3360);
nor U3447 (N_3447,N_3272,N_3252);
nand U3448 (N_3448,N_3242,N_3207);
and U3449 (N_3449,N_3399,N_3378);
nand U3450 (N_3450,N_3342,N_3206);
or U3451 (N_3451,N_3323,N_3270);
and U3452 (N_3452,N_3222,N_3383);
xor U3453 (N_3453,N_3329,N_3372);
and U3454 (N_3454,N_3263,N_3377);
and U3455 (N_3455,N_3211,N_3215);
nand U3456 (N_3456,N_3371,N_3208);
or U3457 (N_3457,N_3220,N_3385);
nand U3458 (N_3458,N_3249,N_3302);
nor U3459 (N_3459,N_3310,N_3376);
nor U3460 (N_3460,N_3203,N_3234);
or U3461 (N_3461,N_3321,N_3325);
or U3462 (N_3462,N_3350,N_3231);
and U3463 (N_3463,N_3229,N_3341);
xor U3464 (N_3464,N_3237,N_3352);
nand U3465 (N_3465,N_3301,N_3307);
nand U3466 (N_3466,N_3262,N_3253);
nand U3467 (N_3467,N_3397,N_3273);
xnor U3468 (N_3468,N_3250,N_3287);
nand U3469 (N_3469,N_3269,N_3313);
and U3470 (N_3470,N_3297,N_3355);
nor U3471 (N_3471,N_3356,N_3361);
or U3472 (N_3472,N_3227,N_3236);
nand U3473 (N_3473,N_3213,N_3204);
nor U3474 (N_3474,N_3339,N_3338);
or U3475 (N_3475,N_3392,N_3322);
and U3476 (N_3476,N_3298,N_3292);
nand U3477 (N_3477,N_3390,N_3367);
and U3478 (N_3478,N_3243,N_3363);
or U3479 (N_3479,N_3349,N_3255);
nand U3480 (N_3480,N_3288,N_3311);
nand U3481 (N_3481,N_3202,N_3294);
nand U3482 (N_3482,N_3293,N_3238);
and U3483 (N_3483,N_3381,N_3217);
or U3484 (N_3484,N_3336,N_3347);
or U3485 (N_3485,N_3267,N_3279);
or U3486 (N_3486,N_3245,N_3314);
and U3487 (N_3487,N_3209,N_3362);
nand U3488 (N_3488,N_3248,N_3290);
nand U3489 (N_3489,N_3393,N_3205);
and U3490 (N_3490,N_3369,N_3326);
and U3491 (N_3491,N_3332,N_3232);
and U3492 (N_3492,N_3328,N_3327);
or U3493 (N_3493,N_3280,N_3319);
nor U3494 (N_3494,N_3330,N_3368);
nor U3495 (N_3495,N_3366,N_3306);
or U3496 (N_3496,N_3300,N_3219);
nor U3497 (N_3497,N_3221,N_3240);
nand U3498 (N_3498,N_3320,N_3331);
and U3499 (N_3499,N_3268,N_3375);
and U3500 (N_3500,N_3339,N_3372);
nand U3501 (N_3501,N_3205,N_3318);
and U3502 (N_3502,N_3330,N_3346);
nor U3503 (N_3503,N_3343,N_3248);
nand U3504 (N_3504,N_3391,N_3353);
nor U3505 (N_3505,N_3392,N_3206);
nor U3506 (N_3506,N_3310,N_3366);
or U3507 (N_3507,N_3278,N_3376);
or U3508 (N_3508,N_3376,N_3210);
and U3509 (N_3509,N_3357,N_3313);
nor U3510 (N_3510,N_3319,N_3220);
and U3511 (N_3511,N_3342,N_3217);
nor U3512 (N_3512,N_3324,N_3226);
nor U3513 (N_3513,N_3229,N_3398);
or U3514 (N_3514,N_3337,N_3264);
nor U3515 (N_3515,N_3320,N_3392);
nor U3516 (N_3516,N_3207,N_3310);
nand U3517 (N_3517,N_3254,N_3256);
nor U3518 (N_3518,N_3391,N_3304);
nand U3519 (N_3519,N_3222,N_3376);
nand U3520 (N_3520,N_3252,N_3214);
nor U3521 (N_3521,N_3398,N_3295);
or U3522 (N_3522,N_3254,N_3284);
or U3523 (N_3523,N_3214,N_3299);
and U3524 (N_3524,N_3216,N_3365);
and U3525 (N_3525,N_3326,N_3320);
nor U3526 (N_3526,N_3346,N_3259);
and U3527 (N_3527,N_3385,N_3376);
nand U3528 (N_3528,N_3334,N_3217);
nand U3529 (N_3529,N_3292,N_3219);
nand U3530 (N_3530,N_3269,N_3280);
and U3531 (N_3531,N_3295,N_3226);
or U3532 (N_3532,N_3201,N_3319);
and U3533 (N_3533,N_3316,N_3345);
or U3534 (N_3534,N_3213,N_3216);
and U3535 (N_3535,N_3357,N_3254);
and U3536 (N_3536,N_3225,N_3394);
nor U3537 (N_3537,N_3296,N_3214);
and U3538 (N_3538,N_3367,N_3282);
nor U3539 (N_3539,N_3251,N_3304);
nand U3540 (N_3540,N_3341,N_3326);
nor U3541 (N_3541,N_3224,N_3254);
and U3542 (N_3542,N_3319,N_3271);
or U3543 (N_3543,N_3389,N_3238);
xnor U3544 (N_3544,N_3246,N_3381);
nand U3545 (N_3545,N_3257,N_3398);
nor U3546 (N_3546,N_3290,N_3238);
xor U3547 (N_3547,N_3247,N_3273);
nand U3548 (N_3548,N_3216,N_3239);
nor U3549 (N_3549,N_3202,N_3383);
nand U3550 (N_3550,N_3376,N_3313);
xor U3551 (N_3551,N_3288,N_3227);
nor U3552 (N_3552,N_3222,N_3357);
and U3553 (N_3553,N_3326,N_3286);
nor U3554 (N_3554,N_3319,N_3252);
nor U3555 (N_3555,N_3209,N_3307);
nand U3556 (N_3556,N_3341,N_3306);
and U3557 (N_3557,N_3359,N_3334);
and U3558 (N_3558,N_3268,N_3319);
or U3559 (N_3559,N_3314,N_3207);
nand U3560 (N_3560,N_3364,N_3295);
and U3561 (N_3561,N_3237,N_3327);
xnor U3562 (N_3562,N_3391,N_3266);
or U3563 (N_3563,N_3298,N_3246);
nor U3564 (N_3564,N_3334,N_3261);
nand U3565 (N_3565,N_3239,N_3399);
nand U3566 (N_3566,N_3290,N_3207);
or U3567 (N_3567,N_3305,N_3211);
nand U3568 (N_3568,N_3238,N_3258);
xor U3569 (N_3569,N_3276,N_3250);
nand U3570 (N_3570,N_3374,N_3348);
and U3571 (N_3571,N_3346,N_3308);
nand U3572 (N_3572,N_3371,N_3278);
and U3573 (N_3573,N_3349,N_3269);
and U3574 (N_3574,N_3316,N_3242);
nor U3575 (N_3575,N_3344,N_3390);
nor U3576 (N_3576,N_3237,N_3273);
nand U3577 (N_3577,N_3228,N_3300);
and U3578 (N_3578,N_3302,N_3248);
nor U3579 (N_3579,N_3216,N_3269);
or U3580 (N_3580,N_3204,N_3263);
nand U3581 (N_3581,N_3219,N_3318);
and U3582 (N_3582,N_3229,N_3364);
nand U3583 (N_3583,N_3282,N_3324);
and U3584 (N_3584,N_3211,N_3346);
nand U3585 (N_3585,N_3309,N_3345);
and U3586 (N_3586,N_3340,N_3248);
nand U3587 (N_3587,N_3228,N_3202);
nand U3588 (N_3588,N_3269,N_3340);
nor U3589 (N_3589,N_3257,N_3306);
nor U3590 (N_3590,N_3275,N_3352);
or U3591 (N_3591,N_3352,N_3207);
and U3592 (N_3592,N_3209,N_3231);
and U3593 (N_3593,N_3346,N_3315);
nor U3594 (N_3594,N_3340,N_3301);
and U3595 (N_3595,N_3272,N_3367);
xor U3596 (N_3596,N_3285,N_3201);
nor U3597 (N_3597,N_3338,N_3244);
xnor U3598 (N_3598,N_3358,N_3275);
xnor U3599 (N_3599,N_3286,N_3299);
or U3600 (N_3600,N_3575,N_3526);
or U3601 (N_3601,N_3408,N_3412);
nor U3602 (N_3602,N_3481,N_3509);
or U3603 (N_3603,N_3537,N_3416);
nor U3604 (N_3604,N_3572,N_3402);
or U3605 (N_3605,N_3593,N_3518);
nand U3606 (N_3606,N_3429,N_3542);
and U3607 (N_3607,N_3425,N_3550);
or U3608 (N_3608,N_3442,N_3553);
or U3609 (N_3609,N_3534,N_3592);
and U3610 (N_3610,N_3434,N_3557);
or U3611 (N_3611,N_3414,N_3454);
nor U3612 (N_3612,N_3552,N_3480);
nor U3613 (N_3613,N_3587,N_3490);
nor U3614 (N_3614,N_3532,N_3515);
or U3615 (N_3615,N_3535,N_3413);
nand U3616 (N_3616,N_3584,N_3500);
nor U3617 (N_3617,N_3488,N_3496);
or U3618 (N_3618,N_3574,N_3486);
nor U3619 (N_3619,N_3428,N_3440);
and U3620 (N_3620,N_3502,N_3560);
nor U3621 (N_3621,N_3436,N_3512);
and U3622 (N_3622,N_3471,N_3426);
and U3623 (N_3623,N_3459,N_3523);
or U3624 (N_3624,N_3571,N_3499);
or U3625 (N_3625,N_3430,N_3498);
xor U3626 (N_3626,N_3415,N_3458);
nor U3627 (N_3627,N_3541,N_3507);
nand U3628 (N_3628,N_3448,N_3524);
and U3629 (N_3629,N_3452,N_3595);
nor U3630 (N_3630,N_3439,N_3576);
and U3631 (N_3631,N_3463,N_3545);
and U3632 (N_3632,N_3464,N_3418);
or U3633 (N_3633,N_3599,N_3438);
nor U3634 (N_3634,N_3483,N_3527);
nand U3635 (N_3635,N_3549,N_3585);
and U3636 (N_3636,N_3521,N_3403);
nor U3637 (N_3637,N_3479,N_3437);
xnor U3638 (N_3638,N_3462,N_3580);
nand U3639 (N_3639,N_3538,N_3495);
nand U3640 (N_3640,N_3525,N_3457);
and U3641 (N_3641,N_3531,N_3445);
or U3642 (N_3642,N_3563,N_3533);
nor U3643 (N_3643,N_3564,N_3485);
or U3644 (N_3644,N_3583,N_3513);
and U3645 (N_3645,N_3597,N_3594);
and U3646 (N_3646,N_3506,N_3422);
nand U3647 (N_3647,N_3472,N_3424);
xnor U3648 (N_3648,N_3474,N_3477);
or U3649 (N_3649,N_3579,N_3517);
and U3650 (N_3650,N_3450,N_3559);
nand U3651 (N_3651,N_3561,N_3590);
or U3652 (N_3652,N_3432,N_3591);
or U3653 (N_3653,N_3582,N_3484);
and U3654 (N_3654,N_3494,N_3562);
and U3655 (N_3655,N_3470,N_3455);
and U3656 (N_3656,N_3478,N_3501);
nor U3657 (N_3657,N_3514,N_3406);
nor U3658 (N_3658,N_3530,N_3508);
or U3659 (N_3659,N_3570,N_3420);
and U3660 (N_3660,N_3404,N_3573);
and U3661 (N_3661,N_3577,N_3447);
xor U3662 (N_3662,N_3578,N_3421);
or U3663 (N_3663,N_3473,N_3487);
or U3664 (N_3664,N_3551,N_3558);
or U3665 (N_3665,N_3407,N_3504);
nand U3666 (N_3666,N_3493,N_3453);
nor U3667 (N_3667,N_3423,N_3466);
xnor U3668 (N_3668,N_3548,N_3546);
or U3669 (N_3669,N_3443,N_3409);
and U3670 (N_3670,N_3411,N_3433);
or U3671 (N_3671,N_3461,N_3468);
nand U3672 (N_3672,N_3446,N_3555);
nor U3673 (N_3673,N_3544,N_3522);
or U3674 (N_3674,N_3581,N_3503);
nor U3675 (N_3675,N_3475,N_3569);
and U3676 (N_3676,N_3510,N_3511);
nor U3677 (N_3677,N_3519,N_3489);
nor U3678 (N_3678,N_3505,N_3482);
or U3679 (N_3679,N_3540,N_3543);
and U3680 (N_3680,N_3491,N_3539);
or U3681 (N_3681,N_3417,N_3410);
nor U3682 (N_3682,N_3431,N_3456);
or U3683 (N_3683,N_3405,N_3401);
and U3684 (N_3684,N_3451,N_3528);
nand U3685 (N_3685,N_3467,N_3427);
xnor U3686 (N_3686,N_3596,N_3435);
and U3687 (N_3687,N_3566,N_3419);
or U3688 (N_3688,N_3516,N_3476);
or U3689 (N_3689,N_3465,N_3520);
and U3690 (N_3690,N_3529,N_3547);
and U3691 (N_3691,N_3589,N_3441);
or U3692 (N_3692,N_3556,N_3444);
and U3693 (N_3693,N_3400,N_3588);
nand U3694 (N_3694,N_3536,N_3565);
nor U3695 (N_3695,N_3449,N_3497);
nand U3696 (N_3696,N_3460,N_3598);
or U3697 (N_3697,N_3586,N_3554);
or U3698 (N_3698,N_3567,N_3492);
and U3699 (N_3699,N_3469,N_3568);
and U3700 (N_3700,N_3423,N_3412);
nor U3701 (N_3701,N_3405,N_3503);
or U3702 (N_3702,N_3570,N_3457);
or U3703 (N_3703,N_3544,N_3436);
nand U3704 (N_3704,N_3498,N_3451);
nor U3705 (N_3705,N_3565,N_3431);
nand U3706 (N_3706,N_3470,N_3521);
xnor U3707 (N_3707,N_3532,N_3412);
and U3708 (N_3708,N_3464,N_3554);
nand U3709 (N_3709,N_3415,N_3563);
and U3710 (N_3710,N_3542,N_3569);
xnor U3711 (N_3711,N_3544,N_3536);
nand U3712 (N_3712,N_3416,N_3522);
nor U3713 (N_3713,N_3570,N_3573);
or U3714 (N_3714,N_3445,N_3527);
or U3715 (N_3715,N_3420,N_3478);
nand U3716 (N_3716,N_3543,N_3515);
nand U3717 (N_3717,N_3456,N_3458);
nand U3718 (N_3718,N_3490,N_3536);
nand U3719 (N_3719,N_3587,N_3577);
nor U3720 (N_3720,N_3490,N_3512);
nor U3721 (N_3721,N_3547,N_3412);
nand U3722 (N_3722,N_3491,N_3577);
or U3723 (N_3723,N_3591,N_3559);
and U3724 (N_3724,N_3445,N_3459);
or U3725 (N_3725,N_3437,N_3504);
nor U3726 (N_3726,N_3526,N_3532);
nor U3727 (N_3727,N_3551,N_3502);
or U3728 (N_3728,N_3501,N_3529);
and U3729 (N_3729,N_3495,N_3569);
xor U3730 (N_3730,N_3594,N_3472);
nor U3731 (N_3731,N_3406,N_3553);
nor U3732 (N_3732,N_3547,N_3432);
nor U3733 (N_3733,N_3409,N_3501);
nand U3734 (N_3734,N_3483,N_3496);
and U3735 (N_3735,N_3512,N_3478);
xnor U3736 (N_3736,N_3460,N_3426);
or U3737 (N_3737,N_3481,N_3429);
or U3738 (N_3738,N_3446,N_3509);
nand U3739 (N_3739,N_3483,N_3534);
nand U3740 (N_3740,N_3401,N_3537);
nand U3741 (N_3741,N_3466,N_3475);
and U3742 (N_3742,N_3596,N_3444);
or U3743 (N_3743,N_3584,N_3574);
xnor U3744 (N_3744,N_3473,N_3486);
xnor U3745 (N_3745,N_3492,N_3543);
and U3746 (N_3746,N_3484,N_3444);
nand U3747 (N_3747,N_3444,N_3535);
nand U3748 (N_3748,N_3549,N_3403);
or U3749 (N_3749,N_3537,N_3566);
nor U3750 (N_3750,N_3515,N_3409);
nand U3751 (N_3751,N_3499,N_3556);
or U3752 (N_3752,N_3531,N_3577);
or U3753 (N_3753,N_3472,N_3496);
and U3754 (N_3754,N_3558,N_3593);
nand U3755 (N_3755,N_3517,N_3483);
nand U3756 (N_3756,N_3478,N_3541);
nand U3757 (N_3757,N_3405,N_3544);
and U3758 (N_3758,N_3561,N_3562);
nand U3759 (N_3759,N_3429,N_3521);
or U3760 (N_3760,N_3459,N_3458);
nand U3761 (N_3761,N_3506,N_3456);
nand U3762 (N_3762,N_3444,N_3429);
nor U3763 (N_3763,N_3564,N_3406);
nand U3764 (N_3764,N_3507,N_3519);
or U3765 (N_3765,N_3466,N_3524);
and U3766 (N_3766,N_3554,N_3569);
or U3767 (N_3767,N_3429,N_3407);
xor U3768 (N_3768,N_3598,N_3556);
and U3769 (N_3769,N_3423,N_3527);
nor U3770 (N_3770,N_3484,N_3485);
nor U3771 (N_3771,N_3458,N_3407);
nand U3772 (N_3772,N_3547,N_3425);
nand U3773 (N_3773,N_3560,N_3562);
or U3774 (N_3774,N_3427,N_3407);
nand U3775 (N_3775,N_3468,N_3485);
nor U3776 (N_3776,N_3590,N_3481);
and U3777 (N_3777,N_3524,N_3400);
nand U3778 (N_3778,N_3482,N_3580);
xnor U3779 (N_3779,N_3586,N_3489);
and U3780 (N_3780,N_3511,N_3503);
and U3781 (N_3781,N_3580,N_3491);
nand U3782 (N_3782,N_3427,N_3590);
nand U3783 (N_3783,N_3482,N_3587);
xor U3784 (N_3784,N_3425,N_3599);
nor U3785 (N_3785,N_3522,N_3422);
nor U3786 (N_3786,N_3533,N_3593);
and U3787 (N_3787,N_3400,N_3578);
and U3788 (N_3788,N_3519,N_3547);
xor U3789 (N_3789,N_3496,N_3574);
nand U3790 (N_3790,N_3508,N_3443);
and U3791 (N_3791,N_3464,N_3476);
nand U3792 (N_3792,N_3409,N_3484);
and U3793 (N_3793,N_3410,N_3496);
or U3794 (N_3794,N_3462,N_3525);
nand U3795 (N_3795,N_3568,N_3572);
and U3796 (N_3796,N_3423,N_3428);
and U3797 (N_3797,N_3545,N_3407);
and U3798 (N_3798,N_3438,N_3595);
nand U3799 (N_3799,N_3446,N_3420);
and U3800 (N_3800,N_3608,N_3747);
or U3801 (N_3801,N_3750,N_3668);
and U3802 (N_3802,N_3791,N_3799);
nor U3803 (N_3803,N_3624,N_3636);
or U3804 (N_3804,N_3725,N_3775);
nor U3805 (N_3805,N_3789,N_3715);
xnor U3806 (N_3806,N_3759,N_3797);
or U3807 (N_3807,N_3626,N_3634);
nor U3808 (N_3808,N_3704,N_3712);
nor U3809 (N_3809,N_3758,N_3613);
and U3810 (N_3810,N_3690,N_3697);
nand U3811 (N_3811,N_3693,N_3784);
and U3812 (N_3812,N_3744,N_3787);
and U3813 (N_3813,N_3792,N_3681);
nand U3814 (N_3814,N_3749,N_3772);
nand U3815 (N_3815,N_3615,N_3600);
or U3816 (N_3816,N_3644,N_3620);
nand U3817 (N_3817,N_3798,N_3723);
nand U3818 (N_3818,N_3657,N_3713);
and U3819 (N_3819,N_3619,N_3766);
and U3820 (N_3820,N_3689,N_3622);
nand U3821 (N_3821,N_3655,N_3780);
and U3822 (N_3822,N_3760,N_3762);
and U3823 (N_3823,N_3763,N_3631);
or U3824 (N_3824,N_3732,N_3633);
and U3825 (N_3825,N_3796,N_3670);
and U3826 (N_3826,N_3669,N_3625);
and U3827 (N_3827,N_3771,N_3745);
or U3828 (N_3828,N_3640,N_3730);
xor U3829 (N_3829,N_3793,N_3676);
nor U3830 (N_3830,N_3601,N_3649);
and U3831 (N_3831,N_3687,N_3646);
nor U3832 (N_3832,N_3653,N_3768);
or U3833 (N_3833,N_3662,N_3779);
or U3834 (N_3834,N_3785,N_3647);
nand U3835 (N_3835,N_3674,N_3656);
nand U3836 (N_3836,N_3694,N_3781);
and U3837 (N_3837,N_3686,N_3642);
or U3838 (N_3838,N_3628,N_3663);
nand U3839 (N_3839,N_3664,N_3773);
or U3840 (N_3840,N_3609,N_3714);
or U3841 (N_3841,N_3707,N_3765);
nor U3842 (N_3842,N_3729,N_3722);
and U3843 (N_3843,N_3795,N_3726);
nor U3844 (N_3844,N_3740,N_3691);
or U3845 (N_3845,N_3743,N_3685);
or U3846 (N_3846,N_3692,N_3724);
and U3847 (N_3847,N_3643,N_3737);
nor U3848 (N_3848,N_3777,N_3651);
xor U3849 (N_3849,N_3679,N_3720);
or U3850 (N_3850,N_3728,N_3705);
or U3851 (N_3851,N_3774,N_3736);
nor U3852 (N_3852,N_3614,N_3621);
and U3853 (N_3853,N_3683,N_3731);
or U3854 (N_3854,N_3635,N_3700);
or U3855 (N_3855,N_3672,N_3603);
and U3856 (N_3856,N_3639,N_3710);
nor U3857 (N_3857,N_3719,N_3671);
nand U3858 (N_3858,N_3755,N_3682);
nand U3859 (N_3859,N_3703,N_3660);
and U3860 (N_3860,N_3778,N_3733);
nand U3861 (N_3861,N_3654,N_3767);
nor U3862 (N_3862,N_3673,N_3742);
nand U3863 (N_3863,N_3716,N_3718);
or U3864 (N_3864,N_3616,N_3738);
and U3865 (N_3865,N_3790,N_3698);
or U3866 (N_3866,N_3680,N_3727);
or U3867 (N_3867,N_3623,N_3627);
nor U3868 (N_3868,N_3607,N_3666);
or U3869 (N_3869,N_3786,N_3699);
and U3870 (N_3870,N_3734,N_3610);
and U3871 (N_3871,N_3788,N_3641);
nand U3872 (N_3872,N_3688,N_3761);
and U3873 (N_3873,N_3783,N_3630);
xor U3874 (N_3874,N_3675,N_3648);
or U3875 (N_3875,N_3604,N_3770);
or U3876 (N_3876,N_3739,N_3708);
and U3877 (N_3877,N_3632,N_3752);
and U3878 (N_3878,N_3717,N_3618);
nand U3879 (N_3879,N_3606,N_3782);
nor U3880 (N_3880,N_3794,N_3735);
nor U3881 (N_3881,N_3711,N_3611);
nand U3882 (N_3882,N_3605,N_3695);
nand U3883 (N_3883,N_3677,N_3652);
nor U3884 (N_3884,N_3764,N_3701);
or U3885 (N_3885,N_3706,N_3741);
or U3886 (N_3886,N_3684,N_3667);
nand U3887 (N_3887,N_3721,N_3665);
or U3888 (N_3888,N_3638,N_3637);
or U3889 (N_3889,N_3661,N_3746);
nor U3890 (N_3890,N_3658,N_3748);
or U3891 (N_3891,N_3709,N_3696);
or U3892 (N_3892,N_3659,N_3612);
nand U3893 (N_3893,N_3629,N_3754);
nand U3894 (N_3894,N_3650,N_3776);
nor U3895 (N_3895,N_3702,N_3769);
nand U3896 (N_3896,N_3617,N_3678);
nand U3897 (N_3897,N_3756,N_3602);
nand U3898 (N_3898,N_3757,N_3753);
nor U3899 (N_3899,N_3645,N_3751);
nor U3900 (N_3900,N_3775,N_3741);
and U3901 (N_3901,N_3757,N_3612);
or U3902 (N_3902,N_3686,N_3666);
and U3903 (N_3903,N_3646,N_3623);
or U3904 (N_3904,N_3678,N_3707);
nand U3905 (N_3905,N_3679,N_3601);
nor U3906 (N_3906,N_3707,N_3737);
or U3907 (N_3907,N_3701,N_3694);
and U3908 (N_3908,N_3604,N_3789);
nor U3909 (N_3909,N_3613,N_3649);
or U3910 (N_3910,N_3672,N_3740);
or U3911 (N_3911,N_3745,N_3755);
nor U3912 (N_3912,N_3664,N_3742);
or U3913 (N_3913,N_3733,N_3704);
or U3914 (N_3914,N_3605,N_3701);
or U3915 (N_3915,N_3682,N_3616);
or U3916 (N_3916,N_3614,N_3688);
nand U3917 (N_3917,N_3718,N_3768);
and U3918 (N_3918,N_3773,N_3665);
nor U3919 (N_3919,N_3710,N_3614);
or U3920 (N_3920,N_3763,N_3738);
nand U3921 (N_3921,N_3695,N_3673);
and U3922 (N_3922,N_3632,N_3698);
nor U3923 (N_3923,N_3756,N_3685);
and U3924 (N_3924,N_3781,N_3730);
and U3925 (N_3925,N_3718,N_3695);
and U3926 (N_3926,N_3710,N_3758);
and U3927 (N_3927,N_3702,N_3663);
nand U3928 (N_3928,N_3619,N_3753);
xor U3929 (N_3929,N_3667,N_3666);
and U3930 (N_3930,N_3786,N_3728);
xnor U3931 (N_3931,N_3624,N_3629);
nand U3932 (N_3932,N_3769,N_3666);
and U3933 (N_3933,N_3673,N_3717);
or U3934 (N_3934,N_3668,N_3665);
xnor U3935 (N_3935,N_3783,N_3600);
xor U3936 (N_3936,N_3709,N_3610);
nor U3937 (N_3937,N_3642,N_3756);
or U3938 (N_3938,N_3607,N_3618);
or U3939 (N_3939,N_3627,N_3699);
nor U3940 (N_3940,N_3793,N_3753);
or U3941 (N_3941,N_3651,N_3634);
and U3942 (N_3942,N_3601,N_3617);
or U3943 (N_3943,N_3678,N_3611);
or U3944 (N_3944,N_3644,N_3757);
and U3945 (N_3945,N_3728,N_3635);
and U3946 (N_3946,N_3658,N_3721);
and U3947 (N_3947,N_3600,N_3618);
or U3948 (N_3948,N_3637,N_3668);
nand U3949 (N_3949,N_3726,N_3687);
xnor U3950 (N_3950,N_3769,N_3740);
nand U3951 (N_3951,N_3716,N_3733);
nand U3952 (N_3952,N_3632,N_3654);
or U3953 (N_3953,N_3674,N_3749);
xor U3954 (N_3954,N_3785,N_3612);
nand U3955 (N_3955,N_3696,N_3796);
nor U3956 (N_3956,N_3765,N_3767);
or U3957 (N_3957,N_3711,N_3609);
and U3958 (N_3958,N_3715,N_3795);
or U3959 (N_3959,N_3642,N_3782);
nand U3960 (N_3960,N_3629,N_3652);
nand U3961 (N_3961,N_3631,N_3625);
or U3962 (N_3962,N_3688,N_3635);
or U3963 (N_3963,N_3628,N_3783);
nand U3964 (N_3964,N_3780,N_3751);
or U3965 (N_3965,N_3625,N_3682);
nor U3966 (N_3966,N_3703,N_3602);
nand U3967 (N_3967,N_3763,N_3760);
xor U3968 (N_3968,N_3767,N_3644);
or U3969 (N_3969,N_3729,N_3672);
nor U3970 (N_3970,N_3772,N_3624);
nor U3971 (N_3971,N_3770,N_3753);
xnor U3972 (N_3972,N_3776,N_3640);
and U3973 (N_3973,N_3705,N_3768);
or U3974 (N_3974,N_3797,N_3752);
or U3975 (N_3975,N_3649,N_3679);
nand U3976 (N_3976,N_3701,N_3712);
or U3977 (N_3977,N_3743,N_3714);
and U3978 (N_3978,N_3698,N_3644);
xor U3979 (N_3979,N_3653,N_3722);
xor U3980 (N_3980,N_3734,N_3760);
nor U3981 (N_3981,N_3641,N_3647);
and U3982 (N_3982,N_3750,N_3737);
nor U3983 (N_3983,N_3684,N_3648);
nand U3984 (N_3984,N_3771,N_3678);
nor U3985 (N_3985,N_3628,N_3730);
and U3986 (N_3986,N_3758,N_3675);
nor U3987 (N_3987,N_3619,N_3686);
nor U3988 (N_3988,N_3738,N_3629);
nor U3989 (N_3989,N_3644,N_3771);
xor U3990 (N_3990,N_3636,N_3776);
nand U3991 (N_3991,N_3731,N_3768);
xnor U3992 (N_3992,N_3684,N_3688);
xnor U3993 (N_3993,N_3795,N_3745);
nor U3994 (N_3994,N_3651,N_3711);
or U3995 (N_3995,N_3700,N_3611);
and U3996 (N_3996,N_3782,N_3647);
nor U3997 (N_3997,N_3785,N_3733);
nand U3998 (N_3998,N_3675,N_3634);
nor U3999 (N_3999,N_3631,N_3603);
nand U4000 (N_4000,N_3868,N_3813);
and U4001 (N_4001,N_3841,N_3968);
and U4002 (N_4002,N_3983,N_3904);
and U4003 (N_4003,N_3817,N_3892);
nor U4004 (N_4004,N_3917,N_3828);
nand U4005 (N_4005,N_3862,N_3914);
and U4006 (N_4006,N_3824,N_3972);
nor U4007 (N_4007,N_3891,N_3937);
or U4008 (N_4008,N_3884,N_3926);
nor U4009 (N_4009,N_3975,N_3872);
nor U4010 (N_4010,N_3910,N_3913);
or U4011 (N_4011,N_3846,N_3850);
nor U4012 (N_4012,N_3903,N_3920);
nand U4013 (N_4013,N_3958,N_3804);
nor U4014 (N_4014,N_3946,N_3848);
nor U4015 (N_4015,N_3854,N_3949);
or U4016 (N_4016,N_3996,N_3927);
or U4017 (N_4017,N_3833,N_3918);
or U4018 (N_4018,N_3830,N_3901);
nor U4019 (N_4019,N_3998,N_3896);
nor U4020 (N_4020,N_3948,N_3974);
xor U4021 (N_4021,N_3823,N_3870);
nand U4022 (N_4022,N_3963,N_3933);
xnor U4023 (N_4023,N_3905,N_3831);
nor U4024 (N_4024,N_3907,N_3849);
xor U4025 (N_4025,N_3809,N_3990);
nand U4026 (N_4026,N_3919,N_3827);
or U4027 (N_4027,N_3940,N_3924);
nor U4028 (N_4028,N_3985,N_3880);
nand U4029 (N_4029,N_3886,N_3806);
nor U4030 (N_4030,N_3935,N_3947);
or U4031 (N_4031,N_3925,N_3954);
nand U4032 (N_4032,N_3962,N_3931);
and U4033 (N_4033,N_3936,N_3911);
nand U4034 (N_4034,N_3863,N_3888);
and U4035 (N_4035,N_3916,N_3982);
and U4036 (N_4036,N_3944,N_3842);
nand U4037 (N_4037,N_3825,N_3984);
nand U4038 (N_4038,N_3898,N_3932);
xnor U4039 (N_4039,N_3969,N_3909);
nand U4040 (N_4040,N_3822,N_3875);
xor U4041 (N_4041,N_3882,N_3897);
xor U4042 (N_4042,N_3836,N_3816);
and U4043 (N_4043,N_3808,N_3908);
nor U4044 (N_4044,N_3953,N_3885);
xor U4045 (N_4045,N_3820,N_3902);
nand U4046 (N_4046,N_3801,N_3877);
and U4047 (N_4047,N_3921,N_3859);
nor U4048 (N_4048,N_3802,N_3950);
or U4049 (N_4049,N_3895,N_3951);
nor U4050 (N_4050,N_3923,N_3930);
xnor U4051 (N_4051,N_3807,N_3894);
nand U4052 (N_4052,N_3855,N_3890);
nor U4053 (N_4053,N_3874,N_3964);
nor U4054 (N_4054,N_3873,N_3865);
or U4055 (N_4055,N_3960,N_3881);
or U4056 (N_4056,N_3893,N_3928);
and U4057 (N_4057,N_3956,N_3973);
nand U4058 (N_4058,N_3976,N_3845);
xor U4059 (N_4059,N_3821,N_3815);
nand U4060 (N_4060,N_3812,N_3826);
and U4061 (N_4061,N_3819,N_3997);
and U4062 (N_4062,N_3803,N_3995);
nand U4063 (N_4063,N_3837,N_3858);
nor U4064 (N_4064,N_3860,N_3853);
and U4065 (N_4065,N_3899,N_3942);
nor U4066 (N_4066,N_3967,N_3867);
or U4067 (N_4067,N_3988,N_3994);
and U4068 (N_4068,N_3987,N_3939);
or U4069 (N_4069,N_3945,N_3887);
nor U4070 (N_4070,N_3943,N_3999);
and U4071 (N_4071,N_3941,N_3957);
or U4072 (N_4072,N_3843,N_3906);
nand U4073 (N_4073,N_3986,N_3800);
nor U4074 (N_4074,N_3856,N_3844);
and U4075 (N_4075,N_3981,N_3915);
nand U4076 (N_4076,N_3955,N_3811);
or U4077 (N_4077,N_3971,N_3991);
and U4078 (N_4078,N_3889,N_3829);
nand U4079 (N_4079,N_3970,N_3834);
or U4080 (N_4080,N_3878,N_3851);
or U4081 (N_4081,N_3832,N_3838);
xor U4082 (N_4082,N_3861,N_3883);
nor U4083 (N_4083,N_3938,N_3929);
or U4084 (N_4084,N_3966,N_3852);
xnor U4085 (N_4085,N_3818,N_3980);
nor U4086 (N_4086,N_3847,N_3805);
nand U4087 (N_4087,N_3869,N_3961);
and U4088 (N_4088,N_3814,N_3839);
or U4089 (N_4089,N_3989,N_3857);
and U4090 (N_4090,N_3900,N_3934);
or U4091 (N_4091,N_3977,N_3835);
or U4092 (N_4092,N_3840,N_3810);
and U4093 (N_4093,N_3866,N_3864);
nand U4094 (N_4094,N_3912,N_3952);
nand U4095 (N_4095,N_3922,N_3993);
xor U4096 (N_4096,N_3965,N_3979);
and U4097 (N_4097,N_3959,N_3879);
nand U4098 (N_4098,N_3876,N_3992);
nand U4099 (N_4099,N_3978,N_3871);
and U4100 (N_4100,N_3893,N_3944);
nor U4101 (N_4101,N_3900,N_3857);
or U4102 (N_4102,N_3940,N_3823);
and U4103 (N_4103,N_3826,N_3807);
nand U4104 (N_4104,N_3947,N_3890);
or U4105 (N_4105,N_3807,N_3870);
nand U4106 (N_4106,N_3800,N_3990);
and U4107 (N_4107,N_3978,N_3852);
nor U4108 (N_4108,N_3973,N_3940);
nor U4109 (N_4109,N_3903,N_3942);
or U4110 (N_4110,N_3836,N_3916);
nor U4111 (N_4111,N_3951,N_3820);
nand U4112 (N_4112,N_3873,N_3994);
nand U4113 (N_4113,N_3965,N_3948);
nor U4114 (N_4114,N_3802,N_3927);
and U4115 (N_4115,N_3985,N_3922);
xor U4116 (N_4116,N_3848,N_3997);
and U4117 (N_4117,N_3953,N_3966);
xnor U4118 (N_4118,N_3999,N_3916);
nand U4119 (N_4119,N_3846,N_3913);
and U4120 (N_4120,N_3895,N_3908);
xnor U4121 (N_4121,N_3975,N_3878);
and U4122 (N_4122,N_3827,N_3974);
xnor U4123 (N_4123,N_3994,N_3984);
xnor U4124 (N_4124,N_3856,N_3931);
nor U4125 (N_4125,N_3829,N_3947);
nor U4126 (N_4126,N_3939,N_3833);
nor U4127 (N_4127,N_3855,N_3879);
nor U4128 (N_4128,N_3989,N_3816);
or U4129 (N_4129,N_3806,N_3964);
nand U4130 (N_4130,N_3814,N_3907);
nand U4131 (N_4131,N_3983,N_3918);
nor U4132 (N_4132,N_3813,N_3819);
nand U4133 (N_4133,N_3968,N_3860);
and U4134 (N_4134,N_3930,N_3863);
and U4135 (N_4135,N_3841,N_3969);
and U4136 (N_4136,N_3966,N_3849);
nand U4137 (N_4137,N_3932,N_3852);
nor U4138 (N_4138,N_3891,N_3835);
nand U4139 (N_4139,N_3974,N_3907);
nor U4140 (N_4140,N_3820,N_3828);
and U4141 (N_4141,N_3981,N_3892);
or U4142 (N_4142,N_3924,N_3991);
xor U4143 (N_4143,N_3811,N_3923);
and U4144 (N_4144,N_3827,N_3920);
nor U4145 (N_4145,N_3938,N_3964);
nand U4146 (N_4146,N_3867,N_3880);
and U4147 (N_4147,N_3858,N_3900);
nor U4148 (N_4148,N_3833,N_3973);
nand U4149 (N_4149,N_3861,N_3895);
nand U4150 (N_4150,N_3872,N_3846);
nand U4151 (N_4151,N_3925,N_3909);
or U4152 (N_4152,N_3960,N_3856);
and U4153 (N_4153,N_3801,N_3850);
xnor U4154 (N_4154,N_3951,N_3925);
and U4155 (N_4155,N_3937,N_3855);
and U4156 (N_4156,N_3916,N_3814);
or U4157 (N_4157,N_3944,N_3869);
and U4158 (N_4158,N_3895,N_3932);
and U4159 (N_4159,N_3999,N_3859);
and U4160 (N_4160,N_3833,N_3912);
and U4161 (N_4161,N_3828,N_3850);
and U4162 (N_4162,N_3983,N_3825);
and U4163 (N_4163,N_3851,N_3986);
nand U4164 (N_4164,N_3918,N_3876);
or U4165 (N_4165,N_3843,N_3877);
or U4166 (N_4166,N_3848,N_3875);
and U4167 (N_4167,N_3906,N_3979);
or U4168 (N_4168,N_3826,N_3916);
nor U4169 (N_4169,N_3909,N_3849);
or U4170 (N_4170,N_3929,N_3821);
nor U4171 (N_4171,N_3830,N_3960);
nand U4172 (N_4172,N_3863,N_3989);
nand U4173 (N_4173,N_3967,N_3966);
nor U4174 (N_4174,N_3946,N_3893);
and U4175 (N_4175,N_3904,N_3848);
and U4176 (N_4176,N_3915,N_3913);
xor U4177 (N_4177,N_3893,N_3978);
nor U4178 (N_4178,N_3865,N_3900);
xnor U4179 (N_4179,N_3960,N_3966);
nand U4180 (N_4180,N_3870,N_3827);
and U4181 (N_4181,N_3879,N_3915);
or U4182 (N_4182,N_3877,N_3814);
and U4183 (N_4183,N_3864,N_3966);
nand U4184 (N_4184,N_3817,N_3862);
nand U4185 (N_4185,N_3956,N_3972);
and U4186 (N_4186,N_3973,N_3805);
and U4187 (N_4187,N_3881,N_3980);
or U4188 (N_4188,N_3985,N_3863);
nand U4189 (N_4189,N_3854,N_3842);
nor U4190 (N_4190,N_3847,N_3839);
and U4191 (N_4191,N_3897,N_3973);
nand U4192 (N_4192,N_3973,N_3802);
nand U4193 (N_4193,N_3954,N_3984);
and U4194 (N_4194,N_3955,N_3834);
nor U4195 (N_4195,N_3812,N_3974);
nor U4196 (N_4196,N_3802,N_3846);
nor U4197 (N_4197,N_3917,N_3915);
and U4198 (N_4198,N_3902,N_3999);
nor U4199 (N_4199,N_3893,N_3860);
and U4200 (N_4200,N_4111,N_4162);
nand U4201 (N_4201,N_4160,N_4090);
and U4202 (N_4202,N_4018,N_4194);
or U4203 (N_4203,N_4186,N_4150);
nor U4204 (N_4204,N_4098,N_4197);
nand U4205 (N_4205,N_4172,N_4178);
nand U4206 (N_4206,N_4155,N_4142);
and U4207 (N_4207,N_4121,N_4123);
and U4208 (N_4208,N_4112,N_4017);
nor U4209 (N_4209,N_4159,N_4041);
and U4210 (N_4210,N_4161,N_4045);
or U4211 (N_4211,N_4181,N_4184);
nor U4212 (N_4212,N_4087,N_4007);
nor U4213 (N_4213,N_4029,N_4019);
or U4214 (N_4214,N_4156,N_4149);
nand U4215 (N_4215,N_4167,N_4137);
nor U4216 (N_4216,N_4109,N_4026);
and U4217 (N_4217,N_4070,N_4131);
or U4218 (N_4218,N_4085,N_4036);
and U4219 (N_4219,N_4063,N_4073);
and U4220 (N_4220,N_4028,N_4148);
and U4221 (N_4221,N_4116,N_4187);
or U4222 (N_4222,N_4086,N_4147);
xor U4223 (N_4223,N_4152,N_4047);
and U4224 (N_4224,N_4180,N_4190);
nand U4225 (N_4225,N_4127,N_4157);
or U4226 (N_4226,N_4177,N_4032);
or U4227 (N_4227,N_4113,N_4080);
nor U4228 (N_4228,N_4035,N_4074);
and U4229 (N_4229,N_4005,N_4143);
xor U4230 (N_4230,N_4023,N_4075);
nor U4231 (N_4231,N_4058,N_4015);
and U4232 (N_4232,N_4096,N_4014);
nor U4233 (N_4233,N_4012,N_4170);
nor U4234 (N_4234,N_4097,N_4013);
or U4235 (N_4235,N_4044,N_4082);
or U4236 (N_4236,N_4061,N_4000);
or U4237 (N_4237,N_4078,N_4198);
or U4238 (N_4238,N_4049,N_4072);
nand U4239 (N_4239,N_4037,N_4105);
nor U4240 (N_4240,N_4101,N_4196);
and U4241 (N_4241,N_4077,N_4006);
and U4242 (N_4242,N_4089,N_4110);
or U4243 (N_4243,N_4169,N_4158);
nand U4244 (N_4244,N_4002,N_4144);
or U4245 (N_4245,N_4140,N_4107);
nand U4246 (N_4246,N_4125,N_4188);
nand U4247 (N_4247,N_4092,N_4171);
and U4248 (N_4248,N_4192,N_4165);
nor U4249 (N_4249,N_4195,N_4027);
and U4250 (N_4250,N_4146,N_4083);
nor U4251 (N_4251,N_4064,N_4128);
or U4252 (N_4252,N_4053,N_4185);
nor U4253 (N_4253,N_4145,N_4003);
nand U4254 (N_4254,N_4182,N_4135);
nand U4255 (N_4255,N_4183,N_4071);
and U4256 (N_4256,N_4016,N_4062);
nand U4257 (N_4257,N_4054,N_4132);
nor U4258 (N_4258,N_4009,N_4199);
or U4259 (N_4259,N_4091,N_4130);
nor U4260 (N_4260,N_4114,N_4104);
nor U4261 (N_4261,N_4118,N_4001);
or U4262 (N_4262,N_4034,N_4081);
nor U4263 (N_4263,N_4164,N_4066);
nor U4264 (N_4264,N_4057,N_4033);
nand U4265 (N_4265,N_4176,N_4069);
nand U4266 (N_4266,N_4154,N_4193);
nand U4267 (N_4267,N_4039,N_4065);
nor U4268 (N_4268,N_4011,N_4052);
nor U4269 (N_4269,N_4040,N_4100);
nor U4270 (N_4270,N_4084,N_4068);
nor U4271 (N_4271,N_4099,N_4067);
and U4272 (N_4272,N_4139,N_4103);
and U4273 (N_4273,N_4129,N_4094);
and U4274 (N_4274,N_4048,N_4166);
or U4275 (N_4275,N_4031,N_4175);
or U4276 (N_4276,N_4060,N_4189);
or U4277 (N_4277,N_4051,N_4010);
nand U4278 (N_4278,N_4022,N_4136);
nand U4279 (N_4279,N_4025,N_4059);
nand U4280 (N_4280,N_4076,N_4115);
nor U4281 (N_4281,N_4163,N_4038);
and U4282 (N_4282,N_4138,N_4042);
nor U4283 (N_4283,N_4179,N_4151);
and U4284 (N_4284,N_4043,N_4106);
or U4285 (N_4285,N_4119,N_4050);
xor U4286 (N_4286,N_4168,N_4004);
nand U4287 (N_4287,N_4124,N_4055);
xnor U4288 (N_4288,N_4020,N_4191);
nor U4289 (N_4289,N_4095,N_4117);
nand U4290 (N_4290,N_4153,N_4173);
nand U4291 (N_4291,N_4174,N_4120);
nand U4292 (N_4292,N_4021,N_4133);
nor U4293 (N_4293,N_4046,N_4093);
nand U4294 (N_4294,N_4056,N_4141);
or U4295 (N_4295,N_4134,N_4024);
and U4296 (N_4296,N_4102,N_4126);
nand U4297 (N_4297,N_4088,N_4030);
nand U4298 (N_4298,N_4122,N_4079);
nor U4299 (N_4299,N_4008,N_4108);
xnor U4300 (N_4300,N_4086,N_4050);
or U4301 (N_4301,N_4175,N_4138);
and U4302 (N_4302,N_4110,N_4016);
and U4303 (N_4303,N_4094,N_4102);
nand U4304 (N_4304,N_4043,N_4089);
or U4305 (N_4305,N_4004,N_4012);
or U4306 (N_4306,N_4156,N_4143);
and U4307 (N_4307,N_4046,N_4156);
and U4308 (N_4308,N_4059,N_4162);
or U4309 (N_4309,N_4164,N_4128);
nand U4310 (N_4310,N_4122,N_4139);
and U4311 (N_4311,N_4005,N_4168);
or U4312 (N_4312,N_4086,N_4018);
nand U4313 (N_4313,N_4044,N_4195);
nor U4314 (N_4314,N_4163,N_4174);
nor U4315 (N_4315,N_4141,N_4134);
nor U4316 (N_4316,N_4015,N_4194);
nor U4317 (N_4317,N_4088,N_4032);
xor U4318 (N_4318,N_4121,N_4166);
or U4319 (N_4319,N_4059,N_4173);
nand U4320 (N_4320,N_4068,N_4128);
and U4321 (N_4321,N_4091,N_4028);
and U4322 (N_4322,N_4012,N_4040);
nor U4323 (N_4323,N_4024,N_4085);
or U4324 (N_4324,N_4096,N_4030);
and U4325 (N_4325,N_4165,N_4080);
and U4326 (N_4326,N_4085,N_4171);
xnor U4327 (N_4327,N_4121,N_4086);
or U4328 (N_4328,N_4162,N_4034);
nand U4329 (N_4329,N_4098,N_4103);
or U4330 (N_4330,N_4189,N_4165);
or U4331 (N_4331,N_4188,N_4076);
or U4332 (N_4332,N_4054,N_4031);
or U4333 (N_4333,N_4003,N_4064);
or U4334 (N_4334,N_4163,N_4063);
and U4335 (N_4335,N_4136,N_4033);
or U4336 (N_4336,N_4171,N_4134);
or U4337 (N_4337,N_4007,N_4132);
and U4338 (N_4338,N_4038,N_4059);
xor U4339 (N_4339,N_4098,N_4075);
nor U4340 (N_4340,N_4148,N_4070);
or U4341 (N_4341,N_4139,N_4127);
and U4342 (N_4342,N_4073,N_4088);
or U4343 (N_4343,N_4001,N_4190);
or U4344 (N_4344,N_4031,N_4014);
nand U4345 (N_4345,N_4076,N_4192);
nand U4346 (N_4346,N_4040,N_4131);
and U4347 (N_4347,N_4143,N_4104);
nand U4348 (N_4348,N_4194,N_4115);
and U4349 (N_4349,N_4111,N_4010);
nor U4350 (N_4350,N_4131,N_4013);
nor U4351 (N_4351,N_4197,N_4155);
or U4352 (N_4352,N_4042,N_4188);
and U4353 (N_4353,N_4003,N_4150);
nor U4354 (N_4354,N_4039,N_4071);
nor U4355 (N_4355,N_4141,N_4001);
nor U4356 (N_4356,N_4067,N_4136);
nand U4357 (N_4357,N_4173,N_4055);
nand U4358 (N_4358,N_4173,N_4031);
nand U4359 (N_4359,N_4141,N_4078);
and U4360 (N_4360,N_4130,N_4034);
and U4361 (N_4361,N_4168,N_4062);
xnor U4362 (N_4362,N_4013,N_4108);
or U4363 (N_4363,N_4066,N_4184);
nand U4364 (N_4364,N_4125,N_4164);
xnor U4365 (N_4365,N_4173,N_4050);
or U4366 (N_4366,N_4064,N_4026);
or U4367 (N_4367,N_4029,N_4002);
nor U4368 (N_4368,N_4103,N_4001);
nor U4369 (N_4369,N_4139,N_4111);
or U4370 (N_4370,N_4131,N_4018);
nor U4371 (N_4371,N_4158,N_4167);
and U4372 (N_4372,N_4153,N_4137);
nand U4373 (N_4373,N_4085,N_4082);
nand U4374 (N_4374,N_4027,N_4031);
or U4375 (N_4375,N_4034,N_4177);
nand U4376 (N_4376,N_4062,N_4097);
or U4377 (N_4377,N_4199,N_4032);
nand U4378 (N_4378,N_4053,N_4008);
nor U4379 (N_4379,N_4116,N_4081);
or U4380 (N_4380,N_4191,N_4143);
or U4381 (N_4381,N_4112,N_4127);
xnor U4382 (N_4382,N_4147,N_4038);
nor U4383 (N_4383,N_4181,N_4152);
or U4384 (N_4384,N_4058,N_4071);
or U4385 (N_4385,N_4013,N_4015);
nor U4386 (N_4386,N_4002,N_4075);
and U4387 (N_4387,N_4083,N_4135);
nor U4388 (N_4388,N_4062,N_4125);
or U4389 (N_4389,N_4185,N_4055);
or U4390 (N_4390,N_4028,N_4041);
nor U4391 (N_4391,N_4067,N_4131);
or U4392 (N_4392,N_4179,N_4146);
and U4393 (N_4393,N_4056,N_4170);
nor U4394 (N_4394,N_4027,N_4183);
nand U4395 (N_4395,N_4125,N_4095);
nand U4396 (N_4396,N_4162,N_4099);
and U4397 (N_4397,N_4134,N_4194);
or U4398 (N_4398,N_4136,N_4090);
nor U4399 (N_4399,N_4066,N_4068);
and U4400 (N_4400,N_4233,N_4387);
and U4401 (N_4401,N_4250,N_4211);
or U4402 (N_4402,N_4252,N_4321);
or U4403 (N_4403,N_4202,N_4208);
nand U4404 (N_4404,N_4254,N_4222);
nor U4405 (N_4405,N_4209,N_4299);
nor U4406 (N_4406,N_4324,N_4303);
and U4407 (N_4407,N_4337,N_4332);
nor U4408 (N_4408,N_4284,N_4291);
xor U4409 (N_4409,N_4357,N_4334);
or U4410 (N_4410,N_4226,N_4305);
nand U4411 (N_4411,N_4336,N_4393);
or U4412 (N_4412,N_4231,N_4281);
and U4413 (N_4413,N_4272,N_4280);
and U4414 (N_4414,N_4259,N_4388);
or U4415 (N_4415,N_4239,N_4282);
nand U4416 (N_4416,N_4374,N_4394);
nand U4417 (N_4417,N_4316,N_4382);
xor U4418 (N_4418,N_4359,N_4245);
or U4419 (N_4419,N_4351,N_4356);
nand U4420 (N_4420,N_4344,N_4224);
nor U4421 (N_4421,N_4318,N_4269);
or U4422 (N_4422,N_4215,N_4230);
nor U4423 (N_4423,N_4362,N_4327);
nand U4424 (N_4424,N_4273,N_4225);
and U4425 (N_4425,N_4341,N_4349);
and U4426 (N_4426,N_4360,N_4219);
or U4427 (N_4427,N_4329,N_4300);
xnor U4428 (N_4428,N_4377,N_4384);
and U4429 (N_4429,N_4277,N_4320);
nand U4430 (N_4430,N_4255,N_4256);
and U4431 (N_4431,N_4283,N_4307);
or U4432 (N_4432,N_4287,N_4237);
xor U4433 (N_4433,N_4368,N_4392);
and U4434 (N_4434,N_4375,N_4217);
and U4435 (N_4435,N_4385,N_4306);
and U4436 (N_4436,N_4353,N_4347);
xnor U4437 (N_4437,N_4348,N_4354);
or U4438 (N_4438,N_4240,N_4397);
and U4439 (N_4439,N_4396,N_4228);
nor U4440 (N_4440,N_4345,N_4270);
or U4441 (N_4441,N_4301,N_4298);
or U4442 (N_4442,N_4371,N_4263);
and U4443 (N_4443,N_4313,N_4232);
and U4444 (N_4444,N_4244,N_4220);
and U4445 (N_4445,N_4214,N_4361);
nand U4446 (N_4446,N_4285,N_4370);
or U4447 (N_4447,N_4248,N_4261);
nand U4448 (N_4448,N_4213,N_4204);
nor U4449 (N_4449,N_4363,N_4247);
and U4450 (N_4450,N_4381,N_4216);
nand U4451 (N_4451,N_4331,N_4258);
nor U4452 (N_4452,N_4367,N_4365);
and U4453 (N_4453,N_4358,N_4304);
nand U4454 (N_4454,N_4201,N_4235);
nor U4455 (N_4455,N_4319,N_4262);
nand U4456 (N_4456,N_4333,N_4257);
nand U4457 (N_4457,N_4205,N_4246);
xnor U4458 (N_4458,N_4203,N_4266);
and U4459 (N_4459,N_4340,N_4311);
nand U4460 (N_4460,N_4339,N_4352);
xnor U4461 (N_4461,N_4317,N_4379);
and U4462 (N_4462,N_4315,N_4293);
nor U4463 (N_4463,N_4200,N_4253);
or U4464 (N_4464,N_4391,N_4346);
nand U4465 (N_4465,N_4310,N_4227);
nor U4466 (N_4466,N_4288,N_4335);
nor U4467 (N_4467,N_4308,N_4229);
nand U4468 (N_4468,N_4274,N_4212);
or U4469 (N_4469,N_4390,N_4342);
or U4470 (N_4470,N_4312,N_4326);
and U4471 (N_4471,N_4265,N_4218);
xor U4472 (N_4472,N_4290,N_4323);
xor U4473 (N_4473,N_4395,N_4383);
and U4474 (N_4474,N_4289,N_4297);
and U4475 (N_4475,N_4242,N_4366);
and U4476 (N_4476,N_4236,N_4343);
or U4477 (N_4477,N_4221,N_4364);
nand U4478 (N_4478,N_4249,N_4292);
nand U4479 (N_4479,N_4398,N_4286);
nor U4480 (N_4480,N_4372,N_4223);
nor U4481 (N_4481,N_4275,N_4325);
and U4482 (N_4482,N_4243,N_4338);
nand U4483 (N_4483,N_4276,N_4241);
and U4484 (N_4484,N_4355,N_4260);
nand U4485 (N_4485,N_4302,N_4279);
or U4486 (N_4486,N_4267,N_4386);
nand U4487 (N_4487,N_4296,N_4350);
nor U4488 (N_4488,N_4309,N_4271);
and U4489 (N_4489,N_4210,N_4328);
or U4490 (N_4490,N_4380,N_4330);
xor U4491 (N_4491,N_4294,N_4278);
or U4492 (N_4492,N_4268,N_4369);
xnor U4493 (N_4493,N_4251,N_4399);
nand U4494 (N_4494,N_4314,N_4234);
and U4495 (N_4495,N_4389,N_4206);
or U4496 (N_4496,N_4378,N_4295);
and U4497 (N_4497,N_4373,N_4238);
nor U4498 (N_4498,N_4264,N_4322);
nor U4499 (N_4499,N_4376,N_4207);
and U4500 (N_4500,N_4365,N_4300);
nand U4501 (N_4501,N_4394,N_4316);
nor U4502 (N_4502,N_4342,N_4284);
nand U4503 (N_4503,N_4395,N_4306);
and U4504 (N_4504,N_4361,N_4261);
and U4505 (N_4505,N_4387,N_4281);
and U4506 (N_4506,N_4363,N_4303);
or U4507 (N_4507,N_4338,N_4341);
and U4508 (N_4508,N_4334,N_4356);
nand U4509 (N_4509,N_4218,N_4229);
and U4510 (N_4510,N_4319,N_4246);
nand U4511 (N_4511,N_4392,N_4366);
nor U4512 (N_4512,N_4363,N_4271);
and U4513 (N_4513,N_4368,N_4380);
xor U4514 (N_4514,N_4358,N_4336);
xor U4515 (N_4515,N_4321,N_4378);
and U4516 (N_4516,N_4232,N_4244);
nor U4517 (N_4517,N_4222,N_4305);
and U4518 (N_4518,N_4265,N_4305);
or U4519 (N_4519,N_4321,N_4208);
nor U4520 (N_4520,N_4397,N_4360);
and U4521 (N_4521,N_4320,N_4262);
nor U4522 (N_4522,N_4242,N_4391);
nor U4523 (N_4523,N_4311,N_4293);
and U4524 (N_4524,N_4364,N_4300);
nand U4525 (N_4525,N_4279,N_4356);
or U4526 (N_4526,N_4204,N_4327);
nor U4527 (N_4527,N_4284,N_4201);
nor U4528 (N_4528,N_4271,N_4303);
and U4529 (N_4529,N_4236,N_4388);
or U4530 (N_4530,N_4247,N_4394);
or U4531 (N_4531,N_4399,N_4278);
and U4532 (N_4532,N_4201,N_4368);
nand U4533 (N_4533,N_4378,N_4289);
nor U4534 (N_4534,N_4395,N_4380);
or U4535 (N_4535,N_4288,N_4298);
nor U4536 (N_4536,N_4326,N_4394);
and U4537 (N_4537,N_4223,N_4269);
and U4538 (N_4538,N_4257,N_4338);
and U4539 (N_4539,N_4264,N_4251);
or U4540 (N_4540,N_4344,N_4299);
xor U4541 (N_4541,N_4312,N_4221);
xor U4542 (N_4542,N_4375,N_4206);
and U4543 (N_4543,N_4378,N_4386);
nand U4544 (N_4544,N_4320,N_4202);
xnor U4545 (N_4545,N_4219,N_4350);
nor U4546 (N_4546,N_4211,N_4333);
or U4547 (N_4547,N_4352,N_4240);
and U4548 (N_4548,N_4301,N_4322);
nand U4549 (N_4549,N_4209,N_4382);
and U4550 (N_4550,N_4254,N_4286);
or U4551 (N_4551,N_4366,N_4294);
nand U4552 (N_4552,N_4263,N_4340);
and U4553 (N_4553,N_4240,N_4223);
nand U4554 (N_4554,N_4305,N_4254);
nor U4555 (N_4555,N_4323,N_4200);
and U4556 (N_4556,N_4292,N_4232);
nor U4557 (N_4557,N_4325,N_4304);
nor U4558 (N_4558,N_4243,N_4359);
or U4559 (N_4559,N_4275,N_4366);
and U4560 (N_4560,N_4226,N_4372);
nand U4561 (N_4561,N_4367,N_4386);
or U4562 (N_4562,N_4385,N_4378);
nand U4563 (N_4563,N_4248,N_4317);
and U4564 (N_4564,N_4234,N_4376);
or U4565 (N_4565,N_4368,N_4275);
nand U4566 (N_4566,N_4352,N_4227);
nand U4567 (N_4567,N_4221,N_4330);
nor U4568 (N_4568,N_4286,N_4368);
nand U4569 (N_4569,N_4371,N_4232);
nand U4570 (N_4570,N_4368,N_4383);
nor U4571 (N_4571,N_4368,N_4336);
or U4572 (N_4572,N_4284,N_4356);
or U4573 (N_4573,N_4238,N_4257);
nand U4574 (N_4574,N_4340,N_4348);
and U4575 (N_4575,N_4253,N_4204);
and U4576 (N_4576,N_4312,N_4314);
nor U4577 (N_4577,N_4298,N_4332);
nand U4578 (N_4578,N_4388,N_4209);
nand U4579 (N_4579,N_4287,N_4306);
or U4580 (N_4580,N_4243,N_4309);
or U4581 (N_4581,N_4375,N_4377);
xnor U4582 (N_4582,N_4382,N_4330);
or U4583 (N_4583,N_4357,N_4258);
nand U4584 (N_4584,N_4361,N_4201);
or U4585 (N_4585,N_4371,N_4349);
or U4586 (N_4586,N_4381,N_4212);
nand U4587 (N_4587,N_4329,N_4341);
nand U4588 (N_4588,N_4364,N_4290);
and U4589 (N_4589,N_4394,N_4343);
and U4590 (N_4590,N_4281,N_4389);
nand U4591 (N_4591,N_4365,N_4204);
and U4592 (N_4592,N_4286,N_4285);
nor U4593 (N_4593,N_4200,N_4229);
or U4594 (N_4594,N_4359,N_4389);
and U4595 (N_4595,N_4250,N_4226);
or U4596 (N_4596,N_4330,N_4242);
nand U4597 (N_4597,N_4238,N_4366);
or U4598 (N_4598,N_4295,N_4201);
xor U4599 (N_4599,N_4221,N_4339);
and U4600 (N_4600,N_4557,N_4594);
and U4601 (N_4601,N_4488,N_4511);
or U4602 (N_4602,N_4560,N_4415);
or U4603 (N_4603,N_4521,N_4548);
nand U4604 (N_4604,N_4501,N_4570);
and U4605 (N_4605,N_4582,N_4485);
and U4606 (N_4606,N_4470,N_4430);
xnor U4607 (N_4607,N_4536,N_4425);
xor U4608 (N_4608,N_4450,N_4418);
and U4609 (N_4609,N_4503,N_4432);
nor U4610 (N_4610,N_4481,N_4408);
nor U4611 (N_4611,N_4522,N_4444);
and U4612 (N_4612,N_4553,N_4471);
nand U4613 (N_4613,N_4585,N_4437);
and U4614 (N_4614,N_4498,N_4458);
or U4615 (N_4615,N_4568,N_4545);
nor U4616 (N_4616,N_4475,N_4480);
and U4617 (N_4617,N_4505,N_4493);
and U4618 (N_4618,N_4581,N_4530);
nor U4619 (N_4619,N_4452,N_4448);
or U4620 (N_4620,N_4526,N_4517);
or U4621 (N_4621,N_4416,N_4589);
nor U4622 (N_4622,N_4479,N_4424);
and U4623 (N_4623,N_4463,N_4457);
or U4624 (N_4624,N_4532,N_4518);
nand U4625 (N_4625,N_4510,N_4461);
xnor U4626 (N_4626,N_4549,N_4588);
or U4627 (N_4627,N_4508,N_4476);
nand U4628 (N_4628,N_4519,N_4593);
and U4629 (N_4629,N_4514,N_4564);
nor U4630 (N_4630,N_4591,N_4486);
or U4631 (N_4631,N_4576,N_4406);
or U4632 (N_4632,N_4421,N_4489);
nand U4633 (N_4633,N_4523,N_4410);
nor U4634 (N_4634,N_4401,N_4567);
and U4635 (N_4635,N_4512,N_4573);
and U4636 (N_4636,N_4419,N_4533);
xnor U4637 (N_4637,N_4469,N_4453);
xor U4638 (N_4638,N_4537,N_4596);
nor U4639 (N_4639,N_4451,N_4467);
or U4640 (N_4640,N_4566,N_4525);
and U4641 (N_4641,N_4500,N_4482);
and U4642 (N_4642,N_4506,N_4414);
and U4643 (N_4643,N_4527,N_4590);
nor U4644 (N_4644,N_4428,N_4413);
nand U4645 (N_4645,N_4587,N_4539);
and U4646 (N_4646,N_4561,N_4562);
or U4647 (N_4647,N_4455,N_4595);
and U4648 (N_4648,N_4447,N_4487);
or U4649 (N_4649,N_4534,N_4563);
or U4650 (N_4650,N_4565,N_4528);
nand U4651 (N_4651,N_4550,N_4541);
and U4652 (N_4652,N_4520,N_4438);
and U4653 (N_4653,N_4547,N_4441);
and U4654 (N_4654,N_4551,N_4572);
xor U4655 (N_4655,N_4507,N_4509);
nand U4656 (N_4656,N_4423,N_4446);
and U4657 (N_4657,N_4569,N_4409);
nor U4658 (N_4658,N_4578,N_4478);
and U4659 (N_4659,N_4542,N_4577);
and U4660 (N_4660,N_4449,N_4599);
and U4661 (N_4661,N_4504,N_4554);
and U4662 (N_4662,N_4427,N_4556);
xor U4663 (N_4663,N_4442,N_4473);
and U4664 (N_4664,N_4496,N_4460);
and U4665 (N_4665,N_4559,N_4580);
and U4666 (N_4666,N_4484,N_4574);
and U4667 (N_4667,N_4544,N_4490);
xnor U4668 (N_4668,N_4492,N_4495);
nor U4669 (N_4669,N_4404,N_4417);
nand U4670 (N_4670,N_4497,N_4405);
nand U4671 (N_4671,N_4538,N_4454);
nand U4672 (N_4672,N_4435,N_4529);
and U4673 (N_4673,N_4597,N_4472);
nor U4674 (N_4674,N_4494,N_4400);
nor U4675 (N_4675,N_4513,N_4402);
and U4676 (N_4676,N_4422,N_4403);
or U4677 (N_4677,N_4477,N_4439);
or U4678 (N_4678,N_4462,N_4468);
or U4679 (N_4679,N_4445,N_4426);
xor U4680 (N_4680,N_4502,N_4440);
nand U4681 (N_4681,N_4584,N_4552);
xnor U4682 (N_4682,N_4466,N_4546);
or U4683 (N_4683,N_4433,N_4555);
and U4684 (N_4684,N_4558,N_4459);
nor U4685 (N_4685,N_4515,N_4575);
and U4686 (N_4686,N_4598,N_4491);
nand U4687 (N_4687,N_4434,N_4540);
nor U4688 (N_4688,N_4571,N_4579);
and U4689 (N_4689,N_4524,N_4583);
nor U4690 (N_4690,N_4411,N_4464);
nor U4691 (N_4691,N_4483,N_4543);
xor U4692 (N_4692,N_4592,N_4465);
nor U4693 (N_4693,N_4474,N_4412);
or U4694 (N_4694,N_4420,N_4456);
xor U4695 (N_4695,N_4499,N_4586);
xnor U4696 (N_4696,N_4443,N_4531);
and U4697 (N_4697,N_4407,N_4431);
or U4698 (N_4698,N_4535,N_4436);
nor U4699 (N_4699,N_4516,N_4429);
nand U4700 (N_4700,N_4465,N_4402);
or U4701 (N_4701,N_4587,N_4471);
and U4702 (N_4702,N_4480,N_4416);
nor U4703 (N_4703,N_4403,N_4440);
xor U4704 (N_4704,N_4557,N_4597);
and U4705 (N_4705,N_4514,N_4544);
nand U4706 (N_4706,N_4529,N_4546);
nand U4707 (N_4707,N_4598,N_4588);
and U4708 (N_4708,N_4462,N_4467);
nand U4709 (N_4709,N_4586,N_4496);
or U4710 (N_4710,N_4578,N_4486);
nor U4711 (N_4711,N_4594,N_4552);
nor U4712 (N_4712,N_4513,N_4485);
or U4713 (N_4713,N_4406,N_4428);
and U4714 (N_4714,N_4504,N_4541);
xnor U4715 (N_4715,N_4464,N_4597);
nand U4716 (N_4716,N_4576,N_4533);
or U4717 (N_4717,N_4540,N_4508);
or U4718 (N_4718,N_4511,N_4401);
nand U4719 (N_4719,N_4411,N_4483);
nor U4720 (N_4720,N_4536,N_4581);
nand U4721 (N_4721,N_4579,N_4582);
and U4722 (N_4722,N_4415,N_4563);
nand U4723 (N_4723,N_4448,N_4409);
or U4724 (N_4724,N_4574,N_4567);
or U4725 (N_4725,N_4436,N_4493);
and U4726 (N_4726,N_4406,N_4540);
or U4727 (N_4727,N_4587,N_4485);
nor U4728 (N_4728,N_4594,N_4472);
and U4729 (N_4729,N_4546,N_4576);
and U4730 (N_4730,N_4406,N_4505);
nand U4731 (N_4731,N_4582,N_4446);
nand U4732 (N_4732,N_4530,N_4564);
nand U4733 (N_4733,N_4588,N_4446);
xor U4734 (N_4734,N_4424,N_4495);
nand U4735 (N_4735,N_4514,N_4541);
or U4736 (N_4736,N_4548,N_4583);
nand U4737 (N_4737,N_4510,N_4579);
and U4738 (N_4738,N_4566,N_4477);
nor U4739 (N_4739,N_4443,N_4480);
and U4740 (N_4740,N_4474,N_4506);
nor U4741 (N_4741,N_4502,N_4491);
xor U4742 (N_4742,N_4599,N_4426);
nand U4743 (N_4743,N_4404,N_4513);
nor U4744 (N_4744,N_4529,N_4434);
nor U4745 (N_4745,N_4593,N_4599);
or U4746 (N_4746,N_4571,N_4442);
and U4747 (N_4747,N_4453,N_4417);
and U4748 (N_4748,N_4412,N_4480);
or U4749 (N_4749,N_4518,N_4576);
nand U4750 (N_4750,N_4413,N_4583);
nor U4751 (N_4751,N_4412,N_4453);
or U4752 (N_4752,N_4552,N_4448);
nor U4753 (N_4753,N_4566,N_4453);
nand U4754 (N_4754,N_4455,N_4514);
and U4755 (N_4755,N_4532,N_4579);
xnor U4756 (N_4756,N_4433,N_4422);
xnor U4757 (N_4757,N_4593,N_4412);
and U4758 (N_4758,N_4455,N_4587);
or U4759 (N_4759,N_4548,N_4516);
and U4760 (N_4760,N_4580,N_4572);
nand U4761 (N_4761,N_4537,N_4536);
or U4762 (N_4762,N_4509,N_4568);
nand U4763 (N_4763,N_4557,N_4516);
and U4764 (N_4764,N_4509,N_4574);
or U4765 (N_4765,N_4552,N_4572);
nand U4766 (N_4766,N_4444,N_4591);
nor U4767 (N_4767,N_4577,N_4468);
or U4768 (N_4768,N_4425,N_4401);
and U4769 (N_4769,N_4452,N_4480);
nand U4770 (N_4770,N_4407,N_4424);
or U4771 (N_4771,N_4572,N_4447);
nand U4772 (N_4772,N_4501,N_4557);
or U4773 (N_4773,N_4597,N_4429);
and U4774 (N_4774,N_4535,N_4457);
and U4775 (N_4775,N_4569,N_4429);
and U4776 (N_4776,N_4508,N_4425);
xnor U4777 (N_4777,N_4565,N_4449);
and U4778 (N_4778,N_4440,N_4457);
nand U4779 (N_4779,N_4501,N_4432);
and U4780 (N_4780,N_4552,N_4538);
nor U4781 (N_4781,N_4446,N_4506);
and U4782 (N_4782,N_4597,N_4475);
nor U4783 (N_4783,N_4455,N_4464);
and U4784 (N_4784,N_4488,N_4507);
or U4785 (N_4785,N_4475,N_4464);
and U4786 (N_4786,N_4531,N_4540);
xor U4787 (N_4787,N_4573,N_4414);
nand U4788 (N_4788,N_4513,N_4470);
nand U4789 (N_4789,N_4420,N_4550);
or U4790 (N_4790,N_4476,N_4550);
nand U4791 (N_4791,N_4576,N_4499);
nand U4792 (N_4792,N_4407,N_4551);
and U4793 (N_4793,N_4487,N_4506);
nor U4794 (N_4794,N_4435,N_4423);
nand U4795 (N_4795,N_4558,N_4472);
and U4796 (N_4796,N_4472,N_4484);
nand U4797 (N_4797,N_4432,N_4472);
and U4798 (N_4798,N_4491,N_4501);
and U4799 (N_4799,N_4434,N_4417);
nand U4800 (N_4800,N_4725,N_4772);
or U4801 (N_4801,N_4705,N_4697);
nor U4802 (N_4802,N_4632,N_4634);
and U4803 (N_4803,N_4774,N_4761);
nand U4804 (N_4804,N_4680,N_4733);
or U4805 (N_4805,N_4780,N_4678);
or U4806 (N_4806,N_4721,N_4650);
nor U4807 (N_4807,N_4645,N_4676);
xnor U4808 (N_4808,N_4717,N_4627);
nand U4809 (N_4809,N_4698,N_4703);
xnor U4810 (N_4810,N_4699,N_4769);
nand U4811 (N_4811,N_4667,N_4601);
nor U4812 (N_4812,N_4784,N_4706);
xnor U4813 (N_4813,N_4791,N_4639);
nand U4814 (N_4814,N_4630,N_4765);
and U4815 (N_4815,N_4600,N_4677);
nor U4816 (N_4816,N_4716,N_4607);
or U4817 (N_4817,N_4685,N_4662);
and U4818 (N_4818,N_4798,N_4665);
and U4819 (N_4819,N_4760,N_4658);
xor U4820 (N_4820,N_4776,N_4758);
or U4821 (N_4821,N_4693,N_4731);
or U4822 (N_4822,N_4711,N_4694);
and U4823 (N_4823,N_4686,N_4747);
and U4824 (N_4824,N_4740,N_4738);
or U4825 (N_4825,N_4604,N_4709);
and U4826 (N_4826,N_4787,N_4696);
and U4827 (N_4827,N_4622,N_4771);
and U4828 (N_4828,N_4628,N_4666);
and U4829 (N_4829,N_4661,N_4657);
nor U4830 (N_4830,N_4736,N_4644);
and U4831 (N_4831,N_4757,N_4767);
or U4832 (N_4832,N_4663,N_4766);
xnor U4833 (N_4833,N_4633,N_4718);
nand U4834 (N_4834,N_4789,N_4602);
or U4835 (N_4835,N_4681,N_4742);
and U4836 (N_4836,N_4625,N_4669);
nor U4837 (N_4837,N_4701,N_4750);
or U4838 (N_4838,N_4689,N_4673);
or U4839 (N_4839,N_4682,N_4660);
nor U4840 (N_4840,N_4623,N_4744);
nand U4841 (N_4841,N_4732,N_4704);
nand U4842 (N_4842,N_4668,N_4754);
or U4843 (N_4843,N_4722,N_4752);
or U4844 (N_4844,N_4656,N_4653);
and U4845 (N_4845,N_4786,N_4788);
and U4846 (N_4846,N_4618,N_4683);
and U4847 (N_4847,N_4641,N_4692);
and U4848 (N_4848,N_4664,N_4794);
and U4849 (N_4849,N_4640,N_4652);
nor U4850 (N_4850,N_4715,N_4700);
nor U4851 (N_4851,N_4615,N_4672);
nor U4852 (N_4852,N_4755,N_4726);
xor U4853 (N_4853,N_4624,N_4714);
and U4854 (N_4854,N_4734,N_4720);
or U4855 (N_4855,N_4708,N_4603);
xor U4856 (N_4856,N_4614,N_4647);
and U4857 (N_4857,N_4759,N_4783);
or U4858 (N_4858,N_4728,N_4764);
nand U4859 (N_4859,N_4773,N_4775);
and U4860 (N_4860,N_4671,N_4636);
or U4861 (N_4861,N_4629,N_4620);
nor U4862 (N_4862,N_4631,N_4749);
nor U4863 (N_4863,N_4710,N_4730);
nand U4864 (N_4864,N_4702,N_4611);
and U4865 (N_4865,N_4610,N_4638);
or U4866 (N_4866,N_4690,N_4687);
nor U4867 (N_4867,N_4763,N_4617);
or U4868 (N_4868,N_4727,N_4743);
and U4869 (N_4869,N_4659,N_4635);
or U4870 (N_4870,N_4621,N_4608);
or U4871 (N_4871,N_4762,N_4790);
nand U4872 (N_4872,N_4713,N_4792);
nand U4873 (N_4873,N_4719,N_4712);
or U4874 (N_4874,N_4735,N_4648);
nand U4875 (N_4875,N_4651,N_4748);
and U4876 (N_4876,N_4684,N_4654);
or U4877 (N_4877,N_4751,N_4670);
and U4878 (N_4878,N_4679,N_4777);
and U4879 (N_4879,N_4729,N_4655);
nand U4880 (N_4880,N_4723,N_4741);
nand U4881 (N_4881,N_4675,N_4753);
xnor U4882 (N_4882,N_4612,N_4707);
nor U4883 (N_4883,N_4785,N_4781);
and U4884 (N_4884,N_4779,N_4626);
or U4885 (N_4885,N_4770,N_4695);
and U4886 (N_4886,N_4674,N_4605);
nor U4887 (N_4887,N_4616,N_4619);
nand U4888 (N_4888,N_4756,N_4739);
nand U4889 (N_4889,N_4799,N_4745);
and U4890 (N_4890,N_4795,N_4609);
xor U4891 (N_4891,N_4724,N_4746);
nand U4892 (N_4892,N_4737,N_4643);
or U4893 (N_4893,N_4793,N_4637);
and U4894 (N_4894,N_4606,N_4642);
nor U4895 (N_4895,N_4649,N_4778);
or U4896 (N_4896,N_4797,N_4688);
or U4897 (N_4897,N_4613,N_4796);
or U4898 (N_4898,N_4691,N_4646);
nor U4899 (N_4899,N_4782,N_4768);
nor U4900 (N_4900,N_4679,N_4677);
nand U4901 (N_4901,N_4720,N_4660);
or U4902 (N_4902,N_4725,N_4732);
or U4903 (N_4903,N_4795,N_4633);
nor U4904 (N_4904,N_4760,N_4731);
and U4905 (N_4905,N_4734,N_4731);
xnor U4906 (N_4906,N_4661,N_4635);
and U4907 (N_4907,N_4757,N_4768);
nor U4908 (N_4908,N_4717,N_4728);
or U4909 (N_4909,N_4664,N_4752);
or U4910 (N_4910,N_4756,N_4684);
or U4911 (N_4911,N_4717,N_4605);
or U4912 (N_4912,N_4616,N_4721);
xnor U4913 (N_4913,N_4618,N_4696);
and U4914 (N_4914,N_4615,N_4688);
nor U4915 (N_4915,N_4614,N_4666);
xnor U4916 (N_4916,N_4704,N_4757);
nand U4917 (N_4917,N_4615,N_4705);
xor U4918 (N_4918,N_4641,N_4607);
and U4919 (N_4919,N_4691,N_4639);
and U4920 (N_4920,N_4763,N_4722);
nor U4921 (N_4921,N_4796,N_4742);
or U4922 (N_4922,N_4795,N_4780);
nand U4923 (N_4923,N_4619,N_4770);
and U4924 (N_4924,N_4741,N_4677);
and U4925 (N_4925,N_4719,N_4741);
or U4926 (N_4926,N_4642,N_4629);
nand U4927 (N_4927,N_4651,N_4650);
nand U4928 (N_4928,N_4628,N_4611);
or U4929 (N_4929,N_4641,N_4749);
nand U4930 (N_4930,N_4724,N_4659);
and U4931 (N_4931,N_4766,N_4671);
nand U4932 (N_4932,N_4724,N_4747);
xor U4933 (N_4933,N_4641,N_4798);
or U4934 (N_4934,N_4729,N_4777);
or U4935 (N_4935,N_4737,N_4727);
nor U4936 (N_4936,N_4764,N_4788);
nor U4937 (N_4937,N_4606,N_4686);
nand U4938 (N_4938,N_4632,N_4742);
and U4939 (N_4939,N_4774,N_4770);
or U4940 (N_4940,N_4689,N_4724);
xor U4941 (N_4941,N_4784,N_4788);
and U4942 (N_4942,N_4771,N_4695);
nand U4943 (N_4943,N_4692,N_4615);
and U4944 (N_4944,N_4730,N_4775);
nor U4945 (N_4945,N_4766,N_4694);
xnor U4946 (N_4946,N_4717,N_4673);
nand U4947 (N_4947,N_4660,N_4755);
xor U4948 (N_4948,N_4765,N_4700);
nor U4949 (N_4949,N_4797,N_4606);
nor U4950 (N_4950,N_4722,N_4644);
nor U4951 (N_4951,N_4641,N_4600);
and U4952 (N_4952,N_4735,N_4677);
or U4953 (N_4953,N_4633,N_4717);
or U4954 (N_4954,N_4626,N_4785);
xor U4955 (N_4955,N_4765,N_4729);
and U4956 (N_4956,N_4684,N_4607);
and U4957 (N_4957,N_4718,N_4642);
nand U4958 (N_4958,N_4737,N_4648);
nor U4959 (N_4959,N_4622,N_4603);
or U4960 (N_4960,N_4626,N_4655);
and U4961 (N_4961,N_4736,N_4689);
nand U4962 (N_4962,N_4657,N_4651);
and U4963 (N_4963,N_4635,N_4753);
nand U4964 (N_4964,N_4602,N_4778);
and U4965 (N_4965,N_4673,N_4790);
nand U4966 (N_4966,N_4620,N_4787);
xor U4967 (N_4967,N_4613,N_4793);
nor U4968 (N_4968,N_4641,N_4737);
xnor U4969 (N_4969,N_4743,N_4631);
nand U4970 (N_4970,N_4629,N_4767);
nand U4971 (N_4971,N_4731,N_4755);
or U4972 (N_4972,N_4706,N_4660);
nand U4973 (N_4973,N_4709,N_4767);
nand U4974 (N_4974,N_4723,N_4622);
and U4975 (N_4975,N_4664,N_4726);
and U4976 (N_4976,N_4773,N_4618);
or U4977 (N_4977,N_4644,N_4709);
nor U4978 (N_4978,N_4698,N_4792);
or U4979 (N_4979,N_4604,N_4661);
nor U4980 (N_4980,N_4780,N_4700);
nand U4981 (N_4981,N_4650,N_4626);
nor U4982 (N_4982,N_4668,N_4650);
and U4983 (N_4983,N_4726,N_4605);
and U4984 (N_4984,N_4794,N_4648);
xor U4985 (N_4985,N_4692,N_4732);
nor U4986 (N_4986,N_4729,N_4744);
nor U4987 (N_4987,N_4777,N_4668);
nand U4988 (N_4988,N_4784,N_4713);
or U4989 (N_4989,N_4613,N_4650);
and U4990 (N_4990,N_4761,N_4625);
nor U4991 (N_4991,N_4708,N_4709);
or U4992 (N_4992,N_4666,N_4635);
and U4993 (N_4993,N_4731,N_4748);
nor U4994 (N_4994,N_4653,N_4797);
nor U4995 (N_4995,N_4621,N_4750);
nand U4996 (N_4996,N_4691,N_4722);
or U4997 (N_4997,N_4699,N_4752);
xor U4998 (N_4998,N_4713,N_4633);
nand U4999 (N_4999,N_4623,N_4726);
and U5000 (N_5000,N_4938,N_4905);
and U5001 (N_5001,N_4870,N_4858);
and U5002 (N_5002,N_4990,N_4881);
nand U5003 (N_5003,N_4878,N_4963);
and U5004 (N_5004,N_4898,N_4959);
nand U5005 (N_5005,N_4843,N_4912);
nand U5006 (N_5006,N_4889,N_4901);
nand U5007 (N_5007,N_4880,N_4997);
nor U5008 (N_5008,N_4874,N_4929);
nor U5009 (N_5009,N_4988,N_4975);
nor U5010 (N_5010,N_4926,N_4810);
or U5011 (N_5011,N_4869,N_4845);
or U5012 (N_5012,N_4834,N_4882);
nor U5013 (N_5013,N_4921,N_4837);
or U5014 (N_5014,N_4925,N_4839);
or U5015 (N_5015,N_4978,N_4814);
nand U5016 (N_5016,N_4866,N_4983);
and U5017 (N_5017,N_4941,N_4893);
xor U5018 (N_5018,N_4856,N_4977);
and U5019 (N_5019,N_4826,N_4917);
nor U5020 (N_5020,N_4823,N_4920);
nor U5021 (N_5021,N_4969,N_4999);
or U5022 (N_5022,N_4935,N_4993);
and U5023 (N_5023,N_4800,N_4821);
nand U5024 (N_5024,N_4867,N_4960);
nor U5025 (N_5025,N_4994,N_4918);
nor U5026 (N_5026,N_4970,N_4954);
nor U5027 (N_5027,N_4952,N_4979);
nor U5028 (N_5028,N_4853,N_4903);
nor U5029 (N_5029,N_4808,N_4916);
nor U5030 (N_5030,N_4884,N_4961);
and U5031 (N_5031,N_4896,N_4817);
xor U5032 (N_5032,N_4995,N_4827);
and U5033 (N_5033,N_4863,N_4982);
nor U5034 (N_5034,N_4847,N_4949);
nor U5035 (N_5035,N_4980,N_4849);
nor U5036 (N_5036,N_4965,N_4985);
or U5037 (N_5037,N_4865,N_4908);
and U5038 (N_5038,N_4820,N_4835);
or U5039 (N_5039,N_4859,N_4976);
or U5040 (N_5040,N_4934,N_4840);
or U5041 (N_5041,N_4887,N_4940);
nand U5042 (N_5042,N_4996,N_4836);
nor U5043 (N_5043,N_4950,N_4933);
or U5044 (N_5044,N_4894,N_4939);
nor U5045 (N_5045,N_4850,N_4822);
or U5046 (N_5046,N_4953,N_4928);
or U5047 (N_5047,N_4875,N_4832);
or U5048 (N_5048,N_4981,N_4915);
or U5049 (N_5049,N_4909,N_4913);
and U5050 (N_5050,N_4992,N_4809);
and U5051 (N_5051,N_4966,N_4904);
nand U5052 (N_5052,N_4973,N_4911);
nand U5053 (N_5053,N_4816,N_4892);
nor U5054 (N_5054,N_4919,N_4824);
nor U5055 (N_5055,N_4885,N_4806);
and U5056 (N_5056,N_4924,N_4900);
nand U5057 (N_5057,N_4956,N_4937);
xnor U5058 (N_5058,N_4944,N_4895);
or U5059 (N_5059,N_4931,N_4812);
nand U5060 (N_5060,N_4968,N_4890);
or U5061 (N_5061,N_4828,N_4852);
nor U5062 (N_5062,N_4801,N_4802);
or U5063 (N_5063,N_4833,N_4972);
nand U5064 (N_5064,N_4811,N_4902);
nor U5065 (N_5065,N_4842,N_4910);
and U5066 (N_5066,N_4948,N_4971);
or U5067 (N_5067,N_4803,N_4838);
nand U5068 (N_5068,N_4888,N_4897);
or U5069 (N_5069,N_4964,N_4805);
nor U5070 (N_5070,N_4804,N_4922);
or U5071 (N_5071,N_4958,N_4942);
or U5072 (N_5072,N_4848,N_4923);
and U5073 (N_5073,N_4989,N_4857);
nand U5074 (N_5074,N_4914,N_4936);
and U5075 (N_5075,N_4830,N_4861);
nor U5076 (N_5076,N_4955,N_4932);
and U5077 (N_5077,N_4855,N_4851);
or U5078 (N_5078,N_4951,N_4871);
nand U5079 (N_5079,N_4876,N_4813);
and U5080 (N_5080,N_4860,N_4883);
or U5081 (N_5081,N_4907,N_4946);
nand U5082 (N_5082,N_4962,N_4877);
or U5083 (N_5083,N_4815,N_4967);
and U5084 (N_5084,N_4868,N_4886);
and U5085 (N_5085,N_4986,N_4807);
and U5086 (N_5086,N_4974,N_4829);
nor U5087 (N_5087,N_4947,N_4987);
or U5088 (N_5088,N_4984,N_4998);
nor U5089 (N_5089,N_4872,N_4846);
and U5090 (N_5090,N_4831,N_4945);
xnor U5091 (N_5091,N_4906,N_4891);
nor U5092 (N_5092,N_4825,N_4862);
and U5093 (N_5093,N_4818,N_4943);
nand U5094 (N_5094,N_4930,N_4819);
nor U5095 (N_5095,N_4873,N_4927);
nor U5096 (N_5096,N_4854,N_4841);
and U5097 (N_5097,N_4991,N_4844);
nor U5098 (N_5098,N_4879,N_4864);
or U5099 (N_5099,N_4957,N_4899);
nand U5100 (N_5100,N_4812,N_4875);
xnor U5101 (N_5101,N_4830,N_4933);
and U5102 (N_5102,N_4966,N_4802);
nor U5103 (N_5103,N_4930,N_4978);
nor U5104 (N_5104,N_4871,N_4973);
and U5105 (N_5105,N_4834,N_4842);
and U5106 (N_5106,N_4828,N_4881);
and U5107 (N_5107,N_4905,N_4993);
and U5108 (N_5108,N_4907,N_4882);
nor U5109 (N_5109,N_4903,N_4840);
and U5110 (N_5110,N_4823,N_4953);
and U5111 (N_5111,N_4950,N_4965);
or U5112 (N_5112,N_4861,N_4804);
nor U5113 (N_5113,N_4928,N_4974);
and U5114 (N_5114,N_4894,N_4901);
nor U5115 (N_5115,N_4998,N_4845);
xor U5116 (N_5116,N_4862,N_4913);
and U5117 (N_5117,N_4800,N_4987);
and U5118 (N_5118,N_4866,N_4913);
xor U5119 (N_5119,N_4973,N_4828);
or U5120 (N_5120,N_4858,N_4952);
and U5121 (N_5121,N_4866,N_4973);
nand U5122 (N_5122,N_4905,N_4992);
nand U5123 (N_5123,N_4869,N_4848);
and U5124 (N_5124,N_4849,N_4957);
nor U5125 (N_5125,N_4938,N_4800);
nor U5126 (N_5126,N_4806,N_4816);
xnor U5127 (N_5127,N_4896,N_4987);
xor U5128 (N_5128,N_4957,N_4883);
nand U5129 (N_5129,N_4818,N_4804);
nand U5130 (N_5130,N_4968,N_4962);
and U5131 (N_5131,N_4831,N_4829);
nand U5132 (N_5132,N_4860,N_4892);
nand U5133 (N_5133,N_4832,N_4846);
nor U5134 (N_5134,N_4916,N_4957);
xor U5135 (N_5135,N_4921,N_4826);
or U5136 (N_5136,N_4805,N_4991);
or U5137 (N_5137,N_4973,N_4819);
or U5138 (N_5138,N_4897,N_4898);
nand U5139 (N_5139,N_4961,N_4993);
or U5140 (N_5140,N_4964,N_4982);
and U5141 (N_5141,N_4931,N_4935);
nand U5142 (N_5142,N_4804,N_4908);
nand U5143 (N_5143,N_4848,N_4872);
or U5144 (N_5144,N_4910,N_4803);
and U5145 (N_5145,N_4910,N_4801);
and U5146 (N_5146,N_4952,N_4947);
and U5147 (N_5147,N_4868,N_4822);
xor U5148 (N_5148,N_4874,N_4828);
or U5149 (N_5149,N_4849,N_4973);
xnor U5150 (N_5150,N_4801,N_4884);
and U5151 (N_5151,N_4970,N_4941);
xnor U5152 (N_5152,N_4878,N_4996);
and U5153 (N_5153,N_4930,N_4807);
nor U5154 (N_5154,N_4927,N_4989);
xor U5155 (N_5155,N_4812,N_4973);
xor U5156 (N_5156,N_4922,N_4984);
xnor U5157 (N_5157,N_4862,N_4919);
nand U5158 (N_5158,N_4871,N_4947);
or U5159 (N_5159,N_4812,N_4835);
nor U5160 (N_5160,N_4920,N_4839);
or U5161 (N_5161,N_4952,N_4804);
and U5162 (N_5162,N_4925,N_4947);
nor U5163 (N_5163,N_4891,N_4986);
nor U5164 (N_5164,N_4855,N_4991);
nor U5165 (N_5165,N_4816,N_4921);
nor U5166 (N_5166,N_4978,N_4969);
xnor U5167 (N_5167,N_4904,N_4873);
nand U5168 (N_5168,N_4941,N_4852);
nand U5169 (N_5169,N_4968,N_4927);
nor U5170 (N_5170,N_4973,N_4964);
or U5171 (N_5171,N_4875,N_4904);
nand U5172 (N_5172,N_4989,N_4884);
nor U5173 (N_5173,N_4807,N_4999);
and U5174 (N_5174,N_4990,N_4895);
xnor U5175 (N_5175,N_4949,N_4939);
and U5176 (N_5176,N_4930,N_4881);
or U5177 (N_5177,N_4847,N_4971);
xor U5178 (N_5178,N_4907,N_4856);
and U5179 (N_5179,N_4826,N_4893);
or U5180 (N_5180,N_4940,N_4847);
and U5181 (N_5181,N_4812,N_4936);
nor U5182 (N_5182,N_4893,N_4951);
nor U5183 (N_5183,N_4877,N_4955);
nand U5184 (N_5184,N_4999,N_4979);
nor U5185 (N_5185,N_4876,N_4856);
and U5186 (N_5186,N_4878,N_4889);
nor U5187 (N_5187,N_4980,N_4868);
and U5188 (N_5188,N_4950,N_4898);
or U5189 (N_5189,N_4806,N_4912);
xor U5190 (N_5190,N_4894,N_4968);
nor U5191 (N_5191,N_4940,N_4914);
and U5192 (N_5192,N_4851,N_4828);
nor U5193 (N_5193,N_4836,N_4989);
or U5194 (N_5194,N_4849,N_4974);
nor U5195 (N_5195,N_4880,N_4946);
or U5196 (N_5196,N_4805,N_4949);
or U5197 (N_5197,N_4807,N_4924);
or U5198 (N_5198,N_4976,N_4868);
xor U5199 (N_5199,N_4883,N_4822);
nor U5200 (N_5200,N_5046,N_5188);
or U5201 (N_5201,N_5048,N_5158);
or U5202 (N_5202,N_5053,N_5164);
xor U5203 (N_5203,N_5161,N_5022);
nor U5204 (N_5204,N_5075,N_5185);
and U5205 (N_5205,N_5043,N_5124);
or U5206 (N_5206,N_5119,N_5165);
nor U5207 (N_5207,N_5105,N_5091);
or U5208 (N_5208,N_5088,N_5147);
and U5209 (N_5209,N_5171,N_5100);
nor U5210 (N_5210,N_5012,N_5107);
or U5211 (N_5211,N_5047,N_5057);
and U5212 (N_5212,N_5019,N_5156);
nand U5213 (N_5213,N_5140,N_5112);
or U5214 (N_5214,N_5077,N_5060);
nand U5215 (N_5215,N_5086,N_5170);
nand U5216 (N_5216,N_5005,N_5143);
and U5217 (N_5217,N_5067,N_5013);
nor U5218 (N_5218,N_5194,N_5039);
and U5219 (N_5219,N_5154,N_5009);
and U5220 (N_5220,N_5065,N_5036);
nor U5221 (N_5221,N_5142,N_5080);
nand U5222 (N_5222,N_5095,N_5081);
xor U5223 (N_5223,N_5179,N_5078);
nor U5224 (N_5224,N_5035,N_5045);
nor U5225 (N_5225,N_5061,N_5177);
or U5226 (N_5226,N_5071,N_5189);
or U5227 (N_5227,N_5197,N_5054);
and U5228 (N_5228,N_5002,N_5087);
or U5229 (N_5229,N_5120,N_5102);
nor U5230 (N_5230,N_5074,N_5122);
nand U5231 (N_5231,N_5130,N_5050);
xor U5232 (N_5232,N_5098,N_5199);
nor U5233 (N_5233,N_5192,N_5195);
nor U5234 (N_5234,N_5163,N_5052);
nor U5235 (N_5235,N_5092,N_5108);
and U5236 (N_5236,N_5094,N_5167);
xor U5237 (N_5237,N_5090,N_5141);
nand U5238 (N_5238,N_5134,N_5187);
xor U5239 (N_5239,N_5051,N_5117);
nand U5240 (N_5240,N_5162,N_5111);
or U5241 (N_5241,N_5008,N_5157);
xnor U5242 (N_5242,N_5076,N_5184);
and U5243 (N_5243,N_5084,N_5186);
nand U5244 (N_5244,N_5059,N_5042);
or U5245 (N_5245,N_5068,N_5083);
xnor U5246 (N_5246,N_5183,N_5031);
and U5247 (N_5247,N_5181,N_5144);
nor U5248 (N_5248,N_5150,N_5064);
and U5249 (N_5249,N_5113,N_5041);
nand U5250 (N_5250,N_5137,N_5000);
xnor U5251 (N_5251,N_5127,N_5003);
nand U5252 (N_5252,N_5044,N_5079);
nor U5253 (N_5253,N_5097,N_5070);
or U5254 (N_5254,N_5160,N_5037);
or U5255 (N_5255,N_5106,N_5015);
and U5256 (N_5256,N_5175,N_5073);
nand U5257 (N_5257,N_5025,N_5026);
or U5258 (N_5258,N_5028,N_5126);
or U5259 (N_5259,N_5193,N_5159);
nor U5260 (N_5260,N_5146,N_5001);
or U5261 (N_5261,N_5114,N_5085);
or U5262 (N_5262,N_5089,N_5138);
nor U5263 (N_5263,N_5125,N_5020);
xnor U5264 (N_5264,N_5118,N_5024);
or U5265 (N_5265,N_5023,N_5033);
or U5266 (N_5266,N_5069,N_5072);
and U5267 (N_5267,N_5018,N_5135);
and U5268 (N_5268,N_5017,N_5007);
and U5269 (N_5269,N_5139,N_5196);
nand U5270 (N_5270,N_5038,N_5133);
nor U5271 (N_5271,N_5166,N_5176);
or U5272 (N_5272,N_5109,N_5149);
nand U5273 (N_5273,N_5191,N_5178);
xor U5274 (N_5274,N_5021,N_5198);
and U5275 (N_5275,N_5103,N_5016);
or U5276 (N_5276,N_5131,N_5190);
nor U5277 (N_5277,N_5129,N_5066);
and U5278 (N_5278,N_5169,N_5096);
xnor U5279 (N_5279,N_5040,N_5173);
nand U5280 (N_5280,N_5128,N_5010);
or U5281 (N_5281,N_5172,N_5148);
or U5282 (N_5282,N_5029,N_5174);
and U5283 (N_5283,N_5145,N_5055);
nand U5284 (N_5284,N_5006,N_5110);
nor U5285 (N_5285,N_5123,N_5032);
nor U5286 (N_5286,N_5151,N_5180);
and U5287 (N_5287,N_5063,N_5153);
or U5288 (N_5288,N_5101,N_5056);
or U5289 (N_5289,N_5121,N_5014);
nand U5290 (N_5290,N_5168,N_5182);
nor U5291 (N_5291,N_5082,N_5004);
nand U5292 (N_5292,N_5093,N_5058);
nand U5293 (N_5293,N_5099,N_5104);
nand U5294 (N_5294,N_5155,N_5152);
and U5295 (N_5295,N_5030,N_5136);
nand U5296 (N_5296,N_5062,N_5027);
and U5297 (N_5297,N_5034,N_5011);
or U5298 (N_5298,N_5115,N_5116);
and U5299 (N_5299,N_5049,N_5132);
nor U5300 (N_5300,N_5193,N_5016);
nand U5301 (N_5301,N_5020,N_5091);
nor U5302 (N_5302,N_5007,N_5018);
nor U5303 (N_5303,N_5182,N_5039);
and U5304 (N_5304,N_5056,N_5075);
nand U5305 (N_5305,N_5062,N_5074);
nor U5306 (N_5306,N_5189,N_5041);
nor U5307 (N_5307,N_5180,N_5160);
and U5308 (N_5308,N_5145,N_5024);
nor U5309 (N_5309,N_5154,N_5018);
nand U5310 (N_5310,N_5027,N_5109);
nor U5311 (N_5311,N_5109,N_5057);
nor U5312 (N_5312,N_5179,N_5014);
nand U5313 (N_5313,N_5062,N_5197);
nand U5314 (N_5314,N_5141,N_5001);
nor U5315 (N_5315,N_5032,N_5152);
or U5316 (N_5316,N_5153,N_5057);
and U5317 (N_5317,N_5107,N_5062);
or U5318 (N_5318,N_5067,N_5189);
nor U5319 (N_5319,N_5084,N_5181);
or U5320 (N_5320,N_5036,N_5074);
and U5321 (N_5321,N_5057,N_5029);
and U5322 (N_5322,N_5000,N_5174);
and U5323 (N_5323,N_5083,N_5127);
nand U5324 (N_5324,N_5005,N_5138);
xnor U5325 (N_5325,N_5179,N_5029);
or U5326 (N_5326,N_5169,N_5018);
nor U5327 (N_5327,N_5024,N_5134);
and U5328 (N_5328,N_5178,N_5139);
or U5329 (N_5329,N_5088,N_5093);
nand U5330 (N_5330,N_5012,N_5187);
nand U5331 (N_5331,N_5098,N_5164);
nand U5332 (N_5332,N_5066,N_5048);
and U5333 (N_5333,N_5190,N_5120);
nand U5334 (N_5334,N_5183,N_5194);
nand U5335 (N_5335,N_5156,N_5036);
nor U5336 (N_5336,N_5091,N_5168);
nand U5337 (N_5337,N_5052,N_5169);
and U5338 (N_5338,N_5101,N_5143);
nor U5339 (N_5339,N_5135,N_5071);
and U5340 (N_5340,N_5013,N_5173);
and U5341 (N_5341,N_5073,N_5184);
nand U5342 (N_5342,N_5084,N_5139);
nand U5343 (N_5343,N_5001,N_5156);
nor U5344 (N_5344,N_5151,N_5149);
or U5345 (N_5345,N_5060,N_5107);
nand U5346 (N_5346,N_5181,N_5029);
or U5347 (N_5347,N_5199,N_5148);
or U5348 (N_5348,N_5039,N_5068);
nand U5349 (N_5349,N_5162,N_5093);
nor U5350 (N_5350,N_5188,N_5054);
nor U5351 (N_5351,N_5073,N_5030);
and U5352 (N_5352,N_5168,N_5134);
and U5353 (N_5353,N_5152,N_5109);
or U5354 (N_5354,N_5107,N_5053);
nand U5355 (N_5355,N_5113,N_5112);
and U5356 (N_5356,N_5173,N_5151);
and U5357 (N_5357,N_5015,N_5110);
and U5358 (N_5358,N_5063,N_5081);
nor U5359 (N_5359,N_5167,N_5021);
or U5360 (N_5360,N_5171,N_5136);
nor U5361 (N_5361,N_5010,N_5109);
nand U5362 (N_5362,N_5134,N_5123);
nor U5363 (N_5363,N_5102,N_5111);
or U5364 (N_5364,N_5105,N_5083);
nor U5365 (N_5365,N_5162,N_5184);
and U5366 (N_5366,N_5197,N_5127);
or U5367 (N_5367,N_5188,N_5127);
nand U5368 (N_5368,N_5051,N_5192);
and U5369 (N_5369,N_5139,N_5142);
nand U5370 (N_5370,N_5175,N_5155);
and U5371 (N_5371,N_5087,N_5100);
or U5372 (N_5372,N_5081,N_5141);
nor U5373 (N_5373,N_5082,N_5010);
and U5374 (N_5374,N_5113,N_5119);
or U5375 (N_5375,N_5059,N_5192);
or U5376 (N_5376,N_5192,N_5108);
nor U5377 (N_5377,N_5073,N_5098);
or U5378 (N_5378,N_5166,N_5182);
and U5379 (N_5379,N_5022,N_5039);
nand U5380 (N_5380,N_5122,N_5105);
nor U5381 (N_5381,N_5126,N_5164);
nor U5382 (N_5382,N_5041,N_5106);
nand U5383 (N_5383,N_5045,N_5034);
or U5384 (N_5384,N_5067,N_5062);
nand U5385 (N_5385,N_5138,N_5053);
or U5386 (N_5386,N_5131,N_5143);
nor U5387 (N_5387,N_5162,N_5045);
or U5388 (N_5388,N_5188,N_5139);
and U5389 (N_5389,N_5179,N_5033);
nand U5390 (N_5390,N_5142,N_5179);
or U5391 (N_5391,N_5033,N_5095);
nor U5392 (N_5392,N_5194,N_5182);
nand U5393 (N_5393,N_5091,N_5186);
and U5394 (N_5394,N_5135,N_5176);
and U5395 (N_5395,N_5138,N_5104);
and U5396 (N_5396,N_5013,N_5144);
or U5397 (N_5397,N_5198,N_5086);
or U5398 (N_5398,N_5083,N_5110);
or U5399 (N_5399,N_5044,N_5013);
nand U5400 (N_5400,N_5390,N_5307);
and U5401 (N_5401,N_5215,N_5279);
xor U5402 (N_5402,N_5320,N_5270);
or U5403 (N_5403,N_5380,N_5218);
nor U5404 (N_5404,N_5353,N_5206);
nand U5405 (N_5405,N_5399,N_5316);
and U5406 (N_5406,N_5385,N_5364);
nand U5407 (N_5407,N_5255,N_5318);
nand U5408 (N_5408,N_5291,N_5295);
and U5409 (N_5409,N_5321,N_5313);
or U5410 (N_5410,N_5303,N_5372);
or U5411 (N_5411,N_5297,N_5214);
or U5412 (N_5412,N_5360,N_5301);
or U5413 (N_5413,N_5217,N_5312);
and U5414 (N_5414,N_5322,N_5266);
or U5415 (N_5415,N_5314,N_5249);
xnor U5416 (N_5416,N_5205,N_5377);
nand U5417 (N_5417,N_5248,N_5337);
nand U5418 (N_5418,N_5379,N_5355);
nand U5419 (N_5419,N_5317,N_5326);
nand U5420 (N_5420,N_5272,N_5392);
nor U5421 (N_5421,N_5290,N_5260);
nand U5422 (N_5422,N_5244,N_5376);
and U5423 (N_5423,N_5370,N_5245);
or U5424 (N_5424,N_5367,N_5247);
or U5425 (N_5425,N_5258,N_5327);
nand U5426 (N_5426,N_5226,N_5207);
or U5427 (N_5427,N_5257,N_5391);
or U5428 (N_5428,N_5275,N_5243);
nand U5429 (N_5429,N_5242,N_5287);
nor U5430 (N_5430,N_5342,N_5292);
nor U5431 (N_5431,N_5282,N_5267);
nand U5432 (N_5432,N_5262,N_5296);
nand U5433 (N_5433,N_5373,N_5365);
nor U5434 (N_5434,N_5371,N_5277);
or U5435 (N_5435,N_5265,N_5237);
nand U5436 (N_5436,N_5200,N_5231);
nor U5437 (N_5437,N_5341,N_5302);
or U5438 (N_5438,N_5223,N_5246);
or U5439 (N_5439,N_5288,N_5294);
and U5440 (N_5440,N_5201,N_5340);
or U5441 (N_5441,N_5230,N_5368);
nor U5442 (N_5442,N_5210,N_5259);
nor U5443 (N_5443,N_5203,N_5256);
nand U5444 (N_5444,N_5343,N_5239);
nor U5445 (N_5445,N_5209,N_5236);
and U5446 (N_5446,N_5232,N_5253);
or U5447 (N_5447,N_5273,N_5235);
nand U5448 (N_5448,N_5208,N_5336);
nand U5449 (N_5449,N_5361,N_5350);
nand U5450 (N_5450,N_5286,N_5252);
or U5451 (N_5451,N_5268,N_5284);
or U5452 (N_5452,N_5397,N_5234);
xor U5453 (N_5453,N_5227,N_5211);
or U5454 (N_5454,N_5333,N_5324);
and U5455 (N_5455,N_5228,N_5363);
xor U5456 (N_5456,N_5304,N_5358);
or U5457 (N_5457,N_5306,N_5384);
and U5458 (N_5458,N_5359,N_5354);
nor U5459 (N_5459,N_5369,N_5383);
nor U5460 (N_5460,N_5389,N_5261);
nor U5461 (N_5461,N_5381,N_5348);
xor U5462 (N_5462,N_5393,N_5281);
and U5463 (N_5463,N_5329,N_5331);
and U5464 (N_5464,N_5366,N_5349);
and U5465 (N_5465,N_5351,N_5222);
or U5466 (N_5466,N_5219,N_5356);
or U5467 (N_5467,N_5319,N_5305);
or U5468 (N_5468,N_5285,N_5308);
xor U5469 (N_5469,N_5240,N_5334);
nand U5470 (N_5470,N_5309,N_5221);
or U5471 (N_5471,N_5298,N_5338);
nor U5472 (N_5472,N_5212,N_5269);
nand U5473 (N_5473,N_5300,N_5204);
nand U5474 (N_5474,N_5345,N_5271);
nor U5475 (N_5475,N_5293,N_5332);
nor U5476 (N_5476,N_5225,N_5299);
xnor U5477 (N_5477,N_5330,N_5283);
or U5478 (N_5478,N_5362,N_5276);
nand U5479 (N_5479,N_5382,N_5386);
and U5480 (N_5480,N_5387,N_5310);
and U5481 (N_5481,N_5263,N_5344);
nor U5482 (N_5482,N_5346,N_5238);
nor U5483 (N_5483,N_5251,N_5394);
or U5484 (N_5484,N_5233,N_5325);
and U5485 (N_5485,N_5202,N_5339);
and U5486 (N_5486,N_5347,N_5315);
nor U5487 (N_5487,N_5278,N_5311);
nand U5488 (N_5488,N_5323,N_5396);
nor U5489 (N_5489,N_5220,N_5398);
nor U5490 (N_5490,N_5328,N_5241);
nand U5491 (N_5491,N_5274,N_5224);
nor U5492 (N_5492,N_5357,N_5213);
nor U5493 (N_5493,N_5229,N_5374);
or U5494 (N_5494,N_5250,N_5216);
or U5495 (N_5495,N_5289,N_5375);
nand U5496 (N_5496,N_5388,N_5395);
nand U5497 (N_5497,N_5378,N_5335);
nor U5498 (N_5498,N_5254,N_5264);
nor U5499 (N_5499,N_5352,N_5280);
or U5500 (N_5500,N_5276,N_5338);
nand U5501 (N_5501,N_5321,N_5243);
nand U5502 (N_5502,N_5231,N_5326);
nand U5503 (N_5503,N_5218,N_5370);
or U5504 (N_5504,N_5348,N_5340);
and U5505 (N_5505,N_5369,N_5321);
or U5506 (N_5506,N_5229,N_5252);
nand U5507 (N_5507,N_5322,N_5393);
or U5508 (N_5508,N_5217,N_5234);
nor U5509 (N_5509,N_5278,N_5246);
or U5510 (N_5510,N_5298,N_5220);
nand U5511 (N_5511,N_5211,N_5383);
nand U5512 (N_5512,N_5347,N_5398);
nand U5513 (N_5513,N_5372,N_5326);
and U5514 (N_5514,N_5382,N_5261);
nand U5515 (N_5515,N_5285,N_5331);
and U5516 (N_5516,N_5252,N_5308);
and U5517 (N_5517,N_5323,N_5214);
xor U5518 (N_5518,N_5306,N_5322);
nand U5519 (N_5519,N_5242,N_5382);
or U5520 (N_5520,N_5396,N_5290);
nand U5521 (N_5521,N_5321,N_5215);
and U5522 (N_5522,N_5238,N_5226);
xor U5523 (N_5523,N_5345,N_5264);
nand U5524 (N_5524,N_5241,N_5318);
nor U5525 (N_5525,N_5386,N_5319);
and U5526 (N_5526,N_5213,N_5353);
nor U5527 (N_5527,N_5379,N_5222);
xor U5528 (N_5528,N_5259,N_5246);
or U5529 (N_5529,N_5240,N_5337);
nand U5530 (N_5530,N_5369,N_5312);
or U5531 (N_5531,N_5232,N_5292);
or U5532 (N_5532,N_5344,N_5208);
or U5533 (N_5533,N_5344,N_5273);
or U5534 (N_5534,N_5338,N_5362);
nand U5535 (N_5535,N_5291,N_5357);
or U5536 (N_5536,N_5250,N_5252);
nor U5537 (N_5537,N_5383,N_5273);
xnor U5538 (N_5538,N_5327,N_5324);
or U5539 (N_5539,N_5257,N_5313);
and U5540 (N_5540,N_5356,N_5209);
nor U5541 (N_5541,N_5281,N_5395);
and U5542 (N_5542,N_5253,N_5369);
nor U5543 (N_5543,N_5386,N_5353);
xnor U5544 (N_5544,N_5278,N_5250);
and U5545 (N_5545,N_5313,N_5293);
or U5546 (N_5546,N_5282,N_5396);
nand U5547 (N_5547,N_5264,N_5220);
nand U5548 (N_5548,N_5273,N_5312);
or U5549 (N_5549,N_5379,N_5322);
or U5550 (N_5550,N_5217,N_5275);
and U5551 (N_5551,N_5378,N_5215);
nor U5552 (N_5552,N_5255,N_5258);
nor U5553 (N_5553,N_5214,N_5258);
nand U5554 (N_5554,N_5370,N_5389);
or U5555 (N_5555,N_5365,N_5230);
nand U5556 (N_5556,N_5321,N_5242);
nor U5557 (N_5557,N_5305,N_5318);
or U5558 (N_5558,N_5329,N_5360);
nor U5559 (N_5559,N_5230,N_5229);
xnor U5560 (N_5560,N_5331,N_5384);
or U5561 (N_5561,N_5276,N_5249);
nor U5562 (N_5562,N_5394,N_5380);
nor U5563 (N_5563,N_5313,N_5258);
and U5564 (N_5564,N_5362,N_5223);
nor U5565 (N_5565,N_5214,N_5203);
nand U5566 (N_5566,N_5236,N_5342);
nand U5567 (N_5567,N_5247,N_5279);
and U5568 (N_5568,N_5246,N_5358);
nand U5569 (N_5569,N_5331,N_5284);
or U5570 (N_5570,N_5375,N_5279);
and U5571 (N_5571,N_5354,N_5271);
nand U5572 (N_5572,N_5379,N_5275);
nand U5573 (N_5573,N_5235,N_5385);
or U5574 (N_5574,N_5271,N_5258);
and U5575 (N_5575,N_5206,N_5331);
and U5576 (N_5576,N_5230,N_5253);
nor U5577 (N_5577,N_5256,N_5213);
and U5578 (N_5578,N_5235,N_5216);
nand U5579 (N_5579,N_5243,N_5382);
or U5580 (N_5580,N_5280,N_5329);
xor U5581 (N_5581,N_5332,N_5229);
nand U5582 (N_5582,N_5203,N_5358);
xnor U5583 (N_5583,N_5397,N_5262);
and U5584 (N_5584,N_5388,N_5346);
or U5585 (N_5585,N_5282,N_5200);
nand U5586 (N_5586,N_5366,N_5326);
or U5587 (N_5587,N_5347,N_5243);
and U5588 (N_5588,N_5346,N_5281);
nand U5589 (N_5589,N_5317,N_5383);
nand U5590 (N_5590,N_5361,N_5329);
nand U5591 (N_5591,N_5309,N_5344);
xnor U5592 (N_5592,N_5221,N_5396);
and U5593 (N_5593,N_5307,N_5356);
or U5594 (N_5594,N_5241,N_5226);
nand U5595 (N_5595,N_5396,N_5359);
nand U5596 (N_5596,N_5366,N_5368);
and U5597 (N_5597,N_5324,N_5202);
or U5598 (N_5598,N_5304,N_5303);
or U5599 (N_5599,N_5250,N_5334);
nand U5600 (N_5600,N_5543,N_5551);
or U5601 (N_5601,N_5411,N_5546);
xnor U5602 (N_5602,N_5522,N_5405);
nor U5603 (N_5603,N_5418,N_5417);
and U5604 (N_5604,N_5459,N_5413);
nand U5605 (N_5605,N_5565,N_5483);
and U5606 (N_5606,N_5503,N_5554);
nand U5607 (N_5607,N_5429,N_5523);
nor U5608 (N_5608,N_5545,N_5457);
nor U5609 (N_5609,N_5514,N_5557);
or U5610 (N_5610,N_5473,N_5492);
nor U5611 (N_5611,N_5590,N_5531);
nand U5612 (N_5612,N_5427,N_5499);
or U5613 (N_5613,N_5437,N_5535);
or U5614 (N_5614,N_5506,N_5401);
or U5615 (N_5615,N_5453,N_5436);
nor U5616 (N_5616,N_5480,N_5454);
nor U5617 (N_5617,N_5526,N_5441);
or U5618 (N_5618,N_5442,N_5493);
nand U5619 (N_5619,N_5567,N_5451);
nand U5620 (N_5620,N_5450,N_5577);
nand U5621 (N_5621,N_5564,N_5532);
nand U5622 (N_5622,N_5484,N_5595);
nor U5623 (N_5623,N_5434,N_5485);
xor U5624 (N_5624,N_5525,N_5561);
xor U5625 (N_5625,N_5544,N_5537);
and U5626 (N_5626,N_5589,N_5460);
xor U5627 (N_5627,N_5425,N_5416);
nand U5628 (N_5628,N_5443,N_5599);
nor U5629 (N_5629,N_5432,N_5540);
and U5630 (N_5630,N_5422,N_5482);
and U5631 (N_5631,N_5448,N_5475);
nor U5632 (N_5632,N_5500,N_5410);
or U5633 (N_5633,N_5515,N_5556);
nor U5634 (N_5634,N_5445,N_5517);
nor U5635 (N_5635,N_5471,N_5518);
or U5636 (N_5636,N_5596,N_5539);
or U5637 (N_5637,N_5468,N_5547);
nor U5638 (N_5638,N_5406,N_5513);
and U5639 (N_5639,N_5456,N_5400);
nand U5640 (N_5640,N_5516,N_5527);
nor U5641 (N_5641,N_5553,N_5494);
or U5642 (N_5642,N_5466,N_5541);
and U5643 (N_5643,N_5594,N_5458);
and U5644 (N_5644,N_5412,N_5433);
nor U5645 (N_5645,N_5404,N_5470);
and U5646 (N_5646,N_5461,N_5569);
or U5647 (N_5647,N_5428,N_5440);
xnor U5648 (N_5648,N_5402,N_5414);
xnor U5649 (N_5649,N_5464,N_5487);
xor U5650 (N_5650,N_5449,N_5498);
nor U5651 (N_5651,N_5528,N_5568);
or U5652 (N_5652,N_5519,N_5566);
xnor U5653 (N_5653,N_5585,N_5420);
nand U5654 (N_5654,N_5421,N_5455);
nor U5655 (N_5655,N_5511,N_5444);
nand U5656 (N_5656,N_5530,N_5572);
and U5657 (N_5657,N_5550,N_5476);
or U5658 (N_5658,N_5534,N_5552);
nor U5659 (N_5659,N_5587,N_5533);
nor U5660 (N_5660,N_5469,N_5593);
nand U5661 (N_5661,N_5521,N_5580);
or U5662 (N_5662,N_5562,N_5463);
or U5663 (N_5663,N_5598,N_5581);
and U5664 (N_5664,N_5520,N_5472);
nor U5665 (N_5665,N_5446,N_5510);
nand U5666 (N_5666,N_5426,N_5555);
or U5667 (N_5667,N_5502,N_5586);
nand U5668 (N_5668,N_5549,N_5559);
nand U5669 (N_5669,N_5579,N_5462);
nand U5670 (N_5670,N_5542,N_5508);
nor U5671 (N_5671,N_5486,N_5576);
or U5672 (N_5672,N_5496,N_5465);
nand U5673 (N_5673,N_5512,N_5538);
nand U5674 (N_5674,N_5439,N_5573);
nand U5675 (N_5675,N_5430,N_5438);
nand U5676 (N_5676,N_5488,N_5431);
nand U5677 (N_5677,N_5447,N_5505);
nor U5678 (N_5678,N_5419,N_5582);
or U5679 (N_5679,N_5479,N_5504);
nand U5680 (N_5680,N_5558,N_5490);
nand U5681 (N_5681,N_5588,N_5524);
and U5682 (N_5682,N_5574,N_5584);
and U5683 (N_5683,N_5583,N_5507);
nor U5684 (N_5684,N_5501,N_5563);
or U5685 (N_5685,N_5403,N_5478);
and U5686 (N_5686,N_5423,N_5415);
or U5687 (N_5687,N_5536,N_5452);
or U5688 (N_5688,N_5560,N_5467);
xor U5689 (N_5689,N_5408,N_5591);
nand U5690 (N_5690,N_5509,N_5575);
and U5691 (N_5691,N_5571,N_5489);
nor U5692 (N_5692,N_5578,N_5477);
or U5693 (N_5693,N_5548,N_5474);
nand U5694 (N_5694,N_5491,N_5435);
and U5695 (N_5695,N_5424,N_5497);
or U5696 (N_5696,N_5409,N_5592);
nand U5697 (N_5697,N_5597,N_5495);
nor U5698 (N_5698,N_5407,N_5481);
and U5699 (N_5699,N_5529,N_5570);
nand U5700 (N_5700,N_5573,N_5489);
or U5701 (N_5701,N_5482,N_5506);
nor U5702 (N_5702,N_5455,N_5405);
or U5703 (N_5703,N_5478,N_5531);
nand U5704 (N_5704,N_5524,N_5523);
nand U5705 (N_5705,N_5550,N_5590);
nor U5706 (N_5706,N_5553,N_5575);
and U5707 (N_5707,N_5527,N_5537);
nor U5708 (N_5708,N_5548,N_5520);
nand U5709 (N_5709,N_5485,N_5409);
nor U5710 (N_5710,N_5476,N_5572);
nor U5711 (N_5711,N_5433,N_5492);
or U5712 (N_5712,N_5520,N_5418);
and U5713 (N_5713,N_5487,N_5465);
nand U5714 (N_5714,N_5483,N_5415);
or U5715 (N_5715,N_5538,N_5570);
or U5716 (N_5716,N_5475,N_5424);
nand U5717 (N_5717,N_5492,N_5567);
xor U5718 (N_5718,N_5576,N_5485);
nor U5719 (N_5719,N_5443,N_5573);
nor U5720 (N_5720,N_5468,N_5594);
and U5721 (N_5721,N_5547,N_5466);
xor U5722 (N_5722,N_5537,N_5429);
and U5723 (N_5723,N_5520,N_5542);
nor U5724 (N_5724,N_5557,N_5551);
or U5725 (N_5725,N_5435,N_5494);
nor U5726 (N_5726,N_5590,N_5417);
xnor U5727 (N_5727,N_5558,N_5454);
nand U5728 (N_5728,N_5561,N_5544);
nand U5729 (N_5729,N_5410,N_5472);
or U5730 (N_5730,N_5541,N_5550);
nand U5731 (N_5731,N_5515,N_5546);
nand U5732 (N_5732,N_5543,N_5531);
nand U5733 (N_5733,N_5403,N_5581);
and U5734 (N_5734,N_5511,N_5490);
xnor U5735 (N_5735,N_5485,N_5441);
and U5736 (N_5736,N_5462,N_5539);
nor U5737 (N_5737,N_5593,N_5420);
nor U5738 (N_5738,N_5405,N_5461);
nor U5739 (N_5739,N_5412,N_5475);
or U5740 (N_5740,N_5590,N_5585);
or U5741 (N_5741,N_5524,N_5579);
nand U5742 (N_5742,N_5519,N_5469);
and U5743 (N_5743,N_5582,N_5576);
nor U5744 (N_5744,N_5503,N_5596);
and U5745 (N_5745,N_5454,N_5536);
nor U5746 (N_5746,N_5558,N_5516);
nand U5747 (N_5747,N_5550,N_5533);
or U5748 (N_5748,N_5551,N_5432);
nand U5749 (N_5749,N_5593,N_5437);
nor U5750 (N_5750,N_5552,N_5425);
nand U5751 (N_5751,N_5441,N_5556);
nor U5752 (N_5752,N_5531,N_5424);
xnor U5753 (N_5753,N_5412,N_5587);
nand U5754 (N_5754,N_5400,N_5592);
and U5755 (N_5755,N_5431,N_5444);
nand U5756 (N_5756,N_5582,N_5571);
nand U5757 (N_5757,N_5423,N_5541);
or U5758 (N_5758,N_5462,N_5505);
xor U5759 (N_5759,N_5427,N_5519);
and U5760 (N_5760,N_5566,N_5531);
nor U5761 (N_5761,N_5430,N_5500);
or U5762 (N_5762,N_5468,N_5578);
nor U5763 (N_5763,N_5577,N_5522);
nor U5764 (N_5764,N_5481,N_5429);
xnor U5765 (N_5765,N_5464,N_5585);
nor U5766 (N_5766,N_5450,N_5555);
nor U5767 (N_5767,N_5526,N_5420);
nor U5768 (N_5768,N_5536,N_5438);
or U5769 (N_5769,N_5593,N_5554);
and U5770 (N_5770,N_5468,N_5588);
nand U5771 (N_5771,N_5493,N_5424);
and U5772 (N_5772,N_5457,N_5459);
nand U5773 (N_5773,N_5567,N_5566);
nand U5774 (N_5774,N_5432,N_5543);
and U5775 (N_5775,N_5405,N_5504);
xnor U5776 (N_5776,N_5529,N_5583);
nand U5777 (N_5777,N_5561,N_5542);
xnor U5778 (N_5778,N_5400,N_5588);
or U5779 (N_5779,N_5525,N_5529);
nand U5780 (N_5780,N_5450,N_5480);
and U5781 (N_5781,N_5480,N_5561);
and U5782 (N_5782,N_5420,N_5543);
nand U5783 (N_5783,N_5469,N_5496);
and U5784 (N_5784,N_5511,N_5585);
and U5785 (N_5785,N_5558,N_5588);
and U5786 (N_5786,N_5588,N_5543);
nand U5787 (N_5787,N_5477,N_5435);
nand U5788 (N_5788,N_5507,N_5560);
or U5789 (N_5789,N_5440,N_5523);
or U5790 (N_5790,N_5418,N_5464);
and U5791 (N_5791,N_5428,N_5576);
nand U5792 (N_5792,N_5455,N_5569);
nor U5793 (N_5793,N_5559,N_5545);
or U5794 (N_5794,N_5463,N_5540);
and U5795 (N_5795,N_5566,N_5443);
nor U5796 (N_5796,N_5479,N_5539);
nand U5797 (N_5797,N_5450,N_5563);
xor U5798 (N_5798,N_5585,N_5463);
nand U5799 (N_5799,N_5408,N_5476);
or U5800 (N_5800,N_5617,N_5795);
or U5801 (N_5801,N_5608,N_5743);
nor U5802 (N_5802,N_5771,N_5615);
nor U5803 (N_5803,N_5616,N_5643);
and U5804 (N_5804,N_5669,N_5630);
xor U5805 (N_5805,N_5611,N_5726);
nand U5806 (N_5806,N_5605,N_5622);
nand U5807 (N_5807,N_5702,N_5654);
nor U5808 (N_5808,N_5704,N_5618);
and U5809 (N_5809,N_5635,N_5679);
and U5810 (N_5810,N_5609,N_5728);
nand U5811 (N_5811,N_5751,N_5778);
nor U5812 (N_5812,N_5690,N_5723);
and U5813 (N_5813,N_5683,N_5668);
and U5814 (N_5814,N_5745,N_5652);
and U5815 (N_5815,N_5787,N_5730);
or U5816 (N_5816,N_5767,N_5686);
or U5817 (N_5817,N_5716,N_5684);
and U5818 (N_5818,N_5748,N_5670);
nor U5819 (N_5819,N_5760,N_5680);
nor U5820 (N_5820,N_5759,N_5665);
xor U5821 (N_5821,N_5762,N_5604);
nor U5822 (N_5822,N_5674,N_5629);
nand U5823 (N_5823,N_5644,N_5747);
nand U5824 (N_5824,N_5734,N_5736);
and U5825 (N_5825,N_5638,N_5648);
or U5826 (N_5826,N_5664,N_5688);
or U5827 (N_5827,N_5793,N_5667);
and U5828 (N_5828,N_5756,N_5636);
nor U5829 (N_5829,N_5695,N_5676);
nor U5830 (N_5830,N_5752,N_5722);
nand U5831 (N_5831,N_5639,N_5719);
nand U5832 (N_5832,N_5602,N_5773);
xnor U5833 (N_5833,N_5632,N_5768);
nor U5834 (N_5834,N_5625,N_5701);
nor U5835 (N_5835,N_5753,N_5682);
nor U5836 (N_5836,N_5749,N_5784);
xnor U5837 (N_5837,N_5781,N_5610);
nand U5838 (N_5838,N_5746,N_5698);
nand U5839 (N_5839,N_5685,N_5754);
nor U5840 (N_5840,N_5614,N_5789);
and U5841 (N_5841,N_5623,N_5717);
or U5842 (N_5842,N_5631,N_5764);
nor U5843 (N_5843,N_5647,N_5708);
and U5844 (N_5844,N_5713,N_5656);
or U5845 (N_5845,N_5799,N_5653);
nor U5846 (N_5846,N_5740,N_5655);
and U5847 (N_5847,N_5696,N_5687);
xor U5848 (N_5848,N_5732,N_5720);
nor U5849 (N_5849,N_5779,N_5729);
and U5850 (N_5850,N_5731,N_5738);
or U5851 (N_5851,N_5606,N_5645);
nand U5852 (N_5852,N_5774,N_5607);
or U5853 (N_5853,N_5763,N_5703);
xnor U5854 (N_5854,N_5785,N_5733);
nor U5855 (N_5855,N_5727,N_5601);
nor U5856 (N_5856,N_5775,N_5673);
nor U5857 (N_5857,N_5699,N_5714);
nor U5858 (N_5858,N_5626,N_5711);
nor U5859 (N_5859,N_5661,N_5624);
nand U5860 (N_5860,N_5666,N_5649);
nand U5861 (N_5861,N_5659,N_5788);
nor U5862 (N_5862,N_5692,N_5650);
xnor U5863 (N_5863,N_5671,N_5757);
nor U5864 (N_5864,N_5697,N_5613);
nor U5865 (N_5865,N_5721,N_5707);
xnor U5866 (N_5866,N_5797,N_5766);
nand U5867 (N_5867,N_5741,N_5627);
nor U5868 (N_5868,N_5678,N_5709);
and U5869 (N_5869,N_5640,N_5663);
nand U5870 (N_5870,N_5735,N_5628);
and U5871 (N_5871,N_5657,N_5621);
or U5872 (N_5872,N_5700,N_5742);
nor U5873 (N_5873,N_5782,N_5710);
and U5874 (N_5874,N_5770,N_5786);
or U5875 (N_5875,N_5637,N_5681);
or U5876 (N_5876,N_5705,N_5744);
or U5877 (N_5877,N_5769,N_5694);
nor U5878 (N_5878,N_5798,N_5725);
nand U5879 (N_5879,N_5758,N_5691);
xnor U5880 (N_5880,N_5612,N_5672);
nor U5881 (N_5881,N_5737,N_5658);
nor U5882 (N_5882,N_5794,N_5796);
or U5883 (N_5883,N_5633,N_5780);
or U5884 (N_5884,N_5750,N_5755);
and U5885 (N_5885,N_5660,N_5724);
nand U5886 (N_5886,N_5791,N_5718);
or U5887 (N_5887,N_5646,N_5772);
nand U5888 (N_5888,N_5600,N_5739);
and U5889 (N_5889,N_5777,N_5689);
nand U5890 (N_5890,N_5603,N_5790);
and U5891 (N_5891,N_5792,N_5620);
xnor U5892 (N_5892,N_5675,N_5642);
or U5893 (N_5893,N_5776,N_5619);
nor U5894 (N_5894,N_5715,N_5634);
nand U5895 (N_5895,N_5651,N_5761);
nand U5896 (N_5896,N_5693,N_5712);
and U5897 (N_5897,N_5641,N_5706);
and U5898 (N_5898,N_5783,N_5677);
nand U5899 (N_5899,N_5765,N_5662);
xor U5900 (N_5900,N_5782,N_5671);
or U5901 (N_5901,N_5638,N_5777);
xor U5902 (N_5902,N_5621,N_5780);
nor U5903 (N_5903,N_5623,N_5720);
nor U5904 (N_5904,N_5675,N_5605);
nor U5905 (N_5905,N_5736,N_5785);
and U5906 (N_5906,N_5738,N_5606);
nand U5907 (N_5907,N_5782,N_5681);
nor U5908 (N_5908,N_5656,N_5614);
nand U5909 (N_5909,N_5692,N_5608);
and U5910 (N_5910,N_5743,N_5742);
and U5911 (N_5911,N_5704,N_5727);
nand U5912 (N_5912,N_5773,N_5646);
nand U5913 (N_5913,N_5775,N_5693);
nor U5914 (N_5914,N_5787,N_5607);
nand U5915 (N_5915,N_5798,N_5709);
or U5916 (N_5916,N_5672,N_5789);
nor U5917 (N_5917,N_5693,N_5617);
and U5918 (N_5918,N_5706,N_5623);
or U5919 (N_5919,N_5609,N_5696);
nor U5920 (N_5920,N_5678,N_5602);
nor U5921 (N_5921,N_5662,N_5723);
nand U5922 (N_5922,N_5762,N_5770);
nor U5923 (N_5923,N_5738,N_5788);
nor U5924 (N_5924,N_5674,N_5791);
and U5925 (N_5925,N_5769,N_5670);
nor U5926 (N_5926,N_5716,N_5607);
nand U5927 (N_5927,N_5784,N_5729);
or U5928 (N_5928,N_5746,N_5740);
and U5929 (N_5929,N_5638,N_5747);
and U5930 (N_5930,N_5704,N_5708);
nand U5931 (N_5931,N_5702,N_5643);
and U5932 (N_5932,N_5799,N_5663);
or U5933 (N_5933,N_5753,N_5770);
or U5934 (N_5934,N_5675,N_5648);
nor U5935 (N_5935,N_5603,N_5718);
nand U5936 (N_5936,N_5656,N_5703);
or U5937 (N_5937,N_5613,N_5781);
nand U5938 (N_5938,N_5672,N_5601);
nand U5939 (N_5939,N_5690,N_5643);
nor U5940 (N_5940,N_5798,N_5771);
or U5941 (N_5941,N_5772,N_5634);
nor U5942 (N_5942,N_5782,N_5715);
and U5943 (N_5943,N_5698,N_5710);
and U5944 (N_5944,N_5728,N_5793);
nor U5945 (N_5945,N_5679,N_5761);
nand U5946 (N_5946,N_5796,N_5681);
and U5947 (N_5947,N_5727,N_5723);
or U5948 (N_5948,N_5664,N_5731);
or U5949 (N_5949,N_5626,N_5755);
and U5950 (N_5950,N_5704,N_5639);
or U5951 (N_5951,N_5669,N_5785);
nor U5952 (N_5952,N_5644,N_5653);
nor U5953 (N_5953,N_5699,N_5677);
or U5954 (N_5954,N_5698,N_5773);
xor U5955 (N_5955,N_5657,N_5662);
and U5956 (N_5956,N_5794,N_5775);
or U5957 (N_5957,N_5643,N_5689);
nand U5958 (N_5958,N_5766,N_5799);
nor U5959 (N_5959,N_5680,N_5728);
nor U5960 (N_5960,N_5783,N_5776);
or U5961 (N_5961,N_5662,N_5798);
and U5962 (N_5962,N_5790,N_5703);
xnor U5963 (N_5963,N_5759,N_5701);
and U5964 (N_5964,N_5636,N_5648);
and U5965 (N_5965,N_5654,N_5738);
nand U5966 (N_5966,N_5744,N_5762);
xor U5967 (N_5967,N_5701,N_5622);
and U5968 (N_5968,N_5731,N_5709);
nor U5969 (N_5969,N_5699,N_5710);
xnor U5970 (N_5970,N_5675,N_5609);
nor U5971 (N_5971,N_5782,N_5758);
or U5972 (N_5972,N_5602,N_5667);
or U5973 (N_5973,N_5797,N_5717);
nand U5974 (N_5974,N_5755,N_5661);
or U5975 (N_5975,N_5682,N_5787);
and U5976 (N_5976,N_5715,N_5659);
or U5977 (N_5977,N_5614,N_5778);
or U5978 (N_5978,N_5783,N_5638);
nor U5979 (N_5979,N_5660,N_5672);
or U5980 (N_5980,N_5726,N_5723);
and U5981 (N_5981,N_5638,N_5770);
and U5982 (N_5982,N_5642,N_5622);
nand U5983 (N_5983,N_5694,N_5756);
nor U5984 (N_5984,N_5629,N_5687);
and U5985 (N_5985,N_5775,N_5777);
nor U5986 (N_5986,N_5615,N_5783);
and U5987 (N_5987,N_5748,N_5686);
and U5988 (N_5988,N_5767,N_5749);
or U5989 (N_5989,N_5746,N_5749);
nor U5990 (N_5990,N_5785,N_5727);
and U5991 (N_5991,N_5718,N_5633);
nand U5992 (N_5992,N_5792,N_5712);
nand U5993 (N_5993,N_5627,N_5702);
or U5994 (N_5994,N_5786,N_5692);
or U5995 (N_5995,N_5666,N_5690);
or U5996 (N_5996,N_5644,N_5779);
and U5997 (N_5997,N_5607,N_5722);
and U5998 (N_5998,N_5779,N_5673);
nor U5999 (N_5999,N_5746,N_5683);
or U6000 (N_6000,N_5970,N_5988);
nor U6001 (N_6001,N_5800,N_5856);
xor U6002 (N_6002,N_5893,N_5839);
and U6003 (N_6003,N_5904,N_5853);
nor U6004 (N_6004,N_5876,N_5941);
nor U6005 (N_6005,N_5946,N_5892);
nor U6006 (N_6006,N_5801,N_5850);
and U6007 (N_6007,N_5938,N_5875);
xnor U6008 (N_6008,N_5939,N_5991);
nand U6009 (N_6009,N_5819,N_5914);
and U6010 (N_6010,N_5895,N_5882);
and U6011 (N_6011,N_5982,N_5865);
nand U6012 (N_6012,N_5950,N_5960);
and U6013 (N_6013,N_5944,N_5905);
nand U6014 (N_6014,N_5985,N_5930);
and U6015 (N_6015,N_5820,N_5841);
nand U6016 (N_6016,N_5927,N_5986);
or U6017 (N_6017,N_5869,N_5842);
nand U6018 (N_6018,N_5890,N_5874);
xor U6019 (N_6019,N_5908,N_5872);
nand U6020 (N_6020,N_5824,N_5866);
nand U6021 (N_6021,N_5952,N_5848);
or U6022 (N_6022,N_5851,N_5928);
and U6023 (N_6023,N_5843,N_5812);
nor U6024 (N_6024,N_5947,N_5911);
or U6025 (N_6025,N_5807,N_5955);
or U6026 (N_6026,N_5997,N_5864);
and U6027 (N_6027,N_5883,N_5836);
or U6028 (N_6028,N_5860,N_5958);
nand U6029 (N_6029,N_5959,N_5937);
and U6030 (N_6030,N_5825,N_5983);
xor U6031 (N_6031,N_5867,N_5802);
and U6032 (N_6032,N_5898,N_5921);
nor U6033 (N_6033,N_5925,N_5870);
xor U6034 (N_6034,N_5894,N_5844);
xor U6035 (N_6035,N_5940,N_5976);
or U6036 (N_6036,N_5971,N_5981);
and U6037 (N_6037,N_5957,N_5840);
or U6038 (N_6038,N_5979,N_5859);
xor U6039 (N_6039,N_5936,N_5810);
and U6040 (N_6040,N_5920,N_5877);
nand U6041 (N_6041,N_5934,N_5815);
nand U6042 (N_6042,N_5931,N_5821);
nor U6043 (N_6043,N_5961,N_5951);
nor U6044 (N_6044,N_5832,N_5873);
and U6045 (N_6045,N_5868,N_5980);
nor U6046 (N_6046,N_5863,N_5910);
nand U6047 (N_6047,N_5846,N_5969);
nor U6048 (N_6048,N_5932,N_5949);
nor U6049 (N_6049,N_5984,N_5915);
and U6050 (N_6050,N_5833,N_5923);
or U6051 (N_6051,N_5954,N_5818);
or U6052 (N_6052,N_5896,N_5964);
and U6053 (N_6053,N_5912,N_5900);
xnor U6054 (N_6054,N_5855,N_5805);
and U6055 (N_6055,N_5916,N_5885);
and U6056 (N_6056,N_5968,N_5978);
nand U6057 (N_6057,N_5956,N_5871);
or U6058 (N_6058,N_5834,N_5933);
nand U6059 (N_6059,N_5830,N_5826);
nand U6060 (N_6060,N_5816,N_5858);
and U6061 (N_6061,N_5889,N_5822);
and U6062 (N_6062,N_5935,N_5881);
or U6063 (N_6063,N_5823,N_5854);
xor U6064 (N_6064,N_5977,N_5919);
nor U6065 (N_6065,N_5994,N_5922);
or U6066 (N_6066,N_5887,N_5967);
or U6067 (N_6067,N_5913,N_5897);
or U6068 (N_6068,N_5879,N_5861);
and U6069 (N_6069,N_5829,N_5993);
or U6070 (N_6070,N_5992,N_5998);
nor U6071 (N_6071,N_5972,N_5929);
nand U6072 (N_6072,N_5886,N_5862);
xor U6073 (N_6073,N_5909,N_5803);
nor U6074 (N_6074,N_5999,N_5995);
or U6075 (N_6075,N_5888,N_5852);
nand U6076 (N_6076,N_5847,N_5903);
nor U6077 (N_6077,N_5814,N_5845);
and U6078 (N_6078,N_5948,N_5884);
nand U6079 (N_6079,N_5990,N_5907);
or U6080 (N_6080,N_5831,N_5987);
nand U6081 (N_6081,N_5817,N_5974);
or U6082 (N_6082,N_5891,N_5880);
nor U6083 (N_6083,N_5827,N_5943);
nand U6084 (N_6084,N_5918,N_5963);
or U6085 (N_6085,N_5901,N_5813);
or U6086 (N_6086,N_5945,N_5924);
and U6087 (N_6087,N_5806,N_5962);
xor U6088 (N_6088,N_5808,N_5849);
or U6089 (N_6089,N_5942,N_5809);
and U6090 (N_6090,N_5857,N_5804);
or U6091 (N_6091,N_5973,N_5996);
and U6092 (N_6092,N_5902,N_5917);
nand U6093 (N_6093,N_5838,N_5811);
or U6094 (N_6094,N_5828,N_5966);
nand U6095 (N_6095,N_5953,N_5835);
or U6096 (N_6096,N_5906,N_5975);
nor U6097 (N_6097,N_5837,N_5926);
or U6098 (N_6098,N_5878,N_5965);
nor U6099 (N_6099,N_5899,N_5989);
and U6100 (N_6100,N_5997,N_5937);
nor U6101 (N_6101,N_5940,N_5964);
and U6102 (N_6102,N_5998,N_5918);
and U6103 (N_6103,N_5866,N_5928);
nor U6104 (N_6104,N_5843,N_5807);
nor U6105 (N_6105,N_5888,N_5996);
nand U6106 (N_6106,N_5891,N_5974);
nand U6107 (N_6107,N_5881,N_5993);
nand U6108 (N_6108,N_5933,N_5918);
and U6109 (N_6109,N_5943,N_5882);
and U6110 (N_6110,N_5962,N_5979);
nand U6111 (N_6111,N_5857,N_5970);
or U6112 (N_6112,N_5896,N_5850);
xnor U6113 (N_6113,N_5861,N_5823);
nor U6114 (N_6114,N_5967,N_5843);
nand U6115 (N_6115,N_5834,N_5864);
xnor U6116 (N_6116,N_5938,N_5803);
or U6117 (N_6117,N_5901,N_5920);
and U6118 (N_6118,N_5838,N_5898);
nor U6119 (N_6119,N_5882,N_5951);
nand U6120 (N_6120,N_5923,N_5857);
or U6121 (N_6121,N_5997,N_5874);
nor U6122 (N_6122,N_5977,N_5980);
or U6123 (N_6123,N_5932,N_5927);
nand U6124 (N_6124,N_5970,N_5803);
nand U6125 (N_6125,N_5927,N_5979);
and U6126 (N_6126,N_5875,N_5909);
or U6127 (N_6127,N_5834,N_5858);
xor U6128 (N_6128,N_5890,N_5837);
nand U6129 (N_6129,N_5914,N_5844);
nand U6130 (N_6130,N_5912,N_5890);
nand U6131 (N_6131,N_5914,N_5852);
or U6132 (N_6132,N_5888,N_5802);
nor U6133 (N_6133,N_5861,N_5860);
nand U6134 (N_6134,N_5948,N_5949);
and U6135 (N_6135,N_5916,N_5970);
nand U6136 (N_6136,N_5988,N_5955);
nand U6137 (N_6137,N_5861,N_5920);
xor U6138 (N_6138,N_5877,N_5816);
xor U6139 (N_6139,N_5892,N_5988);
nor U6140 (N_6140,N_5955,N_5869);
nor U6141 (N_6141,N_5830,N_5825);
and U6142 (N_6142,N_5912,N_5837);
nor U6143 (N_6143,N_5941,N_5818);
and U6144 (N_6144,N_5967,N_5908);
nor U6145 (N_6145,N_5953,N_5940);
nor U6146 (N_6146,N_5874,N_5941);
nand U6147 (N_6147,N_5869,N_5846);
nor U6148 (N_6148,N_5966,N_5904);
or U6149 (N_6149,N_5908,N_5873);
or U6150 (N_6150,N_5883,N_5887);
or U6151 (N_6151,N_5895,N_5989);
or U6152 (N_6152,N_5995,N_5903);
or U6153 (N_6153,N_5970,N_5887);
nor U6154 (N_6154,N_5957,N_5894);
xnor U6155 (N_6155,N_5892,N_5856);
or U6156 (N_6156,N_5996,N_5852);
and U6157 (N_6157,N_5932,N_5969);
nand U6158 (N_6158,N_5840,N_5891);
and U6159 (N_6159,N_5806,N_5854);
nor U6160 (N_6160,N_5985,N_5904);
xor U6161 (N_6161,N_5900,N_5922);
or U6162 (N_6162,N_5894,N_5816);
nor U6163 (N_6163,N_5870,N_5907);
and U6164 (N_6164,N_5963,N_5862);
nor U6165 (N_6165,N_5982,N_5967);
xor U6166 (N_6166,N_5898,N_5956);
nor U6167 (N_6167,N_5992,N_5979);
or U6168 (N_6168,N_5978,N_5818);
or U6169 (N_6169,N_5915,N_5844);
or U6170 (N_6170,N_5866,N_5963);
or U6171 (N_6171,N_5943,N_5865);
or U6172 (N_6172,N_5928,N_5887);
or U6173 (N_6173,N_5840,N_5930);
and U6174 (N_6174,N_5948,N_5985);
nor U6175 (N_6175,N_5934,N_5919);
nand U6176 (N_6176,N_5977,N_5848);
or U6177 (N_6177,N_5950,N_5902);
nor U6178 (N_6178,N_5849,N_5894);
and U6179 (N_6179,N_5814,N_5960);
nor U6180 (N_6180,N_5820,N_5952);
nand U6181 (N_6181,N_5961,N_5982);
nor U6182 (N_6182,N_5950,N_5835);
xnor U6183 (N_6183,N_5828,N_5829);
or U6184 (N_6184,N_5976,N_5957);
or U6185 (N_6185,N_5880,N_5956);
nor U6186 (N_6186,N_5948,N_5858);
and U6187 (N_6187,N_5888,N_5831);
xor U6188 (N_6188,N_5924,N_5836);
or U6189 (N_6189,N_5867,N_5907);
nor U6190 (N_6190,N_5828,N_5999);
and U6191 (N_6191,N_5859,N_5997);
or U6192 (N_6192,N_5816,N_5935);
and U6193 (N_6193,N_5971,N_5952);
nor U6194 (N_6194,N_5991,N_5938);
nand U6195 (N_6195,N_5904,N_5928);
nand U6196 (N_6196,N_5966,N_5821);
nand U6197 (N_6197,N_5804,N_5800);
nor U6198 (N_6198,N_5957,N_5962);
or U6199 (N_6199,N_5965,N_5916);
nand U6200 (N_6200,N_6143,N_6044);
or U6201 (N_6201,N_6130,N_6029);
nand U6202 (N_6202,N_6092,N_6064);
nor U6203 (N_6203,N_6008,N_6131);
or U6204 (N_6204,N_6129,N_6073);
nand U6205 (N_6205,N_6163,N_6014);
or U6206 (N_6206,N_6063,N_6159);
nand U6207 (N_6207,N_6108,N_6102);
and U6208 (N_6208,N_6082,N_6089);
or U6209 (N_6209,N_6038,N_6118);
and U6210 (N_6210,N_6070,N_6048);
or U6211 (N_6211,N_6036,N_6154);
and U6212 (N_6212,N_6157,N_6181);
or U6213 (N_6213,N_6085,N_6121);
nor U6214 (N_6214,N_6147,N_6018);
or U6215 (N_6215,N_6066,N_6027);
or U6216 (N_6216,N_6031,N_6145);
nor U6217 (N_6217,N_6171,N_6197);
and U6218 (N_6218,N_6065,N_6193);
or U6219 (N_6219,N_6061,N_6053);
or U6220 (N_6220,N_6125,N_6043);
or U6221 (N_6221,N_6128,N_6059);
or U6222 (N_6222,N_6175,N_6034);
and U6223 (N_6223,N_6123,N_6094);
or U6224 (N_6224,N_6106,N_6137);
nor U6225 (N_6225,N_6049,N_6192);
and U6226 (N_6226,N_6114,N_6052);
nand U6227 (N_6227,N_6168,N_6153);
nand U6228 (N_6228,N_6001,N_6032);
nor U6229 (N_6229,N_6013,N_6051);
and U6230 (N_6230,N_6188,N_6156);
or U6231 (N_6231,N_6030,N_6062);
or U6232 (N_6232,N_6133,N_6182);
xnor U6233 (N_6233,N_6150,N_6100);
and U6234 (N_6234,N_6004,N_6149);
xnor U6235 (N_6235,N_6041,N_6095);
or U6236 (N_6236,N_6119,N_6050);
nor U6237 (N_6237,N_6115,N_6009);
nand U6238 (N_6238,N_6086,N_6170);
nor U6239 (N_6239,N_6028,N_6151);
nor U6240 (N_6240,N_6164,N_6037);
nand U6241 (N_6241,N_6067,N_6080);
or U6242 (N_6242,N_6198,N_6057);
and U6243 (N_6243,N_6103,N_6173);
nor U6244 (N_6244,N_6176,N_6007);
and U6245 (N_6245,N_6180,N_6040);
or U6246 (N_6246,N_6167,N_6039);
nand U6247 (N_6247,N_6113,N_6177);
and U6248 (N_6248,N_6005,N_6186);
xnor U6249 (N_6249,N_6071,N_6010);
nor U6250 (N_6250,N_6148,N_6132);
nand U6251 (N_6251,N_6104,N_6111);
nor U6252 (N_6252,N_6074,N_6017);
nor U6253 (N_6253,N_6047,N_6011);
and U6254 (N_6254,N_6090,N_6088);
and U6255 (N_6255,N_6023,N_6161);
and U6256 (N_6256,N_6190,N_6194);
nor U6257 (N_6257,N_6058,N_6019);
nor U6258 (N_6258,N_6120,N_6166);
and U6259 (N_6259,N_6022,N_6000);
nand U6260 (N_6260,N_6136,N_6075);
xor U6261 (N_6261,N_6116,N_6155);
xor U6262 (N_6262,N_6183,N_6117);
and U6263 (N_6263,N_6184,N_6024);
or U6264 (N_6264,N_6134,N_6172);
xor U6265 (N_6265,N_6109,N_6165);
and U6266 (N_6266,N_6126,N_6093);
or U6267 (N_6267,N_6187,N_6160);
nor U6268 (N_6268,N_6191,N_6179);
and U6269 (N_6269,N_6079,N_6185);
nor U6270 (N_6270,N_6122,N_6015);
xnor U6271 (N_6271,N_6189,N_6098);
and U6272 (N_6272,N_6196,N_6020);
nor U6273 (N_6273,N_6142,N_6084);
xnor U6274 (N_6274,N_6097,N_6158);
nand U6275 (N_6275,N_6139,N_6169);
xnor U6276 (N_6276,N_6112,N_6146);
nor U6277 (N_6277,N_6006,N_6042);
nor U6278 (N_6278,N_6127,N_6096);
nand U6279 (N_6279,N_6199,N_6077);
or U6280 (N_6280,N_6140,N_6138);
nand U6281 (N_6281,N_6003,N_6099);
or U6282 (N_6282,N_6012,N_6162);
xnor U6283 (N_6283,N_6069,N_6055);
and U6284 (N_6284,N_6078,N_6035);
and U6285 (N_6285,N_6101,N_6025);
or U6286 (N_6286,N_6081,N_6124);
and U6287 (N_6287,N_6174,N_6033);
nand U6288 (N_6288,N_6144,N_6054);
or U6289 (N_6289,N_6135,N_6152);
xor U6290 (N_6290,N_6068,N_6107);
xor U6291 (N_6291,N_6178,N_6016);
nor U6292 (N_6292,N_6087,N_6076);
or U6293 (N_6293,N_6002,N_6072);
xnor U6294 (N_6294,N_6046,N_6105);
or U6295 (N_6295,N_6110,N_6141);
and U6296 (N_6296,N_6026,N_6083);
xor U6297 (N_6297,N_6060,N_6021);
nor U6298 (N_6298,N_6091,N_6195);
xnor U6299 (N_6299,N_6056,N_6045);
nor U6300 (N_6300,N_6028,N_6044);
nor U6301 (N_6301,N_6145,N_6157);
or U6302 (N_6302,N_6163,N_6162);
nor U6303 (N_6303,N_6005,N_6166);
and U6304 (N_6304,N_6030,N_6129);
or U6305 (N_6305,N_6154,N_6132);
xnor U6306 (N_6306,N_6132,N_6076);
xnor U6307 (N_6307,N_6135,N_6082);
nor U6308 (N_6308,N_6003,N_6080);
nand U6309 (N_6309,N_6030,N_6098);
nand U6310 (N_6310,N_6164,N_6010);
nor U6311 (N_6311,N_6111,N_6168);
nand U6312 (N_6312,N_6109,N_6000);
nor U6313 (N_6313,N_6033,N_6106);
nor U6314 (N_6314,N_6021,N_6112);
nand U6315 (N_6315,N_6030,N_6168);
or U6316 (N_6316,N_6007,N_6017);
nand U6317 (N_6317,N_6102,N_6060);
and U6318 (N_6318,N_6108,N_6140);
or U6319 (N_6319,N_6110,N_6002);
nor U6320 (N_6320,N_6005,N_6006);
nand U6321 (N_6321,N_6128,N_6146);
or U6322 (N_6322,N_6048,N_6020);
and U6323 (N_6323,N_6091,N_6122);
or U6324 (N_6324,N_6193,N_6126);
or U6325 (N_6325,N_6163,N_6090);
nor U6326 (N_6326,N_6047,N_6052);
nand U6327 (N_6327,N_6169,N_6177);
nor U6328 (N_6328,N_6196,N_6070);
nand U6329 (N_6329,N_6037,N_6034);
or U6330 (N_6330,N_6029,N_6132);
or U6331 (N_6331,N_6012,N_6118);
nor U6332 (N_6332,N_6154,N_6130);
xnor U6333 (N_6333,N_6040,N_6195);
xor U6334 (N_6334,N_6140,N_6179);
nor U6335 (N_6335,N_6116,N_6191);
nor U6336 (N_6336,N_6011,N_6149);
xor U6337 (N_6337,N_6021,N_6121);
or U6338 (N_6338,N_6132,N_6047);
and U6339 (N_6339,N_6126,N_6051);
nor U6340 (N_6340,N_6196,N_6147);
nor U6341 (N_6341,N_6029,N_6060);
or U6342 (N_6342,N_6034,N_6075);
nor U6343 (N_6343,N_6112,N_6099);
nor U6344 (N_6344,N_6025,N_6190);
and U6345 (N_6345,N_6123,N_6117);
xnor U6346 (N_6346,N_6065,N_6187);
nand U6347 (N_6347,N_6194,N_6189);
and U6348 (N_6348,N_6003,N_6067);
or U6349 (N_6349,N_6159,N_6071);
nor U6350 (N_6350,N_6126,N_6022);
nor U6351 (N_6351,N_6068,N_6112);
nand U6352 (N_6352,N_6086,N_6115);
nor U6353 (N_6353,N_6069,N_6106);
xnor U6354 (N_6354,N_6051,N_6090);
nand U6355 (N_6355,N_6097,N_6095);
and U6356 (N_6356,N_6014,N_6179);
nor U6357 (N_6357,N_6145,N_6125);
xnor U6358 (N_6358,N_6038,N_6140);
or U6359 (N_6359,N_6143,N_6112);
nor U6360 (N_6360,N_6021,N_6105);
xnor U6361 (N_6361,N_6163,N_6113);
nand U6362 (N_6362,N_6174,N_6021);
or U6363 (N_6363,N_6018,N_6007);
and U6364 (N_6364,N_6100,N_6142);
or U6365 (N_6365,N_6199,N_6109);
and U6366 (N_6366,N_6120,N_6029);
nor U6367 (N_6367,N_6116,N_6088);
and U6368 (N_6368,N_6116,N_6115);
nand U6369 (N_6369,N_6097,N_6083);
or U6370 (N_6370,N_6147,N_6047);
or U6371 (N_6371,N_6170,N_6151);
xor U6372 (N_6372,N_6192,N_6189);
and U6373 (N_6373,N_6161,N_6149);
and U6374 (N_6374,N_6143,N_6033);
and U6375 (N_6375,N_6108,N_6026);
nor U6376 (N_6376,N_6136,N_6191);
nand U6377 (N_6377,N_6038,N_6078);
nor U6378 (N_6378,N_6123,N_6183);
or U6379 (N_6379,N_6024,N_6149);
nor U6380 (N_6380,N_6025,N_6198);
xnor U6381 (N_6381,N_6153,N_6107);
nand U6382 (N_6382,N_6155,N_6124);
or U6383 (N_6383,N_6049,N_6171);
or U6384 (N_6384,N_6056,N_6078);
or U6385 (N_6385,N_6108,N_6173);
or U6386 (N_6386,N_6164,N_6006);
nor U6387 (N_6387,N_6019,N_6016);
and U6388 (N_6388,N_6179,N_6190);
nand U6389 (N_6389,N_6040,N_6112);
or U6390 (N_6390,N_6005,N_6071);
nand U6391 (N_6391,N_6163,N_6053);
xnor U6392 (N_6392,N_6094,N_6185);
or U6393 (N_6393,N_6171,N_6045);
or U6394 (N_6394,N_6145,N_6013);
or U6395 (N_6395,N_6097,N_6115);
nand U6396 (N_6396,N_6096,N_6028);
or U6397 (N_6397,N_6098,N_6027);
or U6398 (N_6398,N_6004,N_6150);
and U6399 (N_6399,N_6178,N_6005);
nor U6400 (N_6400,N_6396,N_6369);
or U6401 (N_6401,N_6203,N_6275);
nor U6402 (N_6402,N_6364,N_6386);
xor U6403 (N_6403,N_6293,N_6272);
or U6404 (N_6404,N_6294,N_6223);
nor U6405 (N_6405,N_6377,N_6276);
and U6406 (N_6406,N_6297,N_6385);
nor U6407 (N_6407,N_6217,N_6389);
nor U6408 (N_6408,N_6344,N_6277);
nor U6409 (N_6409,N_6285,N_6397);
nand U6410 (N_6410,N_6374,N_6288);
nor U6411 (N_6411,N_6330,N_6218);
xor U6412 (N_6412,N_6229,N_6201);
nand U6413 (N_6413,N_6289,N_6352);
nand U6414 (N_6414,N_6300,N_6209);
or U6415 (N_6415,N_6345,N_6232);
xor U6416 (N_6416,N_6304,N_6360);
xnor U6417 (N_6417,N_6350,N_6376);
or U6418 (N_6418,N_6329,N_6343);
nor U6419 (N_6419,N_6205,N_6328);
or U6420 (N_6420,N_6383,N_6380);
nand U6421 (N_6421,N_6214,N_6313);
nand U6422 (N_6422,N_6332,N_6358);
or U6423 (N_6423,N_6333,N_6357);
nand U6424 (N_6424,N_6335,N_6245);
or U6425 (N_6425,N_6391,N_6341);
nor U6426 (N_6426,N_6219,N_6227);
nand U6427 (N_6427,N_6267,N_6225);
or U6428 (N_6428,N_6254,N_6353);
nor U6429 (N_6429,N_6286,N_6368);
nand U6430 (N_6430,N_6247,N_6371);
and U6431 (N_6431,N_6256,N_6257);
nor U6432 (N_6432,N_6381,N_6216);
nor U6433 (N_6433,N_6261,N_6338);
or U6434 (N_6434,N_6390,N_6239);
nor U6435 (N_6435,N_6316,N_6298);
nor U6436 (N_6436,N_6367,N_6248);
nor U6437 (N_6437,N_6321,N_6244);
and U6438 (N_6438,N_6237,N_6236);
nand U6439 (N_6439,N_6359,N_6246);
and U6440 (N_6440,N_6273,N_6312);
and U6441 (N_6441,N_6331,N_6399);
nor U6442 (N_6442,N_6342,N_6283);
xor U6443 (N_6443,N_6266,N_6280);
nor U6444 (N_6444,N_6392,N_6238);
nor U6445 (N_6445,N_6215,N_6263);
nor U6446 (N_6446,N_6210,N_6361);
or U6447 (N_6447,N_6222,N_6281);
or U6448 (N_6448,N_6325,N_6271);
or U6449 (N_6449,N_6398,N_6296);
nor U6450 (N_6450,N_6303,N_6307);
nor U6451 (N_6451,N_6395,N_6234);
nand U6452 (N_6452,N_6258,N_6240);
xor U6453 (N_6453,N_6260,N_6362);
xor U6454 (N_6454,N_6235,N_6327);
nor U6455 (N_6455,N_6299,N_6379);
nor U6456 (N_6456,N_6268,N_6306);
nand U6457 (N_6457,N_6259,N_6202);
xnor U6458 (N_6458,N_6317,N_6382);
and U6459 (N_6459,N_6243,N_6274);
nand U6460 (N_6460,N_6365,N_6284);
nor U6461 (N_6461,N_6340,N_6233);
and U6462 (N_6462,N_6208,N_6388);
nand U6463 (N_6463,N_6373,N_6270);
nand U6464 (N_6464,N_6290,N_6220);
or U6465 (N_6465,N_6242,N_6302);
nor U6466 (N_6466,N_6206,N_6320);
or U6467 (N_6467,N_6308,N_6253);
nor U6468 (N_6468,N_6322,N_6230);
nand U6469 (N_6469,N_6212,N_6250);
and U6470 (N_6470,N_6213,N_6228);
and U6471 (N_6471,N_6323,N_6346);
or U6472 (N_6472,N_6318,N_6375);
and U6473 (N_6473,N_6372,N_6249);
or U6474 (N_6474,N_6292,N_6334);
or U6475 (N_6475,N_6337,N_6310);
or U6476 (N_6476,N_6349,N_6269);
and U6477 (N_6477,N_6394,N_6311);
xnor U6478 (N_6478,N_6351,N_6291);
and U6479 (N_6479,N_6252,N_6378);
nand U6480 (N_6480,N_6265,N_6314);
nand U6481 (N_6481,N_6315,N_6295);
nor U6482 (N_6482,N_6282,N_6356);
and U6483 (N_6483,N_6301,N_6326);
or U6484 (N_6484,N_6255,N_6309);
nor U6485 (N_6485,N_6324,N_6348);
and U6486 (N_6486,N_6224,N_6278);
and U6487 (N_6487,N_6231,N_6264);
and U6488 (N_6488,N_6370,N_6393);
nor U6489 (N_6489,N_6354,N_6387);
nor U6490 (N_6490,N_6262,N_6305);
and U6491 (N_6491,N_6200,N_6384);
and U6492 (N_6492,N_6251,N_6363);
and U6493 (N_6493,N_6204,N_6226);
xor U6494 (N_6494,N_6221,N_6355);
nand U6495 (N_6495,N_6366,N_6336);
nor U6496 (N_6496,N_6287,N_6279);
nand U6497 (N_6497,N_6241,N_6347);
nand U6498 (N_6498,N_6207,N_6211);
nand U6499 (N_6499,N_6339,N_6319);
nand U6500 (N_6500,N_6388,N_6348);
or U6501 (N_6501,N_6237,N_6393);
and U6502 (N_6502,N_6325,N_6253);
and U6503 (N_6503,N_6318,N_6211);
or U6504 (N_6504,N_6324,N_6354);
or U6505 (N_6505,N_6301,N_6371);
and U6506 (N_6506,N_6363,N_6348);
nand U6507 (N_6507,N_6310,N_6324);
or U6508 (N_6508,N_6256,N_6398);
xor U6509 (N_6509,N_6258,N_6244);
nor U6510 (N_6510,N_6224,N_6341);
xnor U6511 (N_6511,N_6356,N_6258);
or U6512 (N_6512,N_6316,N_6349);
or U6513 (N_6513,N_6323,N_6328);
xor U6514 (N_6514,N_6310,N_6372);
nand U6515 (N_6515,N_6248,N_6241);
nor U6516 (N_6516,N_6253,N_6317);
nand U6517 (N_6517,N_6388,N_6399);
xnor U6518 (N_6518,N_6254,N_6285);
nor U6519 (N_6519,N_6208,N_6306);
nor U6520 (N_6520,N_6235,N_6332);
and U6521 (N_6521,N_6240,N_6283);
nor U6522 (N_6522,N_6263,N_6273);
nor U6523 (N_6523,N_6375,N_6229);
and U6524 (N_6524,N_6242,N_6210);
nand U6525 (N_6525,N_6257,N_6269);
nor U6526 (N_6526,N_6338,N_6280);
or U6527 (N_6527,N_6330,N_6342);
nand U6528 (N_6528,N_6348,N_6209);
nor U6529 (N_6529,N_6212,N_6340);
xnor U6530 (N_6530,N_6356,N_6343);
or U6531 (N_6531,N_6350,N_6326);
xor U6532 (N_6532,N_6323,N_6217);
nand U6533 (N_6533,N_6321,N_6238);
xor U6534 (N_6534,N_6320,N_6210);
xnor U6535 (N_6535,N_6358,N_6308);
or U6536 (N_6536,N_6298,N_6369);
nor U6537 (N_6537,N_6351,N_6397);
nand U6538 (N_6538,N_6220,N_6369);
xnor U6539 (N_6539,N_6356,N_6214);
or U6540 (N_6540,N_6205,N_6360);
nor U6541 (N_6541,N_6318,N_6264);
nand U6542 (N_6542,N_6215,N_6312);
and U6543 (N_6543,N_6334,N_6333);
and U6544 (N_6544,N_6286,N_6225);
nor U6545 (N_6545,N_6355,N_6286);
and U6546 (N_6546,N_6367,N_6234);
xnor U6547 (N_6547,N_6355,N_6324);
nor U6548 (N_6548,N_6271,N_6395);
and U6549 (N_6549,N_6364,N_6286);
or U6550 (N_6550,N_6251,N_6270);
and U6551 (N_6551,N_6212,N_6201);
or U6552 (N_6552,N_6352,N_6309);
nor U6553 (N_6553,N_6336,N_6278);
xnor U6554 (N_6554,N_6340,N_6248);
nand U6555 (N_6555,N_6311,N_6360);
nand U6556 (N_6556,N_6216,N_6252);
nand U6557 (N_6557,N_6272,N_6277);
or U6558 (N_6558,N_6362,N_6226);
and U6559 (N_6559,N_6247,N_6270);
nor U6560 (N_6560,N_6289,N_6398);
nor U6561 (N_6561,N_6209,N_6308);
nand U6562 (N_6562,N_6366,N_6398);
xnor U6563 (N_6563,N_6285,N_6394);
or U6564 (N_6564,N_6293,N_6281);
and U6565 (N_6565,N_6302,N_6332);
nand U6566 (N_6566,N_6334,N_6313);
and U6567 (N_6567,N_6324,N_6206);
and U6568 (N_6568,N_6282,N_6224);
or U6569 (N_6569,N_6236,N_6222);
or U6570 (N_6570,N_6209,N_6281);
and U6571 (N_6571,N_6288,N_6393);
nand U6572 (N_6572,N_6269,N_6300);
and U6573 (N_6573,N_6294,N_6284);
nand U6574 (N_6574,N_6226,N_6234);
xor U6575 (N_6575,N_6397,N_6226);
nor U6576 (N_6576,N_6202,N_6383);
nand U6577 (N_6577,N_6383,N_6254);
or U6578 (N_6578,N_6291,N_6285);
nand U6579 (N_6579,N_6356,N_6265);
nor U6580 (N_6580,N_6294,N_6316);
nand U6581 (N_6581,N_6232,N_6346);
nor U6582 (N_6582,N_6235,N_6264);
nor U6583 (N_6583,N_6261,N_6295);
or U6584 (N_6584,N_6378,N_6359);
nor U6585 (N_6585,N_6355,N_6238);
or U6586 (N_6586,N_6360,N_6365);
xnor U6587 (N_6587,N_6236,N_6342);
nor U6588 (N_6588,N_6284,N_6229);
and U6589 (N_6589,N_6239,N_6275);
nor U6590 (N_6590,N_6324,N_6205);
and U6591 (N_6591,N_6234,N_6206);
or U6592 (N_6592,N_6290,N_6311);
nand U6593 (N_6593,N_6248,N_6208);
or U6594 (N_6594,N_6262,N_6380);
or U6595 (N_6595,N_6256,N_6233);
or U6596 (N_6596,N_6235,N_6256);
and U6597 (N_6597,N_6376,N_6388);
and U6598 (N_6598,N_6311,N_6373);
or U6599 (N_6599,N_6287,N_6379);
nor U6600 (N_6600,N_6488,N_6575);
or U6601 (N_6601,N_6478,N_6454);
or U6602 (N_6602,N_6428,N_6576);
and U6603 (N_6603,N_6542,N_6494);
and U6604 (N_6604,N_6541,N_6501);
and U6605 (N_6605,N_6487,N_6432);
and U6606 (N_6606,N_6439,N_6555);
or U6607 (N_6607,N_6544,N_6512);
or U6608 (N_6608,N_6458,N_6513);
or U6609 (N_6609,N_6414,N_6580);
or U6610 (N_6610,N_6571,N_6453);
xnor U6611 (N_6611,N_6531,N_6450);
nor U6612 (N_6612,N_6586,N_6509);
or U6613 (N_6613,N_6517,N_6493);
nor U6614 (N_6614,N_6524,N_6441);
nor U6615 (N_6615,N_6537,N_6416);
or U6616 (N_6616,N_6594,N_6538);
and U6617 (N_6617,N_6449,N_6521);
and U6618 (N_6618,N_6406,N_6446);
and U6619 (N_6619,N_6456,N_6448);
or U6620 (N_6620,N_6426,N_6577);
or U6621 (N_6621,N_6435,N_6569);
nand U6622 (N_6622,N_6582,N_6529);
or U6623 (N_6623,N_6472,N_6503);
nor U6624 (N_6624,N_6451,N_6452);
nor U6625 (N_6625,N_6411,N_6417);
nand U6626 (N_6626,N_6405,N_6430);
nand U6627 (N_6627,N_6408,N_6560);
nand U6628 (N_6628,N_6404,N_6547);
or U6629 (N_6629,N_6465,N_6518);
and U6630 (N_6630,N_6588,N_6590);
nor U6631 (N_6631,N_6522,N_6457);
nor U6632 (N_6632,N_6539,N_6563);
nor U6633 (N_6633,N_6418,N_6483);
nor U6634 (N_6634,N_6486,N_6573);
nand U6635 (N_6635,N_6477,N_6445);
and U6636 (N_6636,N_6553,N_6427);
or U6637 (N_6637,N_6479,N_6419);
nand U6638 (N_6638,N_6460,N_6533);
nand U6639 (N_6639,N_6403,N_6402);
or U6640 (N_6640,N_6497,N_6559);
nor U6641 (N_6641,N_6558,N_6548);
or U6642 (N_6642,N_6455,N_6429);
xnor U6643 (N_6643,N_6506,N_6420);
and U6644 (N_6644,N_6526,N_6489);
or U6645 (N_6645,N_6587,N_6421);
or U6646 (N_6646,N_6438,N_6413);
xnor U6647 (N_6647,N_6476,N_6469);
nor U6648 (N_6648,N_6543,N_6474);
or U6649 (N_6649,N_6401,N_6583);
nand U6650 (N_6650,N_6515,N_6546);
xnor U6651 (N_6651,N_6447,N_6440);
and U6652 (N_6652,N_6527,N_6500);
nor U6653 (N_6653,N_6570,N_6484);
and U6654 (N_6654,N_6581,N_6467);
nand U6655 (N_6655,N_6572,N_6585);
nor U6656 (N_6656,N_6562,N_6597);
xor U6657 (N_6657,N_6525,N_6596);
xnor U6658 (N_6658,N_6473,N_6595);
and U6659 (N_6659,N_6519,N_6566);
and U6660 (N_6660,N_6498,N_6495);
and U6661 (N_6661,N_6514,N_6400);
nor U6662 (N_6662,N_6552,N_6464);
nand U6663 (N_6663,N_6584,N_6540);
and U6664 (N_6664,N_6530,N_6431);
xor U6665 (N_6665,N_6412,N_6567);
nor U6666 (N_6666,N_6554,N_6496);
and U6667 (N_6667,N_6545,N_6504);
nand U6668 (N_6668,N_6523,N_6511);
and U6669 (N_6669,N_6502,N_6499);
nand U6670 (N_6670,N_6550,N_6434);
nand U6671 (N_6671,N_6536,N_6425);
nor U6672 (N_6672,N_6437,N_6444);
or U6673 (N_6673,N_6507,N_6557);
or U6674 (N_6674,N_6564,N_6598);
and U6675 (N_6675,N_6505,N_6480);
nand U6676 (N_6676,N_6532,N_6459);
or U6677 (N_6677,N_6510,N_6466);
nor U6678 (N_6678,N_6574,N_6565);
nor U6679 (N_6679,N_6556,N_6520);
nand U6680 (N_6680,N_6599,N_6422);
nand U6681 (N_6681,N_6409,N_6485);
or U6682 (N_6682,N_6475,N_6463);
or U6683 (N_6683,N_6551,N_6508);
or U6684 (N_6684,N_6568,N_6535);
or U6685 (N_6685,N_6592,N_6462);
xor U6686 (N_6686,N_6491,N_6423);
and U6687 (N_6687,N_6415,N_6407);
xnor U6688 (N_6688,N_6516,N_6579);
nand U6689 (N_6689,N_6470,N_6468);
and U6690 (N_6690,N_6578,N_6482);
nand U6691 (N_6691,N_6589,N_6549);
or U6692 (N_6692,N_6436,N_6534);
nand U6693 (N_6693,N_6433,N_6410);
and U6694 (N_6694,N_6490,N_6492);
nor U6695 (N_6695,N_6471,N_6442);
nand U6696 (N_6696,N_6528,N_6424);
or U6697 (N_6697,N_6591,N_6461);
and U6698 (N_6698,N_6443,N_6481);
xor U6699 (N_6699,N_6593,N_6561);
or U6700 (N_6700,N_6429,N_6509);
nor U6701 (N_6701,N_6538,N_6491);
and U6702 (N_6702,N_6564,N_6553);
nor U6703 (N_6703,N_6573,N_6451);
nand U6704 (N_6704,N_6522,N_6431);
xor U6705 (N_6705,N_6464,N_6498);
nor U6706 (N_6706,N_6481,N_6462);
nor U6707 (N_6707,N_6418,N_6456);
nand U6708 (N_6708,N_6406,N_6545);
nand U6709 (N_6709,N_6421,N_6411);
and U6710 (N_6710,N_6495,N_6505);
nor U6711 (N_6711,N_6436,N_6525);
nor U6712 (N_6712,N_6482,N_6500);
or U6713 (N_6713,N_6468,N_6509);
or U6714 (N_6714,N_6416,N_6551);
xnor U6715 (N_6715,N_6503,N_6555);
nor U6716 (N_6716,N_6407,N_6591);
nand U6717 (N_6717,N_6574,N_6492);
or U6718 (N_6718,N_6493,N_6525);
nor U6719 (N_6719,N_6435,N_6430);
nand U6720 (N_6720,N_6535,N_6539);
nand U6721 (N_6721,N_6550,N_6566);
and U6722 (N_6722,N_6402,N_6512);
and U6723 (N_6723,N_6416,N_6577);
nor U6724 (N_6724,N_6538,N_6544);
nand U6725 (N_6725,N_6504,N_6543);
and U6726 (N_6726,N_6585,N_6546);
nor U6727 (N_6727,N_6476,N_6561);
or U6728 (N_6728,N_6468,N_6452);
nand U6729 (N_6729,N_6594,N_6485);
nor U6730 (N_6730,N_6595,N_6437);
nand U6731 (N_6731,N_6445,N_6557);
and U6732 (N_6732,N_6528,N_6445);
nor U6733 (N_6733,N_6410,N_6503);
nor U6734 (N_6734,N_6553,N_6425);
nor U6735 (N_6735,N_6412,N_6486);
or U6736 (N_6736,N_6486,N_6482);
and U6737 (N_6737,N_6435,N_6516);
nand U6738 (N_6738,N_6505,N_6463);
nand U6739 (N_6739,N_6581,N_6512);
or U6740 (N_6740,N_6514,N_6435);
or U6741 (N_6741,N_6416,N_6435);
or U6742 (N_6742,N_6516,N_6455);
or U6743 (N_6743,N_6428,N_6596);
nand U6744 (N_6744,N_6554,N_6411);
nand U6745 (N_6745,N_6423,N_6524);
nand U6746 (N_6746,N_6524,N_6543);
and U6747 (N_6747,N_6562,N_6576);
and U6748 (N_6748,N_6466,N_6443);
or U6749 (N_6749,N_6445,N_6543);
xor U6750 (N_6750,N_6466,N_6486);
nor U6751 (N_6751,N_6551,N_6481);
nor U6752 (N_6752,N_6584,N_6594);
nand U6753 (N_6753,N_6509,N_6427);
nor U6754 (N_6754,N_6511,N_6591);
nand U6755 (N_6755,N_6421,N_6557);
or U6756 (N_6756,N_6453,N_6515);
and U6757 (N_6757,N_6521,N_6552);
or U6758 (N_6758,N_6569,N_6414);
nand U6759 (N_6759,N_6464,N_6426);
or U6760 (N_6760,N_6451,N_6471);
nor U6761 (N_6761,N_6574,N_6543);
nand U6762 (N_6762,N_6498,N_6429);
or U6763 (N_6763,N_6407,N_6590);
or U6764 (N_6764,N_6450,N_6537);
nand U6765 (N_6765,N_6496,N_6426);
and U6766 (N_6766,N_6423,N_6509);
or U6767 (N_6767,N_6598,N_6462);
and U6768 (N_6768,N_6520,N_6584);
or U6769 (N_6769,N_6454,N_6518);
nor U6770 (N_6770,N_6489,N_6473);
nand U6771 (N_6771,N_6427,N_6578);
nor U6772 (N_6772,N_6541,N_6419);
and U6773 (N_6773,N_6519,N_6482);
or U6774 (N_6774,N_6507,N_6541);
nor U6775 (N_6775,N_6567,N_6425);
and U6776 (N_6776,N_6551,N_6512);
nor U6777 (N_6777,N_6468,N_6483);
nor U6778 (N_6778,N_6492,N_6445);
nor U6779 (N_6779,N_6487,N_6544);
or U6780 (N_6780,N_6557,N_6591);
or U6781 (N_6781,N_6581,N_6571);
nand U6782 (N_6782,N_6586,N_6493);
or U6783 (N_6783,N_6482,N_6401);
or U6784 (N_6784,N_6475,N_6505);
and U6785 (N_6785,N_6526,N_6556);
nand U6786 (N_6786,N_6528,N_6565);
xor U6787 (N_6787,N_6503,N_6445);
xor U6788 (N_6788,N_6436,N_6533);
nor U6789 (N_6789,N_6568,N_6419);
and U6790 (N_6790,N_6461,N_6415);
and U6791 (N_6791,N_6493,N_6432);
nand U6792 (N_6792,N_6528,N_6413);
nor U6793 (N_6793,N_6511,N_6595);
or U6794 (N_6794,N_6428,N_6475);
or U6795 (N_6795,N_6443,N_6520);
and U6796 (N_6796,N_6532,N_6405);
nor U6797 (N_6797,N_6513,N_6461);
or U6798 (N_6798,N_6421,N_6524);
or U6799 (N_6799,N_6445,N_6420);
nor U6800 (N_6800,N_6753,N_6745);
or U6801 (N_6801,N_6773,N_6762);
or U6802 (N_6802,N_6694,N_6658);
and U6803 (N_6803,N_6603,N_6643);
nand U6804 (N_6804,N_6626,N_6737);
nand U6805 (N_6805,N_6713,N_6648);
and U6806 (N_6806,N_6647,N_6724);
and U6807 (N_6807,N_6665,N_6661);
and U6808 (N_6808,N_6707,N_6664);
nor U6809 (N_6809,N_6675,N_6611);
or U6810 (N_6810,N_6761,N_6621);
nor U6811 (N_6811,N_6774,N_6788);
nor U6812 (N_6812,N_6620,N_6715);
or U6813 (N_6813,N_6652,N_6623);
or U6814 (N_6814,N_6628,N_6786);
and U6815 (N_6815,N_6627,N_6601);
nand U6816 (N_6816,N_6784,N_6711);
and U6817 (N_6817,N_6638,N_6792);
and U6818 (N_6818,N_6738,N_6624);
or U6819 (N_6819,N_6654,N_6755);
or U6820 (N_6820,N_6723,N_6785);
xnor U6821 (N_6821,N_6746,N_6653);
nand U6822 (N_6822,N_6789,N_6778);
xnor U6823 (N_6823,N_6633,N_6776);
nor U6824 (N_6824,N_6607,N_6717);
nor U6825 (N_6825,N_6646,N_6709);
nor U6826 (N_6826,N_6677,N_6605);
and U6827 (N_6827,N_6615,N_6725);
and U6828 (N_6828,N_6769,N_6649);
nor U6829 (N_6829,N_6610,N_6650);
or U6830 (N_6830,N_6671,N_6760);
nor U6831 (N_6831,N_6766,N_6606);
and U6832 (N_6832,N_6759,N_6630);
and U6833 (N_6833,N_6747,N_6680);
or U6834 (N_6834,N_6749,N_6732);
and U6835 (N_6835,N_6667,N_6701);
nor U6836 (N_6836,N_6678,N_6689);
and U6837 (N_6837,N_6696,N_6683);
or U6838 (N_6838,N_6673,N_6632);
nand U6839 (N_6839,N_6756,N_6791);
nor U6840 (N_6840,N_6794,N_6736);
xor U6841 (N_6841,N_6614,N_6674);
nor U6842 (N_6842,N_6750,N_6751);
or U6843 (N_6843,N_6693,N_6681);
nand U6844 (N_6844,N_6655,N_6799);
nand U6845 (N_6845,N_6763,N_6739);
and U6846 (N_6846,N_6775,N_6619);
or U6847 (N_6847,N_6625,N_6727);
xnor U6848 (N_6848,N_6734,N_6631);
nor U6849 (N_6849,N_6612,N_6783);
and U6850 (N_6850,N_6659,N_6741);
and U6851 (N_6851,N_6604,N_6795);
xnor U6852 (N_6852,N_6733,N_6726);
or U6853 (N_6853,N_6702,N_6682);
or U6854 (N_6854,N_6634,N_6771);
or U6855 (N_6855,N_6704,N_6719);
nand U6856 (N_6856,N_6728,N_6768);
xor U6857 (N_6857,N_6714,N_6635);
nand U6858 (N_6858,N_6748,N_6669);
or U6859 (N_6859,N_6642,N_6720);
or U6860 (N_6860,N_6796,N_6740);
and U6861 (N_6861,N_6797,N_6721);
and U6862 (N_6862,N_6687,N_6684);
nand U6863 (N_6863,N_6645,N_6699);
nand U6864 (N_6864,N_6765,N_6668);
nor U6865 (N_6865,N_6608,N_6698);
nor U6866 (N_6866,N_6708,N_6676);
and U6867 (N_6867,N_6657,N_6764);
and U6868 (N_6868,N_6710,N_6793);
or U6869 (N_6869,N_6690,N_6757);
nor U6870 (N_6870,N_6729,N_6618);
or U6871 (N_6871,N_6679,N_6718);
or U6872 (N_6872,N_6735,N_6644);
and U6873 (N_6873,N_6666,N_6656);
or U6874 (N_6874,N_6706,N_6613);
or U6875 (N_6875,N_6617,N_6744);
nor U6876 (N_6876,N_6663,N_6782);
nor U6877 (N_6877,N_6798,N_6700);
nand U6878 (N_6878,N_6742,N_6754);
nand U6879 (N_6879,N_6790,N_6780);
and U6880 (N_6880,N_6767,N_6770);
nor U6881 (N_6881,N_6705,N_6730);
or U6882 (N_6882,N_6772,N_6672);
xnor U6883 (N_6883,N_6660,N_6692);
nand U6884 (N_6884,N_6688,N_6691);
or U6885 (N_6885,N_6651,N_6777);
xnor U6886 (N_6886,N_6722,N_6602);
and U6887 (N_6887,N_6758,N_6712);
nor U6888 (N_6888,N_6752,N_6670);
nand U6889 (N_6889,N_6686,N_6781);
nor U6890 (N_6890,N_6616,N_6609);
or U6891 (N_6891,N_6743,N_6622);
xnor U6892 (N_6892,N_6731,N_6641);
xnor U6893 (N_6893,N_6695,N_6787);
xnor U6894 (N_6894,N_6640,N_6779);
xor U6895 (N_6895,N_6600,N_6639);
nand U6896 (N_6896,N_6637,N_6662);
nand U6897 (N_6897,N_6636,N_6697);
or U6898 (N_6898,N_6716,N_6629);
or U6899 (N_6899,N_6685,N_6703);
and U6900 (N_6900,N_6739,N_6760);
nand U6901 (N_6901,N_6659,N_6695);
xnor U6902 (N_6902,N_6603,N_6660);
nand U6903 (N_6903,N_6679,N_6603);
nand U6904 (N_6904,N_6718,N_6716);
nand U6905 (N_6905,N_6627,N_6701);
and U6906 (N_6906,N_6790,N_6728);
nor U6907 (N_6907,N_6676,N_6771);
and U6908 (N_6908,N_6663,N_6778);
and U6909 (N_6909,N_6646,N_6688);
nand U6910 (N_6910,N_6663,N_6787);
or U6911 (N_6911,N_6787,N_6777);
and U6912 (N_6912,N_6656,N_6700);
nor U6913 (N_6913,N_6675,N_6729);
nand U6914 (N_6914,N_6635,N_6660);
or U6915 (N_6915,N_6632,N_6694);
nor U6916 (N_6916,N_6741,N_6714);
or U6917 (N_6917,N_6732,N_6700);
nor U6918 (N_6918,N_6653,N_6754);
and U6919 (N_6919,N_6714,N_6697);
and U6920 (N_6920,N_6733,N_6620);
nor U6921 (N_6921,N_6783,N_6608);
and U6922 (N_6922,N_6736,N_6601);
and U6923 (N_6923,N_6718,N_6696);
or U6924 (N_6924,N_6795,N_6741);
xor U6925 (N_6925,N_6615,N_6742);
nand U6926 (N_6926,N_6637,N_6779);
nand U6927 (N_6927,N_6718,N_6684);
nor U6928 (N_6928,N_6778,N_6620);
nand U6929 (N_6929,N_6767,N_6751);
or U6930 (N_6930,N_6764,N_6625);
nand U6931 (N_6931,N_6760,N_6619);
nand U6932 (N_6932,N_6670,N_6644);
or U6933 (N_6933,N_6654,N_6649);
or U6934 (N_6934,N_6708,N_6667);
nand U6935 (N_6935,N_6669,N_6666);
nand U6936 (N_6936,N_6660,N_6661);
or U6937 (N_6937,N_6720,N_6699);
or U6938 (N_6938,N_6676,N_6680);
nor U6939 (N_6939,N_6675,N_6766);
nor U6940 (N_6940,N_6675,N_6776);
nor U6941 (N_6941,N_6621,N_6693);
xnor U6942 (N_6942,N_6628,N_6662);
or U6943 (N_6943,N_6773,N_6797);
nor U6944 (N_6944,N_6669,N_6798);
and U6945 (N_6945,N_6782,N_6728);
nor U6946 (N_6946,N_6682,N_6759);
or U6947 (N_6947,N_6778,N_6603);
nand U6948 (N_6948,N_6632,N_6601);
or U6949 (N_6949,N_6793,N_6693);
nand U6950 (N_6950,N_6642,N_6794);
and U6951 (N_6951,N_6646,N_6729);
and U6952 (N_6952,N_6643,N_6669);
and U6953 (N_6953,N_6744,N_6761);
xor U6954 (N_6954,N_6783,N_6703);
or U6955 (N_6955,N_6763,N_6729);
or U6956 (N_6956,N_6618,N_6680);
nor U6957 (N_6957,N_6627,N_6635);
nand U6958 (N_6958,N_6682,N_6730);
nor U6959 (N_6959,N_6610,N_6612);
or U6960 (N_6960,N_6770,N_6785);
and U6961 (N_6961,N_6742,N_6698);
or U6962 (N_6962,N_6725,N_6787);
or U6963 (N_6963,N_6639,N_6667);
nand U6964 (N_6964,N_6776,N_6638);
and U6965 (N_6965,N_6748,N_6730);
nor U6966 (N_6966,N_6692,N_6646);
or U6967 (N_6967,N_6798,N_6727);
nor U6968 (N_6968,N_6797,N_6710);
and U6969 (N_6969,N_6780,N_6797);
and U6970 (N_6970,N_6785,N_6694);
nor U6971 (N_6971,N_6718,N_6773);
and U6972 (N_6972,N_6656,N_6789);
nand U6973 (N_6973,N_6729,N_6792);
nor U6974 (N_6974,N_6611,N_6780);
or U6975 (N_6975,N_6767,N_6600);
nor U6976 (N_6976,N_6651,N_6731);
nor U6977 (N_6977,N_6661,N_6606);
nand U6978 (N_6978,N_6668,N_6730);
and U6979 (N_6979,N_6722,N_6762);
nand U6980 (N_6980,N_6793,N_6774);
xnor U6981 (N_6981,N_6770,N_6769);
xnor U6982 (N_6982,N_6650,N_6755);
nor U6983 (N_6983,N_6623,N_6757);
xnor U6984 (N_6984,N_6622,N_6707);
nor U6985 (N_6985,N_6671,N_6759);
nor U6986 (N_6986,N_6749,N_6648);
nor U6987 (N_6987,N_6613,N_6795);
and U6988 (N_6988,N_6695,N_6771);
or U6989 (N_6989,N_6679,N_6684);
nor U6990 (N_6990,N_6750,N_6743);
nor U6991 (N_6991,N_6607,N_6671);
or U6992 (N_6992,N_6607,N_6767);
xor U6993 (N_6993,N_6607,N_6694);
nor U6994 (N_6994,N_6795,N_6699);
nand U6995 (N_6995,N_6630,N_6699);
nor U6996 (N_6996,N_6716,N_6796);
xnor U6997 (N_6997,N_6768,N_6688);
or U6998 (N_6998,N_6606,N_6754);
or U6999 (N_6999,N_6662,N_6654);
xnor U7000 (N_7000,N_6875,N_6893);
or U7001 (N_7001,N_6911,N_6931);
nand U7002 (N_7002,N_6936,N_6957);
nand U7003 (N_7003,N_6853,N_6953);
nor U7004 (N_7004,N_6909,N_6955);
nand U7005 (N_7005,N_6995,N_6878);
nand U7006 (N_7006,N_6806,N_6982);
and U7007 (N_7007,N_6869,N_6981);
xnor U7008 (N_7008,N_6857,N_6938);
nand U7009 (N_7009,N_6898,N_6983);
nor U7010 (N_7010,N_6821,N_6824);
and U7011 (N_7011,N_6901,N_6833);
and U7012 (N_7012,N_6926,N_6977);
and U7013 (N_7013,N_6949,N_6876);
or U7014 (N_7014,N_6945,N_6894);
nand U7015 (N_7015,N_6888,N_6944);
and U7016 (N_7016,N_6823,N_6819);
and U7017 (N_7017,N_6854,N_6850);
nor U7018 (N_7018,N_6808,N_6810);
and U7019 (N_7019,N_6979,N_6951);
and U7020 (N_7020,N_6848,N_6803);
nand U7021 (N_7021,N_6969,N_6891);
nand U7022 (N_7022,N_6826,N_6907);
nand U7023 (N_7023,N_6834,N_6801);
or U7024 (N_7024,N_6851,N_6975);
xnor U7025 (N_7025,N_6974,N_6813);
nor U7026 (N_7026,N_6948,N_6989);
nand U7027 (N_7027,N_6871,N_6914);
or U7028 (N_7028,N_6943,N_6861);
nor U7029 (N_7029,N_6809,N_6913);
nand U7030 (N_7030,N_6965,N_6908);
and U7031 (N_7031,N_6916,N_6929);
or U7032 (N_7032,N_6877,N_6827);
nand U7033 (N_7033,N_6815,N_6902);
nor U7034 (N_7034,N_6988,N_6831);
xnor U7035 (N_7035,N_6959,N_6941);
or U7036 (N_7036,N_6889,N_6807);
or U7037 (N_7037,N_6840,N_6990);
nor U7038 (N_7038,N_6912,N_6855);
nor U7039 (N_7039,N_6884,N_6994);
nor U7040 (N_7040,N_6997,N_6930);
nor U7041 (N_7041,N_6906,N_6814);
nor U7042 (N_7042,N_6865,N_6842);
or U7043 (N_7043,N_6946,N_6958);
and U7044 (N_7044,N_6895,N_6844);
nor U7045 (N_7045,N_6852,N_6887);
nor U7046 (N_7046,N_6919,N_6973);
xor U7047 (N_7047,N_6918,N_6942);
nand U7048 (N_7048,N_6830,N_6890);
nor U7049 (N_7049,N_6934,N_6999);
xnor U7050 (N_7050,N_6864,N_6950);
or U7051 (N_7051,N_6804,N_6952);
nand U7052 (N_7052,N_6874,N_6935);
and U7053 (N_7053,N_6885,N_6835);
nand U7054 (N_7054,N_6863,N_6825);
or U7055 (N_7055,N_6921,N_6928);
nor U7056 (N_7056,N_6933,N_6984);
nor U7057 (N_7057,N_6968,N_6961);
xor U7058 (N_7058,N_6978,N_6883);
xnor U7059 (N_7059,N_6829,N_6882);
and U7060 (N_7060,N_6956,N_6910);
and U7061 (N_7061,N_6881,N_6980);
nor U7062 (N_7062,N_6828,N_6860);
nor U7063 (N_7063,N_6986,N_6837);
or U7064 (N_7064,N_6900,N_6971);
or U7065 (N_7065,N_6904,N_6866);
and U7066 (N_7066,N_6976,N_6924);
nor U7067 (N_7067,N_6917,N_6856);
and U7068 (N_7068,N_6870,N_6843);
or U7069 (N_7069,N_6873,N_6925);
nand U7070 (N_7070,N_6927,N_6880);
and U7071 (N_7071,N_6940,N_6817);
xor U7072 (N_7072,N_6872,N_6964);
nor U7073 (N_7073,N_6838,N_6867);
or U7074 (N_7074,N_6845,N_6998);
nand U7075 (N_7075,N_6841,N_6996);
or U7076 (N_7076,N_6915,N_6954);
or U7077 (N_7077,N_6920,N_6816);
and U7078 (N_7078,N_6993,N_6822);
nor U7079 (N_7079,N_6939,N_6947);
nand U7080 (N_7080,N_6839,N_6820);
nor U7081 (N_7081,N_6897,N_6987);
and U7082 (N_7082,N_6905,N_6991);
nor U7083 (N_7083,N_6862,N_6892);
or U7084 (N_7084,N_6992,N_6818);
xor U7085 (N_7085,N_6879,N_6812);
or U7086 (N_7086,N_6847,N_6858);
and U7087 (N_7087,N_6868,N_6849);
nor U7088 (N_7088,N_6937,N_6923);
and U7089 (N_7089,N_6811,N_6899);
xor U7090 (N_7090,N_6967,N_6960);
nand U7091 (N_7091,N_6896,N_6859);
and U7092 (N_7092,N_6903,N_6962);
and U7093 (N_7093,N_6922,N_6805);
or U7094 (N_7094,N_6846,N_6972);
nor U7095 (N_7095,N_6836,N_6985);
nand U7096 (N_7096,N_6966,N_6963);
nor U7097 (N_7097,N_6800,N_6832);
and U7098 (N_7098,N_6970,N_6932);
nand U7099 (N_7099,N_6802,N_6886);
and U7100 (N_7100,N_6893,N_6870);
nand U7101 (N_7101,N_6898,N_6997);
or U7102 (N_7102,N_6946,N_6939);
xnor U7103 (N_7103,N_6942,N_6919);
nand U7104 (N_7104,N_6814,N_6868);
nor U7105 (N_7105,N_6900,N_6929);
or U7106 (N_7106,N_6976,N_6979);
nand U7107 (N_7107,N_6954,N_6841);
nand U7108 (N_7108,N_6843,N_6881);
nand U7109 (N_7109,N_6949,N_6852);
and U7110 (N_7110,N_6917,N_6999);
and U7111 (N_7111,N_6877,N_6985);
nor U7112 (N_7112,N_6856,N_6925);
or U7113 (N_7113,N_6816,N_6917);
and U7114 (N_7114,N_6809,N_6999);
nand U7115 (N_7115,N_6911,N_6926);
xnor U7116 (N_7116,N_6906,N_6981);
nand U7117 (N_7117,N_6976,N_6948);
or U7118 (N_7118,N_6987,N_6880);
and U7119 (N_7119,N_6961,N_6819);
and U7120 (N_7120,N_6841,N_6979);
nor U7121 (N_7121,N_6910,N_6899);
and U7122 (N_7122,N_6843,N_6912);
and U7123 (N_7123,N_6922,N_6873);
nand U7124 (N_7124,N_6881,N_6926);
xnor U7125 (N_7125,N_6872,N_6885);
and U7126 (N_7126,N_6842,N_6961);
or U7127 (N_7127,N_6829,N_6854);
nand U7128 (N_7128,N_6888,N_6866);
nand U7129 (N_7129,N_6801,N_6822);
and U7130 (N_7130,N_6925,N_6853);
nand U7131 (N_7131,N_6802,N_6990);
and U7132 (N_7132,N_6921,N_6981);
and U7133 (N_7133,N_6862,N_6878);
nand U7134 (N_7134,N_6992,N_6843);
xor U7135 (N_7135,N_6839,N_6805);
or U7136 (N_7136,N_6935,N_6886);
nor U7137 (N_7137,N_6836,N_6875);
nand U7138 (N_7138,N_6929,N_6837);
nor U7139 (N_7139,N_6976,N_6827);
and U7140 (N_7140,N_6852,N_6846);
xor U7141 (N_7141,N_6957,N_6810);
or U7142 (N_7142,N_6935,N_6966);
and U7143 (N_7143,N_6879,N_6945);
or U7144 (N_7144,N_6944,N_6831);
and U7145 (N_7145,N_6834,N_6927);
or U7146 (N_7146,N_6965,N_6849);
or U7147 (N_7147,N_6916,N_6924);
nand U7148 (N_7148,N_6894,N_6985);
or U7149 (N_7149,N_6927,N_6975);
nor U7150 (N_7150,N_6821,N_6839);
and U7151 (N_7151,N_6923,N_6834);
nor U7152 (N_7152,N_6918,N_6896);
xor U7153 (N_7153,N_6957,N_6972);
nand U7154 (N_7154,N_6994,N_6984);
nor U7155 (N_7155,N_6842,N_6932);
and U7156 (N_7156,N_6800,N_6855);
or U7157 (N_7157,N_6991,N_6913);
nor U7158 (N_7158,N_6950,N_6973);
and U7159 (N_7159,N_6972,N_6922);
nor U7160 (N_7160,N_6893,N_6966);
or U7161 (N_7161,N_6971,N_6931);
or U7162 (N_7162,N_6852,N_6939);
or U7163 (N_7163,N_6919,N_6926);
or U7164 (N_7164,N_6979,N_6872);
nor U7165 (N_7165,N_6897,N_6953);
and U7166 (N_7166,N_6999,N_6828);
or U7167 (N_7167,N_6929,N_6986);
and U7168 (N_7168,N_6934,N_6919);
and U7169 (N_7169,N_6882,N_6804);
and U7170 (N_7170,N_6915,N_6822);
nor U7171 (N_7171,N_6941,N_6927);
nand U7172 (N_7172,N_6846,N_6917);
and U7173 (N_7173,N_6947,N_6865);
and U7174 (N_7174,N_6859,N_6909);
and U7175 (N_7175,N_6900,N_6844);
and U7176 (N_7176,N_6931,N_6807);
or U7177 (N_7177,N_6846,N_6847);
nand U7178 (N_7178,N_6872,N_6909);
or U7179 (N_7179,N_6908,N_6987);
xnor U7180 (N_7180,N_6900,N_6842);
or U7181 (N_7181,N_6812,N_6917);
xor U7182 (N_7182,N_6834,N_6950);
nand U7183 (N_7183,N_6866,N_6917);
or U7184 (N_7184,N_6886,N_6894);
and U7185 (N_7185,N_6842,N_6846);
nor U7186 (N_7186,N_6991,N_6963);
or U7187 (N_7187,N_6856,N_6997);
xor U7188 (N_7188,N_6975,N_6918);
nand U7189 (N_7189,N_6889,N_6981);
xor U7190 (N_7190,N_6930,N_6884);
nor U7191 (N_7191,N_6981,N_6888);
nand U7192 (N_7192,N_6819,N_6907);
or U7193 (N_7193,N_6887,N_6918);
nand U7194 (N_7194,N_6832,N_6850);
xor U7195 (N_7195,N_6985,N_6815);
nor U7196 (N_7196,N_6887,N_6925);
nand U7197 (N_7197,N_6917,N_6901);
nand U7198 (N_7198,N_6957,N_6953);
nor U7199 (N_7199,N_6823,N_6942);
and U7200 (N_7200,N_7199,N_7028);
xor U7201 (N_7201,N_7018,N_7169);
nand U7202 (N_7202,N_7163,N_7086);
nand U7203 (N_7203,N_7145,N_7031);
nor U7204 (N_7204,N_7139,N_7006);
or U7205 (N_7205,N_7111,N_7188);
nand U7206 (N_7206,N_7122,N_7143);
nand U7207 (N_7207,N_7036,N_7053);
xor U7208 (N_7208,N_7083,N_7013);
nand U7209 (N_7209,N_7003,N_7118);
or U7210 (N_7210,N_7116,N_7007);
xor U7211 (N_7211,N_7101,N_7113);
and U7212 (N_7212,N_7121,N_7161);
and U7213 (N_7213,N_7150,N_7021);
nand U7214 (N_7214,N_7195,N_7187);
and U7215 (N_7215,N_7160,N_7008);
xnor U7216 (N_7216,N_7148,N_7173);
xnor U7217 (N_7217,N_7040,N_7076);
xor U7218 (N_7218,N_7000,N_7067);
nand U7219 (N_7219,N_7016,N_7181);
nand U7220 (N_7220,N_7012,N_7130);
and U7221 (N_7221,N_7092,N_7105);
and U7222 (N_7222,N_7142,N_7140);
and U7223 (N_7223,N_7131,N_7029);
and U7224 (N_7224,N_7175,N_7151);
nor U7225 (N_7225,N_7049,N_7055);
nor U7226 (N_7226,N_7088,N_7011);
nand U7227 (N_7227,N_7048,N_7179);
nor U7228 (N_7228,N_7002,N_7112);
nor U7229 (N_7229,N_7058,N_7107);
nor U7230 (N_7230,N_7196,N_7070);
nor U7231 (N_7231,N_7198,N_7068);
and U7232 (N_7232,N_7132,N_7156);
nor U7233 (N_7233,N_7126,N_7050);
or U7234 (N_7234,N_7004,N_7194);
nor U7235 (N_7235,N_7104,N_7197);
nand U7236 (N_7236,N_7165,N_7082);
nand U7237 (N_7237,N_7157,N_7158);
and U7238 (N_7238,N_7176,N_7017);
or U7239 (N_7239,N_7174,N_7026);
xnor U7240 (N_7240,N_7098,N_7046);
nand U7241 (N_7241,N_7103,N_7167);
nor U7242 (N_7242,N_7091,N_7193);
nand U7243 (N_7243,N_7095,N_7071);
or U7244 (N_7244,N_7035,N_7033);
or U7245 (N_7245,N_7001,N_7037);
and U7246 (N_7246,N_7185,N_7152);
and U7247 (N_7247,N_7032,N_7009);
nor U7248 (N_7248,N_7024,N_7099);
nor U7249 (N_7249,N_7062,N_7154);
and U7250 (N_7250,N_7030,N_7178);
nor U7251 (N_7251,N_7138,N_7072);
nor U7252 (N_7252,N_7096,N_7190);
nor U7253 (N_7253,N_7078,N_7124);
nor U7254 (N_7254,N_7061,N_7084);
and U7255 (N_7255,N_7039,N_7019);
nor U7256 (N_7256,N_7162,N_7100);
or U7257 (N_7257,N_7115,N_7109);
nor U7258 (N_7258,N_7051,N_7184);
and U7259 (N_7259,N_7022,N_7056);
or U7260 (N_7260,N_7075,N_7054);
nand U7261 (N_7261,N_7135,N_7020);
nand U7262 (N_7262,N_7066,N_7166);
nand U7263 (N_7263,N_7117,N_7069);
nand U7264 (N_7264,N_7114,N_7047);
nand U7265 (N_7265,N_7044,N_7159);
xnor U7266 (N_7266,N_7149,N_7106);
or U7267 (N_7267,N_7010,N_7129);
nor U7268 (N_7268,N_7125,N_7089);
and U7269 (N_7269,N_7063,N_7171);
or U7270 (N_7270,N_7041,N_7141);
nand U7271 (N_7271,N_7186,N_7108);
nand U7272 (N_7272,N_7043,N_7128);
nor U7273 (N_7273,N_7042,N_7177);
or U7274 (N_7274,N_7064,N_7081);
and U7275 (N_7275,N_7182,N_7133);
and U7276 (N_7276,N_7085,N_7180);
nor U7277 (N_7277,N_7155,N_7144);
and U7278 (N_7278,N_7090,N_7102);
nor U7279 (N_7279,N_7015,N_7183);
nor U7280 (N_7280,N_7060,N_7038);
nand U7281 (N_7281,N_7025,N_7170);
nand U7282 (N_7282,N_7059,N_7146);
or U7283 (N_7283,N_7168,N_7034);
and U7284 (N_7284,N_7110,N_7191);
nor U7285 (N_7285,N_7087,N_7014);
nor U7286 (N_7286,N_7123,N_7192);
nor U7287 (N_7287,N_7045,N_7093);
or U7288 (N_7288,N_7052,N_7134);
or U7289 (N_7289,N_7080,N_7074);
or U7290 (N_7290,N_7094,N_7065);
xor U7291 (N_7291,N_7120,N_7077);
nor U7292 (N_7292,N_7189,N_7136);
and U7293 (N_7293,N_7005,N_7153);
or U7294 (N_7294,N_7023,N_7147);
nand U7295 (N_7295,N_7119,N_7127);
and U7296 (N_7296,N_7097,N_7073);
nor U7297 (N_7297,N_7057,N_7172);
xnor U7298 (N_7298,N_7164,N_7137);
and U7299 (N_7299,N_7027,N_7079);
nor U7300 (N_7300,N_7076,N_7068);
or U7301 (N_7301,N_7027,N_7090);
nand U7302 (N_7302,N_7012,N_7095);
nor U7303 (N_7303,N_7023,N_7007);
and U7304 (N_7304,N_7092,N_7193);
nor U7305 (N_7305,N_7092,N_7143);
and U7306 (N_7306,N_7152,N_7183);
nor U7307 (N_7307,N_7172,N_7166);
nor U7308 (N_7308,N_7173,N_7143);
nand U7309 (N_7309,N_7113,N_7029);
and U7310 (N_7310,N_7096,N_7018);
or U7311 (N_7311,N_7080,N_7086);
nand U7312 (N_7312,N_7119,N_7107);
or U7313 (N_7313,N_7174,N_7017);
nand U7314 (N_7314,N_7132,N_7040);
nand U7315 (N_7315,N_7049,N_7022);
nor U7316 (N_7316,N_7055,N_7097);
and U7317 (N_7317,N_7015,N_7111);
nor U7318 (N_7318,N_7189,N_7098);
xnor U7319 (N_7319,N_7196,N_7045);
nor U7320 (N_7320,N_7078,N_7009);
nand U7321 (N_7321,N_7176,N_7138);
nor U7322 (N_7322,N_7197,N_7113);
nand U7323 (N_7323,N_7193,N_7103);
xnor U7324 (N_7324,N_7107,N_7100);
nor U7325 (N_7325,N_7139,N_7197);
and U7326 (N_7326,N_7112,N_7101);
nand U7327 (N_7327,N_7173,N_7038);
or U7328 (N_7328,N_7078,N_7125);
xnor U7329 (N_7329,N_7013,N_7085);
and U7330 (N_7330,N_7028,N_7122);
and U7331 (N_7331,N_7126,N_7143);
or U7332 (N_7332,N_7042,N_7135);
or U7333 (N_7333,N_7008,N_7017);
nor U7334 (N_7334,N_7165,N_7023);
nor U7335 (N_7335,N_7066,N_7021);
or U7336 (N_7336,N_7108,N_7194);
xnor U7337 (N_7337,N_7175,N_7178);
nand U7338 (N_7338,N_7001,N_7040);
nor U7339 (N_7339,N_7199,N_7033);
xnor U7340 (N_7340,N_7082,N_7034);
or U7341 (N_7341,N_7128,N_7049);
or U7342 (N_7342,N_7117,N_7081);
nor U7343 (N_7343,N_7134,N_7010);
nand U7344 (N_7344,N_7165,N_7043);
or U7345 (N_7345,N_7063,N_7169);
nand U7346 (N_7346,N_7108,N_7138);
nand U7347 (N_7347,N_7125,N_7084);
and U7348 (N_7348,N_7155,N_7027);
and U7349 (N_7349,N_7081,N_7123);
or U7350 (N_7350,N_7100,N_7194);
and U7351 (N_7351,N_7093,N_7028);
nand U7352 (N_7352,N_7072,N_7152);
nand U7353 (N_7353,N_7153,N_7108);
xor U7354 (N_7354,N_7015,N_7069);
and U7355 (N_7355,N_7063,N_7099);
and U7356 (N_7356,N_7005,N_7195);
nand U7357 (N_7357,N_7172,N_7198);
nand U7358 (N_7358,N_7120,N_7107);
nor U7359 (N_7359,N_7001,N_7195);
nand U7360 (N_7360,N_7077,N_7102);
or U7361 (N_7361,N_7184,N_7045);
nand U7362 (N_7362,N_7053,N_7136);
nor U7363 (N_7363,N_7087,N_7156);
nand U7364 (N_7364,N_7058,N_7129);
nor U7365 (N_7365,N_7000,N_7196);
or U7366 (N_7366,N_7075,N_7027);
and U7367 (N_7367,N_7066,N_7065);
and U7368 (N_7368,N_7179,N_7169);
nand U7369 (N_7369,N_7013,N_7090);
nor U7370 (N_7370,N_7023,N_7168);
nor U7371 (N_7371,N_7116,N_7135);
or U7372 (N_7372,N_7170,N_7074);
nand U7373 (N_7373,N_7041,N_7147);
or U7374 (N_7374,N_7062,N_7045);
and U7375 (N_7375,N_7141,N_7107);
nor U7376 (N_7376,N_7080,N_7131);
or U7377 (N_7377,N_7149,N_7105);
nor U7378 (N_7378,N_7084,N_7141);
and U7379 (N_7379,N_7044,N_7137);
nor U7380 (N_7380,N_7094,N_7187);
and U7381 (N_7381,N_7115,N_7185);
or U7382 (N_7382,N_7073,N_7050);
nand U7383 (N_7383,N_7115,N_7193);
nand U7384 (N_7384,N_7000,N_7086);
and U7385 (N_7385,N_7049,N_7141);
and U7386 (N_7386,N_7152,N_7102);
and U7387 (N_7387,N_7040,N_7004);
or U7388 (N_7388,N_7165,N_7084);
nand U7389 (N_7389,N_7094,N_7177);
or U7390 (N_7390,N_7151,N_7125);
or U7391 (N_7391,N_7031,N_7156);
or U7392 (N_7392,N_7190,N_7050);
xnor U7393 (N_7393,N_7117,N_7127);
xor U7394 (N_7394,N_7119,N_7050);
or U7395 (N_7395,N_7086,N_7109);
and U7396 (N_7396,N_7030,N_7054);
nor U7397 (N_7397,N_7077,N_7083);
nand U7398 (N_7398,N_7043,N_7046);
or U7399 (N_7399,N_7015,N_7157);
nor U7400 (N_7400,N_7287,N_7281);
and U7401 (N_7401,N_7343,N_7324);
or U7402 (N_7402,N_7375,N_7360);
or U7403 (N_7403,N_7294,N_7354);
nand U7404 (N_7404,N_7239,N_7278);
nand U7405 (N_7405,N_7233,N_7369);
nor U7406 (N_7406,N_7336,N_7262);
or U7407 (N_7407,N_7248,N_7225);
or U7408 (N_7408,N_7203,N_7328);
and U7409 (N_7409,N_7379,N_7384);
and U7410 (N_7410,N_7265,N_7200);
nand U7411 (N_7411,N_7297,N_7329);
nand U7412 (N_7412,N_7269,N_7220);
xnor U7413 (N_7413,N_7394,N_7256);
xnor U7414 (N_7414,N_7386,N_7353);
nor U7415 (N_7415,N_7208,N_7267);
and U7416 (N_7416,N_7361,N_7259);
nor U7417 (N_7417,N_7289,N_7243);
nor U7418 (N_7418,N_7363,N_7230);
and U7419 (N_7419,N_7214,N_7245);
nor U7420 (N_7420,N_7215,N_7309);
or U7421 (N_7421,N_7295,N_7226);
or U7422 (N_7422,N_7204,N_7284);
or U7423 (N_7423,N_7249,N_7366);
nand U7424 (N_7424,N_7356,N_7345);
nand U7425 (N_7425,N_7320,N_7342);
nand U7426 (N_7426,N_7219,N_7382);
or U7427 (N_7427,N_7319,N_7338);
and U7428 (N_7428,N_7307,N_7283);
nor U7429 (N_7429,N_7397,N_7252);
and U7430 (N_7430,N_7352,N_7251);
nand U7431 (N_7431,N_7270,N_7376);
nor U7432 (N_7432,N_7247,N_7257);
and U7433 (N_7433,N_7272,N_7276);
and U7434 (N_7434,N_7395,N_7367);
nand U7435 (N_7435,N_7346,N_7237);
nor U7436 (N_7436,N_7303,N_7349);
or U7437 (N_7437,N_7286,N_7339);
nand U7438 (N_7438,N_7337,N_7313);
nor U7439 (N_7439,N_7322,N_7254);
and U7440 (N_7440,N_7365,N_7305);
nor U7441 (N_7441,N_7327,N_7378);
xnor U7442 (N_7442,N_7323,N_7300);
nor U7443 (N_7443,N_7236,N_7334);
and U7444 (N_7444,N_7315,N_7302);
or U7445 (N_7445,N_7383,N_7316);
xor U7446 (N_7446,N_7250,N_7273);
nand U7447 (N_7447,N_7240,N_7209);
and U7448 (N_7448,N_7341,N_7304);
or U7449 (N_7449,N_7351,N_7340);
nand U7450 (N_7450,N_7282,N_7314);
nand U7451 (N_7451,N_7235,N_7372);
and U7452 (N_7452,N_7234,N_7211);
or U7453 (N_7453,N_7393,N_7333);
or U7454 (N_7454,N_7399,N_7350);
or U7455 (N_7455,N_7373,N_7202);
nor U7456 (N_7456,N_7244,N_7210);
nand U7457 (N_7457,N_7310,N_7398);
nand U7458 (N_7458,N_7325,N_7261);
nor U7459 (N_7459,N_7370,N_7321);
and U7460 (N_7460,N_7222,N_7255);
and U7461 (N_7461,N_7238,N_7385);
or U7462 (N_7462,N_7392,N_7308);
nand U7463 (N_7463,N_7277,N_7330);
nor U7464 (N_7464,N_7292,N_7205);
or U7465 (N_7465,N_7280,N_7227);
xor U7466 (N_7466,N_7298,N_7357);
xor U7467 (N_7467,N_7306,N_7231);
nor U7468 (N_7468,N_7279,N_7263);
nand U7469 (N_7469,N_7387,N_7266);
nor U7470 (N_7470,N_7258,N_7260);
or U7471 (N_7471,N_7213,N_7396);
nor U7472 (N_7472,N_7331,N_7296);
and U7473 (N_7473,N_7317,N_7347);
nand U7474 (N_7474,N_7207,N_7246);
and U7475 (N_7475,N_7206,N_7374);
and U7476 (N_7476,N_7264,N_7301);
xor U7477 (N_7477,N_7344,N_7218);
and U7478 (N_7478,N_7275,N_7326);
xnor U7479 (N_7479,N_7253,N_7293);
xnor U7480 (N_7480,N_7364,N_7299);
and U7481 (N_7481,N_7242,N_7223);
nor U7482 (N_7482,N_7201,N_7368);
nor U7483 (N_7483,N_7362,N_7271);
nor U7484 (N_7484,N_7377,N_7358);
xor U7485 (N_7485,N_7216,N_7380);
or U7486 (N_7486,N_7285,N_7348);
nor U7487 (N_7487,N_7389,N_7228);
or U7488 (N_7488,N_7390,N_7217);
and U7489 (N_7489,N_7388,N_7381);
or U7490 (N_7490,N_7288,N_7312);
nand U7491 (N_7491,N_7291,N_7332);
nand U7492 (N_7492,N_7274,N_7268);
nor U7493 (N_7493,N_7318,N_7241);
nor U7494 (N_7494,N_7355,N_7224);
nor U7495 (N_7495,N_7359,N_7371);
and U7496 (N_7496,N_7232,N_7391);
nor U7497 (N_7497,N_7221,N_7290);
and U7498 (N_7498,N_7212,N_7335);
nand U7499 (N_7499,N_7311,N_7229);
and U7500 (N_7500,N_7301,N_7246);
or U7501 (N_7501,N_7299,N_7241);
or U7502 (N_7502,N_7392,N_7330);
nand U7503 (N_7503,N_7379,N_7215);
xnor U7504 (N_7504,N_7243,N_7248);
or U7505 (N_7505,N_7282,N_7288);
nand U7506 (N_7506,N_7353,N_7313);
nand U7507 (N_7507,N_7229,N_7374);
xor U7508 (N_7508,N_7233,N_7271);
xnor U7509 (N_7509,N_7291,N_7200);
nor U7510 (N_7510,N_7306,N_7364);
and U7511 (N_7511,N_7299,N_7217);
nand U7512 (N_7512,N_7362,N_7299);
nor U7513 (N_7513,N_7223,N_7364);
nor U7514 (N_7514,N_7227,N_7283);
nor U7515 (N_7515,N_7345,N_7341);
and U7516 (N_7516,N_7296,N_7227);
or U7517 (N_7517,N_7273,N_7301);
nor U7518 (N_7518,N_7284,N_7317);
and U7519 (N_7519,N_7272,N_7279);
nand U7520 (N_7520,N_7261,N_7364);
nand U7521 (N_7521,N_7214,N_7269);
and U7522 (N_7522,N_7354,N_7395);
nor U7523 (N_7523,N_7363,N_7357);
and U7524 (N_7524,N_7375,N_7323);
nor U7525 (N_7525,N_7330,N_7349);
or U7526 (N_7526,N_7323,N_7330);
or U7527 (N_7527,N_7373,N_7384);
and U7528 (N_7528,N_7351,N_7238);
or U7529 (N_7529,N_7366,N_7292);
xnor U7530 (N_7530,N_7383,N_7278);
xor U7531 (N_7531,N_7368,N_7375);
nor U7532 (N_7532,N_7222,N_7330);
xor U7533 (N_7533,N_7228,N_7363);
nor U7534 (N_7534,N_7274,N_7350);
nand U7535 (N_7535,N_7269,N_7325);
nand U7536 (N_7536,N_7292,N_7270);
xor U7537 (N_7537,N_7306,N_7255);
nor U7538 (N_7538,N_7275,N_7277);
and U7539 (N_7539,N_7218,N_7293);
or U7540 (N_7540,N_7387,N_7242);
or U7541 (N_7541,N_7327,N_7330);
or U7542 (N_7542,N_7224,N_7385);
nand U7543 (N_7543,N_7212,N_7373);
or U7544 (N_7544,N_7373,N_7342);
nor U7545 (N_7545,N_7201,N_7271);
or U7546 (N_7546,N_7331,N_7214);
nand U7547 (N_7547,N_7397,N_7217);
xnor U7548 (N_7548,N_7254,N_7334);
and U7549 (N_7549,N_7230,N_7369);
nand U7550 (N_7550,N_7386,N_7240);
xor U7551 (N_7551,N_7320,N_7344);
and U7552 (N_7552,N_7328,N_7314);
nand U7553 (N_7553,N_7261,N_7358);
or U7554 (N_7554,N_7204,N_7333);
and U7555 (N_7555,N_7252,N_7253);
nor U7556 (N_7556,N_7320,N_7387);
and U7557 (N_7557,N_7309,N_7210);
nand U7558 (N_7558,N_7323,N_7318);
nor U7559 (N_7559,N_7364,N_7355);
and U7560 (N_7560,N_7370,N_7264);
or U7561 (N_7561,N_7287,N_7223);
xor U7562 (N_7562,N_7254,N_7239);
nand U7563 (N_7563,N_7224,N_7344);
and U7564 (N_7564,N_7326,N_7354);
nand U7565 (N_7565,N_7233,N_7211);
nor U7566 (N_7566,N_7343,N_7330);
and U7567 (N_7567,N_7229,N_7387);
nand U7568 (N_7568,N_7278,N_7326);
and U7569 (N_7569,N_7236,N_7371);
nand U7570 (N_7570,N_7207,N_7253);
nand U7571 (N_7571,N_7235,N_7385);
xor U7572 (N_7572,N_7379,N_7257);
and U7573 (N_7573,N_7282,N_7273);
or U7574 (N_7574,N_7351,N_7221);
nand U7575 (N_7575,N_7308,N_7272);
nand U7576 (N_7576,N_7241,N_7388);
nand U7577 (N_7577,N_7215,N_7262);
or U7578 (N_7578,N_7293,N_7251);
or U7579 (N_7579,N_7285,N_7344);
nand U7580 (N_7580,N_7292,N_7254);
nand U7581 (N_7581,N_7218,N_7372);
and U7582 (N_7582,N_7203,N_7304);
nand U7583 (N_7583,N_7377,N_7343);
or U7584 (N_7584,N_7279,N_7221);
xnor U7585 (N_7585,N_7317,N_7283);
nor U7586 (N_7586,N_7260,N_7230);
nand U7587 (N_7587,N_7213,N_7223);
and U7588 (N_7588,N_7317,N_7311);
nand U7589 (N_7589,N_7385,N_7296);
and U7590 (N_7590,N_7247,N_7327);
or U7591 (N_7591,N_7370,N_7278);
or U7592 (N_7592,N_7305,N_7309);
and U7593 (N_7593,N_7307,N_7217);
nand U7594 (N_7594,N_7232,N_7352);
xor U7595 (N_7595,N_7344,N_7383);
or U7596 (N_7596,N_7242,N_7335);
or U7597 (N_7597,N_7341,N_7205);
nand U7598 (N_7598,N_7327,N_7394);
nor U7599 (N_7599,N_7373,N_7375);
nand U7600 (N_7600,N_7534,N_7527);
or U7601 (N_7601,N_7519,N_7428);
or U7602 (N_7602,N_7543,N_7593);
and U7603 (N_7603,N_7469,N_7541);
nand U7604 (N_7604,N_7410,N_7438);
nor U7605 (N_7605,N_7451,N_7506);
nor U7606 (N_7606,N_7565,N_7520);
nand U7607 (N_7607,N_7457,N_7580);
and U7608 (N_7608,N_7406,N_7424);
and U7609 (N_7609,N_7422,N_7532);
nand U7610 (N_7610,N_7596,N_7552);
or U7611 (N_7611,N_7550,N_7515);
and U7612 (N_7612,N_7456,N_7569);
nor U7613 (N_7613,N_7579,N_7407);
nor U7614 (N_7614,N_7590,N_7510);
xor U7615 (N_7615,N_7467,N_7546);
and U7616 (N_7616,N_7439,N_7553);
and U7617 (N_7617,N_7591,N_7431);
nand U7618 (N_7618,N_7521,N_7533);
and U7619 (N_7619,N_7577,N_7417);
nand U7620 (N_7620,N_7524,N_7516);
nand U7621 (N_7621,N_7465,N_7414);
and U7622 (N_7622,N_7459,N_7528);
and U7623 (N_7623,N_7471,N_7595);
or U7624 (N_7624,N_7436,N_7567);
and U7625 (N_7625,N_7599,N_7586);
xnor U7626 (N_7626,N_7560,N_7500);
nand U7627 (N_7627,N_7462,N_7453);
or U7628 (N_7628,N_7574,N_7537);
or U7629 (N_7629,N_7425,N_7556);
nor U7630 (N_7630,N_7484,N_7478);
xor U7631 (N_7631,N_7493,N_7589);
and U7632 (N_7632,N_7508,N_7404);
nand U7633 (N_7633,N_7423,N_7522);
nand U7634 (N_7634,N_7566,N_7432);
and U7635 (N_7635,N_7557,N_7400);
nor U7636 (N_7636,N_7443,N_7473);
or U7637 (N_7637,N_7507,N_7578);
or U7638 (N_7638,N_7433,N_7446);
nand U7639 (N_7639,N_7549,N_7488);
xnor U7640 (N_7640,N_7409,N_7497);
nand U7641 (N_7641,N_7504,N_7444);
xnor U7642 (N_7642,N_7536,N_7517);
or U7643 (N_7643,N_7430,N_7491);
nor U7644 (N_7644,N_7477,N_7450);
nor U7645 (N_7645,N_7480,N_7494);
and U7646 (N_7646,N_7470,N_7492);
and U7647 (N_7647,N_7572,N_7585);
nand U7648 (N_7648,N_7452,N_7518);
or U7649 (N_7649,N_7476,N_7481);
nor U7650 (N_7650,N_7511,N_7525);
nor U7651 (N_7651,N_7495,N_7402);
or U7652 (N_7652,N_7499,N_7435);
xnor U7653 (N_7653,N_7485,N_7412);
or U7654 (N_7654,N_7460,N_7454);
xnor U7655 (N_7655,N_7496,N_7475);
nor U7656 (N_7656,N_7598,N_7555);
and U7657 (N_7657,N_7461,N_7415);
nand U7658 (N_7658,N_7582,N_7539);
or U7659 (N_7659,N_7530,N_7570);
nor U7660 (N_7660,N_7526,N_7535);
and U7661 (N_7661,N_7583,N_7540);
or U7662 (N_7662,N_7408,N_7498);
and U7663 (N_7663,N_7573,N_7483);
and U7664 (N_7664,N_7420,N_7513);
or U7665 (N_7665,N_7437,N_7501);
nor U7666 (N_7666,N_7575,N_7581);
xor U7667 (N_7667,N_7474,N_7564);
nand U7668 (N_7668,N_7531,N_7448);
nor U7669 (N_7669,N_7486,N_7421);
nor U7670 (N_7670,N_7568,N_7403);
nand U7671 (N_7671,N_7449,N_7455);
and U7672 (N_7672,N_7487,N_7529);
xor U7673 (N_7673,N_7561,N_7463);
nor U7674 (N_7674,N_7547,N_7514);
or U7675 (N_7675,N_7418,N_7479);
and U7676 (N_7676,N_7490,N_7551);
and U7677 (N_7677,N_7405,N_7597);
nand U7678 (N_7678,N_7559,N_7512);
and U7679 (N_7679,N_7466,N_7538);
or U7680 (N_7680,N_7440,N_7468);
or U7681 (N_7681,N_7502,N_7509);
or U7682 (N_7682,N_7503,N_7558);
or U7683 (N_7683,N_7413,N_7472);
or U7684 (N_7684,N_7505,N_7401);
nor U7685 (N_7685,N_7542,N_7587);
nor U7686 (N_7686,N_7442,N_7426);
or U7687 (N_7687,N_7445,N_7458);
or U7688 (N_7688,N_7554,N_7544);
nor U7689 (N_7689,N_7482,N_7427);
and U7690 (N_7690,N_7464,N_7419);
or U7691 (N_7691,N_7416,N_7434);
nand U7692 (N_7692,N_7594,N_7429);
or U7693 (N_7693,N_7523,N_7545);
or U7694 (N_7694,N_7588,N_7441);
nor U7695 (N_7695,N_7592,N_7571);
xor U7696 (N_7696,N_7548,N_7411);
nand U7697 (N_7697,N_7489,N_7447);
or U7698 (N_7698,N_7576,N_7584);
nand U7699 (N_7699,N_7562,N_7563);
nor U7700 (N_7700,N_7436,N_7540);
and U7701 (N_7701,N_7521,N_7587);
nor U7702 (N_7702,N_7483,N_7464);
nor U7703 (N_7703,N_7452,N_7483);
nor U7704 (N_7704,N_7458,N_7532);
nand U7705 (N_7705,N_7403,N_7563);
and U7706 (N_7706,N_7448,N_7433);
or U7707 (N_7707,N_7590,N_7598);
nand U7708 (N_7708,N_7464,N_7478);
and U7709 (N_7709,N_7491,N_7435);
nor U7710 (N_7710,N_7573,N_7452);
nand U7711 (N_7711,N_7441,N_7528);
nor U7712 (N_7712,N_7599,N_7423);
nand U7713 (N_7713,N_7409,N_7531);
or U7714 (N_7714,N_7591,N_7448);
or U7715 (N_7715,N_7465,N_7494);
or U7716 (N_7716,N_7529,N_7480);
nand U7717 (N_7717,N_7578,N_7531);
and U7718 (N_7718,N_7544,N_7528);
nand U7719 (N_7719,N_7452,N_7555);
nor U7720 (N_7720,N_7579,N_7545);
or U7721 (N_7721,N_7420,N_7475);
xnor U7722 (N_7722,N_7442,N_7579);
nand U7723 (N_7723,N_7530,N_7424);
and U7724 (N_7724,N_7544,N_7580);
xnor U7725 (N_7725,N_7482,N_7580);
and U7726 (N_7726,N_7520,N_7517);
nand U7727 (N_7727,N_7564,N_7549);
nor U7728 (N_7728,N_7524,N_7473);
nor U7729 (N_7729,N_7580,N_7536);
nor U7730 (N_7730,N_7520,N_7494);
or U7731 (N_7731,N_7426,N_7479);
nor U7732 (N_7732,N_7557,N_7405);
or U7733 (N_7733,N_7449,N_7568);
nor U7734 (N_7734,N_7419,N_7410);
and U7735 (N_7735,N_7421,N_7465);
or U7736 (N_7736,N_7516,N_7598);
or U7737 (N_7737,N_7535,N_7573);
nand U7738 (N_7738,N_7561,N_7472);
nor U7739 (N_7739,N_7492,N_7444);
nand U7740 (N_7740,N_7411,N_7455);
and U7741 (N_7741,N_7522,N_7488);
nand U7742 (N_7742,N_7416,N_7537);
or U7743 (N_7743,N_7573,N_7595);
and U7744 (N_7744,N_7460,N_7474);
nor U7745 (N_7745,N_7483,N_7503);
nor U7746 (N_7746,N_7491,N_7470);
nand U7747 (N_7747,N_7520,N_7480);
xnor U7748 (N_7748,N_7498,N_7454);
and U7749 (N_7749,N_7430,N_7555);
nand U7750 (N_7750,N_7545,N_7531);
nor U7751 (N_7751,N_7580,N_7407);
xnor U7752 (N_7752,N_7571,N_7420);
nand U7753 (N_7753,N_7507,N_7469);
nor U7754 (N_7754,N_7404,N_7504);
xnor U7755 (N_7755,N_7401,N_7455);
or U7756 (N_7756,N_7401,N_7468);
nor U7757 (N_7757,N_7523,N_7509);
nor U7758 (N_7758,N_7476,N_7440);
xor U7759 (N_7759,N_7522,N_7476);
or U7760 (N_7760,N_7512,N_7514);
nor U7761 (N_7761,N_7521,N_7565);
nand U7762 (N_7762,N_7507,N_7459);
nand U7763 (N_7763,N_7506,N_7414);
or U7764 (N_7764,N_7447,N_7461);
or U7765 (N_7765,N_7452,N_7429);
nor U7766 (N_7766,N_7518,N_7469);
nand U7767 (N_7767,N_7540,N_7570);
nand U7768 (N_7768,N_7445,N_7410);
nand U7769 (N_7769,N_7460,N_7587);
and U7770 (N_7770,N_7421,N_7417);
xnor U7771 (N_7771,N_7516,N_7562);
and U7772 (N_7772,N_7539,N_7552);
nand U7773 (N_7773,N_7529,N_7430);
nor U7774 (N_7774,N_7513,N_7480);
nor U7775 (N_7775,N_7465,N_7502);
or U7776 (N_7776,N_7476,N_7431);
nand U7777 (N_7777,N_7577,N_7468);
nor U7778 (N_7778,N_7443,N_7521);
xnor U7779 (N_7779,N_7548,N_7429);
and U7780 (N_7780,N_7409,N_7567);
xnor U7781 (N_7781,N_7438,N_7564);
and U7782 (N_7782,N_7560,N_7404);
nor U7783 (N_7783,N_7486,N_7449);
nor U7784 (N_7784,N_7473,N_7432);
nor U7785 (N_7785,N_7546,N_7559);
nor U7786 (N_7786,N_7577,N_7551);
nand U7787 (N_7787,N_7531,N_7573);
and U7788 (N_7788,N_7502,N_7478);
and U7789 (N_7789,N_7599,N_7416);
nand U7790 (N_7790,N_7541,N_7502);
or U7791 (N_7791,N_7408,N_7421);
nand U7792 (N_7792,N_7564,N_7425);
and U7793 (N_7793,N_7478,N_7476);
and U7794 (N_7794,N_7552,N_7554);
nand U7795 (N_7795,N_7422,N_7550);
nor U7796 (N_7796,N_7518,N_7434);
nor U7797 (N_7797,N_7545,N_7421);
or U7798 (N_7798,N_7479,N_7502);
nand U7799 (N_7799,N_7467,N_7429);
nor U7800 (N_7800,N_7732,N_7662);
nand U7801 (N_7801,N_7785,N_7646);
and U7802 (N_7802,N_7682,N_7759);
xor U7803 (N_7803,N_7642,N_7729);
and U7804 (N_7804,N_7799,N_7680);
or U7805 (N_7805,N_7654,N_7723);
or U7806 (N_7806,N_7612,N_7798);
nor U7807 (N_7807,N_7624,N_7692);
nand U7808 (N_7808,N_7766,N_7748);
or U7809 (N_7809,N_7647,N_7629);
nor U7810 (N_7810,N_7669,N_7733);
or U7811 (N_7811,N_7797,N_7606);
or U7812 (N_7812,N_7790,N_7701);
nor U7813 (N_7813,N_7764,N_7730);
xnor U7814 (N_7814,N_7725,N_7779);
nand U7815 (N_7815,N_7602,N_7696);
and U7816 (N_7816,N_7713,N_7721);
nor U7817 (N_7817,N_7716,N_7683);
nor U7818 (N_7818,N_7690,N_7728);
nor U7819 (N_7819,N_7621,N_7638);
xnor U7820 (N_7820,N_7755,N_7739);
or U7821 (N_7821,N_7639,N_7743);
nand U7822 (N_7822,N_7636,N_7780);
nor U7823 (N_7823,N_7640,N_7633);
xor U7824 (N_7824,N_7758,N_7783);
nor U7825 (N_7825,N_7668,N_7695);
xor U7826 (N_7826,N_7742,N_7684);
nand U7827 (N_7827,N_7671,N_7751);
and U7828 (N_7828,N_7617,N_7698);
xor U7829 (N_7829,N_7618,N_7605);
nand U7830 (N_7830,N_7632,N_7762);
nor U7831 (N_7831,N_7767,N_7637);
or U7832 (N_7832,N_7664,N_7649);
nor U7833 (N_7833,N_7774,N_7709);
and U7834 (N_7834,N_7643,N_7674);
nand U7835 (N_7835,N_7699,N_7641);
or U7836 (N_7836,N_7737,N_7675);
nor U7837 (N_7837,N_7765,N_7736);
nor U7838 (N_7838,N_7651,N_7719);
nand U7839 (N_7839,N_7622,N_7724);
or U7840 (N_7840,N_7689,N_7650);
nand U7841 (N_7841,N_7672,N_7685);
nor U7842 (N_7842,N_7776,N_7753);
and U7843 (N_7843,N_7673,N_7628);
nor U7844 (N_7844,N_7760,N_7784);
nand U7845 (N_7845,N_7796,N_7772);
xor U7846 (N_7846,N_7666,N_7626);
or U7847 (N_7847,N_7773,N_7793);
nand U7848 (N_7848,N_7611,N_7686);
nand U7849 (N_7849,N_7603,N_7738);
nand U7850 (N_7850,N_7634,N_7787);
or U7851 (N_7851,N_7704,N_7794);
xnor U7852 (N_7852,N_7714,N_7769);
or U7853 (N_7853,N_7744,N_7731);
or U7854 (N_7854,N_7763,N_7677);
and U7855 (N_7855,N_7754,N_7705);
or U7856 (N_7856,N_7613,N_7741);
and U7857 (N_7857,N_7726,N_7619);
nor U7858 (N_7858,N_7608,N_7777);
nor U7859 (N_7859,N_7691,N_7708);
nor U7860 (N_7860,N_7717,N_7778);
and U7861 (N_7861,N_7782,N_7610);
nand U7862 (N_7862,N_7715,N_7718);
nand U7863 (N_7863,N_7687,N_7630);
or U7864 (N_7864,N_7735,N_7609);
nor U7865 (N_7865,N_7614,N_7703);
and U7866 (N_7866,N_7625,N_7600);
xor U7867 (N_7867,N_7688,N_7655);
nor U7868 (N_7868,N_7694,N_7720);
nand U7869 (N_7869,N_7663,N_7702);
and U7870 (N_7870,N_7659,N_7706);
nand U7871 (N_7871,N_7757,N_7679);
nor U7872 (N_7872,N_7670,N_7652);
nand U7873 (N_7873,N_7771,N_7749);
nand U7874 (N_7874,N_7707,N_7745);
nor U7875 (N_7875,N_7786,N_7620);
nand U7876 (N_7876,N_7660,N_7700);
and U7877 (N_7877,N_7601,N_7756);
nor U7878 (N_7878,N_7775,N_7788);
and U7879 (N_7879,N_7747,N_7734);
nand U7880 (N_7880,N_7681,N_7722);
or U7881 (N_7881,N_7789,N_7665);
nor U7882 (N_7882,N_7727,N_7607);
nand U7883 (N_7883,N_7750,N_7746);
nand U7884 (N_7884,N_7791,N_7658);
and U7885 (N_7885,N_7792,N_7615);
and U7886 (N_7886,N_7678,N_7661);
or U7887 (N_7887,N_7768,N_7645);
nor U7888 (N_7888,N_7676,N_7740);
or U7889 (N_7889,N_7616,N_7761);
nor U7890 (N_7890,N_7648,N_7644);
and U7891 (N_7891,N_7631,N_7697);
nand U7892 (N_7892,N_7667,N_7623);
xor U7893 (N_7893,N_7693,N_7712);
and U7894 (N_7894,N_7604,N_7627);
and U7895 (N_7895,N_7635,N_7795);
or U7896 (N_7896,N_7752,N_7653);
or U7897 (N_7897,N_7710,N_7656);
nor U7898 (N_7898,N_7770,N_7657);
nand U7899 (N_7899,N_7711,N_7781);
and U7900 (N_7900,N_7688,N_7788);
and U7901 (N_7901,N_7763,N_7701);
or U7902 (N_7902,N_7733,N_7766);
nand U7903 (N_7903,N_7622,N_7735);
or U7904 (N_7904,N_7666,N_7682);
and U7905 (N_7905,N_7628,N_7602);
or U7906 (N_7906,N_7647,N_7639);
nand U7907 (N_7907,N_7731,N_7663);
or U7908 (N_7908,N_7600,N_7761);
nor U7909 (N_7909,N_7630,N_7663);
nand U7910 (N_7910,N_7725,N_7688);
and U7911 (N_7911,N_7653,N_7627);
xor U7912 (N_7912,N_7741,N_7605);
xnor U7913 (N_7913,N_7672,N_7690);
nor U7914 (N_7914,N_7755,N_7700);
nor U7915 (N_7915,N_7660,N_7707);
xor U7916 (N_7916,N_7764,N_7701);
and U7917 (N_7917,N_7792,N_7772);
nand U7918 (N_7918,N_7671,N_7663);
xor U7919 (N_7919,N_7624,N_7632);
and U7920 (N_7920,N_7675,N_7695);
or U7921 (N_7921,N_7689,N_7615);
or U7922 (N_7922,N_7625,N_7650);
and U7923 (N_7923,N_7704,N_7670);
and U7924 (N_7924,N_7668,N_7622);
xor U7925 (N_7925,N_7791,N_7742);
nor U7926 (N_7926,N_7614,N_7689);
or U7927 (N_7927,N_7698,N_7754);
nor U7928 (N_7928,N_7782,N_7706);
xor U7929 (N_7929,N_7671,N_7602);
nand U7930 (N_7930,N_7758,N_7680);
nor U7931 (N_7931,N_7794,N_7753);
nand U7932 (N_7932,N_7789,N_7643);
and U7933 (N_7933,N_7794,N_7636);
nor U7934 (N_7934,N_7748,N_7726);
and U7935 (N_7935,N_7666,N_7721);
nor U7936 (N_7936,N_7785,N_7762);
and U7937 (N_7937,N_7780,N_7695);
nor U7938 (N_7938,N_7707,N_7686);
or U7939 (N_7939,N_7755,N_7741);
and U7940 (N_7940,N_7700,N_7704);
nand U7941 (N_7941,N_7621,N_7643);
nand U7942 (N_7942,N_7712,N_7751);
nand U7943 (N_7943,N_7735,N_7645);
nor U7944 (N_7944,N_7667,N_7760);
and U7945 (N_7945,N_7667,N_7712);
nand U7946 (N_7946,N_7649,N_7655);
and U7947 (N_7947,N_7736,N_7685);
nor U7948 (N_7948,N_7773,N_7684);
or U7949 (N_7949,N_7724,N_7601);
or U7950 (N_7950,N_7735,N_7644);
and U7951 (N_7951,N_7709,N_7793);
xor U7952 (N_7952,N_7620,N_7658);
nand U7953 (N_7953,N_7704,N_7673);
or U7954 (N_7954,N_7710,N_7630);
nor U7955 (N_7955,N_7751,N_7740);
nand U7956 (N_7956,N_7641,N_7775);
and U7957 (N_7957,N_7731,N_7749);
nand U7958 (N_7958,N_7778,N_7690);
nor U7959 (N_7959,N_7603,N_7799);
nor U7960 (N_7960,N_7676,N_7748);
xnor U7961 (N_7961,N_7676,N_7712);
or U7962 (N_7962,N_7602,N_7611);
nor U7963 (N_7963,N_7787,N_7773);
and U7964 (N_7964,N_7784,N_7743);
and U7965 (N_7965,N_7709,N_7787);
nor U7966 (N_7966,N_7635,N_7604);
and U7967 (N_7967,N_7659,N_7679);
or U7968 (N_7968,N_7685,N_7693);
and U7969 (N_7969,N_7672,N_7744);
xnor U7970 (N_7970,N_7685,N_7715);
nor U7971 (N_7971,N_7769,N_7780);
or U7972 (N_7972,N_7767,N_7759);
and U7973 (N_7973,N_7625,N_7762);
nand U7974 (N_7974,N_7743,N_7654);
and U7975 (N_7975,N_7639,N_7659);
and U7976 (N_7976,N_7798,N_7755);
and U7977 (N_7977,N_7600,N_7708);
nand U7978 (N_7978,N_7629,N_7678);
and U7979 (N_7979,N_7639,N_7687);
nor U7980 (N_7980,N_7610,N_7600);
nand U7981 (N_7981,N_7708,N_7627);
nor U7982 (N_7982,N_7770,N_7677);
nand U7983 (N_7983,N_7747,N_7679);
or U7984 (N_7984,N_7625,N_7787);
xor U7985 (N_7985,N_7721,N_7744);
or U7986 (N_7986,N_7738,N_7790);
nand U7987 (N_7987,N_7719,N_7799);
and U7988 (N_7988,N_7720,N_7716);
nor U7989 (N_7989,N_7743,N_7791);
or U7990 (N_7990,N_7724,N_7767);
nor U7991 (N_7991,N_7607,N_7786);
and U7992 (N_7992,N_7604,N_7774);
or U7993 (N_7993,N_7643,N_7642);
or U7994 (N_7994,N_7660,N_7778);
and U7995 (N_7995,N_7639,N_7790);
or U7996 (N_7996,N_7643,N_7703);
xnor U7997 (N_7997,N_7727,N_7657);
nor U7998 (N_7998,N_7728,N_7631);
nand U7999 (N_7999,N_7621,N_7603);
or U8000 (N_8000,N_7803,N_7860);
or U8001 (N_8001,N_7918,N_7958);
or U8002 (N_8002,N_7930,N_7966);
nor U8003 (N_8003,N_7983,N_7962);
nand U8004 (N_8004,N_7824,N_7915);
nand U8005 (N_8005,N_7831,N_7972);
nor U8006 (N_8006,N_7991,N_7899);
and U8007 (N_8007,N_7920,N_7973);
nor U8008 (N_8008,N_7861,N_7961);
and U8009 (N_8009,N_7892,N_7932);
or U8010 (N_8010,N_7891,N_7828);
nor U8011 (N_8011,N_7989,N_7801);
and U8012 (N_8012,N_7808,N_7936);
nand U8013 (N_8013,N_7894,N_7996);
nand U8014 (N_8014,N_7922,N_7858);
or U8015 (N_8015,N_7848,N_7825);
or U8016 (N_8016,N_7965,N_7970);
nand U8017 (N_8017,N_7883,N_7866);
xnor U8018 (N_8018,N_7947,N_7907);
or U8019 (N_8019,N_7869,N_7941);
and U8020 (N_8020,N_7968,N_7971);
xnor U8021 (N_8021,N_7893,N_7827);
nand U8022 (N_8022,N_7806,N_7921);
or U8023 (N_8023,N_7999,N_7951);
nor U8024 (N_8024,N_7993,N_7826);
nor U8025 (N_8025,N_7815,N_7872);
nand U8026 (N_8026,N_7810,N_7800);
or U8027 (N_8027,N_7953,N_7917);
nor U8028 (N_8028,N_7855,N_7854);
nor U8029 (N_8029,N_7863,N_7885);
xnor U8030 (N_8030,N_7986,N_7844);
or U8031 (N_8031,N_7955,N_7868);
or U8032 (N_8032,N_7846,N_7839);
or U8033 (N_8033,N_7814,N_7981);
nor U8034 (N_8034,N_7865,N_7823);
and U8035 (N_8035,N_7985,N_7913);
nor U8036 (N_8036,N_7939,N_7964);
nand U8037 (N_8037,N_7959,N_7910);
and U8038 (N_8038,N_7895,N_7940);
nor U8039 (N_8039,N_7929,N_7925);
nor U8040 (N_8040,N_7919,N_7805);
and U8041 (N_8041,N_7926,N_7998);
or U8042 (N_8042,N_7813,N_7841);
nor U8043 (N_8043,N_7987,N_7931);
nor U8044 (N_8044,N_7845,N_7909);
nor U8045 (N_8045,N_7852,N_7994);
and U8046 (N_8046,N_7820,N_7954);
or U8047 (N_8047,N_7832,N_7904);
nand U8048 (N_8048,N_7949,N_7992);
nor U8049 (N_8049,N_7889,N_7906);
xor U8050 (N_8050,N_7916,N_7873);
xor U8051 (N_8051,N_7963,N_7842);
and U8052 (N_8052,N_7816,N_7829);
nand U8053 (N_8053,N_7967,N_7881);
or U8054 (N_8054,N_7830,N_7807);
or U8055 (N_8055,N_7818,N_7902);
or U8056 (N_8056,N_7938,N_7838);
xnor U8057 (N_8057,N_7979,N_7923);
nand U8058 (N_8058,N_7911,N_7851);
or U8059 (N_8059,N_7875,N_7990);
nor U8060 (N_8060,N_7853,N_7952);
nor U8061 (N_8061,N_7975,N_7819);
nor U8062 (N_8062,N_7944,N_7984);
nand U8063 (N_8063,N_7859,N_7980);
or U8064 (N_8064,N_7876,N_7802);
xor U8065 (N_8065,N_7847,N_7978);
xor U8066 (N_8066,N_7943,N_7884);
nor U8067 (N_8067,N_7879,N_7809);
xnor U8068 (N_8068,N_7969,N_7878);
nand U8069 (N_8069,N_7977,N_7864);
nand U8070 (N_8070,N_7942,N_7812);
nand U8071 (N_8071,N_7982,N_7882);
nand U8072 (N_8072,N_7886,N_7946);
and U8073 (N_8073,N_7880,N_7837);
and U8074 (N_8074,N_7817,N_7871);
or U8075 (N_8075,N_7905,N_7950);
and U8076 (N_8076,N_7935,N_7997);
nand U8077 (N_8077,N_7908,N_7927);
and U8078 (N_8078,N_7811,N_7857);
and U8079 (N_8079,N_7901,N_7840);
and U8080 (N_8080,N_7928,N_7960);
and U8081 (N_8081,N_7937,N_7896);
or U8082 (N_8082,N_7934,N_7897);
nand U8083 (N_8083,N_7821,N_7924);
nor U8084 (N_8084,N_7862,N_7870);
nor U8085 (N_8085,N_7903,N_7912);
and U8086 (N_8086,N_7835,N_7945);
nor U8087 (N_8087,N_7898,N_7874);
nor U8088 (N_8088,N_7914,N_7957);
nand U8089 (N_8089,N_7995,N_7804);
nand U8090 (N_8090,N_7834,N_7843);
nor U8091 (N_8091,N_7948,N_7833);
nor U8092 (N_8092,N_7849,N_7888);
or U8093 (N_8093,N_7890,N_7956);
nand U8094 (N_8094,N_7887,N_7974);
or U8095 (N_8095,N_7988,N_7900);
nor U8096 (N_8096,N_7976,N_7867);
or U8097 (N_8097,N_7856,N_7836);
or U8098 (N_8098,N_7933,N_7850);
and U8099 (N_8099,N_7877,N_7822);
nand U8100 (N_8100,N_7924,N_7889);
and U8101 (N_8101,N_7923,N_7814);
nand U8102 (N_8102,N_7942,N_7921);
or U8103 (N_8103,N_7811,N_7882);
xor U8104 (N_8104,N_7983,N_7850);
and U8105 (N_8105,N_7809,N_7812);
xnor U8106 (N_8106,N_7838,N_7891);
or U8107 (N_8107,N_7998,N_7902);
xor U8108 (N_8108,N_7929,N_7899);
nor U8109 (N_8109,N_7841,N_7970);
and U8110 (N_8110,N_7802,N_7973);
nor U8111 (N_8111,N_7821,N_7813);
nor U8112 (N_8112,N_7841,N_7932);
nor U8113 (N_8113,N_7985,N_7842);
and U8114 (N_8114,N_7827,N_7836);
nand U8115 (N_8115,N_7835,N_7954);
nor U8116 (N_8116,N_7975,N_7980);
nor U8117 (N_8117,N_7808,N_7939);
nand U8118 (N_8118,N_7841,N_7900);
nor U8119 (N_8119,N_7921,N_7869);
xor U8120 (N_8120,N_7885,N_7821);
and U8121 (N_8121,N_7848,N_7840);
xor U8122 (N_8122,N_7931,N_7965);
and U8123 (N_8123,N_7804,N_7854);
and U8124 (N_8124,N_7902,N_7882);
nand U8125 (N_8125,N_7817,N_7933);
or U8126 (N_8126,N_7917,N_7825);
xnor U8127 (N_8127,N_7859,N_7944);
and U8128 (N_8128,N_7940,N_7886);
and U8129 (N_8129,N_7887,N_7855);
nor U8130 (N_8130,N_7986,N_7885);
xor U8131 (N_8131,N_7971,N_7841);
nor U8132 (N_8132,N_7939,N_7942);
nand U8133 (N_8133,N_7936,N_7818);
or U8134 (N_8134,N_7806,N_7871);
xnor U8135 (N_8135,N_7816,N_7805);
or U8136 (N_8136,N_7886,N_7845);
nand U8137 (N_8137,N_7975,N_7835);
or U8138 (N_8138,N_7836,N_7868);
or U8139 (N_8139,N_7912,N_7822);
xor U8140 (N_8140,N_7835,N_7904);
nor U8141 (N_8141,N_7910,N_7815);
nor U8142 (N_8142,N_7895,N_7849);
nor U8143 (N_8143,N_7899,N_7803);
or U8144 (N_8144,N_7824,N_7896);
nand U8145 (N_8145,N_7830,N_7999);
or U8146 (N_8146,N_7815,N_7941);
or U8147 (N_8147,N_7946,N_7970);
nand U8148 (N_8148,N_7874,N_7838);
or U8149 (N_8149,N_7938,N_7999);
and U8150 (N_8150,N_7973,N_7948);
nand U8151 (N_8151,N_7915,N_7913);
xnor U8152 (N_8152,N_7949,N_7838);
xnor U8153 (N_8153,N_7951,N_7967);
xnor U8154 (N_8154,N_7819,N_7910);
nor U8155 (N_8155,N_7812,N_7888);
nor U8156 (N_8156,N_7963,N_7816);
nor U8157 (N_8157,N_7890,N_7964);
nor U8158 (N_8158,N_7821,N_7996);
and U8159 (N_8159,N_7888,N_7948);
xor U8160 (N_8160,N_7971,N_7871);
nand U8161 (N_8161,N_7912,N_7876);
nand U8162 (N_8162,N_7958,N_7963);
nand U8163 (N_8163,N_7999,N_7973);
and U8164 (N_8164,N_7885,N_7890);
nor U8165 (N_8165,N_7825,N_7860);
nand U8166 (N_8166,N_7866,N_7845);
and U8167 (N_8167,N_7989,N_7828);
or U8168 (N_8168,N_7832,N_7930);
xnor U8169 (N_8169,N_7857,N_7821);
nand U8170 (N_8170,N_7949,N_7807);
xnor U8171 (N_8171,N_7830,N_7988);
or U8172 (N_8172,N_7857,N_7874);
xnor U8173 (N_8173,N_7922,N_7814);
and U8174 (N_8174,N_7886,N_7805);
nor U8175 (N_8175,N_7958,N_7923);
nand U8176 (N_8176,N_7834,N_7898);
nor U8177 (N_8177,N_7842,N_7991);
or U8178 (N_8178,N_7850,N_7932);
nand U8179 (N_8179,N_7927,N_7809);
nor U8180 (N_8180,N_7950,N_7955);
and U8181 (N_8181,N_7983,N_7912);
or U8182 (N_8182,N_7838,N_7863);
or U8183 (N_8183,N_7933,N_7953);
nand U8184 (N_8184,N_7874,N_7876);
nor U8185 (N_8185,N_7803,N_7850);
and U8186 (N_8186,N_7801,N_7905);
xnor U8187 (N_8187,N_7812,N_7902);
and U8188 (N_8188,N_7906,N_7831);
or U8189 (N_8189,N_7856,N_7805);
nand U8190 (N_8190,N_7898,N_7828);
or U8191 (N_8191,N_7878,N_7931);
nand U8192 (N_8192,N_7858,N_7903);
and U8193 (N_8193,N_7861,N_7929);
or U8194 (N_8194,N_7959,N_7899);
and U8195 (N_8195,N_7833,N_7848);
nor U8196 (N_8196,N_7966,N_7860);
or U8197 (N_8197,N_7916,N_7922);
nand U8198 (N_8198,N_7908,N_7916);
or U8199 (N_8199,N_7916,N_7904);
and U8200 (N_8200,N_8066,N_8120);
xor U8201 (N_8201,N_8019,N_8079);
or U8202 (N_8202,N_8115,N_8102);
nor U8203 (N_8203,N_8002,N_8058);
or U8204 (N_8204,N_8095,N_8062);
nand U8205 (N_8205,N_8064,N_8128);
nor U8206 (N_8206,N_8109,N_8007);
nand U8207 (N_8207,N_8088,N_8103);
nor U8208 (N_8208,N_8187,N_8146);
nand U8209 (N_8209,N_8046,N_8040);
nor U8210 (N_8210,N_8168,N_8092);
nand U8211 (N_8211,N_8196,N_8060);
or U8212 (N_8212,N_8094,N_8086);
nand U8213 (N_8213,N_8181,N_8003);
and U8214 (N_8214,N_8018,N_8188);
nand U8215 (N_8215,N_8084,N_8148);
and U8216 (N_8216,N_8175,N_8123);
or U8217 (N_8217,N_8156,N_8093);
nor U8218 (N_8218,N_8192,N_8020);
nor U8219 (N_8219,N_8035,N_8159);
or U8220 (N_8220,N_8143,N_8068);
nor U8221 (N_8221,N_8053,N_8169);
or U8222 (N_8222,N_8043,N_8185);
nand U8223 (N_8223,N_8042,N_8033);
nand U8224 (N_8224,N_8063,N_8098);
and U8225 (N_8225,N_8154,N_8107);
or U8226 (N_8226,N_8172,N_8073);
or U8227 (N_8227,N_8097,N_8199);
or U8228 (N_8228,N_8089,N_8129);
nand U8229 (N_8229,N_8160,N_8125);
nand U8230 (N_8230,N_8044,N_8183);
and U8231 (N_8231,N_8024,N_8069);
and U8232 (N_8232,N_8155,N_8171);
nor U8233 (N_8233,N_8141,N_8126);
and U8234 (N_8234,N_8030,N_8174);
xor U8235 (N_8235,N_8057,N_8051);
and U8236 (N_8236,N_8015,N_8076);
nand U8237 (N_8237,N_8165,N_8081);
and U8238 (N_8238,N_8118,N_8186);
xor U8239 (N_8239,N_8184,N_8179);
nand U8240 (N_8240,N_8005,N_8072);
nand U8241 (N_8241,N_8149,N_8108);
or U8242 (N_8242,N_8134,N_8119);
nor U8243 (N_8243,N_8009,N_8090);
nor U8244 (N_8244,N_8133,N_8099);
nor U8245 (N_8245,N_8194,N_8191);
and U8246 (N_8246,N_8082,N_8147);
and U8247 (N_8247,N_8180,N_8193);
nand U8248 (N_8248,N_8113,N_8167);
nand U8249 (N_8249,N_8130,N_8027);
nand U8250 (N_8250,N_8152,N_8121);
xor U8251 (N_8251,N_8173,N_8023);
nor U8252 (N_8252,N_8177,N_8056);
nor U8253 (N_8253,N_8132,N_8162);
and U8254 (N_8254,N_8111,N_8189);
nor U8255 (N_8255,N_8047,N_8163);
nor U8256 (N_8256,N_8085,N_8144);
nand U8257 (N_8257,N_8045,N_8112);
nand U8258 (N_8258,N_8190,N_8050);
and U8259 (N_8259,N_8140,N_8070);
nor U8260 (N_8260,N_8198,N_8074);
and U8261 (N_8261,N_8182,N_8105);
nor U8262 (N_8262,N_8061,N_8011);
or U8263 (N_8263,N_8054,N_8131);
or U8264 (N_8264,N_8135,N_8096);
nand U8265 (N_8265,N_8022,N_8151);
nand U8266 (N_8266,N_8158,N_8176);
xor U8267 (N_8267,N_8145,N_8136);
or U8268 (N_8268,N_8041,N_8104);
or U8269 (N_8269,N_8106,N_8036);
or U8270 (N_8270,N_8137,N_8116);
nand U8271 (N_8271,N_8055,N_8157);
nor U8272 (N_8272,N_8161,N_8100);
nand U8273 (N_8273,N_8150,N_8166);
nand U8274 (N_8274,N_8048,N_8122);
nand U8275 (N_8275,N_8078,N_8016);
or U8276 (N_8276,N_8037,N_8014);
nand U8277 (N_8277,N_8065,N_8049);
nor U8278 (N_8278,N_8142,N_8153);
and U8279 (N_8279,N_8091,N_8031);
nor U8280 (N_8280,N_8114,N_8170);
nor U8281 (N_8281,N_8026,N_8195);
or U8282 (N_8282,N_8197,N_8029);
or U8283 (N_8283,N_8110,N_8080);
and U8284 (N_8284,N_8028,N_8017);
nand U8285 (N_8285,N_8021,N_8001);
and U8286 (N_8286,N_8101,N_8010);
or U8287 (N_8287,N_8052,N_8083);
nor U8288 (N_8288,N_8127,N_8178);
xnor U8289 (N_8289,N_8067,N_8006);
nand U8290 (N_8290,N_8139,N_8039);
nor U8291 (N_8291,N_8004,N_8075);
nand U8292 (N_8292,N_8038,N_8000);
nand U8293 (N_8293,N_8071,N_8124);
or U8294 (N_8294,N_8164,N_8117);
nor U8295 (N_8295,N_8034,N_8012);
nand U8296 (N_8296,N_8008,N_8025);
xnor U8297 (N_8297,N_8087,N_8059);
xnor U8298 (N_8298,N_8077,N_8032);
nor U8299 (N_8299,N_8013,N_8138);
nor U8300 (N_8300,N_8031,N_8178);
or U8301 (N_8301,N_8076,N_8165);
nor U8302 (N_8302,N_8022,N_8100);
nand U8303 (N_8303,N_8040,N_8059);
xor U8304 (N_8304,N_8106,N_8013);
nor U8305 (N_8305,N_8045,N_8172);
nor U8306 (N_8306,N_8178,N_8098);
nor U8307 (N_8307,N_8104,N_8189);
nor U8308 (N_8308,N_8086,N_8115);
or U8309 (N_8309,N_8114,N_8132);
and U8310 (N_8310,N_8022,N_8016);
nor U8311 (N_8311,N_8189,N_8053);
xor U8312 (N_8312,N_8052,N_8137);
nand U8313 (N_8313,N_8050,N_8114);
and U8314 (N_8314,N_8112,N_8083);
and U8315 (N_8315,N_8084,N_8126);
and U8316 (N_8316,N_8144,N_8035);
nand U8317 (N_8317,N_8021,N_8107);
and U8318 (N_8318,N_8041,N_8029);
and U8319 (N_8319,N_8019,N_8169);
xnor U8320 (N_8320,N_8144,N_8124);
nor U8321 (N_8321,N_8148,N_8165);
and U8322 (N_8322,N_8136,N_8062);
nand U8323 (N_8323,N_8044,N_8145);
nor U8324 (N_8324,N_8009,N_8132);
and U8325 (N_8325,N_8093,N_8153);
nor U8326 (N_8326,N_8176,N_8135);
nor U8327 (N_8327,N_8006,N_8195);
xnor U8328 (N_8328,N_8028,N_8025);
nor U8329 (N_8329,N_8182,N_8126);
nand U8330 (N_8330,N_8128,N_8091);
or U8331 (N_8331,N_8179,N_8195);
or U8332 (N_8332,N_8127,N_8187);
nand U8333 (N_8333,N_8135,N_8001);
nand U8334 (N_8334,N_8114,N_8081);
nor U8335 (N_8335,N_8034,N_8188);
and U8336 (N_8336,N_8156,N_8016);
nor U8337 (N_8337,N_8062,N_8064);
nand U8338 (N_8338,N_8017,N_8107);
and U8339 (N_8339,N_8005,N_8167);
nor U8340 (N_8340,N_8089,N_8140);
and U8341 (N_8341,N_8141,N_8050);
nand U8342 (N_8342,N_8193,N_8189);
xor U8343 (N_8343,N_8135,N_8166);
nor U8344 (N_8344,N_8103,N_8017);
and U8345 (N_8345,N_8088,N_8102);
and U8346 (N_8346,N_8132,N_8090);
and U8347 (N_8347,N_8177,N_8033);
or U8348 (N_8348,N_8132,N_8036);
or U8349 (N_8349,N_8022,N_8002);
nand U8350 (N_8350,N_8118,N_8021);
nor U8351 (N_8351,N_8183,N_8022);
nor U8352 (N_8352,N_8032,N_8153);
nand U8353 (N_8353,N_8174,N_8191);
or U8354 (N_8354,N_8031,N_8056);
nand U8355 (N_8355,N_8001,N_8169);
nand U8356 (N_8356,N_8089,N_8039);
or U8357 (N_8357,N_8059,N_8037);
or U8358 (N_8358,N_8119,N_8160);
nand U8359 (N_8359,N_8085,N_8160);
or U8360 (N_8360,N_8038,N_8170);
or U8361 (N_8361,N_8125,N_8180);
or U8362 (N_8362,N_8019,N_8025);
or U8363 (N_8363,N_8138,N_8004);
nand U8364 (N_8364,N_8119,N_8065);
nand U8365 (N_8365,N_8105,N_8151);
or U8366 (N_8366,N_8035,N_8197);
nor U8367 (N_8367,N_8183,N_8043);
nor U8368 (N_8368,N_8110,N_8096);
or U8369 (N_8369,N_8137,N_8053);
and U8370 (N_8370,N_8024,N_8039);
nor U8371 (N_8371,N_8111,N_8043);
or U8372 (N_8372,N_8050,N_8194);
nor U8373 (N_8373,N_8122,N_8054);
nor U8374 (N_8374,N_8064,N_8179);
nor U8375 (N_8375,N_8159,N_8101);
nand U8376 (N_8376,N_8174,N_8156);
xnor U8377 (N_8377,N_8195,N_8084);
nor U8378 (N_8378,N_8036,N_8080);
nand U8379 (N_8379,N_8154,N_8185);
nor U8380 (N_8380,N_8015,N_8018);
nand U8381 (N_8381,N_8122,N_8068);
nand U8382 (N_8382,N_8035,N_8088);
or U8383 (N_8383,N_8047,N_8087);
nor U8384 (N_8384,N_8010,N_8128);
nor U8385 (N_8385,N_8106,N_8089);
nand U8386 (N_8386,N_8117,N_8170);
and U8387 (N_8387,N_8031,N_8042);
nand U8388 (N_8388,N_8092,N_8040);
nor U8389 (N_8389,N_8150,N_8098);
nand U8390 (N_8390,N_8033,N_8048);
or U8391 (N_8391,N_8156,N_8066);
and U8392 (N_8392,N_8127,N_8067);
nand U8393 (N_8393,N_8029,N_8116);
nand U8394 (N_8394,N_8199,N_8120);
nor U8395 (N_8395,N_8043,N_8163);
nand U8396 (N_8396,N_8197,N_8111);
nor U8397 (N_8397,N_8063,N_8041);
and U8398 (N_8398,N_8073,N_8114);
or U8399 (N_8399,N_8028,N_8152);
and U8400 (N_8400,N_8239,N_8316);
xor U8401 (N_8401,N_8203,N_8354);
nand U8402 (N_8402,N_8388,N_8228);
nand U8403 (N_8403,N_8301,N_8399);
nor U8404 (N_8404,N_8295,N_8314);
or U8405 (N_8405,N_8333,N_8241);
and U8406 (N_8406,N_8214,N_8355);
nor U8407 (N_8407,N_8327,N_8273);
nor U8408 (N_8408,N_8356,N_8221);
and U8409 (N_8409,N_8227,N_8230);
and U8410 (N_8410,N_8282,N_8300);
and U8411 (N_8411,N_8217,N_8215);
nor U8412 (N_8412,N_8260,N_8237);
or U8413 (N_8413,N_8313,N_8322);
and U8414 (N_8414,N_8271,N_8247);
nand U8415 (N_8415,N_8339,N_8398);
nand U8416 (N_8416,N_8392,N_8384);
or U8417 (N_8417,N_8320,N_8341);
and U8418 (N_8418,N_8397,N_8340);
nand U8419 (N_8419,N_8298,N_8249);
and U8420 (N_8420,N_8378,N_8382);
or U8421 (N_8421,N_8229,N_8274);
and U8422 (N_8422,N_8281,N_8268);
or U8423 (N_8423,N_8279,N_8343);
nor U8424 (N_8424,N_8346,N_8350);
or U8425 (N_8425,N_8272,N_8297);
nand U8426 (N_8426,N_8380,N_8304);
xor U8427 (N_8427,N_8293,N_8323);
or U8428 (N_8428,N_8370,N_8210);
nor U8429 (N_8429,N_8289,N_8294);
nor U8430 (N_8430,N_8387,N_8222);
and U8431 (N_8431,N_8201,N_8232);
nor U8432 (N_8432,N_8362,N_8235);
xor U8433 (N_8433,N_8280,N_8256);
nand U8434 (N_8434,N_8347,N_8288);
xnor U8435 (N_8435,N_8325,N_8269);
xor U8436 (N_8436,N_8376,N_8352);
and U8437 (N_8437,N_8357,N_8286);
nor U8438 (N_8438,N_8225,N_8359);
xor U8439 (N_8439,N_8213,N_8226);
or U8440 (N_8440,N_8396,N_8265);
and U8441 (N_8441,N_8264,N_8263);
xor U8442 (N_8442,N_8231,N_8332);
or U8443 (N_8443,N_8367,N_8312);
or U8444 (N_8444,N_8205,N_8363);
nand U8445 (N_8445,N_8338,N_8248);
or U8446 (N_8446,N_8218,N_8360);
nand U8447 (N_8447,N_8216,N_8324);
nand U8448 (N_8448,N_8345,N_8250);
nor U8449 (N_8449,N_8329,N_8285);
and U8450 (N_8450,N_8374,N_8266);
nand U8451 (N_8451,N_8318,N_8385);
and U8452 (N_8452,N_8317,N_8344);
or U8453 (N_8453,N_8233,N_8254);
and U8454 (N_8454,N_8200,N_8259);
or U8455 (N_8455,N_8326,N_8365);
and U8456 (N_8456,N_8244,N_8207);
nor U8457 (N_8457,N_8276,N_8358);
nand U8458 (N_8458,N_8212,N_8277);
or U8459 (N_8459,N_8373,N_8394);
nor U8460 (N_8460,N_8262,N_8349);
xor U8461 (N_8461,N_8284,N_8219);
xor U8462 (N_8462,N_8389,N_8278);
xor U8463 (N_8463,N_8368,N_8283);
or U8464 (N_8464,N_8246,N_8255);
nor U8465 (N_8465,N_8240,N_8224);
and U8466 (N_8466,N_8234,N_8302);
nor U8467 (N_8467,N_8209,N_8202);
nand U8468 (N_8468,N_8330,N_8275);
and U8469 (N_8469,N_8310,N_8361);
nand U8470 (N_8470,N_8348,N_8292);
xor U8471 (N_8471,N_8334,N_8377);
or U8472 (N_8472,N_8242,N_8383);
or U8473 (N_8473,N_8303,N_8395);
or U8474 (N_8474,N_8267,N_8342);
and U8475 (N_8475,N_8353,N_8296);
xnor U8476 (N_8476,N_8366,N_8364);
nand U8477 (N_8477,N_8308,N_8252);
and U8478 (N_8478,N_8206,N_8258);
nand U8479 (N_8479,N_8386,N_8335);
nand U8480 (N_8480,N_8390,N_8238);
and U8481 (N_8481,N_8223,N_8245);
nor U8482 (N_8482,N_8381,N_8270);
nor U8483 (N_8483,N_8306,N_8211);
nor U8484 (N_8484,N_8220,N_8251);
or U8485 (N_8485,N_8287,N_8379);
nor U8486 (N_8486,N_8319,N_8371);
nand U8487 (N_8487,N_8305,N_8243);
and U8488 (N_8488,N_8299,N_8351);
nand U8489 (N_8489,N_8393,N_8369);
nand U8490 (N_8490,N_8331,N_8309);
nand U8491 (N_8491,N_8337,N_8236);
nand U8492 (N_8492,N_8208,N_8307);
nor U8493 (N_8493,N_8204,N_8328);
or U8494 (N_8494,N_8372,N_8391);
xnor U8495 (N_8495,N_8290,N_8375);
or U8496 (N_8496,N_8261,N_8321);
and U8497 (N_8497,N_8311,N_8253);
and U8498 (N_8498,N_8257,N_8336);
or U8499 (N_8499,N_8291,N_8315);
and U8500 (N_8500,N_8208,N_8246);
xor U8501 (N_8501,N_8397,N_8331);
xor U8502 (N_8502,N_8275,N_8300);
nor U8503 (N_8503,N_8300,N_8242);
nor U8504 (N_8504,N_8251,N_8364);
or U8505 (N_8505,N_8299,N_8270);
and U8506 (N_8506,N_8291,N_8369);
or U8507 (N_8507,N_8200,N_8237);
xor U8508 (N_8508,N_8370,N_8326);
or U8509 (N_8509,N_8231,N_8202);
or U8510 (N_8510,N_8221,N_8215);
nor U8511 (N_8511,N_8218,N_8216);
nor U8512 (N_8512,N_8236,N_8397);
or U8513 (N_8513,N_8364,N_8291);
xnor U8514 (N_8514,N_8249,N_8393);
or U8515 (N_8515,N_8226,N_8246);
and U8516 (N_8516,N_8326,N_8235);
or U8517 (N_8517,N_8391,N_8239);
and U8518 (N_8518,N_8208,N_8248);
or U8519 (N_8519,N_8387,N_8335);
or U8520 (N_8520,N_8200,N_8389);
nor U8521 (N_8521,N_8252,N_8379);
and U8522 (N_8522,N_8327,N_8268);
xnor U8523 (N_8523,N_8289,N_8357);
nand U8524 (N_8524,N_8217,N_8228);
nor U8525 (N_8525,N_8288,N_8341);
and U8526 (N_8526,N_8255,N_8288);
and U8527 (N_8527,N_8337,N_8392);
nor U8528 (N_8528,N_8347,N_8313);
nor U8529 (N_8529,N_8202,N_8381);
xor U8530 (N_8530,N_8367,N_8225);
xnor U8531 (N_8531,N_8303,N_8363);
or U8532 (N_8532,N_8271,N_8320);
and U8533 (N_8533,N_8256,N_8270);
nand U8534 (N_8534,N_8270,N_8266);
nand U8535 (N_8535,N_8261,N_8310);
nand U8536 (N_8536,N_8396,N_8255);
xnor U8537 (N_8537,N_8311,N_8263);
and U8538 (N_8538,N_8270,N_8293);
nand U8539 (N_8539,N_8234,N_8225);
xnor U8540 (N_8540,N_8258,N_8343);
and U8541 (N_8541,N_8346,N_8224);
and U8542 (N_8542,N_8379,N_8201);
nand U8543 (N_8543,N_8224,N_8306);
and U8544 (N_8544,N_8373,N_8384);
and U8545 (N_8545,N_8351,N_8267);
or U8546 (N_8546,N_8236,N_8386);
nor U8547 (N_8547,N_8269,N_8366);
nor U8548 (N_8548,N_8223,N_8227);
nor U8549 (N_8549,N_8269,N_8354);
nand U8550 (N_8550,N_8325,N_8260);
and U8551 (N_8551,N_8375,N_8306);
nand U8552 (N_8552,N_8387,N_8357);
and U8553 (N_8553,N_8271,N_8329);
nor U8554 (N_8554,N_8308,N_8355);
and U8555 (N_8555,N_8342,N_8221);
nor U8556 (N_8556,N_8359,N_8370);
nor U8557 (N_8557,N_8312,N_8363);
nand U8558 (N_8558,N_8365,N_8257);
and U8559 (N_8559,N_8371,N_8342);
nor U8560 (N_8560,N_8247,N_8313);
or U8561 (N_8561,N_8276,N_8287);
or U8562 (N_8562,N_8326,N_8262);
nand U8563 (N_8563,N_8230,N_8290);
xnor U8564 (N_8564,N_8327,N_8292);
nor U8565 (N_8565,N_8269,N_8389);
nand U8566 (N_8566,N_8308,N_8307);
nand U8567 (N_8567,N_8355,N_8254);
nand U8568 (N_8568,N_8393,N_8268);
nand U8569 (N_8569,N_8259,N_8235);
or U8570 (N_8570,N_8224,N_8266);
or U8571 (N_8571,N_8255,N_8384);
nor U8572 (N_8572,N_8256,N_8295);
or U8573 (N_8573,N_8214,N_8242);
xor U8574 (N_8574,N_8361,N_8206);
nor U8575 (N_8575,N_8334,N_8258);
or U8576 (N_8576,N_8364,N_8242);
or U8577 (N_8577,N_8328,N_8205);
and U8578 (N_8578,N_8269,N_8232);
or U8579 (N_8579,N_8229,N_8349);
or U8580 (N_8580,N_8379,N_8376);
or U8581 (N_8581,N_8298,N_8315);
and U8582 (N_8582,N_8391,N_8236);
nand U8583 (N_8583,N_8245,N_8244);
nand U8584 (N_8584,N_8389,N_8275);
and U8585 (N_8585,N_8358,N_8345);
and U8586 (N_8586,N_8343,N_8346);
nor U8587 (N_8587,N_8380,N_8277);
or U8588 (N_8588,N_8351,N_8359);
nand U8589 (N_8589,N_8245,N_8318);
and U8590 (N_8590,N_8314,N_8393);
or U8591 (N_8591,N_8261,N_8269);
or U8592 (N_8592,N_8385,N_8260);
nand U8593 (N_8593,N_8370,N_8297);
nor U8594 (N_8594,N_8217,N_8378);
xnor U8595 (N_8595,N_8235,N_8389);
or U8596 (N_8596,N_8387,N_8274);
nand U8597 (N_8597,N_8205,N_8355);
nand U8598 (N_8598,N_8353,N_8286);
nor U8599 (N_8599,N_8293,N_8211);
or U8600 (N_8600,N_8409,N_8485);
xnor U8601 (N_8601,N_8447,N_8508);
nor U8602 (N_8602,N_8595,N_8519);
nand U8603 (N_8603,N_8599,N_8449);
and U8604 (N_8604,N_8428,N_8510);
or U8605 (N_8605,N_8443,N_8507);
nor U8606 (N_8606,N_8451,N_8582);
nand U8607 (N_8607,N_8520,N_8453);
nand U8608 (N_8608,N_8536,N_8413);
xnor U8609 (N_8609,N_8432,N_8506);
and U8610 (N_8610,N_8526,N_8579);
nand U8611 (N_8611,N_8516,N_8544);
xnor U8612 (N_8612,N_8465,N_8406);
xor U8613 (N_8613,N_8431,N_8515);
or U8614 (N_8614,N_8546,N_8484);
nand U8615 (N_8615,N_8521,N_8437);
nand U8616 (N_8616,N_8532,N_8542);
nand U8617 (N_8617,N_8573,N_8466);
or U8618 (N_8618,N_8498,N_8421);
nand U8619 (N_8619,N_8505,N_8408);
and U8620 (N_8620,N_8429,N_8486);
or U8621 (N_8621,N_8407,N_8514);
nand U8622 (N_8622,N_8540,N_8558);
nand U8623 (N_8623,N_8524,N_8561);
xor U8624 (N_8624,N_8433,N_8403);
and U8625 (N_8625,N_8400,N_8441);
or U8626 (N_8626,N_8489,N_8559);
nand U8627 (N_8627,N_8473,N_8461);
or U8628 (N_8628,N_8446,N_8477);
nand U8629 (N_8629,N_8412,N_8419);
or U8630 (N_8630,N_8490,N_8450);
and U8631 (N_8631,N_8464,N_8454);
or U8632 (N_8632,N_8550,N_8530);
xnor U8633 (N_8633,N_8534,N_8469);
and U8634 (N_8634,N_8590,N_8493);
nand U8635 (N_8635,N_8455,N_8497);
nand U8636 (N_8636,N_8523,N_8420);
nor U8637 (N_8637,N_8517,N_8492);
and U8638 (N_8638,N_8404,N_8525);
or U8639 (N_8639,N_8456,N_8488);
or U8640 (N_8640,N_8528,N_8538);
or U8641 (N_8641,N_8541,N_8402);
and U8642 (N_8642,N_8576,N_8584);
xnor U8643 (N_8643,N_8462,N_8448);
nor U8644 (N_8644,N_8480,N_8504);
nand U8645 (N_8645,N_8598,N_8591);
or U8646 (N_8646,N_8487,N_8416);
nor U8647 (N_8647,N_8569,N_8588);
nor U8648 (N_8648,N_8518,N_8439);
nand U8649 (N_8649,N_8557,N_8499);
nand U8650 (N_8650,N_8460,N_8470);
or U8651 (N_8651,N_8452,N_8405);
nand U8652 (N_8652,N_8549,N_8483);
nor U8653 (N_8653,N_8552,N_8430);
xnor U8654 (N_8654,N_8537,N_8572);
and U8655 (N_8655,N_8543,N_8425);
and U8656 (N_8656,N_8539,N_8435);
nand U8657 (N_8657,N_8568,N_8442);
nand U8658 (N_8658,N_8494,N_8501);
or U8659 (N_8659,N_8424,N_8445);
nand U8660 (N_8660,N_8545,N_8596);
nand U8661 (N_8661,N_8531,N_8468);
and U8662 (N_8662,N_8535,N_8575);
nand U8663 (N_8663,N_8580,N_8463);
or U8664 (N_8664,N_8556,N_8597);
and U8665 (N_8665,N_8411,N_8555);
or U8666 (N_8666,N_8586,N_8589);
nand U8667 (N_8667,N_8417,N_8512);
nor U8668 (N_8668,N_8423,N_8436);
nor U8669 (N_8669,N_8482,N_8458);
xnor U8670 (N_8670,N_8566,N_8562);
or U8671 (N_8671,N_8410,N_8427);
and U8672 (N_8672,N_8503,N_8509);
xnor U8673 (N_8673,N_8592,N_8476);
or U8674 (N_8674,N_8438,N_8481);
nand U8675 (N_8675,N_8472,N_8583);
nand U8676 (N_8676,N_8511,N_8457);
or U8677 (N_8677,N_8578,N_8585);
and U8678 (N_8678,N_8444,N_8587);
nand U8679 (N_8679,N_8554,N_8434);
and U8680 (N_8680,N_8567,N_8467);
nor U8681 (N_8681,N_8522,N_8594);
or U8682 (N_8682,N_8414,N_8529);
and U8683 (N_8683,N_8496,N_8547);
nor U8684 (N_8684,N_8574,N_8495);
or U8685 (N_8685,N_8513,N_8564);
nand U8686 (N_8686,N_8581,N_8563);
or U8687 (N_8687,N_8593,N_8415);
nor U8688 (N_8688,N_8502,N_8565);
or U8689 (N_8689,N_8475,N_8570);
and U8690 (N_8690,N_8551,N_8533);
nor U8691 (N_8691,N_8479,N_8571);
and U8692 (N_8692,N_8418,N_8459);
xor U8693 (N_8693,N_8471,N_8440);
nor U8694 (N_8694,N_8548,N_8500);
nand U8695 (N_8695,N_8553,N_8491);
xnor U8696 (N_8696,N_8560,N_8478);
nand U8697 (N_8697,N_8401,N_8422);
nand U8698 (N_8698,N_8426,N_8474);
nand U8699 (N_8699,N_8527,N_8577);
nor U8700 (N_8700,N_8569,N_8538);
and U8701 (N_8701,N_8551,N_8528);
and U8702 (N_8702,N_8472,N_8475);
xor U8703 (N_8703,N_8564,N_8586);
nand U8704 (N_8704,N_8479,N_8568);
or U8705 (N_8705,N_8547,N_8555);
xnor U8706 (N_8706,N_8498,N_8439);
or U8707 (N_8707,N_8533,N_8538);
nor U8708 (N_8708,N_8500,N_8524);
and U8709 (N_8709,N_8554,N_8414);
nand U8710 (N_8710,N_8593,N_8579);
nor U8711 (N_8711,N_8511,N_8509);
and U8712 (N_8712,N_8512,N_8582);
nor U8713 (N_8713,N_8497,N_8450);
and U8714 (N_8714,N_8453,N_8561);
nand U8715 (N_8715,N_8563,N_8409);
nand U8716 (N_8716,N_8573,N_8550);
xor U8717 (N_8717,N_8433,N_8595);
nor U8718 (N_8718,N_8560,N_8584);
and U8719 (N_8719,N_8532,N_8545);
xor U8720 (N_8720,N_8512,N_8446);
nand U8721 (N_8721,N_8409,N_8535);
nor U8722 (N_8722,N_8502,N_8597);
or U8723 (N_8723,N_8558,N_8429);
or U8724 (N_8724,N_8507,N_8432);
and U8725 (N_8725,N_8594,N_8527);
or U8726 (N_8726,N_8543,N_8563);
and U8727 (N_8727,N_8427,N_8593);
nor U8728 (N_8728,N_8478,N_8481);
xor U8729 (N_8729,N_8570,N_8487);
nand U8730 (N_8730,N_8484,N_8463);
or U8731 (N_8731,N_8545,N_8444);
and U8732 (N_8732,N_8503,N_8464);
or U8733 (N_8733,N_8537,N_8418);
xnor U8734 (N_8734,N_8410,N_8423);
and U8735 (N_8735,N_8415,N_8466);
nand U8736 (N_8736,N_8521,N_8461);
xnor U8737 (N_8737,N_8454,N_8492);
or U8738 (N_8738,N_8496,N_8454);
and U8739 (N_8739,N_8518,N_8406);
and U8740 (N_8740,N_8508,N_8527);
nand U8741 (N_8741,N_8598,N_8434);
nand U8742 (N_8742,N_8464,N_8431);
or U8743 (N_8743,N_8411,N_8446);
and U8744 (N_8744,N_8478,N_8409);
nand U8745 (N_8745,N_8405,N_8420);
or U8746 (N_8746,N_8507,N_8470);
nor U8747 (N_8747,N_8415,N_8426);
nand U8748 (N_8748,N_8518,N_8420);
nand U8749 (N_8749,N_8455,N_8427);
xor U8750 (N_8750,N_8582,N_8401);
xor U8751 (N_8751,N_8459,N_8432);
or U8752 (N_8752,N_8577,N_8438);
nand U8753 (N_8753,N_8550,N_8406);
or U8754 (N_8754,N_8567,N_8579);
nor U8755 (N_8755,N_8569,N_8408);
nor U8756 (N_8756,N_8512,N_8485);
xor U8757 (N_8757,N_8481,N_8480);
nor U8758 (N_8758,N_8533,N_8436);
nor U8759 (N_8759,N_8413,N_8505);
or U8760 (N_8760,N_8510,N_8508);
nor U8761 (N_8761,N_8574,N_8483);
nor U8762 (N_8762,N_8599,N_8563);
or U8763 (N_8763,N_8561,N_8547);
nor U8764 (N_8764,N_8486,N_8572);
or U8765 (N_8765,N_8468,N_8599);
nor U8766 (N_8766,N_8566,N_8548);
nand U8767 (N_8767,N_8598,N_8510);
and U8768 (N_8768,N_8576,N_8482);
or U8769 (N_8769,N_8482,N_8418);
and U8770 (N_8770,N_8538,N_8522);
nand U8771 (N_8771,N_8553,N_8442);
xnor U8772 (N_8772,N_8539,N_8586);
and U8773 (N_8773,N_8427,N_8516);
nor U8774 (N_8774,N_8442,N_8428);
and U8775 (N_8775,N_8544,N_8534);
xor U8776 (N_8776,N_8509,N_8455);
nand U8777 (N_8777,N_8560,N_8470);
and U8778 (N_8778,N_8439,N_8536);
nand U8779 (N_8779,N_8593,N_8598);
nor U8780 (N_8780,N_8428,N_8597);
or U8781 (N_8781,N_8558,N_8482);
nor U8782 (N_8782,N_8580,N_8548);
nand U8783 (N_8783,N_8558,N_8566);
and U8784 (N_8784,N_8440,N_8439);
xor U8785 (N_8785,N_8459,N_8458);
nand U8786 (N_8786,N_8511,N_8561);
and U8787 (N_8787,N_8599,N_8439);
or U8788 (N_8788,N_8565,N_8409);
or U8789 (N_8789,N_8587,N_8530);
or U8790 (N_8790,N_8569,N_8472);
xnor U8791 (N_8791,N_8435,N_8544);
nor U8792 (N_8792,N_8519,N_8590);
and U8793 (N_8793,N_8552,N_8536);
or U8794 (N_8794,N_8575,N_8476);
nand U8795 (N_8795,N_8572,N_8544);
nand U8796 (N_8796,N_8425,N_8481);
nor U8797 (N_8797,N_8445,N_8550);
and U8798 (N_8798,N_8496,N_8539);
and U8799 (N_8799,N_8430,N_8410);
nand U8800 (N_8800,N_8745,N_8629);
and U8801 (N_8801,N_8677,N_8656);
nor U8802 (N_8802,N_8681,N_8647);
and U8803 (N_8803,N_8796,N_8726);
or U8804 (N_8804,N_8604,N_8756);
or U8805 (N_8805,N_8637,N_8746);
nor U8806 (N_8806,N_8760,N_8625);
nand U8807 (N_8807,N_8739,N_8742);
and U8808 (N_8808,N_8612,N_8731);
or U8809 (N_8809,N_8725,N_8697);
and U8810 (N_8810,N_8732,N_8646);
nand U8811 (N_8811,N_8668,N_8722);
nor U8812 (N_8812,N_8737,N_8605);
nor U8813 (N_8813,N_8696,N_8684);
xnor U8814 (N_8814,N_8617,N_8773);
nand U8815 (N_8815,N_8702,N_8657);
nor U8816 (N_8816,N_8601,N_8782);
nand U8817 (N_8817,N_8688,N_8627);
nor U8818 (N_8818,N_8631,N_8609);
nor U8819 (N_8819,N_8633,N_8636);
nand U8820 (N_8820,N_8680,N_8664);
and U8821 (N_8821,N_8772,N_8670);
nor U8822 (N_8822,N_8744,N_8717);
nand U8823 (N_8823,N_8660,N_8706);
nor U8824 (N_8824,N_8761,N_8762);
xor U8825 (N_8825,N_8768,N_8751);
nand U8826 (N_8826,N_8630,N_8614);
xor U8827 (N_8827,N_8603,N_8775);
and U8828 (N_8828,N_8683,N_8623);
xnor U8829 (N_8829,N_8784,N_8735);
or U8830 (N_8830,N_8634,N_8749);
or U8831 (N_8831,N_8750,N_8776);
nand U8832 (N_8832,N_8606,N_8618);
nand U8833 (N_8833,N_8686,N_8723);
nor U8834 (N_8834,N_8610,N_8771);
and U8835 (N_8835,N_8619,N_8705);
nor U8836 (N_8836,N_8758,N_8797);
or U8837 (N_8837,N_8753,N_8778);
or U8838 (N_8838,N_8695,N_8724);
nor U8839 (N_8839,N_8691,N_8645);
or U8840 (N_8840,N_8767,N_8755);
nand U8841 (N_8841,N_8651,N_8792);
xor U8842 (N_8842,N_8653,N_8798);
nor U8843 (N_8843,N_8787,N_8626);
or U8844 (N_8844,N_8632,N_8710);
nor U8845 (N_8845,N_8790,N_8788);
nor U8846 (N_8846,N_8665,N_8766);
and U8847 (N_8847,N_8687,N_8678);
xnor U8848 (N_8848,N_8716,N_8712);
xnor U8849 (N_8849,N_8639,N_8689);
nor U8850 (N_8850,N_8765,N_8690);
or U8851 (N_8851,N_8714,N_8621);
nand U8852 (N_8852,N_8780,N_8770);
nor U8853 (N_8853,N_8611,N_8613);
xor U8854 (N_8854,N_8764,N_8779);
nor U8855 (N_8855,N_8707,N_8703);
nor U8856 (N_8856,N_8777,N_8669);
or U8857 (N_8857,N_8718,N_8640);
nand U8858 (N_8858,N_8786,N_8644);
or U8859 (N_8859,N_8781,N_8659);
xor U8860 (N_8860,N_8715,N_8700);
or U8861 (N_8861,N_8728,N_8704);
or U8862 (N_8862,N_8616,N_8622);
and U8863 (N_8863,N_8675,N_8738);
and U8864 (N_8864,N_8602,N_8789);
xnor U8865 (N_8865,N_8662,N_8661);
nor U8866 (N_8866,N_8763,N_8673);
xnor U8867 (N_8867,N_8729,N_8628);
or U8868 (N_8868,N_8600,N_8711);
nand U8869 (N_8869,N_8652,N_8692);
or U8870 (N_8870,N_8783,N_8672);
or U8871 (N_8871,N_8685,N_8655);
and U8872 (N_8872,N_8709,N_8733);
xnor U8873 (N_8873,N_8795,N_8720);
nor U8874 (N_8874,N_8701,N_8615);
nor U8875 (N_8875,N_8693,N_8757);
nor U8876 (N_8876,N_8769,N_8649);
or U8877 (N_8877,N_8747,N_8667);
or U8878 (N_8878,N_8740,N_8799);
nor U8879 (N_8879,N_8791,N_8643);
and U8880 (N_8880,N_8794,N_8793);
or U8881 (N_8881,N_8620,N_8694);
nor U8882 (N_8882,N_8642,N_8682);
nand U8883 (N_8883,N_8650,N_8727);
or U8884 (N_8884,N_8759,N_8785);
nand U8885 (N_8885,N_8607,N_8699);
and U8886 (N_8886,N_8721,N_8736);
nor U8887 (N_8887,N_8635,N_8654);
or U8888 (N_8888,N_8679,N_8658);
and U8889 (N_8889,N_8752,N_8641);
nand U8890 (N_8890,N_8719,N_8754);
or U8891 (N_8891,N_8730,N_8741);
nor U8892 (N_8892,N_8666,N_8676);
nor U8893 (N_8893,N_8663,N_8608);
and U8894 (N_8894,N_8698,N_8648);
nand U8895 (N_8895,N_8743,N_8748);
or U8896 (N_8896,N_8734,N_8638);
nor U8897 (N_8897,N_8671,N_8674);
nand U8898 (N_8898,N_8708,N_8713);
and U8899 (N_8899,N_8624,N_8774);
and U8900 (N_8900,N_8758,N_8780);
nand U8901 (N_8901,N_8742,N_8759);
nand U8902 (N_8902,N_8674,N_8799);
nor U8903 (N_8903,N_8773,N_8629);
and U8904 (N_8904,N_8672,N_8671);
and U8905 (N_8905,N_8696,N_8765);
and U8906 (N_8906,N_8615,N_8734);
nor U8907 (N_8907,N_8686,N_8617);
nor U8908 (N_8908,N_8710,N_8649);
nand U8909 (N_8909,N_8756,N_8628);
nor U8910 (N_8910,N_8779,N_8677);
nand U8911 (N_8911,N_8692,N_8623);
or U8912 (N_8912,N_8737,N_8728);
or U8913 (N_8913,N_8692,N_8723);
nand U8914 (N_8914,N_8642,N_8746);
nand U8915 (N_8915,N_8708,N_8718);
or U8916 (N_8916,N_8731,N_8661);
nand U8917 (N_8917,N_8630,N_8618);
and U8918 (N_8918,N_8751,N_8680);
or U8919 (N_8919,N_8756,N_8702);
and U8920 (N_8920,N_8723,N_8713);
xor U8921 (N_8921,N_8678,N_8755);
nor U8922 (N_8922,N_8637,N_8788);
nor U8923 (N_8923,N_8730,N_8700);
xnor U8924 (N_8924,N_8771,N_8743);
nand U8925 (N_8925,N_8616,N_8777);
and U8926 (N_8926,N_8795,N_8721);
nor U8927 (N_8927,N_8793,N_8614);
nor U8928 (N_8928,N_8699,N_8788);
and U8929 (N_8929,N_8695,N_8723);
nor U8930 (N_8930,N_8746,N_8748);
nor U8931 (N_8931,N_8714,N_8623);
nor U8932 (N_8932,N_8713,N_8734);
and U8933 (N_8933,N_8607,N_8787);
and U8934 (N_8934,N_8776,N_8723);
nand U8935 (N_8935,N_8702,N_8757);
nand U8936 (N_8936,N_8727,N_8776);
or U8937 (N_8937,N_8617,N_8731);
nand U8938 (N_8938,N_8669,N_8795);
and U8939 (N_8939,N_8620,N_8708);
xnor U8940 (N_8940,N_8674,N_8751);
nor U8941 (N_8941,N_8699,N_8700);
or U8942 (N_8942,N_8788,N_8666);
and U8943 (N_8943,N_8603,N_8633);
nand U8944 (N_8944,N_8758,N_8793);
or U8945 (N_8945,N_8662,N_8632);
or U8946 (N_8946,N_8795,N_8772);
or U8947 (N_8947,N_8731,N_8649);
nor U8948 (N_8948,N_8784,N_8606);
or U8949 (N_8949,N_8654,N_8600);
nor U8950 (N_8950,N_8768,N_8747);
nand U8951 (N_8951,N_8704,N_8662);
and U8952 (N_8952,N_8708,N_8645);
nor U8953 (N_8953,N_8759,N_8772);
nand U8954 (N_8954,N_8664,N_8704);
and U8955 (N_8955,N_8645,N_8760);
xor U8956 (N_8956,N_8630,N_8612);
xor U8957 (N_8957,N_8632,N_8732);
nand U8958 (N_8958,N_8633,N_8662);
and U8959 (N_8959,N_8739,N_8609);
or U8960 (N_8960,N_8730,N_8793);
xor U8961 (N_8961,N_8726,N_8673);
xor U8962 (N_8962,N_8700,N_8681);
xnor U8963 (N_8963,N_8691,N_8667);
nor U8964 (N_8964,N_8626,N_8768);
nand U8965 (N_8965,N_8725,N_8617);
nor U8966 (N_8966,N_8781,N_8726);
nand U8967 (N_8967,N_8676,N_8724);
nand U8968 (N_8968,N_8796,N_8636);
and U8969 (N_8969,N_8756,N_8796);
nand U8970 (N_8970,N_8677,N_8654);
xnor U8971 (N_8971,N_8770,N_8718);
and U8972 (N_8972,N_8775,N_8654);
or U8973 (N_8973,N_8789,N_8675);
nor U8974 (N_8974,N_8756,N_8754);
nor U8975 (N_8975,N_8705,N_8656);
nand U8976 (N_8976,N_8710,N_8739);
nand U8977 (N_8977,N_8746,N_8738);
or U8978 (N_8978,N_8719,N_8627);
nor U8979 (N_8979,N_8707,N_8749);
and U8980 (N_8980,N_8784,N_8778);
nor U8981 (N_8981,N_8648,N_8711);
or U8982 (N_8982,N_8721,N_8603);
nand U8983 (N_8983,N_8613,N_8796);
or U8984 (N_8984,N_8659,N_8622);
or U8985 (N_8985,N_8612,N_8655);
nor U8986 (N_8986,N_8696,N_8640);
and U8987 (N_8987,N_8689,N_8779);
nor U8988 (N_8988,N_8639,N_8649);
nor U8989 (N_8989,N_8799,N_8615);
and U8990 (N_8990,N_8634,N_8707);
nand U8991 (N_8991,N_8732,N_8758);
and U8992 (N_8992,N_8775,N_8688);
and U8993 (N_8993,N_8724,N_8704);
and U8994 (N_8994,N_8684,N_8660);
nand U8995 (N_8995,N_8667,N_8692);
and U8996 (N_8996,N_8644,N_8654);
xor U8997 (N_8997,N_8691,N_8799);
and U8998 (N_8998,N_8706,N_8762);
or U8999 (N_8999,N_8712,N_8679);
xor U9000 (N_9000,N_8990,N_8959);
and U9001 (N_9001,N_8930,N_8865);
or U9002 (N_9002,N_8879,N_8999);
nand U9003 (N_9003,N_8881,N_8978);
and U9004 (N_9004,N_8892,N_8972);
or U9005 (N_9005,N_8920,N_8962);
nand U9006 (N_9006,N_8989,N_8973);
nand U9007 (N_9007,N_8827,N_8897);
nand U9008 (N_9008,N_8885,N_8853);
or U9009 (N_9009,N_8835,N_8814);
nand U9010 (N_9010,N_8900,N_8954);
or U9011 (N_9011,N_8826,N_8913);
xnor U9012 (N_9012,N_8816,N_8822);
or U9013 (N_9013,N_8910,N_8833);
or U9014 (N_9014,N_8874,N_8926);
or U9015 (N_9015,N_8950,N_8902);
nor U9016 (N_9016,N_8915,N_8958);
and U9017 (N_9017,N_8880,N_8831);
nor U9018 (N_9018,N_8832,N_8839);
nor U9019 (N_9019,N_8936,N_8840);
or U9020 (N_9020,N_8801,N_8849);
xnor U9021 (N_9021,N_8825,N_8955);
and U9022 (N_9022,N_8875,N_8838);
nand U9023 (N_9023,N_8993,N_8951);
and U9024 (N_9024,N_8846,N_8809);
or U9025 (N_9025,N_8909,N_8906);
nor U9026 (N_9026,N_8983,N_8802);
and U9027 (N_9027,N_8903,N_8981);
or U9028 (N_9028,N_8933,N_8937);
nand U9029 (N_9029,N_8922,N_8995);
nor U9030 (N_9030,N_8997,N_8883);
nor U9031 (N_9031,N_8800,N_8948);
nand U9032 (N_9032,N_8975,N_8908);
nand U9033 (N_9033,N_8985,N_8867);
nor U9034 (N_9034,N_8970,N_8817);
nand U9035 (N_9035,N_8858,N_8977);
xnor U9036 (N_9036,N_8842,N_8984);
or U9037 (N_9037,N_8851,N_8919);
nor U9038 (N_9038,N_8843,N_8847);
or U9039 (N_9039,N_8864,N_8859);
and U9040 (N_9040,N_8890,N_8956);
or U9041 (N_9041,N_8886,N_8911);
or U9042 (N_9042,N_8819,N_8882);
or U9043 (N_9043,N_8841,N_8961);
nor U9044 (N_9044,N_8855,N_8828);
nor U9045 (N_9045,N_8845,N_8872);
and U9046 (N_9046,N_8953,N_8812);
nand U9047 (N_9047,N_8969,N_8918);
nand U9048 (N_9048,N_8870,N_8974);
nand U9049 (N_9049,N_8965,N_8979);
nand U9050 (N_9050,N_8894,N_8863);
nand U9051 (N_9051,N_8952,N_8830);
or U9052 (N_9052,N_8884,N_8996);
nor U9053 (N_9053,N_8824,N_8813);
and U9054 (N_9054,N_8935,N_8986);
and U9055 (N_9055,N_8928,N_8807);
or U9056 (N_9056,N_8940,N_8980);
nand U9057 (N_9057,N_8811,N_8857);
and U9058 (N_9058,N_8925,N_8854);
nor U9059 (N_9059,N_8896,N_8901);
nand U9060 (N_9060,N_8806,N_8895);
and U9061 (N_9061,N_8967,N_8820);
or U9062 (N_9062,N_8907,N_8808);
xor U9063 (N_9063,N_8941,N_8861);
nor U9064 (N_9064,N_8866,N_8868);
xnor U9065 (N_9065,N_8850,N_8914);
nand U9066 (N_9066,N_8942,N_8966);
nor U9067 (N_9067,N_8960,N_8963);
xor U9068 (N_9068,N_8834,N_8932);
nor U9069 (N_9069,N_8804,N_8904);
xor U9070 (N_9070,N_8924,N_8994);
and U9071 (N_9071,N_8916,N_8887);
or U9072 (N_9072,N_8964,N_8856);
nor U9073 (N_9073,N_8899,N_8998);
nor U9074 (N_9074,N_8889,N_8823);
nand U9075 (N_9075,N_8957,N_8931);
xnor U9076 (N_9076,N_8905,N_8988);
or U9077 (N_9077,N_8876,N_8921);
nand U9078 (N_9078,N_8844,N_8968);
and U9079 (N_9079,N_8945,N_8992);
nor U9080 (N_9080,N_8938,N_8891);
and U9081 (N_9081,N_8982,N_8912);
and U9082 (N_9082,N_8943,N_8934);
nand U9083 (N_9083,N_8848,N_8818);
nand U9084 (N_9084,N_8987,N_8877);
or U9085 (N_9085,N_8991,N_8949);
nand U9086 (N_9086,N_8803,N_8927);
and U9087 (N_9087,N_8871,N_8946);
nand U9088 (N_9088,N_8829,N_8929);
and U9089 (N_9089,N_8810,N_8893);
xor U9090 (N_9090,N_8888,N_8878);
and U9091 (N_9091,N_8821,N_8923);
nor U9092 (N_9092,N_8971,N_8815);
xnor U9093 (N_9093,N_8939,N_8805);
and U9094 (N_9094,N_8917,N_8862);
or U9095 (N_9095,N_8869,N_8944);
xnor U9096 (N_9096,N_8873,N_8852);
or U9097 (N_9097,N_8860,N_8836);
or U9098 (N_9098,N_8898,N_8837);
xor U9099 (N_9099,N_8947,N_8976);
xor U9100 (N_9100,N_8822,N_8890);
xor U9101 (N_9101,N_8826,N_8951);
and U9102 (N_9102,N_8889,N_8992);
nand U9103 (N_9103,N_8910,N_8863);
nor U9104 (N_9104,N_8984,N_8880);
or U9105 (N_9105,N_8804,N_8999);
nand U9106 (N_9106,N_8864,N_8964);
nand U9107 (N_9107,N_8812,N_8887);
xor U9108 (N_9108,N_8802,N_8850);
nand U9109 (N_9109,N_8898,N_8882);
or U9110 (N_9110,N_8935,N_8808);
xor U9111 (N_9111,N_8960,N_8991);
or U9112 (N_9112,N_8900,N_8813);
or U9113 (N_9113,N_8894,N_8996);
xnor U9114 (N_9114,N_8881,N_8844);
or U9115 (N_9115,N_8954,N_8856);
or U9116 (N_9116,N_8990,N_8880);
nand U9117 (N_9117,N_8801,N_8810);
nand U9118 (N_9118,N_8845,N_8997);
nand U9119 (N_9119,N_8877,N_8988);
or U9120 (N_9120,N_8827,N_8842);
or U9121 (N_9121,N_8963,N_8866);
nor U9122 (N_9122,N_8945,N_8920);
and U9123 (N_9123,N_8842,N_8887);
or U9124 (N_9124,N_8805,N_8831);
nand U9125 (N_9125,N_8964,N_8851);
and U9126 (N_9126,N_8959,N_8921);
nand U9127 (N_9127,N_8918,N_8895);
nand U9128 (N_9128,N_8962,N_8963);
nor U9129 (N_9129,N_8847,N_8807);
and U9130 (N_9130,N_8907,N_8906);
or U9131 (N_9131,N_8837,N_8852);
and U9132 (N_9132,N_8949,N_8888);
nand U9133 (N_9133,N_8827,N_8880);
or U9134 (N_9134,N_8827,N_8919);
nand U9135 (N_9135,N_8821,N_8872);
nor U9136 (N_9136,N_8967,N_8823);
nand U9137 (N_9137,N_8962,N_8874);
and U9138 (N_9138,N_8873,N_8853);
xor U9139 (N_9139,N_8920,N_8805);
xnor U9140 (N_9140,N_8935,N_8800);
nor U9141 (N_9141,N_8980,N_8955);
and U9142 (N_9142,N_8940,N_8868);
nor U9143 (N_9143,N_8949,N_8994);
and U9144 (N_9144,N_8837,N_8873);
nor U9145 (N_9145,N_8820,N_8831);
and U9146 (N_9146,N_8951,N_8811);
and U9147 (N_9147,N_8862,N_8923);
xor U9148 (N_9148,N_8853,N_8825);
and U9149 (N_9149,N_8961,N_8908);
nand U9150 (N_9150,N_8853,N_8903);
or U9151 (N_9151,N_8995,N_8902);
or U9152 (N_9152,N_8848,N_8992);
nor U9153 (N_9153,N_8889,N_8951);
and U9154 (N_9154,N_8812,N_8840);
nor U9155 (N_9155,N_8946,N_8956);
nand U9156 (N_9156,N_8876,N_8936);
xor U9157 (N_9157,N_8898,N_8815);
nand U9158 (N_9158,N_8932,N_8960);
nor U9159 (N_9159,N_8948,N_8932);
and U9160 (N_9160,N_8852,N_8903);
nor U9161 (N_9161,N_8874,N_8916);
or U9162 (N_9162,N_8844,N_8987);
nand U9163 (N_9163,N_8804,N_8952);
nor U9164 (N_9164,N_8991,N_8889);
and U9165 (N_9165,N_8942,N_8890);
and U9166 (N_9166,N_8919,N_8964);
or U9167 (N_9167,N_8852,N_8861);
nor U9168 (N_9168,N_8896,N_8830);
or U9169 (N_9169,N_8807,N_8919);
or U9170 (N_9170,N_8862,N_8899);
nand U9171 (N_9171,N_8969,N_8919);
nand U9172 (N_9172,N_8903,N_8951);
and U9173 (N_9173,N_8885,N_8858);
nor U9174 (N_9174,N_8851,N_8812);
or U9175 (N_9175,N_8868,N_8852);
nor U9176 (N_9176,N_8997,N_8924);
nand U9177 (N_9177,N_8995,N_8934);
nand U9178 (N_9178,N_8862,N_8834);
nand U9179 (N_9179,N_8942,N_8897);
nor U9180 (N_9180,N_8983,N_8835);
nand U9181 (N_9181,N_8935,N_8882);
nand U9182 (N_9182,N_8900,N_8972);
xor U9183 (N_9183,N_8938,N_8846);
and U9184 (N_9184,N_8800,N_8896);
and U9185 (N_9185,N_8904,N_8828);
nand U9186 (N_9186,N_8903,N_8945);
and U9187 (N_9187,N_8910,N_8942);
nand U9188 (N_9188,N_8925,N_8832);
and U9189 (N_9189,N_8853,N_8921);
nor U9190 (N_9190,N_8839,N_8920);
and U9191 (N_9191,N_8803,N_8832);
nand U9192 (N_9192,N_8873,N_8818);
nor U9193 (N_9193,N_8950,N_8917);
and U9194 (N_9194,N_8856,N_8916);
nor U9195 (N_9195,N_8934,N_8834);
or U9196 (N_9196,N_8979,N_8947);
nand U9197 (N_9197,N_8947,N_8928);
and U9198 (N_9198,N_8953,N_8991);
and U9199 (N_9199,N_8897,N_8904);
xnor U9200 (N_9200,N_9158,N_9036);
or U9201 (N_9201,N_9092,N_9051);
and U9202 (N_9202,N_9166,N_9170);
xnor U9203 (N_9203,N_9186,N_9146);
and U9204 (N_9204,N_9098,N_9175);
or U9205 (N_9205,N_9193,N_9058);
or U9206 (N_9206,N_9142,N_9052);
nor U9207 (N_9207,N_9147,N_9129);
and U9208 (N_9208,N_9085,N_9014);
and U9209 (N_9209,N_9078,N_9178);
nor U9210 (N_9210,N_9019,N_9015);
and U9211 (N_9211,N_9114,N_9090);
or U9212 (N_9212,N_9160,N_9150);
xnor U9213 (N_9213,N_9159,N_9096);
or U9214 (N_9214,N_9057,N_9094);
and U9215 (N_9215,N_9174,N_9180);
nor U9216 (N_9216,N_9028,N_9105);
and U9217 (N_9217,N_9054,N_9034);
and U9218 (N_9218,N_9133,N_9115);
xor U9219 (N_9219,N_9177,N_9189);
and U9220 (N_9220,N_9139,N_9016);
or U9221 (N_9221,N_9012,N_9010);
nor U9222 (N_9222,N_9192,N_9125);
nor U9223 (N_9223,N_9006,N_9153);
nand U9224 (N_9224,N_9076,N_9070);
and U9225 (N_9225,N_9042,N_9065);
and U9226 (N_9226,N_9113,N_9097);
nand U9227 (N_9227,N_9009,N_9195);
nand U9228 (N_9228,N_9038,N_9182);
nand U9229 (N_9229,N_9173,N_9077);
and U9230 (N_9230,N_9049,N_9087);
nand U9231 (N_9231,N_9069,N_9055);
xor U9232 (N_9232,N_9183,N_9063);
nor U9233 (N_9233,N_9086,N_9068);
and U9234 (N_9234,N_9040,N_9020);
and U9235 (N_9235,N_9024,N_9171);
nor U9236 (N_9236,N_9141,N_9035);
or U9237 (N_9237,N_9145,N_9110);
or U9238 (N_9238,N_9001,N_9127);
nor U9239 (N_9239,N_9047,N_9167);
nand U9240 (N_9240,N_9067,N_9156);
or U9241 (N_9241,N_9190,N_9030);
or U9242 (N_9242,N_9025,N_9041);
and U9243 (N_9243,N_9196,N_9128);
nand U9244 (N_9244,N_9043,N_9199);
xor U9245 (N_9245,N_9108,N_9059);
or U9246 (N_9246,N_9187,N_9074);
or U9247 (N_9247,N_9168,N_9007);
nor U9248 (N_9248,N_9060,N_9053);
and U9249 (N_9249,N_9046,N_9045);
nand U9250 (N_9250,N_9002,N_9130);
or U9251 (N_9251,N_9037,N_9029);
or U9252 (N_9252,N_9104,N_9080);
and U9253 (N_9253,N_9138,N_9102);
xor U9254 (N_9254,N_9137,N_9197);
xor U9255 (N_9255,N_9164,N_9048);
nand U9256 (N_9256,N_9033,N_9152);
nor U9257 (N_9257,N_9022,N_9005);
nor U9258 (N_9258,N_9044,N_9120);
nand U9259 (N_9259,N_9000,N_9154);
nor U9260 (N_9260,N_9194,N_9091);
nor U9261 (N_9261,N_9017,N_9132);
and U9262 (N_9262,N_9191,N_9082);
nor U9263 (N_9263,N_9072,N_9172);
or U9264 (N_9264,N_9003,N_9032);
nand U9265 (N_9265,N_9123,N_9185);
xnor U9266 (N_9266,N_9008,N_9165);
nor U9267 (N_9267,N_9100,N_9026);
and U9268 (N_9268,N_9131,N_9179);
and U9269 (N_9269,N_9148,N_9103);
or U9270 (N_9270,N_9188,N_9136);
nor U9271 (N_9271,N_9056,N_9198);
nand U9272 (N_9272,N_9073,N_9140);
or U9273 (N_9273,N_9011,N_9089);
and U9274 (N_9274,N_9149,N_9004);
and U9275 (N_9275,N_9107,N_9101);
and U9276 (N_9276,N_9151,N_9112);
nand U9277 (N_9277,N_9181,N_9106);
nand U9278 (N_9278,N_9018,N_9162);
nor U9279 (N_9279,N_9117,N_9084);
and U9280 (N_9280,N_9121,N_9111);
and U9281 (N_9281,N_9116,N_9119);
nor U9282 (N_9282,N_9071,N_9050);
or U9283 (N_9283,N_9079,N_9013);
nor U9284 (N_9284,N_9161,N_9081);
or U9285 (N_9285,N_9031,N_9083);
nor U9286 (N_9286,N_9134,N_9066);
nor U9287 (N_9287,N_9155,N_9184);
and U9288 (N_9288,N_9144,N_9169);
nand U9289 (N_9289,N_9088,N_9118);
or U9290 (N_9290,N_9163,N_9099);
nor U9291 (N_9291,N_9109,N_9095);
or U9292 (N_9292,N_9126,N_9027);
nor U9293 (N_9293,N_9135,N_9124);
xnor U9294 (N_9294,N_9064,N_9176);
nor U9295 (N_9295,N_9061,N_9122);
and U9296 (N_9296,N_9062,N_9143);
and U9297 (N_9297,N_9157,N_9039);
or U9298 (N_9298,N_9021,N_9023);
or U9299 (N_9299,N_9075,N_9093);
or U9300 (N_9300,N_9056,N_9075);
nand U9301 (N_9301,N_9016,N_9081);
and U9302 (N_9302,N_9112,N_9001);
and U9303 (N_9303,N_9011,N_9149);
nor U9304 (N_9304,N_9147,N_9154);
nor U9305 (N_9305,N_9173,N_9110);
nor U9306 (N_9306,N_9184,N_9134);
or U9307 (N_9307,N_9161,N_9162);
xnor U9308 (N_9308,N_9078,N_9058);
nor U9309 (N_9309,N_9123,N_9012);
xor U9310 (N_9310,N_9032,N_9151);
and U9311 (N_9311,N_9139,N_9151);
nor U9312 (N_9312,N_9141,N_9156);
nand U9313 (N_9313,N_9145,N_9046);
or U9314 (N_9314,N_9010,N_9093);
and U9315 (N_9315,N_9018,N_9193);
and U9316 (N_9316,N_9140,N_9145);
nor U9317 (N_9317,N_9195,N_9180);
and U9318 (N_9318,N_9077,N_9115);
and U9319 (N_9319,N_9084,N_9154);
and U9320 (N_9320,N_9018,N_9087);
or U9321 (N_9321,N_9124,N_9187);
nor U9322 (N_9322,N_9106,N_9054);
nand U9323 (N_9323,N_9012,N_9058);
or U9324 (N_9324,N_9080,N_9052);
xnor U9325 (N_9325,N_9033,N_9092);
nor U9326 (N_9326,N_9100,N_9098);
or U9327 (N_9327,N_9122,N_9046);
or U9328 (N_9328,N_9049,N_9023);
nand U9329 (N_9329,N_9183,N_9114);
nand U9330 (N_9330,N_9170,N_9018);
or U9331 (N_9331,N_9098,N_9115);
xor U9332 (N_9332,N_9074,N_9001);
nand U9333 (N_9333,N_9096,N_9020);
and U9334 (N_9334,N_9193,N_9098);
or U9335 (N_9335,N_9117,N_9020);
nand U9336 (N_9336,N_9093,N_9005);
and U9337 (N_9337,N_9148,N_9170);
nor U9338 (N_9338,N_9072,N_9164);
or U9339 (N_9339,N_9055,N_9085);
and U9340 (N_9340,N_9196,N_9051);
or U9341 (N_9341,N_9130,N_9075);
nand U9342 (N_9342,N_9010,N_9187);
and U9343 (N_9343,N_9192,N_9188);
nor U9344 (N_9344,N_9066,N_9075);
nor U9345 (N_9345,N_9040,N_9013);
nor U9346 (N_9346,N_9049,N_9179);
nor U9347 (N_9347,N_9053,N_9127);
or U9348 (N_9348,N_9091,N_9096);
nor U9349 (N_9349,N_9044,N_9080);
nor U9350 (N_9350,N_9099,N_9094);
nor U9351 (N_9351,N_9194,N_9110);
or U9352 (N_9352,N_9151,N_9138);
nor U9353 (N_9353,N_9023,N_9197);
nor U9354 (N_9354,N_9076,N_9051);
nor U9355 (N_9355,N_9059,N_9105);
nor U9356 (N_9356,N_9148,N_9078);
nand U9357 (N_9357,N_9032,N_9016);
or U9358 (N_9358,N_9178,N_9183);
and U9359 (N_9359,N_9084,N_9040);
or U9360 (N_9360,N_9142,N_9176);
nor U9361 (N_9361,N_9031,N_9016);
or U9362 (N_9362,N_9184,N_9070);
and U9363 (N_9363,N_9135,N_9000);
or U9364 (N_9364,N_9034,N_9021);
and U9365 (N_9365,N_9025,N_9099);
nor U9366 (N_9366,N_9171,N_9195);
and U9367 (N_9367,N_9090,N_9016);
nor U9368 (N_9368,N_9087,N_9021);
xnor U9369 (N_9369,N_9041,N_9114);
and U9370 (N_9370,N_9134,N_9190);
or U9371 (N_9371,N_9077,N_9102);
or U9372 (N_9372,N_9164,N_9029);
or U9373 (N_9373,N_9174,N_9113);
nand U9374 (N_9374,N_9182,N_9104);
or U9375 (N_9375,N_9199,N_9154);
nand U9376 (N_9376,N_9053,N_9031);
nor U9377 (N_9377,N_9078,N_9014);
nor U9378 (N_9378,N_9040,N_9089);
nor U9379 (N_9379,N_9021,N_9163);
xnor U9380 (N_9380,N_9073,N_9052);
nor U9381 (N_9381,N_9179,N_9132);
nor U9382 (N_9382,N_9097,N_9091);
and U9383 (N_9383,N_9068,N_9159);
nand U9384 (N_9384,N_9123,N_9089);
xor U9385 (N_9385,N_9069,N_9045);
nand U9386 (N_9386,N_9196,N_9126);
and U9387 (N_9387,N_9154,N_9021);
or U9388 (N_9388,N_9158,N_9006);
and U9389 (N_9389,N_9076,N_9129);
xnor U9390 (N_9390,N_9128,N_9153);
nand U9391 (N_9391,N_9198,N_9045);
nand U9392 (N_9392,N_9057,N_9120);
xor U9393 (N_9393,N_9046,N_9124);
or U9394 (N_9394,N_9059,N_9197);
nor U9395 (N_9395,N_9037,N_9011);
and U9396 (N_9396,N_9186,N_9181);
and U9397 (N_9397,N_9140,N_9179);
and U9398 (N_9398,N_9020,N_9079);
xor U9399 (N_9399,N_9057,N_9030);
nor U9400 (N_9400,N_9322,N_9359);
xnor U9401 (N_9401,N_9270,N_9287);
and U9402 (N_9402,N_9386,N_9341);
xnor U9403 (N_9403,N_9210,N_9246);
and U9404 (N_9404,N_9297,N_9244);
nand U9405 (N_9405,N_9200,N_9222);
xnor U9406 (N_9406,N_9312,N_9294);
and U9407 (N_9407,N_9350,N_9230);
nand U9408 (N_9408,N_9353,N_9319);
and U9409 (N_9409,N_9371,N_9286);
and U9410 (N_9410,N_9311,N_9368);
or U9411 (N_9411,N_9226,N_9340);
nor U9412 (N_9412,N_9370,N_9225);
or U9413 (N_9413,N_9273,N_9292);
nand U9414 (N_9414,N_9289,N_9211);
xnor U9415 (N_9415,N_9253,N_9245);
or U9416 (N_9416,N_9261,N_9250);
or U9417 (N_9417,N_9399,N_9334);
nor U9418 (N_9418,N_9325,N_9260);
or U9419 (N_9419,N_9335,N_9393);
and U9420 (N_9420,N_9336,N_9252);
or U9421 (N_9421,N_9395,N_9299);
xor U9422 (N_9422,N_9378,N_9276);
nand U9423 (N_9423,N_9259,N_9229);
nor U9424 (N_9424,N_9362,N_9376);
nor U9425 (N_9425,N_9274,N_9249);
and U9426 (N_9426,N_9327,N_9218);
xnor U9427 (N_9427,N_9243,N_9234);
nor U9428 (N_9428,N_9381,N_9262);
xor U9429 (N_9429,N_9308,N_9313);
nand U9430 (N_9430,N_9347,N_9231);
and U9431 (N_9431,N_9221,N_9291);
nor U9432 (N_9432,N_9397,N_9365);
or U9433 (N_9433,N_9330,N_9387);
and U9434 (N_9434,N_9258,N_9235);
nand U9435 (N_9435,N_9254,N_9293);
and U9436 (N_9436,N_9315,N_9206);
and U9437 (N_9437,N_9236,N_9209);
nand U9438 (N_9438,N_9278,N_9346);
or U9439 (N_9439,N_9318,N_9317);
and U9440 (N_9440,N_9396,N_9267);
and U9441 (N_9441,N_9256,N_9279);
and U9442 (N_9442,N_9298,N_9323);
nor U9443 (N_9443,N_9329,N_9208);
or U9444 (N_9444,N_9344,N_9366);
nor U9445 (N_9445,N_9349,N_9382);
nor U9446 (N_9446,N_9374,N_9309);
nand U9447 (N_9447,N_9247,N_9272);
nand U9448 (N_9448,N_9332,N_9342);
or U9449 (N_9449,N_9338,N_9216);
nor U9450 (N_9450,N_9326,N_9324);
nand U9451 (N_9451,N_9392,N_9280);
and U9452 (N_9452,N_9360,N_9305);
xnor U9453 (N_9453,N_9288,N_9345);
nor U9454 (N_9454,N_9320,N_9214);
nor U9455 (N_9455,N_9224,N_9290);
and U9456 (N_9456,N_9277,N_9339);
nand U9457 (N_9457,N_9333,N_9390);
and U9458 (N_9458,N_9356,N_9275);
nor U9459 (N_9459,N_9369,N_9240);
or U9460 (N_9460,N_9331,N_9241);
or U9461 (N_9461,N_9266,N_9357);
xor U9462 (N_9462,N_9352,N_9358);
nand U9463 (N_9463,N_9367,N_9379);
nand U9464 (N_9464,N_9233,N_9373);
and U9465 (N_9465,N_9238,N_9219);
or U9466 (N_9466,N_9215,N_9377);
nor U9467 (N_9467,N_9282,N_9201);
nand U9468 (N_9468,N_9248,N_9296);
xnor U9469 (N_9469,N_9239,N_9316);
nand U9470 (N_9470,N_9281,N_9202);
nor U9471 (N_9471,N_9295,N_9394);
nor U9472 (N_9472,N_9355,N_9361);
xor U9473 (N_9473,N_9203,N_9284);
xor U9474 (N_9474,N_9337,N_9363);
and U9475 (N_9475,N_9265,N_9205);
nand U9476 (N_9476,N_9354,N_9237);
nor U9477 (N_9477,N_9257,N_9255);
xor U9478 (N_9478,N_9300,N_9398);
nand U9479 (N_9479,N_9391,N_9321);
nand U9480 (N_9480,N_9343,N_9271);
and U9481 (N_9481,N_9283,N_9348);
xor U9482 (N_9482,N_9372,N_9227);
nand U9483 (N_9483,N_9307,N_9306);
and U9484 (N_9484,N_9228,N_9213);
or U9485 (N_9485,N_9251,N_9351);
and U9486 (N_9486,N_9383,N_9328);
nor U9487 (N_9487,N_9384,N_9204);
xnor U9488 (N_9488,N_9310,N_9304);
xnor U9489 (N_9489,N_9223,N_9388);
xor U9490 (N_9490,N_9264,N_9385);
and U9491 (N_9491,N_9220,N_9301);
or U9492 (N_9492,N_9242,N_9232);
and U9493 (N_9493,N_9207,N_9302);
xor U9494 (N_9494,N_9389,N_9269);
or U9495 (N_9495,N_9217,N_9263);
and U9496 (N_9496,N_9364,N_9268);
nor U9497 (N_9497,N_9380,N_9303);
or U9498 (N_9498,N_9375,N_9314);
nand U9499 (N_9499,N_9212,N_9285);
nor U9500 (N_9500,N_9291,N_9378);
xor U9501 (N_9501,N_9335,N_9214);
nand U9502 (N_9502,N_9357,N_9271);
or U9503 (N_9503,N_9212,N_9395);
or U9504 (N_9504,N_9247,N_9239);
or U9505 (N_9505,N_9300,N_9307);
and U9506 (N_9506,N_9262,N_9320);
nor U9507 (N_9507,N_9292,N_9323);
xor U9508 (N_9508,N_9236,N_9363);
nand U9509 (N_9509,N_9226,N_9339);
nand U9510 (N_9510,N_9223,N_9363);
nor U9511 (N_9511,N_9261,N_9247);
and U9512 (N_9512,N_9298,N_9363);
nand U9513 (N_9513,N_9254,N_9233);
or U9514 (N_9514,N_9255,N_9352);
or U9515 (N_9515,N_9235,N_9307);
nand U9516 (N_9516,N_9359,N_9284);
nor U9517 (N_9517,N_9390,N_9257);
nor U9518 (N_9518,N_9398,N_9333);
nor U9519 (N_9519,N_9329,N_9211);
and U9520 (N_9520,N_9346,N_9358);
and U9521 (N_9521,N_9322,N_9278);
and U9522 (N_9522,N_9324,N_9397);
and U9523 (N_9523,N_9226,N_9236);
nand U9524 (N_9524,N_9215,N_9278);
xnor U9525 (N_9525,N_9304,N_9232);
or U9526 (N_9526,N_9231,N_9325);
or U9527 (N_9527,N_9330,N_9236);
and U9528 (N_9528,N_9349,N_9354);
nor U9529 (N_9529,N_9331,N_9232);
or U9530 (N_9530,N_9321,N_9294);
or U9531 (N_9531,N_9239,N_9360);
nor U9532 (N_9532,N_9268,N_9335);
and U9533 (N_9533,N_9348,N_9258);
and U9534 (N_9534,N_9351,N_9284);
and U9535 (N_9535,N_9315,N_9319);
nor U9536 (N_9536,N_9285,N_9272);
nand U9537 (N_9537,N_9235,N_9342);
nand U9538 (N_9538,N_9318,N_9311);
nor U9539 (N_9539,N_9245,N_9378);
or U9540 (N_9540,N_9351,N_9287);
nor U9541 (N_9541,N_9377,N_9385);
and U9542 (N_9542,N_9390,N_9227);
nor U9543 (N_9543,N_9239,N_9300);
or U9544 (N_9544,N_9223,N_9330);
or U9545 (N_9545,N_9393,N_9311);
nand U9546 (N_9546,N_9361,N_9222);
nor U9547 (N_9547,N_9351,N_9223);
nor U9548 (N_9548,N_9217,N_9270);
and U9549 (N_9549,N_9370,N_9368);
nor U9550 (N_9550,N_9217,N_9367);
and U9551 (N_9551,N_9359,N_9200);
nor U9552 (N_9552,N_9315,N_9379);
nor U9553 (N_9553,N_9340,N_9311);
and U9554 (N_9554,N_9288,N_9289);
or U9555 (N_9555,N_9287,N_9309);
or U9556 (N_9556,N_9372,N_9314);
or U9557 (N_9557,N_9225,N_9205);
nand U9558 (N_9558,N_9350,N_9254);
or U9559 (N_9559,N_9393,N_9278);
and U9560 (N_9560,N_9319,N_9261);
nor U9561 (N_9561,N_9277,N_9374);
nor U9562 (N_9562,N_9319,N_9284);
or U9563 (N_9563,N_9334,N_9331);
or U9564 (N_9564,N_9286,N_9378);
nand U9565 (N_9565,N_9341,N_9263);
or U9566 (N_9566,N_9378,N_9338);
nand U9567 (N_9567,N_9285,N_9208);
nand U9568 (N_9568,N_9360,N_9345);
nand U9569 (N_9569,N_9337,N_9357);
nand U9570 (N_9570,N_9326,N_9219);
xnor U9571 (N_9571,N_9369,N_9273);
or U9572 (N_9572,N_9377,N_9210);
nand U9573 (N_9573,N_9322,N_9337);
and U9574 (N_9574,N_9304,N_9221);
xnor U9575 (N_9575,N_9336,N_9239);
or U9576 (N_9576,N_9303,N_9342);
nor U9577 (N_9577,N_9294,N_9220);
or U9578 (N_9578,N_9258,N_9280);
nor U9579 (N_9579,N_9383,N_9243);
or U9580 (N_9580,N_9397,N_9316);
nand U9581 (N_9581,N_9274,N_9302);
nand U9582 (N_9582,N_9365,N_9217);
or U9583 (N_9583,N_9206,N_9385);
and U9584 (N_9584,N_9392,N_9272);
or U9585 (N_9585,N_9298,N_9320);
nand U9586 (N_9586,N_9387,N_9382);
nor U9587 (N_9587,N_9222,N_9226);
nor U9588 (N_9588,N_9267,N_9214);
and U9589 (N_9589,N_9393,N_9282);
nand U9590 (N_9590,N_9326,N_9305);
and U9591 (N_9591,N_9248,N_9250);
nand U9592 (N_9592,N_9251,N_9227);
nand U9593 (N_9593,N_9242,N_9207);
and U9594 (N_9594,N_9376,N_9388);
and U9595 (N_9595,N_9356,N_9369);
nand U9596 (N_9596,N_9350,N_9351);
and U9597 (N_9597,N_9398,N_9244);
or U9598 (N_9598,N_9383,N_9253);
and U9599 (N_9599,N_9322,N_9368);
xor U9600 (N_9600,N_9576,N_9435);
nand U9601 (N_9601,N_9565,N_9464);
xnor U9602 (N_9602,N_9506,N_9553);
xnor U9603 (N_9603,N_9561,N_9546);
and U9604 (N_9604,N_9491,N_9405);
xor U9605 (N_9605,N_9585,N_9407);
nor U9606 (N_9606,N_9467,N_9412);
or U9607 (N_9607,N_9566,N_9510);
nor U9608 (N_9608,N_9448,N_9595);
and U9609 (N_9609,N_9486,N_9423);
nor U9610 (N_9610,N_9589,N_9461);
xor U9611 (N_9611,N_9481,N_9430);
or U9612 (N_9612,N_9477,N_9426);
and U9613 (N_9613,N_9579,N_9493);
xor U9614 (N_9614,N_9413,N_9571);
and U9615 (N_9615,N_9534,N_9526);
or U9616 (N_9616,N_9568,N_9583);
nand U9617 (N_9617,N_9427,N_9508);
or U9618 (N_9618,N_9521,N_9530);
nor U9619 (N_9619,N_9485,N_9403);
xor U9620 (N_9620,N_9466,N_9476);
nand U9621 (N_9621,N_9545,N_9544);
or U9622 (N_9622,N_9540,N_9460);
and U9623 (N_9623,N_9560,N_9563);
nand U9624 (N_9624,N_9590,N_9524);
nand U9625 (N_9625,N_9452,N_9482);
and U9626 (N_9626,N_9578,N_9528);
or U9627 (N_9627,N_9444,N_9402);
nor U9628 (N_9628,N_9539,N_9475);
or U9629 (N_9629,N_9443,N_9411);
nand U9630 (N_9630,N_9419,N_9529);
and U9631 (N_9631,N_9410,N_9598);
and U9632 (N_9632,N_9518,N_9494);
nand U9633 (N_9633,N_9454,N_9478);
and U9634 (N_9634,N_9449,N_9570);
or U9635 (N_9635,N_9536,N_9502);
nand U9636 (N_9636,N_9501,N_9512);
xor U9637 (N_9637,N_9465,N_9555);
and U9638 (N_9638,N_9581,N_9514);
or U9639 (N_9639,N_9447,N_9591);
nor U9640 (N_9640,N_9562,N_9489);
or U9641 (N_9641,N_9520,N_9543);
nor U9642 (N_9642,N_9455,N_9445);
nor U9643 (N_9643,N_9437,N_9597);
nor U9644 (N_9644,N_9505,N_9586);
and U9645 (N_9645,N_9422,N_9468);
or U9646 (N_9646,N_9569,N_9469);
nand U9647 (N_9647,N_9541,N_9432);
and U9648 (N_9648,N_9434,N_9474);
nor U9649 (N_9649,N_9527,N_9440);
nand U9650 (N_9650,N_9479,N_9480);
and U9651 (N_9651,N_9532,N_9593);
or U9652 (N_9652,N_9458,N_9439);
or U9653 (N_9653,N_9451,N_9492);
nor U9654 (N_9654,N_9418,N_9472);
and U9655 (N_9655,N_9580,N_9457);
nor U9656 (N_9656,N_9497,N_9533);
nand U9657 (N_9657,N_9441,N_9424);
nand U9658 (N_9658,N_9408,N_9421);
and U9659 (N_9659,N_9406,N_9401);
or U9660 (N_9660,N_9429,N_9573);
nor U9661 (N_9661,N_9525,N_9596);
and U9662 (N_9662,N_9509,N_9577);
or U9663 (N_9663,N_9517,N_9436);
and U9664 (N_9664,N_9484,N_9446);
or U9665 (N_9665,N_9409,N_9516);
or U9666 (N_9666,N_9572,N_9498);
nor U9667 (N_9667,N_9416,N_9428);
or U9668 (N_9668,N_9552,N_9442);
nor U9669 (N_9669,N_9537,N_9549);
nand U9670 (N_9670,N_9574,N_9483);
nand U9671 (N_9671,N_9515,N_9456);
nand U9672 (N_9672,N_9535,N_9558);
xnor U9673 (N_9673,N_9556,N_9522);
nand U9674 (N_9674,N_9415,N_9417);
or U9675 (N_9675,N_9551,N_9500);
nand U9676 (N_9676,N_9420,N_9414);
nor U9677 (N_9677,N_9453,N_9490);
nand U9678 (N_9678,N_9459,N_9567);
and U9679 (N_9679,N_9550,N_9557);
or U9680 (N_9680,N_9496,N_9488);
nor U9681 (N_9681,N_9404,N_9473);
and U9682 (N_9682,N_9584,N_9564);
nand U9683 (N_9683,N_9511,N_9554);
or U9684 (N_9684,N_9575,N_9463);
nand U9685 (N_9685,N_9548,N_9531);
and U9686 (N_9686,N_9504,N_9433);
nor U9687 (N_9687,N_9538,N_9542);
nor U9688 (N_9688,N_9588,N_9438);
and U9689 (N_9689,N_9499,N_9431);
nor U9690 (N_9690,N_9471,N_9599);
xor U9691 (N_9691,N_9513,N_9462);
nor U9692 (N_9692,N_9587,N_9495);
or U9693 (N_9693,N_9400,N_9425);
nand U9694 (N_9694,N_9582,N_9592);
nand U9695 (N_9695,N_9519,N_9547);
or U9696 (N_9696,N_9594,N_9487);
or U9697 (N_9697,N_9559,N_9470);
nand U9698 (N_9698,N_9523,N_9507);
nand U9699 (N_9699,N_9503,N_9450);
nand U9700 (N_9700,N_9485,N_9454);
and U9701 (N_9701,N_9445,N_9599);
nor U9702 (N_9702,N_9539,N_9418);
nand U9703 (N_9703,N_9423,N_9584);
or U9704 (N_9704,N_9470,N_9595);
nand U9705 (N_9705,N_9469,N_9456);
xor U9706 (N_9706,N_9536,N_9455);
nand U9707 (N_9707,N_9515,N_9570);
nor U9708 (N_9708,N_9500,N_9411);
or U9709 (N_9709,N_9506,N_9407);
and U9710 (N_9710,N_9573,N_9458);
nor U9711 (N_9711,N_9564,N_9469);
or U9712 (N_9712,N_9452,N_9566);
xnor U9713 (N_9713,N_9563,N_9445);
nand U9714 (N_9714,N_9594,N_9506);
nor U9715 (N_9715,N_9527,N_9406);
nand U9716 (N_9716,N_9512,N_9529);
and U9717 (N_9717,N_9495,N_9446);
or U9718 (N_9718,N_9400,N_9411);
nor U9719 (N_9719,N_9432,N_9487);
nand U9720 (N_9720,N_9400,N_9532);
or U9721 (N_9721,N_9560,N_9413);
nor U9722 (N_9722,N_9438,N_9518);
xor U9723 (N_9723,N_9553,N_9454);
or U9724 (N_9724,N_9421,N_9539);
and U9725 (N_9725,N_9425,N_9426);
and U9726 (N_9726,N_9547,N_9506);
or U9727 (N_9727,N_9421,N_9417);
xor U9728 (N_9728,N_9470,N_9410);
nor U9729 (N_9729,N_9513,N_9445);
or U9730 (N_9730,N_9563,N_9565);
nor U9731 (N_9731,N_9546,N_9524);
or U9732 (N_9732,N_9592,N_9544);
nor U9733 (N_9733,N_9500,N_9420);
nor U9734 (N_9734,N_9594,N_9437);
or U9735 (N_9735,N_9410,N_9558);
nor U9736 (N_9736,N_9549,N_9530);
and U9737 (N_9737,N_9404,N_9553);
or U9738 (N_9738,N_9578,N_9431);
or U9739 (N_9739,N_9502,N_9501);
or U9740 (N_9740,N_9421,N_9452);
xor U9741 (N_9741,N_9428,N_9465);
nor U9742 (N_9742,N_9440,N_9501);
and U9743 (N_9743,N_9544,N_9464);
and U9744 (N_9744,N_9437,N_9503);
nand U9745 (N_9745,N_9524,N_9530);
or U9746 (N_9746,N_9493,N_9480);
or U9747 (N_9747,N_9561,N_9563);
or U9748 (N_9748,N_9424,N_9532);
or U9749 (N_9749,N_9505,N_9464);
or U9750 (N_9750,N_9455,N_9562);
nand U9751 (N_9751,N_9553,N_9595);
and U9752 (N_9752,N_9550,N_9455);
nor U9753 (N_9753,N_9477,N_9535);
nor U9754 (N_9754,N_9485,N_9545);
or U9755 (N_9755,N_9534,N_9402);
or U9756 (N_9756,N_9455,N_9545);
xnor U9757 (N_9757,N_9481,N_9441);
nor U9758 (N_9758,N_9518,N_9461);
nor U9759 (N_9759,N_9450,N_9525);
or U9760 (N_9760,N_9547,N_9403);
or U9761 (N_9761,N_9404,N_9440);
xnor U9762 (N_9762,N_9450,N_9452);
or U9763 (N_9763,N_9510,N_9577);
xor U9764 (N_9764,N_9402,N_9416);
nor U9765 (N_9765,N_9572,N_9598);
or U9766 (N_9766,N_9599,N_9561);
or U9767 (N_9767,N_9556,N_9500);
and U9768 (N_9768,N_9515,N_9433);
xnor U9769 (N_9769,N_9594,N_9449);
nor U9770 (N_9770,N_9537,N_9520);
and U9771 (N_9771,N_9459,N_9535);
or U9772 (N_9772,N_9463,N_9550);
xor U9773 (N_9773,N_9546,N_9499);
nor U9774 (N_9774,N_9514,N_9477);
or U9775 (N_9775,N_9585,N_9429);
nand U9776 (N_9776,N_9457,N_9419);
xnor U9777 (N_9777,N_9530,N_9480);
and U9778 (N_9778,N_9560,N_9503);
or U9779 (N_9779,N_9430,N_9549);
xnor U9780 (N_9780,N_9455,N_9496);
and U9781 (N_9781,N_9419,N_9525);
nand U9782 (N_9782,N_9511,N_9597);
xnor U9783 (N_9783,N_9433,N_9537);
or U9784 (N_9784,N_9473,N_9447);
and U9785 (N_9785,N_9529,N_9504);
nand U9786 (N_9786,N_9475,N_9402);
nand U9787 (N_9787,N_9402,N_9449);
nand U9788 (N_9788,N_9565,N_9541);
xor U9789 (N_9789,N_9436,N_9526);
and U9790 (N_9790,N_9489,N_9539);
nand U9791 (N_9791,N_9437,N_9556);
or U9792 (N_9792,N_9422,N_9580);
nand U9793 (N_9793,N_9507,N_9583);
nand U9794 (N_9794,N_9463,N_9435);
nor U9795 (N_9795,N_9497,N_9506);
xor U9796 (N_9796,N_9407,N_9489);
nor U9797 (N_9797,N_9580,N_9590);
nor U9798 (N_9798,N_9485,N_9590);
nand U9799 (N_9799,N_9450,N_9428);
and U9800 (N_9800,N_9749,N_9787);
nand U9801 (N_9801,N_9768,N_9786);
nor U9802 (N_9802,N_9718,N_9777);
or U9803 (N_9803,N_9646,N_9674);
and U9804 (N_9804,N_9626,N_9637);
and U9805 (N_9805,N_9723,N_9776);
nor U9806 (N_9806,N_9794,N_9700);
and U9807 (N_9807,N_9650,N_9672);
and U9808 (N_9808,N_9609,N_9633);
nand U9809 (N_9809,N_9616,N_9704);
and U9810 (N_9810,N_9601,N_9632);
nor U9811 (N_9811,N_9654,N_9613);
nor U9812 (N_9812,N_9683,N_9722);
xnor U9813 (N_9813,N_9756,N_9747);
or U9814 (N_9814,N_9769,N_9717);
nand U9815 (N_9815,N_9778,N_9746);
or U9816 (N_9816,N_9640,N_9635);
nor U9817 (N_9817,N_9793,N_9663);
xnor U9818 (N_9818,N_9711,N_9682);
nor U9819 (N_9819,N_9623,N_9799);
xnor U9820 (N_9820,N_9785,N_9686);
or U9821 (N_9821,N_9779,N_9752);
and U9822 (N_9822,N_9606,N_9741);
xor U9823 (N_9823,N_9617,N_9610);
xor U9824 (N_9824,N_9630,N_9761);
or U9825 (N_9825,N_9784,N_9668);
and U9826 (N_9826,N_9659,N_9662);
nand U9827 (N_9827,N_9618,N_9671);
and U9828 (N_9828,N_9602,N_9677);
or U9829 (N_9829,N_9636,N_9760);
nand U9830 (N_9830,N_9763,N_9762);
nand U9831 (N_9831,N_9608,N_9667);
nand U9832 (N_9832,N_9754,N_9745);
nor U9833 (N_9833,N_9721,N_9669);
nor U9834 (N_9834,N_9713,N_9702);
and U9835 (N_9835,N_9692,N_9736);
and U9836 (N_9836,N_9706,N_9724);
and U9837 (N_9837,N_9797,N_9649);
nand U9838 (N_9838,N_9730,N_9791);
nand U9839 (N_9839,N_9684,N_9651);
or U9840 (N_9840,N_9679,N_9638);
and U9841 (N_9841,N_9751,N_9789);
or U9842 (N_9842,N_9703,N_9603);
and U9843 (N_9843,N_9664,N_9676);
and U9844 (N_9844,N_9631,N_9775);
or U9845 (N_9845,N_9658,N_9643);
xor U9846 (N_9846,N_9710,N_9782);
and U9847 (N_9847,N_9641,N_9687);
nand U9848 (N_9848,N_9605,N_9712);
nor U9849 (N_9849,N_9781,N_9726);
and U9850 (N_9850,N_9689,N_9690);
xnor U9851 (N_9851,N_9696,N_9657);
nand U9852 (N_9852,N_9620,N_9621);
nor U9853 (N_9853,N_9691,N_9733);
nor U9854 (N_9854,N_9701,N_9666);
nand U9855 (N_9855,N_9728,N_9656);
nor U9856 (N_9856,N_9628,N_9739);
nor U9857 (N_9857,N_9719,N_9709);
and U9858 (N_9858,N_9788,N_9773);
or U9859 (N_9859,N_9645,N_9619);
nand U9860 (N_9860,N_9744,N_9735);
nor U9861 (N_9861,N_9665,N_9795);
or U9862 (N_9862,N_9660,N_9648);
nor U9863 (N_9863,N_9790,N_9653);
nand U9864 (N_9864,N_9715,N_9771);
or U9865 (N_9865,N_9738,N_9681);
and U9866 (N_9866,N_9767,N_9698);
xnor U9867 (N_9867,N_9780,N_9743);
xnor U9868 (N_9868,N_9720,N_9731);
and U9869 (N_9869,N_9644,N_9624);
or U9870 (N_9870,N_9629,N_9675);
or U9871 (N_9871,N_9614,N_9707);
and U9872 (N_9872,N_9611,N_9766);
nor U9873 (N_9873,N_9725,N_9764);
and U9874 (N_9874,N_9647,N_9607);
nor U9875 (N_9875,N_9688,N_9655);
nor U9876 (N_9876,N_9634,N_9625);
or U9877 (N_9877,N_9772,N_9661);
nand U9878 (N_9878,N_9798,N_9705);
nor U9879 (N_9879,N_9783,N_9770);
nor U9880 (N_9880,N_9695,N_9753);
nor U9881 (N_9881,N_9796,N_9729);
nor U9882 (N_9882,N_9642,N_9680);
xor U9883 (N_9883,N_9600,N_9615);
nor U9884 (N_9884,N_9758,N_9697);
or U9885 (N_9885,N_9732,N_9714);
and U9886 (N_9886,N_9716,N_9694);
nand U9887 (N_9887,N_9774,N_9612);
nor U9888 (N_9888,N_9652,N_9670);
nor U9889 (N_9889,N_9748,N_9693);
or U9890 (N_9890,N_9742,N_9737);
nor U9891 (N_9891,N_9740,N_9627);
nor U9892 (N_9892,N_9792,N_9750);
or U9893 (N_9893,N_9755,N_9708);
nor U9894 (N_9894,N_9622,N_9699);
nand U9895 (N_9895,N_9727,N_9734);
and U9896 (N_9896,N_9673,N_9639);
nor U9897 (N_9897,N_9678,N_9685);
nand U9898 (N_9898,N_9759,N_9757);
and U9899 (N_9899,N_9604,N_9765);
nand U9900 (N_9900,N_9694,N_9723);
nand U9901 (N_9901,N_9733,N_9718);
xnor U9902 (N_9902,N_9668,N_9617);
or U9903 (N_9903,N_9681,N_9754);
xnor U9904 (N_9904,N_9601,N_9776);
and U9905 (N_9905,N_9792,N_9797);
xnor U9906 (N_9906,N_9741,N_9686);
and U9907 (N_9907,N_9771,N_9704);
xnor U9908 (N_9908,N_9695,N_9670);
nor U9909 (N_9909,N_9775,N_9639);
and U9910 (N_9910,N_9685,N_9657);
nor U9911 (N_9911,N_9651,N_9725);
nor U9912 (N_9912,N_9667,N_9780);
and U9913 (N_9913,N_9644,N_9770);
or U9914 (N_9914,N_9605,N_9781);
or U9915 (N_9915,N_9775,N_9664);
nand U9916 (N_9916,N_9682,N_9742);
and U9917 (N_9917,N_9764,N_9752);
nor U9918 (N_9918,N_9692,N_9668);
or U9919 (N_9919,N_9789,N_9602);
xnor U9920 (N_9920,N_9677,N_9744);
nand U9921 (N_9921,N_9770,N_9656);
nand U9922 (N_9922,N_9631,N_9788);
and U9923 (N_9923,N_9669,N_9723);
or U9924 (N_9924,N_9795,N_9650);
nand U9925 (N_9925,N_9799,N_9750);
nor U9926 (N_9926,N_9623,N_9614);
or U9927 (N_9927,N_9708,N_9644);
nor U9928 (N_9928,N_9752,N_9735);
nand U9929 (N_9929,N_9706,N_9611);
and U9930 (N_9930,N_9611,N_9642);
nand U9931 (N_9931,N_9635,N_9755);
or U9932 (N_9932,N_9796,N_9704);
nor U9933 (N_9933,N_9786,N_9715);
nor U9934 (N_9934,N_9664,N_9730);
or U9935 (N_9935,N_9666,N_9642);
or U9936 (N_9936,N_9716,N_9611);
nand U9937 (N_9937,N_9674,N_9641);
and U9938 (N_9938,N_9708,N_9790);
or U9939 (N_9939,N_9748,N_9794);
xnor U9940 (N_9940,N_9752,N_9713);
or U9941 (N_9941,N_9750,N_9705);
or U9942 (N_9942,N_9764,N_9661);
nand U9943 (N_9943,N_9746,N_9706);
or U9944 (N_9944,N_9775,N_9643);
and U9945 (N_9945,N_9662,N_9673);
nor U9946 (N_9946,N_9697,N_9669);
and U9947 (N_9947,N_9656,N_9776);
nand U9948 (N_9948,N_9650,N_9716);
nand U9949 (N_9949,N_9694,N_9617);
or U9950 (N_9950,N_9778,N_9701);
and U9951 (N_9951,N_9610,N_9673);
and U9952 (N_9952,N_9625,N_9612);
nand U9953 (N_9953,N_9608,N_9642);
xnor U9954 (N_9954,N_9743,N_9714);
and U9955 (N_9955,N_9679,N_9613);
and U9956 (N_9956,N_9784,N_9741);
and U9957 (N_9957,N_9700,N_9777);
and U9958 (N_9958,N_9605,N_9623);
xor U9959 (N_9959,N_9619,N_9654);
and U9960 (N_9960,N_9644,N_9709);
nor U9961 (N_9961,N_9681,N_9713);
nand U9962 (N_9962,N_9721,N_9728);
nor U9963 (N_9963,N_9797,N_9772);
nand U9964 (N_9964,N_9721,N_9763);
xnor U9965 (N_9965,N_9730,N_9737);
nor U9966 (N_9966,N_9615,N_9663);
and U9967 (N_9967,N_9712,N_9678);
nor U9968 (N_9968,N_9790,N_9764);
and U9969 (N_9969,N_9775,N_9767);
nand U9970 (N_9970,N_9701,N_9703);
nor U9971 (N_9971,N_9772,N_9738);
nor U9972 (N_9972,N_9703,N_9678);
xnor U9973 (N_9973,N_9614,N_9741);
nor U9974 (N_9974,N_9742,N_9798);
or U9975 (N_9975,N_9659,N_9693);
xor U9976 (N_9976,N_9635,N_9617);
and U9977 (N_9977,N_9790,N_9792);
and U9978 (N_9978,N_9672,N_9724);
nor U9979 (N_9979,N_9667,N_9635);
nor U9980 (N_9980,N_9735,N_9696);
or U9981 (N_9981,N_9778,N_9762);
and U9982 (N_9982,N_9653,N_9620);
nand U9983 (N_9983,N_9764,N_9758);
xor U9984 (N_9984,N_9768,N_9799);
nand U9985 (N_9985,N_9654,N_9796);
nand U9986 (N_9986,N_9625,N_9606);
nor U9987 (N_9987,N_9744,N_9676);
nand U9988 (N_9988,N_9619,N_9673);
and U9989 (N_9989,N_9608,N_9665);
and U9990 (N_9990,N_9786,N_9746);
or U9991 (N_9991,N_9663,N_9738);
nor U9992 (N_9992,N_9792,N_9713);
nand U9993 (N_9993,N_9728,N_9667);
nor U9994 (N_9994,N_9786,N_9652);
xnor U9995 (N_9995,N_9661,N_9714);
xnor U9996 (N_9996,N_9748,N_9702);
nor U9997 (N_9997,N_9646,N_9687);
nand U9998 (N_9998,N_9621,N_9756);
and U9999 (N_9999,N_9769,N_9613);
or U10000 (N_10000,N_9862,N_9981);
nand U10001 (N_10001,N_9945,N_9993);
or U10002 (N_10002,N_9974,N_9806);
nor U10003 (N_10003,N_9984,N_9911);
and U10004 (N_10004,N_9858,N_9834);
xor U10005 (N_10005,N_9953,N_9920);
nor U10006 (N_10006,N_9961,N_9941);
nand U10007 (N_10007,N_9899,N_9983);
xnor U10008 (N_10008,N_9880,N_9876);
nand U10009 (N_10009,N_9817,N_9969);
nand U10010 (N_10010,N_9922,N_9937);
or U10011 (N_10011,N_9927,N_9923);
and U10012 (N_10012,N_9943,N_9888);
nor U10013 (N_10013,N_9979,N_9833);
and U10014 (N_10014,N_9925,N_9869);
and U10015 (N_10015,N_9976,N_9843);
nand U10016 (N_10016,N_9801,N_9818);
and U10017 (N_10017,N_9828,N_9965);
nand U10018 (N_10018,N_9950,N_9855);
and U10019 (N_10019,N_9936,N_9972);
xor U10020 (N_10020,N_9990,N_9831);
nor U10021 (N_10021,N_9918,N_9816);
nand U10022 (N_10022,N_9852,N_9890);
xor U10023 (N_10023,N_9842,N_9939);
or U10024 (N_10024,N_9924,N_9998);
nand U10025 (N_10025,N_9865,N_9975);
nand U10026 (N_10026,N_9809,N_9883);
or U10027 (N_10027,N_9882,N_9934);
xnor U10028 (N_10028,N_9861,N_9970);
or U10029 (N_10029,N_9854,N_9906);
nor U10030 (N_10030,N_9938,N_9803);
or U10031 (N_10031,N_9824,N_9957);
nor U10032 (N_10032,N_9859,N_9966);
nand U10033 (N_10033,N_9850,N_9994);
xnor U10034 (N_10034,N_9832,N_9905);
xor U10035 (N_10035,N_9825,N_9992);
nor U10036 (N_10036,N_9830,N_9837);
or U10037 (N_10037,N_9914,N_9968);
or U10038 (N_10038,N_9985,N_9933);
and U10039 (N_10039,N_9962,N_9844);
nand U10040 (N_10040,N_9813,N_9947);
or U10041 (N_10041,N_9804,N_9967);
and U10042 (N_10042,N_9912,N_9805);
or U10043 (N_10043,N_9874,N_9935);
or U10044 (N_10044,N_9978,N_9900);
nor U10045 (N_10045,N_9903,N_9839);
nand U10046 (N_10046,N_9864,N_9949);
or U10047 (N_10047,N_9897,N_9988);
nand U10048 (N_10048,N_9848,N_9849);
nand U10049 (N_10049,N_9860,N_9977);
nand U10050 (N_10050,N_9960,N_9995);
and U10051 (N_10051,N_9986,N_9836);
xor U10052 (N_10052,N_9889,N_9958);
and U10053 (N_10053,N_9971,N_9902);
xor U10054 (N_10054,N_9991,N_9893);
nor U10055 (N_10055,N_9931,N_9908);
and U10056 (N_10056,N_9867,N_9901);
nand U10057 (N_10057,N_9808,N_9815);
and U10058 (N_10058,N_9907,N_9819);
nand U10059 (N_10059,N_9853,N_9851);
or U10060 (N_10060,N_9807,N_9870);
nor U10061 (N_10061,N_9951,N_9847);
nor U10062 (N_10062,N_9946,N_9871);
nor U10063 (N_10063,N_9826,N_9838);
xnor U10064 (N_10064,N_9845,N_9840);
or U10065 (N_10065,N_9878,N_9915);
nand U10066 (N_10066,N_9980,N_9963);
nor U10067 (N_10067,N_9875,N_9898);
xnor U10068 (N_10068,N_9812,N_9948);
xor U10069 (N_10069,N_9891,N_9954);
and U10070 (N_10070,N_9802,N_9884);
or U10071 (N_10071,N_9823,N_9822);
nor U10072 (N_10072,N_9944,N_9879);
nor U10073 (N_10073,N_9863,N_9896);
or U10074 (N_10074,N_9873,N_9810);
nand U10075 (N_10075,N_9904,N_9895);
nor U10076 (N_10076,N_9913,N_9930);
or U10077 (N_10077,N_9926,N_9917);
nor U10078 (N_10078,N_9814,N_9866);
or U10079 (N_10079,N_9959,N_9868);
or U10080 (N_10080,N_9885,N_9919);
xnor U10081 (N_10081,N_9921,N_9856);
nand U10082 (N_10082,N_9997,N_9987);
nor U10083 (N_10083,N_9820,N_9929);
nor U10084 (N_10084,N_9955,N_9964);
or U10085 (N_10085,N_9800,N_9989);
or U10086 (N_10086,N_9846,N_9857);
or U10087 (N_10087,N_9881,N_9877);
and U10088 (N_10088,N_9829,N_9886);
or U10089 (N_10089,N_9872,N_9999);
or U10090 (N_10090,N_9916,N_9841);
nand U10091 (N_10091,N_9996,N_9811);
nor U10092 (N_10092,N_9982,N_9932);
and U10093 (N_10093,N_9835,N_9894);
or U10094 (N_10094,N_9928,N_9973);
nand U10095 (N_10095,N_9887,N_9892);
or U10096 (N_10096,N_9952,N_9909);
nor U10097 (N_10097,N_9827,N_9910);
nor U10098 (N_10098,N_9956,N_9942);
nor U10099 (N_10099,N_9940,N_9821);
nand U10100 (N_10100,N_9906,N_9846);
nand U10101 (N_10101,N_9996,N_9892);
nor U10102 (N_10102,N_9825,N_9896);
and U10103 (N_10103,N_9862,N_9985);
nand U10104 (N_10104,N_9998,N_9820);
nand U10105 (N_10105,N_9942,N_9909);
or U10106 (N_10106,N_9868,N_9982);
or U10107 (N_10107,N_9905,N_9861);
nor U10108 (N_10108,N_9878,N_9828);
nand U10109 (N_10109,N_9857,N_9949);
nand U10110 (N_10110,N_9960,N_9828);
and U10111 (N_10111,N_9819,N_9832);
or U10112 (N_10112,N_9802,N_9828);
or U10113 (N_10113,N_9974,N_9846);
and U10114 (N_10114,N_9980,N_9810);
or U10115 (N_10115,N_9812,N_9805);
nand U10116 (N_10116,N_9955,N_9912);
nor U10117 (N_10117,N_9867,N_9934);
nand U10118 (N_10118,N_9975,N_9806);
and U10119 (N_10119,N_9935,N_9816);
nor U10120 (N_10120,N_9856,N_9868);
or U10121 (N_10121,N_9996,N_9886);
and U10122 (N_10122,N_9980,N_9931);
xnor U10123 (N_10123,N_9877,N_9845);
and U10124 (N_10124,N_9883,N_9864);
and U10125 (N_10125,N_9849,N_9935);
or U10126 (N_10126,N_9827,N_9912);
and U10127 (N_10127,N_9933,N_9991);
nor U10128 (N_10128,N_9830,N_9934);
or U10129 (N_10129,N_9954,N_9884);
or U10130 (N_10130,N_9960,N_9809);
or U10131 (N_10131,N_9897,N_9977);
and U10132 (N_10132,N_9836,N_9817);
nor U10133 (N_10133,N_9936,N_9965);
or U10134 (N_10134,N_9881,N_9931);
or U10135 (N_10135,N_9808,N_9875);
nand U10136 (N_10136,N_9982,N_9928);
nor U10137 (N_10137,N_9980,N_9968);
nor U10138 (N_10138,N_9983,N_9965);
nand U10139 (N_10139,N_9867,N_9893);
xnor U10140 (N_10140,N_9958,N_9978);
and U10141 (N_10141,N_9867,N_9971);
nor U10142 (N_10142,N_9968,N_9840);
nand U10143 (N_10143,N_9815,N_9911);
nand U10144 (N_10144,N_9890,N_9867);
nand U10145 (N_10145,N_9950,N_9910);
and U10146 (N_10146,N_9944,N_9996);
and U10147 (N_10147,N_9880,N_9809);
or U10148 (N_10148,N_9958,N_9909);
nand U10149 (N_10149,N_9881,N_9826);
nor U10150 (N_10150,N_9885,N_9824);
or U10151 (N_10151,N_9941,N_9931);
and U10152 (N_10152,N_9852,N_9940);
nor U10153 (N_10153,N_9868,N_9955);
or U10154 (N_10154,N_9852,N_9904);
and U10155 (N_10155,N_9804,N_9940);
nor U10156 (N_10156,N_9950,N_9936);
or U10157 (N_10157,N_9991,N_9941);
nand U10158 (N_10158,N_9934,N_9989);
and U10159 (N_10159,N_9863,N_9928);
nor U10160 (N_10160,N_9812,N_9825);
or U10161 (N_10161,N_9830,N_9859);
or U10162 (N_10162,N_9910,N_9994);
and U10163 (N_10163,N_9899,N_9912);
and U10164 (N_10164,N_9932,N_9879);
nor U10165 (N_10165,N_9957,N_9805);
nand U10166 (N_10166,N_9819,N_9893);
nand U10167 (N_10167,N_9929,N_9998);
and U10168 (N_10168,N_9805,N_9904);
nand U10169 (N_10169,N_9894,N_9922);
or U10170 (N_10170,N_9949,N_9980);
or U10171 (N_10171,N_9867,N_9826);
xor U10172 (N_10172,N_9819,N_9910);
nand U10173 (N_10173,N_9818,N_9844);
and U10174 (N_10174,N_9906,N_9948);
and U10175 (N_10175,N_9811,N_9810);
or U10176 (N_10176,N_9820,N_9972);
xnor U10177 (N_10177,N_9921,N_9989);
and U10178 (N_10178,N_9898,N_9890);
or U10179 (N_10179,N_9946,N_9939);
nor U10180 (N_10180,N_9813,N_9814);
nand U10181 (N_10181,N_9824,N_9918);
xor U10182 (N_10182,N_9847,N_9870);
nand U10183 (N_10183,N_9962,N_9922);
nand U10184 (N_10184,N_9872,N_9809);
nor U10185 (N_10185,N_9801,N_9889);
or U10186 (N_10186,N_9972,N_9858);
or U10187 (N_10187,N_9802,N_9890);
and U10188 (N_10188,N_9981,N_9827);
and U10189 (N_10189,N_9851,N_9889);
and U10190 (N_10190,N_9959,N_9915);
nand U10191 (N_10191,N_9997,N_9955);
nand U10192 (N_10192,N_9951,N_9948);
nand U10193 (N_10193,N_9854,N_9813);
nor U10194 (N_10194,N_9973,N_9858);
nor U10195 (N_10195,N_9924,N_9989);
xnor U10196 (N_10196,N_9980,N_9905);
nor U10197 (N_10197,N_9889,N_9915);
or U10198 (N_10198,N_9881,N_9920);
or U10199 (N_10199,N_9868,N_9976);
nor U10200 (N_10200,N_10109,N_10159);
nor U10201 (N_10201,N_10171,N_10104);
and U10202 (N_10202,N_10108,N_10166);
or U10203 (N_10203,N_10001,N_10184);
or U10204 (N_10204,N_10066,N_10127);
or U10205 (N_10205,N_10071,N_10052);
and U10206 (N_10206,N_10048,N_10189);
nand U10207 (N_10207,N_10086,N_10140);
xnor U10208 (N_10208,N_10195,N_10000);
and U10209 (N_10209,N_10064,N_10050);
nand U10210 (N_10210,N_10042,N_10096);
or U10211 (N_10211,N_10107,N_10095);
and U10212 (N_10212,N_10017,N_10158);
nand U10213 (N_10213,N_10046,N_10136);
and U10214 (N_10214,N_10130,N_10010);
or U10215 (N_10215,N_10105,N_10074);
nand U10216 (N_10216,N_10162,N_10067);
xor U10217 (N_10217,N_10072,N_10125);
or U10218 (N_10218,N_10009,N_10097);
nor U10219 (N_10219,N_10045,N_10060);
or U10220 (N_10220,N_10079,N_10141);
nor U10221 (N_10221,N_10178,N_10118);
nand U10222 (N_10222,N_10156,N_10008);
nand U10223 (N_10223,N_10021,N_10185);
nor U10224 (N_10224,N_10035,N_10179);
nand U10225 (N_10225,N_10006,N_10142);
or U10226 (N_10226,N_10055,N_10139);
xor U10227 (N_10227,N_10049,N_10034);
nor U10228 (N_10228,N_10092,N_10199);
or U10229 (N_10229,N_10033,N_10085);
nor U10230 (N_10230,N_10084,N_10038);
nand U10231 (N_10231,N_10183,N_10099);
and U10232 (N_10232,N_10011,N_10093);
and U10233 (N_10233,N_10015,N_10146);
nand U10234 (N_10234,N_10098,N_10082);
nand U10235 (N_10235,N_10116,N_10012);
or U10236 (N_10236,N_10163,N_10115);
or U10237 (N_10237,N_10083,N_10110);
nand U10238 (N_10238,N_10040,N_10028);
nand U10239 (N_10239,N_10090,N_10056);
nand U10240 (N_10240,N_10023,N_10111);
nor U10241 (N_10241,N_10182,N_10148);
and U10242 (N_10242,N_10054,N_10153);
nor U10243 (N_10243,N_10143,N_10133);
or U10244 (N_10244,N_10106,N_10170);
and U10245 (N_10245,N_10131,N_10165);
nand U10246 (N_10246,N_10102,N_10036);
and U10247 (N_10247,N_10191,N_10144);
and U10248 (N_10248,N_10103,N_10168);
nand U10249 (N_10249,N_10177,N_10147);
nand U10250 (N_10250,N_10117,N_10152);
and U10251 (N_10251,N_10100,N_10120);
or U10252 (N_10252,N_10194,N_10004);
nand U10253 (N_10253,N_10018,N_10081);
and U10254 (N_10254,N_10078,N_10047);
nor U10255 (N_10255,N_10197,N_10062);
nor U10256 (N_10256,N_10080,N_10073);
nor U10257 (N_10257,N_10128,N_10173);
and U10258 (N_10258,N_10186,N_10167);
nand U10259 (N_10259,N_10174,N_10029);
and U10260 (N_10260,N_10007,N_10016);
and U10261 (N_10261,N_10119,N_10039);
xnor U10262 (N_10262,N_10161,N_10031);
or U10263 (N_10263,N_10134,N_10058);
or U10264 (N_10264,N_10091,N_10005);
nor U10265 (N_10265,N_10043,N_10041);
nor U10266 (N_10266,N_10188,N_10070);
and U10267 (N_10267,N_10063,N_10175);
or U10268 (N_10268,N_10114,N_10172);
or U10269 (N_10269,N_10138,N_10187);
nand U10270 (N_10270,N_10003,N_10069);
nand U10271 (N_10271,N_10181,N_10160);
nor U10272 (N_10272,N_10024,N_10059);
or U10273 (N_10273,N_10124,N_10089);
nor U10274 (N_10274,N_10019,N_10087);
or U10275 (N_10275,N_10126,N_10014);
nor U10276 (N_10276,N_10025,N_10020);
nand U10277 (N_10277,N_10151,N_10137);
or U10278 (N_10278,N_10198,N_10002);
or U10279 (N_10279,N_10129,N_10061);
nor U10280 (N_10280,N_10057,N_10192);
or U10281 (N_10281,N_10154,N_10135);
and U10282 (N_10282,N_10026,N_10032);
nand U10283 (N_10283,N_10101,N_10196);
and U10284 (N_10284,N_10150,N_10027);
or U10285 (N_10285,N_10030,N_10053);
nand U10286 (N_10286,N_10180,N_10122);
or U10287 (N_10287,N_10132,N_10176);
nand U10288 (N_10288,N_10155,N_10121);
nand U10289 (N_10289,N_10075,N_10190);
or U10290 (N_10290,N_10088,N_10044);
nor U10291 (N_10291,N_10013,N_10068);
nor U10292 (N_10292,N_10164,N_10051);
or U10293 (N_10293,N_10094,N_10037);
nor U10294 (N_10294,N_10145,N_10193);
or U10295 (N_10295,N_10112,N_10022);
and U10296 (N_10296,N_10065,N_10077);
and U10297 (N_10297,N_10169,N_10157);
or U10298 (N_10298,N_10149,N_10113);
nor U10299 (N_10299,N_10123,N_10076);
nor U10300 (N_10300,N_10172,N_10002);
nand U10301 (N_10301,N_10168,N_10185);
nor U10302 (N_10302,N_10040,N_10144);
or U10303 (N_10303,N_10099,N_10194);
xnor U10304 (N_10304,N_10080,N_10052);
or U10305 (N_10305,N_10034,N_10197);
nor U10306 (N_10306,N_10186,N_10096);
nand U10307 (N_10307,N_10155,N_10007);
nand U10308 (N_10308,N_10122,N_10164);
nand U10309 (N_10309,N_10068,N_10124);
or U10310 (N_10310,N_10094,N_10087);
xnor U10311 (N_10311,N_10196,N_10177);
nand U10312 (N_10312,N_10117,N_10030);
and U10313 (N_10313,N_10053,N_10016);
nor U10314 (N_10314,N_10147,N_10126);
nor U10315 (N_10315,N_10068,N_10023);
or U10316 (N_10316,N_10051,N_10052);
or U10317 (N_10317,N_10008,N_10027);
nor U10318 (N_10318,N_10176,N_10192);
and U10319 (N_10319,N_10107,N_10063);
or U10320 (N_10320,N_10105,N_10164);
xnor U10321 (N_10321,N_10186,N_10043);
or U10322 (N_10322,N_10000,N_10153);
xnor U10323 (N_10323,N_10078,N_10093);
nand U10324 (N_10324,N_10092,N_10148);
nor U10325 (N_10325,N_10046,N_10027);
xor U10326 (N_10326,N_10064,N_10008);
and U10327 (N_10327,N_10096,N_10164);
or U10328 (N_10328,N_10091,N_10148);
xor U10329 (N_10329,N_10094,N_10181);
or U10330 (N_10330,N_10193,N_10132);
and U10331 (N_10331,N_10053,N_10087);
or U10332 (N_10332,N_10160,N_10037);
nor U10333 (N_10333,N_10041,N_10020);
or U10334 (N_10334,N_10029,N_10060);
nor U10335 (N_10335,N_10019,N_10038);
nor U10336 (N_10336,N_10096,N_10151);
and U10337 (N_10337,N_10149,N_10002);
nand U10338 (N_10338,N_10034,N_10118);
xnor U10339 (N_10339,N_10191,N_10008);
nor U10340 (N_10340,N_10118,N_10031);
and U10341 (N_10341,N_10095,N_10091);
or U10342 (N_10342,N_10050,N_10175);
nor U10343 (N_10343,N_10166,N_10146);
xor U10344 (N_10344,N_10022,N_10120);
xnor U10345 (N_10345,N_10112,N_10180);
nand U10346 (N_10346,N_10077,N_10034);
nor U10347 (N_10347,N_10185,N_10152);
or U10348 (N_10348,N_10078,N_10159);
nor U10349 (N_10349,N_10094,N_10149);
xor U10350 (N_10350,N_10147,N_10025);
nor U10351 (N_10351,N_10040,N_10115);
nor U10352 (N_10352,N_10062,N_10060);
and U10353 (N_10353,N_10070,N_10112);
and U10354 (N_10354,N_10153,N_10196);
xnor U10355 (N_10355,N_10197,N_10153);
or U10356 (N_10356,N_10081,N_10065);
nor U10357 (N_10357,N_10074,N_10011);
nor U10358 (N_10358,N_10163,N_10032);
or U10359 (N_10359,N_10180,N_10053);
and U10360 (N_10360,N_10002,N_10020);
nand U10361 (N_10361,N_10087,N_10130);
nand U10362 (N_10362,N_10029,N_10101);
and U10363 (N_10363,N_10014,N_10055);
and U10364 (N_10364,N_10106,N_10158);
nor U10365 (N_10365,N_10147,N_10190);
or U10366 (N_10366,N_10094,N_10046);
or U10367 (N_10367,N_10117,N_10114);
or U10368 (N_10368,N_10057,N_10194);
xnor U10369 (N_10369,N_10100,N_10181);
and U10370 (N_10370,N_10192,N_10009);
xnor U10371 (N_10371,N_10051,N_10188);
xor U10372 (N_10372,N_10064,N_10023);
xor U10373 (N_10373,N_10177,N_10041);
nor U10374 (N_10374,N_10153,N_10112);
nor U10375 (N_10375,N_10008,N_10176);
nor U10376 (N_10376,N_10106,N_10041);
xor U10377 (N_10377,N_10078,N_10112);
nor U10378 (N_10378,N_10128,N_10094);
or U10379 (N_10379,N_10146,N_10110);
xor U10380 (N_10380,N_10132,N_10161);
nand U10381 (N_10381,N_10057,N_10000);
and U10382 (N_10382,N_10124,N_10040);
nand U10383 (N_10383,N_10152,N_10008);
or U10384 (N_10384,N_10050,N_10097);
and U10385 (N_10385,N_10076,N_10178);
nor U10386 (N_10386,N_10075,N_10189);
and U10387 (N_10387,N_10073,N_10055);
or U10388 (N_10388,N_10091,N_10069);
nor U10389 (N_10389,N_10049,N_10033);
nand U10390 (N_10390,N_10020,N_10126);
nand U10391 (N_10391,N_10129,N_10078);
nor U10392 (N_10392,N_10103,N_10153);
nor U10393 (N_10393,N_10187,N_10010);
nand U10394 (N_10394,N_10046,N_10078);
nand U10395 (N_10395,N_10043,N_10141);
nand U10396 (N_10396,N_10142,N_10007);
nand U10397 (N_10397,N_10041,N_10067);
nand U10398 (N_10398,N_10081,N_10000);
xor U10399 (N_10399,N_10154,N_10038);
or U10400 (N_10400,N_10267,N_10248);
or U10401 (N_10401,N_10391,N_10276);
xor U10402 (N_10402,N_10324,N_10275);
nand U10403 (N_10403,N_10366,N_10369);
and U10404 (N_10404,N_10382,N_10330);
nor U10405 (N_10405,N_10339,N_10387);
nor U10406 (N_10406,N_10396,N_10301);
and U10407 (N_10407,N_10348,N_10380);
or U10408 (N_10408,N_10311,N_10341);
and U10409 (N_10409,N_10260,N_10328);
or U10410 (N_10410,N_10255,N_10247);
xnor U10411 (N_10411,N_10256,N_10266);
and U10412 (N_10412,N_10308,N_10385);
xnor U10413 (N_10413,N_10281,N_10338);
or U10414 (N_10414,N_10347,N_10390);
and U10415 (N_10415,N_10222,N_10240);
nor U10416 (N_10416,N_10329,N_10351);
or U10417 (N_10417,N_10395,N_10210);
or U10418 (N_10418,N_10272,N_10268);
nor U10419 (N_10419,N_10340,N_10350);
nor U10420 (N_10420,N_10249,N_10357);
and U10421 (N_10421,N_10213,N_10282);
xor U10422 (N_10422,N_10365,N_10394);
nand U10423 (N_10423,N_10321,N_10343);
and U10424 (N_10424,N_10283,N_10388);
or U10425 (N_10425,N_10274,N_10393);
xor U10426 (N_10426,N_10236,N_10383);
or U10427 (N_10427,N_10270,N_10367);
xor U10428 (N_10428,N_10207,N_10242);
nor U10429 (N_10429,N_10309,N_10314);
or U10430 (N_10430,N_10293,N_10320);
nor U10431 (N_10431,N_10335,N_10319);
or U10432 (N_10432,N_10299,N_10262);
nor U10433 (N_10433,N_10397,N_10305);
nand U10434 (N_10434,N_10306,N_10278);
and U10435 (N_10435,N_10368,N_10287);
nor U10436 (N_10436,N_10392,N_10244);
nand U10437 (N_10437,N_10219,N_10336);
xor U10438 (N_10438,N_10310,N_10300);
nor U10439 (N_10439,N_10334,N_10215);
nand U10440 (N_10440,N_10379,N_10239);
and U10441 (N_10441,N_10211,N_10326);
nor U10442 (N_10442,N_10398,N_10220);
or U10443 (N_10443,N_10234,N_10232);
and U10444 (N_10444,N_10245,N_10360);
and U10445 (N_10445,N_10307,N_10227);
nand U10446 (N_10446,N_10359,N_10363);
or U10447 (N_10447,N_10246,N_10323);
or U10448 (N_10448,N_10304,N_10374);
nor U10449 (N_10449,N_10203,N_10201);
or U10450 (N_10450,N_10288,N_10233);
xnor U10451 (N_10451,N_10370,N_10204);
nor U10452 (N_10452,N_10237,N_10251);
or U10453 (N_10453,N_10355,N_10231);
or U10454 (N_10454,N_10280,N_10228);
nand U10455 (N_10455,N_10250,N_10208);
nor U10456 (N_10456,N_10290,N_10223);
or U10457 (N_10457,N_10354,N_10361);
nand U10458 (N_10458,N_10342,N_10346);
nand U10459 (N_10459,N_10316,N_10322);
or U10460 (N_10460,N_10298,N_10271);
nor U10461 (N_10461,N_10284,N_10344);
nor U10462 (N_10462,N_10303,N_10263);
or U10463 (N_10463,N_10362,N_10285);
nand U10464 (N_10464,N_10241,N_10399);
nand U10465 (N_10465,N_10212,N_10206);
nand U10466 (N_10466,N_10381,N_10225);
nor U10467 (N_10467,N_10292,N_10315);
or U10468 (N_10468,N_10230,N_10345);
nand U10469 (N_10469,N_10318,N_10377);
or U10470 (N_10470,N_10337,N_10229);
xor U10471 (N_10471,N_10356,N_10226);
nor U10472 (N_10472,N_10235,N_10325);
or U10473 (N_10473,N_10218,N_10312);
or U10474 (N_10474,N_10375,N_10384);
or U10475 (N_10475,N_10202,N_10243);
or U10476 (N_10476,N_10261,N_10297);
and U10477 (N_10477,N_10286,N_10371);
nor U10478 (N_10478,N_10209,N_10252);
or U10479 (N_10479,N_10264,N_10205);
nor U10480 (N_10480,N_10352,N_10238);
nand U10481 (N_10481,N_10302,N_10378);
nand U10482 (N_10482,N_10389,N_10258);
xnor U10483 (N_10483,N_10224,N_10265);
nand U10484 (N_10484,N_10279,N_10200);
and U10485 (N_10485,N_10358,N_10259);
and U10486 (N_10486,N_10269,N_10254);
or U10487 (N_10487,N_10257,N_10289);
or U10488 (N_10488,N_10372,N_10295);
nand U10489 (N_10489,N_10353,N_10331);
nor U10490 (N_10490,N_10333,N_10294);
nand U10491 (N_10491,N_10317,N_10216);
or U10492 (N_10492,N_10291,N_10273);
or U10493 (N_10493,N_10214,N_10386);
nand U10494 (N_10494,N_10217,N_10327);
nor U10495 (N_10495,N_10221,N_10313);
nand U10496 (N_10496,N_10373,N_10253);
and U10497 (N_10497,N_10277,N_10364);
nand U10498 (N_10498,N_10349,N_10332);
nand U10499 (N_10499,N_10376,N_10296);
nand U10500 (N_10500,N_10294,N_10372);
xor U10501 (N_10501,N_10323,N_10354);
nand U10502 (N_10502,N_10309,N_10227);
nand U10503 (N_10503,N_10366,N_10260);
nand U10504 (N_10504,N_10322,N_10332);
and U10505 (N_10505,N_10264,N_10329);
and U10506 (N_10506,N_10389,N_10373);
xor U10507 (N_10507,N_10320,N_10233);
and U10508 (N_10508,N_10304,N_10301);
nand U10509 (N_10509,N_10310,N_10304);
nor U10510 (N_10510,N_10284,N_10307);
nor U10511 (N_10511,N_10250,N_10351);
nand U10512 (N_10512,N_10340,N_10239);
xnor U10513 (N_10513,N_10362,N_10234);
nor U10514 (N_10514,N_10363,N_10399);
or U10515 (N_10515,N_10349,N_10352);
or U10516 (N_10516,N_10340,N_10360);
nand U10517 (N_10517,N_10229,N_10233);
or U10518 (N_10518,N_10281,N_10332);
and U10519 (N_10519,N_10303,N_10396);
xnor U10520 (N_10520,N_10237,N_10364);
nand U10521 (N_10521,N_10355,N_10358);
nor U10522 (N_10522,N_10355,N_10356);
nand U10523 (N_10523,N_10204,N_10231);
xnor U10524 (N_10524,N_10351,N_10354);
nand U10525 (N_10525,N_10267,N_10374);
and U10526 (N_10526,N_10231,N_10289);
xnor U10527 (N_10527,N_10382,N_10395);
or U10528 (N_10528,N_10320,N_10272);
or U10529 (N_10529,N_10312,N_10318);
nand U10530 (N_10530,N_10212,N_10204);
and U10531 (N_10531,N_10293,N_10210);
nand U10532 (N_10532,N_10248,N_10229);
and U10533 (N_10533,N_10259,N_10337);
nor U10534 (N_10534,N_10337,N_10319);
nand U10535 (N_10535,N_10201,N_10367);
nor U10536 (N_10536,N_10292,N_10205);
or U10537 (N_10537,N_10214,N_10251);
nor U10538 (N_10538,N_10361,N_10394);
xnor U10539 (N_10539,N_10388,N_10325);
or U10540 (N_10540,N_10217,N_10203);
xor U10541 (N_10541,N_10321,N_10398);
or U10542 (N_10542,N_10293,N_10260);
nor U10543 (N_10543,N_10260,N_10237);
or U10544 (N_10544,N_10358,N_10271);
xnor U10545 (N_10545,N_10242,N_10270);
xnor U10546 (N_10546,N_10306,N_10201);
or U10547 (N_10547,N_10290,N_10341);
xnor U10548 (N_10548,N_10384,N_10292);
nor U10549 (N_10549,N_10373,N_10348);
and U10550 (N_10550,N_10282,N_10229);
or U10551 (N_10551,N_10234,N_10202);
or U10552 (N_10552,N_10328,N_10390);
nand U10553 (N_10553,N_10243,N_10340);
and U10554 (N_10554,N_10245,N_10332);
or U10555 (N_10555,N_10269,N_10323);
or U10556 (N_10556,N_10364,N_10361);
or U10557 (N_10557,N_10374,N_10226);
nand U10558 (N_10558,N_10382,N_10374);
nor U10559 (N_10559,N_10375,N_10238);
nor U10560 (N_10560,N_10250,N_10249);
nor U10561 (N_10561,N_10366,N_10230);
nand U10562 (N_10562,N_10321,N_10332);
nand U10563 (N_10563,N_10296,N_10262);
or U10564 (N_10564,N_10330,N_10246);
and U10565 (N_10565,N_10285,N_10365);
and U10566 (N_10566,N_10387,N_10274);
nand U10567 (N_10567,N_10354,N_10206);
nand U10568 (N_10568,N_10309,N_10251);
and U10569 (N_10569,N_10350,N_10314);
or U10570 (N_10570,N_10206,N_10337);
nor U10571 (N_10571,N_10245,N_10397);
nand U10572 (N_10572,N_10354,N_10287);
or U10573 (N_10573,N_10201,N_10381);
xnor U10574 (N_10574,N_10315,N_10233);
nand U10575 (N_10575,N_10215,N_10274);
nor U10576 (N_10576,N_10370,N_10348);
nand U10577 (N_10577,N_10351,N_10337);
nand U10578 (N_10578,N_10282,N_10301);
nand U10579 (N_10579,N_10329,N_10389);
or U10580 (N_10580,N_10362,N_10259);
xnor U10581 (N_10581,N_10200,N_10324);
nand U10582 (N_10582,N_10250,N_10278);
nor U10583 (N_10583,N_10269,N_10390);
nand U10584 (N_10584,N_10259,N_10379);
or U10585 (N_10585,N_10272,N_10369);
or U10586 (N_10586,N_10272,N_10359);
or U10587 (N_10587,N_10201,N_10332);
nor U10588 (N_10588,N_10311,N_10349);
xnor U10589 (N_10589,N_10322,N_10340);
nor U10590 (N_10590,N_10334,N_10274);
xor U10591 (N_10591,N_10229,N_10383);
nor U10592 (N_10592,N_10330,N_10387);
nand U10593 (N_10593,N_10361,N_10244);
nand U10594 (N_10594,N_10234,N_10228);
nor U10595 (N_10595,N_10232,N_10340);
nand U10596 (N_10596,N_10242,N_10217);
nor U10597 (N_10597,N_10340,N_10357);
xor U10598 (N_10598,N_10300,N_10322);
nand U10599 (N_10599,N_10204,N_10366);
or U10600 (N_10600,N_10538,N_10422);
or U10601 (N_10601,N_10565,N_10402);
nand U10602 (N_10602,N_10504,N_10427);
nand U10603 (N_10603,N_10542,N_10451);
or U10604 (N_10604,N_10516,N_10497);
nor U10605 (N_10605,N_10463,N_10597);
or U10606 (N_10606,N_10583,N_10540);
nor U10607 (N_10607,N_10466,N_10455);
nand U10608 (N_10608,N_10421,N_10522);
and U10609 (N_10609,N_10564,N_10493);
or U10610 (N_10610,N_10409,N_10444);
nand U10611 (N_10611,N_10595,N_10535);
and U10612 (N_10612,N_10438,N_10481);
nor U10613 (N_10613,N_10556,N_10460);
xor U10614 (N_10614,N_10419,N_10532);
or U10615 (N_10615,N_10501,N_10590);
nand U10616 (N_10616,N_10521,N_10571);
or U10617 (N_10617,N_10489,N_10592);
nand U10618 (N_10618,N_10468,N_10533);
or U10619 (N_10619,N_10491,N_10560);
nand U10620 (N_10620,N_10472,N_10513);
nand U10621 (N_10621,N_10569,N_10440);
or U10622 (N_10622,N_10584,N_10567);
nor U10623 (N_10623,N_10408,N_10410);
nor U10624 (N_10624,N_10514,N_10439);
or U10625 (N_10625,N_10598,N_10568);
nand U10626 (N_10626,N_10487,N_10517);
and U10627 (N_10627,N_10518,N_10539);
nor U10628 (N_10628,N_10586,N_10495);
nor U10629 (N_10629,N_10418,N_10519);
xor U10630 (N_10630,N_10411,N_10488);
and U10631 (N_10631,N_10483,N_10482);
or U10632 (N_10632,N_10423,N_10449);
or U10633 (N_10633,N_10545,N_10446);
xnor U10634 (N_10634,N_10434,N_10580);
and U10635 (N_10635,N_10558,N_10471);
nor U10636 (N_10636,N_10480,N_10534);
xor U10637 (N_10637,N_10429,N_10541);
nor U10638 (N_10638,N_10403,N_10476);
xnor U10639 (N_10639,N_10511,N_10551);
and U10640 (N_10640,N_10515,N_10561);
xor U10641 (N_10641,N_10576,N_10536);
nor U10642 (N_10642,N_10459,N_10526);
nor U10643 (N_10643,N_10442,N_10413);
nand U10644 (N_10644,N_10525,N_10553);
nand U10645 (N_10645,N_10407,N_10436);
nand U10646 (N_10646,N_10432,N_10485);
nor U10647 (N_10647,N_10461,N_10548);
nor U10648 (N_10648,N_10450,N_10524);
nor U10649 (N_10649,N_10554,N_10550);
nor U10650 (N_10650,N_10498,N_10428);
nand U10651 (N_10651,N_10454,N_10531);
or U10652 (N_10652,N_10574,N_10508);
nand U10653 (N_10653,N_10547,N_10430);
or U10654 (N_10654,N_10435,N_10464);
or U10655 (N_10655,N_10557,N_10443);
nor U10656 (N_10656,N_10477,N_10552);
xor U10657 (N_10657,N_10591,N_10543);
nor U10658 (N_10658,N_10506,N_10473);
nand U10659 (N_10659,N_10507,N_10404);
and U10660 (N_10660,N_10503,N_10500);
xor U10661 (N_10661,N_10484,N_10475);
or U10662 (N_10662,N_10520,N_10502);
nor U10663 (N_10663,N_10585,N_10425);
xnor U10664 (N_10664,N_10523,N_10424);
and U10665 (N_10665,N_10499,N_10570);
or U10666 (N_10666,N_10456,N_10596);
or U10667 (N_10667,N_10465,N_10492);
xor U10668 (N_10668,N_10566,N_10406);
nor U10669 (N_10669,N_10420,N_10415);
or U10670 (N_10670,N_10416,N_10562);
nor U10671 (N_10671,N_10469,N_10588);
xnor U10672 (N_10672,N_10582,N_10453);
or U10673 (N_10673,N_10433,N_10412);
or U10674 (N_10674,N_10457,N_10470);
and U10675 (N_10675,N_10462,N_10530);
nor U10676 (N_10676,N_10490,N_10505);
and U10677 (N_10677,N_10577,N_10528);
and U10678 (N_10678,N_10537,N_10445);
nor U10679 (N_10679,N_10448,N_10546);
and U10680 (N_10680,N_10400,N_10599);
nand U10681 (N_10681,N_10589,N_10510);
and U10682 (N_10682,N_10544,N_10401);
nand U10683 (N_10683,N_10494,N_10593);
or U10684 (N_10684,N_10496,N_10437);
nand U10685 (N_10685,N_10431,N_10426);
nor U10686 (N_10686,N_10458,N_10405);
nand U10687 (N_10687,N_10452,N_10467);
xnor U10688 (N_10688,N_10447,N_10478);
nor U10689 (N_10689,N_10594,N_10417);
or U10690 (N_10690,N_10414,N_10527);
or U10691 (N_10691,N_10587,N_10486);
xor U10692 (N_10692,N_10509,N_10479);
xor U10693 (N_10693,N_10559,N_10512);
or U10694 (N_10694,N_10549,N_10575);
and U10695 (N_10695,N_10578,N_10563);
nand U10696 (N_10696,N_10572,N_10579);
and U10697 (N_10697,N_10529,N_10581);
nor U10698 (N_10698,N_10474,N_10555);
nand U10699 (N_10699,N_10441,N_10573);
xnor U10700 (N_10700,N_10430,N_10536);
and U10701 (N_10701,N_10565,N_10551);
or U10702 (N_10702,N_10565,N_10457);
xnor U10703 (N_10703,N_10514,N_10418);
or U10704 (N_10704,N_10528,N_10583);
and U10705 (N_10705,N_10407,N_10596);
nor U10706 (N_10706,N_10583,N_10452);
nor U10707 (N_10707,N_10572,N_10584);
and U10708 (N_10708,N_10400,N_10465);
nand U10709 (N_10709,N_10401,N_10431);
nand U10710 (N_10710,N_10537,N_10580);
or U10711 (N_10711,N_10485,N_10510);
nand U10712 (N_10712,N_10443,N_10403);
and U10713 (N_10713,N_10412,N_10552);
or U10714 (N_10714,N_10552,N_10430);
nor U10715 (N_10715,N_10452,N_10573);
nor U10716 (N_10716,N_10582,N_10464);
nand U10717 (N_10717,N_10508,N_10423);
xor U10718 (N_10718,N_10564,N_10433);
or U10719 (N_10719,N_10435,N_10572);
nor U10720 (N_10720,N_10560,N_10478);
or U10721 (N_10721,N_10433,N_10470);
or U10722 (N_10722,N_10504,N_10559);
xor U10723 (N_10723,N_10503,N_10473);
or U10724 (N_10724,N_10480,N_10548);
or U10725 (N_10725,N_10404,N_10501);
nand U10726 (N_10726,N_10525,N_10477);
nor U10727 (N_10727,N_10471,N_10404);
and U10728 (N_10728,N_10410,N_10453);
nor U10729 (N_10729,N_10441,N_10545);
or U10730 (N_10730,N_10421,N_10534);
and U10731 (N_10731,N_10433,N_10441);
nor U10732 (N_10732,N_10593,N_10446);
or U10733 (N_10733,N_10500,N_10429);
or U10734 (N_10734,N_10502,N_10456);
xnor U10735 (N_10735,N_10595,N_10404);
or U10736 (N_10736,N_10537,N_10591);
or U10737 (N_10737,N_10435,N_10590);
nor U10738 (N_10738,N_10424,N_10561);
nand U10739 (N_10739,N_10524,N_10481);
nand U10740 (N_10740,N_10491,N_10422);
and U10741 (N_10741,N_10577,N_10588);
or U10742 (N_10742,N_10527,N_10575);
and U10743 (N_10743,N_10415,N_10460);
xnor U10744 (N_10744,N_10434,N_10504);
and U10745 (N_10745,N_10479,N_10550);
xnor U10746 (N_10746,N_10588,N_10451);
xnor U10747 (N_10747,N_10442,N_10479);
nor U10748 (N_10748,N_10582,N_10573);
or U10749 (N_10749,N_10417,N_10576);
and U10750 (N_10750,N_10518,N_10486);
nor U10751 (N_10751,N_10544,N_10445);
nor U10752 (N_10752,N_10536,N_10434);
nand U10753 (N_10753,N_10453,N_10523);
nand U10754 (N_10754,N_10404,N_10535);
or U10755 (N_10755,N_10459,N_10431);
nand U10756 (N_10756,N_10431,N_10491);
or U10757 (N_10757,N_10510,N_10528);
and U10758 (N_10758,N_10585,N_10438);
nor U10759 (N_10759,N_10570,N_10592);
nor U10760 (N_10760,N_10510,N_10526);
or U10761 (N_10761,N_10561,N_10517);
or U10762 (N_10762,N_10492,N_10520);
or U10763 (N_10763,N_10587,N_10510);
and U10764 (N_10764,N_10592,N_10594);
nand U10765 (N_10765,N_10597,N_10483);
nand U10766 (N_10766,N_10519,N_10551);
nor U10767 (N_10767,N_10578,N_10446);
or U10768 (N_10768,N_10539,N_10573);
or U10769 (N_10769,N_10487,N_10568);
and U10770 (N_10770,N_10536,N_10476);
or U10771 (N_10771,N_10414,N_10592);
and U10772 (N_10772,N_10457,N_10530);
or U10773 (N_10773,N_10470,N_10435);
and U10774 (N_10774,N_10447,N_10589);
nand U10775 (N_10775,N_10539,N_10410);
and U10776 (N_10776,N_10491,N_10487);
and U10777 (N_10777,N_10555,N_10404);
or U10778 (N_10778,N_10564,N_10425);
and U10779 (N_10779,N_10502,N_10411);
nand U10780 (N_10780,N_10535,N_10572);
or U10781 (N_10781,N_10539,N_10554);
xor U10782 (N_10782,N_10418,N_10438);
nor U10783 (N_10783,N_10501,N_10413);
and U10784 (N_10784,N_10577,N_10466);
nand U10785 (N_10785,N_10438,N_10433);
and U10786 (N_10786,N_10599,N_10463);
or U10787 (N_10787,N_10530,N_10468);
nor U10788 (N_10788,N_10403,N_10498);
nor U10789 (N_10789,N_10533,N_10508);
nand U10790 (N_10790,N_10511,N_10506);
or U10791 (N_10791,N_10512,N_10595);
and U10792 (N_10792,N_10489,N_10413);
and U10793 (N_10793,N_10533,N_10416);
nand U10794 (N_10794,N_10575,N_10518);
nor U10795 (N_10795,N_10426,N_10567);
nor U10796 (N_10796,N_10428,N_10471);
nand U10797 (N_10797,N_10459,N_10509);
nand U10798 (N_10798,N_10542,N_10445);
and U10799 (N_10799,N_10459,N_10466);
nand U10800 (N_10800,N_10652,N_10683);
and U10801 (N_10801,N_10694,N_10687);
and U10802 (N_10802,N_10656,N_10738);
nand U10803 (N_10803,N_10788,N_10624);
and U10804 (N_10804,N_10756,N_10716);
nand U10805 (N_10805,N_10718,N_10782);
or U10806 (N_10806,N_10696,N_10795);
and U10807 (N_10807,N_10721,N_10762);
or U10808 (N_10808,N_10761,N_10744);
or U10809 (N_10809,N_10711,N_10771);
or U10810 (N_10810,N_10612,N_10606);
nor U10811 (N_10811,N_10631,N_10659);
nand U10812 (N_10812,N_10660,N_10746);
nor U10813 (N_10813,N_10726,N_10641);
nand U10814 (N_10814,N_10786,N_10627);
or U10815 (N_10815,N_10698,N_10715);
nor U10816 (N_10816,N_10610,N_10642);
and U10817 (N_10817,N_10603,N_10789);
or U10818 (N_10818,N_10630,N_10697);
nand U10819 (N_10819,N_10668,N_10604);
nor U10820 (N_10820,N_10619,N_10614);
or U10821 (N_10821,N_10628,N_10702);
xor U10822 (N_10822,N_10763,N_10663);
and U10823 (N_10823,N_10722,N_10773);
nand U10824 (N_10824,N_10649,N_10787);
and U10825 (N_10825,N_10772,N_10766);
nand U10826 (N_10826,N_10775,N_10684);
nor U10827 (N_10827,N_10617,N_10770);
and U10828 (N_10828,N_10677,N_10602);
nand U10829 (N_10829,N_10749,N_10752);
nor U10830 (N_10830,N_10751,N_10760);
nand U10831 (N_10831,N_10730,N_10713);
and U10832 (N_10832,N_10759,N_10701);
or U10833 (N_10833,N_10705,N_10758);
nand U10834 (N_10834,N_10618,N_10785);
or U10835 (N_10835,N_10662,N_10664);
nand U10836 (N_10836,N_10736,N_10676);
nor U10837 (N_10837,N_10647,N_10689);
and U10838 (N_10838,N_10710,N_10797);
or U10839 (N_10839,N_10693,N_10757);
and U10840 (N_10840,N_10737,N_10613);
and U10841 (N_10841,N_10682,N_10674);
and U10842 (N_10842,N_10699,N_10622);
nand U10843 (N_10843,N_10670,N_10767);
nor U10844 (N_10844,N_10626,N_10608);
and U10845 (N_10845,N_10796,N_10672);
nand U10846 (N_10846,N_10743,N_10679);
nand U10847 (N_10847,N_10655,N_10720);
nor U10848 (N_10848,N_10725,N_10667);
nor U10849 (N_10849,N_10779,N_10791);
or U10850 (N_10850,N_10723,N_10724);
or U10851 (N_10851,N_10629,N_10755);
or U10852 (N_10852,N_10704,N_10768);
nand U10853 (N_10853,N_10707,N_10638);
and U10854 (N_10854,N_10690,N_10609);
or U10855 (N_10855,N_10792,N_10793);
nand U10856 (N_10856,N_10644,N_10776);
nor U10857 (N_10857,N_10794,N_10769);
nor U10858 (N_10858,N_10681,N_10728);
nor U10859 (N_10859,N_10798,N_10633);
nor U10860 (N_10860,N_10675,N_10637);
or U10861 (N_10861,N_10727,N_10712);
xor U10862 (N_10862,N_10623,N_10734);
nor U10863 (N_10863,N_10739,N_10600);
nor U10864 (N_10864,N_10735,N_10784);
and U10865 (N_10865,N_10777,N_10607);
xor U10866 (N_10866,N_10780,N_10601);
or U10867 (N_10867,N_10666,N_10673);
or U10868 (N_10868,N_10790,N_10625);
and U10869 (N_10869,N_10653,N_10616);
and U10870 (N_10870,N_10733,N_10651);
nand U10871 (N_10871,N_10717,N_10732);
xnor U10872 (N_10872,N_10740,N_10658);
nand U10873 (N_10873,N_10764,N_10605);
nand U10874 (N_10874,N_10695,N_10703);
nand U10875 (N_10875,N_10706,N_10748);
nand U10876 (N_10876,N_10731,N_10661);
or U10877 (N_10877,N_10708,N_10635);
nor U10878 (N_10878,N_10700,N_10781);
nor U10879 (N_10879,N_10778,N_10799);
nor U10880 (N_10880,N_10680,N_10742);
and U10881 (N_10881,N_10639,N_10691);
and U10882 (N_10882,N_10671,N_10615);
nor U10883 (N_10883,N_10640,N_10774);
nand U10884 (N_10884,N_10692,N_10750);
or U10885 (N_10885,N_10669,N_10665);
or U10886 (N_10886,N_10719,N_10688);
xor U10887 (N_10887,N_10648,N_10611);
or U10888 (N_10888,N_10646,N_10783);
xor U10889 (N_10889,N_10741,N_10753);
or U10890 (N_10890,N_10636,N_10709);
nor U10891 (N_10891,N_10765,N_10729);
nand U10892 (N_10892,N_10678,N_10754);
nor U10893 (N_10893,N_10632,N_10643);
and U10894 (N_10894,N_10620,N_10747);
or U10895 (N_10895,N_10745,N_10685);
nor U10896 (N_10896,N_10686,N_10621);
or U10897 (N_10897,N_10645,N_10714);
nand U10898 (N_10898,N_10654,N_10657);
nor U10899 (N_10899,N_10634,N_10650);
xnor U10900 (N_10900,N_10766,N_10692);
and U10901 (N_10901,N_10731,N_10768);
nand U10902 (N_10902,N_10756,N_10629);
nand U10903 (N_10903,N_10715,N_10727);
nand U10904 (N_10904,N_10762,N_10610);
and U10905 (N_10905,N_10746,N_10724);
nor U10906 (N_10906,N_10792,N_10660);
and U10907 (N_10907,N_10605,N_10766);
or U10908 (N_10908,N_10693,N_10666);
nor U10909 (N_10909,N_10609,N_10619);
or U10910 (N_10910,N_10722,N_10650);
and U10911 (N_10911,N_10762,N_10664);
nor U10912 (N_10912,N_10741,N_10711);
and U10913 (N_10913,N_10682,N_10613);
and U10914 (N_10914,N_10771,N_10609);
or U10915 (N_10915,N_10772,N_10680);
nand U10916 (N_10916,N_10693,N_10605);
or U10917 (N_10917,N_10633,N_10704);
or U10918 (N_10918,N_10716,N_10637);
and U10919 (N_10919,N_10770,N_10669);
nor U10920 (N_10920,N_10613,N_10707);
and U10921 (N_10921,N_10685,N_10628);
or U10922 (N_10922,N_10618,N_10629);
nor U10923 (N_10923,N_10690,N_10644);
and U10924 (N_10924,N_10679,N_10710);
nor U10925 (N_10925,N_10649,N_10679);
and U10926 (N_10926,N_10701,N_10789);
nand U10927 (N_10927,N_10635,N_10734);
nand U10928 (N_10928,N_10704,N_10695);
nand U10929 (N_10929,N_10728,N_10642);
xnor U10930 (N_10930,N_10764,N_10606);
or U10931 (N_10931,N_10606,N_10768);
nor U10932 (N_10932,N_10602,N_10617);
or U10933 (N_10933,N_10742,N_10633);
and U10934 (N_10934,N_10627,N_10621);
xor U10935 (N_10935,N_10766,N_10695);
and U10936 (N_10936,N_10621,N_10718);
and U10937 (N_10937,N_10670,N_10602);
and U10938 (N_10938,N_10721,N_10742);
nand U10939 (N_10939,N_10686,N_10776);
nor U10940 (N_10940,N_10605,N_10623);
nand U10941 (N_10941,N_10713,N_10644);
or U10942 (N_10942,N_10719,N_10769);
nand U10943 (N_10943,N_10676,N_10628);
xnor U10944 (N_10944,N_10604,N_10728);
and U10945 (N_10945,N_10645,N_10636);
nand U10946 (N_10946,N_10668,N_10694);
xnor U10947 (N_10947,N_10655,N_10656);
and U10948 (N_10948,N_10755,N_10645);
nor U10949 (N_10949,N_10625,N_10653);
or U10950 (N_10950,N_10665,N_10639);
nor U10951 (N_10951,N_10784,N_10660);
nand U10952 (N_10952,N_10720,N_10694);
or U10953 (N_10953,N_10752,N_10691);
nand U10954 (N_10954,N_10715,N_10721);
nor U10955 (N_10955,N_10637,N_10686);
or U10956 (N_10956,N_10759,N_10786);
nor U10957 (N_10957,N_10784,N_10670);
or U10958 (N_10958,N_10668,N_10766);
or U10959 (N_10959,N_10796,N_10726);
or U10960 (N_10960,N_10768,N_10692);
and U10961 (N_10961,N_10685,N_10774);
or U10962 (N_10962,N_10783,N_10749);
and U10963 (N_10963,N_10733,N_10616);
or U10964 (N_10964,N_10759,N_10666);
and U10965 (N_10965,N_10754,N_10758);
or U10966 (N_10966,N_10748,N_10665);
nand U10967 (N_10967,N_10788,N_10740);
and U10968 (N_10968,N_10776,N_10785);
and U10969 (N_10969,N_10649,N_10678);
nand U10970 (N_10970,N_10664,N_10733);
nand U10971 (N_10971,N_10674,N_10642);
nand U10972 (N_10972,N_10796,N_10605);
and U10973 (N_10973,N_10712,N_10660);
nand U10974 (N_10974,N_10679,N_10685);
or U10975 (N_10975,N_10756,N_10683);
and U10976 (N_10976,N_10619,N_10783);
and U10977 (N_10977,N_10703,N_10779);
nor U10978 (N_10978,N_10754,N_10642);
nand U10979 (N_10979,N_10663,N_10625);
and U10980 (N_10980,N_10740,N_10610);
nand U10981 (N_10981,N_10657,N_10653);
nand U10982 (N_10982,N_10705,N_10707);
and U10983 (N_10983,N_10785,N_10781);
nand U10984 (N_10984,N_10637,N_10741);
xnor U10985 (N_10985,N_10649,N_10669);
nand U10986 (N_10986,N_10640,N_10703);
or U10987 (N_10987,N_10712,N_10731);
nor U10988 (N_10988,N_10759,N_10716);
nand U10989 (N_10989,N_10701,N_10714);
or U10990 (N_10990,N_10669,N_10607);
nand U10991 (N_10991,N_10777,N_10651);
and U10992 (N_10992,N_10753,N_10616);
xor U10993 (N_10993,N_10600,N_10643);
nand U10994 (N_10994,N_10686,N_10707);
nor U10995 (N_10995,N_10677,N_10766);
nand U10996 (N_10996,N_10667,N_10744);
and U10997 (N_10997,N_10656,N_10606);
and U10998 (N_10998,N_10698,N_10617);
and U10999 (N_10999,N_10613,N_10698);
nand U11000 (N_11000,N_10873,N_10911);
xnor U11001 (N_11001,N_10923,N_10986);
nand U11002 (N_11002,N_10890,N_10973);
and U11003 (N_11003,N_10983,N_10945);
nand U11004 (N_11004,N_10866,N_10994);
nor U11005 (N_11005,N_10906,N_10925);
nand U11006 (N_11006,N_10965,N_10903);
nand U11007 (N_11007,N_10932,N_10860);
xnor U11008 (N_11008,N_10868,N_10908);
nand U11009 (N_11009,N_10912,N_10820);
and U11010 (N_11010,N_10982,N_10807);
and U11011 (N_11011,N_10926,N_10905);
nor U11012 (N_11012,N_10990,N_10872);
or U11013 (N_11013,N_10825,N_10991);
or U11014 (N_11014,N_10985,N_10839);
and U11015 (N_11015,N_10850,N_10957);
nand U11016 (N_11016,N_10929,N_10917);
and U11017 (N_11017,N_10933,N_10819);
nand U11018 (N_11018,N_10884,N_10801);
nor U11019 (N_11019,N_10888,N_10913);
nor U11020 (N_11020,N_10992,N_10811);
nor U11021 (N_11021,N_10845,N_10855);
nor U11022 (N_11022,N_10821,N_10892);
and U11023 (N_11023,N_10854,N_10924);
and U11024 (N_11024,N_10998,N_10812);
and U11025 (N_11025,N_10987,N_10838);
nor U11026 (N_11026,N_10975,N_10803);
or U11027 (N_11027,N_10830,N_10919);
or U11028 (N_11028,N_10877,N_10804);
and U11029 (N_11029,N_10887,N_10995);
and U11030 (N_11030,N_10802,N_10953);
nor U11031 (N_11031,N_10902,N_10893);
nor U11032 (N_11032,N_10993,N_10837);
or U11033 (N_11033,N_10823,N_10907);
nor U11034 (N_11034,N_10954,N_10824);
and U11035 (N_11035,N_10897,N_10808);
nand U11036 (N_11036,N_10881,N_10978);
nor U11037 (N_11037,N_10891,N_10922);
and U11038 (N_11038,N_10843,N_10878);
and U11039 (N_11039,N_10840,N_10856);
nand U11040 (N_11040,N_10870,N_10981);
nand U11041 (N_11041,N_10876,N_10951);
and U11042 (N_11042,N_10832,N_10946);
nand U11043 (N_11043,N_10949,N_10880);
and U11044 (N_11044,N_10875,N_10955);
nand U11045 (N_11045,N_10950,N_10961);
nor U11046 (N_11046,N_10970,N_10871);
nor U11047 (N_11047,N_10916,N_10846);
nor U11048 (N_11048,N_10861,N_10827);
or U11049 (N_11049,N_10937,N_10952);
nand U11050 (N_11050,N_10867,N_10869);
and U11051 (N_11051,N_10989,N_10968);
or U11052 (N_11052,N_10901,N_10938);
or U11053 (N_11053,N_10900,N_10805);
and U11054 (N_11054,N_10883,N_10822);
and U11055 (N_11055,N_10962,N_10814);
or U11056 (N_11056,N_10806,N_10918);
nand U11057 (N_11057,N_10818,N_10979);
or U11058 (N_11058,N_10874,N_10879);
xnor U11059 (N_11059,N_10800,N_10841);
nand U11060 (N_11060,N_10859,N_10936);
nand U11061 (N_11061,N_10935,N_10966);
nor U11062 (N_11062,N_10960,N_10842);
xnor U11063 (N_11063,N_10921,N_10943);
nand U11064 (N_11064,N_10894,N_10964);
nand U11065 (N_11065,N_10828,N_10984);
or U11066 (N_11066,N_10858,N_10977);
nor U11067 (N_11067,N_10864,N_10996);
and U11068 (N_11068,N_10959,N_10909);
nor U11069 (N_11069,N_10980,N_10956);
or U11070 (N_11070,N_10930,N_10847);
nand U11071 (N_11071,N_10810,N_10809);
nand U11072 (N_11072,N_10829,N_10857);
and U11073 (N_11073,N_10836,N_10853);
and U11074 (N_11074,N_10849,N_10988);
or U11075 (N_11075,N_10835,N_10948);
nor U11076 (N_11076,N_10815,N_10972);
nor U11077 (N_11077,N_10851,N_10831);
nand U11078 (N_11078,N_10844,N_10941);
xnor U11079 (N_11079,N_10947,N_10963);
or U11080 (N_11080,N_10886,N_10976);
xor U11081 (N_11081,N_10826,N_10813);
nand U11082 (N_11082,N_10885,N_10817);
nand U11083 (N_11083,N_10999,N_10971);
or U11084 (N_11084,N_10931,N_10889);
nor U11085 (N_11085,N_10852,N_10904);
and U11086 (N_11086,N_10833,N_10914);
or U11087 (N_11087,N_10939,N_10862);
or U11088 (N_11088,N_10895,N_10898);
or U11089 (N_11089,N_10899,N_10896);
nand U11090 (N_11090,N_10834,N_10863);
and U11091 (N_11091,N_10974,N_10944);
xor U11092 (N_11092,N_10816,N_10882);
and U11093 (N_11093,N_10934,N_10927);
nand U11094 (N_11094,N_10940,N_10928);
or U11095 (N_11095,N_10958,N_10848);
nor U11096 (N_11096,N_10942,N_10915);
xnor U11097 (N_11097,N_10967,N_10865);
nand U11098 (N_11098,N_10910,N_10997);
and U11099 (N_11099,N_10920,N_10969);
nor U11100 (N_11100,N_10978,N_10940);
nor U11101 (N_11101,N_10984,N_10931);
nand U11102 (N_11102,N_10998,N_10932);
nor U11103 (N_11103,N_10824,N_10896);
and U11104 (N_11104,N_10904,N_10866);
or U11105 (N_11105,N_10801,N_10921);
nand U11106 (N_11106,N_10823,N_10948);
xor U11107 (N_11107,N_10959,N_10933);
and U11108 (N_11108,N_10919,N_10927);
nor U11109 (N_11109,N_10971,N_10977);
or U11110 (N_11110,N_10976,N_10892);
nand U11111 (N_11111,N_10899,N_10913);
xor U11112 (N_11112,N_10985,N_10923);
xor U11113 (N_11113,N_10927,N_10816);
nand U11114 (N_11114,N_10944,N_10863);
and U11115 (N_11115,N_10878,N_10927);
nor U11116 (N_11116,N_10976,N_10846);
or U11117 (N_11117,N_10817,N_10862);
nand U11118 (N_11118,N_10889,N_10816);
nor U11119 (N_11119,N_10973,N_10959);
xnor U11120 (N_11120,N_10816,N_10973);
nor U11121 (N_11121,N_10904,N_10978);
and U11122 (N_11122,N_10913,N_10803);
and U11123 (N_11123,N_10864,N_10984);
nand U11124 (N_11124,N_10903,N_10982);
or U11125 (N_11125,N_10975,N_10878);
and U11126 (N_11126,N_10814,N_10977);
xnor U11127 (N_11127,N_10883,N_10893);
or U11128 (N_11128,N_10901,N_10961);
or U11129 (N_11129,N_10833,N_10991);
or U11130 (N_11130,N_10811,N_10827);
and U11131 (N_11131,N_10848,N_10827);
or U11132 (N_11132,N_10868,N_10944);
and U11133 (N_11133,N_10868,N_10801);
nand U11134 (N_11134,N_10898,N_10825);
nand U11135 (N_11135,N_10976,N_10862);
xor U11136 (N_11136,N_10946,N_10893);
nand U11137 (N_11137,N_10982,N_10979);
or U11138 (N_11138,N_10880,N_10809);
and U11139 (N_11139,N_10805,N_10931);
and U11140 (N_11140,N_10914,N_10942);
nor U11141 (N_11141,N_10879,N_10995);
nand U11142 (N_11142,N_10976,N_10951);
or U11143 (N_11143,N_10842,N_10870);
nor U11144 (N_11144,N_10897,N_10912);
nor U11145 (N_11145,N_10939,N_10867);
nor U11146 (N_11146,N_10840,N_10825);
nor U11147 (N_11147,N_10995,N_10987);
and U11148 (N_11148,N_10834,N_10846);
or U11149 (N_11149,N_10878,N_10872);
xor U11150 (N_11150,N_10823,N_10843);
xnor U11151 (N_11151,N_10895,N_10981);
nand U11152 (N_11152,N_10960,N_10966);
or U11153 (N_11153,N_10800,N_10961);
xnor U11154 (N_11154,N_10808,N_10900);
xnor U11155 (N_11155,N_10912,N_10805);
nand U11156 (N_11156,N_10913,N_10875);
nor U11157 (N_11157,N_10910,N_10946);
nor U11158 (N_11158,N_10951,N_10882);
or U11159 (N_11159,N_10819,N_10872);
nor U11160 (N_11160,N_10881,N_10985);
nor U11161 (N_11161,N_10809,N_10849);
nand U11162 (N_11162,N_10805,N_10942);
xor U11163 (N_11163,N_10828,N_10800);
xor U11164 (N_11164,N_10964,N_10849);
and U11165 (N_11165,N_10826,N_10884);
nor U11166 (N_11166,N_10874,N_10933);
nor U11167 (N_11167,N_10866,N_10876);
and U11168 (N_11168,N_10933,N_10938);
nand U11169 (N_11169,N_10912,N_10860);
or U11170 (N_11170,N_10954,N_10967);
nand U11171 (N_11171,N_10948,N_10867);
xnor U11172 (N_11172,N_10855,N_10846);
and U11173 (N_11173,N_10865,N_10909);
xor U11174 (N_11174,N_10815,N_10997);
xnor U11175 (N_11175,N_10875,N_10930);
xnor U11176 (N_11176,N_10834,N_10977);
or U11177 (N_11177,N_10808,N_10813);
nand U11178 (N_11178,N_10865,N_10886);
or U11179 (N_11179,N_10883,N_10957);
and U11180 (N_11180,N_10892,N_10896);
nor U11181 (N_11181,N_10996,N_10808);
and U11182 (N_11182,N_10944,N_10952);
nor U11183 (N_11183,N_10805,N_10926);
nor U11184 (N_11184,N_10985,N_10851);
nor U11185 (N_11185,N_10807,N_10947);
xor U11186 (N_11186,N_10801,N_10962);
nand U11187 (N_11187,N_10922,N_10913);
and U11188 (N_11188,N_10878,N_10819);
and U11189 (N_11189,N_10983,N_10972);
nor U11190 (N_11190,N_10961,N_10956);
xnor U11191 (N_11191,N_10810,N_10989);
nor U11192 (N_11192,N_10949,N_10863);
or U11193 (N_11193,N_10951,N_10921);
nor U11194 (N_11194,N_10905,N_10963);
nor U11195 (N_11195,N_10990,N_10897);
and U11196 (N_11196,N_10813,N_10935);
and U11197 (N_11197,N_10842,N_10823);
and U11198 (N_11198,N_10960,N_10809);
nor U11199 (N_11199,N_10974,N_10991);
and U11200 (N_11200,N_11100,N_11169);
and U11201 (N_11201,N_11016,N_11126);
nand U11202 (N_11202,N_11021,N_11103);
or U11203 (N_11203,N_11076,N_11085);
nor U11204 (N_11204,N_11051,N_11041);
nor U11205 (N_11205,N_11143,N_11149);
nand U11206 (N_11206,N_11023,N_11158);
nor U11207 (N_11207,N_11001,N_11039);
or U11208 (N_11208,N_11013,N_11119);
nand U11209 (N_11209,N_11186,N_11132);
nand U11210 (N_11210,N_11179,N_11114);
nor U11211 (N_11211,N_11134,N_11115);
and U11212 (N_11212,N_11092,N_11160);
or U11213 (N_11213,N_11060,N_11043);
nor U11214 (N_11214,N_11002,N_11022);
nand U11215 (N_11215,N_11064,N_11157);
nor U11216 (N_11216,N_11019,N_11101);
nand U11217 (N_11217,N_11156,N_11094);
or U11218 (N_11218,N_11097,N_11127);
nand U11219 (N_11219,N_11151,N_11141);
nand U11220 (N_11220,N_11144,N_11189);
nand U11221 (N_11221,N_11018,N_11099);
or U11222 (N_11222,N_11024,N_11140);
and U11223 (N_11223,N_11117,N_11010);
nand U11224 (N_11224,N_11004,N_11185);
or U11225 (N_11225,N_11130,N_11125);
nor U11226 (N_11226,N_11148,N_11145);
nand U11227 (N_11227,N_11164,N_11083);
and U11228 (N_11228,N_11086,N_11098);
xnor U11229 (N_11229,N_11007,N_11011);
and U11230 (N_11230,N_11102,N_11034);
nand U11231 (N_11231,N_11135,N_11162);
nand U11232 (N_11232,N_11014,N_11072);
and U11233 (N_11233,N_11123,N_11163);
nor U11234 (N_11234,N_11167,N_11192);
nor U11235 (N_11235,N_11009,N_11178);
xor U11236 (N_11236,N_11069,N_11059);
and U11237 (N_11237,N_11046,N_11177);
nor U11238 (N_11238,N_11070,N_11031);
nand U11239 (N_11239,N_11017,N_11173);
nand U11240 (N_11240,N_11142,N_11065);
and U11241 (N_11241,N_11029,N_11066);
or U11242 (N_11242,N_11030,N_11105);
nand U11243 (N_11243,N_11188,N_11068);
and U11244 (N_11244,N_11147,N_11104);
nand U11245 (N_11245,N_11184,N_11063);
or U11246 (N_11246,N_11080,N_11047);
nor U11247 (N_11247,N_11079,N_11109);
xnor U11248 (N_11248,N_11042,N_11054);
nor U11249 (N_11249,N_11195,N_11074);
nand U11250 (N_11250,N_11035,N_11000);
nand U11251 (N_11251,N_11095,N_11111);
and U11252 (N_11252,N_11187,N_11137);
and U11253 (N_11253,N_11058,N_11071);
nor U11254 (N_11254,N_11120,N_11174);
nand U11255 (N_11255,N_11067,N_11045);
and U11256 (N_11256,N_11028,N_11052);
nor U11257 (N_11257,N_11182,N_11027);
or U11258 (N_11258,N_11183,N_11176);
nor U11259 (N_11259,N_11049,N_11012);
and U11260 (N_11260,N_11131,N_11062);
or U11261 (N_11261,N_11138,N_11044);
nor U11262 (N_11262,N_11033,N_11146);
nor U11263 (N_11263,N_11025,N_11166);
and U11264 (N_11264,N_11078,N_11161);
or U11265 (N_11265,N_11088,N_11038);
nand U11266 (N_11266,N_11053,N_11168);
and U11267 (N_11267,N_11118,N_11129);
nand U11268 (N_11268,N_11006,N_11198);
or U11269 (N_11269,N_11003,N_11026);
xnor U11270 (N_11270,N_11048,N_11108);
and U11271 (N_11271,N_11170,N_11128);
or U11272 (N_11272,N_11180,N_11171);
xnor U11273 (N_11273,N_11159,N_11084);
nand U11274 (N_11274,N_11110,N_11077);
and U11275 (N_11275,N_11175,N_11193);
xor U11276 (N_11276,N_11008,N_11112);
xor U11277 (N_11277,N_11106,N_11122);
and U11278 (N_11278,N_11096,N_11090);
and U11279 (N_11279,N_11089,N_11032);
nor U11280 (N_11280,N_11020,N_11121);
nand U11281 (N_11281,N_11036,N_11197);
nor U11282 (N_11282,N_11194,N_11165);
or U11283 (N_11283,N_11107,N_11091);
and U11284 (N_11284,N_11154,N_11015);
nor U11285 (N_11285,N_11093,N_11124);
and U11286 (N_11286,N_11081,N_11040);
and U11287 (N_11287,N_11191,N_11116);
nor U11288 (N_11288,N_11136,N_11075);
and U11289 (N_11289,N_11082,N_11133);
nor U11290 (N_11290,N_11153,N_11190);
and U11291 (N_11291,N_11172,N_11139);
nand U11292 (N_11292,N_11150,N_11152);
and U11293 (N_11293,N_11181,N_11155);
nor U11294 (N_11294,N_11055,N_11113);
or U11295 (N_11295,N_11050,N_11199);
nor U11296 (N_11296,N_11073,N_11087);
nor U11297 (N_11297,N_11061,N_11056);
or U11298 (N_11298,N_11057,N_11005);
and U11299 (N_11299,N_11196,N_11037);
and U11300 (N_11300,N_11170,N_11049);
nand U11301 (N_11301,N_11194,N_11182);
and U11302 (N_11302,N_11049,N_11048);
nand U11303 (N_11303,N_11023,N_11060);
and U11304 (N_11304,N_11004,N_11151);
nand U11305 (N_11305,N_11145,N_11120);
nand U11306 (N_11306,N_11175,N_11192);
nor U11307 (N_11307,N_11125,N_11020);
or U11308 (N_11308,N_11118,N_11106);
nor U11309 (N_11309,N_11011,N_11076);
nand U11310 (N_11310,N_11184,N_11008);
nor U11311 (N_11311,N_11053,N_11001);
xor U11312 (N_11312,N_11124,N_11117);
or U11313 (N_11313,N_11002,N_11028);
or U11314 (N_11314,N_11165,N_11115);
nor U11315 (N_11315,N_11037,N_11099);
nor U11316 (N_11316,N_11137,N_11194);
or U11317 (N_11317,N_11096,N_11047);
nor U11318 (N_11318,N_11019,N_11141);
nor U11319 (N_11319,N_11058,N_11098);
nor U11320 (N_11320,N_11177,N_11150);
nand U11321 (N_11321,N_11096,N_11057);
xor U11322 (N_11322,N_11130,N_11071);
nor U11323 (N_11323,N_11042,N_11192);
nor U11324 (N_11324,N_11194,N_11086);
or U11325 (N_11325,N_11026,N_11048);
xnor U11326 (N_11326,N_11027,N_11043);
nor U11327 (N_11327,N_11069,N_11097);
or U11328 (N_11328,N_11171,N_11046);
nor U11329 (N_11329,N_11182,N_11199);
and U11330 (N_11330,N_11165,N_11138);
and U11331 (N_11331,N_11140,N_11117);
nor U11332 (N_11332,N_11167,N_11098);
or U11333 (N_11333,N_11185,N_11101);
nor U11334 (N_11334,N_11168,N_11026);
xnor U11335 (N_11335,N_11104,N_11196);
and U11336 (N_11336,N_11154,N_11197);
nor U11337 (N_11337,N_11044,N_11101);
nand U11338 (N_11338,N_11160,N_11033);
or U11339 (N_11339,N_11055,N_11193);
nand U11340 (N_11340,N_11062,N_11179);
or U11341 (N_11341,N_11030,N_11156);
and U11342 (N_11342,N_11005,N_11113);
or U11343 (N_11343,N_11118,N_11002);
and U11344 (N_11344,N_11138,N_11154);
xnor U11345 (N_11345,N_11108,N_11044);
nor U11346 (N_11346,N_11113,N_11081);
or U11347 (N_11347,N_11145,N_11187);
and U11348 (N_11348,N_11118,N_11070);
nor U11349 (N_11349,N_11190,N_11054);
nand U11350 (N_11350,N_11017,N_11066);
xnor U11351 (N_11351,N_11006,N_11160);
nor U11352 (N_11352,N_11163,N_11093);
nand U11353 (N_11353,N_11067,N_11061);
xor U11354 (N_11354,N_11185,N_11003);
xnor U11355 (N_11355,N_11158,N_11166);
nor U11356 (N_11356,N_11063,N_11143);
xnor U11357 (N_11357,N_11010,N_11195);
or U11358 (N_11358,N_11070,N_11037);
and U11359 (N_11359,N_11180,N_11159);
nor U11360 (N_11360,N_11119,N_11014);
nor U11361 (N_11361,N_11106,N_11000);
or U11362 (N_11362,N_11012,N_11134);
nor U11363 (N_11363,N_11126,N_11093);
nor U11364 (N_11364,N_11000,N_11193);
nand U11365 (N_11365,N_11071,N_11127);
nand U11366 (N_11366,N_11072,N_11147);
and U11367 (N_11367,N_11068,N_11055);
or U11368 (N_11368,N_11141,N_11108);
or U11369 (N_11369,N_11004,N_11006);
and U11370 (N_11370,N_11094,N_11138);
nand U11371 (N_11371,N_11064,N_11175);
nand U11372 (N_11372,N_11006,N_11175);
or U11373 (N_11373,N_11034,N_11118);
or U11374 (N_11374,N_11085,N_11054);
nor U11375 (N_11375,N_11048,N_11017);
nor U11376 (N_11376,N_11159,N_11156);
and U11377 (N_11377,N_11004,N_11146);
nor U11378 (N_11378,N_11106,N_11194);
nor U11379 (N_11379,N_11069,N_11144);
nand U11380 (N_11380,N_11110,N_11096);
nor U11381 (N_11381,N_11067,N_11186);
nand U11382 (N_11382,N_11098,N_11165);
and U11383 (N_11383,N_11037,N_11030);
nand U11384 (N_11384,N_11033,N_11092);
or U11385 (N_11385,N_11104,N_11085);
nor U11386 (N_11386,N_11113,N_11095);
xnor U11387 (N_11387,N_11196,N_11123);
xor U11388 (N_11388,N_11002,N_11031);
or U11389 (N_11389,N_11034,N_11082);
and U11390 (N_11390,N_11145,N_11168);
or U11391 (N_11391,N_11121,N_11019);
and U11392 (N_11392,N_11003,N_11190);
nand U11393 (N_11393,N_11190,N_11065);
or U11394 (N_11394,N_11021,N_11049);
nor U11395 (N_11395,N_11035,N_11086);
and U11396 (N_11396,N_11089,N_11181);
or U11397 (N_11397,N_11189,N_11180);
xor U11398 (N_11398,N_11059,N_11056);
and U11399 (N_11399,N_11189,N_11016);
or U11400 (N_11400,N_11248,N_11304);
nand U11401 (N_11401,N_11209,N_11277);
nand U11402 (N_11402,N_11308,N_11256);
and U11403 (N_11403,N_11371,N_11245);
or U11404 (N_11404,N_11294,N_11384);
nor U11405 (N_11405,N_11335,N_11303);
nor U11406 (N_11406,N_11390,N_11330);
or U11407 (N_11407,N_11306,N_11229);
nor U11408 (N_11408,N_11301,N_11244);
xnor U11409 (N_11409,N_11310,N_11313);
nor U11410 (N_11410,N_11269,N_11379);
nor U11411 (N_11411,N_11297,N_11341);
or U11412 (N_11412,N_11359,N_11385);
and U11413 (N_11413,N_11361,N_11287);
xor U11414 (N_11414,N_11273,N_11374);
nand U11415 (N_11415,N_11372,N_11261);
xnor U11416 (N_11416,N_11276,N_11227);
nand U11417 (N_11417,N_11238,N_11346);
and U11418 (N_11418,N_11201,N_11316);
nand U11419 (N_11419,N_11302,N_11397);
or U11420 (N_11420,N_11251,N_11311);
and U11421 (N_11421,N_11350,N_11319);
nor U11422 (N_11422,N_11228,N_11215);
xor U11423 (N_11423,N_11265,N_11236);
or U11424 (N_11424,N_11280,N_11250);
nor U11425 (N_11425,N_11231,N_11362);
nand U11426 (N_11426,N_11283,N_11324);
nand U11427 (N_11427,N_11300,N_11249);
nor U11428 (N_11428,N_11366,N_11377);
or U11429 (N_11429,N_11327,N_11355);
nand U11430 (N_11430,N_11381,N_11368);
nand U11431 (N_11431,N_11392,N_11360);
xnor U11432 (N_11432,N_11352,N_11275);
or U11433 (N_11433,N_11334,N_11376);
xnor U11434 (N_11434,N_11223,N_11246);
or U11435 (N_11435,N_11240,N_11378);
or U11436 (N_11436,N_11337,N_11203);
xor U11437 (N_11437,N_11382,N_11317);
and U11438 (N_11438,N_11290,N_11255);
and U11439 (N_11439,N_11260,N_11237);
nand U11440 (N_11440,N_11340,N_11314);
xnor U11441 (N_11441,N_11272,N_11218);
and U11442 (N_11442,N_11307,N_11387);
or U11443 (N_11443,N_11211,N_11270);
nor U11444 (N_11444,N_11295,N_11345);
nor U11445 (N_11445,N_11214,N_11296);
or U11446 (N_11446,N_11399,N_11204);
or U11447 (N_11447,N_11239,N_11386);
nor U11448 (N_11448,N_11282,N_11286);
nor U11449 (N_11449,N_11252,N_11291);
nand U11450 (N_11450,N_11370,N_11293);
nand U11451 (N_11451,N_11338,N_11348);
nand U11452 (N_11452,N_11358,N_11383);
or U11453 (N_11453,N_11267,N_11354);
and U11454 (N_11454,N_11257,N_11369);
nand U11455 (N_11455,N_11247,N_11225);
and U11456 (N_11456,N_11309,N_11343);
and U11457 (N_11457,N_11234,N_11339);
nor U11458 (N_11458,N_11226,N_11391);
or U11459 (N_11459,N_11213,N_11393);
and U11460 (N_11460,N_11388,N_11259);
or U11461 (N_11461,N_11318,N_11230);
and U11462 (N_11462,N_11274,N_11312);
or U11463 (N_11463,N_11298,N_11373);
xnor U11464 (N_11464,N_11342,N_11288);
xnor U11465 (N_11465,N_11212,N_11305);
and U11466 (N_11466,N_11266,N_11326);
or U11467 (N_11467,N_11241,N_11207);
or U11468 (N_11468,N_11353,N_11232);
or U11469 (N_11469,N_11216,N_11278);
or U11470 (N_11470,N_11221,N_11271);
xor U11471 (N_11471,N_11351,N_11323);
nand U11472 (N_11472,N_11364,N_11222);
and U11473 (N_11473,N_11285,N_11208);
and U11474 (N_11474,N_11263,N_11220);
nor U11475 (N_11475,N_11356,N_11320);
or U11476 (N_11476,N_11210,N_11344);
or U11477 (N_11477,N_11394,N_11332);
xor U11478 (N_11478,N_11268,N_11328);
and U11479 (N_11479,N_11380,N_11235);
nor U11480 (N_11480,N_11329,N_11347);
nor U11481 (N_11481,N_11331,N_11264);
and U11482 (N_11482,N_11205,N_11262);
and U11483 (N_11483,N_11224,N_11395);
nand U11484 (N_11484,N_11363,N_11333);
nor U11485 (N_11485,N_11292,N_11322);
or U11486 (N_11486,N_11281,N_11202);
or U11487 (N_11487,N_11284,N_11315);
nand U11488 (N_11488,N_11321,N_11279);
or U11489 (N_11489,N_11398,N_11258);
or U11490 (N_11490,N_11336,N_11242);
or U11491 (N_11491,N_11253,N_11325);
or U11492 (N_11492,N_11254,N_11375);
nand U11493 (N_11493,N_11349,N_11243);
and U11494 (N_11494,N_11219,N_11396);
or U11495 (N_11495,N_11217,N_11289);
nand U11496 (N_11496,N_11299,N_11206);
nand U11497 (N_11497,N_11367,N_11200);
nand U11498 (N_11498,N_11233,N_11389);
nor U11499 (N_11499,N_11365,N_11357);
or U11500 (N_11500,N_11203,N_11397);
xnor U11501 (N_11501,N_11363,N_11209);
nand U11502 (N_11502,N_11314,N_11363);
nand U11503 (N_11503,N_11257,N_11279);
nand U11504 (N_11504,N_11311,N_11391);
xor U11505 (N_11505,N_11218,N_11279);
nand U11506 (N_11506,N_11389,N_11216);
nor U11507 (N_11507,N_11256,N_11364);
and U11508 (N_11508,N_11227,N_11305);
or U11509 (N_11509,N_11212,N_11296);
or U11510 (N_11510,N_11212,N_11276);
nor U11511 (N_11511,N_11330,N_11265);
or U11512 (N_11512,N_11315,N_11376);
and U11513 (N_11513,N_11396,N_11326);
nor U11514 (N_11514,N_11264,N_11362);
or U11515 (N_11515,N_11279,N_11375);
and U11516 (N_11516,N_11339,N_11211);
nand U11517 (N_11517,N_11309,N_11347);
nand U11518 (N_11518,N_11271,N_11386);
nor U11519 (N_11519,N_11255,N_11329);
or U11520 (N_11520,N_11254,N_11274);
and U11521 (N_11521,N_11342,N_11211);
or U11522 (N_11522,N_11326,N_11397);
and U11523 (N_11523,N_11210,N_11225);
nor U11524 (N_11524,N_11328,N_11237);
and U11525 (N_11525,N_11222,N_11338);
or U11526 (N_11526,N_11263,N_11290);
or U11527 (N_11527,N_11332,N_11302);
nor U11528 (N_11528,N_11319,N_11232);
xnor U11529 (N_11529,N_11307,N_11205);
nor U11530 (N_11530,N_11329,N_11285);
or U11531 (N_11531,N_11295,N_11271);
or U11532 (N_11532,N_11207,N_11397);
nand U11533 (N_11533,N_11380,N_11213);
nor U11534 (N_11534,N_11256,N_11338);
or U11535 (N_11535,N_11277,N_11347);
or U11536 (N_11536,N_11352,N_11297);
and U11537 (N_11537,N_11275,N_11209);
nor U11538 (N_11538,N_11320,N_11369);
and U11539 (N_11539,N_11264,N_11271);
or U11540 (N_11540,N_11314,N_11294);
nor U11541 (N_11541,N_11349,N_11236);
nor U11542 (N_11542,N_11388,N_11340);
xnor U11543 (N_11543,N_11207,N_11372);
nand U11544 (N_11544,N_11338,N_11233);
or U11545 (N_11545,N_11380,N_11324);
nor U11546 (N_11546,N_11357,N_11319);
and U11547 (N_11547,N_11367,N_11379);
nand U11548 (N_11548,N_11273,N_11258);
and U11549 (N_11549,N_11356,N_11369);
and U11550 (N_11550,N_11332,N_11254);
or U11551 (N_11551,N_11306,N_11262);
and U11552 (N_11552,N_11360,N_11287);
or U11553 (N_11553,N_11323,N_11240);
or U11554 (N_11554,N_11247,N_11392);
or U11555 (N_11555,N_11215,N_11253);
nand U11556 (N_11556,N_11234,N_11305);
or U11557 (N_11557,N_11203,N_11278);
nor U11558 (N_11558,N_11393,N_11386);
nor U11559 (N_11559,N_11334,N_11257);
nor U11560 (N_11560,N_11284,N_11309);
or U11561 (N_11561,N_11297,N_11295);
nor U11562 (N_11562,N_11352,N_11343);
and U11563 (N_11563,N_11213,N_11229);
nand U11564 (N_11564,N_11323,N_11228);
or U11565 (N_11565,N_11241,N_11254);
nor U11566 (N_11566,N_11213,N_11338);
nor U11567 (N_11567,N_11322,N_11234);
nor U11568 (N_11568,N_11320,N_11247);
or U11569 (N_11569,N_11387,N_11343);
and U11570 (N_11570,N_11399,N_11385);
nand U11571 (N_11571,N_11317,N_11261);
xnor U11572 (N_11572,N_11210,N_11343);
and U11573 (N_11573,N_11201,N_11204);
or U11574 (N_11574,N_11209,N_11362);
and U11575 (N_11575,N_11237,N_11228);
nand U11576 (N_11576,N_11386,N_11295);
or U11577 (N_11577,N_11301,N_11354);
and U11578 (N_11578,N_11214,N_11308);
nor U11579 (N_11579,N_11355,N_11345);
nor U11580 (N_11580,N_11360,N_11300);
nand U11581 (N_11581,N_11273,N_11267);
nand U11582 (N_11582,N_11379,N_11243);
or U11583 (N_11583,N_11266,N_11269);
and U11584 (N_11584,N_11386,N_11353);
nand U11585 (N_11585,N_11330,N_11203);
or U11586 (N_11586,N_11370,N_11357);
and U11587 (N_11587,N_11284,N_11251);
nor U11588 (N_11588,N_11233,N_11344);
nor U11589 (N_11589,N_11230,N_11341);
and U11590 (N_11590,N_11396,N_11379);
nor U11591 (N_11591,N_11326,N_11318);
or U11592 (N_11592,N_11243,N_11232);
nor U11593 (N_11593,N_11343,N_11257);
nand U11594 (N_11594,N_11309,N_11250);
xor U11595 (N_11595,N_11215,N_11234);
or U11596 (N_11596,N_11341,N_11265);
nor U11597 (N_11597,N_11296,N_11213);
or U11598 (N_11598,N_11220,N_11384);
nor U11599 (N_11599,N_11207,N_11278);
or U11600 (N_11600,N_11579,N_11401);
or U11601 (N_11601,N_11531,N_11416);
or U11602 (N_11602,N_11493,N_11452);
or U11603 (N_11603,N_11571,N_11422);
or U11604 (N_11604,N_11428,N_11582);
nor U11605 (N_11605,N_11457,N_11491);
nor U11606 (N_11606,N_11554,N_11507);
nand U11607 (N_11607,N_11541,N_11408);
and U11608 (N_11608,N_11536,N_11477);
xor U11609 (N_11609,N_11538,N_11566);
and U11610 (N_11610,N_11503,N_11470);
or U11611 (N_11611,N_11599,N_11504);
or U11612 (N_11612,N_11456,N_11551);
nand U11613 (N_11613,N_11447,N_11440);
and U11614 (N_11614,N_11468,N_11596);
and U11615 (N_11615,N_11437,N_11450);
xor U11616 (N_11616,N_11574,N_11515);
xor U11617 (N_11617,N_11523,N_11542);
nand U11618 (N_11618,N_11407,N_11451);
or U11619 (N_11619,N_11575,N_11402);
xnor U11620 (N_11620,N_11587,N_11500);
nor U11621 (N_11621,N_11425,N_11563);
nand U11622 (N_11622,N_11537,N_11584);
xnor U11623 (N_11623,N_11530,N_11589);
or U11624 (N_11624,N_11454,N_11521);
and U11625 (N_11625,N_11446,N_11486);
nand U11626 (N_11626,N_11592,N_11558);
or U11627 (N_11627,N_11580,N_11476);
nor U11628 (N_11628,N_11581,N_11540);
xnor U11629 (N_11629,N_11525,N_11427);
and U11630 (N_11630,N_11505,N_11502);
and U11631 (N_11631,N_11562,N_11565);
nand U11632 (N_11632,N_11495,N_11412);
and U11633 (N_11633,N_11522,N_11552);
nor U11634 (N_11634,N_11550,N_11460);
xnor U11635 (N_11635,N_11473,N_11547);
or U11636 (N_11636,N_11442,N_11479);
or U11637 (N_11637,N_11519,N_11585);
nor U11638 (N_11638,N_11480,N_11561);
or U11639 (N_11639,N_11438,N_11484);
nor U11640 (N_11640,N_11597,N_11458);
nand U11641 (N_11641,N_11489,N_11508);
or U11642 (N_11642,N_11475,N_11492);
nor U11643 (N_11643,N_11570,N_11573);
or U11644 (N_11644,N_11429,N_11462);
and U11645 (N_11645,N_11514,N_11430);
nand U11646 (N_11646,N_11595,N_11481);
nand U11647 (N_11647,N_11545,N_11411);
or U11648 (N_11648,N_11487,N_11439);
nor U11649 (N_11649,N_11516,N_11586);
nand U11650 (N_11650,N_11583,N_11449);
and U11651 (N_11651,N_11443,N_11555);
nand U11652 (N_11652,N_11418,N_11461);
and U11653 (N_11653,N_11403,N_11572);
nand U11654 (N_11654,N_11578,N_11472);
and U11655 (N_11655,N_11478,N_11529);
nor U11656 (N_11656,N_11512,N_11445);
and U11657 (N_11657,N_11534,N_11497);
nor U11658 (N_11658,N_11432,N_11567);
xor U11659 (N_11659,N_11419,N_11517);
or U11660 (N_11660,N_11501,N_11448);
nand U11661 (N_11661,N_11406,N_11436);
or U11662 (N_11662,N_11494,N_11420);
nor U11663 (N_11663,N_11509,N_11421);
nor U11664 (N_11664,N_11576,N_11482);
or U11665 (N_11665,N_11539,N_11593);
or U11666 (N_11666,N_11548,N_11474);
nand U11667 (N_11667,N_11455,N_11498);
nor U11668 (N_11668,N_11591,N_11533);
nor U11669 (N_11669,N_11535,N_11490);
nand U11670 (N_11670,N_11471,N_11417);
nor U11671 (N_11671,N_11485,N_11549);
nand U11672 (N_11672,N_11496,N_11559);
or U11673 (N_11673,N_11441,N_11409);
xnor U11674 (N_11674,N_11444,N_11415);
xnor U11675 (N_11675,N_11590,N_11528);
or U11676 (N_11676,N_11543,N_11598);
xor U11677 (N_11677,N_11518,N_11553);
or U11678 (N_11678,N_11499,N_11511);
nand U11679 (N_11679,N_11594,N_11465);
or U11680 (N_11680,N_11544,N_11426);
and U11681 (N_11681,N_11424,N_11467);
nand U11682 (N_11682,N_11459,N_11560);
xnor U11683 (N_11683,N_11404,N_11588);
and U11684 (N_11684,N_11520,N_11556);
or U11685 (N_11685,N_11414,N_11513);
or U11686 (N_11686,N_11463,N_11510);
nor U11687 (N_11687,N_11568,N_11577);
xnor U11688 (N_11688,N_11423,N_11433);
and U11689 (N_11689,N_11400,N_11526);
and U11690 (N_11690,N_11434,N_11564);
and U11691 (N_11691,N_11435,N_11410);
and U11692 (N_11692,N_11532,N_11527);
and U11693 (N_11693,N_11488,N_11431);
and U11694 (N_11694,N_11405,N_11546);
or U11695 (N_11695,N_11524,N_11483);
nand U11696 (N_11696,N_11466,N_11469);
nor U11697 (N_11697,N_11569,N_11413);
nand U11698 (N_11698,N_11453,N_11557);
nor U11699 (N_11699,N_11464,N_11506);
nor U11700 (N_11700,N_11592,N_11483);
nor U11701 (N_11701,N_11549,N_11566);
nor U11702 (N_11702,N_11587,N_11524);
nor U11703 (N_11703,N_11467,N_11540);
nor U11704 (N_11704,N_11586,N_11517);
nor U11705 (N_11705,N_11551,N_11532);
or U11706 (N_11706,N_11517,N_11583);
and U11707 (N_11707,N_11592,N_11498);
or U11708 (N_11708,N_11478,N_11548);
nand U11709 (N_11709,N_11420,N_11552);
or U11710 (N_11710,N_11477,N_11508);
xnor U11711 (N_11711,N_11590,N_11405);
nor U11712 (N_11712,N_11400,N_11462);
nand U11713 (N_11713,N_11449,N_11470);
nand U11714 (N_11714,N_11484,N_11571);
nor U11715 (N_11715,N_11425,N_11505);
and U11716 (N_11716,N_11592,N_11490);
nor U11717 (N_11717,N_11523,N_11555);
xor U11718 (N_11718,N_11440,N_11485);
nor U11719 (N_11719,N_11548,N_11528);
nand U11720 (N_11720,N_11563,N_11592);
or U11721 (N_11721,N_11518,N_11567);
and U11722 (N_11722,N_11401,N_11448);
xor U11723 (N_11723,N_11502,N_11560);
nor U11724 (N_11724,N_11503,N_11528);
nor U11725 (N_11725,N_11578,N_11504);
nand U11726 (N_11726,N_11576,N_11544);
nand U11727 (N_11727,N_11550,N_11440);
xnor U11728 (N_11728,N_11503,N_11475);
xnor U11729 (N_11729,N_11442,N_11448);
nand U11730 (N_11730,N_11488,N_11575);
nand U11731 (N_11731,N_11518,N_11586);
or U11732 (N_11732,N_11426,N_11434);
nand U11733 (N_11733,N_11454,N_11582);
and U11734 (N_11734,N_11520,N_11476);
nand U11735 (N_11735,N_11597,N_11431);
or U11736 (N_11736,N_11488,N_11430);
nand U11737 (N_11737,N_11406,N_11484);
nor U11738 (N_11738,N_11430,N_11476);
or U11739 (N_11739,N_11428,N_11469);
or U11740 (N_11740,N_11460,N_11576);
xor U11741 (N_11741,N_11500,N_11454);
or U11742 (N_11742,N_11470,N_11516);
and U11743 (N_11743,N_11594,N_11562);
and U11744 (N_11744,N_11578,N_11413);
nor U11745 (N_11745,N_11528,N_11498);
or U11746 (N_11746,N_11592,N_11494);
nand U11747 (N_11747,N_11499,N_11487);
nand U11748 (N_11748,N_11449,N_11557);
xor U11749 (N_11749,N_11567,N_11413);
xor U11750 (N_11750,N_11400,N_11421);
nor U11751 (N_11751,N_11576,N_11435);
xnor U11752 (N_11752,N_11462,N_11547);
nand U11753 (N_11753,N_11453,N_11444);
nand U11754 (N_11754,N_11417,N_11490);
nor U11755 (N_11755,N_11545,N_11447);
or U11756 (N_11756,N_11534,N_11574);
or U11757 (N_11757,N_11401,N_11558);
nand U11758 (N_11758,N_11436,N_11460);
and U11759 (N_11759,N_11515,N_11408);
nand U11760 (N_11760,N_11457,N_11484);
or U11761 (N_11761,N_11437,N_11571);
or U11762 (N_11762,N_11444,N_11426);
nor U11763 (N_11763,N_11499,N_11573);
and U11764 (N_11764,N_11538,N_11470);
nor U11765 (N_11765,N_11474,N_11523);
nor U11766 (N_11766,N_11488,N_11554);
and U11767 (N_11767,N_11420,N_11461);
xnor U11768 (N_11768,N_11561,N_11586);
and U11769 (N_11769,N_11485,N_11517);
nand U11770 (N_11770,N_11578,N_11570);
and U11771 (N_11771,N_11464,N_11599);
nand U11772 (N_11772,N_11408,N_11516);
or U11773 (N_11773,N_11430,N_11535);
xor U11774 (N_11774,N_11532,N_11429);
or U11775 (N_11775,N_11595,N_11456);
nor U11776 (N_11776,N_11506,N_11476);
and U11777 (N_11777,N_11550,N_11552);
nand U11778 (N_11778,N_11513,N_11537);
xnor U11779 (N_11779,N_11537,N_11472);
xor U11780 (N_11780,N_11544,N_11560);
nor U11781 (N_11781,N_11428,N_11476);
nor U11782 (N_11782,N_11532,N_11522);
xor U11783 (N_11783,N_11466,N_11580);
nand U11784 (N_11784,N_11447,N_11459);
xnor U11785 (N_11785,N_11448,N_11578);
or U11786 (N_11786,N_11470,N_11454);
nand U11787 (N_11787,N_11522,N_11476);
and U11788 (N_11788,N_11496,N_11435);
nand U11789 (N_11789,N_11592,N_11458);
or U11790 (N_11790,N_11403,N_11469);
xor U11791 (N_11791,N_11409,N_11566);
and U11792 (N_11792,N_11594,N_11514);
or U11793 (N_11793,N_11558,N_11452);
xnor U11794 (N_11794,N_11402,N_11583);
or U11795 (N_11795,N_11535,N_11512);
and U11796 (N_11796,N_11463,N_11438);
nand U11797 (N_11797,N_11440,N_11572);
nor U11798 (N_11798,N_11573,N_11433);
nor U11799 (N_11799,N_11499,N_11405);
nand U11800 (N_11800,N_11616,N_11614);
xnor U11801 (N_11801,N_11755,N_11785);
and U11802 (N_11802,N_11753,N_11776);
nand U11803 (N_11803,N_11612,N_11771);
or U11804 (N_11804,N_11726,N_11627);
nand U11805 (N_11805,N_11672,N_11754);
nand U11806 (N_11806,N_11784,N_11604);
nand U11807 (N_11807,N_11611,N_11671);
or U11808 (N_11808,N_11623,N_11622);
or U11809 (N_11809,N_11643,N_11648);
xnor U11810 (N_11810,N_11781,N_11798);
nand U11811 (N_11811,N_11710,N_11630);
and U11812 (N_11812,N_11675,N_11748);
nand U11813 (N_11813,N_11724,N_11795);
and U11814 (N_11814,N_11751,N_11769);
and U11815 (N_11815,N_11716,N_11609);
or U11816 (N_11816,N_11629,N_11693);
and U11817 (N_11817,N_11688,N_11796);
or U11818 (N_11818,N_11793,N_11750);
or U11819 (N_11819,N_11770,N_11686);
nand U11820 (N_11820,N_11735,N_11658);
or U11821 (N_11821,N_11676,N_11737);
nand U11822 (N_11822,N_11783,N_11677);
and U11823 (N_11823,N_11764,N_11746);
nor U11824 (N_11824,N_11702,N_11624);
nor U11825 (N_11825,N_11666,N_11720);
or U11826 (N_11826,N_11778,N_11664);
and U11827 (N_11827,N_11714,N_11767);
or U11828 (N_11828,N_11628,N_11617);
xor U11829 (N_11829,N_11749,N_11739);
nor U11830 (N_11830,N_11696,N_11773);
or U11831 (N_11831,N_11745,N_11657);
nor U11832 (N_11832,N_11794,N_11670);
nor U11833 (N_11833,N_11621,N_11752);
or U11834 (N_11834,N_11756,N_11734);
nor U11835 (N_11835,N_11690,N_11711);
or U11836 (N_11836,N_11650,N_11790);
or U11837 (N_11837,N_11717,N_11636);
and U11838 (N_11838,N_11642,N_11603);
nor U11839 (N_11839,N_11681,N_11774);
and U11840 (N_11840,N_11740,N_11639);
or U11841 (N_11841,N_11730,N_11652);
nor U11842 (N_11842,N_11626,N_11674);
or U11843 (N_11843,N_11610,N_11731);
or U11844 (N_11844,N_11760,N_11718);
xnor U11845 (N_11845,N_11728,N_11685);
nor U11846 (N_11846,N_11691,N_11655);
xnor U11847 (N_11847,N_11600,N_11659);
or U11848 (N_11848,N_11665,N_11692);
and U11849 (N_11849,N_11641,N_11732);
nor U11850 (N_11850,N_11741,N_11687);
xor U11851 (N_11851,N_11683,N_11680);
and U11852 (N_11852,N_11761,N_11789);
or U11853 (N_11853,N_11743,N_11775);
or U11854 (N_11854,N_11763,N_11721);
or U11855 (N_11855,N_11608,N_11733);
and U11856 (N_11856,N_11679,N_11701);
nand U11857 (N_11857,N_11765,N_11619);
and U11858 (N_11858,N_11637,N_11613);
nor U11859 (N_11859,N_11644,N_11725);
nand U11860 (N_11860,N_11601,N_11631);
or U11861 (N_11861,N_11780,N_11708);
or U11862 (N_11862,N_11649,N_11712);
and U11863 (N_11863,N_11606,N_11668);
nor U11864 (N_11864,N_11633,N_11736);
nand U11865 (N_11865,N_11620,N_11719);
nand U11866 (N_11866,N_11615,N_11722);
or U11867 (N_11867,N_11766,N_11705);
nor U11868 (N_11868,N_11747,N_11667);
nand U11869 (N_11869,N_11707,N_11738);
nand U11870 (N_11870,N_11786,N_11713);
nand U11871 (N_11871,N_11787,N_11646);
and U11872 (N_11872,N_11715,N_11704);
nand U11873 (N_11873,N_11634,N_11792);
and U11874 (N_11874,N_11654,N_11723);
nor U11875 (N_11875,N_11703,N_11799);
nand U11876 (N_11876,N_11684,N_11660);
and U11877 (N_11877,N_11673,N_11699);
nand U11878 (N_11878,N_11694,N_11663);
nand U11879 (N_11879,N_11653,N_11706);
nand U11880 (N_11880,N_11662,N_11682);
or U11881 (N_11881,N_11788,N_11640);
or U11882 (N_11882,N_11638,N_11645);
xor U11883 (N_11883,N_11758,N_11772);
nand U11884 (N_11884,N_11625,N_11762);
or U11885 (N_11885,N_11777,N_11727);
or U11886 (N_11886,N_11782,N_11709);
or U11887 (N_11887,N_11651,N_11744);
xnor U11888 (N_11888,N_11768,N_11759);
nor U11889 (N_11889,N_11656,N_11698);
and U11890 (N_11890,N_11607,N_11695);
nor U11891 (N_11891,N_11779,N_11602);
or U11892 (N_11892,N_11689,N_11605);
and U11893 (N_11893,N_11742,N_11635);
or U11894 (N_11894,N_11669,N_11661);
nand U11895 (N_11895,N_11700,N_11678);
nand U11896 (N_11896,N_11797,N_11647);
nand U11897 (N_11897,N_11729,N_11632);
or U11898 (N_11898,N_11618,N_11697);
nand U11899 (N_11899,N_11757,N_11791);
nor U11900 (N_11900,N_11759,N_11776);
and U11901 (N_11901,N_11689,N_11772);
and U11902 (N_11902,N_11671,N_11693);
xor U11903 (N_11903,N_11720,N_11648);
or U11904 (N_11904,N_11665,N_11617);
nor U11905 (N_11905,N_11672,N_11799);
or U11906 (N_11906,N_11661,N_11773);
nor U11907 (N_11907,N_11671,N_11632);
or U11908 (N_11908,N_11647,N_11715);
nand U11909 (N_11909,N_11625,N_11676);
or U11910 (N_11910,N_11687,N_11693);
nand U11911 (N_11911,N_11717,N_11794);
nor U11912 (N_11912,N_11678,N_11732);
nor U11913 (N_11913,N_11724,N_11684);
and U11914 (N_11914,N_11792,N_11603);
and U11915 (N_11915,N_11798,N_11659);
and U11916 (N_11916,N_11688,N_11706);
nand U11917 (N_11917,N_11707,N_11637);
and U11918 (N_11918,N_11649,N_11786);
and U11919 (N_11919,N_11602,N_11700);
and U11920 (N_11920,N_11708,N_11649);
nor U11921 (N_11921,N_11672,N_11629);
or U11922 (N_11922,N_11648,N_11662);
or U11923 (N_11923,N_11670,N_11734);
or U11924 (N_11924,N_11600,N_11708);
or U11925 (N_11925,N_11756,N_11724);
xnor U11926 (N_11926,N_11758,N_11655);
and U11927 (N_11927,N_11671,N_11787);
or U11928 (N_11928,N_11655,N_11674);
or U11929 (N_11929,N_11702,N_11792);
xor U11930 (N_11930,N_11671,N_11757);
nor U11931 (N_11931,N_11627,N_11654);
xor U11932 (N_11932,N_11615,N_11619);
or U11933 (N_11933,N_11645,N_11699);
and U11934 (N_11934,N_11645,N_11620);
nor U11935 (N_11935,N_11736,N_11659);
nor U11936 (N_11936,N_11718,N_11677);
or U11937 (N_11937,N_11715,N_11770);
nor U11938 (N_11938,N_11734,N_11678);
or U11939 (N_11939,N_11629,N_11785);
nand U11940 (N_11940,N_11624,N_11705);
and U11941 (N_11941,N_11652,N_11720);
and U11942 (N_11942,N_11760,N_11780);
or U11943 (N_11943,N_11700,N_11778);
or U11944 (N_11944,N_11669,N_11691);
xnor U11945 (N_11945,N_11783,N_11621);
nand U11946 (N_11946,N_11748,N_11789);
nand U11947 (N_11947,N_11767,N_11646);
or U11948 (N_11948,N_11792,N_11795);
nor U11949 (N_11949,N_11709,N_11621);
nand U11950 (N_11950,N_11781,N_11652);
nor U11951 (N_11951,N_11699,N_11799);
and U11952 (N_11952,N_11678,N_11719);
xor U11953 (N_11953,N_11671,N_11656);
and U11954 (N_11954,N_11691,N_11766);
or U11955 (N_11955,N_11692,N_11756);
or U11956 (N_11956,N_11793,N_11748);
xnor U11957 (N_11957,N_11719,N_11791);
nand U11958 (N_11958,N_11688,N_11674);
xor U11959 (N_11959,N_11648,N_11795);
and U11960 (N_11960,N_11637,N_11671);
or U11961 (N_11961,N_11773,N_11666);
xor U11962 (N_11962,N_11710,N_11662);
nand U11963 (N_11963,N_11785,N_11681);
nand U11964 (N_11964,N_11721,N_11754);
nand U11965 (N_11965,N_11633,N_11798);
and U11966 (N_11966,N_11651,N_11608);
nand U11967 (N_11967,N_11606,N_11783);
nand U11968 (N_11968,N_11793,N_11731);
nand U11969 (N_11969,N_11645,N_11713);
nand U11970 (N_11970,N_11754,N_11770);
nand U11971 (N_11971,N_11628,N_11735);
and U11972 (N_11972,N_11671,N_11630);
nand U11973 (N_11973,N_11602,N_11603);
and U11974 (N_11974,N_11778,N_11658);
or U11975 (N_11975,N_11688,N_11658);
nor U11976 (N_11976,N_11608,N_11751);
nor U11977 (N_11977,N_11725,N_11611);
and U11978 (N_11978,N_11776,N_11614);
nand U11979 (N_11979,N_11798,N_11696);
and U11980 (N_11980,N_11630,N_11698);
nor U11981 (N_11981,N_11613,N_11787);
nand U11982 (N_11982,N_11743,N_11739);
or U11983 (N_11983,N_11786,N_11670);
or U11984 (N_11984,N_11734,N_11620);
and U11985 (N_11985,N_11762,N_11786);
or U11986 (N_11986,N_11655,N_11756);
xnor U11987 (N_11987,N_11630,N_11605);
nand U11988 (N_11988,N_11692,N_11786);
or U11989 (N_11989,N_11705,N_11769);
nor U11990 (N_11990,N_11770,N_11697);
xnor U11991 (N_11991,N_11676,N_11613);
nand U11992 (N_11992,N_11661,N_11671);
nand U11993 (N_11993,N_11737,N_11668);
nor U11994 (N_11994,N_11672,N_11689);
or U11995 (N_11995,N_11724,N_11773);
nand U11996 (N_11996,N_11760,N_11733);
xnor U11997 (N_11997,N_11649,N_11691);
nand U11998 (N_11998,N_11659,N_11648);
nand U11999 (N_11999,N_11696,N_11776);
nor U12000 (N_12000,N_11911,N_11922);
nor U12001 (N_12001,N_11865,N_11900);
nand U12002 (N_12002,N_11830,N_11808);
nand U12003 (N_12003,N_11973,N_11864);
xnor U12004 (N_12004,N_11915,N_11807);
and U12005 (N_12005,N_11932,N_11925);
and U12006 (N_12006,N_11926,N_11951);
and U12007 (N_12007,N_11953,N_11941);
nand U12008 (N_12008,N_11820,N_11905);
nand U12009 (N_12009,N_11816,N_11867);
and U12010 (N_12010,N_11938,N_11800);
nor U12011 (N_12011,N_11838,N_11997);
nand U12012 (N_12012,N_11980,N_11892);
nand U12013 (N_12013,N_11948,N_11921);
xnor U12014 (N_12014,N_11869,N_11904);
nand U12015 (N_12015,N_11883,N_11914);
nor U12016 (N_12016,N_11918,N_11955);
and U12017 (N_12017,N_11977,N_11887);
nand U12018 (N_12018,N_11861,N_11821);
and U12019 (N_12019,N_11964,N_11875);
or U12020 (N_12020,N_11959,N_11809);
nand U12021 (N_12021,N_11814,N_11802);
or U12022 (N_12022,N_11901,N_11913);
or U12023 (N_12023,N_11954,N_11939);
nand U12024 (N_12024,N_11972,N_11920);
nor U12025 (N_12025,N_11849,N_11858);
nand U12026 (N_12026,N_11813,N_11819);
nand U12027 (N_12027,N_11854,N_11818);
and U12028 (N_12028,N_11855,N_11804);
nor U12029 (N_12029,N_11945,N_11963);
nor U12030 (N_12030,N_11936,N_11958);
xor U12031 (N_12031,N_11898,N_11880);
xnor U12032 (N_12032,N_11896,N_11975);
nor U12033 (N_12033,N_11886,N_11851);
nand U12034 (N_12034,N_11903,N_11873);
nor U12035 (N_12035,N_11840,N_11987);
nor U12036 (N_12036,N_11871,N_11970);
nand U12037 (N_12037,N_11872,N_11862);
and U12038 (N_12038,N_11989,N_11908);
or U12039 (N_12039,N_11811,N_11995);
nor U12040 (N_12040,N_11931,N_11877);
xnor U12041 (N_12041,N_11823,N_11923);
or U12042 (N_12042,N_11965,N_11952);
nor U12043 (N_12043,N_11993,N_11859);
nor U12044 (N_12044,N_11888,N_11950);
nor U12045 (N_12045,N_11996,N_11839);
nor U12046 (N_12046,N_11897,N_11909);
or U12047 (N_12047,N_11876,N_11826);
nor U12048 (N_12048,N_11836,N_11890);
nand U12049 (N_12049,N_11917,N_11815);
nand U12050 (N_12050,N_11962,N_11837);
and U12051 (N_12051,N_11860,N_11934);
nand U12052 (N_12052,N_11899,N_11998);
nand U12053 (N_12053,N_11831,N_11805);
nor U12054 (N_12054,N_11878,N_11933);
nand U12055 (N_12055,N_11969,N_11848);
nor U12056 (N_12056,N_11866,N_11912);
nand U12057 (N_12057,N_11884,N_11919);
and U12058 (N_12058,N_11979,N_11885);
nand U12059 (N_12059,N_11806,N_11895);
and U12060 (N_12060,N_11874,N_11845);
nor U12061 (N_12061,N_11927,N_11961);
xor U12062 (N_12062,N_11990,N_11852);
nand U12063 (N_12063,N_11832,N_11985);
or U12064 (N_12064,N_11981,N_11930);
nor U12065 (N_12065,N_11846,N_11827);
and U12066 (N_12066,N_11928,N_11956);
nand U12067 (N_12067,N_11902,N_11894);
and U12068 (N_12068,N_11944,N_11817);
nor U12069 (N_12069,N_11803,N_11863);
and U12070 (N_12070,N_11957,N_11882);
nand U12071 (N_12071,N_11850,N_11968);
nor U12072 (N_12072,N_11976,N_11935);
xnor U12073 (N_12073,N_11893,N_11889);
or U12074 (N_12074,N_11828,N_11916);
and U12075 (N_12075,N_11966,N_11857);
or U12076 (N_12076,N_11801,N_11824);
nor U12077 (N_12077,N_11999,N_11835);
and U12078 (N_12078,N_11943,N_11856);
or U12079 (N_12079,N_11906,N_11910);
nand U12080 (N_12080,N_11988,N_11822);
or U12081 (N_12081,N_11924,N_11971);
or U12082 (N_12082,N_11994,N_11974);
or U12083 (N_12083,N_11870,N_11991);
and U12084 (N_12084,N_11937,N_11984);
nor U12085 (N_12085,N_11829,N_11812);
nand U12086 (N_12086,N_11978,N_11940);
or U12087 (N_12087,N_11844,N_11907);
nor U12088 (N_12088,N_11983,N_11929);
xnor U12089 (N_12089,N_11853,N_11842);
nand U12090 (N_12090,N_11982,N_11841);
or U12091 (N_12091,N_11847,N_11942);
nand U12092 (N_12092,N_11833,N_11881);
and U12093 (N_12093,N_11986,N_11967);
nor U12094 (N_12094,N_11992,N_11947);
nand U12095 (N_12095,N_11843,N_11834);
and U12096 (N_12096,N_11810,N_11960);
or U12097 (N_12097,N_11946,N_11891);
or U12098 (N_12098,N_11879,N_11868);
xnor U12099 (N_12099,N_11949,N_11825);
nand U12100 (N_12100,N_11876,N_11837);
nand U12101 (N_12101,N_11834,N_11902);
and U12102 (N_12102,N_11974,N_11848);
or U12103 (N_12103,N_11895,N_11918);
xnor U12104 (N_12104,N_11967,N_11815);
xor U12105 (N_12105,N_11810,N_11844);
nor U12106 (N_12106,N_11999,N_11955);
nor U12107 (N_12107,N_11975,N_11925);
and U12108 (N_12108,N_11971,N_11862);
xor U12109 (N_12109,N_11889,N_11813);
xnor U12110 (N_12110,N_11932,N_11905);
nor U12111 (N_12111,N_11956,N_11824);
and U12112 (N_12112,N_11876,N_11888);
or U12113 (N_12113,N_11946,N_11840);
and U12114 (N_12114,N_11909,N_11801);
or U12115 (N_12115,N_11937,N_11805);
or U12116 (N_12116,N_11834,N_11911);
nor U12117 (N_12117,N_11894,N_11940);
or U12118 (N_12118,N_11807,N_11844);
and U12119 (N_12119,N_11821,N_11889);
nand U12120 (N_12120,N_11909,N_11891);
or U12121 (N_12121,N_11813,N_11890);
or U12122 (N_12122,N_11905,N_11924);
or U12123 (N_12123,N_11964,N_11929);
nand U12124 (N_12124,N_11805,N_11827);
nor U12125 (N_12125,N_11843,N_11897);
or U12126 (N_12126,N_11830,N_11849);
or U12127 (N_12127,N_11901,N_11811);
and U12128 (N_12128,N_11867,N_11977);
nand U12129 (N_12129,N_11947,N_11959);
and U12130 (N_12130,N_11902,N_11945);
or U12131 (N_12131,N_11828,N_11817);
or U12132 (N_12132,N_11802,N_11936);
or U12133 (N_12133,N_11881,N_11859);
or U12134 (N_12134,N_11887,N_11862);
nand U12135 (N_12135,N_11806,N_11908);
and U12136 (N_12136,N_11937,N_11845);
and U12137 (N_12137,N_11920,N_11988);
or U12138 (N_12138,N_11896,N_11907);
nand U12139 (N_12139,N_11848,N_11817);
xnor U12140 (N_12140,N_11814,N_11855);
nand U12141 (N_12141,N_11869,N_11976);
nand U12142 (N_12142,N_11879,N_11928);
nor U12143 (N_12143,N_11883,N_11989);
nand U12144 (N_12144,N_11994,N_11982);
and U12145 (N_12145,N_11898,N_11913);
nor U12146 (N_12146,N_11939,N_11865);
or U12147 (N_12147,N_11915,N_11809);
nor U12148 (N_12148,N_11858,N_11944);
xnor U12149 (N_12149,N_11837,N_11948);
nand U12150 (N_12150,N_11844,N_11840);
nor U12151 (N_12151,N_11820,N_11938);
nor U12152 (N_12152,N_11986,N_11873);
nand U12153 (N_12153,N_11988,N_11842);
nand U12154 (N_12154,N_11821,N_11991);
nand U12155 (N_12155,N_11994,N_11902);
nand U12156 (N_12156,N_11870,N_11867);
or U12157 (N_12157,N_11928,N_11930);
nor U12158 (N_12158,N_11858,N_11884);
nor U12159 (N_12159,N_11810,N_11893);
and U12160 (N_12160,N_11820,N_11914);
or U12161 (N_12161,N_11871,N_11879);
or U12162 (N_12162,N_11945,N_11983);
nor U12163 (N_12163,N_11839,N_11835);
nor U12164 (N_12164,N_11846,N_11859);
and U12165 (N_12165,N_11832,N_11838);
xnor U12166 (N_12166,N_11818,N_11872);
nor U12167 (N_12167,N_11959,N_11875);
and U12168 (N_12168,N_11928,N_11924);
nor U12169 (N_12169,N_11820,N_11869);
or U12170 (N_12170,N_11914,N_11855);
or U12171 (N_12171,N_11871,N_11976);
nor U12172 (N_12172,N_11960,N_11827);
or U12173 (N_12173,N_11861,N_11907);
nand U12174 (N_12174,N_11898,N_11960);
and U12175 (N_12175,N_11907,N_11865);
nor U12176 (N_12176,N_11932,N_11803);
nand U12177 (N_12177,N_11873,N_11845);
or U12178 (N_12178,N_11804,N_11873);
nand U12179 (N_12179,N_11944,N_11929);
or U12180 (N_12180,N_11885,N_11874);
and U12181 (N_12181,N_11972,N_11870);
and U12182 (N_12182,N_11920,N_11983);
xor U12183 (N_12183,N_11975,N_11848);
nor U12184 (N_12184,N_11812,N_11917);
or U12185 (N_12185,N_11850,N_11980);
or U12186 (N_12186,N_11916,N_11800);
or U12187 (N_12187,N_11967,N_11877);
nand U12188 (N_12188,N_11949,N_11829);
nor U12189 (N_12189,N_11801,N_11968);
nor U12190 (N_12190,N_11818,N_11920);
or U12191 (N_12191,N_11957,N_11894);
nand U12192 (N_12192,N_11846,N_11864);
nand U12193 (N_12193,N_11880,N_11895);
nor U12194 (N_12194,N_11936,N_11925);
nand U12195 (N_12195,N_11897,N_11893);
xnor U12196 (N_12196,N_11906,N_11809);
or U12197 (N_12197,N_11828,N_11866);
nand U12198 (N_12198,N_11994,N_11943);
or U12199 (N_12199,N_11979,N_11880);
or U12200 (N_12200,N_12167,N_12190);
or U12201 (N_12201,N_12094,N_12077);
nand U12202 (N_12202,N_12090,N_12041);
or U12203 (N_12203,N_12115,N_12089);
and U12204 (N_12204,N_12174,N_12079);
nand U12205 (N_12205,N_12178,N_12035);
and U12206 (N_12206,N_12019,N_12160);
and U12207 (N_12207,N_12068,N_12112);
or U12208 (N_12208,N_12165,N_12063);
nor U12209 (N_12209,N_12100,N_12097);
nor U12210 (N_12210,N_12034,N_12030);
or U12211 (N_12211,N_12187,N_12168);
and U12212 (N_12212,N_12101,N_12136);
nor U12213 (N_12213,N_12051,N_12109);
nand U12214 (N_12214,N_12135,N_12123);
xor U12215 (N_12215,N_12175,N_12129);
nand U12216 (N_12216,N_12042,N_12131);
or U12217 (N_12217,N_12196,N_12155);
xor U12218 (N_12218,N_12009,N_12141);
nand U12219 (N_12219,N_12182,N_12189);
nor U12220 (N_12220,N_12184,N_12173);
xor U12221 (N_12221,N_12065,N_12044);
or U12222 (N_12222,N_12134,N_12029);
nor U12223 (N_12223,N_12043,N_12006);
nor U12224 (N_12224,N_12075,N_12194);
nand U12225 (N_12225,N_12003,N_12085);
xor U12226 (N_12226,N_12152,N_12110);
nor U12227 (N_12227,N_12002,N_12053);
or U12228 (N_12228,N_12171,N_12073);
or U12229 (N_12229,N_12143,N_12142);
nor U12230 (N_12230,N_12172,N_12151);
or U12231 (N_12231,N_12026,N_12170);
nor U12232 (N_12232,N_12098,N_12177);
nor U12233 (N_12233,N_12126,N_12088);
nor U12234 (N_12234,N_12074,N_12145);
nand U12235 (N_12235,N_12199,N_12137);
and U12236 (N_12236,N_12188,N_12004);
or U12237 (N_12237,N_12095,N_12133);
xnor U12238 (N_12238,N_12021,N_12010);
and U12239 (N_12239,N_12067,N_12076);
nand U12240 (N_12240,N_12001,N_12037);
and U12241 (N_12241,N_12185,N_12128);
and U12242 (N_12242,N_12124,N_12081);
nor U12243 (N_12243,N_12096,N_12122);
xor U12244 (N_12244,N_12061,N_12183);
or U12245 (N_12245,N_12139,N_12055);
and U12246 (N_12246,N_12119,N_12186);
or U12247 (N_12247,N_12058,N_12025);
nor U12248 (N_12248,N_12020,N_12092);
or U12249 (N_12249,N_12193,N_12070);
xor U12250 (N_12250,N_12080,N_12024);
nand U12251 (N_12251,N_12039,N_12031);
or U12252 (N_12252,N_12176,N_12103);
nand U12253 (N_12253,N_12011,N_12169);
nand U12254 (N_12254,N_12104,N_12147);
nor U12255 (N_12255,N_12153,N_12078);
nor U12256 (N_12256,N_12192,N_12059);
nor U12257 (N_12257,N_12052,N_12179);
nor U12258 (N_12258,N_12040,N_12140);
or U12259 (N_12259,N_12191,N_12099);
or U12260 (N_12260,N_12148,N_12164);
nand U12261 (N_12261,N_12132,N_12159);
nand U12262 (N_12262,N_12102,N_12197);
nand U12263 (N_12263,N_12195,N_12125);
and U12264 (N_12264,N_12083,N_12086);
or U12265 (N_12265,N_12036,N_12054);
nor U12266 (N_12266,N_12033,N_12007);
xor U12267 (N_12267,N_12107,N_12038);
xnor U12268 (N_12268,N_12049,N_12162);
xor U12269 (N_12269,N_12105,N_12000);
nand U12270 (N_12270,N_12013,N_12056);
and U12271 (N_12271,N_12072,N_12091);
or U12272 (N_12272,N_12113,N_12008);
nand U12273 (N_12273,N_12047,N_12028);
nand U12274 (N_12274,N_12118,N_12108);
and U12275 (N_12275,N_12015,N_12005);
or U12276 (N_12276,N_12018,N_12045);
or U12277 (N_12277,N_12014,N_12166);
nand U12278 (N_12278,N_12050,N_12027);
nor U12279 (N_12279,N_12062,N_12154);
xnor U12280 (N_12280,N_12127,N_12163);
nand U12281 (N_12281,N_12120,N_12071);
nor U12282 (N_12282,N_12017,N_12082);
nor U12283 (N_12283,N_12057,N_12111);
xnor U12284 (N_12284,N_12121,N_12161);
or U12285 (N_12285,N_12198,N_12087);
nand U12286 (N_12286,N_12060,N_12149);
or U12287 (N_12287,N_12069,N_12138);
or U12288 (N_12288,N_12023,N_12066);
or U12289 (N_12289,N_12158,N_12144);
or U12290 (N_12290,N_12156,N_12157);
nand U12291 (N_12291,N_12150,N_12130);
and U12292 (N_12292,N_12106,N_12117);
and U12293 (N_12293,N_12012,N_12084);
nor U12294 (N_12294,N_12016,N_12180);
or U12295 (N_12295,N_12116,N_12093);
nor U12296 (N_12296,N_12022,N_12181);
or U12297 (N_12297,N_12046,N_12114);
nor U12298 (N_12298,N_12032,N_12146);
and U12299 (N_12299,N_12048,N_12064);
nand U12300 (N_12300,N_12091,N_12040);
nand U12301 (N_12301,N_12185,N_12089);
nor U12302 (N_12302,N_12078,N_12141);
nand U12303 (N_12303,N_12145,N_12044);
nor U12304 (N_12304,N_12123,N_12196);
and U12305 (N_12305,N_12040,N_12162);
or U12306 (N_12306,N_12185,N_12118);
nand U12307 (N_12307,N_12183,N_12080);
nand U12308 (N_12308,N_12183,N_12129);
and U12309 (N_12309,N_12124,N_12030);
nand U12310 (N_12310,N_12195,N_12171);
or U12311 (N_12311,N_12036,N_12007);
or U12312 (N_12312,N_12035,N_12032);
and U12313 (N_12313,N_12188,N_12002);
xnor U12314 (N_12314,N_12040,N_12152);
and U12315 (N_12315,N_12035,N_12021);
nand U12316 (N_12316,N_12164,N_12162);
xor U12317 (N_12317,N_12064,N_12122);
or U12318 (N_12318,N_12128,N_12101);
nand U12319 (N_12319,N_12028,N_12051);
nor U12320 (N_12320,N_12112,N_12049);
nor U12321 (N_12321,N_12027,N_12036);
xnor U12322 (N_12322,N_12021,N_12002);
nor U12323 (N_12323,N_12101,N_12051);
nand U12324 (N_12324,N_12128,N_12166);
or U12325 (N_12325,N_12007,N_12098);
nand U12326 (N_12326,N_12057,N_12153);
or U12327 (N_12327,N_12190,N_12029);
and U12328 (N_12328,N_12110,N_12064);
nor U12329 (N_12329,N_12136,N_12159);
nor U12330 (N_12330,N_12150,N_12088);
nand U12331 (N_12331,N_12070,N_12186);
or U12332 (N_12332,N_12126,N_12185);
nand U12333 (N_12333,N_12176,N_12108);
nor U12334 (N_12334,N_12090,N_12084);
xnor U12335 (N_12335,N_12184,N_12117);
and U12336 (N_12336,N_12068,N_12059);
xnor U12337 (N_12337,N_12137,N_12126);
and U12338 (N_12338,N_12040,N_12192);
or U12339 (N_12339,N_12164,N_12197);
xor U12340 (N_12340,N_12088,N_12119);
or U12341 (N_12341,N_12116,N_12004);
and U12342 (N_12342,N_12103,N_12069);
nand U12343 (N_12343,N_12061,N_12062);
or U12344 (N_12344,N_12042,N_12124);
xor U12345 (N_12345,N_12039,N_12121);
and U12346 (N_12346,N_12124,N_12035);
nor U12347 (N_12347,N_12038,N_12047);
xnor U12348 (N_12348,N_12031,N_12027);
and U12349 (N_12349,N_12058,N_12157);
nor U12350 (N_12350,N_12179,N_12128);
nand U12351 (N_12351,N_12057,N_12199);
xor U12352 (N_12352,N_12191,N_12040);
or U12353 (N_12353,N_12150,N_12148);
or U12354 (N_12354,N_12054,N_12189);
or U12355 (N_12355,N_12181,N_12176);
nand U12356 (N_12356,N_12108,N_12013);
nand U12357 (N_12357,N_12012,N_12102);
or U12358 (N_12358,N_12038,N_12001);
or U12359 (N_12359,N_12048,N_12111);
and U12360 (N_12360,N_12034,N_12117);
nand U12361 (N_12361,N_12058,N_12099);
nand U12362 (N_12362,N_12008,N_12119);
nor U12363 (N_12363,N_12045,N_12024);
and U12364 (N_12364,N_12112,N_12190);
nor U12365 (N_12365,N_12119,N_12000);
xnor U12366 (N_12366,N_12051,N_12008);
or U12367 (N_12367,N_12008,N_12065);
or U12368 (N_12368,N_12063,N_12095);
nor U12369 (N_12369,N_12084,N_12077);
xor U12370 (N_12370,N_12033,N_12017);
and U12371 (N_12371,N_12096,N_12009);
and U12372 (N_12372,N_12043,N_12032);
or U12373 (N_12373,N_12109,N_12175);
nand U12374 (N_12374,N_12095,N_12116);
or U12375 (N_12375,N_12181,N_12046);
xnor U12376 (N_12376,N_12122,N_12060);
xnor U12377 (N_12377,N_12143,N_12111);
or U12378 (N_12378,N_12113,N_12187);
nor U12379 (N_12379,N_12073,N_12111);
or U12380 (N_12380,N_12110,N_12097);
nor U12381 (N_12381,N_12181,N_12157);
nor U12382 (N_12382,N_12158,N_12195);
and U12383 (N_12383,N_12189,N_12090);
or U12384 (N_12384,N_12088,N_12117);
or U12385 (N_12385,N_12129,N_12008);
nand U12386 (N_12386,N_12036,N_12087);
nor U12387 (N_12387,N_12173,N_12041);
and U12388 (N_12388,N_12153,N_12005);
or U12389 (N_12389,N_12023,N_12049);
and U12390 (N_12390,N_12085,N_12026);
nor U12391 (N_12391,N_12139,N_12159);
and U12392 (N_12392,N_12036,N_12097);
nor U12393 (N_12393,N_12128,N_12030);
or U12394 (N_12394,N_12096,N_12112);
or U12395 (N_12395,N_12167,N_12068);
and U12396 (N_12396,N_12163,N_12124);
nand U12397 (N_12397,N_12087,N_12188);
nand U12398 (N_12398,N_12005,N_12133);
or U12399 (N_12399,N_12017,N_12007);
and U12400 (N_12400,N_12321,N_12386);
nor U12401 (N_12401,N_12371,N_12310);
nor U12402 (N_12402,N_12355,N_12356);
nor U12403 (N_12403,N_12364,N_12227);
or U12404 (N_12404,N_12305,N_12398);
nor U12405 (N_12405,N_12255,N_12312);
and U12406 (N_12406,N_12368,N_12228);
nor U12407 (N_12407,N_12346,N_12351);
nand U12408 (N_12408,N_12348,N_12277);
or U12409 (N_12409,N_12328,N_12311);
and U12410 (N_12410,N_12275,N_12218);
nor U12411 (N_12411,N_12204,N_12376);
nor U12412 (N_12412,N_12257,N_12265);
nor U12413 (N_12413,N_12387,N_12217);
xnor U12414 (N_12414,N_12307,N_12350);
nand U12415 (N_12415,N_12273,N_12211);
and U12416 (N_12416,N_12300,N_12222);
and U12417 (N_12417,N_12278,N_12287);
nand U12418 (N_12418,N_12269,N_12261);
nor U12419 (N_12419,N_12392,N_12323);
xor U12420 (N_12420,N_12393,N_12345);
and U12421 (N_12421,N_12389,N_12253);
xnor U12422 (N_12422,N_12259,N_12324);
and U12423 (N_12423,N_12317,N_12358);
or U12424 (N_12424,N_12375,N_12240);
and U12425 (N_12425,N_12374,N_12224);
nor U12426 (N_12426,N_12238,N_12266);
nor U12427 (N_12427,N_12303,N_12232);
or U12428 (N_12428,N_12363,N_12388);
nor U12429 (N_12429,N_12314,N_12272);
xnor U12430 (N_12430,N_12315,N_12316);
nand U12431 (N_12431,N_12234,N_12339);
xor U12432 (N_12432,N_12254,N_12396);
and U12433 (N_12433,N_12366,N_12225);
nand U12434 (N_12434,N_12208,N_12294);
and U12435 (N_12435,N_12214,N_12251);
or U12436 (N_12436,N_12216,N_12397);
and U12437 (N_12437,N_12209,N_12258);
and U12438 (N_12438,N_12248,N_12332);
nor U12439 (N_12439,N_12384,N_12354);
nor U12440 (N_12440,N_12377,N_12286);
nor U12441 (N_12441,N_12373,N_12243);
xnor U12442 (N_12442,N_12206,N_12349);
xnor U12443 (N_12443,N_12288,N_12365);
or U12444 (N_12444,N_12244,N_12270);
or U12445 (N_12445,N_12304,N_12229);
nand U12446 (N_12446,N_12337,N_12291);
nor U12447 (N_12447,N_12353,N_12241);
and U12448 (N_12448,N_12296,N_12325);
or U12449 (N_12449,N_12362,N_12359);
nand U12450 (N_12450,N_12200,N_12338);
nor U12451 (N_12451,N_12247,N_12347);
nand U12452 (N_12452,N_12308,N_12309);
nand U12453 (N_12453,N_12342,N_12221);
and U12454 (N_12454,N_12226,N_12249);
or U12455 (N_12455,N_12378,N_12382);
nor U12456 (N_12456,N_12395,N_12399);
nor U12457 (N_12457,N_12220,N_12301);
or U12458 (N_12458,N_12239,N_12381);
and U12459 (N_12459,N_12246,N_12213);
nor U12460 (N_12460,N_12335,N_12330);
or U12461 (N_12461,N_12279,N_12219);
nand U12462 (N_12462,N_12360,N_12370);
nand U12463 (N_12463,N_12380,N_12215);
xnor U12464 (N_12464,N_12242,N_12340);
or U12465 (N_12465,N_12341,N_12283);
nor U12466 (N_12466,N_12383,N_12271);
nor U12467 (N_12467,N_12267,N_12306);
nor U12468 (N_12468,N_12385,N_12329);
xnor U12469 (N_12469,N_12367,N_12318);
and U12470 (N_12470,N_12289,N_12297);
and U12471 (N_12471,N_12352,N_12235);
or U12472 (N_12472,N_12326,N_12256);
or U12473 (N_12473,N_12357,N_12262);
or U12474 (N_12474,N_12343,N_12298);
xor U12475 (N_12475,N_12202,N_12236);
nand U12476 (N_12476,N_12203,N_12231);
or U12477 (N_12477,N_12293,N_12333);
or U12478 (N_12478,N_12274,N_12268);
and U12479 (N_12479,N_12336,N_12295);
or U12480 (N_12480,N_12210,N_12212);
nor U12481 (N_12481,N_12281,N_12230);
nand U12482 (N_12482,N_12245,N_12299);
and U12483 (N_12483,N_12290,N_12250);
or U12484 (N_12484,N_12313,N_12331);
nor U12485 (N_12485,N_12372,N_12361);
nand U12486 (N_12486,N_12205,N_12260);
and U12487 (N_12487,N_12319,N_12263);
and U12488 (N_12488,N_12201,N_12276);
nor U12489 (N_12489,N_12369,N_12237);
or U12490 (N_12490,N_12390,N_12302);
nand U12491 (N_12491,N_12344,N_12284);
xnor U12492 (N_12492,N_12252,N_12285);
nand U12493 (N_12493,N_12394,N_12322);
nand U12494 (N_12494,N_12223,N_12207);
and U12495 (N_12495,N_12233,N_12334);
and U12496 (N_12496,N_12320,N_12264);
nor U12497 (N_12497,N_12327,N_12282);
and U12498 (N_12498,N_12391,N_12292);
nor U12499 (N_12499,N_12280,N_12379);
nor U12500 (N_12500,N_12227,N_12209);
xnor U12501 (N_12501,N_12322,N_12266);
nand U12502 (N_12502,N_12225,N_12274);
or U12503 (N_12503,N_12259,N_12205);
xnor U12504 (N_12504,N_12322,N_12312);
nand U12505 (N_12505,N_12225,N_12292);
nand U12506 (N_12506,N_12224,N_12371);
nand U12507 (N_12507,N_12300,N_12250);
nor U12508 (N_12508,N_12344,N_12282);
nor U12509 (N_12509,N_12344,N_12259);
nor U12510 (N_12510,N_12323,N_12263);
or U12511 (N_12511,N_12340,N_12219);
nor U12512 (N_12512,N_12202,N_12244);
or U12513 (N_12513,N_12318,N_12293);
nor U12514 (N_12514,N_12348,N_12215);
or U12515 (N_12515,N_12314,N_12366);
and U12516 (N_12516,N_12390,N_12266);
xnor U12517 (N_12517,N_12307,N_12344);
or U12518 (N_12518,N_12213,N_12375);
nand U12519 (N_12519,N_12244,N_12350);
nor U12520 (N_12520,N_12234,N_12250);
nand U12521 (N_12521,N_12384,N_12299);
and U12522 (N_12522,N_12234,N_12222);
or U12523 (N_12523,N_12358,N_12398);
or U12524 (N_12524,N_12212,N_12345);
nor U12525 (N_12525,N_12311,N_12253);
and U12526 (N_12526,N_12215,N_12317);
or U12527 (N_12527,N_12385,N_12341);
or U12528 (N_12528,N_12388,N_12205);
nor U12529 (N_12529,N_12398,N_12292);
nand U12530 (N_12530,N_12275,N_12240);
nand U12531 (N_12531,N_12251,N_12229);
or U12532 (N_12532,N_12371,N_12278);
nor U12533 (N_12533,N_12264,N_12314);
and U12534 (N_12534,N_12276,N_12380);
and U12535 (N_12535,N_12275,N_12254);
nand U12536 (N_12536,N_12359,N_12340);
xor U12537 (N_12537,N_12220,N_12377);
or U12538 (N_12538,N_12342,N_12344);
nor U12539 (N_12539,N_12285,N_12343);
nor U12540 (N_12540,N_12248,N_12230);
and U12541 (N_12541,N_12238,N_12261);
nor U12542 (N_12542,N_12221,N_12349);
xor U12543 (N_12543,N_12329,N_12357);
or U12544 (N_12544,N_12223,N_12398);
and U12545 (N_12545,N_12281,N_12378);
and U12546 (N_12546,N_12346,N_12225);
or U12547 (N_12547,N_12377,N_12258);
nor U12548 (N_12548,N_12350,N_12328);
nor U12549 (N_12549,N_12210,N_12229);
nand U12550 (N_12550,N_12319,N_12361);
nor U12551 (N_12551,N_12336,N_12296);
or U12552 (N_12552,N_12329,N_12256);
and U12553 (N_12553,N_12323,N_12385);
and U12554 (N_12554,N_12234,N_12392);
nand U12555 (N_12555,N_12335,N_12209);
or U12556 (N_12556,N_12221,N_12318);
or U12557 (N_12557,N_12245,N_12289);
nand U12558 (N_12558,N_12398,N_12364);
xnor U12559 (N_12559,N_12206,N_12236);
nor U12560 (N_12560,N_12241,N_12388);
nor U12561 (N_12561,N_12265,N_12310);
nand U12562 (N_12562,N_12380,N_12396);
nor U12563 (N_12563,N_12267,N_12316);
and U12564 (N_12564,N_12270,N_12212);
nor U12565 (N_12565,N_12300,N_12354);
or U12566 (N_12566,N_12337,N_12374);
or U12567 (N_12567,N_12397,N_12304);
and U12568 (N_12568,N_12296,N_12274);
nand U12569 (N_12569,N_12215,N_12332);
nor U12570 (N_12570,N_12385,N_12261);
and U12571 (N_12571,N_12357,N_12233);
and U12572 (N_12572,N_12214,N_12346);
xnor U12573 (N_12573,N_12272,N_12251);
nor U12574 (N_12574,N_12352,N_12367);
or U12575 (N_12575,N_12248,N_12316);
nor U12576 (N_12576,N_12369,N_12227);
nor U12577 (N_12577,N_12265,N_12364);
nand U12578 (N_12578,N_12381,N_12301);
xor U12579 (N_12579,N_12316,N_12331);
nand U12580 (N_12580,N_12230,N_12214);
and U12581 (N_12581,N_12308,N_12329);
xor U12582 (N_12582,N_12299,N_12278);
nor U12583 (N_12583,N_12209,N_12304);
and U12584 (N_12584,N_12336,N_12324);
nor U12585 (N_12585,N_12260,N_12362);
nand U12586 (N_12586,N_12366,N_12364);
and U12587 (N_12587,N_12303,N_12375);
nor U12588 (N_12588,N_12386,N_12260);
and U12589 (N_12589,N_12268,N_12232);
or U12590 (N_12590,N_12220,N_12249);
or U12591 (N_12591,N_12318,N_12253);
or U12592 (N_12592,N_12276,N_12264);
xnor U12593 (N_12593,N_12251,N_12369);
and U12594 (N_12594,N_12239,N_12271);
or U12595 (N_12595,N_12329,N_12306);
xnor U12596 (N_12596,N_12218,N_12242);
or U12597 (N_12597,N_12303,N_12356);
xor U12598 (N_12598,N_12228,N_12355);
or U12599 (N_12599,N_12212,N_12226);
xnor U12600 (N_12600,N_12531,N_12422);
and U12601 (N_12601,N_12408,N_12517);
nand U12602 (N_12602,N_12568,N_12485);
nand U12603 (N_12603,N_12409,N_12405);
and U12604 (N_12604,N_12579,N_12525);
and U12605 (N_12605,N_12501,N_12562);
nand U12606 (N_12606,N_12539,N_12441);
nor U12607 (N_12607,N_12466,N_12553);
or U12608 (N_12608,N_12592,N_12492);
nand U12609 (N_12609,N_12499,N_12563);
and U12610 (N_12610,N_12494,N_12464);
and U12611 (N_12611,N_12488,N_12576);
or U12612 (N_12612,N_12570,N_12419);
nor U12613 (N_12613,N_12478,N_12515);
xor U12614 (N_12614,N_12575,N_12402);
xor U12615 (N_12615,N_12439,N_12493);
and U12616 (N_12616,N_12430,N_12523);
or U12617 (N_12617,N_12588,N_12487);
and U12618 (N_12618,N_12471,N_12428);
xor U12619 (N_12619,N_12503,N_12470);
xnor U12620 (N_12620,N_12458,N_12489);
and U12621 (N_12621,N_12537,N_12583);
nor U12622 (N_12622,N_12532,N_12473);
nand U12623 (N_12623,N_12444,N_12585);
or U12624 (N_12624,N_12536,N_12593);
or U12625 (N_12625,N_12463,N_12502);
or U12626 (N_12626,N_12521,N_12508);
nor U12627 (N_12627,N_12555,N_12497);
and U12628 (N_12628,N_12433,N_12512);
and U12629 (N_12629,N_12567,N_12407);
and U12630 (N_12630,N_12545,N_12528);
and U12631 (N_12631,N_12560,N_12454);
and U12632 (N_12632,N_12417,N_12406);
nand U12633 (N_12633,N_12414,N_12462);
nand U12634 (N_12634,N_12477,N_12572);
xor U12635 (N_12635,N_12442,N_12460);
nand U12636 (N_12636,N_12578,N_12582);
xor U12637 (N_12637,N_12519,N_12586);
or U12638 (N_12638,N_12418,N_12561);
or U12639 (N_12639,N_12451,N_12518);
or U12640 (N_12640,N_12510,N_12479);
nor U12641 (N_12641,N_12429,N_12504);
nor U12642 (N_12642,N_12569,N_12557);
nand U12643 (N_12643,N_12558,N_12413);
nor U12644 (N_12644,N_12538,N_12544);
nor U12645 (N_12645,N_12410,N_12484);
or U12646 (N_12646,N_12411,N_12500);
nor U12647 (N_12647,N_12434,N_12581);
and U12648 (N_12648,N_12587,N_12415);
nor U12649 (N_12649,N_12595,N_12547);
nand U12650 (N_12650,N_12549,N_12527);
or U12651 (N_12651,N_12486,N_12573);
and U12652 (N_12652,N_12426,N_12421);
xnor U12653 (N_12653,N_12483,N_12534);
and U12654 (N_12654,N_12496,N_12565);
and U12655 (N_12655,N_12453,N_12450);
nor U12656 (N_12656,N_12548,N_12505);
or U12657 (N_12657,N_12580,N_12590);
nand U12658 (N_12658,N_12566,N_12491);
or U12659 (N_12659,N_12440,N_12481);
and U12660 (N_12660,N_12506,N_12447);
nand U12661 (N_12661,N_12541,N_12400);
nand U12662 (N_12662,N_12457,N_12514);
nand U12663 (N_12663,N_12507,N_12445);
nor U12664 (N_12664,N_12509,N_12596);
nor U12665 (N_12665,N_12472,N_12564);
nand U12666 (N_12666,N_12490,N_12533);
and U12667 (N_12667,N_12540,N_12516);
nor U12668 (N_12668,N_12546,N_12552);
or U12669 (N_12669,N_12467,N_12443);
and U12670 (N_12670,N_12543,N_12438);
or U12671 (N_12671,N_12449,N_12574);
and U12672 (N_12672,N_12577,N_12571);
nor U12673 (N_12673,N_12522,N_12431);
and U12674 (N_12674,N_12475,N_12403);
nand U12675 (N_12675,N_12459,N_12495);
or U12676 (N_12676,N_12551,N_12401);
nand U12677 (N_12677,N_12424,N_12556);
or U12678 (N_12678,N_12594,N_12529);
and U12679 (N_12679,N_12511,N_12456);
nand U12680 (N_12680,N_12436,N_12498);
and U12681 (N_12681,N_12530,N_12432);
xor U12682 (N_12682,N_12404,N_12423);
or U12683 (N_12683,N_12455,N_12437);
and U12684 (N_12684,N_12524,N_12448);
xor U12685 (N_12685,N_12598,N_12584);
nor U12686 (N_12686,N_12435,N_12589);
and U12687 (N_12687,N_12520,N_12474);
or U12688 (N_12688,N_12412,N_12446);
nor U12689 (N_12689,N_12476,N_12599);
or U12690 (N_12690,N_12559,N_12480);
nand U12691 (N_12691,N_12427,N_12461);
and U12692 (N_12692,N_12513,N_12535);
nor U12693 (N_12693,N_12416,N_12468);
nor U12694 (N_12694,N_12542,N_12482);
nor U12695 (N_12695,N_12465,N_12469);
and U12696 (N_12696,N_12526,N_12420);
xnor U12697 (N_12697,N_12554,N_12550);
or U12698 (N_12698,N_12425,N_12591);
nand U12699 (N_12699,N_12597,N_12452);
and U12700 (N_12700,N_12591,N_12408);
and U12701 (N_12701,N_12409,N_12436);
and U12702 (N_12702,N_12492,N_12511);
nor U12703 (N_12703,N_12560,N_12510);
or U12704 (N_12704,N_12533,N_12413);
nor U12705 (N_12705,N_12490,N_12581);
nor U12706 (N_12706,N_12412,N_12417);
nor U12707 (N_12707,N_12443,N_12440);
or U12708 (N_12708,N_12451,N_12519);
nand U12709 (N_12709,N_12401,N_12588);
nor U12710 (N_12710,N_12483,N_12400);
nor U12711 (N_12711,N_12527,N_12427);
and U12712 (N_12712,N_12470,N_12539);
nand U12713 (N_12713,N_12595,N_12476);
or U12714 (N_12714,N_12559,N_12434);
and U12715 (N_12715,N_12432,N_12570);
nor U12716 (N_12716,N_12434,N_12462);
nand U12717 (N_12717,N_12483,N_12560);
nor U12718 (N_12718,N_12573,N_12553);
or U12719 (N_12719,N_12584,N_12581);
and U12720 (N_12720,N_12512,N_12511);
nor U12721 (N_12721,N_12578,N_12491);
nor U12722 (N_12722,N_12588,N_12523);
nor U12723 (N_12723,N_12501,N_12475);
nor U12724 (N_12724,N_12518,N_12566);
nor U12725 (N_12725,N_12446,N_12489);
nor U12726 (N_12726,N_12570,N_12513);
or U12727 (N_12727,N_12465,N_12553);
and U12728 (N_12728,N_12413,N_12541);
xor U12729 (N_12729,N_12469,N_12409);
nor U12730 (N_12730,N_12465,N_12509);
nor U12731 (N_12731,N_12407,N_12503);
or U12732 (N_12732,N_12475,N_12525);
or U12733 (N_12733,N_12592,N_12446);
nand U12734 (N_12734,N_12537,N_12513);
or U12735 (N_12735,N_12508,N_12473);
nor U12736 (N_12736,N_12519,N_12498);
and U12737 (N_12737,N_12482,N_12505);
or U12738 (N_12738,N_12595,N_12511);
xnor U12739 (N_12739,N_12422,N_12493);
nand U12740 (N_12740,N_12493,N_12438);
nand U12741 (N_12741,N_12484,N_12429);
or U12742 (N_12742,N_12583,N_12467);
or U12743 (N_12743,N_12589,N_12424);
and U12744 (N_12744,N_12461,N_12408);
nand U12745 (N_12745,N_12515,N_12404);
or U12746 (N_12746,N_12484,N_12481);
nor U12747 (N_12747,N_12418,N_12589);
and U12748 (N_12748,N_12477,N_12595);
and U12749 (N_12749,N_12535,N_12502);
or U12750 (N_12750,N_12520,N_12597);
or U12751 (N_12751,N_12512,N_12480);
nand U12752 (N_12752,N_12457,N_12448);
and U12753 (N_12753,N_12591,N_12550);
nor U12754 (N_12754,N_12463,N_12431);
or U12755 (N_12755,N_12495,N_12491);
and U12756 (N_12756,N_12571,N_12441);
and U12757 (N_12757,N_12473,N_12548);
nand U12758 (N_12758,N_12501,N_12566);
or U12759 (N_12759,N_12469,N_12509);
or U12760 (N_12760,N_12520,N_12576);
nor U12761 (N_12761,N_12550,N_12476);
or U12762 (N_12762,N_12467,N_12561);
nand U12763 (N_12763,N_12579,N_12439);
nor U12764 (N_12764,N_12583,N_12598);
nand U12765 (N_12765,N_12557,N_12532);
or U12766 (N_12766,N_12506,N_12552);
nand U12767 (N_12767,N_12497,N_12462);
and U12768 (N_12768,N_12519,N_12541);
nor U12769 (N_12769,N_12405,N_12471);
or U12770 (N_12770,N_12549,N_12590);
nor U12771 (N_12771,N_12499,N_12418);
xor U12772 (N_12772,N_12533,N_12424);
nand U12773 (N_12773,N_12402,N_12586);
nand U12774 (N_12774,N_12545,N_12410);
and U12775 (N_12775,N_12422,N_12507);
nand U12776 (N_12776,N_12415,N_12448);
or U12777 (N_12777,N_12567,N_12525);
or U12778 (N_12778,N_12528,N_12513);
nor U12779 (N_12779,N_12579,N_12437);
nand U12780 (N_12780,N_12482,N_12560);
nor U12781 (N_12781,N_12558,N_12507);
nand U12782 (N_12782,N_12458,N_12587);
and U12783 (N_12783,N_12499,N_12491);
nand U12784 (N_12784,N_12432,N_12464);
or U12785 (N_12785,N_12520,N_12528);
nor U12786 (N_12786,N_12552,N_12499);
nand U12787 (N_12787,N_12516,N_12524);
nor U12788 (N_12788,N_12591,N_12411);
or U12789 (N_12789,N_12442,N_12583);
nand U12790 (N_12790,N_12481,N_12554);
nor U12791 (N_12791,N_12455,N_12554);
nor U12792 (N_12792,N_12586,N_12467);
nor U12793 (N_12793,N_12414,N_12575);
nand U12794 (N_12794,N_12522,N_12432);
or U12795 (N_12795,N_12417,N_12501);
nand U12796 (N_12796,N_12413,N_12425);
nand U12797 (N_12797,N_12434,N_12522);
nor U12798 (N_12798,N_12463,N_12434);
nand U12799 (N_12799,N_12543,N_12572);
or U12800 (N_12800,N_12677,N_12608);
and U12801 (N_12801,N_12708,N_12675);
or U12802 (N_12802,N_12663,N_12694);
or U12803 (N_12803,N_12793,N_12788);
nand U12804 (N_12804,N_12640,N_12783);
nand U12805 (N_12805,N_12693,N_12773);
or U12806 (N_12806,N_12723,N_12705);
or U12807 (N_12807,N_12776,N_12636);
and U12808 (N_12808,N_12797,N_12735);
and U12809 (N_12809,N_12777,N_12633);
and U12810 (N_12810,N_12734,N_12618);
nand U12811 (N_12811,N_12753,N_12645);
nor U12812 (N_12812,N_12648,N_12678);
or U12813 (N_12813,N_12738,N_12750);
xnor U12814 (N_12814,N_12626,N_12711);
nand U12815 (N_12815,N_12623,N_12765);
nor U12816 (N_12816,N_12722,N_12762);
or U12817 (N_12817,N_12644,N_12674);
nor U12818 (N_12818,N_12775,N_12712);
and U12819 (N_12819,N_12666,N_12649);
and U12820 (N_12820,N_12771,N_12763);
or U12821 (N_12821,N_12689,N_12690);
and U12822 (N_12822,N_12707,N_12770);
xor U12823 (N_12823,N_12761,N_12670);
or U12824 (N_12824,N_12661,N_12620);
nand U12825 (N_12825,N_12652,N_12791);
and U12826 (N_12826,N_12673,N_12628);
nor U12827 (N_12827,N_12601,N_12609);
or U12828 (N_12828,N_12726,N_12728);
and U12829 (N_12829,N_12660,N_12641);
nor U12830 (N_12830,N_12725,N_12758);
or U12831 (N_12831,N_12631,N_12716);
or U12832 (N_12832,N_12785,N_12606);
nand U12833 (N_12833,N_12779,N_12695);
or U12834 (N_12834,N_12732,N_12787);
xor U12835 (N_12835,N_12639,N_12752);
or U12836 (N_12836,N_12766,N_12704);
and U12837 (N_12837,N_12603,N_12701);
or U12838 (N_12838,N_12600,N_12730);
or U12839 (N_12839,N_12688,N_12676);
nand U12840 (N_12840,N_12746,N_12720);
and U12841 (N_12841,N_12622,N_12630);
or U12842 (N_12842,N_12602,N_12760);
or U12843 (N_12843,N_12627,N_12756);
nor U12844 (N_12844,N_12672,N_12792);
and U12845 (N_12845,N_12625,N_12768);
nand U12846 (N_12846,N_12796,N_12658);
nor U12847 (N_12847,N_12629,N_12615);
and U12848 (N_12848,N_12604,N_12710);
or U12849 (N_12849,N_12611,N_12780);
nand U12850 (N_12850,N_12664,N_12655);
nand U12851 (N_12851,N_12653,N_12782);
nand U12852 (N_12852,N_12715,N_12733);
nor U12853 (N_12853,N_12650,N_12698);
nor U12854 (N_12854,N_12621,N_12643);
nand U12855 (N_12855,N_12651,N_12743);
and U12856 (N_12856,N_12646,N_12772);
nor U12857 (N_12857,N_12786,N_12784);
and U12858 (N_12858,N_12709,N_12696);
nor U12859 (N_12859,N_12731,N_12617);
or U12860 (N_12860,N_12634,N_12749);
nand U12861 (N_12861,N_12635,N_12691);
nor U12862 (N_12862,N_12647,N_12665);
nand U12863 (N_12863,N_12745,N_12642);
and U12864 (N_12864,N_12607,N_12714);
nor U12865 (N_12865,N_12684,N_12702);
or U12866 (N_12866,N_12742,N_12703);
and U12867 (N_12867,N_12719,N_12736);
xnor U12868 (N_12868,N_12679,N_12795);
or U12869 (N_12869,N_12721,N_12748);
xor U12870 (N_12870,N_12619,N_12741);
or U12871 (N_12871,N_12683,N_12724);
nor U12872 (N_12872,N_12713,N_12790);
xnor U12873 (N_12873,N_12799,N_12789);
or U12874 (N_12874,N_12767,N_12632);
nand U12875 (N_12875,N_12605,N_12754);
nand U12876 (N_12876,N_12681,N_12668);
nor U12877 (N_12877,N_12798,N_12737);
nand U12878 (N_12878,N_12769,N_12637);
nor U12879 (N_12879,N_12751,N_12654);
or U12880 (N_12880,N_12781,N_12662);
and U12881 (N_12881,N_12682,N_12667);
or U12882 (N_12882,N_12692,N_12757);
nand U12883 (N_12883,N_12612,N_12613);
or U12884 (N_12884,N_12685,N_12669);
nor U12885 (N_12885,N_12614,N_12739);
and U12886 (N_12886,N_12755,N_12729);
and U12887 (N_12887,N_12624,N_12764);
and U12888 (N_12888,N_12656,N_12671);
and U12889 (N_12889,N_12778,N_12659);
or U12890 (N_12890,N_12700,N_12727);
and U12891 (N_12891,N_12747,N_12686);
nor U12892 (N_12892,N_12680,N_12616);
or U12893 (N_12893,N_12706,N_12657);
nand U12894 (N_12894,N_12610,N_12699);
or U12895 (N_12895,N_12638,N_12718);
nor U12896 (N_12896,N_12740,N_12794);
or U12897 (N_12897,N_12697,N_12744);
or U12898 (N_12898,N_12774,N_12687);
nand U12899 (N_12899,N_12717,N_12759);
nand U12900 (N_12900,N_12633,N_12608);
nor U12901 (N_12901,N_12752,N_12666);
and U12902 (N_12902,N_12742,N_12631);
or U12903 (N_12903,N_12625,N_12603);
and U12904 (N_12904,N_12796,N_12731);
nor U12905 (N_12905,N_12725,N_12741);
and U12906 (N_12906,N_12724,N_12633);
nand U12907 (N_12907,N_12705,N_12633);
nor U12908 (N_12908,N_12610,N_12790);
and U12909 (N_12909,N_12608,N_12734);
or U12910 (N_12910,N_12658,N_12623);
or U12911 (N_12911,N_12767,N_12782);
nand U12912 (N_12912,N_12760,N_12735);
nand U12913 (N_12913,N_12656,N_12659);
nor U12914 (N_12914,N_12678,N_12779);
or U12915 (N_12915,N_12748,N_12653);
nand U12916 (N_12916,N_12625,N_12711);
nand U12917 (N_12917,N_12709,N_12640);
nand U12918 (N_12918,N_12619,N_12778);
or U12919 (N_12919,N_12617,N_12616);
nor U12920 (N_12920,N_12654,N_12708);
or U12921 (N_12921,N_12627,N_12654);
or U12922 (N_12922,N_12638,N_12725);
nor U12923 (N_12923,N_12799,N_12668);
nor U12924 (N_12924,N_12635,N_12659);
or U12925 (N_12925,N_12745,N_12628);
nor U12926 (N_12926,N_12675,N_12700);
or U12927 (N_12927,N_12602,N_12609);
and U12928 (N_12928,N_12623,N_12655);
nor U12929 (N_12929,N_12644,N_12719);
and U12930 (N_12930,N_12710,N_12636);
nor U12931 (N_12931,N_12627,N_12783);
or U12932 (N_12932,N_12785,N_12775);
nand U12933 (N_12933,N_12642,N_12738);
nor U12934 (N_12934,N_12628,N_12693);
and U12935 (N_12935,N_12712,N_12765);
nand U12936 (N_12936,N_12600,N_12753);
and U12937 (N_12937,N_12699,N_12621);
and U12938 (N_12938,N_12696,N_12723);
nand U12939 (N_12939,N_12789,N_12655);
xor U12940 (N_12940,N_12710,N_12768);
nor U12941 (N_12941,N_12659,N_12700);
nor U12942 (N_12942,N_12710,N_12746);
nand U12943 (N_12943,N_12764,N_12674);
and U12944 (N_12944,N_12759,N_12715);
and U12945 (N_12945,N_12620,N_12781);
nand U12946 (N_12946,N_12653,N_12789);
nor U12947 (N_12947,N_12654,N_12775);
or U12948 (N_12948,N_12793,N_12711);
nand U12949 (N_12949,N_12651,N_12734);
and U12950 (N_12950,N_12747,N_12799);
or U12951 (N_12951,N_12738,N_12643);
and U12952 (N_12952,N_12651,N_12729);
or U12953 (N_12953,N_12609,N_12607);
nor U12954 (N_12954,N_12634,N_12630);
nor U12955 (N_12955,N_12758,N_12798);
nor U12956 (N_12956,N_12684,N_12647);
nand U12957 (N_12957,N_12753,N_12752);
nor U12958 (N_12958,N_12719,N_12743);
and U12959 (N_12959,N_12671,N_12634);
nor U12960 (N_12960,N_12698,N_12695);
nand U12961 (N_12961,N_12753,N_12713);
or U12962 (N_12962,N_12729,N_12764);
nand U12963 (N_12963,N_12641,N_12637);
and U12964 (N_12964,N_12602,N_12673);
or U12965 (N_12965,N_12741,N_12637);
nand U12966 (N_12966,N_12705,N_12645);
nand U12967 (N_12967,N_12711,N_12694);
or U12968 (N_12968,N_12650,N_12726);
and U12969 (N_12969,N_12699,N_12744);
and U12970 (N_12970,N_12797,N_12678);
and U12971 (N_12971,N_12639,N_12720);
nand U12972 (N_12972,N_12639,N_12646);
and U12973 (N_12973,N_12752,N_12668);
or U12974 (N_12974,N_12749,N_12666);
xor U12975 (N_12975,N_12730,N_12683);
and U12976 (N_12976,N_12707,N_12687);
and U12977 (N_12977,N_12654,N_12784);
and U12978 (N_12978,N_12692,N_12677);
and U12979 (N_12979,N_12739,N_12653);
xnor U12980 (N_12980,N_12623,N_12760);
nor U12981 (N_12981,N_12613,N_12636);
nor U12982 (N_12982,N_12711,N_12799);
nor U12983 (N_12983,N_12650,N_12652);
and U12984 (N_12984,N_12664,N_12722);
xnor U12985 (N_12985,N_12763,N_12719);
nand U12986 (N_12986,N_12751,N_12610);
and U12987 (N_12987,N_12751,N_12653);
nor U12988 (N_12988,N_12686,N_12749);
nand U12989 (N_12989,N_12645,N_12626);
nand U12990 (N_12990,N_12750,N_12623);
nand U12991 (N_12991,N_12717,N_12736);
and U12992 (N_12992,N_12663,N_12604);
or U12993 (N_12993,N_12672,N_12754);
and U12994 (N_12994,N_12634,N_12665);
or U12995 (N_12995,N_12781,N_12600);
nand U12996 (N_12996,N_12734,N_12792);
or U12997 (N_12997,N_12727,N_12627);
nor U12998 (N_12998,N_12704,N_12681);
and U12999 (N_12999,N_12692,N_12790);
or U13000 (N_13000,N_12883,N_12923);
nand U13001 (N_13001,N_12992,N_12853);
or U13002 (N_13002,N_12944,N_12899);
nor U13003 (N_13003,N_12814,N_12806);
or U13004 (N_13004,N_12967,N_12975);
nor U13005 (N_13005,N_12848,N_12864);
xnor U13006 (N_13006,N_12912,N_12926);
nand U13007 (N_13007,N_12935,N_12805);
nor U13008 (N_13008,N_12934,N_12979);
xnor U13009 (N_13009,N_12894,N_12955);
nand U13010 (N_13010,N_12933,N_12841);
nand U13011 (N_13011,N_12986,N_12873);
nand U13012 (N_13012,N_12844,N_12990);
nor U13013 (N_13013,N_12905,N_12801);
nand U13014 (N_13014,N_12968,N_12974);
and U13015 (N_13015,N_12834,N_12982);
or U13016 (N_13016,N_12915,N_12959);
or U13017 (N_13017,N_12983,N_12849);
nor U13018 (N_13018,N_12846,N_12838);
nor U13019 (N_13019,N_12895,N_12859);
and U13020 (N_13020,N_12800,N_12994);
or U13021 (N_13021,N_12962,N_12917);
nor U13022 (N_13022,N_12941,N_12939);
nand U13023 (N_13023,N_12845,N_12901);
or U13024 (N_13024,N_12900,N_12916);
nor U13025 (N_13025,N_12958,N_12854);
nor U13026 (N_13026,N_12987,N_12950);
xnor U13027 (N_13027,N_12808,N_12811);
nand U13028 (N_13028,N_12822,N_12981);
nor U13029 (N_13029,N_12932,N_12971);
nor U13030 (N_13030,N_12988,N_12888);
and U13031 (N_13031,N_12946,N_12833);
or U13032 (N_13032,N_12837,N_12884);
nor U13033 (N_13033,N_12831,N_12869);
nand U13034 (N_13034,N_12972,N_12898);
nor U13035 (N_13035,N_12855,N_12928);
and U13036 (N_13036,N_12824,N_12889);
nor U13037 (N_13037,N_12902,N_12871);
nor U13038 (N_13038,N_12861,N_12887);
or U13039 (N_13039,N_12879,N_12892);
xnor U13040 (N_13040,N_12862,N_12910);
nor U13041 (N_13041,N_12999,N_12815);
nor U13042 (N_13042,N_12809,N_12947);
or U13043 (N_13043,N_12847,N_12828);
or U13044 (N_13044,N_12995,N_12819);
or U13045 (N_13045,N_12872,N_12961);
or U13046 (N_13046,N_12909,N_12842);
nor U13047 (N_13047,N_12891,N_12970);
and U13048 (N_13048,N_12817,N_12852);
nand U13049 (N_13049,N_12818,N_12810);
nor U13050 (N_13050,N_12963,N_12940);
and U13051 (N_13051,N_12851,N_12973);
and U13052 (N_13052,N_12965,N_12870);
nand U13053 (N_13053,N_12922,N_12936);
nand U13054 (N_13054,N_12943,N_12913);
and U13055 (N_13055,N_12840,N_12813);
nor U13056 (N_13056,N_12969,N_12906);
and U13057 (N_13057,N_12893,N_12966);
or U13058 (N_13058,N_12911,N_12868);
and U13059 (N_13059,N_12985,N_12897);
xor U13060 (N_13060,N_12850,N_12803);
nand U13061 (N_13061,N_12825,N_12839);
nand U13062 (N_13062,N_12948,N_12949);
nand U13063 (N_13063,N_12832,N_12816);
and U13064 (N_13064,N_12802,N_12980);
nand U13065 (N_13065,N_12924,N_12881);
nand U13066 (N_13066,N_12952,N_12860);
nand U13067 (N_13067,N_12856,N_12938);
and U13068 (N_13068,N_12976,N_12823);
nand U13069 (N_13069,N_12836,N_12977);
xnor U13070 (N_13070,N_12921,N_12993);
nand U13071 (N_13071,N_12920,N_12914);
nand U13072 (N_13072,N_12827,N_12877);
xor U13073 (N_13073,N_12821,N_12953);
or U13074 (N_13074,N_12942,N_12907);
or U13075 (N_13075,N_12876,N_12991);
nor U13076 (N_13076,N_12951,N_12896);
and U13077 (N_13077,N_12996,N_12954);
or U13078 (N_13078,N_12880,N_12829);
and U13079 (N_13079,N_12804,N_12807);
nand U13080 (N_13080,N_12904,N_12886);
nand U13081 (N_13081,N_12960,N_12927);
or U13082 (N_13082,N_12903,N_12866);
or U13083 (N_13083,N_12882,N_12835);
nor U13084 (N_13084,N_12919,N_12875);
and U13085 (N_13085,N_12957,N_12858);
nand U13086 (N_13086,N_12978,N_12931);
and U13087 (N_13087,N_12929,N_12890);
or U13088 (N_13088,N_12830,N_12874);
and U13089 (N_13089,N_12878,N_12984);
and U13090 (N_13090,N_12857,N_12908);
nand U13091 (N_13091,N_12918,N_12865);
or U13092 (N_13092,N_12843,N_12863);
and U13093 (N_13093,N_12997,N_12826);
nor U13094 (N_13094,N_12925,N_12867);
nand U13095 (N_13095,N_12945,N_12956);
nor U13096 (N_13096,N_12964,N_12998);
and U13097 (N_13097,N_12812,N_12885);
nand U13098 (N_13098,N_12989,N_12930);
and U13099 (N_13099,N_12937,N_12820);
nand U13100 (N_13100,N_12945,N_12868);
or U13101 (N_13101,N_12966,N_12830);
nor U13102 (N_13102,N_12880,N_12864);
nor U13103 (N_13103,N_12904,N_12848);
and U13104 (N_13104,N_12832,N_12882);
nand U13105 (N_13105,N_12809,N_12885);
nand U13106 (N_13106,N_12956,N_12891);
or U13107 (N_13107,N_12932,N_12924);
nor U13108 (N_13108,N_12844,N_12861);
nor U13109 (N_13109,N_12886,N_12901);
nor U13110 (N_13110,N_12831,N_12832);
or U13111 (N_13111,N_12846,N_12952);
nor U13112 (N_13112,N_12838,N_12929);
or U13113 (N_13113,N_12950,N_12991);
nand U13114 (N_13114,N_12880,N_12940);
nand U13115 (N_13115,N_12810,N_12907);
and U13116 (N_13116,N_12823,N_12902);
nor U13117 (N_13117,N_12813,N_12968);
nor U13118 (N_13118,N_12931,N_12973);
nand U13119 (N_13119,N_12974,N_12883);
and U13120 (N_13120,N_12899,N_12955);
and U13121 (N_13121,N_12822,N_12884);
and U13122 (N_13122,N_12964,N_12822);
and U13123 (N_13123,N_12826,N_12999);
nand U13124 (N_13124,N_12885,N_12944);
and U13125 (N_13125,N_12805,N_12816);
or U13126 (N_13126,N_12859,N_12981);
or U13127 (N_13127,N_12988,N_12885);
nor U13128 (N_13128,N_12868,N_12867);
and U13129 (N_13129,N_12973,N_12845);
nand U13130 (N_13130,N_12928,N_12831);
or U13131 (N_13131,N_12908,N_12957);
nor U13132 (N_13132,N_12975,N_12818);
or U13133 (N_13133,N_12916,N_12869);
nor U13134 (N_13134,N_12921,N_12900);
and U13135 (N_13135,N_12820,N_12901);
or U13136 (N_13136,N_12983,N_12985);
and U13137 (N_13137,N_12863,N_12998);
nor U13138 (N_13138,N_12986,N_12822);
and U13139 (N_13139,N_12801,N_12985);
and U13140 (N_13140,N_12960,N_12911);
nor U13141 (N_13141,N_12953,N_12853);
xor U13142 (N_13142,N_12908,N_12890);
and U13143 (N_13143,N_12870,N_12860);
xor U13144 (N_13144,N_12949,N_12990);
or U13145 (N_13145,N_12819,N_12843);
and U13146 (N_13146,N_12814,N_12828);
nand U13147 (N_13147,N_12856,N_12862);
nand U13148 (N_13148,N_12915,N_12836);
or U13149 (N_13149,N_12995,N_12829);
nor U13150 (N_13150,N_12867,N_12932);
nand U13151 (N_13151,N_12941,N_12827);
nand U13152 (N_13152,N_12814,N_12835);
or U13153 (N_13153,N_12807,N_12922);
nor U13154 (N_13154,N_12936,N_12941);
xnor U13155 (N_13155,N_12925,N_12946);
nand U13156 (N_13156,N_12916,N_12811);
nor U13157 (N_13157,N_12919,N_12847);
xnor U13158 (N_13158,N_12818,N_12977);
and U13159 (N_13159,N_12803,N_12973);
or U13160 (N_13160,N_12824,N_12811);
or U13161 (N_13161,N_12839,N_12991);
nor U13162 (N_13162,N_12977,N_12940);
nor U13163 (N_13163,N_12953,N_12805);
or U13164 (N_13164,N_12801,N_12936);
nand U13165 (N_13165,N_12873,N_12840);
or U13166 (N_13166,N_12846,N_12949);
and U13167 (N_13167,N_12989,N_12904);
and U13168 (N_13168,N_12899,N_12965);
nor U13169 (N_13169,N_12965,N_12969);
and U13170 (N_13170,N_12900,N_12973);
nand U13171 (N_13171,N_12931,N_12917);
nand U13172 (N_13172,N_12809,N_12987);
or U13173 (N_13173,N_12831,N_12824);
and U13174 (N_13174,N_12946,N_12835);
nand U13175 (N_13175,N_12916,N_12887);
and U13176 (N_13176,N_12910,N_12981);
xnor U13177 (N_13177,N_12986,N_12945);
nor U13178 (N_13178,N_12972,N_12927);
nand U13179 (N_13179,N_12807,N_12860);
or U13180 (N_13180,N_12899,N_12850);
nand U13181 (N_13181,N_12935,N_12897);
nand U13182 (N_13182,N_12919,N_12944);
nor U13183 (N_13183,N_12895,N_12829);
xor U13184 (N_13184,N_12836,N_12822);
nand U13185 (N_13185,N_12805,N_12982);
nand U13186 (N_13186,N_12981,N_12811);
nand U13187 (N_13187,N_12824,N_12961);
or U13188 (N_13188,N_12957,N_12892);
xor U13189 (N_13189,N_12833,N_12981);
or U13190 (N_13190,N_12801,N_12944);
nand U13191 (N_13191,N_12993,N_12814);
or U13192 (N_13192,N_12934,N_12835);
and U13193 (N_13193,N_12956,N_12899);
and U13194 (N_13194,N_12836,N_12926);
nor U13195 (N_13195,N_12919,N_12996);
nor U13196 (N_13196,N_12993,N_12892);
nand U13197 (N_13197,N_12882,N_12841);
or U13198 (N_13198,N_12992,N_12860);
nor U13199 (N_13199,N_12914,N_12892);
nor U13200 (N_13200,N_13128,N_13014);
and U13201 (N_13201,N_13162,N_13035);
nand U13202 (N_13202,N_13199,N_13030);
or U13203 (N_13203,N_13023,N_13032);
or U13204 (N_13204,N_13187,N_13140);
nand U13205 (N_13205,N_13018,N_13011);
nand U13206 (N_13206,N_13053,N_13034);
or U13207 (N_13207,N_13136,N_13055);
or U13208 (N_13208,N_13193,N_13078);
xnor U13209 (N_13209,N_13067,N_13194);
nor U13210 (N_13210,N_13144,N_13121);
and U13211 (N_13211,N_13197,N_13098);
nor U13212 (N_13212,N_13024,N_13045);
or U13213 (N_13213,N_13108,N_13182);
or U13214 (N_13214,N_13026,N_13189);
nand U13215 (N_13215,N_13104,N_13184);
nor U13216 (N_13216,N_13083,N_13036);
and U13217 (N_13217,N_13129,N_13050);
nand U13218 (N_13218,N_13179,N_13052);
and U13219 (N_13219,N_13141,N_13151);
or U13220 (N_13220,N_13090,N_13132);
nand U13221 (N_13221,N_13016,N_13178);
nor U13222 (N_13222,N_13019,N_13073);
nand U13223 (N_13223,N_13080,N_13123);
nor U13224 (N_13224,N_13106,N_13093);
or U13225 (N_13225,N_13038,N_13049);
or U13226 (N_13226,N_13153,N_13095);
or U13227 (N_13227,N_13092,N_13099);
and U13228 (N_13228,N_13075,N_13008);
and U13229 (N_13229,N_13111,N_13029);
nor U13230 (N_13230,N_13116,N_13041);
xor U13231 (N_13231,N_13154,N_13198);
and U13232 (N_13232,N_13148,N_13031);
or U13233 (N_13233,N_13020,N_13022);
xor U13234 (N_13234,N_13040,N_13059);
nand U13235 (N_13235,N_13159,N_13192);
xnor U13236 (N_13236,N_13068,N_13046);
xnor U13237 (N_13237,N_13190,N_13088);
nand U13238 (N_13238,N_13165,N_13065);
or U13239 (N_13239,N_13183,N_13064);
and U13240 (N_13240,N_13180,N_13004);
nand U13241 (N_13241,N_13058,N_13101);
or U13242 (N_13242,N_13155,N_13146);
nand U13243 (N_13243,N_13118,N_13051);
xor U13244 (N_13244,N_13085,N_13074);
nor U13245 (N_13245,N_13094,N_13196);
or U13246 (N_13246,N_13027,N_13077);
nand U13247 (N_13247,N_13097,N_13164);
nand U13248 (N_13248,N_13168,N_13010);
nor U13249 (N_13249,N_13115,N_13100);
xnor U13250 (N_13250,N_13042,N_13131);
nand U13251 (N_13251,N_13125,N_13086);
xor U13252 (N_13252,N_13066,N_13127);
nor U13253 (N_13253,N_13166,N_13005);
nor U13254 (N_13254,N_13114,N_13013);
or U13255 (N_13255,N_13175,N_13057);
and U13256 (N_13256,N_13001,N_13170);
xnor U13257 (N_13257,N_13134,N_13149);
or U13258 (N_13258,N_13137,N_13033);
nand U13259 (N_13259,N_13007,N_13188);
nor U13260 (N_13260,N_13173,N_13181);
or U13261 (N_13261,N_13039,N_13124);
nand U13262 (N_13262,N_13069,N_13156);
nor U13263 (N_13263,N_13070,N_13126);
and U13264 (N_13264,N_13002,N_13109);
nand U13265 (N_13265,N_13091,N_13143);
and U13266 (N_13266,N_13087,N_13147);
xor U13267 (N_13267,N_13006,N_13195);
or U13268 (N_13268,N_13186,N_13072);
nand U13269 (N_13269,N_13163,N_13105);
or U13270 (N_13270,N_13120,N_13139);
nand U13271 (N_13271,N_13044,N_13102);
or U13272 (N_13272,N_13062,N_13060);
nor U13273 (N_13273,N_13160,N_13110);
nor U13274 (N_13274,N_13169,N_13113);
xnor U13275 (N_13275,N_13135,N_13015);
or U13276 (N_13276,N_13082,N_13047);
nor U13277 (N_13277,N_13043,N_13054);
or U13278 (N_13278,N_13112,N_13103);
nor U13279 (N_13279,N_13071,N_13056);
and U13280 (N_13280,N_13176,N_13081);
and U13281 (N_13281,N_13076,N_13119);
nor U13282 (N_13282,N_13117,N_13009);
nand U13283 (N_13283,N_13133,N_13171);
and U13284 (N_13284,N_13003,N_13167);
nand U13285 (N_13285,N_13048,N_13089);
xnor U13286 (N_13286,N_13161,N_13130);
and U13287 (N_13287,N_13122,N_13174);
or U13288 (N_13288,N_13021,N_13138);
and U13289 (N_13289,N_13028,N_13079);
or U13290 (N_13290,N_13000,N_13152);
or U13291 (N_13291,N_13145,N_13061);
xnor U13292 (N_13292,N_13150,N_13177);
nor U13293 (N_13293,N_13037,N_13142);
and U13294 (N_13294,N_13191,N_13096);
nor U13295 (N_13295,N_13063,N_13157);
or U13296 (N_13296,N_13025,N_13017);
nand U13297 (N_13297,N_13172,N_13084);
xor U13298 (N_13298,N_13107,N_13012);
nor U13299 (N_13299,N_13185,N_13158);
and U13300 (N_13300,N_13042,N_13045);
or U13301 (N_13301,N_13146,N_13123);
xnor U13302 (N_13302,N_13076,N_13140);
nor U13303 (N_13303,N_13064,N_13096);
nand U13304 (N_13304,N_13182,N_13142);
nand U13305 (N_13305,N_13131,N_13128);
nor U13306 (N_13306,N_13116,N_13016);
or U13307 (N_13307,N_13141,N_13199);
nor U13308 (N_13308,N_13172,N_13087);
nor U13309 (N_13309,N_13174,N_13083);
nand U13310 (N_13310,N_13129,N_13116);
or U13311 (N_13311,N_13185,N_13115);
and U13312 (N_13312,N_13117,N_13042);
nor U13313 (N_13313,N_13128,N_13052);
nor U13314 (N_13314,N_13172,N_13112);
and U13315 (N_13315,N_13165,N_13188);
and U13316 (N_13316,N_13150,N_13029);
xor U13317 (N_13317,N_13193,N_13093);
or U13318 (N_13318,N_13141,N_13015);
and U13319 (N_13319,N_13073,N_13148);
or U13320 (N_13320,N_13119,N_13172);
and U13321 (N_13321,N_13078,N_13157);
or U13322 (N_13322,N_13058,N_13008);
nand U13323 (N_13323,N_13063,N_13182);
and U13324 (N_13324,N_13183,N_13099);
nor U13325 (N_13325,N_13108,N_13157);
xor U13326 (N_13326,N_13082,N_13120);
nor U13327 (N_13327,N_13138,N_13120);
nor U13328 (N_13328,N_13024,N_13093);
nand U13329 (N_13329,N_13174,N_13075);
xor U13330 (N_13330,N_13112,N_13007);
nand U13331 (N_13331,N_13124,N_13097);
or U13332 (N_13332,N_13155,N_13079);
and U13333 (N_13333,N_13125,N_13162);
or U13334 (N_13334,N_13125,N_13184);
and U13335 (N_13335,N_13109,N_13101);
nand U13336 (N_13336,N_13060,N_13155);
nor U13337 (N_13337,N_13018,N_13169);
nor U13338 (N_13338,N_13011,N_13044);
nor U13339 (N_13339,N_13020,N_13110);
and U13340 (N_13340,N_13031,N_13098);
nor U13341 (N_13341,N_13107,N_13169);
nand U13342 (N_13342,N_13161,N_13141);
or U13343 (N_13343,N_13188,N_13143);
or U13344 (N_13344,N_13119,N_13008);
nand U13345 (N_13345,N_13021,N_13168);
and U13346 (N_13346,N_13003,N_13063);
xor U13347 (N_13347,N_13007,N_13018);
nor U13348 (N_13348,N_13066,N_13196);
and U13349 (N_13349,N_13088,N_13124);
and U13350 (N_13350,N_13184,N_13064);
or U13351 (N_13351,N_13072,N_13045);
and U13352 (N_13352,N_13025,N_13011);
nand U13353 (N_13353,N_13025,N_13056);
nand U13354 (N_13354,N_13169,N_13164);
or U13355 (N_13355,N_13123,N_13010);
nand U13356 (N_13356,N_13044,N_13115);
nand U13357 (N_13357,N_13125,N_13192);
xor U13358 (N_13358,N_13178,N_13127);
nand U13359 (N_13359,N_13035,N_13128);
and U13360 (N_13360,N_13042,N_13094);
nand U13361 (N_13361,N_13060,N_13110);
and U13362 (N_13362,N_13077,N_13086);
nand U13363 (N_13363,N_13191,N_13144);
or U13364 (N_13364,N_13129,N_13143);
nand U13365 (N_13365,N_13165,N_13105);
xnor U13366 (N_13366,N_13197,N_13068);
and U13367 (N_13367,N_13017,N_13117);
and U13368 (N_13368,N_13053,N_13181);
nand U13369 (N_13369,N_13159,N_13161);
or U13370 (N_13370,N_13042,N_13063);
nand U13371 (N_13371,N_13027,N_13097);
nand U13372 (N_13372,N_13180,N_13127);
nor U13373 (N_13373,N_13157,N_13113);
or U13374 (N_13374,N_13055,N_13077);
nor U13375 (N_13375,N_13176,N_13021);
nor U13376 (N_13376,N_13085,N_13141);
nand U13377 (N_13377,N_13025,N_13023);
and U13378 (N_13378,N_13197,N_13039);
and U13379 (N_13379,N_13073,N_13071);
nor U13380 (N_13380,N_13077,N_13186);
nor U13381 (N_13381,N_13185,N_13109);
nand U13382 (N_13382,N_13187,N_13090);
or U13383 (N_13383,N_13139,N_13160);
or U13384 (N_13384,N_13151,N_13003);
or U13385 (N_13385,N_13093,N_13056);
nand U13386 (N_13386,N_13198,N_13153);
xnor U13387 (N_13387,N_13049,N_13177);
nor U13388 (N_13388,N_13020,N_13106);
nand U13389 (N_13389,N_13170,N_13114);
or U13390 (N_13390,N_13118,N_13114);
and U13391 (N_13391,N_13025,N_13102);
nand U13392 (N_13392,N_13159,N_13125);
nor U13393 (N_13393,N_13030,N_13014);
or U13394 (N_13394,N_13194,N_13121);
or U13395 (N_13395,N_13030,N_13182);
or U13396 (N_13396,N_13147,N_13105);
and U13397 (N_13397,N_13103,N_13024);
nand U13398 (N_13398,N_13099,N_13166);
nor U13399 (N_13399,N_13199,N_13064);
xnor U13400 (N_13400,N_13371,N_13214);
and U13401 (N_13401,N_13373,N_13314);
xor U13402 (N_13402,N_13346,N_13228);
and U13403 (N_13403,N_13353,N_13354);
or U13404 (N_13404,N_13399,N_13238);
or U13405 (N_13405,N_13394,N_13279);
or U13406 (N_13406,N_13215,N_13285);
and U13407 (N_13407,N_13218,N_13391);
and U13408 (N_13408,N_13395,N_13256);
nor U13409 (N_13409,N_13249,N_13323);
and U13410 (N_13410,N_13207,N_13339);
or U13411 (N_13411,N_13363,N_13345);
xnor U13412 (N_13412,N_13334,N_13216);
nor U13413 (N_13413,N_13310,N_13302);
nand U13414 (N_13414,N_13356,N_13389);
nand U13415 (N_13415,N_13393,N_13270);
and U13416 (N_13416,N_13269,N_13222);
nor U13417 (N_13417,N_13255,N_13397);
or U13418 (N_13418,N_13376,N_13331);
or U13419 (N_13419,N_13358,N_13266);
nand U13420 (N_13420,N_13299,N_13326);
or U13421 (N_13421,N_13227,N_13337);
or U13422 (N_13422,N_13303,N_13246);
nor U13423 (N_13423,N_13308,N_13368);
nor U13424 (N_13424,N_13300,N_13250);
and U13425 (N_13425,N_13289,N_13386);
nor U13426 (N_13426,N_13262,N_13297);
nor U13427 (N_13427,N_13240,N_13280);
nor U13428 (N_13428,N_13294,N_13208);
nor U13429 (N_13429,N_13224,N_13298);
nor U13430 (N_13430,N_13281,N_13319);
nand U13431 (N_13431,N_13315,N_13237);
xnor U13432 (N_13432,N_13210,N_13313);
nand U13433 (N_13433,N_13234,N_13387);
xor U13434 (N_13434,N_13351,N_13388);
or U13435 (N_13435,N_13295,N_13322);
and U13436 (N_13436,N_13350,N_13321);
and U13437 (N_13437,N_13252,N_13336);
and U13438 (N_13438,N_13332,N_13384);
nor U13439 (N_13439,N_13248,N_13204);
xor U13440 (N_13440,N_13292,N_13272);
or U13441 (N_13441,N_13277,N_13268);
and U13442 (N_13442,N_13284,N_13372);
and U13443 (N_13443,N_13309,N_13293);
nand U13444 (N_13444,N_13328,N_13283);
or U13445 (N_13445,N_13347,N_13366);
nor U13446 (N_13446,N_13317,N_13352);
nand U13447 (N_13447,N_13273,N_13264);
nor U13448 (N_13448,N_13385,N_13349);
and U13449 (N_13449,N_13392,N_13367);
or U13450 (N_13450,N_13217,N_13236);
xor U13451 (N_13451,N_13235,N_13370);
and U13452 (N_13452,N_13390,N_13343);
nand U13453 (N_13453,N_13338,N_13211);
or U13454 (N_13454,N_13398,N_13374);
nor U13455 (N_13455,N_13301,N_13383);
and U13456 (N_13456,N_13274,N_13325);
and U13457 (N_13457,N_13306,N_13231);
nand U13458 (N_13458,N_13239,N_13260);
nand U13459 (N_13459,N_13205,N_13307);
nor U13460 (N_13460,N_13271,N_13267);
nand U13461 (N_13461,N_13232,N_13379);
nand U13462 (N_13462,N_13258,N_13335);
and U13463 (N_13463,N_13226,N_13396);
nor U13464 (N_13464,N_13242,N_13265);
or U13465 (N_13465,N_13381,N_13359);
nand U13466 (N_13466,N_13378,N_13330);
and U13467 (N_13467,N_13369,N_13247);
xor U13468 (N_13468,N_13342,N_13275);
nor U13469 (N_13469,N_13253,N_13221);
and U13470 (N_13470,N_13223,N_13219);
or U13471 (N_13471,N_13305,N_13202);
nor U13472 (N_13472,N_13327,N_13229);
nor U13473 (N_13473,N_13324,N_13209);
or U13474 (N_13474,N_13361,N_13341);
xnor U13475 (N_13475,N_13312,N_13344);
xnor U13476 (N_13476,N_13329,N_13318);
nand U13477 (N_13477,N_13200,N_13320);
nand U13478 (N_13478,N_13257,N_13278);
xnor U13479 (N_13479,N_13348,N_13316);
nand U13480 (N_13480,N_13263,N_13304);
xnor U13481 (N_13481,N_13254,N_13212);
nor U13482 (N_13482,N_13261,N_13244);
and U13483 (N_13483,N_13225,N_13251);
nand U13484 (N_13484,N_13245,N_13206);
nand U13485 (N_13485,N_13243,N_13241);
and U13486 (N_13486,N_13362,N_13333);
and U13487 (N_13487,N_13364,N_13375);
and U13488 (N_13488,N_13282,N_13290);
nand U13489 (N_13489,N_13382,N_13201);
and U13490 (N_13490,N_13220,N_13296);
and U13491 (N_13491,N_13213,N_13203);
nor U13492 (N_13492,N_13357,N_13365);
nor U13493 (N_13493,N_13311,N_13286);
xnor U13494 (N_13494,N_13291,N_13287);
or U13495 (N_13495,N_13360,N_13288);
nor U13496 (N_13496,N_13259,N_13377);
or U13497 (N_13497,N_13230,N_13380);
and U13498 (N_13498,N_13233,N_13355);
or U13499 (N_13499,N_13276,N_13340);
nor U13500 (N_13500,N_13226,N_13229);
or U13501 (N_13501,N_13345,N_13366);
nand U13502 (N_13502,N_13317,N_13294);
nand U13503 (N_13503,N_13297,N_13258);
nand U13504 (N_13504,N_13296,N_13218);
and U13505 (N_13505,N_13203,N_13327);
and U13506 (N_13506,N_13230,N_13261);
nor U13507 (N_13507,N_13264,N_13263);
nor U13508 (N_13508,N_13326,N_13298);
xnor U13509 (N_13509,N_13356,N_13263);
or U13510 (N_13510,N_13229,N_13388);
or U13511 (N_13511,N_13300,N_13215);
or U13512 (N_13512,N_13384,N_13255);
or U13513 (N_13513,N_13234,N_13394);
nand U13514 (N_13514,N_13330,N_13237);
or U13515 (N_13515,N_13252,N_13221);
nand U13516 (N_13516,N_13304,N_13372);
and U13517 (N_13517,N_13347,N_13229);
nor U13518 (N_13518,N_13307,N_13362);
nand U13519 (N_13519,N_13397,N_13358);
and U13520 (N_13520,N_13254,N_13269);
nand U13521 (N_13521,N_13284,N_13244);
and U13522 (N_13522,N_13330,N_13202);
and U13523 (N_13523,N_13329,N_13233);
or U13524 (N_13524,N_13344,N_13302);
and U13525 (N_13525,N_13302,N_13346);
and U13526 (N_13526,N_13258,N_13372);
and U13527 (N_13527,N_13216,N_13315);
and U13528 (N_13528,N_13218,N_13367);
and U13529 (N_13529,N_13349,N_13281);
nand U13530 (N_13530,N_13355,N_13259);
and U13531 (N_13531,N_13299,N_13360);
nand U13532 (N_13532,N_13220,N_13302);
and U13533 (N_13533,N_13231,N_13202);
or U13534 (N_13534,N_13244,N_13255);
nor U13535 (N_13535,N_13331,N_13310);
nand U13536 (N_13536,N_13392,N_13325);
xnor U13537 (N_13537,N_13379,N_13243);
nand U13538 (N_13538,N_13321,N_13251);
nor U13539 (N_13539,N_13329,N_13369);
and U13540 (N_13540,N_13349,N_13271);
or U13541 (N_13541,N_13241,N_13229);
and U13542 (N_13542,N_13228,N_13333);
nand U13543 (N_13543,N_13332,N_13225);
nor U13544 (N_13544,N_13286,N_13361);
and U13545 (N_13545,N_13235,N_13380);
nand U13546 (N_13546,N_13348,N_13346);
nand U13547 (N_13547,N_13397,N_13289);
or U13548 (N_13548,N_13346,N_13318);
nand U13549 (N_13549,N_13337,N_13397);
nor U13550 (N_13550,N_13237,N_13399);
nand U13551 (N_13551,N_13398,N_13355);
and U13552 (N_13552,N_13315,N_13368);
and U13553 (N_13553,N_13285,N_13305);
nor U13554 (N_13554,N_13254,N_13285);
nor U13555 (N_13555,N_13293,N_13221);
nor U13556 (N_13556,N_13242,N_13216);
nand U13557 (N_13557,N_13334,N_13243);
xnor U13558 (N_13558,N_13398,N_13307);
or U13559 (N_13559,N_13245,N_13368);
nor U13560 (N_13560,N_13307,N_13265);
nand U13561 (N_13561,N_13368,N_13318);
xnor U13562 (N_13562,N_13305,N_13330);
or U13563 (N_13563,N_13384,N_13215);
nand U13564 (N_13564,N_13229,N_13280);
and U13565 (N_13565,N_13360,N_13222);
nand U13566 (N_13566,N_13322,N_13222);
and U13567 (N_13567,N_13294,N_13226);
nand U13568 (N_13568,N_13220,N_13370);
nand U13569 (N_13569,N_13259,N_13200);
or U13570 (N_13570,N_13335,N_13354);
xnor U13571 (N_13571,N_13201,N_13384);
nor U13572 (N_13572,N_13388,N_13393);
nor U13573 (N_13573,N_13204,N_13268);
nor U13574 (N_13574,N_13381,N_13346);
or U13575 (N_13575,N_13344,N_13263);
or U13576 (N_13576,N_13299,N_13316);
and U13577 (N_13577,N_13253,N_13388);
nand U13578 (N_13578,N_13223,N_13366);
and U13579 (N_13579,N_13277,N_13279);
nor U13580 (N_13580,N_13359,N_13323);
or U13581 (N_13581,N_13260,N_13215);
or U13582 (N_13582,N_13326,N_13220);
and U13583 (N_13583,N_13203,N_13386);
xor U13584 (N_13584,N_13255,N_13297);
and U13585 (N_13585,N_13243,N_13372);
or U13586 (N_13586,N_13251,N_13301);
and U13587 (N_13587,N_13325,N_13228);
and U13588 (N_13588,N_13210,N_13234);
or U13589 (N_13589,N_13283,N_13370);
or U13590 (N_13590,N_13371,N_13278);
xnor U13591 (N_13591,N_13382,N_13208);
nand U13592 (N_13592,N_13364,N_13260);
and U13593 (N_13593,N_13311,N_13290);
nor U13594 (N_13594,N_13366,N_13276);
nor U13595 (N_13595,N_13340,N_13318);
or U13596 (N_13596,N_13371,N_13207);
xnor U13597 (N_13597,N_13321,N_13303);
and U13598 (N_13598,N_13389,N_13220);
or U13599 (N_13599,N_13279,N_13297);
xnor U13600 (N_13600,N_13509,N_13419);
and U13601 (N_13601,N_13449,N_13573);
xor U13602 (N_13602,N_13426,N_13587);
xor U13603 (N_13603,N_13497,N_13536);
or U13604 (N_13604,N_13579,N_13468);
or U13605 (N_13605,N_13423,N_13567);
and U13606 (N_13606,N_13492,N_13576);
or U13607 (N_13607,N_13584,N_13564);
xnor U13608 (N_13608,N_13515,N_13531);
nor U13609 (N_13609,N_13432,N_13568);
nand U13610 (N_13610,N_13476,N_13465);
or U13611 (N_13611,N_13496,N_13519);
nor U13612 (N_13612,N_13535,N_13439);
nor U13613 (N_13613,N_13478,N_13598);
xor U13614 (N_13614,N_13434,N_13469);
and U13615 (N_13615,N_13402,N_13408);
or U13616 (N_13616,N_13498,N_13559);
nand U13617 (N_13617,N_13597,N_13590);
and U13618 (N_13618,N_13425,N_13595);
nor U13619 (N_13619,N_13473,N_13405);
nor U13620 (N_13620,N_13480,N_13448);
and U13621 (N_13621,N_13470,N_13504);
nor U13622 (N_13622,N_13451,N_13547);
xnor U13623 (N_13623,N_13577,N_13460);
and U13624 (N_13624,N_13548,N_13532);
nand U13625 (N_13625,N_13540,N_13482);
xnor U13626 (N_13626,N_13420,N_13461);
nor U13627 (N_13627,N_13485,N_13544);
and U13628 (N_13628,N_13513,N_13455);
nor U13629 (N_13629,N_13524,N_13593);
nor U13630 (N_13630,N_13569,N_13542);
nor U13631 (N_13631,N_13447,N_13488);
and U13632 (N_13632,N_13436,N_13570);
xor U13633 (N_13633,N_13407,N_13516);
or U13634 (N_13634,N_13546,N_13493);
nor U13635 (N_13635,N_13464,N_13404);
or U13636 (N_13636,N_13526,N_13518);
or U13637 (N_13637,N_13545,N_13591);
xor U13638 (N_13638,N_13517,N_13522);
nor U13639 (N_13639,N_13429,N_13533);
nand U13640 (N_13640,N_13539,N_13512);
and U13641 (N_13641,N_13537,N_13444);
nand U13642 (N_13642,N_13416,N_13400);
and U13643 (N_13643,N_13543,N_13502);
nand U13644 (N_13644,N_13491,N_13463);
and U13645 (N_13645,N_13445,N_13552);
or U13646 (N_13646,N_13521,N_13410);
nand U13647 (N_13647,N_13467,N_13452);
or U13648 (N_13648,N_13549,N_13443);
or U13649 (N_13649,N_13594,N_13553);
and U13650 (N_13650,N_13511,N_13538);
or U13651 (N_13651,N_13421,N_13555);
nor U13652 (N_13652,N_13599,N_13588);
and U13653 (N_13653,N_13474,N_13486);
or U13654 (N_13654,N_13471,N_13574);
nor U13655 (N_13655,N_13582,N_13453);
or U13656 (N_13656,N_13417,N_13572);
nand U13657 (N_13657,N_13575,N_13418);
or U13658 (N_13658,N_13412,N_13438);
or U13659 (N_13659,N_13456,N_13413);
nand U13660 (N_13660,N_13446,N_13437);
nor U13661 (N_13661,N_13483,N_13490);
or U13662 (N_13662,N_13583,N_13571);
and U13663 (N_13663,N_13523,N_13528);
and U13664 (N_13664,N_13581,N_13501);
nand U13665 (N_13665,N_13578,N_13435);
xnor U13666 (N_13666,N_13508,N_13565);
nand U13667 (N_13667,N_13529,N_13563);
and U13668 (N_13668,N_13477,N_13457);
and U13669 (N_13669,N_13494,N_13415);
and U13670 (N_13670,N_13514,N_13550);
xor U13671 (N_13671,N_13414,N_13585);
nand U13672 (N_13672,N_13479,N_13558);
and U13673 (N_13673,N_13454,N_13505);
or U13674 (N_13674,N_13527,N_13442);
nand U13675 (N_13675,N_13431,N_13566);
xor U13676 (N_13676,N_13433,N_13541);
and U13677 (N_13677,N_13458,N_13589);
xnor U13678 (N_13678,N_13520,N_13462);
nor U13679 (N_13679,N_13551,N_13510);
nor U13680 (N_13680,N_13554,N_13409);
and U13681 (N_13681,N_13596,N_13489);
xor U13682 (N_13682,N_13401,N_13561);
xor U13683 (N_13683,N_13411,N_13481);
or U13684 (N_13684,N_13427,N_13495);
and U13685 (N_13685,N_13534,N_13484);
or U13686 (N_13686,N_13450,N_13586);
xnor U13687 (N_13687,N_13406,N_13503);
xnor U13688 (N_13688,N_13440,N_13530);
nor U13689 (N_13689,N_13506,N_13592);
and U13690 (N_13690,N_13499,N_13459);
nand U13691 (N_13691,N_13580,N_13441);
xor U13692 (N_13692,N_13424,N_13487);
nor U13693 (N_13693,N_13475,N_13525);
and U13694 (N_13694,N_13562,N_13428);
nand U13695 (N_13695,N_13403,N_13557);
nor U13696 (N_13696,N_13500,N_13472);
and U13697 (N_13697,N_13556,N_13560);
nand U13698 (N_13698,N_13422,N_13466);
and U13699 (N_13699,N_13507,N_13430);
and U13700 (N_13700,N_13547,N_13452);
and U13701 (N_13701,N_13515,N_13525);
and U13702 (N_13702,N_13587,N_13507);
xor U13703 (N_13703,N_13514,N_13560);
and U13704 (N_13704,N_13567,N_13525);
nand U13705 (N_13705,N_13499,N_13445);
nor U13706 (N_13706,N_13526,N_13535);
or U13707 (N_13707,N_13526,N_13540);
nor U13708 (N_13708,N_13479,N_13546);
or U13709 (N_13709,N_13501,N_13552);
xnor U13710 (N_13710,N_13501,N_13458);
or U13711 (N_13711,N_13426,N_13434);
or U13712 (N_13712,N_13561,N_13468);
nand U13713 (N_13713,N_13414,N_13438);
nor U13714 (N_13714,N_13478,N_13534);
nor U13715 (N_13715,N_13418,N_13507);
nand U13716 (N_13716,N_13486,N_13480);
nand U13717 (N_13717,N_13501,N_13404);
nor U13718 (N_13718,N_13431,N_13447);
or U13719 (N_13719,N_13560,N_13527);
and U13720 (N_13720,N_13527,N_13464);
nor U13721 (N_13721,N_13582,N_13591);
nor U13722 (N_13722,N_13562,N_13432);
nand U13723 (N_13723,N_13428,N_13408);
or U13724 (N_13724,N_13598,N_13564);
or U13725 (N_13725,N_13442,N_13559);
and U13726 (N_13726,N_13595,N_13496);
nand U13727 (N_13727,N_13440,N_13497);
or U13728 (N_13728,N_13425,N_13465);
and U13729 (N_13729,N_13491,N_13530);
nor U13730 (N_13730,N_13452,N_13490);
xnor U13731 (N_13731,N_13589,N_13548);
nand U13732 (N_13732,N_13539,N_13533);
nor U13733 (N_13733,N_13553,N_13468);
and U13734 (N_13734,N_13530,N_13497);
and U13735 (N_13735,N_13560,N_13454);
nand U13736 (N_13736,N_13417,N_13405);
or U13737 (N_13737,N_13516,N_13421);
and U13738 (N_13738,N_13473,N_13577);
nor U13739 (N_13739,N_13496,N_13511);
and U13740 (N_13740,N_13550,N_13427);
nor U13741 (N_13741,N_13414,N_13535);
or U13742 (N_13742,N_13563,N_13441);
and U13743 (N_13743,N_13533,N_13415);
or U13744 (N_13744,N_13597,N_13587);
nor U13745 (N_13745,N_13474,N_13566);
and U13746 (N_13746,N_13561,N_13515);
or U13747 (N_13747,N_13497,N_13408);
xnor U13748 (N_13748,N_13476,N_13471);
nand U13749 (N_13749,N_13557,N_13503);
nor U13750 (N_13750,N_13474,N_13572);
nor U13751 (N_13751,N_13498,N_13530);
or U13752 (N_13752,N_13509,N_13457);
nor U13753 (N_13753,N_13411,N_13476);
or U13754 (N_13754,N_13478,N_13500);
and U13755 (N_13755,N_13552,N_13425);
nand U13756 (N_13756,N_13550,N_13408);
nor U13757 (N_13757,N_13587,N_13434);
nand U13758 (N_13758,N_13483,N_13574);
nand U13759 (N_13759,N_13571,N_13564);
nor U13760 (N_13760,N_13578,N_13580);
and U13761 (N_13761,N_13578,N_13442);
and U13762 (N_13762,N_13591,N_13593);
nor U13763 (N_13763,N_13490,N_13495);
or U13764 (N_13764,N_13459,N_13509);
nor U13765 (N_13765,N_13405,N_13430);
or U13766 (N_13766,N_13577,N_13558);
nand U13767 (N_13767,N_13519,N_13557);
nor U13768 (N_13768,N_13429,N_13454);
nand U13769 (N_13769,N_13515,N_13439);
and U13770 (N_13770,N_13496,N_13477);
nor U13771 (N_13771,N_13567,N_13417);
and U13772 (N_13772,N_13459,N_13559);
nor U13773 (N_13773,N_13418,N_13528);
nor U13774 (N_13774,N_13547,N_13453);
or U13775 (N_13775,N_13586,N_13519);
or U13776 (N_13776,N_13494,N_13483);
and U13777 (N_13777,N_13420,N_13512);
and U13778 (N_13778,N_13509,N_13489);
or U13779 (N_13779,N_13582,N_13540);
nand U13780 (N_13780,N_13595,N_13579);
nand U13781 (N_13781,N_13490,N_13421);
or U13782 (N_13782,N_13458,N_13560);
and U13783 (N_13783,N_13499,N_13477);
nand U13784 (N_13784,N_13419,N_13404);
nand U13785 (N_13785,N_13500,N_13573);
or U13786 (N_13786,N_13515,N_13516);
nor U13787 (N_13787,N_13463,N_13568);
or U13788 (N_13788,N_13508,N_13513);
or U13789 (N_13789,N_13513,N_13495);
nor U13790 (N_13790,N_13511,N_13582);
and U13791 (N_13791,N_13591,N_13434);
nand U13792 (N_13792,N_13499,N_13418);
or U13793 (N_13793,N_13507,N_13452);
or U13794 (N_13794,N_13538,N_13451);
nand U13795 (N_13795,N_13586,N_13549);
nor U13796 (N_13796,N_13526,N_13439);
and U13797 (N_13797,N_13556,N_13526);
nand U13798 (N_13798,N_13544,N_13474);
nor U13799 (N_13799,N_13453,N_13576);
and U13800 (N_13800,N_13774,N_13716);
xor U13801 (N_13801,N_13617,N_13701);
and U13802 (N_13802,N_13642,N_13620);
nand U13803 (N_13803,N_13682,N_13687);
nor U13804 (N_13804,N_13672,N_13768);
nand U13805 (N_13805,N_13700,N_13683);
and U13806 (N_13806,N_13624,N_13669);
nor U13807 (N_13807,N_13798,N_13639);
nand U13808 (N_13808,N_13638,N_13660);
nand U13809 (N_13809,N_13741,N_13753);
nand U13810 (N_13810,N_13732,N_13622);
nor U13811 (N_13811,N_13695,N_13725);
or U13812 (N_13812,N_13750,N_13793);
and U13813 (N_13813,N_13608,N_13693);
xnor U13814 (N_13814,N_13627,N_13677);
nor U13815 (N_13815,N_13663,N_13796);
nand U13816 (N_13816,N_13717,N_13618);
and U13817 (N_13817,N_13604,N_13742);
and U13818 (N_13818,N_13715,N_13654);
nor U13819 (N_13819,N_13691,N_13727);
nand U13820 (N_13820,N_13760,N_13605);
and U13821 (N_13821,N_13799,N_13646);
or U13822 (N_13822,N_13662,N_13752);
or U13823 (N_13823,N_13771,N_13671);
or U13824 (N_13824,N_13609,N_13712);
or U13825 (N_13825,N_13761,N_13785);
xnor U13826 (N_13826,N_13759,N_13783);
nand U13827 (N_13827,N_13674,N_13643);
nor U13828 (N_13828,N_13626,N_13612);
and U13829 (N_13829,N_13737,N_13724);
nor U13830 (N_13830,N_13728,N_13644);
and U13831 (N_13831,N_13762,N_13603);
xnor U13832 (N_13832,N_13679,N_13681);
xnor U13833 (N_13833,N_13630,N_13794);
nor U13834 (N_13834,N_13777,N_13778);
or U13835 (N_13835,N_13616,N_13692);
or U13836 (N_13836,N_13703,N_13685);
and U13837 (N_13837,N_13606,N_13659);
and U13838 (N_13838,N_13720,N_13655);
and U13839 (N_13839,N_13614,N_13600);
and U13840 (N_13840,N_13640,N_13673);
and U13841 (N_13841,N_13730,N_13786);
and U13842 (N_13842,N_13754,N_13675);
nor U13843 (N_13843,N_13729,N_13756);
or U13844 (N_13844,N_13686,N_13629);
or U13845 (N_13845,N_13763,N_13628);
nor U13846 (N_13846,N_13775,N_13632);
nand U13847 (N_13847,N_13634,N_13631);
nor U13848 (N_13848,N_13765,N_13792);
and U13849 (N_13849,N_13713,N_13784);
nor U13850 (N_13850,N_13702,N_13667);
nand U13851 (N_13851,N_13748,N_13745);
and U13852 (N_13852,N_13633,N_13647);
and U13853 (N_13853,N_13619,N_13708);
and U13854 (N_13854,N_13688,N_13743);
and U13855 (N_13855,N_13615,N_13607);
nor U13856 (N_13856,N_13719,N_13650);
nand U13857 (N_13857,N_13779,N_13711);
and U13858 (N_13858,N_13689,N_13721);
and U13859 (N_13859,N_13645,N_13714);
nor U13860 (N_13860,N_13731,N_13769);
nor U13861 (N_13861,N_13718,N_13749);
nor U13862 (N_13862,N_13698,N_13623);
nor U13863 (N_13863,N_13770,N_13625);
or U13864 (N_13864,N_13664,N_13736);
nor U13865 (N_13865,N_13795,N_13680);
and U13866 (N_13866,N_13746,N_13641);
or U13867 (N_13867,N_13670,N_13791);
xnor U13868 (N_13868,N_13649,N_13757);
or U13869 (N_13869,N_13772,N_13790);
nand U13870 (N_13870,N_13707,N_13697);
and U13871 (N_13871,N_13788,N_13676);
and U13872 (N_13872,N_13758,N_13658);
nor U13873 (N_13873,N_13723,N_13767);
nor U13874 (N_13874,N_13696,N_13656);
nor U13875 (N_13875,N_13613,N_13665);
nor U13876 (N_13876,N_13709,N_13602);
and U13877 (N_13877,N_13611,N_13747);
or U13878 (N_13878,N_13678,N_13706);
or U13879 (N_13879,N_13652,N_13797);
nor U13880 (N_13880,N_13726,N_13601);
xnor U13881 (N_13881,N_13636,N_13635);
xnor U13882 (N_13882,N_13739,N_13699);
nand U13883 (N_13883,N_13684,N_13735);
nor U13884 (N_13884,N_13648,N_13690);
or U13885 (N_13885,N_13766,N_13637);
nand U13886 (N_13886,N_13734,N_13751);
xor U13887 (N_13887,N_13755,N_13789);
nor U13888 (N_13888,N_13781,N_13651);
xnor U13889 (N_13889,N_13661,N_13738);
and U13890 (N_13890,N_13782,N_13710);
nand U13891 (N_13891,N_13780,N_13668);
xor U13892 (N_13892,N_13773,N_13787);
and U13893 (N_13893,N_13657,N_13764);
and U13894 (N_13894,N_13733,N_13621);
and U13895 (N_13895,N_13666,N_13610);
nor U13896 (N_13896,N_13776,N_13705);
nand U13897 (N_13897,N_13722,N_13704);
or U13898 (N_13898,N_13740,N_13653);
and U13899 (N_13899,N_13694,N_13744);
nor U13900 (N_13900,N_13667,N_13768);
or U13901 (N_13901,N_13767,N_13618);
or U13902 (N_13902,N_13679,N_13633);
and U13903 (N_13903,N_13731,N_13723);
nand U13904 (N_13904,N_13707,N_13726);
nand U13905 (N_13905,N_13721,N_13722);
nand U13906 (N_13906,N_13641,N_13793);
xor U13907 (N_13907,N_13649,N_13784);
and U13908 (N_13908,N_13613,N_13733);
nand U13909 (N_13909,N_13605,N_13631);
nand U13910 (N_13910,N_13734,N_13779);
nor U13911 (N_13911,N_13629,N_13777);
nor U13912 (N_13912,N_13601,N_13618);
nor U13913 (N_13913,N_13741,N_13717);
or U13914 (N_13914,N_13779,N_13692);
xnor U13915 (N_13915,N_13629,N_13794);
and U13916 (N_13916,N_13673,N_13637);
nand U13917 (N_13917,N_13719,N_13759);
xnor U13918 (N_13918,N_13725,N_13786);
and U13919 (N_13919,N_13791,N_13701);
xor U13920 (N_13920,N_13741,N_13618);
or U13921 (N_13921,N_13631,N_13790);
nand U13922 (N_13922,N_13723,N_13774);
or U13923 (N_13923,N_13611,N_13641);
or U13924 (N_13924,N_13648,N_13666);
nand U13925 (N_13925,N_13660,N_13729);
and U13926 (N_13926,N_13621,N_13623);
nor U13927 (N_13927,N_13723,N_13715);
nor U13928 (N_13928,N_13712,N_13720);
and U13929 (N_13929,N_13771,N_13754);
and U13930 (N_13930,N_13627,N_13736);
nor U13931 (N_13931,N_13697,N_13693);
xnor U13932 (N_13932,N_13778,N_13688);
nand U13933 (N_13933,N_13711,N_13614);
or U13934 (N_13934,N_13675,N_13739);
nor U13935 (N_13935,N_13654,N_13747);
nor U13936 (N_13936,N_13728,N_13668);
and U13937 (N_13937,N_13752,N_13729);
nand U13938 (N_13938,N_13663,N_13757);
or U13939 (N_13939,N_13624,N_13751);
nor U13940 (N_13940,N_13711,N_13645);
xor U13941 (N_13941,N_13620,N_13733);
or U13942 (N_13942,N_13665,N_13695);
or U13943 (N_13943,N_13603,N_13742);
nand U13944 (N_13944,N_13627,N_13718);
xor U13945 (N_13945,N_13612,N_13642);
nor U13946 (N_13946,N_13788,N_13614);
and U13947 (N_13947,N_13776,N_13739);
or U13948 (N_13948,N_13721,N_13751);
nand U13949 (N_13949,N_13665,N_13740);
xnor U13950 (N_13950,N_13766,N_13735);
or U13951 (N_13951,N_13795,N_13760);
and U13952 (N_13952,N_13626,N_13750);
nand U13953 (N_13953,N_13684,N_13726);
and U13954 (N_13954,N_13798,N_13789);
or U13955 (N_13955,N_13622,N_13675);
and U13956 (N_13956,N_13640,N_13651);
nor U13957 (N_13957,N_13770,N_13799);
nor U13958 (N_13958,N_13619,N_13731);
and U13959 (N_13959,N_13633,N_13684);
or U13960 (N_13960,N_13642,N_13619);
nand U13961 (N_13961,N_13775,N_13753);
nor U13962 (N_13962,N_13710,N_13770);
nand U13963 (N_13963,N_13747,N_13691);
or U13964 (N_13964,N_13697,N_13701);
nor U13965 (N_13965,N_13725,N_13763);
nand U13966 (N_13966,N_13697,N_13685);
or U13967 (N_13967,N_13784,N_13611);
or U13968 (N_13968,N_13653,N_13646);
nand U13969 (N_13969,N_13660,N_13721);
and U13970 (N_13970,N_13704,N_13777);
nand U13971 (N_13971,N_13767,N_13638);
nand U13972 (N_13972,N_13698,N_13765);
or U13973 (N_13973,N_13782,N_13663);
nor U13974 (N_13974,N_13773,N_13634);
nor U13975 (N_13975,N_13659,N_13728);
nand U13976 (N_13976,N_13782,N_13780);
nand U13977 (N_13977,N_13783,N_13785);
xnor U13978 (N_13978,N_13715,N_13779);
and U13979 (N_13979,N_13702,N_13705);
and U13980 (N_13980,N_13657,N_13694);
or U13981 (N_13981,N_13697,N_13754);
and U13982 (N_13982,N_13753,N_13695);
xor U13983 (N_13983,N_13704,N_13689);
and U13984 (N_13984,N_13788,N_13658);
and U13985 (N_13985,N_13620,N_13649);
and U13986 (N_13986,N_13662,N_13722);
xnor U13987 (N_13987,N_13748,N_13792);
nand U13988 (N_13988,N_13687,N_13619);
or U13989 (N_13989,N_13773,N_13716);
and U13990 (N_13990,N_13631,N_13717);
or U13991 (N_13991,N_13785,N_13688);
or U13992 (N_13992,N_13685,N_13712);
nor U13993 (N_13993,N_13636,N_13695);
or U13994 (N_13994,N_13689,N_13750);
nand U13995 (N_13995,N_13633,N_13641);
and U13996 (N_13996,N_13664,N_13796);
and U13997 (N_13997,N_13620,N_13646);
or U13998 (N_13998,N_13725,N_13735);
and U13999 (N_13999,N_13762,N_13668);
or U14000 (N_14000,N_13816,N_13900);
nor U14001 (N_14001,N_13889,N_13978);
xnor U14002 (N_14002,N_13881,N_13872);
nand U14003 (N_14003,N_13829,N_13932);
or U14004 (N_14004,N_13961,N_13813);
nand U14005 (N_14005,N_13864,N_13967);
nor U14006 (N_14006,N_13937,N_13853);
or U14007 (N_14007,N_13875,N_13976);
or U14008 (N_14008,N_13955,N_13877);
and U14009 (N_14009,N_13847,N_13858);
and U14010 (N_14010,N_13959,N_13926);
and U14011 (N_14011,N_13838,N_13815);
nand U14012 (N_14012,N_13820,N_13998);
and U14013 (N_14013,N_13972,N_13854);
xnor U14014 (N_14014,N_13894,N_13845);
or U14015 (N_14015,N_13859,N_13874);
xor U14016 (N_14016,N_13835,N_13962);
or U14017 (N_14017,N_13928,N_13837);
and U14018 (N_14018,N_13867,N_13819);
and U14019 (N_14019,N_13991,N_13985);
nand U14020 (N_14020,N_13974,N_13933);
and U14021 (N_14021,N_13901,N_13949);
or U14022 (N_14022,N_13929,N_13812);
or U14023 (N_14023,N_13899,N_13860);
or U14024 (N_14024,N_13992,N_13944);
and U14025 (N_14025,N_13965,N_13897);
or U14026 (N_14026,N_13830,N_13996);
nor U14027 (N_14027,N_13927,N_13903);
or U14028 (N_14028,N_13803,N_13869);
and U14029 (N_14029,N_13828,N_13873);
and U14030 (N_14030,N_13841,N_13988);
nand U14031 (N_14031,N_13836,N_13993);
nor U14032 (N_14032,N_13947,N_13910);
nor U14033 (N_14033,N_13811,N_13823);
nor U14034 (N_14034,N_13876,N_13986);
nand U14035 (N_14035,N_13930,N_13878);
or U14036 (N_14036,N_13826,N_13807);
nor U14037 (N_14037,N_13902,N_13895);
and U14038 (N_14038,N_13935,N_13925);
nand U14039 (N_14039,N_13981,N_13865);
nand U14040 (N_14040,N_13920,N_13977);
nor U14041 (N_14041,N_13891,N_13942);
or U14042 (N_14042,N_13863,N_13958);
and U14043 (N_14043,N_13890,N_13801);
nor U14044 (N_14044,N_13952,N_13898);
nor U14045 (N_14045,N_13851,N_13866);
or U14046 (N_14046,N_13934,N_13896);
or U14047 (N_14047,N_13954,N_13808);
nor U14048 (N_14048,N_13999,N_13868);
nor U14049 (N_14049,N_13887,N_13862);
nor U14050 (N_14050,N_13916,N_13906);
nor U14051 (N_14051,N_13914,N_13817);
nand U14052 (N_14052,N_13964,N_13923);
and U14053 (N_14053,N_13907,N_13971);
or U14054 (N_14054,N_13941,N_13884);
xnor U14055 (N_14055,N_13832,N_13982);
or U14056 (N_14056,N_13979,N_13800);
or U14057 (N_14057,N_13886,N_13945);
and U14058 (N_14058,N_13919,N_13973);
nand U14059 (N_14059,N_13905,N_13963);
or U14060 (N_14060,N_13983,N_13844);
nand U14061 (N_14061,N_13822,N_13839);
nand U14062 (N_14062,N_13911,N_13833);
xor U14063 (N_14063,N_13946,N_13805);
or U14064 (N_14064,N_13918,N_13957);
xnor U14065 (N_14065,N_13912,N_13960);
nand U14066 (N_14066,N_13809,N_13968);
nand U14067 (N_14067,N_13825,N_13857);
and U14068 (N_14068,N_13909,N_13931);
xor U14069 (N_14069,N_13850,N_13995);
nand U14070 (N_14070,N_13969,N_13888);
or U14071 (N_14071,N_13938,N_13882);
nand U14072 (N_14072,N_13831,N_13871);
nand U14073 (N_14073,N_13917,N_13943);
or U14074 (N_14074,N_13856,N_13810);
nand U14075 (N_14075,N_13921,N_13843);
nand U14076 (N_14076,N_13870,N_13852);
xor U14077 (N_14077,N_13861,N_13802);
nor U14078 (N_14078,N_13818,N_13885);
and U14079 (N_14079,N_13940,N_13970);
nor U14080 (N_14080,N_13989,N_13994);
xor U14081 (N_14081,N_13879,N_13924);
and U14082 (N_14082,N_13980,N_13827);
nand U14083 (N_14083,N_13922,N_13880);
and U14084 (N_14084,N_13848,N_13990);
nor U14085 (N_14085,N_13953,N_13950);
nand U14086 (N_14086,N_13948,N_13855);
or U14087 (N_14087,N_13956,N_13904);
nor U14088 (N_14088,N_13987,N_13893);
nand U14089 (N_14089,N_13840,N_13915);
nand U14090 (N_14090,N_13939,N_13966);
nand U14091 (N_14091,N_13908,N_13821);
nor U14092 (N_14092,N_13849,N_13834);
or U14093 (N_14093,N_13975,N_13806);
or U14094 (N_14094,N_13814,N_13936);
and U14095 (N_14095,N_13804,N_13984);
nor U14096 (N_14096,N_13997,N_13951);
nand U14097 (N_14097,N_13846,N_13883);
nand U14098 (N_14098,N_13824,N_13842);
nor U14099 (N_14099,N_13892,N_13913);
nor U14100 (N_14100,N_13866,N_13846);
and U14101 (N_14101,N_13815,N_13967);
nand U14102 (N_14102,N_13826,N_13843);
and U14103 (N_14103,N_13864,N_13856);
nor U14104 (N_14104,N_13915,N_13878);
nand U14105 (N_14105,N_13851,N_13902);
and U14106 (N_14106,N_13978,N_13970);
and U14107 (N_14107,N_13886,N_13969);
nand U14108 (N_14108,N_13924,N_13846);
xor U14109 (N_14109,N_13849,N_13922);
nand U14110 (N_14110,N_13918,N_13901);
nor U14111 (N_14111,N_13923,N_13986);
xor U14112 (N_14112,N_13878,N_13920);
nor U14113 (N_14113,N_13843,N_13802);
nor U14114 (N_14114,N_13923,N_13845);
nand U14115 (N_14115,N_13898,N_13922);
nor U14116 (N_14116,N_13842,N_13870);
nor U14117 (N_14117,N_13811,N_13833);
nand U14118 (N_14118,N_13802,N_13999);
nor U14119 (N_14119,N_13871,N_13992);
nand U14120 (N_14120,N_13866,N_13834);
nor U14121 (N_14121,N_13937,N_13913);
nand U14122 (N_14122,N_13904,N_13813);
or U14123 (N_14123,N_13904,N_13880);
nor U14124 (N_14124,N_13865,N_13882);
or U14125 (N_14125,N_13876,N_13971);
nand U14126 (N_14126,N_13863,N_13868);
nand U14127 (N_14127,N_13834,N_13855);
or U14128 (N_14128,N_13892,N_13868);
nor U14129 (N_14129,N_13840,N_13812);
nor U14130 (N_14130,N_13899,N_13820);
nand U14131 (N_14131,N_13889,N_13929);
nor U14132 (N_14132,N_13860,N_13854);
and U14133 (N_14133,N_13893,N_13810);
nor U14134 (N_14134,N_13925,N_13972);
nor U14135 (N_14135,N_13956,N_13909);
and U14136 (N_14136,N_13916,N_13983);
nor U14137 (N_14137,N_13926,N_13850);
xor U14138 (N_14138,N_13928,N_13954);
nand U14139 (N_14139,N_13852,N_13805);
and U14140 (N_14140,N_13989,N_13895);
nor U14141 (N_14141,N_13953,N_13851);
nor U14142 (N_14142,N_13811,N_13880);
nand U14143 (N_14143,N_13839,N_13971);
or U14144 (N_14144,N_13822,N_13901);
nor U14145 (N_14145,N_13860,N_13916);
and U14146 (N_14146,N_13841,N_13809);
or U14147 (N_14147,N_13809,N_13898);
or U14148 (N_14148,N_13855,N_13991);
nor U14149 (N_14149,N_13838,N_13988);
or U14150 (N_14150,N_13897,N_13874);
nand U14151 (N_14151,N_13905,N_13863);
or U14152 (N_14152,N_13902,N_13984);
nor U14153 (N_14153,N_13992,N_13876);
or U14154 (N_14154,N_13947,N_13933);
nand U14155 (N_14155,N_13982,N_13824);
and U14156 (N_14156,N_13943,N_13954);
nand U14157 (N_14157,N_13829,N_13906);
nand U14158 (N_14158,N_13982,N_13921);
nand U14159 (N_14159,N_13980,N_13922);
nand U14160 (N_14160,N_13960,N_13844);
nand U14161 (N_14161,N_13967,N_13883);
or U14162 (N_14162,N_13856,N_13960);
xnor U14163 (N_14163,N_13831,N_13925);
and U14164 (N_14164,N_13960,N_13880);
or U14165 (N_14165,N_13890,N_13850);
or U14166 (N_14166,N_13887,N_13873);
and U14167 (N_14167,N_13971,N_13836);
and U14168 (N_14168,N_13926,N_13810);
nor U14169 (N_14169,N_13897,N_13995);
nor U14170 (N_14170,N_13846,N_13936);
nand U14171 (N_14171,N_13988,N_13980);
or U14172 (N_14172,N_13996,N_13845);
nand U14173 (N_14173,N_13808,N_13826);
or U14174 (N_14174,N_13960,N_13816);
and U14175 (N_14175,N_13816,N_13877);
nand U14176 (N_14176,N_13961,N_13851);
nor U14177 (N_14177,N_13829,N_13925);
and U14178 (N_14178,N_13936,N_13945);
and U14179 (N_14179,N_13871,N_13824);
nor U14180 (N_14180,N_13830,N_13991);
and U14181 (N_14181,N_13889,N_13911);
nand U14182 (N_14182,N_13914,N_13896);
and U14183 (N_14183,N_13876,N_13961);
nor U14184 (N_14184,N_13950,N_13801);
and U14185 (N_14185,N_13970,N_13960);
nor U14186 (N_14186,N_13877,N_13845);
and U14187 (N_14187,N_13894,N_13973);
and U14188 (N_14188,N_13924,N_13959);
and U14189 (N_14189,N_13935,N_13885);
and U14190 (N_14190,N_13956,N_13942);
or U14191 (N_14191,N_13893,N_13885);
or U14192 (N_14192,N_13825,N_13946);
nand U14193 (N_14193,N_13991,N_13929);
nor U14194 (N_14194,N_13852,N_13926);
nor U14195 (N_14195,N_13896,N_13929);
or U14196 (N_14196,N_13897,N_13831);
xor U14197 (N_14197,N_13814,N_13857);
nor U14198 (N_14198,N_13849,N_13815);
xnor U14199 (N_14199,N_13948,N_13972);
nor U14200 (N_14200,N_14162,N_14106);
and U14201 (N_14201,N_14036,N_14142);
or U14202 (N_14202,N_14035,N_14098);
nor U14203 (N_14203,N_14049,N_14050);
nand U14204 (N_14204,N_14132,N_14061);
and U14205 (N_14205,N_14135,N_14021);
nor U14206 (N_14206,N_14187,N_14065);
or U14207 (N_14207,N_14121,N_14034);
xnor U14208 (N_14208,N_14137,N_14066);
xnor U14209 (N_14209,N_14019,N_14198);
and U14210 (N_14210,N_14016,N_14017);
nand U14211 (N_14211,N_14155,N_14192);
and U14212 (N_14212,N_14100,N_14179);
and U14213 (N_14213,N_14060,N_14153);
or U14214 (N_14214,N_14040,N_14150);
nand U14215 (N_14215,N_14174,N_14189);
nand U14216 (N_14216,N_14018,N_14148);
nor U14217 (N_14217,N_14119,N_14003);
and U14218 (N_14218,N_14094,N_14133);
or U14219 (N_14219,N_14127,N_14180);
nand U14220 (N_14220,N_14058,N_14123);
or U14221 (N_14221,N_14023,N_14012);
nand U14222 (N_14222,N_14059,N_14011);
and U14223 (N_14223,N_14159,N_14128);
nand U14224 (N_14224,N_14184,N_14157);
and U14225 (N_14225,N_14062,N_14074);
xnor U14226 (N_14226,N_14197,N_14047);
nand U14227 (N_14227,N_14120,N_14084);
and U14228 (N_14228,N_14130,N_14093);
and U14229 (N_14229,N_14168,N_14196);
nor U14230 (N_14230,N_14090,N_14178);
and U14231 (N_14231,N_14082,N_14113);
and U14232 (N_14232,N_14027,N_14083);
xor U14233 (N_14233,N_14139,N_14185);
and U14234 (N_14234,N_14086,N_14095);
and U14235 (N_14235,N_14020,N_14126);
or U14236 (N_14236,N_14075,N_14158);
or U14237 (N_14237,N_14193,N_14073);
or U14238 (N_14238,N_14048,N_14181);
nor U14239 (N_14239,N_14186,N_14001);
and U14240 (N_14240,N_14068,N_14136);
or U14241 (N_14241,N_14109,N_14134);
nor U14242 (N_14242,N_14164,N_14055);
or U14243 (N_14243,N_14102,N_14144);
xnor U14244 (N_14244,N_14010,N_14039);
nand U14245 (N_14245,N_14097,N_14077);
nand U14246 (N_14246,N_14072,N_14101);
and U14247 (N_14247,N_14007,N_14088);
nand U14248 (N_14248,N_14115,N_14152);
nor U14249 (N_14249,N_14188,N_14052);
nand U14250 (N_14250,N_14080,N_14116);
and U14251 (N_14251,N_14042,N_14037);
nand U14252 (N_14252,N_14167,N_14151);
nor U14253 (N_14253,N_14006,N_14125);
nor U14254 (N_14254,N_14025,N_14044);
nor U14255 (N_14255,N_14004,N_14029);
nor U14256 (N_14256,N_14014,N_14149);
nor U14257 (N_14257,N_14057,N_14046);
nor U14258 (N_14258,N_14013,N_14110);
and U14259 (N_14259,N_14079,N_14063);
nand U14260 (N_14260,N_14026,N_14111);
and U14261 (N_14261,N_14114,N_14096);
nand U14262 (N_14262,N_14173,N_14070);
nor U14263 (N_14263,N_14030,N_14069);
and U14264 (N_14264,N_14032,N_14122);
nand U14265 (N_14265,N_14108,N_14024);
nand U14266 (N_14266,N_14161,N_14031);
or U14267 (N_14267,N_14056,N_14131);
nor U14268 (N_14268,N_14163,N_14118);
and U14269 (N_14269,N_14195,N_14071);
nor U14270 (N_14270,N_14076,N_14022);
nor U14271 (N_14271,N_14138,N_14183);
and U14272 (N_14272,N_14028,N_14087);
and U14273 (N_14273,N_14041,N_14160);
nand U14274 (N_14274,N_14140,N_14091);
nor U14275 (N_14275,N_14085,N_14166);
nand U14276 (N_14276,N_14117,N_14154);
nand U14277 (N_14277,N_14067,N_14043);
nor U14278 (N_14278,N_14182,N_14107);
nand U14279 (N_14279,N_14005,N_14078);
and U14280 (N_14280,N_14143,N_14053);
nor U14281 (N_14281,N_14000,N_14105);
nor U14282 (N_14282,N_14172,N_14176);
and U14283 (N_14283,N_14194,N_14051);
nor U14284 (N_14284,N_14104,N_14015);
or U14285 (N_14285,N_14054,N_14190);
nor U14286 (N_14286,N_14146,N_14169);
nor U14287 (N_14287,N_14177,N_14145);
nor U14288 (N_14288,N_14165,N_14064);
or U14289 (N_14289,N_14175,N_14038);
or U14290 (N_14290,N_14002,N_14099);
xor U14291 (N_14291,N_14170,N_14141);
and U14292 (N_14292,N_14199,N_14129);
nor U14293 (N_14293,N_14191,N_14081);
nor U14294 (N_14294,N_14092,N_14124);
nor U14295 (N_14295,N_14045,N_14008);
or U14296 (N_14296,N_14171,N_14089);
nor U14297 (N_14297,N_14009,N_14147);
and U14298 (N_14298,N_14156,N_14033);
and U14299 (N_14299,N_14112,N_14103);
nand U14300 (N_14300,N_14059,N_14028);
nand U14301 (N_14301,N_14161,N_14140);
or U14302 (N_14302,N_14145,N_14092);
or U14303 (N_14303,N_14126,N_14035);
or U14304 (N_14304,N_14052,N_14135);
or U14305 (N_14305,N_14167,N_14047);
nand U14306 (N_14306,N_14036,N_14132);
nand U14307 (N_14307,N_14175,N_14088);
and U14308 (N_14308,N_14082,N_14019);
xor U14309 (N_14309,N_14131,N_14127);
or U14310 (N_14310,N_14124,N_14105);
xnor U14311 (N_14311,N_14018,N_14058);
xnor U14312 (N_14312,N_14152,N_14055);
and U14313 (N_14313,N_14131,N_14161);
and U14314 (N_14314,N_14046,N_14044);
nor U14315 (N_14315,N_14011,N_14164);
nor U14316 (N_14316,N_14149,N_14197);
or U14317 (N_14317,N_14134,N_14091);
or U14318 (N_14318,N_14053,N_14055);
nand U14319 (N_14319,N_14198,N_14026);
nor U14320 (N_14320,N_14126,N_14181);
xor U14321 (N_14321,N_14148,N_14170);
nand U14322 (N_14322,N_14174,N_14198);
nor U14323 (N_14323,N_14047,N_14038);
and U14324 (N_14324,N_14111,N_14098);
nor U14325 (N_14325,N_14014,N_14199);
or U14326 (N_14326,N_14160,N_14021);
and U14327 (N_14327,N_14104,N_14188);
or U14328 (N_14328,N_14065,N_14038);
and U14329 (N_14329,N_14002,N_14184);
or U14330 (N_14330,N_14191,N_14137);
or U14331 (N_14331,N_14144,N_14075);
or U14332 (N_14332,N_14122,N_14177);
nand U14333 (N_14333,N_14040,N_14016);
or U14334 (N_14334,N_14150,N_14048);
and U14335 (N_14335,N_14025,N_14063);
and U14336 (N_14336,N_14133,N_14046);
and U14337 (N_14337,N_14155,N_14058);
and U14338 (N_14338,N_14007,N_14074);
nor U14339 (N_14339,N_14178,N_14097);
or U14340 (N_14340,N_14191,N_14102);
nand U14341 (N_14341,N_14157,N_14148);
and U14342 (N_14342,N_14016,N_14027);
or U14343 (N_14343,N_14147,N_14197);
nand U14344 (N_14344,N_14187,N_14061);
nand U14345 (N_14345,N_14058,N_14032);
nand U14346 (N_14346,N_14039,N_14107);
nand U14347 (N_14347,N_14171,N_14109);
and U14348 (N_14348,N_14161,N_14067);
and U14349 (N_14349,N_14176,N_14106);
and U14350 (N_14350,N_14061,N_14001);
nand U14351 (N_14351,N_14109,N_14094);
nor U14352 (N_14352,N_14152,N_14086);
and U14353 (N_14353,N_14173,N_14159);
or U14354 (N_14354,N_14053,N_14061);
and U14355 (N_14355,N_14122,N_14064);
nor U14356 (N_14356,N_14040,N_14030);
nor U14357 (N_14357,N_14076,N_14171);
nor U14358 (N_14358,N_14001,N_14134);
nand U14359 (N_14359,N_14089,N_14065);
nand U14360 (N_14360,N_14124,N_14189);
nor U14361 (N_14361,N_14131,N_14145);
nand U14362 (N_14362,N_14053,N_14188);
nor U14363 (N_14363,N_14121,N_14011);
and U14364 (N_14364,N_14086,N_14176);
nor U14365 (N_14365,N_14024,N_14163);
or U14366 (N_14366,N_14173,N_14090);
or U14367 (N_14367,N_14132,N_14000);
xnor U14368 (N_14368,N_14042,N_14065);
nor U14369 (N_14369,N_14097,N_14168);
nor U14370 (N_14370,N_14174,N_14004);
nand U14371 (N_14371,N_14094,N_14051);
and U14372 (N_14372,N_14123,N_14096);
nor U14373 (N_14373,N_14133,N_14103);
and U14374 (N_14374,N_14087,N_14129);
or U14375 (N_14375,N_14051,N_14147);
and U14376 (N_14376,N_14036,N_14153);
nor U14377 (N_14377,N_14038,N_14152);
and U14378 (N_14378,N_14008,N_14081);
nor U14379 (N_14379,N_14144,N_14011);
nor U14380 (N_14380,N_14072,N_14198);
or U14381 (N_14381,N_14121,N_14123);
and U14382 (N_14382,N_14066,N_14055);
or U14383 (N_14383,N_14082,N_14030);
nand U14384 (N_14384,N_14115,N_14039);
nand U14385 (N_14385,N_14009,N_14175);
nor U14386 (N_14386,N_14098,N_14091);
nand U14387 (N_14387,N_14055,N_14143);
and U14388 (N_14388,N_14070,N_14091);
xnor U14389 (N_14389,N_14097,N_14115);
or U14390 (N_14390,N_14097,N_14100);
and U14391 (N_14391,N_14047,N_14065);
or U14392 (N_14392,N_14063,N_14164);
or U14393 (N_14393,N_14027,N_14013);
nor U14394 (N_14394,N_14177,N_14149);
and U14395 (N_14395,N_14019,N_14097);
nor U14396 (N_14396,N_14106,N_14192);
nor U14397 (N_14397,N_14025,N_14097);
xnor U14398 (N_14398,N_14102,N_14183);
nor U14399 (N_14399,N_14135,N_14098);
and U14400 (N_14400,N_14305,N_14214);
or U14401 (N_14401,N_14237,N_14346);
nor U14402 (N_14402,N_14368,N_14349);
xor U14403 (N_14403,N_14225,N_14227);
or U14404 (N_14404,N_14200,N_14257);
nand U14405 (N_14405,N_14209,N_14372);
xnor U14406 (N_14406,N_14256,N_14345);
and U14407 (N_14407,N_14394,N_14347);
nor U14408 (N_14408,N_14269,N_14354);
or U14409 (N_14409,N_14247,N_14218);
or U14410 (N_14410,N_14307,N_14204);
nand U14411 (N_14411,N_14250,N_14369);
and U14412 (N_14412,N_14326,N_14212);
and U14413 (N_14413,N_14378,N_14213);
nand U14414 (N_14414,N_14289,N_14344);
and U14415 (N_14415,N_14252,N_14226);
nand U14416 (N_14416,N_14286,N_14365);
or U14417 (N_14417,N_14355,N_14244);
or U14418 (N_14418,N_14366,N_14284);
nand U14419 (N_14419,N_14332,N_14234);
nor U14420 (N_14420,N_14319,N_14374);
nand U14421 (N_14421,N_14334,N_14275);
xnor U14422 (N_14422,N_14208,N_14393);
or U14423 (N_14423,N_14359,N_14240);
or U14424 (N_14424,N_14310,N_14376);
nand U14425 (N_14425,N_14277,N_14395);
and U14426 (N_14426,N_14251,N_14222);
or U14427 (N_14427,N_14341,N_14296);
xor U14428 (N_14428,N_14322,N_14321);
or U14429 (N_14429,N_14232,N_14300);
nand U14430 (N_14430,N_14268,N_14229);
or U14431 (N_14431,N_14398,N_14301);
or U14432 (N_14432,N_14387,N_14331);
or U14433 (N_14433,N_14337,N_14328);
and U14434 (N_14434,N_14375,N_14302);
and U14435 (N_14435,N_14370,N_14217);
xor U14436 (N_14436,N_14392,N_14293);
or U14437 (N_14437,N_14235,N_14338);
or U14438 (N_14438,N_14228,N_14373);
nand U14439 (N_14439,N_14290,N_14243);
nand U14440 (N_14440,N_14390,N_14263);
nand U14441 (N_14441,N_14385,N_14333);
nor U14442 (N_14442,N_14356,N_14327);
nand U14443 (N_14443,N_14242,N_14340);
or U14444 (N_14444,N_14260,N_14231);
or U14445 (N_14445,N_14265,N_14391);
xnor U14446 (N_14446,N_14283,N_14357);
and U14447 (N_14447,N_14303,N_14274);
and U14448 (N_14448,N_14396,N_14270);
nor U14449 (N_14449,N_14239,N_14255);
nand U14450 (N_14450,N_14267,N_14358);
or U14451 (N_14451,N_14371,N_14313);
or U14452 (N_14452,N_14363,N_14353);
xnor U14453 (N_14453,N_14271,N_14224);
nand U14454 (N_14454,N_14367,N_14264);
or U14455 (N_14455,N_14258,N_14291);
nand U14456 (N_14456,N_14248,N_14287);
or U14457 (N_14457,N_14350,N_14273);
or U14458 (N_14458,N_14397,N_14221);
nor U14459 (N_14459,N_14325,N_14384);
or U14460 (N_14460,N_14254,N_14351);
nand U14461 (N_14461,N_14339,N_14329);
or U14462 (N_14462,N_14206,N_14211);
or U14463 (N_14463,N_14377,N_14317);
nand U14464 (N_14464,N_14262,N_14219);
xor U14465 (N_14465,N_14210,N_14246);
and U14466 (N_14466,N_14389,N_14241);
nand U14467 (N_14467,N_14388,N_14223);
nand U14468 (N_14468,N_14323,N_14342);
and U14469 (N_14469,N_14309,N_14207);
nand U14470 (N_14470,N_14295,N_14288);
nand U14471 (N_14471,N_14306,N_14380);
nor U14472 (N_14472,N_14245,N_14299);
nand U14473 (N_14473,N_14201,N_14216);
and U14474 (N_14474,N_14316,N_14318);
nand U14475 (N_14475,N_14364,N_14238);
and U14476 (N_14476,N_14308,N_14203);
or U14477 (N_14477,N_14266,N_14259);
nor U14478 (N_14478,N_14361,N_14381);
and U14479 (N_14479,N_14399,N_14292);
or U14480 (N_14480,N_14320,N_14336);
and U14481 (N_14481,N_14282,N_14297);
or U14482 (N_14482,N_14311,N_14279);
or U14483 (N_14483,N_14314,N_14281);
nand U14484 (N_14484,N_14343,N_14386);
nor U14485 (N_14485,N_14285,N_14324);
and U14486 (N_14486,N_14276,N_14383);
xor U14487 (N_14487,N_14360,N_14312);
and U14488 (N_14488,N_14335,N_14382);
nor U14489 (N_14489,N_14278,N_14249);
nor U14490 (N_14490,N_14362,N_14379);
and U14491 (N_14491,N_14261,N_14352);
nor U14492 (N_14492,N_14236,N_14294);
and U14493 (N_14493,N_14280,N_14298);
and U14494 (N_14494,N_14205,N_14315);
or U14495 (N_14495,N_14202,N_14348);
nor U14496 (N_14496,N_14215,N_14272);
nor U14497 (N_14497,N_14253,N_14304);
nand U14498 (N_14498,N_14330,N_14220);
xor U14499 (N_14499,N_14233,N_14230);
nor U14500 (N_14500,N_14355,N_14251);
nor U14501 (N_14501,N_14260,N_14269);
xnor U14502 (N_14502,N_14383,N_14290);
or U14503 (N_14503,N_14274,N_14271);
or U14504 (N_14504,N_14240,N_14365);
or U14505 (N_14505,N_14357,N_14263);
and U14506 (N_14506,N_14376,N_14365);
nor U14507 (N_14507,N_14347,N_14216);
nor U14508 (N_14508,N_14245,N_14371);
nor U14509 (N_14509,N_14234,N_14389);
and U14510 (N_14510,N_14247,N_14258);
nor U14511 (N_14511,N_14361,N_14313);
and U14512 (N_14512,N_14326,N_14266);
nand U14513 (N_14513,N_14210,N_14252);
nand U14514 (N_14514,N_14360,N_14345);
nand U14515 (N_14515,N_14328,N_14336);
and U14516 (N_14516,N_14318,N_14346);
nor U14517 (N_14517,N_14283,N_14323);
nand U14518 (N_14518,N_14206,N_14231);
and U14519 (N_14519,N_14302,N_14291);
nand U14520 (N_14520,N_14260,N_14200);
nand U14521 (N_14521,N_14240,N_14284);
and U14522 (N_14522,N_14254,N_14296);
and U14523 (N_14523,N_14383,N_14378);
xnor U14524 (N_14524,N_14331,N_14355);
nand U14525 (N_14525,N_14394,N_14208);
and U14526 (N_14526,N_14211,N_14261);
nor U14527 (N_14527,N_14349,N_14257);
nor U14528 (N_14528,N_14294,N_14347);
xor U14529 (N_14529,N_14367,N_14341);
or U14530 (N_14530,N_14207,N_14254);
and U14531 (N_14531,N_14383,N_14287);
and U14532 (N_14532,N_14388,N_14271);
and U14533 (N_14533,N_14219,N_14238);
nand U14534 (N_14534,N_14348,N_14319);
nor U14535 (N_14535,N_14202,N_14337);
nand U14536 (N_14536,N_14331,N_14244);
nand U14537 (N_14537,N_14353,N_14228);
nand U14538 (N_14538,N_14252,N_14302);
and U14539 (N_14539,N_14284,N_14361);
or U14540 (N_14540,N_14275,N_14241);
or U14541 (N_14541,N_14316,N_14256);
nor U14542 (N_14542,N_14356,N_14215);
nand U14543 (N_14543,N_14393,N_14332);
nor U14544 (N_14544,N_14380,N_14256);
nand U14545 (N_14545,N_14204,N_14397);
or U14546 (N_14546,N_14369,N_14318);
or U14547 (N_14547,N_14365,N_14252);
or U14548 (N_14548,N_14388,N_14236);
nand U14549 (N_14549,N_14334,N_14352);
nand U14550 (N_14550,N_14300,N_14356);
and U14551 (N_14551,N_14216,N_14322);
nor U14552 (N_14552,N_14344,N_14217);
nand U14553 (N_14553,N_14268,N_14211);
nand U14554 (N_14554,N_14230,N_14283);
nor U14555 (N_14555,N_14307,N_14333);
and U14556 (N_14556,N_14255,N_14328);
nor U14557 (N_14557,N_14233,N_14331);
nand U14558 (N_14558,N_14242,N_14232);
nand U14559 (N_14559,N_14234,N_14370);
or U14560 (N_14560,N_14340,N_14319);
and U14561 (N_14561,N_14269,N_14225);
nand U14562 (N_14562,N_14336,N_14342);
xor U14563 (N_14563,N_14335,N_14307);
or U14564 (N_14564,N_14375,N_14348);
nor U14565 (N_14565,N_14210,N_14214);
or U14566 (N_14566,N_14306,N_14223);
nor U14567 (N_14567,N_14338,N_14251);
and U14568 (N_14568,N_14332,N_14359);
nor U14569 (N_14569,N_14338,N_14397);
and U14570 (N_14570,N_14221,N_14280);
nor U14571 (N_14571,N_14295,N_14263);
and U14572 (N_14572,N_14207,N_14347);
nor U14573 (N_14573,N_14330,N_14317);
xor U14574 (N_14574,N_14294,N_14285);
xor U14575 (N_14575,N_14270,N_14204);
and U14576 (N_14576,N_14294,N_14217);
nand U14577 (N_14577,N_14387,N_14225);
nand U14578 (N_14578,N_14336,N_14216);
nand U14579 (N_14579,N_14265,N_14344);
and U14580 (N_14580,N_14371,N_14324);
or U14581 (N_14581,N_14315,N_14313);
nand U14582 (N_14582,N_14217,N_14279);
or U14583 (N_14583,N_14335,N_14373);
nand U14584 (N_14584,N_14352,N_14276);
nand U14585 (N_14585,N_14230,N_14201);
nor U14586 (N_14586,N_14298,N_14364);
nor U14587 (N_14587,N_14284,N_14382);
or U14588 (N_14588,N_14325,N_14205);
nor U14589 (N_14589,N_14225,N_14241);
nand U14590 (N_14590,N_14262,N_14389);
or U14591 (N_14591,N_14210,N_14292);
nand U14592 (N_14592,N_14288,N_14267);
nand U14593 (N_14593,N_14396,N_14265);
or U14594 (N_14594,N_14370,N_14355);
xnor U14595 (N_14595,N_14323,N_14372);
or U14596 (N_14596,N_14328,N_14373);
or U14597 (N_14597,N_14271,N_14307);
and U14598 (N_14598,N_14341,N_14369);
xnor U14599 (N_14599,N_14252,N_14286);
nor U14600 (N_14600,N_14515,N_14422);
nor U14601 (N_14601,N_14433,N_14500);
and U14602 (N_14602,N_14438,N_14566);
xnor U14603 (N_14603,N_14569,N_14442);
nor U14604 (N_14604,N_14448,N_14561);
nand U14605 (N_14605,N_14478,N_14494);
nor U14606 (N_14606,N_14552,N_14462);
and U14607 (N_14607,N_14446,N_14473);
and U14608 (N_14608,N_14437,N_14414);
or U14609 (N_14609,N_14579,N_14472);
and U14610 (N_14610,N_14415,N_14411);
xnor U14611 (N_14611,N_14476,N_14439);
and U14612 (N_14612,N_14556,N_14400);
nor U14613 (N_14613,N_14413,N_14487);
nor U14614 (N_14614,N_14589,N_14490);
xnor U14615 (N_14615,N_14464,N_14555);
nor U14616 (N_14616,N_14477,N_14489);
nand U14617 (N_14617,N_14538,N_14410);
and U14618 (N_14618,N_14595,N_14506);
xor U14619 (N_14619,N_14530,N_14540);
or U14620 (N_14620,N_14504,N_14513);
or U14621 (N_14621,N_14533,N_14429);
nand U14622 (N_14622,N_14403,N_14522);
nand U14623 (N_14623,N_14460,N_14417);
nand U14624 (N_14624,N_14594,N_14434);
or U14625 (N_14625,N_14416,N_14592);
nor U14626 (N_14626,N_14426,N_14586);
nor U14627 (N_14627,N_14551,N_14484);
xnor U14628 (N_14628,N_14465,N_14454);
xor U14629 (N_14629,N_14455,N_14408);
nor U14630 (N_14630,N_14529,N_14432);
nor U14631 (N_14631,N_14423,N_14488);
or U14632 (N_14632,N_14531,N_14445);
and U14633 (N_14633,N_14451,N_14583);
or U14634 (N_14634,N_14511,N_14428);
or U14635 (N_14635,N_14597,N_14449);
nand U14636 (N_14636,N_14587,N_14418);
xnor U14637 (N_14637,N_14499,N_14596);
and U14638 (N_14638,N_14577,N_14542);
nand U14639 (N_14639,N_14461,N_14516);
or U14640 (N_14640,N_14458,N_14444);
xnor U14641 (N_14641,N_14470,N_14520);
nor U14642 (N_14642,N_14525,N_14425);
nor U14643 (N_14643,N_14578,N_14450);
or U14644 (N_14644,N_14559,N_14498);
xnor U14645 (N_14645,N_14492,N_14480);
nor U14646 (N_14646,N_14493,N_14527);
or U14647 (N_14647,N_14553,N_14440);
nor U14648 (N_14648,N_14571,N_14405);
nand U14649 (N_14649,N_14547,N_14471);
and U14650 (N_14650,N_14567,N_14508);
nor U14651 (N_14651,N_14507,N_14562);
and U14652 (N_14652,N_14456,N_14526);
nor U14653 (N_14653,N_14590,N_14543);
and U14654 (N_14654,N_14580,N_14558);
xnor U14655 (N_14655,N_14512,N_14557);
or U14656 (N_14656,N_14402,N_14521);
and U14657 (N_14657,N_14554,N_14501);
nor U14658 (N_14658,N_14485,N_14560);
and U14659 (N_14659,N_14409,N_14514);
xor U14660 (N_14660,N_14441,N_14406);
nand U14661 (N_14661,N_14436,N_14435);
nand U14662 (N_14662,N_14523,N_14496);
or U14663 (N_14663,N_14565,N_14534);
or U14664 (N_14664,N_14572,N_14457);
nor U14665 (N_14665,N_14505,N_14564);
xnor U14666 (N_14666,N_14524,N_14431);
nor U14667 (N_14667,N_14474,N_14575);
and U14668 (N_14668,N_14570,N_14581);
or U14669 (N_14669,N_14412,N_14541);
nand U14670 (N_14670,N_14598,N_14585);
or U14671 (N_14671,N_14459,N_14532);
or U14672 (N_14672,N_14537,N_14549);
nand U14673 (N_14673,N_14528,N_14483);
nand U14674 (N_14674,N_14453,N_14421);
and U14675 (N_14675,N_14481,N_14519);
nor U14676 (N_14676,N_14495,N_14550);
or U14677 (N_14677,N_14486,N_14593);
xor U14678 (N_14678,N_14502,N_14536);
nand U14679 (N_14679,N_14535,N_14563);
and U14680 (N_14680,N_14419,N_14401);
and U14681 (N_14681,N_14407,N_14427);
nand U14682 (N_14682,N_14574,N_14546);
nand U14683 (N_14683,N_14568,N_14582);
or U14684 (N_14684,N_14599,N_14497);
nand U14685 (N_14685,N_14503,N_14420);
nand U14686 (N_14686,N_14517,N_14468);
and U14687 (N_14687,N_14548,N_14509);
nand U14688 (N_14688,N_14510,N_14544);
or U14689 (N_14689,N_14482,N_14518);
and U14690 (N_14690,N_14447,N_14491);
nand U14691 (N_14691,N_14443,N_14584);
or U14692 (N_14692,N_14452,N_14475);
nand U14693 (N_14693,N_14463,N_14591);
nor U14694 (N_14694,N_14466,N_14424);
nand U14695 (N_14695,N_14467,N_14404);
or U14696 (N_14696,N_14545,N_14576);
xnor U14697 (N_14697,N_14430,N_14573);
and U14698 (N_14698,N_14539,N_14479);
and U14699 (N_14699,N_14588,N_14469);
nand U14700 (N_14700,N_14429,N_14581);
or U14701 (N_14701,N_14479,N_14442);
nand U14702 (N_14702,N_14573,N_14449);
xnor U14703 (N_14703,N_14415,N_14473);
or U14704 (N_14704,N_14456,N_14546);
nor U14705 (N_14705,N_14550,N_14426);
and U14706 (N_14706,N_14511,N_14496);
and U14707 (N_14707,N_14444,N_14470);
nor U14708 (N_14708,N_14515,N_14553);
nand U14709 (N_14709,N_14528,N_14574);
and U14710 (N_14710,N_14467,N_14470);
nor U14711 (N_14711,N_14411,N_14541);
nand U14712 (N_14712,N_14436,N_14575);
nor U14713 (N_14713,N_14545,N_14476);
nor U14714 (N_14714,N_14538,N_14583);
nand U14715 (N_14715,N_14534,N_14484);
nor U14716 (N_14716,N_14519,N_14485);
nand U14717 (N_14717,N_14434,N_14538);
or U14718 (N_14718,N_14476,N_14551);
nor U14719 (N_14719,N_14458,N_14493);
or U14720 (N_14720,N_14548,N_14549);
nor U14721 (N_14721,N_14416,N_14528);
xnor U14722 (N_14722,N_14447,N_14516);
and U14723 (N_14723,N_14550,N_14434);
nand U14724 (N_14724,N_14520,N_14588);
nor U14725 (N_14725,N_14476,N_14434);
nor U14726 (N_14726,N_14551,N_14488);
or U14727 (N_14727,N_14447,N_14577);
nand U14728 (N_14728,N_14431,N_14578);
nor U14729 (N_14729,N_14430,N_14463);
nand U14730 (N_14730,N_14431,N_14466);
nor U14731 (N_14731,N_14530,N_14429);
nor U14732 (N_14732,N_14495,N_14492);
xor U14733 (N_14733,N_14565,N_14418);
or U14734 (N_14734,N_14433,N_14509);
and U14735 (N_14735,N_14439,N_14540);
xor U14736 (N_14736,N_14545,N_14439);
nor U14737 (N_14737,N_14596,N_14496);
nor U14738 (N_14738,N_14515,N_14598);
nor U14739 (N_14739,N_14497,N_14542);
and U14740 (N_14740,N_14450,N_14531);
or U14741 (N_14741,N_14558,N_14540);
nor U14742 (N_14742,N_14471,N_14568);
xnor U14743 (N_14743,N_14414,N_14534);
nor U14744 (N_14744,N_14485,N_14523);
or U14745 (N_14745,N_14572,N_14471);
and U14746 (N_14746,N_14454,N_14544);
nand U14747 (N_14747,N_14527,N_14521);
nand U14748 (N_14748,N_14491,N_14590);
or U14749 (N_14749,N_14593,N_14599);
and U14750 (N_14750,N_14582,N_14532);
xnor U14751 (N_14751,N_14490,N_14455);
xor U14752 (N_14752,N_14558,N_14506);
nor U14753 (N_14753,N_14563,N_14514);
and U14754 (N_14754,N_14404,N_14415);
or U14755 (N_14755,N_14589,N_14427);
nor U14756 (N_14756,N_14402,N_14531);
xor U14757 (N_14757,N_14520,N_14516);
nand U14758 (N_14758,N_14502,N_14434);
xor U14759 (N_14759,N_14466,N_14572);
xor U14760 (N_14760,N_14445,N_14458);
xor U14761 (N_14761,N_14480,N_14547);
nor U14762 (N_14762,N_14561,N_14593);
nor U14763 (N_14763,N_14524,N_14536);
or U14764 (N_14764,N_14483,N_14557);
nand U14765 (N_14765,N_14511,N_14414);
nand U14766 (N_14766,N_14541,N_14430);
or U14767 (N_14767,N_14420,N_14511);
nand U14768 (N_14768,N_14528,N_14565);
xor U14769 (N_14769,N_14575,N_14574);
and U14770 (N_14770,N_14567,N_14584);
and U14771 (N_14771,N_14408,N_14459);
nand U14772 (N_14772,N_14527,N_14406);
nor U14773 (N_14773,N_14416,N_14414);
or U14774 (N_14774,N_14431,N_14478);
nand U14775 (N_14775,N_14562,N_14410);
nand U14776 (N_14776,N_14458,N_14578);
xor U14777 (N_14777,N_14427,N_14488);
nand U14778 (N_14778,N_14513,N_14573);
nand U14779 (N_14779,N_14585,N_14504);
nor U14780 (N_14780,N_14530,N_14419);
nand U14781 (N_14781,N_14500,N_14405);
or U14782 (N_14782,N_14449,N_14499);
or U14783 (N_14783,N_14484,N_14488);
nand U14784 (N_14784,N_14420,N_14444);
xnor U14785 (N_14785,N_14544,N_14528);
and U14786 (N_14786,N_14432,N_14555);
or U14787 (N_14787,N_14431,N_14522);
nor U14788 (N_14788,N_14586,N_14482);
and U14789 (N_14789,N_14584,N_14458);
and U14790 (N_14790,N_14546,N_14532);
and U14791 (N_14791,N_14552,N_14590);
nand U14792 (N_14792,N_14584,N_14589);
nand U14793 (N_14793,N_14420,N_14535);
nand U14794 (N_14794,N_14578,N_14550);
and U14795 (N_14795,N_14470,N_14447);
xor U14796 (N_14796,N_14483,N_14538);
and U14797 (N_14797,N_14535,N_14404);
or U14798 (N_14798,N_14441,N_14489);
nor U14799 (N_14799,N_14443,N_14564);
and U14800 (N_14800,N_14790,N_14690);
or U14801 (N_14801,N_14776,N_14641);
or U14802 (N_14802,N_14652,N_14767);
xnor U14803 (N_14803,N_14699,N_14797);
xor U14804 (N_14804,N_14761,N_14609);
nor U14805 (N_14805,N_14734,N_14733);
or U14806 (N_14806,N_14671,N_14756);
xnor U14807 (N_14807,N_14792,N_14616);
or U14808 (N_14808,N_14646,N_14729);
nor U14809 (N_14809,N_14706,N_14694);
nand U14810 (N_14810,N_14781,N_14779);
nand U14811 (N_14811,N_14618,N_14744);
or U14812 (N_14812,N_14784,N_14657);
and U14813 (N_14813,N_14748,N_14786);
or U14814 (N_14814,N_14757,N_14770);
or U14815 (N_14815,N_14638,N_14685);
xor U14816 (N_14816,N_14649,N_14683);
nor U14817 (N_14817,N_14724,N_14725);
xor U14818 (N_14818,N_14680,N_14785);
and U14819 (N_14819,N_14686,N_14763);
or U14820 (N_14820,N_14703,N_14768);
nand U14821 (N_14821,N_14677,N_14600);
and U14822 (N_14822,N_14650,N_14629);
or U14823 (N_14823,N_14645,N_14791);
nor U14824 (N_14824,N_14793,N_14611);
nor U14825 (N_14825,N_14644,N_14764);
or U14826 (N_14826,N_14647,N_14675);
nor U14827 (N_14827,N_14721,N_14717);
or U14828 (N_14828,N_14749,N_14737);
nand U14829 (N_14829,N_14788,N_14606);
nand U14830 (N_14830,N_14613,N_14731);
and U14831 (N_14831,N_14654,N_14607);
nor U14832 (N_14832,N_14745,N_14735);
or U14833 (N_14833,N_14648,N_14777);
and U14834 (N_14834,N_14674,N_14655);
and U14835 (N_14835,N_14614,N_14743);
and U14836 (N_14836,N_14799,N_14700);
nor U14837 (N_14837,N_14665,N_14627);
or U14838 (N_14838,N_14633,N_14653);
nor U14839 (N_14839,N_14634,N_14670);
nor U14840 (N_14840,N_14796,N_14664);
nand U14841 (N_14841,N_14766,N_14662);
nor U14842 (N_14842,N_14762,N_14620);
or U14843 (N_14843,N_14693,N_14751);
xnor U14844 (N_14844,N_14626,N_14730);
or U14845 (N_14845,N_14752,N_14708);
nand U14846 (N_14846,N_14666,N_14715);
nor U14847 (N_14847,N_14719,N_14668);
nor U14848 (N_14848,N_14617,N_14798);
and U14849 (N_14849,N_14782,N_14742);
nor U14850 (N_14850,N_14714,N_14754);
or U14851 (N_14851,N_14636,N_14651);
nor U14852 (N_14852,N_14631,N_14630);
nor U14853 (N_14853,N_14625,N_14624);
xnor U14854 (N_14854,N_14772,N_14679);
xnor U14855 (N_14855,N_14780,N_14695);
or U14856 (N_14856,N_14765,N_14718);
nor U14857 (N_14857,N_14704,N_14661);
nand U14858 (N_14858,N_14682,N_14794);
nand U14859 (N_14859,N_14656,N_14740);
nor U14860 (N_14860,N_14688,N_14603);
and U14861 (N_14861,N_14672,N_14723);
and U14862 (N_14862,N_14619,N_14696);
and U14863 (N_14863,N_14632,N_14623);
and U14864 (N_14864,N_14622,N_14711);
xnor U14865 (N_14865,N_14769,N_14726);
nand U14866 (N_14866,N_14787,N_14750);
xor U14867 (N_14867,N_14771,N_14684);
nand U14868 (N_14868,N_14755,N_14722);
nand U14869 (N_14869,N_14637,N_14741);
nand U14870 (N_14870,N_14747,N_14692);
nand U14871 (N_14871,N_14669,N_14681);
nor U14872 (N_14872,N_14789,N_14659);
and U14873 (N_14873,N_14687,N_14663);
or U14874 (N_14874,N_14760,N_14736);
and U14875 (N_14875,N_14746,N_14678);
xor U14876 (N_14876,N_14732,N_14705);
xnor U14877 (N_14877,N_14709,N_14702);
nand U14878 (N_14878,N_14775,N_14605);
xnor U14879 (N_14879,N_14608,N_14712);
nor U14880 (N_14880,N_14728,N_14640);
and U14881 (N_14881,N_14689,N_14795);
nand U14882 (N_14882,N_14739,N_14643);
nor U14883 (N_14883,N_14658,N_14720);
nand U14884 (N_14884,N_14713,N_14738);
nor U14885 (N_14885,N_14783,N_14773);
nand U14886 (N_14886,N_14753,N_14710);
nor U14887 (N_14887,N_14716,N_14660);
xnor U14888 (N_14888,N_14612,N_14601);
nor U14889 (N_14889,N_14642,N_14701);
and U14890 (N_14890,N_14707,N_14621);
and U14891 (N_14891,N_14691,N_14604);
or U14892 (N_14892,N_14774,N_14610);
or U14893 (N_14893,N_14758,N_14727);
xnor U14894 (N_14894,N_14676,N_14615);
or U14895 (N_14895,N_14778,N_14602);
or U14896 (N_14896,N_14673,N_14667);
and U14897 (N_14897,N_14697,N_14759);
or U14898 (N_14898,N_14698,N_14635);
or U14899 (N_14899,N_14628,N_14639);
xnor U14900 (N_14900,N_14614,N_14656);
nand U14901 (N_14901,N_14651,N_14688);
or U14902 (N_14902,N_14644,N_14678);
or U14903 (N_14903,N_14670,N_14673);
nand U14904 (N_14904,N_14722,N_14735);
nand U14905 (N_14905,N_14684,N_14612);
nand U14906 (N_14906,N_14653,N_14708);
nand U14907 (N_14907,N_14625,N_14643);
xnor U14908 (N_14908,N_14747,N_14640);
nor U14909 (N_14909,N_14678,N_14613);
nor U14910 (N_14910,N_14791,N_14780);
nor U14911 (N_14911,N_14670,N_14707);
and U14912 (N_14912,N_14714,N_14777);
or U14913 (N_14913,N_14703,N_14728);
or U14914 (N_14914,N_14652,N_14722);
and U14915 (N_14915,N_14771,N_14652);
nand U14916 (N_14916,N_14738,N_14728);
or U14917 (N_14917,N_14640,N_14674);
nor U14918 (N_14918,N_14712,N_14785);
or U14919 (N_14919,N_14754,N_14720);
nor U14920 (N_14920,N_14779,N_14730);
nor U14921 (N_14921,N_14601,N_14770);
nor U14922 (N_14922,N_14649,N_14703);
nand U14923 (N_14923,N_14759,N_14659);
nand U14924 (N_14924,N_14779,N_14741);
xor U14925 (N_14925,N_14781,N_14623);
nor U14926 (N_14926,N_14712,N_14683);
and U14927 (N_14927,N_14626,N_14608);
nand U14928 (N_14928,N_14604,N_14678);
nand U14929 (N_14929,N_14784,N_14603);
or U14930 (N_14930,N_14662,N_14622);
xnor U14931 (N_14931,N_14603,N_14787);
nor U14932 (N_14932,N_14675,N_14733);
and U14933 (N_14933,N_14619,N_14627);
nand U14934 (N_14934,N_14788,N_14731);
and U14935 (N_14935,N_14665,N_14614);
and U14936 (N_14936,N_14626,N_14618);
or U14937 (N_14937,N_14764,N_14641);
nand U14938 (N_14938,N_14782,N_14687);
or U14939 (N_14939,N_14689,N_14799);
nor U14940 (N_14940,N_14735,N_14602);
nand U14941 (N_14941,N_14793,N_14745);
and U14942 (N_14942,N_14781,N_14709);
xnor U14943 (N_14943,N_14732,N_14690);
nand U14944 (N_14944,N_14756,N_14766);
or U14945 (N_14945,N_14644,N_14646);
nor U14946 (N_14946,N_14735,N_14719);
or U14947 (N_14947,N_14746,N_14715);
nand U14948 (N_14948,N_14733,N_14684);
nand U14949 (N_14949,N_14626,N_14797);
xnor U14950 (N_14950,N_14690,N_14752);
nor U14951 (N_14951,N_14754,N_14760);
xor U14952 (N_14952,N_14646,N_14746);
nand U14953 (N_14953,N_14621,N_14712);
nand U14954 (N_14954,N_14605,N_14609);
nand U14955 (N_14955,N_14755,N_14694);
xnor U14956 (N_14956,N_14778,N_14611);
or U14957 (N_14957,N_14771,N_14633);
and U14958 (N_14958,N_14654,N_14710);
nand U14959 (N_14959,N_14628,N_14776);
or U14960 (N_14960,N_14772,N_14666);
or U14961 (N_14961,N_14616,N_14701);
or U14962 (N_14962,N_14606,N_14621);
and U14963 (N_14963,N_14616,N_14769);
and U14964 (N_14964,N_14633,N_14708);
or U14965 (N_14965,N_14669,N_14680);
nor U14966 (N_14966,N_14618,N_14610);
or U14967 (N_14967,N_14645,N_14715);
nand U14968 (N_14968,N_14748,N_14697);
or U14969 (N_14969,N_14731,N_14774);
and U14970 (N_14970,N_14685,N_14711);
or U14971 (N_14971,N_14707,N_14795);
or U14972 (N_14972,N_14726,N_14772);
or U14973 (N_14973,N_14746,N_14698);
nor U14974 (N_14974,N_14601,N_14696);
xor U14975 (N_14975,N_14652,N_14727);
or U14976 (N_14976,N_14629,N_14720);
nand U14977 (N_14977,N_14667,N_14691);
or U14978 (N_14978,N_14738,N_14702);
and U14979 (N_14979,N_14753,N_14690);
nand U14980 (N_14980,N_14727,N_14786);
nor U14981 (N_14981,N_14790,N_14700);
nand U14982 (N_14982,N_14665,N_14699);
nor U14983 (N_14983,N_14679,N_14729);
xnor U14984 (N_14984,N_14655,N_14683);
and U14985 (N_14985,N_14639,N_14706);
nor U14986 (N_14986,N_14760,N_14612);
xnor U14987 (N_14987,N_14630,N_14650);
nor U14988 (N_14988,N_14616,N_14745);
and U14989 (N_14989,N_14796,N_14732);
nand U14990 (N_14990,N_14759,N_14708);
or U14991 (N_14991,N_14691,N_14657);
nor U14992 (N_14992,N_14771,N_14762);
and U14993 (N_14993,N_14755,N_14665);
or U14994 (N_14994,N_14625,N_14694);
nand U14995 (N_14995,N_14616,N_14704);
xnor U14996 (N_14996,N_14788,N_14792);
and U14997 (N_14997,N_14610,N_14653);
nor U14998 (N_14998,N_14628,N_14747);
nor U14999 (N_14999,N_14720,N_14686);
nor U15000 (N_15000,N_14901,N_14905);
nor U15001 (N_15001,N_14980,N_14921);
nand U15002 (N_15002,N_14947,N_14995);
or U15003 (N_15003,N_14978,N_14900);
and U15004 (N_15004,N_14969,N_14960);
and U15005 (N_15005,N_14848,N_14805);
nand U15006 (N_15006,N_14836,N_14831);
or U15007 (N_15007,N_14822,N_14890);
nand U15008 (N_15008,N_14989,N_14941);
nor U15009 (N_15009,N_14863,N_14873);
nand U15010 (N_15010,N_14895,N_14830);
or U15011 (N_15011,N_14849,N_14903);
or U15012 (N_15012,N_14883,N_14936);
or U15013 (N_15013,N_14974,N_14855);
or U15014 (N_15014,N_14837,N_14908);
and U15015 (N_15015,N_14891,N_14812);
nor U15016 (N_15016,N_14857,N_14961);
nand U15017 (N_15017,N_14818,N_14819);
or U15018 (N_15018,N_14866,N_14826);
and U15019 (N_15019,N_14840,N_14851);
or U15020 (N_15020,N_14934,N_14981);
xor U15021 (N_15021,N_14957,N_14844);
and U15022 (N_15022,N_14994,N_14897);
xor U15023 (N_15023,N_14976,N_14949);
nor U15024 (N_15024,N_14962,N_14987);
and U15025 (N_15025,N_14892,N_14861);
and U15026 (N_15026,N_14816,N_14867);
and U15027 (N_15027,N_14802,N_14821);
or U15028 (N_15028,N_14927,N_14828);
nand U15029 (N_15029,N_14925,N_14915);
nor U15030 (N_15030,N_14804,N_14999);
nor U15031 (N_15031,N_14965,N_14955);
and U15032 (N_15032,N_14884,N_14803);
or U15033 (N_15033,N_14964,N_14864);
nor U15034 (N_15034,N_14943,N_14870);
and U15035 (N_15035,N_14966,N_14834);
nand U15036 (N_15036,N_14926,N_14919);
or U15037 (N_15037,N_14889,N_14935);
nand U15038 (N_15038,N_14933,N_14833);
and U15039 (N_15039,N_14820,N_14845);
nand U15040 (N_15040,N_14944,N_14879);
or U15041 (N_15041,N_14846,N_14991);
or U15042 (N_15042,N_14854,N_14853);
nand U15043 (N_15043,N_14807,N_14917);
or U15044 (N_15044,N_14817,N_14856);
or U15045 (N_15045,N_14985,N_14885);
and U15046 (N_15046,N_14953,N_14983);
or U15047 (N_15047,N_14852,N_14898);
nor U15048 (N_15048,N_14811,N_14827);
and U15049 (N_15049,N_14971,N_14871);
xor U15050 (N_15050,N_14958,N_14909);
nor U15051 (N_15051,N_14801,N_14975);
or U15052 (N_15052,N_14832,N_14829);
or U15053 (N_15053,N_14923,N_14894);
xor U15054 (N_15054,N_14967,N_14824);
or U15055 (N_15055,N_14937,N_14938);
nor U15056 (N_15056,N_14956,N_14946);
nand U15057 (N_15057,N_14886,N_14977);
nand U15058 (N_15058,N_14841,N_14810);
xnor U15059 (N_15059,N_14951,N_14972);
nand U15060 (N_15060,N_14940,N_14992);
nor U15061 (N_15061,N_14809,N_14868);
nand U15062 (N_15062,N_14874,N_14813);
nand U15063 (N_15063,N_14916,N_14842);
nand U15064 (N_15064,N_14912,N_14948);
nand U15065 (N_15065,N_14952,N_14942);
nor U15066 (N_15066,N_14954,N_14882);
and U15067 (N_15067,N_14996,N_14998);
and U15068 (N_15068,N_14862,N_14929);
or U15069 (N_15069,N_14825,N_14939);
or U15070 (N_15070,N_14878,N_14860);
nor U15071 (N_15071,N_14865,N_14911);
or U15072 (N_15072,N_14869,N_14888);
and U15073 (N_15073,N_14922,N_14950);
nor U15074 (N_15074,N_14910,N_14843);
and U15075 (N_15075,N_14850,N_14968);
nand U15076 (N_15076,N_14924,N_14838);
xor U15077 (N_15077,N_14906,N_14872);
nor U15078 (N_15078,N_14876,N_14823);
nor U15079 (N_15079,N_14881,N_14993);
nor U15080 (N_15080,N_14918,N_14877);
nor U15081 (N_15081,N_14839,N_14880);
nor U15082 (N_15082,N_14988,N_14904);
nand U15083 (N_15083,N_14858,N_14932);
and U15084 (N_15084,N_14945,N_14913);
xnor U15085 (N_15085,N_14970,N_14899);
nand U15086 (N_15086,N_14920,N_14815);
and U15087 (N_15087,N_14896,N_14930);
or U15088 (N_15088,N_14808,N_14907);
and U15089 (N_15089,N_14806,N_14979);
nor U15090 (N_15090,N_14997,N_14835);
or U15091 (N_15091,N_14931,N_14982);
and U15092 (N_15092,N_14800,N_14914);
xnor U15093 (N_15093,N_14986,N_14902);
or U15094 (N_15094,N_14990,N_14847);
and U15095 (N_15095,N_14814,N_14984);
nand U15096 (N_15096,N_14875,N_14959);
and U15097 (N_15097,N_14893,N_14963);
or U15098 (N_15098,N_14928,N_14859);
and U15099 (N_15099,N_14887,N_14973);
nand U15100 (N_15100,N_14864,N_14997);
nor U15101 (N_15101,N_14914,N_14889);
xnor U15102 (N_15102,N_14884,N_14911);
xnor U15103 (N_15103,N_14853,N_14882);
nor U15104 (N_15104,N_14818,N_14920);
xnor U15105 (N_15105,N_14814,N_14903);
or U15106 (N_15106,N_14857,N_14987);
xor U15107 (N_15107,N_14932,N_14875);
nor U15108 (N_15108,N_14986,N_14942);
xor U15109 (N_15109,N_14898,N_14962);
and U15110 (N_15110,N_14970,N_14997);
or U15111 (N_15111,N_14970,N_14954);
and U15112 (N_15112,N_14934,N_14840);
nor U15113 (N_15113,N_14927,N_14872);
and U15114 (N_15114,N_14984,N_14865);
xnor U15115 (N_15115,N_14850,N_14878);
nand U15116 (N_15116,N_14829,N_14999);
nand U15117 (N_15117,N_14995,N_14850);
nand U15118 (N_15118,N_14802,N_14860);
or U15119 (N_15119,N_14845,N_14812);
and U15120 (N_15120,N_14974,N_14955);
and U15121 (N_15121,N_14929,N_14975);
nand U15122 (N_15122,N_14987,N_14967);
and U15123 (N_15123,N_14803,N_14956);
nor U15124 (N_15124,N_14885,N_14970);
and U15125 (N_15125,N_14888,N_14815);
nand U15126 (N_15126,N_14948,N_14837);
nor U15127 (N_15127,N_14921,N_14840);
or U15128 (N_15128,N_14906,N_14810);
nor U15129 (N_15129,N_14895,N_14960);
nand U15130 (N_15130,N_14977,N_14852);
xnor U15131 (N_15131,N_14805,N_14997);
nor U15132 (N_15132,N_14803,N_14843);
xnor U15133 (N_15133,N_14822,N_14808);
and U15134 (N_15134,N_14871,N_14932);
nand U15135 (N_15135,N_14953,N_14849);
xnor U15136 (N_15136,N_14898,N_14989);
or U15137 (N_15137,N_14821,N_14931);
nand U15138 (N_15138,N_14824,N_14946);
nand U15139 (N_15139,N_14935,N_14832);
or U15140 (N_15140,N_14965,N_14970);
or U15141 (N_15141,N_14943,N_14904);
or U15142 (N_15142,N_14968,N_14858);
and U15143 (N_15143,N_14801,N_14883);
xor U15144 (N_15144,N_14955,N_14950);
nor U15145 (N_15145,N_14977,N_14860);
xor U15146 (N_15146,N_14810,N_14981);
or U15147 (N_15147,N_14930,N_14976);
nand U15148 (N_15148,N_14960,N_14849);
and U15149 (N_15149,N_14855,N_14815);
nor U15150 (N_15150,N_14955,N_14838);
or U15151 (N_15151,N_14848,N_14896);
nand U15152 (N_15152,N_14858,N_14838);
or U15153 (N_15153,N_14916,N_14893);
or U15154 (N_15154,N_14855,N_14830);
and U15155 (N_15155,N_14969,N_14839);
nor U15156 (N_15156,N_14862,N_14932);
nor U15157 (N_15157,N_14884,N_14838);
or U15158 (N_15158,N_14814,N_14904);
or U15159 (N_15159,N_14808,N_14883);
xor U15160 (N_15160,N_14883,N_14891);
or U15161 (N_15161,N_14821,N_14908);
nand U15162 (N_15162,N_14895,N_14826);
or U15163 (N_15163,N_14864,N_14969);
nor U15164 (N_15164,N_14903,N_14996);
and U15165 (N_15165,N_14904,N_14818);
or U15166 (N_15166,N_14986,N_14927);
or U15167 (N_15167,N_14962,N_14842);
nand U15168 (N_15168,N_14920,N_14882);
or U15169 (N_15169,N_14829,N_14876);
nand U15170 (N_15170,N_14812,N_14821);
nor U15171 (N_15171,N_14866,N_14870);
or U15172 (N_15172,N_14815,N_14919);
nor U15173 (N_15173,N_14825,N_14981);
nor U15174 (N_15174,N_14968,N_14829);
nand U15175 (N_15175,N_14959,N_14930);
and U15176 (N_15176,N_14820,N_14837);
or U15177 (N_15177,N_14856,N_14833);
or U15178 (N_15178,N_14834,N_14844);
or U15179 (N_15179,N_14974,N_14810);
or U15180 (N_15180,N_14954,N_14926);
or U15181 (N_15181,N_14928,N_14920);
nand U15182 (N_15182,N_14843,N_14977);
nor U15183 (N_15183,N_14870,N_14998);
and U15184 (N_15184,N_14987,N_14926);
xor U15185 (N_15185,N_14940,N_14929);
nor U15186 (N_15186,N_14991,N_14897);
nand U15187 (N_15187,N_14998,N_14893);
or U15188 (N_15188,N_14938,N_14903);
nand U15189 (N_15189,N_14959,N_14882);
nand U15190 (N_15190,N_14949,N_14913);
nor U15191 (N_15191,N_14828,N_14966);
nand U15192 (N_15192,N_14844,N_14983);
and U15193 (N_15193,N_14852,N_14832);
nor U15194 (N_15194,N_14939,N_14833);
xor U15195 (N_15195,N_14845,N_14923);
nor U15196 (N_15196,N_14883,N_14904);
or U15197 (N_15197,N_14939,N_14818);
nor U15198 (N_15198,N_14918,N_14970);
xor U15199 (N_15199,N_14921,N_14863);
and U15200 (N_15200,N_15096,N_15039);
nand U15201 (N_15201,N_15139,N_15074);
and U15202 (N_15202,N_15052,N_15014);
nand U15203 (N_15203,N_15143,N_15149);
nor U15204 (N_15204,N_15084,N_15158);
nand U15205 (N_15205,N_15083,N_15189);
nand U15206 (N_15206,N_15077,N_15064);
or U15207 (N_15207,N_15175,N_15118);
or U15208 (N_15208,N_15188,N_15184);
and U15209 (N_15209,N_15173,N_15193);
or U15210 (N_15210,N_15162,N_15094);
and U15211 (N_15211,N_15043,N_15061);
nand U15212 (N_15212,N_15113,N_15086);
nand U15213 (N_15213,N_15031,N_15106);
or U15214 (N_15214,N_15001,N_15187);
nor U15215 (N_15215,N_15017,N_15199);
nand U15216 (N_15216,N_15057,N_15115);
or U15217 (N_15217,N_15081,N_15024);
nor U15218 (N_15218,N_15037,N_15026);
and U15219 (N_15219,N_15195,N_15132);
nand U15220 (N_15220,N_15140,N_15045);
or U15221 (N_15221,N_15123,N_15110);
nor U15222 (N_15222,N_15145,N_15073);
nand U15223 (N_15223,N_15155,N_15128);
nand U15224 (N_15224,N_15072,N_15133);
and U15225 (N_15225,N_15042,N_15079);
or U15226 (N_15226,N_15018,N_15015);
nand U15227 (N_15227,N_15034,N_15153);
nor U15228 (N_15228,N_15092,N_15154);
or U15229 (N_15229,N_15080,N_15127);
or U15230 (N_15230,N_15150,N_15138);
and U15231 (N_15231,N_15046,N_15020);
nand U15232 (N_15232,N_15055,N_15000);
nand U15233 (N_15233,N_15186,N_15002);
and U15234 (N_15234,N_15169,N_15117);
or U15235 (N_15235,N_15099,N_15035);
and U15236 (N_15236,N_15164,N_15012);
nor U15237 (N_15237,N_15011,N_15144);
or U15238 (N_15238,N_15111,N_15010);
and U15239 (N_15239,N_15168,N_15016);
xnor U15240 (N_15240,N_15059,N_15062);
nor U15241 (N_15241,N_15125,N_15041);
or U15242 (N_15242,N_15109,N_15027);
or U15243 (N_15243,N_15160,N_15167);
nand U15244 (N_15244,N_15178,N_15051);
nand U15245 (N_15245,N_15008,N_15131);
nor U15246 (N_15246,N_15048,N_15182);
nand U15247 (N_15247,N_15044,N_15134);
nand U15248 (N_15248,N_15122,N_15159);
and U15249 (N_15249,N_15068,N_15040);
or U15250 (N_15250,N_15069,N_15198);
and U15251 (N_15251,N_15013,N_15036);
nor U15252 (N_15252,N_15095,N_15075);
and U15253 (N_15253,N_15087,N_15157);
and U15254 (N_15254,N_15019,N_15126);
nand U15255 (N_15255,N_15054,N_15180);
or U15256 (N_15256,N_15033,N_15141);
nor U15257 (N_15257,N_15196,N_15176);
nand U15258 (N_15258,N_15098,N_15171);
or U15259 (N_15259,N_15091,N_15124);
nand U15260 (N_15260,N_15136,N_15119);
xor U15261 (N_15261,N_15082,N_15165);
and U15262 (N_15262,N_15063,N_15104);
or U15263 (N_15263,N_15105,N_15146);
and U15264 (N_15264,N_15148,N_15078);
and U15265 (N_15265,N_15172,N_15056);
nor U15266 (N_15266,N_15005,N_15076);
nor U15267 (N_15267,N_15006,N_15053);
nor U15268 (N_15268,N_15003,N_15114);
or U15269 (N_15269,N_15177,N_15101);
and U15270 (N_15270,N_15004,N_15120);
nand U15271 (N_15271,N_15192,N_15065);
and U15272 (N_15272,N_15121,N_15179);
nand U15273 (N_15273,N_15108,N_15107);
nor U15274 (N_15274,N_15058,N_15030);
xnor U15275 (N_15275,N_15070,N_15151);
or U15276 (N_15276,N_15089,N_15147);
and U15277 (N_15277,N_15007,N_15191);
nand U15278 (N_15278,N_15156,N_15163);
or U15279 (N_15279,N_15197,N_15112);
and U15280 (N_15280,N_15060,N_15085);
and U15281 (N_15281,N_15049,N_15050);
nand U15282 (N_15282,N_15103,N_15166);
and U15283 (N_15283,N_15032,N_15116);
xnor U15284 (N_15284,N_15161,N_15142);
or U15285 (N_15285,N_15152,N_15088);
and U15286 (N_15286,N_15067,N_15135);
xor U15287 (N_15287,N_15023,N_15100);
nor U15288 (N_15288,N_15129,N_15181);
and U15289 (N_15289,N_15130,N_15093);
or U15290 (N_15290,N_15102,N_15022);
nand U15291 (N_15291,N_15028,N_15190);
nor U15292 (N_15292,N_15029,N_15137);
nand U15293 (N_15293,N_15021,N_15170);
nor U15294 (N_15294,N_15009,N_15071);
nor U15295 (N_15295,N_15066,N_15185);
nor U15296 (N_15296,N_15047,N_15025);
nor U15297 (N_15297,N_15183,N_15174);
xnor U15298 (N_15298,N_15038,N_15097);
nor U15299 (N_15299,N_15090,N_15194);
xnor U15300 (N_15300,N_15002,N_15014);
or U15301 (N_15301,N_15193,N_15196);
nand U15302 (N_15302,N_15190,N_15122);
nand U15303 (N_15303,N_15132,N_15057);
nor U15304 (N_15304,N_15127,N_15050);
nand U15305 (N_15305,N_15095,N_15099);
nand U15306 (N_15306,N_15094,N_15116);
and U15307 (N_15307,N_15050,N_15118);
or U15308 (N_15308,N_15075,N_15179);
and U15309 (N_15309,N_15060,N_15064);
and U15310 (N_15310,N_15131,N_15179);
nand U15311 (N_15311,N_15197,N_15142);
nand U15312 (N_15312,N_15078,N_15187);
or U15313 (N_15313,N_15196,N_15184);
nand U15314 (N_15314,N_15067,N_15183);
or U15315 (N_15315,N_15123,N_15072);
nor U15316 (N_15316,N_15032,N_15107);
or U15317 (N_15317,N_15171,N_15055);
nand U15318 (N_15318,N_15085,N_15003);
nor U15319 (N_15319,N_15130,N_15145);
nor U15320 (N_15320,N_15069,N_15074);
and U15321 (N_15321,N_15175,N_15090);
nor U15322 (N_15322,N_15081,N_15048);
xor U15323 (N_15323,N_15166,N_15015);
or U15324 (N_15324,N_15190,N_15046);
or U15325 (N_15325,N_15055,N_15176);
nor U15326 (N_15326,N_15110,N_15039);
nor U15327 (N_15327,N_15166,N_15079);
or U15328 (N_15328,N_15149,N_15075);
nand U15329 (N_15329,N_15167,N_15004);
xor U15330 (N_15330,N_15053,N_15082);
nor U15331 (N_15331,N_15084,N_15003);
nor U15332 (N_15332,N_15068,N_15025);
nor U15333 (N_15333,N_15077,N_15146);
or U15334 (N_15334,N_15112,N_15150);
or U15335 (N_15335,N_15186,N_15034);
nand U15336 (N_15336,N_15117,N_15079);
or U15337 (N_15337,N_15182,N_15012);
and U15338 (N_15338,N_15113,N_15067);
nor U15339 (N_15339,N_15012,N_15103);
nand U15340 (N_15340,N_15078,N_15084);
and U15341 (N_15341,N_15175,N_15153);
nand U15342 (N_15342,N_15053,N_15009);
nand U15343 (N_15343,N_15025,N_15035);
nand U15344 (N_15344,N_15056,N_15064);
or U15345 (N_15345,N_15033,N_15172);
nor U15346 (N_15346,N_15141,N_15053);
and U15347 (N_15347,N_15134,N_15197);
nand U15348 (N_15348,N_15004,N_15176);
xnor U15349 (N_15349,N_15120,N_15033);
or U15350 (N_15350,N_15142,N_15164);
and U15351 (N_15351,N_15098,N_15114);
xor U15352 (N_15352,N_15013,N_15110);
or U15353 (N_15353,N_15194,N_15021);
or U15354 (N_15354,N_15043,N_15015);
nand U15355 (N_15355,N_15097,N_15188);
nand U15356 (N_15356,N_15010,N_15035);
or U15357 (N_15357,N_15056,N_15101);
nand U15358 (N_15358,N_15129,N_15162);
and U15359 (N_15359,N_15054,N_15028);
and U15360 (N_15360,N_15103,N_15117);
or U15361 (N_15361,N_15014,N_15151);
nor U15362 (N_15362,N_15184,N_15008);
or U15363 (N_15363,N_15131,N_15088);
nor U15364 (N_15364,N_15059,N_15036);
nor U15365 (N_15365,N_15079,N_15085);
nor U15366 (N_15366,N_15116,N_15001);
nand U15367 (N_15367,N_15143,N_15135);
nor U15368 (N_15368,N_15019,N_15139);
and U15369 (N_15369,N_15062,N_15171);
nor U15370 (N_15370,N_15062,N_15198);
nor U15371 (N_15371,N_15186,N_15052);
or U15372 (N_15372,N_15135,N_15082);
nor U15373 (N_15373,N_15027,N_15091);
or U15374 (N_15374,N_15037,N_15115);
and U15375 (N_15375,N_15156,N_15067);
nor U15376 (N_15376,N_15059,N_15131);
or U15377 (N_15377,N_15106,N_15182);
xor U15378 (N_15378,N_15095,N_15082);
or U15379 (N_15379,N_15089,N_15188);
or U15380 (N_15380,N_15078,N_15045);
nor U15381 (N_15381,N_15089,N_15154);
nor U15382 (N_15382,N_15146,N_15168);
and U15383 (N_15383,N_15155,N_15055);
and U15384 (N_15384,N_15018,N_15027);
and U15385 (N_15385,N_15037,N_15123);
nor U15386 (N_15386,N_15139,N_15183);
or U15387 (N_15387,N_15184,N_15185);
nor U15388 (N_15388,N_15093,N_15080);
and U15389 (N_15389,N_15087,N_15084);
nor U15390 (N_15390,N_15168,N_15139);
and U15391 (N_15391,N_15192,N_15198);
or U15392 (N_15392,N_15034,N_15035);
nand U15393 (N_15393,N_15161,N_15005);
nand U15394 (N_15394,N_15032,N_15127);
and U15395 (N_15395,N_15026,N_15087);
and U15396 (N_15396,N_15034,N_15051);
and U15397 (N_15397,N_15037,N_15035);
and U15398 (N_15398,N_15191,N_15088);
or U15399 (N_15399,N_15095,N_15001);
or U15400 (N_15400,N_15307,N_15243);
or U15401 (N_15401,N_15341,N_15221);
and U15402 (N_15402,N_15254,N_15263);
and U15403 (N_15403,N_15233,N_15351);
nor U15404 (N_15404,N_15244,N_15332);
nor U15405 (N_15405,N_15348,N_15210);
and U15406 (N_15406,N_15217,N_15329);
and U15407 (N_15407,N_15224,N_15379);
nor U15408 (N_15408,N_15335,N_15320);
xnor U15409 (N_15409,N_15318,N_15285);
xor U15410 (N_15410,N_15368,N_15249);
nand U15411 (N_15411,N_15384,N_15359);
and U15412 (N_15412,N_15353,N_15220);
nand U15413 (N_15413,N_15267,N_15391);
or U15414 (N_15414,N_15317,N_15240);
nor U15415 (N_15415,N_15252,N_15314);
xnor U15416 (N_15416,N_15325,N_15274);
or U15417 (N_15417,N_15346,N_15315);
or U15418 (N_15418,N_15206,N_15246);
xor U15419 (N_15419,N_15251,N_15231);
or U15420 (N_15420,N_15360,N_15275);
and U15421 (N_15421,N_15270,N_15365);
or U15422 (N_15422,N_15260,N_15343);
nand U15423 (N_15423,N_15222,N_15226);
nand U15424 (N_15424,N_15337,N_15395);
or U15425 (N_15425,N_15201,N_15227);
and U15426 (N_15426,N_15380,N_15340);
nand U15427 (N_15427,N_15291,N_15236);
and U15428 (N_15428,N_15383,N_15319);
nand U15429 (N_15429,N_15242,N_15377);
nor U15430 (N_15430,N_15216,N_15279);
and U15431 (N_15431,N_15232,N_15256);
nor U15432 (N_15432,N_15297,N_15373);
xor U15433 (N_15433,N_15396,N_15223);
nand U15434 (N_15434,N_15207,N_15278);
nand U15435 (N_15435,N_15354,N_15266);
or U15436 (N_15436,N_15304,N_15367);
or U15437 (N_15437,N_15238,N_15259);
nor U15438 (N_15438,N_15349,N_15366);
and U15439 (N_15439,N_15288,N_15241);
nor U15440 (N_15440,N_15200,N_15327);
nor U15441 (N_15441,N_15204,N_15338);
nand U15442 (N_15442,N_15281,N_15331);
and U15443 (N_15443,N_15345,N_15294);
nor U15444 (N_15444,N_15305,N_15276);
and U15445 (N_15445,N_15261,N_15203);
nand U15446 (N_15446,N_15328,N_15273);
nand U15447 (N_15447,N_15397,N_15299);
nand U15448 (N_15448,N_15312,N_15311);
nor U15449 (N_15449,N_15316,N_15393);
nand U15450 (N_15450,N_15357,N_15211);
or U15451 (N_15451,N_15292,N_15205);
xor U15452 (N_15452,N_15355,N_15235);
nand U15453 (N_15453,N_15214,N_15284);
nor U15454 (N_15454,N_15280,N_15370);
nor U15455 (N_15455,N_15209,N_15376);
or U15456 (N_15456,N_15213,N_15295);
xnor U15457 (N_15457,N_15363,N_15352);
or U15458 (N_15458,N_15392,N_15289);
or U15459 (N_15459,N_15257,N_15342);
xnor U15460 (N_15460,N_15313,N_15283);
or U15461 (N_15461,N_15301,N_15269);
xnor U15462 (N_15462,N_15290,N_15350);
nand U15463 (N_15463,N_15215,N_15208);
or U15464 (N_15464,N_15386,N_15212);
nor U15465 (N_15465,N_15218,N_15253);
nand U15466 (N_15466,N_15369,N_15394);
and U15467 (N_15467,N_15245,N_15374);
nand U15468 (N_15468,N_15323,N_15258);
and U15469 (N_15469,N_15372,N_15378);
or U15470 (N_15470,N_15262,N_15287);
or U15471 (N_15471,N_15399,N_15361);
and U15472 (N_15472,N_15296,N_15219);
nor U15473 (N_15473,N_15271,N_15326);
and U15474 (N_15474,N_15381,N_15390);
nand U15475 (N_15475,N_15333,N_15303);
and U15476 (N_15476,N_15306,N_15202);
nand U15477 (N_15477,N_15272,N_15225);
or U15478 (N_15478,N_15229,N_15334);
and U15479 (N_15479,N_15339,N_15322);
or U15480 (N_15480,N_15358,N_15298);
nor U15481 (N_15481,N_15398,N_15321);
xor U15482 (N_15482,N_15387,N_15375);
or U15483 (N_15483,N_15255,N_15308);
nor U15484 (N_15484,N_15250,N_15265);
and U15485 (N_15485,N_15268,N_15248);
nand U15486 (N_15486,N_15239,N_15282);
or U15487 (N_15487,N_15264,N_15356);
nand U15488 (N_15488,N_15302,N_15364);
nand U15489 (N_15489,N_15293,N_15389);
nand U15490 (N_15490,N_15230,N_15286);
and U15491 (N_15491,N_15237,N_15277);
or U15492 (N_15492,N_15228,N_15324);
xor U15493 (N_15493,N_15330,N_15382);
xnor U15494 (N_15494,N_15385,N_15344);
nor U15495 (N_15495,N_15347,N_15247);
nor U15496 (N_15496,N_15300,N_15362);
or U15497 (N_15497,N_15309,N_15310);
or U15498 (N_15498,N_15234,N_15336);
and U15499 (N_15499,N_15388,N_15371);
and U15500 (N_15500,N_15391,N_15317);
nand U15501 (N_15501,N_15313,N_15212);
nor U15502 (N_15502,N_15292,N_15355);
nand U15503 (N_15503,N_15208,N_15345);
nand U15504 (N_15504,N_15276,N_15374);
nand U15505 (N_15505,N_15287,N_15299);
or U15506 (N_15506,N_15367,N_15381);
nor U15507 (N_15507,N_15324,N_15302);
or U15508 (N_15508,N_15265,N_15260);
nand U15509 (N_15509,N_15337,N_15321);
nand U15510 (N_15510,N_15316,N_15219);
nor U15511 (N_15511,N_15395,N_15344);
nand U15512 (N_15512,N_15251,N_15365);
nor U15513 (N_15513,N_15326,N_15313);
and U15514 (N_15514,N_15264,N_15326);
nand U15515 (N_15515,N_15354,N_15385);
nand U15516 (N_15516,N_15296,N_15337);
and U15517 (N_15517,N_15368,N_15303);
nor U15518 (N_15518,N_15270,N_15387);
nand U15519 (N_15519,N_15387,N_15237);
or U15520 (N_15520,N_15376,N_15245);
xnor U15521 (N_15521,N_15369,N_15241);
nand U15522 (N_15522,N_15312,N_15320);
or U15523 (N_15523,N_15306,N_15291);
and U15524 (N_15524,N_15262,N_15227);
nor U15525 (N_15525,N_15375,N_15295);
nor U15526 (N_15526,N_15304,N_15384);
and U15527 (N_15527,N_15303,N_15345);
xnor U15528 (N_15528,N_15308,N_15381);
or U15529 (N_15529,N_15386,N_15232);
xnor U15530 (N_15530,N_15354,N_15289);
nor U15531 (N_15531,N_15246,N_15229);
nor U15532 (N_15532,N_15325,N_15235);
and U15533 (N_15533,N_15341,N_15291);
nand U15534 (N_15534,N_15250,N_15212);
xor U15535 (N_15535,N_15311,N_15239);
or U15536 (N_15536,N_15247,N_15315);
and U15537 (N_15537,N_15346,N_15377);
nor U15538 (N_15538,N_15313,N_15356);
xnor U15539 (N_15539,N_15383,N_15333);
nor U15540 (N_15540,N_15346,N_15303);
nand U15541 (N_15541,N_15231,N_15275);
nor U15542 (N_15542,N_15234,N_15348);
and U15543 (N_15543,N_15325,N_15352);
or U15544 (N_15544,N_15389,N_15246);
and U15545 (N_15545,N_15218,N_15318);
and U15546 (N_15546,N_15350,N_15210);
nor U15547 (N_15547,N_15288,N_15374);
or U15548 (N_15548,N_15236,N_15217);
or U15549 (N_15549,N_15214,N_15257);
and U15550 (N_15550,N_15288,N_15255);
xor U15551 (N_15551,N_15388,N_15219);
and U15552 (N_15552,N_15356,N_15306);
nand U15553 (N_15553,N_15280,N_15323);
nor U15554 (N_15554,N_15281,N_15250);
xnor U15555 (N_15555,N_15236,N_15305);
or U15556 (N_15556,N_15219,N_15257);
and U15557 (N_15557,N_15268,N_15365);
nand U15558 (N_15558,N_15308,N_15316);
or U15559 (N_15559,N_15253,N_15242);
or U15560 (N_15560,N_15227,N_15321);
and U15561 (N_15561,N_15265,N_15319);
xnor U15562 (N_15562,N_15301,N_15379);
or U15563 (N_15563,N_15338,N_15266);
nand U15564 (N_15564,N_15313,N_15289);
and U15565 (N_15565,N_15205,N_15378);
nor U15566 (N_15566,N_15364,N_15307);
nor U15567 (N_15567,N_15277,N_15296);
and U15568 (N_15568,N_15331,N_15262);
or U15569 (N_15569,N_15210,N_15305);
and U15570 (N_15570,N_15373,N_15376);
nand U15571 (N_15571,N_15298,N_15341);
or U15572 (N_15572,N_15352,N_15343);
or U15573 (N_15573,N_15271,N_15399);
nand U15574 (N_15574,N_15297,N_15242);
nor U15575 (N_15575,N_15367,N_15255);
and U15576 (N_15576,N_15241,N_15375);
or U15577 (N_15577,N_15382,N_15244);
nand U15578 (N_15578,N_15264,N_15380);
nand U15579 (N_15579,N_15200,N_15345);
and U15580 (N_15580,N_15205,N_15218);
nand U15581 (N_15581,N_15342,N_15275);
and U15582 (N_15582,N_15301,N_15349);
nand U15583 (N_15583,N_15350,N_15377);
and U15584 (N_15584,N_15218,N_15225);
or U15585 (N_15585,N_15274,N_15310);
xnor U15586 (N_15586,N_15219,N_15318);
nor U15587 (N_15587,N_15242,N_15353);
and U15588 (N_15588,N_15261,N_15210);
nand U15589 (N_15589,N_15391,N_15255);
nor U15590 (N_15590,N_15230,N_15345);
nand U15591 (N_15591,N_15263,N_15233);
or U15592 (N_15592,N_15228,N_15347);
nand U15593 (N_15593,N_15312,N_15259);
or U15594 (N_15594,N_15346,N_15229);
xnor U15595 (N_15595,N_15287,N_15355);
xor U15596 (N_15596,N_15230,N_15320);
and U15597 (N_15597,N_15211,N_15347);
or U15598 (N_15598,N_15317,N_15318);
and U15599 (N_15599,N_15206,N_15213);
or U15600 (N_15600,N_15404,N_15424);
or U15601 (N_15601,N_15403,N_15412);
nand U15602 (N_15602,N_15517,N_15579);
or U15603 (N_15603,N_15567,N_15535);
and U15604 (N_15604,N_15529,N_15481);
nand U15605 (N_15605,N_15559,N_15430);
and U15606 (N_15606,N_15452,N_15451);
nand U15607 (N_15607,N_15578,N_15561);
nand U15608 (N_15608,N_15459,N_15520);
xnor U15609 (N_15609,N_15565,N_15486);
and U15610 (N_15610,N_15401,N_15539);
nor U15611 (N_15611,N_15549,N_15457);
and U15612 (N_15612,N_15537,N_15417);
and U15613 (N_15613,N_15489,N_15555);
and U15614 (N_15614,N_15566,N_15463);
or U15615 (N_15615,N_15418,N_15583);
or U15616 (N_15616,N_15536,N_15466);
nor U15617 (N_15617,N_15521,N_15469);
and U15618 (N_15618,N_15470,N_15429);
nand U15619 (N_15619,N_15450,N_15516);
nand U15620 (N_15620,N_15446,N_15534);
nor U15621 (N_15621,N_15485,N_15473);
nand U15622 (N_15622,N_15571,N_15570);
nor U15623 (N_15623,N_15433,N_15484);
nor U15624 (N_15624,N_15453,N_15428);
nor U15625 (N_15625,N_15504,N_15542);
nand U15626 (N_15626,N_15419,N_15501);
xor U15627 (N_15627,N_15414,N_15575);
nor U15628 (N_15628,N_15465,N_15598);
or U15629 (N_15629,N_15462,N_15554);
nor U15630 (N_15630,N_15556,N_15402);
and U15631 (N_15631,N_15441,N_15595);
nor U15632 (N_15632,N_15512,N_15439);
nand U15633 (N_15633,N_15442,N_15492);
nor U15634 (N_15634,N_15478,N_15477);
and U15635 (N_15635,N_15467,N_15448);
nor U15636 (N_15636,N_15438,N_15584);
xnor U15637 (N_15637,N_15490,N_15497);
or U15638 (N_15638,N_15443,N_15527);
nor U15639 (N_15639,N_15423,N_15591);
and U15640 (N_15640,N_15416,N_15456);
or U15641 (N_15641,N_15551,N_15425);
and U15642 (N_15642,N_15586,N_15577);
and U15643 (N_15643,N_15530,N_15408);
xnor U15644 (N_15644,N_15597,N_15500);
nor U15645 (N_15645,N_15580,N_15528);
and U15646 (N_15646,N_15487,N_15547);
nor U15647 (N_15647,N_15407,N_15552);
xor U15648 (N_15648,N_15593,N_15525);
or U15649 (N_15649,N_15494,N_15434);
or U15650 (N_15650,N_15543,N_15522);
and U15651 (N_15651,N_15587,N_15531);
nor U15652 (N_15652,N_15550,N_15576);
and U15653 (N_15653,N_15532,N_15558);
xor U15654 (N_15654,N_15483,N_15572);
nand U15655 (N_15655,N_15589,N_15588);
and U15656 (N_15656,N_15475,N_15585);
nor U15657 (N_15657,N_15503,N_15491);
or U15658 (N_15658,N_15413,N_15523);
nand U15659 (N_15659,N_15410,N_15573);
and U15660 (N_15660,N_15581,N_15464);
nand U15661 (N_15661,N_15422,N_15435);
or U15662 (N_15662,N_15426,N_15474);
xor U15663 (N_15663,N_15415,N_15545);
nor U15664 (N_15664,N_15468,N_15511);
nor U15665 (N_15665,N_15508,N_15569);
nor U15666 (N_15666,N_15524,N_15436);
and U15667 (N_15667,N_15507,N_15562);
or U15668 (N_15668,N_15431,N_15406);
nor U15669 (N_15669,N_15538,N_15482);
nand U15670 (N_15670,N_15599,N_15420);
and U15671 (N_15671,N_15458,N_15460);
nand U15672 (N_15672,N_15488,N_15400);
nor U15673 (N_15673,N_15596,N_15445);
xor U15674 (N_15674,N_15582,N_15553);
or U15675 (N_15675,N_15546,N_15509);
xor U15676 (N_15676,N_15405,N_15505);
nor U15677 (N_15677,N_15495,N_15447);
and U15678 (N_15678,N_15454,N_15592);
nor U15679 (N_15679,N_15590,N_15568);
nor U15680 (N_15680,N_15506,N_15548);
and U15681 (N_15681,N_15515,N_15449);
and U15682 (N_15682,N_15437,N_15533);
nand U15683 (N_15683,N_15421,N_15574);
xor U15684 (N_15684,N_15455,N_15513);
and U15685 (N_15685,N_15498,N_15444);
nand U15686 (N_15686,N_15499,N_15480);
or U15687 (N_15687,N_15541,N_15519);
and U15688 (N_15688,N_15502,N_15476);
nor U15689 (N_15689,N_15563,N_15526);
nand U15690 (N_15690,N_15409,N_15461);
or U15691 (N_15691,N_15471,N_15440);
or U15692 (N_15692,N_15432,N_15510);
nand U15693 (N_15693,N_15496,N_15514);
and U15694 (N_15694,N_15560,N_15544);
nor U15695 (N_15695,N_15557,N_15427);
or U15696 (N_15696,N_15594,N_15540);
nand U15697 (N_15697,N_15472,N_15564);
nor U15698 (N_15698,N_15493,N_15479);
nand U15699 (N_15699,N_15411,N_15518);
or U15700 (N_15700,N_15513,N_15408);
or U15701 (N_15701,N_15513,N_15512);
nand U15702 (N_15702,N_15435,N_15542);
or U15703 (N_15703,N_15410,N_15509);
nor U15704 (N_15704,N_15457,N_15542);
or U15705 (N_15705,N_15524,N_15547);
and U15706 (N_15706,N_15559,N_15411);
and U15707 (N_15707,N_15565,N_15546);
xor U15708 (N_15708,N_15597,N_15438);
and U15709 (N_15709,N_15558,N_15448);
or U15710 (N_15710,N_15400,N_15595);
nor U15711 (N_15711,N_15492,N_15597);
or U15712 (N_15712,N_15481,N_15450);
nand U15713 (N_15713,N_15406,N_15512);
nor U15714 (N_15714,N_15576,N_15546);
nand U15715 (N_15715,N_15454,N_15538);
nand U15716 (N_15716,N_15589,N_15449);
and U15717 (N_15717,N_15560,N_15401);
or U15718 (N_15718,N_15498,N_15413);
nand U15719 (N_15719,N_15481,N_15518);
nor U15720 (N_15720,N_15469,N_15405);
and U15721 (N_15721,N_15525,N_15466);
or U15722 (N_15722,N_15498,N_15448);
nor U15723 (N_15723,N_15421,N_15551);
nand U15724 (N_15724,N_15529,N_15573);
and U15725 (N_15725,N_15567,N_15572);
nor U15726 (N_15726,N_15454,N_15556);
xor U15727 (N_15727,N_15417,N_15571);
or U15728 (N_15728,N_15462,N_15499);
nor U15729 (N_15729,N_15517,N_15498);
nand U15730 (N_15730,N_15433,N_15464);
or U15731 (N_15731,N_15419,N_15590);
nor U15732 (N_15732,N_15528,N_15563);
or U15733 (N_15733,N_15568,N_15418);
and U15734 (N_15734,N_15436,N_15494);
xnor U15735 (N_15735,N_15437,N_15407);
nor U15736 (N_15736,N_15428,N_15578);
or U15737 (N_15737,N_15573,N_15420);
and U15738 (N_15738,N_15401,N_15493);
and U15739 (N_15739,N_15508,N_15458);
and U15740 (N_15740,N_15430,N_15548);
nor U15741 (N_15741,N_15589,N_15479);
or U15742 (N_15742,N_15524,N_15580);
nand U15743 (N_15743,N_15533,N_15593);
nor U15744 (N_15744,N_15465,N_15568);
and U15745 (N_15745,N_15432,N_15545);
nand U15746 (N_15746,N_15546,N_15594);
and U15747 (N_15747,N_15414,N_15446);
and U15748 (N_15748,N_15541,N_15530);
or U15749 (N_15749,N_15419,N_15421);
or U15750 (N_15750,N_15488,N_15534);
nand U15751 (N_15751,N_15484,N_15562);
and U15752 (N_15752,N_15435,N_15403);
nand U15753 (N_15753,N_15512,N_15565);
nand U15754 (N_15754,N_15486,N_15537);
nor U15755 (N_15755,N_15513,N_15463);
or U15756 (N_15756,N_15521,N_15510);
nand U15757 (N_15757,N_15574,N_15554);
xor U15758 (N_15758,N_15564,N_15543);
nor U15759 (N_15759,N_15528,N_15526);
nor U15760 (N_15760,N_15526,N_15534);
and U15761 (N_15761,N_15481,N_15409);
xor U15762 (N_15762,N_15484,N_15535);
nor U15763 (N_15763,N_15400,N_15491);
and U15764 (N_15764,N_15489,N_15459);
or U15765 (N_15765,N_15464,N_15577);
and U15766 (N_15766,N_15544,N_15454);
and U15767 (N_15767,N_15549,N_15584);
or U15768 (N_15768,N_15495,N_15427);
and U15769 (N_15769,N_15509,N_15446);
or U15770 (N_15770,N_15455,N_15488);
and U15771 (N_15771,N_15405,N_15502);
nor U15772 (N_15772,N_15429,N_15527);
and U15773 (N_15773,N_15464,N_15585);
nand U15774 (N_15774,N_15424,N_15409);
nand U15775 (N_15775,N_15548,N_15559);
nor U15776 (N_15776,N_15597,N_15525);
nor U15777 (N_15777,N_15460,N_15566);
or U15778 (N_15778,N_15559,N_15417);
or U15779 (N_15779,N_15492,N_15550);
or U15780 (N_15780,N_15598,N_15556);
xor U15781 (N_15781,N_15404,N_15555);
and U15782 (N_15782,N_15521,N_15418);
nor U15783 (N_15783,N_15461,N_15506);
or U15784 (N_15784,N_15463,N_15591);
or U15785 (N_15785,N_15423,N_15446);
xnor U15786 (N_15786,N_15512,N_15434);
and U15787 (N_15787,N_15463,N_15503);
xnor U15788 (N_15788,N_15506,N_15539);
nor U15789 (N_15789,N_15465,N_15555);
and U15790 (N_15790,N_15567,N_15422);
and U15791 (N_15791,N_15448,N_15582);
xnor U15792 (N_15792,N_15419,N_15567);
nand U15793 (N_15793,N_15405,N_15579);
nor U15794 (N_15794,N_15416,N_15469);
nor U15795 (N_15795,N_15484,N_15587);
xor U15796 (N_15796,N_15536,N_15527);
and U15797 (N_15797,N_15549,N_15583);
nor U15798 (N_15798,N_15408,N_15542);
nand U15799 (N_15799,N_15412,N_15475);
and U15800 (N_15800,N_15673,N_15702);
or U15801 (N_15801,N_15716,N_15765);
and U15802 (N_15802,N_15679,N_15643);
nor U15803 (N_15803,N_15652,N_15737);
nand U15804 (N_15804,N_15777,N_15731);
nor U15805 (N_15805,N_15704,N_15626);
nand U15806 (N_15806,N_15680,N_15784);
nor U15807 (N_15807,N_15634,N_15734);
or U15808 (N_15808,N_15775,N_15674);
nor U15809 (N_15809,N_15705,N_15700);
or U15810 (N_15810,N_15785,N_15615);
nor U15811 (N_15811,N_15742,N_15609);
or U15812 (N_15812,N_15600,N_15712);
or U15813 (N_15813,N_15715,N_15687);
or U15814 (N_15814,N_15616,N_15793);
xnor U15815 (N_15815,N_15695,N_15624);
or U15816 (N_15816,N_15710,N_15744);
nor U15817 (N_15817,N_15662,N_15645);
nor U15818 (N_15818,N_15786,N_15781);
nand U15819 (N_15819,N_15733,N_15641);
or U15820 (N_15820,N_15678,N_15614);
nand U15821 (N_15821,N_15720,N_15648);
and U15822 (N_15822,N_15745,N_15766);
nor U15823 (N_15823,N_15633,N_15669);
nand U15824 (N_15824,N_15711,N_15795);
nand U15825 (N_15825,N_15730,N_15638);
xor U15826 (N_15826,N_15621,N_15651);
nand U15827 (N_15827,N_15664,N_15718);
or U15828 (N_15828,N_15741,N_15639);
nor U15829 (N_15829,N_15725,N_15604);
and U15830 (N_15830,N_15755,N_15617);
or U15831 (N_15831,N_15792,N_15672);
nor U15832 (N_15832,N_15686,N_15757);
or U15833 (N_15833,N_15798,N_15637);
nand U15834 (N_15834,N_15751,N_15618);
nor U15835 (N_15835,N_15722,N_15668);
nand U15836 (N_15836,N_15619,N_15789);
nor U15837 (N_15837,N_15608,N_15706);
xnor U15838 (N_15838,N_15612,N_15732);
and U15839 (N_15839,N_15675,N_15748);
xnor U15840 (N_15840,N_15727,N_15778);
nand U15841 (N_15841,N_15603,N_15723);
nor U15842 (N_15842,N_15613,N_15630);
or U15843 (N_15843,N_15691,N_15709);
nor U15844 (N_15844,N_15759,N_15655);
nor U15845 (N_15845,N_15649,N_15721);
xnor U15846 (N_15846,N_15756,N_15684);
xnor U15847 (N_15847,N_15653,N_15650);
and U15848 (N_15848,N_15625,N_15659);
nand U15849 (N_15849,N_15701,N_15694);
nor U15850 (N_15850,N_15699,N_15644);
nor U15851 (N_15851,N_15717,N_15685);
nor U15852 (N_15852,N_15677,N_15620);
and U15853 (N_15853,N_15703,N_15663);
nand U15854 (N_15854,N_15739,N_15787);
nand U15855 (N_15855,N_15768,N_15676);
and U15856 (N_15856,N_15627,N_15660);
nor U15857 (N_15857,N_15794,N_15797);
or U15858 (N_15858,N_15642,N_15769);
nand U15859 (N_15859,N_15636,N_15767);
nand U15860 (N_15860,N_15607,N_15635);
and U15861 (N_15861,N_15647,N_15796);
nor U15862 (N_15862,N_15779,N_15762);
nand U15863 (N_15863,N_15774,N_15790);
nor U15864 (N_15864,N_15714,N_15601);
nor U15865 (N_15865,N_15656,N_15747);
nand U15866 (N_15866,N_15791,N_15631);
or U15867 (N_15867,N_15692,N_15697);
or U15868 (N_15868,N_15658,N_15782);
nor U15869 (N_15869,N_15764,N_15698);
and U15870 (N_15870,N_15708,N_15772);
or U15871 (N_15871,N_15606,N_15758);
nor U15872 (N_15872,N_15760,N_15681);
and U15873 (N_15873,N_15657,N_15696);
nand U15874 (N_15874,N_15736,N_15646);
nor U15875 (N_15875,N_15735,N_15610);
nor U15876 (N_15876,N_15611,N_15750);
and U15877 (N_15877,N_15661,N_15729);
and U15878 (N_15878,N_15671,N_15761);
nor U15879 (N_15879,N_15602,N_15771);
nor U15880 (N_15880,N_15713,N_15752);
and U15881 (N_15881,N_15788,N_15773);
or U15882 (N_15882,N_15746,N_15743);
and U15883 (N_15883,N_15623,N_15605);
and U15884 (N_15884,N_15683,N_15749);
nand U15885 (N_15885,N_15740,N_15666);
or U15886 (N_15886,N_15654,N_15770);
nor U15887 (N_15887,N_15763,N_15632);
nor U15888 (N_15888,N_15665,N_15670);
and U15889 (N_15889,N_15726,N_15754);
or U15890 (N_15890,N_15707,N_15738);
or U15891 (N_15891,N_15780,N_15783);
or U15892 (N_15892,N_15719,N_15728);
or U15893 (N_15893,N_15640,N_15689);
or U15894 (N_15894,N_15682,N_15628);
nor U15895 (N_15895,N_15753,N_15693);
nand U15896 (N_15896,N_15622,N_15629);
nor U15897 (N_15897,N_15690,N_15688);
or U15898 (N_15898,N_15799,N_15667);
or U15899 (N_15899,N_15776,N_15724);
nand U15900 (N_15900,N_15673,N_15639);
nand U15901 (N_15901,N_15678,N_15671);
nor U15902 (N_15902,N_15754,N_15775);
or U15903 (N_15903,N_15653,N_15766);
nor U15904 (N_15904,N_15712,N_15651);
or U15905 (N_15905,N_15649,N_15611);
or U15906 (N_15906,N_15717,N_15602);
xnor U15907 (N_15907,N_15603,N_15638);
nor U15908 (N_15908,N_15748,N_15631);
nor U15909 (N_15909,N_15612,N_15662);
xor U15910 (N_15910,N_15724,N_15616);
nor U15911 (N_15911,N_15786,N_15648);
nand U15912 (N_15912,N_15680,N_15718);
and U15913 (N_15913,N_15686,N_15647);
nand U15914 (N_15914,N_15758,N_15783);
or U15915 (N_15915,N_15626,N_15623);
xnor U15916 (N_15916,N_15609,N_15658);
nand U15917 (N_15917,N_15635,N_15653);
and U15918 (N_15918,N_15754,N_15699);
and U15919 (N_15919,N_15650,N_15780);
and U15920 (N_15920,N_15640,N_15725);
nor U15921 (N_15921,N_15725,N_15601);
nand U15922 (N_15922,N_15789,N_15622);
and U15923 (N_15923,N_15745,N_15614);
or U15924 (N_15924,N_15729,N_15770);
nand U15925 (N_15925,N_15611,N_15629);
and U15926 (N_15926,N_15733,N_15698);
or U15927 (N_15927,N_15780,N_15773);
or U15928 (N_15928,N_15685,N_15726);
nor U15929 (N_15929,N_15685,N_15712);
nor U15930 (N_15930,N_15608,N_15623);
xor U15931 (N_15931,N_15777,N_15674);
and U15932 (N_15932,N_15696,N_15770);
or U15933 (N_15933,N_15722,N_15729);
nand U15934 (N_15934,N_15734,N_15702);
nand U15935 (N_15935,N_15616,N_15627);
and U15936 (N_15936,N_15677,N_15743);
and U15937 (N_15937,N_15764,N_15663);
or U15938 (N_15938,N_15749,N_15716);
or U15939 (N_15939,N_15742,N_15644);
nor U15940 (N_15940,N_15600,N_15770);
and U15941 (N_15941,N_15704,N_15610);
nand U15942 (N_15942,N_15625,N_15721);
nor U15943 (N_15943,N_15680,N_15770);
and U15944 (N_15944,N_15714,N_15619);
nor U15945 (N_15945,N_15639,N_15782);
and U15946 (N_15946,N_15675,N_15710);
nand U15947 (N_15947,N_15735,N_15685);
nor U15948 (N_15948,N_15639,N_15765);
and U15949 (N_15949,N_15624,N_15664);
nand U15950 (N_15950,N_15697,N_15704);
nand U15951 (N_15951,N_15784,N_15788);
and U15952 (N_15952,N_15690,N_15675);
nand U15953 (N_15953,N_15659,N_15772);
or U15954 (N_15954,N_15624,N_15660);
or U15955 (N_15955,N_15683,N_15642);
xor U15956 (N_15956,N_15604,N_15629);
nor U15957 (N_15957,N_15682,N_15676);
and U15958 (N_15958,N_15653,N_15649);
nor U15959 (N_15959,N_15737,N_15775);
nand U15960 (N_15960,N_15669,N_15768);
and U15961 (N_15961,N_15612,N_15786);
and U15962 (N_15962,N_15614,N_15642);
or U15963 (N_15963,N_15721,N_15678);
xnor U15964 (N_15964,N_15703,N_15790);
and U15965 (N_15965,N_15757,N_15631);
or U15966 (N_15966,N_15714,N_15690);
nand U15967 (N_15967,N_15791,N_15654);
or U15968 (N_15968,N_15618,N_15725);
nor U15969 (N_15969,N_15645,N_15734);
nor U15970 (N_15970,N_15619,N_15777);
nand U15971 (N_15971,N_15726,N_15715);
nor U15972 (N_15972,N_15771,N_15752);
or U15973 (N_15973,N_15724,N_15684);
and U15974 (N_15974,N_15670,N_15655);
nor U15975 (N_15975,N_15658,N_15772);
nor U15976 (N_15976,N_15762,N_15624);
or U15977 (N_15977,N_15607,N_15780);
or U15978 (N_15978,N_15763,N_15741);
nand U15979 (N_15979,N_15651,N_15681);
and U15980 (N_15980,N_15781,N_15797);
xnor U15981 (N_15981,N_15764,N_15796);
nand U15982 (N_15982,N_15647,N_15754);
or U15983 (N_15983,N_15679,N_15642);
or U15984 (N_15984,N_15631,N_15628);
nor U15985 (N_15985,N_15675,N_15684);
nand U15986 (N_15986,N_15605,N_15785);
or U15987 (N_15987,N_15714,N_15685);
nand U15988 (N_15988,N_15722,N_15614);
or U15989 (N_15989,N_15748,N_15658);
nand U15990 (N_15990,N_15743,N_15797);
or U15991 (N_15991,N_15635,N_15715);
nor U15992 (N_15992,N_15771,N_15640);
xnor U15993 (N_15993,N_15730,N_15734);
nand U15994 (N_15994,N_15759,N_15712);
nand U15995 (N_15995,N_15671,N_15762);
or U15996 (N_15996,N_15736,N_15772);
or U15997 (N_15997,N_15706,N_15670);
nor U15998 (N_15998,N_15664,N_15774);
nand U15999 (N_15999,N_15703,N_15614);
and U16000 (N_16000,N_15914,N_15921);
nor U16001 (N_16001,N_15890,N_15971);
nor U16002 (N_16002,N_15961,N_15820);
or U16003 (N_16003,N_15945,N_15982);
or U16004 (N_16004,N_15800,N_15873);
and U16005 (N_16005,N_15845,N_15954);
nor U16006 (N_16006,N_15836,N_15980);
xnor U16007 (N_16007,N_15818,N_15938);
xnor U16008 (N_16008,N_15986,N_15959);
nand U16009 (N_16009,N_15974,N_15956);
nor U16010 (N_16010,N_15856,N_15815);
nor U16011 (N_16011,N_15834,N_15801);
or U16012 (N_16012,N_15908,N_15806);
nand U16013 (N_16013,N_15893,N_15865);
or U16014 (N_16014,N_15897,N_15947);
nor U16015 (N_16015,N_15819,N_15984);
and U16016 (N_16016,N_15880,N_15891);
nand U16017 (N_16017,N_15838,N_15805);
nand U16018 (N_16018,N_15978,N_15902);
or U16019 (N_16019,N_15927,N_15944);
nor U16020 (N_16020,N_15987,N_15807);
xnor U16021 (N_16021,N_15883,N_15851);
and U16022 (N_16022,N_15831,N_15901);
nand U16023 (N_16023,N_15882,N_15861);
or U16024 (N_16024,N_15946,N_15849);
nand U16025 (N_16025,N_15922,N_15965);
or U16026 (N_16026,N_15832,N_15877);
and U16027 (N_16027,N_15903,N_15917);
or U16028 (N_16028,N_15999,N_15892);
nand U16029 (N_16029,N_15846,N_15976);
and U16030 (N_16030,N_15835,N_15934);
nand U16031 (N_16031,N_15829,N_15859);
nor U16032 (N_16032,N_15981,N_15847);
or U16033 (N_16033,N_15952,N_15989);
xor U16034 (N_16034,N_15888,N_15970);
nand U16035 (N_16035,N_15802,N_15833);
nand U16036 (N_16036,N_15853,N_15951);
nand U16037 (N_16037,N_15931,N_15920);
nand U16038 (N_16038,N_15874,N_15864);
and U16039 (N_16039,N_15860,N_15804);
nand U16040 (N_16040,N_15960,N_15948);
or U16041 (N_16041,N_15811,N_15953);
xnor U16042 (N_16042,N_15923,N_15827);
nand U16043 (N_16043,N_15906,N_15943);
or U16044 (N_16044,N_15885,N_15968);
nor U16045 (N_16045,N_15928,N_15866);
nor U16046 (N_16046,N_15949,N_15918);
or U16047 (N_16047,N_15900,N_15909);
or U16048 (N_16048,N_15935,N_15843);
and U16049 (N_16049,N_15994,N_15983);
nor U16050 (N_16050,N_15857,N_15942);
or U16051 (N_16051,N_15979,N_15871);
and U16052 (N_16052,N_15940,N_15904);
and U16053 (N_16053,N_15810,N_15887);
nand U16054 (N_16054,N_15884,N_15854);
nor U16055 (N_16055,N_15870,N_15812);
xnor U16056 (N_16056,N_15896,N_15886);
nor U16057 (N_16057,N_15957,N_15930);
nand U16058 (N_16058,N_15964,N_15958);
nand U16059 (N_16059,N_15899,N_15912);
xor U16060 (N_16060,N_15814,N_15997);
nand U16061 (N_16061,N_15841,N_15821);
and U16062 (N_16062,N_15950,N_15973);
nor U16063 (N_16063,N_15855,N_15867);
and U16064 (N_16064,N_15936,N_15941);
or U16065 (N_16065,N_15966,N_15872);
xor U16066 (N_16066,N_15842,N_15876);
nand U16067 (N_16067,N_15817,N_15910);
or U16068 (N_16068,N_15895,N_15808);
and U16069 (N_16069,N_15868,N_15816);
xor U16070 (N_16070,N_15996,N_15915);
or U16071 (N_16071,N_15911,N_15878);
or U16072 (N_16072,N_15924,N_15905);
nor U16073 (N_16073,N_15848,N_15824);
nor U16074 (N_16074,N_15939,N_15850);
nand U16075 (N_16075,N_15907,N_15916);
nand U16076 (N_16076,N_15963,N_15955);
xor U16077 (N_16077,N_15840,N_15830);
or U16078 (N_16078,N_15858,N_15919);
nand U16079 (N_16079,N_15803,N_15823);
or U16080 (N_16080,N_15975,N_15926);
xor U16081 (N_16081,N_15913,N_15969);
or U16082 (N_16082,N_15809,N_15967);
xnor U16083 (N_16083,N_15875,N_15990);
or U16084 (N_16084,N_15932,N_15929);
xnor U16085 (N_16085,N_15852,N_15937);
and U16086 (N_16086,N_15998,N_15995);
and U16087 (N_16087,N_15985,N_15863);
nor U16088 (N_16088,N_15837,N_15925);
nand U16089 (N_16089,N_15844,N_15898);
or U16090 (N_16090,N_15992,N_15991);
nor U16091 (N_16091,N_15839,N_15993);
nand U16092 (N_16092,N_15894,N_15862);
nand U16093 (N_16093,N_15879,N_15825);
and U16094 (N_16094,N_15972,N_15813);
nand U16095 (N_16095,N_15822,N_15933);
or U16096 (N_16096,N_15889,N_15988);
or U16097 (N_16097,N_15826,N_15962);
or U16098 (N_16098,N_15828,N_15869);
or U16099 (N_16099,N_15977,N_15881);
nand U16100 (N_16100,N_15848,N_15953);
nand U16101 (N_16101,N_15826,N_15948);
and U16102 (N_16102,N_15895,N_15945);
and U16103 (N_16103,N_15883,N_15970);
xnor U16104 (N_16104,N_15894,N_15858);
xnor U16105 (N_16105,N_15844,N_15818);
or U16106 (N_16106,N_15925,N_15955);
and U16107 (N_16107,N_15800,N_15826);
or U16108 (N_16108,N_15864,N_15920);
and U16109 (N_16109,N_15805,N_15825);
or U16110 (N_16110,N_15871,N_15999);
or U16111 (N_16111,N_15982,N_15882);
nor U16112 (N_16112,N_15959,N_15831);
and U16113 (N_16113,N_15984,N_15806);
nor U16114 (N_16114,N_15938,N_15913);
and U16115 (N_16115,N_15889,N_15945);
nor U16116 (N_16116,N_15854,N_15953);
nand U16117 (N_16117,N_15924,N_15875);
xnor U16118 (N_16118,N_15890,N_15891);
nor U16119 (N_16119,N_15890,N_15888);
nand U16120 (N_16120,N_15835,N_15815);
and U16121 (N_16121,N_15945,N_15802);
xnor U16122 (N_16122,N_15933,N_15878);
or U16123 (N_16123,N_15856,N_15837);
and U16124 (N_16124,N_15996,N_15892);
and U16125 (N_16125,N_15980,N_15805);
or U16126 (N_16126,N_15998,N_15941);
or U16127 (N_16127,N_15948,N_15890);
nor U16128 (N_16128,N_15895,N_15842);
or U16129 (N_16129,N_15875,N_15823);
and U16130 (N_16130,N_15878,N_15826);
xor U16131 (N_16131,N_15813,N_15840);
or U16132 (N_16132,N_15981,N_15814);
or U16133 (N_16133,N_15857,N_15841);
and U16134 (N_16134,N_15960,N_15882);
nor U16135 (N_16135,N_15890,N_15942);
nand U16136 (N_16136,N_15958,N_15954);
and U16137 (N_16137,N_15879,N_15827);
or U16138 (N_16138,N_15896,N_15980);
xnor U16139 (N_16139,N_15877,N_15880);
nand U16140 (N_16140,N_15949,N_15832);
nand U16141 (N_16141,N_15939,N_15972);
nor U16142 (N_16142,N_15883,N_15935);
or U16143 (N_16143,N_15840,N_15874);
or U16144 (N_16144,N_15845,N_15809);
xor U16145 (N_16145,N_15843,N_15947);
and U16146 (N_16146,N_15905,N_15816);
or U16147 (N_16147,N_15943,N_15842);
nor U16148 (N_16148,N_15870,N_15889);
nand U16149 (N_16149,N_15809,N_15990);
and U16150 (N_16150,N_15834,N_15920);
or U16151 (N_16151,N_15928,N_15970);
or U16152 (N_16152,N_15908,N_15990);
and U16153 (N_16153,N_15803,N_15813);
or U16154 (N_16154,N_15896,N_15813);
nor U16155 (N_16155,N_15920,N_15959);
nor U16156 (N_16156,N_15987,N_15851);
or U16157 (N_16157,N_15800,N_15940);
xnor U16158 (N_16158,N_15837,N_15801);
nand U16159 (N_16159,N_15981,N_15924);
xor U16160 (N_16160,N_15814,N_15923);
nand U16161 (N_16161,N_15866,N_15978);
nor U16162 (N_16162,N_15844,N_15886);
nor U16163 (N_16163,N_15967,N_15982);
nor U16164 (N_16164,N_15917,N_15839);
nand U16165 (N_16165,N_15865,N_15960);
or U16166 (N_16166,N_15927,N_15847);
and U16167 (N_16167,N_15988,N_15878);
and U16168 (N_16168,N_15979,N_15940);
nor U16169 (N_16169,N_15831,N_15803);
or U16170 (N_16170,N_15929,N_15879);
or U16171 (N_16171,N_15981,N_15906);
and U16172 (N_16172,N_15847,N_15809);
and U16173 (N_16173,N_15826,N_15953);
and U16174 (N_16174,N_15812,N_15926);
nor U16175 (N_16175,N_15861,N_15959);
nand U16176 (N_16176,N_15942,N_15813);
xnor U16177 (N_16177,N_15853,N_15923);
nand U16178 (N_16178,N_15959,N_15921);
and U16179 (N_16179,N_15937,N_15977);
or U16180 (N_16180,N_15952,N_15921);
and U16181 (N_16181,N_15870,N_15839);
nand U16182 (N_16182,N_15983,N_15991);
nand U16183 (N_16183,N_15896,N_15972);
nor U16184 (N_16184,N_15981,N_15800);
xor U16185 (N_16185,N_15944,N_15922);
and U16186 (N_16186,N_15821,N_15878);
nand U16187 (N_16187,N_15922,N_15979);
or U16188 (N_16188,N_15849,N_15866);
nand U16189 (N_16189,N_15820,N_15919);
nor U16190 (N_16190,N_15844,N_15879);
nor U16191 (N_16191,N_15833,N_15979);
and U16192 (N_16192,N_15895,N_15990);
xor U16193 (N_16193,N_15837,N_15850);
and U16194 (N_16194,N_15856,N_15842);
nand U16195 (N_16195,N_15925,N_15899);
or U16196 (N_16196,N_15872,N_15819);
xnor U16197 (N_16197,N_15946,N_15951);
or U16198 (N_16198,N_15936,N_15893);
and U16199 (N_16199,N_15802,N_15922);
nor U16200 (N_16200,N_16058,N_16085);
nand U16201 (N_16201,N_16067,N_16100);
nor U16202 (N_16202,N_16133,N_16170);
xnor U16203 (N_16203,N_16108,N_16126);
and U16204 (N_16204,N_16002,N_16120);
nand U16205 (N_16205,N_16029,N_16148);
and U16206 (N_16206,N_16112,N_16082);
and U16207 (N_16207,N_16071,N_16033);
or U16208 (N_16208,N_16110,N_16046);
and U16209 (N_16209,N_16090,N_16189);
nand U16210 (N_16210,N_16128,N_16124);
and U16211 (N_16211,N_16129,N_16021);
nand U16212 (N_16212,N_16177,N_16106);
xor U16213 (N_16213,N_16079,N_16020);
xnor U16214 (N_16214,N_16045,N_16178);
nor U16215 (N_16215,N_16006,N_16078);
and U16216 (N_16216,N_16003,N_16062);
or U16217 (N_16217,N_16059,N_16144);
and U16218 (N_16218,N_16016,N_16028);
nor U16219 (N_16219,N_16073,N_16012);
xor U16220 (N_16220,N_16165,N_16163);
and U16221 (N_16221,N_16168,N_16096);
and U16222 (N_16222,N_16052,N_16061);
nand U16223 (N_16223,N_16019,N_16191);
or U16224 (N_16224,N_16198,N_16042);
and U16225 (N_16225,N_16195,N_16053);
or U16226 (N_16226,N_16176,N_16169);
and U16227 (N_16227,N_16139,N_16197);
and U16228 (N_16228,N_16075,N_16065);
nor U16229 (N_16229,N_16134,N_16155);
nand U16230 (N_16230,N_16147,N_16009);
xnor U16231 (N_16231,N_16044,N_16080);
nor U16232 (N_16232,N_16086,N_16151);
or U16233 (N_16233,N_16117,N_16121);
nor U16234 (N_16234,N_16063,N_16131);
and U16235 (N_16235,N_16050,N_16187);
nor U16236 (N_16236,N_16066,N_16130);
and U16237 (N_16237,N_16141,N_16060);
nor U16238 (N_16238,N_16055,N_16092);
nand U16239 (N_16239,N_16160,N_16099);
xnor U16240 (N_16240,N_16156,N_16025);
and U16241 (N_16241,N_16011,N_16081);
xnor U16242 (N_16242,N_16109,N_16143);
nor U16243 (N_16243,N_16136,N_16014);
or U16244 (N_16244,N_16153,N_16199);
or U16245 (N_16245,N_16152,N_16119);
nor U16246 (N_16246,N_16135,N_16031);
nand U16247 (N_16247,N_16102,N_16173);
and U16248 (N_16248,N_16007,N_16041);
and U16249 (N_16249,N_16057,N_16008);
and U16250 (N_16250,N_16023,N_16172);
and U16251 (N_16251,N_16024,N_16188);
nor U16252 (N_16252,N_16076,N_16158);
and U16253 (N_16253,N_16038,N_16005);
nor U16254 (N_16254,N_16087,N_16077);
nand U16255 (N_16255,N_16159,N_16018);
nor U16256 (N_16256,N_16069,N_16157);
or U16257 (N_16257,N_16072,N_16182);
or U16258 (N_16258,N_16093,N_16037);
xor U16259 (N_16259,N_16140,N_16013);
xor U16260 (N_16260,N_16196,N_16174);
xor U16261 (N_16261,N_16035,N_16114);
or U16262 (N_16262,N_16084,N_16098);
or U16263 (N_16263,N_16132,N_16004);
nor U16264 (N_16264,N_16027,N_16032);
and U16265 (N_16265,N_16167,N_16162);
or U16266 (N_16266,N_16161,N_16125);
nor U16267 (N_16267,N_16107,N_16104);
nor U16268 (N_16268,N_16115,N_16015);
nand U16269 (N_16269,N_16094,N_16164);
xor U16270 (N_16270,N_16190,N_16175);
and U16271 (N_16271,N_16194,N_16166);
or U16272 (N_16272,N_16001,N_16034);
or U16273 (N_16273,N_16186,N_16146);
and U16274 (N_16274,N_16150,N_16192);
and U16275 (N_16275,N_16049,N_16142);
or U16276 (N_16276,N_16180,N_16123);
xnor U16277 (N_16277,N_16030,N_16101);
and U16278 (N_16278,N_16068,N_16047);
and U16279 (N_16279,N_16051,N_16026);
nand U16280 (N_16280,N_16010,N_16116);
or U16281 (N_16281,N_16056,N_16088);
xor U16282 (N_16282,N_16022,N_16105);
xor U16283 (N_16283,N_16113,N_16181);
nand U16284 (N_16284,N_16048,N_16043);
nand U16285 (N_16285,N_16103,N_16118);
nor U16286 (N_16286,N_16145,N_16000);
nand U16287 (N_16287,N_16036,N_16097);
or U16288 (N_16288,N_16017,N_16091);
and U16289 (N_16289,N_16070,N_16122);
or U16290 (N_16290,N_16095,N_16183);
and U16291 (N_16291,N_16185,N_16171);
xnor U16292 (N_16292,N_16040,N_16149);
nor U16293 (N_16293,N_16154,N_16138);
nand U16294 (N_16294,N_16074,N_16054);
and U16295 (N_16295,N_16039,N_16193);
nor U16296 (N_16296,N_16111,N_16064);
nor U16297 (N_16297,N_16137,N_16127);
xor U16298 (N_16298,N_16184,N_16179);
nand U16299 (N_16299,N_16083,N_16089);
and U16300 (N_16300,N_16043,N_16115);
and U16301 (N_16301,N_16047,N_16074);
nand U16302 (N_16302,N_16130,N_16000);
nor U16303 (N_16303,N_16053,N_16178);
nor U16304 (N_16304,N_16157,N_16173);
and U16305 (N_16305,N_16110,N_16005);
nand U16306 (N_16306,N_16153,N_16080);
or U16307 (N_16307,N_16102,N_16039);
nand U16308 (N_16308,N_16132,N_16017);
nand U16309 (N_16309,N_16174,N_16011);
nor U16310 (N_16310,N_16055,N_16022);
xnor U16311 (N_16311,N_16047,N_16034);
or U16312 (N_16312,N_16009,N_16040);
nor U16313 (N_16313,N_16016,N_16088);
xnor U16314 (N_16314,N_16112,N_16034);
nor U16315 (N_16315,N_16137,N_16173);
xor U16316 (N_16316,N_16104,N_16191);
xor U16317 (N_16317,N_16185,N_16095);
nand U16318 (N_16318,N_16017,N_16048);
nor U16319 (N_16319,N_16167,N_16125);
nor U16320 (N_16320,N_16171,N_16144);
and U16321 (N_16321,N_16191,N_16140);
xor U16322 (N_16322,N_16164,N_16144);
and U16323 (N_16323,N_16053,N_16166);
nand U16324 (N_16324,N_16050,N_16022);
xor U16325 (N_16325,N_16052,N_16175);
nor U16326 (N_16326,N_16129,N_16143);
nand U16327 (N_16327,N_16195,N_16083);
or U16328 (N_16328,N_16180,N_16163);
nor U16329 (N_16329,N_16170,N_16011);
and U16330 (N_16330,N_16113,N_16075);
nor U16331 (N_16331,N_16063,N_16108);
and U16332 (N_16332,N_16193,N_16000);
and U16333 (N_16333,N_16043,N_16075);
nor U16334 (N_16334,N_16138,N_16123);
nand U16335 (N_16335,N_16149,N_16147);
nand U16336 (N_16336,N_16018,N_16111);
and U16337 (N_16337,N_16037,N_16169);
nor U16338 (N_16338,N_16135,N_16015);
nand U16339 (N_16339,N_16054,N_16124);
and U16340 (N_16340,N_16163,N_16074);
nand U16341 (N_16341,N_16090,N_16017);
and U16342 (N_16342,N_16114,N_16127);
and U16343 (N_16343,N_16152,N_16184);
xor U16344 (N_16344,N_16110,N_16018);
nand U16345 (N_16345,N_16028,N_16138);
nand U16346 (N_16346,N_16094,N_16179);
and U16347 (N_16347,N_16094,N_16101);
and U16348 (N_16348,N_16188,N_16043);
nor U16349 (N_16349,N_16183,N_16015);
nand U16350 (N_16350,N_16002,N_16152);
and U16351 (N_16351,N_16150,N_16072);
xor U16352 (N_16352,N_16064,N_16159);
and U16353 (N_16353,N_16102,N_16072);
and U16354 (N_16354,N_16045,N_16098);
or U16355 (N_16355,N_16066,N_16197);
nand U16356 (N_16356,N_16072,N_16011);
nor U16357 (N_16357,N_16034,N_16186);
nor U16358 (N_16358,N_16015,N_16129);
nand U16359 (N_16359,N_16096,N_16123);
nand U16360 (N_16360,N_16014,N_16016);
and U16361 (N_16361,N_16129,N_16008);
and U16362 (N_16362,N_16180,N_16105);
and U16363 (N_16363,N_16124,N_16156);
nand U16364 (N_16364,N_16096,N_16191);
or U16365 (N_16365,N_16059,N_16033);
and U16366 (N_16366,N_16067,N_16133);
nand U16367 (N_16367,N_16152,N_16040);
and U16368 (N_16368,N_16003,N_16058);
and U16369 (N_16369,N_16059,N_16096);
nand U16370 (N_16370,N_16146,N_16195);
and U16371 (N_16371,N_16072,N_16197);
or U16372 (N_16372,N_16031,N_16023);
nand U16373 (N_16373,N_16028,N_16145);
nor U16374 (N_16374,N_16125,N_16179);
nand U16375 (N_16375,N_16144,N_16044);
nand U16376 (N_16376,N_16174,N_16009);
and U16377 (N_16377,N_16048,N_16180);
nand U16378 (N_16378,N_16054,N_16154);
nand U16379 (N_16379,N_16149,N_16065);
and U16380 (N_16380,N_16041,N_16015);
and U16381 (N_16381,N_16097,N_16096);
and U16382 (N_16382,N_16137,N_16035);
nand U16383 (N_16383,N_16197,N_16112);
nor U16384 (N_16384,N_16005,N_16194);
nand U16385 (N_16385,N_16048,N_16137);
or U16386 (N_16386,N_16126,N_16100);
or U16387 (N_16387,N_16020,N_16064);
or U16388 (N_16388,N_16073,N_16100);
nor U16389 (N_16389,N_16173,N_16139);
and U16390 (N_16390,N_16167,N_16092);
nor U16391 (N_16391,N_16176,N_16044);
nand U16392 (N_16392,N_16026,N_16165);
nand U16393 (N_16393,N_16121,N_16164);
nand U16394 (N_16394,N_16009,N_16171);
or U16395 (N_16395,N_16030,N_16102);
xnor U16396 (N_16396,N_16083,N_16076);
nand U16397 (N_16397,N_16113,N_16180);
nand U16398 (N_16398,N_16167,N_16094);
nor U16399 (N_16399,N_16183,N_16121);
xnor U16400 (N_16400,N_16233,N_16227);
and U16401 (N_16401,N_16237,N_16224);
or U16402 (N_16402,N_16250,N_16301);
or U16403 (N_16403,N_16295,N_16275);
and U16404 (N_16404,N_16302,N_16273);
nor U16405 (N_16405,N_16395,N_16365);
nand U16406 (N_16406,N_16288,N_16311);
nor U16407 (N_16407,N_16231,N_16202);
nor U16408 (N_16408,N_16292,N_16289);
nor U16409 (N_16409,N_16286,N_16267);
nor U16410 (N_16410,N_16304,N_16228);
nor U16411 (N_16411,N_16307,N_16278);
nor U16412 (N_16412,N_16217,N_16334);
nor U16413 (N_16413,N_16211,N_16371);
nor U16414 (N_16414,N_16240,N_16283);
nand U16415 (N_16415,N_16399,N_16306);
or U16416 (N_16416,N_16346,N_16372);
nor U16417 (N_16417,N_16298,N_16331);
nand U16418 (N_16418,N_16374,N_16271);
nand U16419 (N_16419,N_16387,N_16248);
xnor U16420 (N_16420,N_16252,N_16245);
nor U16421 (N_16421,N_16251,N_16310);
nand U16422 (N_16422,N_16335,N_16386);
and U16423 (N_16423,N_16380,N_16356);
and U16424 (N_16424,N_16259,N_16316);
nand U16425 (N_16425,N_16327,N_16276);
nand U16426 (N_16426,N_16363,N_16325);
or U16427 (N_16427,N_16370,N_16270);
and U16428 (N_16428,N_16249,N_16254);
and U16429 (N_16429,N_16234,N_16214);
and U16430 (N_16430,N_16367,N_16393);
and U16431 (N_16431,N_16236,N_16253);
nor U16432 (N_16432,N_16205,N_16364);
and U16433 (N_16433,N_16209,N_16391);
and U16434 (N_16434,N_16353,N_16392);
nor U16435 (N_16435,N_16222,N_16305);
nand U16436 (N_16436,N_16394,N_16284);
or U16437 (N_16437,N_16351,N_16225);
nor U16438 (N_16438,N_16243,N_16297);
nor U16439 (N_16439,N_16357,N_16200);
nor U16440 (N_16440,N_16282,N_16376);
nor U16441 (N_16441,N_16294,N_16382);
and U16442 (N_16442,N_16352,N_16373);
nand U16443 (N_16443,N_16384,N_16232);
xor U16444 (N_16444,N_16242,N_16342);
and U16445 (N_16445,N_16355,N_16397);
or U16446 (N_16446,N_16338,N_16258);
or U16447 (N_16447,N_16223,N_16314);
and U16448 (N_16448,N_16287,N_16207);
and U16449 (N_16449,N_16322,N_16318);
or U16450 (N_16450,N_16337,N_16390);
nand U16451 (N_16451,N_16345,N_16215);
or U16452 (N_16452,N_16326,N_16208);
or U16453 (N_16453,N_16350,N_16218);
or U16454 (N_16454,N_16235,N_16272);
nor U16455 (N_16455,N_16246,N_16379);
nand U16456 (N_16456,N_16377,N_16319);
or U16457 (N_16457,N_16320,N_16241);
xnor U16458 (N_16458,N_16280,N_16383);
nor U16459 (N_16459,N_16290,N_16348);
nand U16460 (N_16460,N_16256,N_16255);
and U16461 (N_16461,N_16339,N_16216);
nor U16462 (N_16462,N_16329,N_16277);
and U16463 (N_16463,N_16291,N_16213);
xnor U16464 (N_16464,N_16369,N_16308);
or U16465 (N_16465,N_16201,N_16389);
and U16466 (N_16466,N_16347,N_16260);
or U16467 (N_16467,N_16323,N_16203);
and U16468 (N_16468,N_16332,N_16210);
and U16469 (N_16469,N_16300,N_16349);
and U16470 (N_16470,N_16381,N_16341);
and U16471 (N_16471,N_16362,N_16375);
and U16472 (N_16472,N_16366,N_16343);
xnor U16473 (N_16473,N_16378,N_16279);
nand U16474 (N_16474,N_16396,N_16354);
nor U16475 (N_16475,N_16206,N_16340);
or U16476 (N_16476,N_16360,N_16281);
nor U16477 (N_16477,N_16219,N_16293);
or U16478 (N_16478,N_16303,N_16230);
and U16479 (N_16479,N_16388,N_16262);
and U16480 (N_16480,N_16361,N_16238);
or U16481 (N_16481,N_16330,N_16296);
or U16482 (N_16482,N_16221,N_16321);
nand U16483 (N_16483,N_16368,N_16344);
and U16484 (N_16484,N_16285,N_16269);
nand U16485 (N_16485,N_16274,N_16315);
xor U16486 (N_16486,N_16358,N_16328);
nand U16487 (N_16487,N_16204,N_16261);
nor U16488 (N_16488,N_16264,N_16244);
nand U16489 (N_16489,N_16257,N_16398);
and U16490 (N_16490,N_16309,N_16359);
or U16491 (N_16491,N_16212,N_16324);
nand U16492 (N_16492,N_16312,N_16336);
nand U16493 (N_16493,N_16385,N_16263);
nor U16494 (N_16494,N_16313,N_16265);
nand U16495 (N_16495,N_16226,N_16229);
nand U16496 (N_16496,N_16317,N_16220);
and U16497 (N_16497,N_16247,N_16333);
nand U16498 (N_16498,N_16266,N_16299);
nand U16499 (N_16499,N_16239,N_16268);
and U16500 (N_16500,N_16252,N_16224);
nand U16501 (N_16501,N_16267,N_16391);
nor U16502 (N_16502,N_16233,N_16275);
xnor U16503 (N_16503,N_16320,N_16377);
or U16504 (N_16504,N_16303,N_16355);
nand U16505 (N_16505,N_16220,N_16372);
nand U16506 (N_16506,N_16328,N_16352);
or U16507 (N_16507,N_16336,N_16325);
or U16508 (N_16508,N_16299,N_16291);
or U16509 (N_16509,N_16266,N_16322);
nand U16510 (N_16510,N_16204,N_16398);
nor U16511 (N_16511,N_16201,N_16235);
and U16512 (N_16512,N_16225,N_16339);
nand U16513 (N_16513,N_16311,N_16322);
xor U16514 (N_16514,N_16223,N_16390);
nor U16515 (N_16515,N_16259,N_16219);
or U16516 (N_16516,N_16258,N_16399);
nand U16517 (N_16517,N_16293,N_16356);
nor U16518 (N_16518,N_16263,N_16215);
or U16519 (N_16519,N_16210,N_16215);
xor U16520 (N_16520,N_16323,N_16353);
xnor U16521 (N_16521,N_16317,N_16263);
nor U16522 (N_16522,N_16219,N_16362);
xor U16523 (N_16523,N_16365,N_16204);
and U16524 (N_16524,N_16221,N_16289);
nor U16525 (N_16525,N_16284,N_16313);
or U16526 (N_16526,N_16226,N_16340);
nand U16527 (N_16527,N_16338,N_16355);
nand U16528 (N_16528,N_16361,N_16306);
and U16529 (N_16529,N_16314,N_16309);
or U16530 (N_16530,N_16287,N_16259);
nor U16531 (N_16531,N_16335,N_16354);
nand U16532 (N_16532,N_16397,N_16316);
or U16533 (N_16533,N_16394,N_16255);
nand U16534 (N_16534,N_16236,N_16373);
nor U16535 (N_16535,N_16244,N_16276);
or U16536 (N_16536,N_16213,N_16313);
nand U16537 (N_16537,N_16345,N_16315);
xnor U16538 (N_16538,N_16395,N_16318);
or U16539 (N_16539,N_16307,N_16242);
and U16540 (N_16540,N_16342,N_16363);
nand U16541 (N_16541,N_16395,N_16234);
and U16542 (N_16542,N_16221,N_16367);
and U16543 (N_16543,N_16358,N_16291);
xor U16544 (N_16544,N_16385,N_16296);
nand U16545 (N_16545,N_16266,N_16341);
or U16546 (N_16546,N_16294,N_16217);
nor U16547 (N_16547,N_16308,N_16305);
or U16548 (N_16548,N_16307,N_16265);
or U16549 (N_16549,N_16321,N_16210);
and U16550 (N_16550,N_16358,N_16242);
or U16551 (N_16551,N_16293,N_16303);
and U16552 (N_16552,N_16334,N_16312);
nand U16553 (N_16553,N_16349,N_16291);
nor U16554 (N_16554,N_16331,N_16215);
and U16555 (N_16555,N_16267,N_16389);
xnor U16556 (N_16556,N_16372,N_16232);
nor U16557 (N_16557,N_16241,N_16202);
and U16558 (N_16558,N_16342,N_16243);
nand U16559 (N_16559,N_16228,N_16245);
nor U16560 (N_16560,N_16355,N_16239);
nor U16561 (N_16561,N_16370,N_16383);
nor U16562 (N_16562,N_16286,N_16325);
and U16563 (N_16563,N_16382,N_16380);
or U16564 (N_16564,N_16292,N_16206);
xor U16565 (N_16565,N_16275,N_16247);
nor U16566 (N_16566,N_16201,N_16257);
nor U16567 (N_16567,N_16314,N_16352);
xor U16568 (N_16568,N_16200,N_16337);
or U16569 (N_16569,N_16229,N_16379);
and U16570 (N_16570,N_16348,N_16279);
or U16571 (N_16571,N_16232,N_16281);
and U16572 (N_16572,N_16240,N_16334);
nand U16573 (N_16573,N_16238,N_16336);
or U16574 (N_16574,N_16326,N_16230);
nor U16575 (N_16575,N_16310,N_16301);
nor U16576 (N_16576,N_16320,N_16270);
nand U16577 (N_16577,N_16292,N_16316);
nand U16578 (N_16578,N_16294,N_16359);
or U16579 (N_16579,N_16320,N_16238);
or U16580 (N_16580,N_16390,N_16302);
nor U16581 (N_16581,N_16234,N_16202);
or U16582 (N_16582,N_16343,N_16378);
and U16583 (N_16583,N_16347,N_16258);
xnor U16584 (N_16584,N_16350,N_16389);
nand U16585 (N_16585,N_16315,N_16260);
nor U16586 (N_16586,N_16245,N_16336);
nand U16587 (N_16587,N_16363,N_16353);
nor U16588 (N_16588,N_16367,N_16322);
or U16589 (N_16589,N_16363,N_16233);
or U16590 (N_16590,N_16266,N_16380);
nor U16591 (N_16591,N_16324,N_16227);
or U16592 (N_16592,N_16322,N_16220);
nand U16593 (N_16593,N_16242,N_16356);
or U16594 (N_16594,N_16241,N_16380);
nand U16595 (N_16595,N_16233,N_16218);
or U16596 (N_16596,N_16226,N_16387);
nand U16597 (N_16597,N_16285,N_16315);
nand U16598 (N_16598,N_16226,N_16372);
xnor U16599 (N_16599,N_16347,N_16308);
nand U16600 (N_16600,N_16533,N_16498);
or U16601 (N_16601,N_16512,N_16542);
xor U16602 (N_16602,N_16444,N_16461);
nor U16603 (N_16603,N_16523,N_16529);
and U16604 (N_16604,N_16435,N_16459);
and U16605 (N_16605,N_16552,N_16580);
or U16606 (N_16606,N_16474,N_16460);
nand U16607 (N_16607,N_16518,N_16536);
nor U16608 (N_16608,N_16489,N_16543);
nor U16609 (N_16609,N_16526,N_16451);
and U16610 (N_16610,N_16475,N_16525);
nor U16611 (N_16611,N_16584,N_16559);
nand U16612 (N_16612,N_16456,N_16470);
or U16613 (N_16613,N_16414,N_16484);
and U16614 (N_16614,N_16480,N_16483);
and U16615 (N_16615,N_16415,N_16482);
or U16616 (N_16616,N_16585,N_16572);
nand U16617 (N_16617,N_16551,N_16588);
nor U16618 (N_16618,N_16406,N_16411);
nor U16619 (N_16619,N_16567,N_16453);
nand U16620 (N_16620,N_16424,N_16516);
nor U16621 (N_16621,N_16554,N_16563);
or U16622 (N_16622,N_16566,N_16520);
nand U16623 (N_16623,N_16544,N_16519);
nand U16624 (N_16624,N_16446,N_16582);
nand U16625 (N_16625,N_16509,N_16468);
nor U16626 (N_16626,N_16447,N_16499);
nor U16627 (N_16627,N_16471,N_16502);
nor U16628 (N_16628,N_16402,N_16558);
and U16629 (N_16629,N_16570,N_16467);
xor U16630 (N_16630,N_16524,N_16493);
nand U16631 (N_16631,N_16591,N_16488);
and U16632 (N_16632,N_16527,N_16535);
nand U16633 (N_16633,N_16575,N_16448);
nor U16634 (N_16634,N_16481,N_16500);
nand U16635 (N_16635,N_16515,N_16439);
and U16636 (N_16636,N_16497,N_16574);
and U16637 (N_16637,N_16442,N_16553);
or U16638 (N_16638,N_16419,N_16571);
or U16639 (N_16639,N_16573,N_16568);
and U16640 (N_16640,N_16503,N_16597);
nand U16641 (N_16641,N_16589,N_16583);
and U16642 (N_16642,N_16487,N_16540);
xnor U16643 (N_16643,N_16430,N_16586);
nand U16644 (N_16644,N_16429,N_16464);
nor U16645 (N_16645,N_16562,N_16569);
nor U16646 (N_16646,N_16593,N_16491);
nand U16647 (N_16647,N_16445,N_16521);
and U16648 (N_16648,N_16532,N_16441);
nand U16649 (N_16649,N_16428,N_16437);
or U16650 (N_16650,N_16530,N_16443);
nor U16651 (N_16651,N_16420,N_16560);
and U16652 (N_16652,N_16413,N_16449);
and U16653 (N_16653,N_16465,N_16549);
or U16654 (N_16654,N_16455,N_16517);
nand U16655 (N_16655,N_16462,N_16440);
nand U16656 (N_16656,N_16561,N_16513);
nor U16657 (N_16657,N_16466,N_16564);
xor U16658 (N_16658,N_16458,N_16408);
and U16659 (N_16659,N_16417,N_16452);
nor U16660 (N_16660,N_16478,N_16557);
and U16661 (N_16661,N_16514,N_16412);
and U16662 (N_16662,N_16565,N_16454);
nor U16663 (N_16663,N_16506,N_16538);
nor U16664 (N_16664,N_16409,N_16416);
nor U16665 (N_16665,N_16598,N_16422);
and U16666 (N_16666,N_16463,N_16587);
nor U16667 (N_16667,N_16594,N_16404);
or U16668 (N_16668,N_16528,N_16403);
nor U16669 (N_16669,N_16431,N_16457);
nor U16670 (N_16670,N_16400,N_16541);
and U16671 (N_16671,N_16418,N_16473);
nand U16672 (N_16672,N_16578,N_16596);
nand U16673 (N_16673,N_16423,N_16494);
nand U16674 (N_16674,N_16485,N_16505);
and U16675 (N_16675,N_16496,N_16599);
and U16676 (N_16676,N_16592,N_16511);
nand U16677 (N_16677,N_16546,N_16410);
nor U16678 (N_16678,N_16433,N_16405);
and U16679 (N_16679,N_16577,N_16534);
and U16680 (N_16680,N_16545,N_16479);
nor U16681 (N_16681,N_16595,N_16432);
or U16682 (N_16682,N_16436,N_16426);
and U16683 (N_16683,N_16504,N_16507);
nor U16684 (N_16684,N_16450,N_16486);
nor U16685 (N_16685,N_16537,N_16581);
nor U16686 (N_16686,N_16427,N_16510);
nand U16687 (N_16687,N_16477,N_16539);
nand U16688 (N_16688,N_16548,N_16547);
and U16689 (N_16689,N_16531,N_16522);
xor U16690 (N_16690,N_16472,N_16434);
and U16691 (N_16691,N_16425,N_16421);
nor U16692 (N_16692,N_16492,N_16469);
nor U16693 (N_16693,N_16579,N_16401);
and U16694 (N_16694,N_16407,N_16550);
nor U16695 (N_16695,N_16555,N_16556);
and U16696 (N_16696,N_16438,N_16476);
or U16697 (N_16697,N_16495,N_16590);
nand U16698 (N_16698,N_16490,N_16576);
nand U16699 (N_16699,N_16508,N_16501);
nor U16700 (N_16700,N_16510,N_16563);
nand U16701 (N_16701,N_16528,N_16559);
nand U16702 (N_16702,N_16409,N_16467);
nand U16703 (N_16703,N_16567,N_16467);
or U16704 (N_16704,N_16480,N_16517);
or U16705 (N_16705,N_16563,N_16505);
and U16706 (N_16706,N_16573,N_16536);
or U16707 (N_16707,N_16567,N_16578);
nand U16708 (N_16708,N_16492,N_16414);
and U16709 (N_16709,N_16514,N_16510);
nor U16710 (N_16710,N_16517,N_16599);
nor U16711 (N_16711,N_16425,N_16595);
and U16712 (N_16712,N_16598,N_16585);
nand U16713 (N_16713,N_16553,N_16569);
nor U16714 (N_16714,N_16450,N_16550);
nor U16715 (N_16715,N_16575,N_16455);
and U16716 (N_16716,N_16509,N_16402);
and U16717 (N_16717,N_16562,N_16572);
nand U16718 (N_16718,N_16435,N_16472);
xnor U16719 (N_16719,N_16438,N_16515);
or U16720 (N_16720,N_16443,N_16400);
xor U16721 (N_16721,N_16461,N_16544);
and U16722 (N_16722,N_16546,N_16536);
nor U16723 (N_16723,N_16567,N_16533);
nand U16724 (N_16724,N_16530,N_16576);
nor U16725 (N_16725,N_16478,N_16400);
or U16726 (N_16726,N_16509,N_16594);
nor U16727 (N_16727,N_16435,N_16451);
and U16728 (N_16728,N_16575,N_16535);
and U16729 (N_16729,N_16589,N_16559);
nand U16730 (N_16730,N_16576,N_16404);
xor U16731 (N_16731,N_16581,N_16469);
or U16732 (N_16732,N_16534,N_16579);
nor U16733 (N_16733,N_16478,N_16447);
or U16734 (N_16734,N_16413,N_16410);
nor U16735 (N_16735,N_16595,N_16423);
or U16736 (N_16736,N_16540,N_16542);
nor U16737 (N_16737,N_16428,N_16522);
and U16738 (N_16738,N_16567,N_16458);
or U16739 (N_16739,N_16597,N_16525);
nor U16740 (N_16740,N_16449,N_16441);
nor U16741 (N_16741,N_16595,N_16403);
and U16742 (N_16742,N_16592,N_16417);
nand U16743 (N_16743,N_16531,N_16582);
nor U16744 (N_16744,N_16581,N_16408);
xor U16745 (N_16745,N_16589,N_16468);
nor U16746 (N_16746,N_16441,N_16454);
nor U16747 (N_16747,N_16511,N_16482);
nand U16748 (N_16748,N_16554,N_16582);
and U16749 (N_16749,N_16572,N_16413);
and U16750 (N_16750,N_16468,N_16533);
nand U16751 (N_16751,N_16551,N_16581);
nor U16752 (N_16752,N_16469,N_16571);
or U16753 (N_16753,N_16511,N_16538);
and U16754 (N_16754,N_16532,N_16576);
or U16755 (N_16755,N_16527,N_16472);
or U16756 (N_16756,N_16403,N_16565);
and U16757 (N_16757,N_16465,N_16447);
or U16758 (N_16758,N_16587,N_16431);
nand U16759 (N_16759,N_16514,N_16416);
nand U16760 (N_16760,N_16509,N_16410);
and U16761 (N_16761,N_16426,N_16462);
or U16762 (N_16762,N_16409,N_16495);
and U16763 (N_16763,N_16576,N_16518);
nand U16764 (N_16764,N_16525,N_16584);
and U16765 (N_16765,N_16567,N_16444);
nand U16766 (N_16766,N_16472,N_16440);
and U16767 (N_16767,N_16534,N_16573);
nor U16768 (N_16768,N_16586,N_16573);
and U16769 (N_16769,N_16467,N_16416);
xnor U16770 (N_16770,N_16444,N_16494);
and U16771 (N_16771,N_16531,N_16552);
nor U16772 (N_16772,N_16563,N_16502);
or U16773 (N_16773,N_16514,N_16481);
nor U16774 (N_16774,N_16559,N_16440);
or U16775 (N_16775,N_16418,N_16484);
and U16776 (N_16776,N_16447,N_16488);
and U16777 (N_16777,N_16477,N_16425);
and U16778 (N_16778,N_16464,N_16523);
nor U16779 (N_16779,N_16411,N_16423);
nand U16780 (N_16780,N_16579,N_16406);
and U16781 (N_16781,N_16505,N_16559);
nor U16782 (N_16782,N_16438,N_16449);
or U16783 (N_16783,N_16464,N_16442);
nand U16784 (N_16784,N_16491,N_16521);
xor U16785 (N_16785,N_16571,N_16513);
and U16786 (N_16786,N_16567,N_16569);
nand U16787 (N_16787,N_16538,N_16421);
nand U16788 (N_16788,N_16434,N_16512);
and U16789 (N_16789,N_16598,N_16492);
nor U16790 (N_16790,N_16527,N_16548);
nand U16791 (N_16791,N_16475,N_16498);
or U16792 (N_16792,N_16546,N_16525);
or U16793 (N_16793,N_16541,N_16510);
or U16794 (N_16794,N_16533,N_16505);
xnor U16795 (N_16795,N_16479,N_16558);
nor U16796 (N_16796,N_16599,N_16498);
nor U16797 (N_16797,N_16433,N_16554);
and U16798 (N_16798,N_16488,N_16530);
or U16799 (N_16799,N_16598,N_16515);
nand U16800 (N_16800,N_16709,N_16697);
nand U16801 (N_16801,N_16795,N_16673);
or U16802 (N_16802,N_16603,N_16718);
and U16803 (N_16803,N_16734,N_16632);
nor U16804 (N_16804,N_16616,N_16679);
and U16805 (N_16805,N_16685,N_16725);
nand U16806 (N_16806,N_16783,N_16644);
or U16807 (N_16807,N_16778,N_16676);
and U16808 (N_16808,N_16637,N_16657);
nand U16809 (N_16809,N_16704,N_16664);
xnor U16810 (N_16810,N_16689,N_16640);
nor U16811 (N_16811,N_16730,N_16601);
nand U16812 (N_16812,N_16729,N_16669);
or U16813 (N_16813,N_16757,N_16792);
xor U16814 (N_16814,N_16680,N_16740);
nand U16815 (N_16815,N_16624,N_16706);
nor U16816 (N_16816,N_16708,N_16762);
and U16817 (N_16817,N_16641,N_16798);
nand U16818 (N_16818,N_16776,N_16712);
nand U16819 (N_16819,N_16658,N_16723);
nor U16820 (N_16820,N_16643,N_16797);
nor U16821 (N_16821,N_16671,N_16750);
nand U16822 (N_16822,N_16639,N_16745);
and U16823 (N_16823,N_16736,N_16630);
nand U16824 (N_16824,N_16784,N_16781);
nor U16825 (N_16825,N_16695,N_16646);
nand U16826 (N_16826,N_16608,N_16693);
nand U16827 (N_16827,N_16678,N_16774);
and U16828 (N_16828,N_16636,N_16765);
and U16829 (N_16829,N_16661,N_16620);
or U16830 (N_16830,N_16694,N_16621);
or U16831 (N_16831,N_16748,N_16605);
or U16832 (N_16832,N_16721,N_16717);
and U16833 (N_16833,N_16699,N_16701);
and U16834 (N_16834,N_16780,N_16794);
nor U16835 (N_16835,N_16789,N_16787);
nand U16836 (N_16836,N_16623,N_16618);
and U16837 (N_16837,N_16724,N_16663);
and U16838 (N_16838,N_16650,N_16666);
and U16839 (N_16839,N_16647,N_16681);
nor U16840 (N_16840,N_16754,N_16758);
or U16841 (N_16841,N_16600,N_16775);
and U16842 (N_16842,N_16649,N_16660);
or U16843 (N_16843,N_16767,N_16611);
and U16844 (N_16844,N_16614,N_16799);
or U16845 (N_16845,N_16607,N_16751);
and U16846 (N_16846,N_16627,N_16788);
nor U16847 (N_16847,N_16672,N_16634);
nand U16848 (N_16848,N_16759,N_16642);
and U16849 (N_16849,N_16733,N_16629);
nor U16850 (N_16850,N_16763,N_16756);
nor U16851 (N_16851,N_16737,N_16662);
nand U16852 (N_16852,N_16675,N_16656);
or U16853 (N_16853,N_16692,N_16744);
nand U16854 (N_16854,N_16791,N_16622);
and U16855 (N_16855,N_16728,N_16638);
xnor U16856 (N_16856,N_16682,N_16705);
nor U16857 (N_16857,N_16700,N_16796);
or U16858 (N_16858,N_16654,N_16764);
nor U16859 (N_16859,N_16604,N_16711);
or U16860 (N_16860,N_16619,N_16667);
and U16861 (N_16861,N_16698,N_16768);
nor U16862 (N_16862,N_16777,N_16766);
and U16863 (N_16863,N_16739,N_16779);
nand U16864 (N_16864,N_16720,N_16782);
nor U16865 (N_16865,N_16793,N_16686);
or U16866 (N_16866,N_16746,N_16617);
nand U16867 (N_16867,N_16732,N_16635);
or U16868 (N_16868,N_16665,N_16670);
xor U16869 (N_16869,N_16772,N_16677);
or U16870 (N_16870,N_16684,N_16726);
nor U16871 (N_16871,N_16731,N_16610);
nor U16872 (N_16872,N_16687,N_16702);
nand U16873 (N_16873,N_16633,N_16719);
nand U16874 (N_16874,N_16659,N_16714);
nand U16875 (N_16875,N_16786,N_16749);
and U16876 (N_16876,N_16753,N_16738);
and U16877 (N_16877,N_16747,N_16688);
or U16878 (N_16878,N_16715,N_16674);
nor U16879 (N_16879,N_16651,N_16771);
nand U16880 (N_16880,N_16668,N_16655);
and U16881 (N_16881,N_16683,N_16628);
nor U16882 (N_16882,N_16790,N_16769);
or U16883 (N_16883,N_16752,N_16707);
or U16884 (N_16884,N_16743,N_16722);
and U16885 (N_16885,N_16609,N_16652);
or U16886 (N_16886,N_16613,N_16653);
nand U16887 (N_16887,N_16773,N_16648);
nand U16888 (N_16888,N_16625,N_16626);
and U16889 (N_16889,N_16710,N_16761);
or U16890 (N_16890,N_16785,N_16735);
and U16891 (N_16891,N_16612,N_16631);
or U16892 (N_16892,N_16645,N_16727);
and U16893 (N_16893,N_16696,N_16760);
nor U16894 (N_16894,N_16742,N_16691);
nor U16895 (N_16895,N_16690,N_16755);
and U16896 (N_16896,N_16602,N_16703);
nand U16897 (N_16897,N_16615,N_16770);
nand U16898 (N_16898,N_16741,N_16606);
nand U16899 (N_16899,N_16716,N_16713);
and U16900 (N_16900,N_16630,N_16761);
nand U16901 (N_16901,N_16700,N_16759);
nand U16902 (N_16902,N_16670,N_16727);
or U16903 (N_16903,N_16602,N_16742);
nor U16904 (N_16904,N_16794,N_16667);
and U16905 (N_16905,N_16768,N_16790);
nor U16906 (N_16906,N_16608,N_16781);
nor U16907 (N_16907,N_16672,N_16725);
nand U16908 (N_16908,N_16641,N_16647);
nand U16909 (N_16909,N_16773,N_16671);
or U16910 (N_16910,N_16667,N_16651);
nand U16911 (N_16911,N_16755,N_16766);
and U16912 (N_16912,N_16647,N_16613);
nor U16913 (N_16913,N_16677,N_16670);
nand U16914 (N_16914,N_16696,N_16655);
and U16915 (N_16915,N_16698,N_16790);
or U16916 (N_16916,N_16611,N_16710);
nor U16917 (N_16917,N_16656,N_16623);
or U16918 (N_16918,N_16634,N_16605);
xnor U16919 (N_16919,N_16722,N_16721);
or U16920 (N_16920,N_16757,N_16691);
and U16921 (N_16921,N_16653,N_16666);
nand U16922 (N_16922,N_16657,N_16698);
nor U16923 (N_16923,N_16645,N_16696);
and U16924 (N_16924,N_16628,N_16739);
or U16925 (N_16925,N_16655,N_16699);
nand U16926 (N_16926,N_16655,N_16743);
xor U16927 (N_16927,N_16674,N_16642);
nor U16928 (N_16928,N_16626,N_16706);
or U16929 (N_16929,N_16735,N_16700);
nor U16930 (N_16930,N_16704,N_16737);
xnor U16931 (N_16931,N_16600,N_16644);
and U16932 (N_16932,N_16718,N_16674);
xnor U16933 (N_16933,N_16701,N_16771);
and U16934 (N_16934,N_16762,N_16774);
nand U16935 (N_16935,N_16704,N_16643);
nor U16936 (N_16936,N_16675,N_16664);
nand U16937 (N_16937,N_16796,N_16706);
xor U16938 (N_16938,N_16766,N_16706);
and U16939 (N_16939,N_16757,N_16798);
and U16940 (N_16940,N_16656,N_16784);
nor U16941 (N_16941,N_16770,N_16681);
xnor U16942 (N_16942,N_16661,N_16622);
or U16943 (N_16943,N_16759,N_16751);
or U16944 (N_16944,N_16644,N_16623);
and U16945 (N_16945,N_16767,N_16614);
and U16946 (N_16946,N_16721,N_16745);
and U16947 (N_16947,N_16740,N_16634);
xor U16948 (N_16948,N_16630,N_16624);
or U16949 (N_16949,N_16749,N_16615);
nor U16950 (N_16950,N_16614,N_16685);
nand U16951 (N_16951,N_16639,N_16784);
or U16952 (N_16952,N_16601,N_16643);
nor U16953 (N_16953,N_16776,N_16647);
and U16954 (N_16954,N_16797,N_16733);
or U16955 (N_16955,N_16720,N_16643);
xor U16956 (N_16956,N_16757,N_16711);
and U16957 (N_16957,N_16767,N_16707);
nand U16958 (N_16958,N_16638,N_16631);
xnor U16959 (N_16959,N_16628,N_16624);
nor U16960 (N_16960,N_16635,N_16626);
nor U16961 (N_16961,N_16618,N_16775);
and U16962 (N_16962,N_16660,N_16633);
nor U16963 (N_16963,N_16619,N_16643);
or U16964 (N_16964,N_16646,N_16758);
or U16965 (N_16965,N_16774,N_16798);
or U16966 (N_16966,N_16612,N_16748);
nand U16967 (N_16967,N_16773,N_16758);
nor U16968 (N_16968,N_16793,N_16734);
nand U16969 (N_16969,N_16689,N_16798);
nand U16970 (N_16970,N_16795,N_16612);
nand U16971 (N_16971,N_16763,N_16658);
nand U16972 (N_16972,N_16751,N_16772);
or U16973 (N_16973,N_16645,N_16678);
nand U16974 (N_16974,N_16743,N_16663);
or U16975 (N_16975,N_16724,N_16792);
nor U16976 (N_16976,N_16698,N_16666);
and U16977 (N_16977,N_16634,N_16783);
and U16978 (N_16978,N_16693,N_16688);
nor U16979 (N_16979,N_16773,N_16700);
xnor U16980 (N_16980,N_16764,N_16782);
and U16981 (N_16981,N_16691,N_16760);
or U16982 (N_16982,N_16702,N_16607);
nand U16983 (N_16983,N_16770,N_16614);
or U16984 (N_16984,N_16714,N_16614);
and U16985 (N_16985,N_16612,N_16738);
and U16986 (N_16986,N_16715,N_16621);
nand U16987 (N_16987,N_16628,N_16648);
nor U16988 (N_16988,N_16738,N_16684);
and U16989 (N_16989,N_16778,N_16737);
nand U16990 (N_16990,N_16799,N_16781);
or U16991 (N_16991,N_16691,N_16616);
or U16992 (N_16992,N_16773,N_16705);
nor U16993 (N_16993,N_16666,N_16671);
xor U16994 (N_16994,N_16727,N_16687);
or U16995 (N_16995,N_16784,N_16687);
nor U16996 (N_16996,N_16772,N_16735);
nand U16997 (N_16997,N_16695,N_16652);
and U16998 (N_16998,N_16629,N_16796);
and U16999 (N_16999,N_16632,N_16775);
or U17000 (N_17000,N_16869,N_16852);
and U17001 (N_17001,N_16901,N_16992);
nor U17002 (N_17002,N_16823,N_16844);
nor U17003 (N_17003,N_16906,N_16803);
nor U17004 (N_17004,N_16978,N_16867);
nand U17005 (N_17005,N_16843,N_16878);
nand U17006 (N_17006,N_16857,N_16879);
and U17007 (N_17007,N_16947,N_16824);
nand U17008 (N_17008,N_16806,N_16991);
and U17009 (N_17009,N_16973,N_16986);
nor U17010 (N_17010,N_16854,N_16802);
and U17011 (N_17011,N_16961,N_16940);
or U17012 (N_17012,N_16839,N_16800);
or U17013 (N_17013,N_16866,N_16811);
nor U17014 (N_17014,N_16821,N_16903);
and U17015 (N_17015,N_16909,N_16872);
xnor U17016 (N_17016,N_16972,N_16850);
nand U17017 (N_17017,N_16997,N_16838);
and U17018 (N_17018,N_16842,N_16905);
or U17019 (N_17019,N_16894,N_16976);
nor U17020 (N_17020,N_16952,N_16890);
nand U17021 (N_17021,N_16900,N_16941);
nand U17022 (N_17022,N_16907,N_16829);
and U17023 (N_17023,N_16846,N_16954);
nand U17024 (N_17024,N_16871,N_16882);
nand U17025 (N_17025,N_16913,N_16848);
or U17026 (N_17026,N_16939,N_16831);
nand U17027 (N_17027,N_16902,N_16981);
nand U17028 (N_17028,N_16977,N_16998);
nand U17029 (N_17029,N_16928,N_16861);
and U17030 (N_17030,N_16926,N_16810);
or U17031 (N_17031,N_16856,N_16818);
or U17032 (N_17032,N_16830,N_16817);
nand U17033 (N_17033,N_16891,N_16924);
nand U17034 (N_17034,N_16820,N_16963);
or U17035 (N_17035,N_16971,N_16889);
nand U17036 (N_17036,N_16970,N_16937);
nand U17037 (N_17037,N_16922,N_16950);
nor U17038 (N_17038,N_16925,N_16859);
or U17039 (N_17039,N_16892,N_16904);
and U17040 (N_17040,N_16923,N_16917);
nor U17041 (N_17041,N_16960,N_16876);
nand U17042 (N_17042,N_16833,N_16989);
and U17043 (N_17043,N_16959,N_16916);
nor U17044 (N_17044,N_16858,N_16893);
nand U17045 (N_17045,N_16968,N_16828);
and U17046 (N_17046,N_16919,N_16807);
and U17047 (N_17047,N_16938,N_16915);
nor U17048 (N_17048,N_16816,N_16956);
xnor U17049 (N_17049,N_16966,N_16975);
nand U17050 (N_17050,N_16870,N_16841);
nor U17051 (N_17051,N_16808,N_16942);
or U17052 (N_17052,N_16930,N_16863);
xnor U17053 (N_17053,N_16851,N_16877);
nor U17054 (N_17054,N_16955,N_16865);
and U17055 (N_17055,N_16908,N_16827);
or U17056 (N_17056,N_16862,N_16885);
nor U17057 (N_17057,N_16929,N_16994);
or U17058 (N_17058,N_16813,N_16805);
xor U17059 (N_17059,N_16983,N_16837);
nor U17060 (N_17060,N_16801,N_16962);
and U17061 (N_17061,N_16819,N_16809);
or U17062 (N_17062,N_16855,N_16815);
nand U17063 (N_17063,N_16883,N_16935);
nand U17064 (N_17064,N_16884,N_16965);
or U17065 (N_17065,N_16953,N_16980);
nand U17066 (N_17066,N_16931,N_16918);
and U17067 (N_17067,N_16927,N_16990);
and U17068 (N_17068,N_16969,N_16881);
nor U17069 (N_17069,N_16967,N_16860);
nand U17070 (N_17070,N_16934,N_16920);
xnor U17071 (N_17071,N_16853,N_16995);
or U17072 (N_17072,N_16957,N_16825);
or U17073 (N_17073,N_16873,N_16958);
nand U17074 (N_17074,N_16979,N_16945);
or U17075 (N_17075,N_16993,N_16868);
xor U17076 (N_17076,N_16982,N_16949);
or U17077 (N_17077,N_16880,N_16912);
or U17078 (N_17078,N_16921,N_16875);
xnor U17079 (N_17079,N_16840,N_16984);
nor U17080 (N_17080,N_16910,N_16914);
nand U17081 (N_17081,N_16899,N_16826);
xor U17082 (N_17082,N_16936,N_16886);
nand U17083 (N_17083,N_16887,N_16898);
nand U17084 (N_17084,N_16987,N_16835);
and U17085 (N_17085,N_16822,N_16874);
nor U17086 (N_17086,N_16951,N_16832);
and U17087 (N_17087,N_16847,N_16845);
nand U17088 (N_17088,N_16864,N_16946);
nand U17089 (N_17089,N_16964,N_16812);
nand U17090 (N_17090,N_16944,N_16834);
nand U17091 (N_17091,N_16897,N_16836);
xor U17092 (N_17092,N_16999,N_16804);
and U17093 (N_17093,N_16933,N_16948);
or U17094 (N_17094,N_16985,N_16911);
or U17095 (N_17095,N_16888,N_16988);
nor U17096 (N_17096,N_16849,N_16896);
or U17097 (N_17097,N_16932,N_16895);
xnor U17098 (N_17098,N_16974,N_16814);
and U17099 (N_17099,N_16943,N_16996);
or U17100 (N_17100,N_16862,N_16977);
and U17101 (N_17101,N_16860,N_16861);
and U17102 (N_17102,N_16972,N_16912);
and U17103 (N_17103,N_16905,N_16961);
or U17104 (N_17104,N_16931,N_16946);
and U17105 (N_17105,N_16974,N_16944);
or U17106 (N_17106,N_16858,N_16806);
nand U17107 (N_17107,N_16985,N_16958);
or U17108 (N_17108,N_16905,N_16838);
nand U17109 (N_17109,N_16929,N_16919);
nor U17110 (N_17110,N_16988,N_16995);
or U17111 (N_17111,N_16957,N_16991);
or U17112 (N_17112,N_16801,N_16887);
and U17113 (N_17113,N_16894,N_16911);
nand U17114 (N_17114,N_16957,N_16992);
or U17115 (N_17115,N_16848,N_16862);
nor U17116 (N_17116,N_16993,N_16926);
or U17117 (N_17117,N_16914,N_16974);
nand U17118 (N_17118,N_16928,N_16966);
nand U17119 (N_17119,N_16872,N_16845);
or U17120 (N_17120,N_16931,N_16834);
nand U17121 (N_17121,N_16916,N_16999);
nand U17122 (N_17122,N_16954,N_16973);
nor U17123 (N_17123,N_16848,N_16921);
nor U17124 (N_17124,N_16804,N_16896);
nand U17125 (N_17125,N_16955,N_16800);
and U17126 (N_17126,N_16866,N_16878);
and U17127 (N_17127,N_16881,N_16996);
and U17128 (N_17128,N_16931,N_16887);
nand U17129 (N_17129,N_16886,N_16891);
nor U17130 (N_17130,N_16855,N_16980);
or U17131 (N_17131,N_16873,N_16934);
or U17132 (N_17132,N_16824,N_16820);
and U17133 (N_17133,N_16920,N_16808);
or U17134 (N_17134,N_16868,N_16830);
nand U17135 (N_17135,N_16845,N_16927);
nor U17136 (N_17136,N_16806,N_16925);
nor U17137 (N_17137,N_16804,N_16855);
nand U17138 (N_17138,N_16922,N_16992);
xor U17139 (N_17139,N_16887,N_16864);
and U17140 (N_17140,N_16830,N_16986);
nor U17141 (N_17141,N_16966,N_16912);
nor U17142 (N_17142,N_16995,N_16868);
nand U17143 (N_17143,N_16862,N_16891);
and U17144 (N_17144,N_16832,N_16836);
or U17145 (N_17145,N_16803,N_16944);
xor U17146 (N_17146,N_16981,N_16986);
and U17147 (N_17147,N_16893,N_16826);
and U17148 (N_17148,N_16977,N_16971);
or U17149 (N_17149,N_16804,N_16911);
nor U17150 (N_17150,N_16959,N_16814);
nor U17151 (N_17151,N_16917,N_16826);
nand U17152 (N_17152,N_16988,N_16871);
nand U17153 (N_17153,N_16823,N_16946);
or U17154 (N_17154,N_16934,N_16981);
nor U17155 (N_17155,N_16984,N_16846);
nor U17156 (N_17156,N_16963,N_16961);
xnor U17157 (N_17157,N_16823,N_16832);
nor U17158 (N_17158,N_16903,N_16969);
nor U17159 (N_17159,N_16962,N_16863);
or U17160 (N_17160,N_16967,N_16844);
nand U17161 (N_17161,N_16956,N_16867);
or U17162 (N_17162,N_16973,N_16931);
or U17163 (N_17163,N_16985,N_16824);
nand U17164 (N_17164,N_16938,N_16833);
xnor U17165 (N_17165,N_16963,N_16852);
or U17166 (N_17166,N_16889,N_16818);
and U17167 (N_17167,N_16949,N_16952);
nor U17168 (N_17168,N_16864,N_16858);
nand U17169 (N_17169,N_16872,N_16989);
or U17170 (N_17170,N_16854,N_16850);
nor U17171 (N_17171,N_16909,N_16838);
or U17172 (N_17172,N_16878,N_16905);
and U17173 (N_17173,N_16900,N_16859);
nor U17174 (N_17174,N_16814,N_16847);
and U17175 (N_17175,N_16862,N_16849);
and U17176 (N_17176,N_16983,N_16936);
and U17177 (N_17177,N_16883,N_16865);
and U17178 (N_17178,N_16812,N_16954);
xor U17179 (N_17179,N_16854,N_16868);
or U17180 (N_17180,N_16826,N_16986);
nor U17181 (N_17181,N_16960,N_16840);
nor U17182 (N_17182,N_16868,N_16855);
nand U17183 (N_17183,N_16834,N_16970);
and U17184 (N_17184,N_16806,N_16867);
or U17185 (N_17185,N_16897,N_16829);
or U17186 (N_17186,N_16931,N_16890);
nor U17187 (N_17187,N_16922,N_16897);
nor U17188 (N_17188,N_16994,N_16950);
nand U17189 (N_17189,N_16944,N_16816);
nor U17190 (N_17190,N_16918,N_16876);
or U17191 (N_17191,N_16976,N_16942);
and U17192 (N_17192,N_16984,N_16894);
and U17193 (N_17193,N_16981,N_16800);
and U17194 (N_17194,N_16971,N_16914);
and U17195 (N_17195,N_16968,N_16836);
or U17196 (N_17196,N_16993,N_16974);
or U17197 (N_17197,N_16986,N_16909);
nor U17198 (N_17198,N_16805,N_16871);
nor U17199 (N_17199,N_16875,N_16837);
nor U17200 (N_17200,N_17159,N_17181);
nor U17201 (N_17201,N_17024,N_17080);
and U17202 (N_17202,N_17016,N_17138);
and U17203 (N_17203,N_17120,N_17006);
or U17204 (N_17204,N_17044,N_17009);
or U17205 (N_17205,N_17091,N_17147);
nand U17206 (N_17206,N_17099,N_17022);
nand U17207 (N_17207,N_17032,N_17037);
and U17208 (N_17208,N_17008,N_17130);
or U17209 (N_17209,N_17155,N_17160);
nand U17210 (N_17210,N_17199,N_17167);
nor U17211 (N_17211,N_17154,N_17190);
nor U17212 (N_17212,N_17100,N_17088);
xnor U17213 (N_17213,N_17136,N_17051);
nand U17214 (N_17214,N_17057,N_17065);
or U17215 (N_17215,N_17173,N_17021);
and U17216 (N_17216,N_17036,N_17072);
or U17217 (N_17217,N_17098,N_17046);
and U17218 (N_17218,N_17105,N_17083);
nand U17219 (N_17219,N_17101,N_17188);
nor U17220 (N_17220,N_17000,N_17162);
and U17221 (N_17221,N_17178,N_17187);
or U17222 (N_17222,N_17102,N_17047);
and U17223 (N_17223,N_17125,N_17183);
nand U17224 (N_17224,N_17020,N_17074);
nor U17225 (N_17225,N_17127,N_17109);
nand U17226 (N_17226,N_17180,N_17082);
or U17227 (N_17227,N_17118,N_17104);
nor U17228 (N_17228,N_17132,N_17084);
and U17229 (N_17229,N_17025,N_17066);
nand U17230 (N_17230,N_17157,N_17040);
nor U17231 (N_17231,N_17002,N_17124);
or U17232 (N_17232,N_17061,N_17087);
nand U17233 (N_17233,N_17049,N_17067);
nor U17234 (N_17234,N_17174,N_17054);
or U17235 (N_17235,N_17145,N_17135);
nor U17236 (N_17236,N_17185,N_17112);
or U17237 (N_17237,N_17045,N_17129);
xnor U17238 (N_17238,N_17001,N_17107);
or U17239 (N_17239,N_17148,N_17184);
xor U17240 (N_17240,N_17171,N_17122);
nand U17241 (N_17241,N_17013,N_17041);
xor U17242 (N_17242,N_17175,N_17086);
nor U17243 (N_17243,N_17166,N_17075);
and U17244 (N_17244,N_17177,N_17149);
and U17245 (N_17245,N_17151,N_17034);
nand U17246 (N_17246,N_17038,N_17003);
nand U17247 (N_17247,N_17073,N_17058);
or U17248 (N_17248,N_17062,N_17126);
nor U17249 (N_17249,N_17197,N_17134);
or U17250 (N_17250,N_17131,N_17095);
nor U17251 (N_17251,N_17156,N_17123);
nand U17252 (N_17252,N_17163,N_17059);
nand U17253 (N_17253,N_17055,N_17169);
and U17254 (N_17254,N_17053,N_17116);
and U17255 (N_17255,N_17064,N_17179);
nor U17256 (N_17256,N_17143,N_17023);
nand U17257 (N_17257,N_17121,N_17192);
nor U17258 (N_17258,N_17033,N_17027);
and U17259 (N_17259,N_17015,N_17128);
or U17260 (N_17260,N_17165,N_17077);
and U17261 (N_17261,N_17005,N_17096);
xor U17262 (N_17262,N_17007,N_17018);
or U17263 (N_17263,N_17078,N_17141);
nand U17264 (N_17264,N_17110,N_17170);
nand U17265 (N_17265,N_17029,N_17052);
nor U17266 (N_17266,N_17079,N_17195);
or U17267 (N_17267,N_17164,N_17133);
nand U17268 (N_17268,N_17014,N_17150);
and U17269 (N_17269,N_17193,N_17106);
and U17270 (N_17270,N_17012,N_17198);
and U17271 (N_17271,N_17069,N_17168);
and U17272 (N_17272,N_17030,N_17146);
nor U17273 (N_17273,N_17070,N_17043);
or U17274 (N_17274,N_17186,N_17011);
or U17275 (N_17275,N_17042,N_17111);
or U17276 (N_17276,N_17142,N_17103);
nand U17277 (N_17277,N_17172,N_17035);
nor U17278 (N_17278,N_17076,N_17056);
nand U17279 (N_17279,N_17139,N_17089);
and U17280 (N_17280,N_17140,N_17119);
and U17281 (N_17281,N_17039,N_17182);
nand U17282 (N_17282,N_17152,N_17010);
nor U17283 (N_17283,N_17094,N_17063);
xnor U17284 (N_17284,N_17144,N_17093);
or U17285 (N_17285,N_17097,N_17153);
nand U17286 (N_17286,N_17114,N_17137);
nor U17287 (N_17287,N_17068,N_17090);
nor U17288 (N_17288,N_17117,N_17189);
and U17289 (N_17289,N_17004,N_17194);
or U17290 (N_17290,N_17050,N_17017);
xnor U17291 (N_17291,N_17161,N_17026);
nor U17292 (N_17292,N_17081,N_17158);
and U17293 (N_17293,N_17060,N_17092);
or U17294 (N_17294,N_17019,N_17031);
or U17295 (N_17295,N_17191,N_17115);
xnor U17296 (N_17296,N_17048,N_17028);
and U17297 (N_17297,N_17108,N_17071);
xor U17298 (N_17298,N_17085,N_17176);
or U17299 (N_17299,N_17113,N_17196);
or U17300 (N_17300,N_17083,N_17082);
and U17301 (N_17301,N_17168,N_17182);
nand U17302 (N_17302,N_17126,N_17185);
xnor U17303 (N_17303,N_17030,N_17114);
xnor U17304 (N_17304,N_17060,N_17083);
and U17305 (N_17305,N_17021,N_17199);
or U17306 (N_17306,N_17136,N_17002);
nor U17307 (N_17307,N_17058,N_17169);
nor U17308 (N_17308,N_17184,N_17059);
or U17309 (N_17309,N_17118,N_17092);
and U17310 (N_17310,N_17188,N_17074);
or U17311 (N_17311,N_17134,N_17065);
nor U17312 (N_17312,N_17095,N_17065);
and U17313 (N_17313,N_17188,N_17134);
nor U17314 (N_17314,N_17006,N_17032);
and U17315 (N_17315,N_17106,N_17115);
xor U17316 (N_17316,N_17047,N_17040);
and U17317 (N_17317,N_17083,N_17137);
nand U17318 (N_17318,N_17134,N_17163);
and U17319 (N_17319,N_17193,N_17135);
and U17320 (N_17320,N_17059,N_17107);
xor U17321 (N_17321,N_17146,N_17005);
nand U17322 (N_17322,N_17178,N_17026);
and U17323 (N_17323,N_17019,N_17149);
and U17324 (N_17324,N_17119,N_17115);
or U17325 (N_17325,N_17003,N_17067);
and U17326 (N_17326,N_17031,N_17122);
nor U17327 (N_17327,N_17149,N_17133);
nand U17328 (N_17328,N_17175,N_17139);
xnor U17329 (N_17329,N_17004,N_17081);
nand U17330 (N_17330,N_17152,N_17114);
and U17331 (N_17331,N_17127,N_17144);
and U17332 (N_17332,N_17117,N_17126);
or U17333 (N_17333,N_17193,N_17159);
nor U17334 (N_17334,N_17077,N_17159);
and U17335 (N_17335,N_17063,N_17080);
or U17336 (N_17336,N_17053,N_17111);
nand U17337 (N_17337,N_17031,N_17163);
nor U17338 (N_17338,N_17075,N_17153);
xnor U17339 (N_17339,N_17198,N_17060);
nand U17340 (N_17340,N_17002,N_17029);
xor U17341 (N_17341,N_17004,N_17132);
or U17342 (N_17342,N_17073,N_17070);
xor U17343 (N_17343,N_17030,N_17105);
and U17344 (N_17344,N_17139,N_17035);
nor U17345 (N_17345,N_17156,N_17066);
xnor U17346 (N_17346,N_17088,N_17084);
or U17347 (N_17347,N_17104,N_17153);
xor U17348 (N_17348,N_17126,N_17131);
and U17349 (N_17349,N_17183,N_17064);
or U17350 (N_17350,N_17072,N_17015);
and U17351 (N_17351,N_17007,N_17096);
nand U17352 (N_17352,N_17069,N_17127);
nand U17353 (N_17353,N_17092,N_17054);
nor U17354 (N_17354,N_17122,N_17116);
nor U17355 (N_17355,N_17199,N_17177);
and U17356 (N_17356,N_17159,N_17092);
and U17357 (N_17357,N_17021,N_17154);
nand U17358 (N_17358,N_17021,N_17165);
nand U17359 (N_17359,N_17182,N_17083);
nor U17360 (N_17360,N_17026,N_17177);
or U17361 (N_17361,N_17088,N_17018);
nor U17362 (N_17362,N_17158,N_17117);
or U17363 (N_17363,N_17191,N_17157);
xor U17364 (N_17364,N_17113,N_17117);
nor U17365 (N_17365,N_17195,N_17196);
and U17366 (N_17366,N_17028,N_17006);
xnor U17367 (N_17367,N_17192,N_17040);
or U17368 (N_17368,N_17190,N_17045);
nand U17369 (N_17369,N_17153,N_17126);
nand U17370 (N_17370,N_17120,N_17109);
nand U17371 (N_17371,N_17068,N_17121);
nand U17372 (N_17372,N_17020,N_17143);
nand U17373 (N_17373,N_17121,N_17095);
nor U17374 (N_17374,N_17169,N_17132);
and U17375 (N_17375,N_17034,N_17168);
nor U17376 (N_17376,N_17018,N_17055);
nand U17377 (N_17377,N_17097,N_17065);
or U17378 (N_17378,N_17080,N_17009);
and U17379 (N_17379,N_17076,N_17149);
and U17380 (N_17380,N_17171,N_17139);
nand U17381 (N_17381,N_17052,N_17172);
or U17382 (N_17382,N_17148,N_17139);
and U17383 (N_17383,N_17154,N_17126);
nand U17384 (N_17384,N_17098,N_17042);
and U17385 (N_17385,N_17142,N_17007);
nand U17386 (N_17386,N_17037,N_17022);
and U17387 (N_17387,N_17123,N_17044);
nand U17388 (N_17388,N_17131,N_17050);
nand U17389 (N_17389,N_17192,N_17157);
nor U17390 (N_17390,N_17100,N_17147);
nor U17391 (N_17391,N_17145,N_17120);
nand U17392 (N_17392,N_17182,N_17063);
nand U17393 (N_17393,N_17166,N_17087);
nand U17394 (N_17394,N_17146,N_17184);
and U17395 (N_17395,N_17083,N_17155);
and U17396 (N_17396,N_17117,N_17141);
or U17397 (N_17397,N_17172,N_17040);
xor U17398 (N_17398,N_17099,N_17047);
or U17399 (N_17399,N_17052,N_17038);
nand U17400 (N_17400,N_17300,N_17333);
and U17401 (N_17401,N_17374,N_17242);
nor U17402 (N_17402,N_17275,N_17303);
or U17403 (N_17403,N_17317,N_17320);
nor U17404 (N_17404,N_17246,N_17273);
or U17405 (N_17405,N_17221,N_17205);
or U17406 (N_17406,N_17288,N_17234);
and U17407 (N_17407,N_17352,N_17269);
nand U17408 (N_17408,N_17314,N_17359);
and U17409 (N_17409,N_17321,N_17394);
or U17410 (N_17410,N_17217,N_17290);
xor U17411 (N_17411,N_17305,N_17247);
nor U17412 (N_17412,N_17383,N_17378);
nand U17413 (N_17413,N_17395,N_17235);
and U17414 (N_17414,N_17384,N_17252);
nand U17415 (N_17415,N_17392,N_17295);
xor U17416 (N_17416,N_17310,N_17233);
xnor U17417 (N_17417,N_17302,N_17325);
or U17418 (N_17418,N_17366,N_17228);
and U17419 (N_17419,N_17338,N_17224);
nor U17420 (N_17420,N_17313,N_17268);
nand U17421 (N_17421,N_17311,N_17243);
nand U17422 (N_17422,N_17360,N_17307);
nand U17423 (N_17423,N_17358,N_17340);
or U17424 (N_17424,N_17294,N_17214);
nor U17425 (N_17425,N_17298,N_17336);
nor U17426 (N_17426,N_17272,N_17347);
nor U17427 (N_17427,N_17372,N_17289);
nor U17428 (N_17428,N_17284,N_17276);
and U17429 (N_17429,N_17373,N_17226);
and U17430 (N_17430,N_17361,N_17223);
and U17431 (N_17431,N_17280,N_17260);
nand U17432 (N_17432,N_17350,N_17238);
nand U17433 (N_17433,N_17281,N_17206);
nor U17434 (N_17434,N_17326,N_17362);
xor U17435 (N_17435,N_17299,N_17344);
or U17436 (N_17436,N_17323,N_17351);
nor U17437 (N_17437,N_17356,N_17379);
or U17438 (N_17438,N_17348,N_17262);
nand U17439 (N_17439,N_17375,N_17283);
and U17440 (N_17440,N_17382,N_17390);
nand U17441 (N_17441,N_17377,N_17346);
nor U17442 (N_17442,N_17318,N_17225);
and U17443 (N_17443,N_17259,N_17343);
or U17444 (N_17444,N_17219,N_17345);
and U17445 (N_17445,N_17253,N_17324);
and U17446 (N_17446,N_17385,N_17327);
or U17447 (N_17447,N_17270,N_17236);
nand U17448 (N_17448,N_17251,N_17264);
and U17449 (N_17449,N_17396,N_17287);
nand U17450 (N_17450,N_17368,N_17204);
or U17451 (N_17451,N_17315,N_17337);
and U17452 (N_17452,N_17387,N_17399);
nand U17453 (N_17453,N_17386,N_17200);
and U17454 (N_17454,N_17319,N_17391);
nor U17455 (N_17455,N_17210,N_17255);
nand U17456 (N_17456,N_17263,N_17257);
xnor U17457 (N_17457,N_17208,N_17388);
nor U17458 (N_17458,N_17254,N_17279);
xor U17459 (N_17459,N_17330,N_17258);
xnor U17460 (N_17460,N_17293,N_17371);
xnor U17461 (N_17461,N_17277,N_17370);
or U17462 (N_17462,N_17232,N_17357);
nor U17463 (N_17463,N_17297,N_17278);
nor U17464 (N_17464,N_17355,N_17244);
and U17465 (N_17465,N_17286,N_17237);
or U17466 (N_17466,N_17292,N_17339);
or U17467 (N_17467,N_17349,N_17261);
or U17468 (N_17468,N_17213,N_17265);
and U17469 (N_17469,N_17239,N_17304);
or U17470 (N_17470,N_17354,N_17309);
and U17471 (N_17471,N_17381,N_17249);
nand U17472 (N_17472,N_17222,N_17308);
and U17473 (N_17473,N_17245,N_17291);
nor U17474 (N_17474,N_17398,N_17241);
nor U17475 (N_17475,N_17282,N_17365);
xnor U17476 (N_17476,N_17301,N_17202);
or U17477 (N_17477,N_17363,N_17267);
and U17478 (N_17478,N_17231,N_17329);
xor U17479 (N_17479,N_17216,N_17207);
and U17480 (N_17480,N_17215,N_17389);
nor U17481 (N_17481,N_17201,N_17397);
nand U17482 (N_17482,N_17271,N_17229);
and U17483 (N_17483,N_17230,N_17248);
and U17484 (N_17484,N_17335,N_17250);
or U17485 (N_17485,N_17209,N_17240);
and U17486 (N_17486,N_17285,N_17369);
xnor U17487 (N_17487,N_17331,N_17342);
nand U17488 (N_17488,N_17212,N_17266);
or U17489 (N_17489,N_17353,N_17306);
nor U17490 (N_17490,N_17218,N_17380);
or U17491 (N_17491,N_17393,N_17296);
nor U17492 (N_17492,N_17203,N_17211);
nand U17493 (N_17493,N_17220,N_17328);
or U17494 (N_17494,N_17341,N_17334);
or U17495 (N_17495,N_17256,N_17332);
and U17496 (N_17496,N_17312,N_17227);
nand U17497 (N_17497,N_17316,N_17364);
nor U17498 (N_17498,N_17274,N_17376);
nand U17499 (N_17499,N_17322,N_17367);
nor U17500 (N_17500,N_17377,N_17394);
and U17501 (N_17501,N_17293,N_17325);
nand U17502 (N_17502,N_17202,N_17376);
and U17503 (N_17503,N_17343,N_17366);
or U17504 (N_17504,N_17349,N_17316);
or U17505 (N_17505,N_17273,N_17396);
nor U17506 (N_17506,N_17352,N_17338);
nand U17507 (N_17507,N_17277,N_17329);
xor U17508 (N_17508,N_17336,N_17277);
nand U17509 (N_17509,N_17365,N_17369);
nand U17510 (N_17510,N_17310,N_17226);
nor U17511 (N_17511,N_17335,N_17306);
nor U17512 (N_17512,N_17352,N_17357);
xnor U17513 (N_17513,N_17356,N_17264);
nor U17514 (N_17514,N_17398,N_17201);
and U17515 (N_17515,N_17313,N_17284);
and U17516 (N_17516,N_17382,N_17237);
or U17517 (N_17517,N_17230,N_17206);
xnor U17518 (N_17518,N_17331,N_17286);
nor U17519 (N_17519,N_17283,N_17205);
xor U17520 (N_17520,N_17346,N_17262);
nor U17521 (N_17521,N_17379,N_17322);
nand U17522 (N_17522,N_17202,N_17271);
or U17523 (N_17523,N_17241,N_17349);
nor U17524 (N_17524,N_17268,N_17290);
xnor U17525 (N_17525,N_17283,N_17237);
nor U17526 (N_17526,N_17217,N_17337);
or U17527 (N_17527,N_17310,N_17223);
and U17528 (N_17528,N_17277,N_17294);
nand U17529 (N_17529,N_17279,N_17319);
nor U17530 (N_17530,N_17396,N_17266);
nor U17531 (N_17531,N_17210,N_17243);
or U17532 (N_17532,N_17333,N_17230);
nor U17533 (N_17533,N_17387,N_17324);
xnor U17534 (N_17534,N_17390,N_17252);
and U17535 (N_17535,N_17309,N_17290);
or U17536 (N_17536,N_17283,N_17286);
nand U17537 (N_17537,N_17345,N_17209);
nor U17538 (N_17538,N_17283,N_17374);
nor U17539 (N_17539,N_17256,N_17349);
nor U17540 (N_17540,N_17262,N_17332);
and U17541 (N_17541,N_17225,N_17396);
and U17542 (N_17542,N_17380,N_17341);
and U17543 (N_17543,N_17391,N_17218);
nand U17544 (N_17544,N_17375,N_17277);
or U17545 (N_17545,N_17278,N_17253);
nand U17546 (N_17546,N_17275,N_17374);
or U17547 (N_17547,N_17347,N_17209);
nor U17548 (N_17548,N_17313,N_17220);
nand U17549 (N_17549,N_17209,N_17382);
nand U17550 (N_17550,N_17390,N_17331);
nand U17551 (N_17551,N_17217,N_17358);
xor U17552 (N_17552,N_17311,N_17365);
nand U17553 (N_17553,N_17388,N_17281);
nand U17554 (N_17554,N_17204,N_17391);
xnor U17555 (N_17555,N_17386,N_17290);
or U17556 (N_17556,N_17372,N_17362);
or U17557 (N_17557,N_17389,N_17351);
nor U17558 (N_17558,N_17213,N_17337);
and U17559 (N_17559,N_17283,N_17247);
xnor U17560 (N_17560,N_17244,N_17388);
nand U17561 (N_17561,N_17312,N_17235);
xor U17562 (N_17562,N_17368,N_17244);
and U17563 (N_17563,N_17260,N_17336);
and U17564 (N_17564,N_17384,N_17326);
or U17565 (N_17565,N_17210,N_17357);
or U17566 (N_17566,N_17392,N_17334);
and U17567 (N_17567,N_17243,N_17245);
or U17568 (N_17568,N_17267,N_17227);
and U17569 (N_17569,N_17337,N_17383);
nand U17570 (N_17570,N_17381,N_17371);
nand U17571 (N_17571,N_17367,N_17227);
nor U17572 (N_17572,N_17349,N_17362);
nand U17573 (N_17573,N_17391,N_17345);
nor U17574 (N_17574,N_17343,N_17277);
nand U17575 (N_17575,N_17351,N_17329);
and U17576 (N_17576,N_17207,N_17355);
nand U17577 (N_17577,N_17242,N_17268);
nor U17578 (N_17578,N_17318,N_17395);
and U17579 (N_17579,N_17253,N_17200);
nand U17580 (N_17580,N_17240,N_17320);
or U17581 (N_17581,N_17218,N_17398);
nor U17582 (N_17582,N_17343,N_17391);
nand U17583 (N_17583,N_17237,N_17345);
or U17584 (N_17584,N_17256,N_17357);
nand U17585 (N_17585,N_17384,N_17230);
and U17586 (N_17586,N_17267,N_17318);
or U17587 (N_17587,N_17396,N_17341);
and U17588 (N_17588,N_17248,N_17228);
nand U17589 (N_17589,N_17377,N_17261);
xnor U17590 (N_17590,N_17311,N_17204);
nand U17591 (N_17591,N_17238,N_17226);
nor U17592 (N_17592,N_17326,N_17346);
or U17593 (N_17593,N_17257,N_17383);
and U17594 (N_17594,N_17259,N_17330);
nor U17595 (N_17595,N_17275,N_17373);
nor U17596 (N_17596,N_17229,N_17387);
and U17597 (N_17597,N_17271,N_17367);
nor U17598 (N_17598,N_17375,N_17217);
nand U17599 (N_17599,N_17238,N_17206);
xor U17600 (N_17600,N_17514,N_17467);
and U17601 (N_17601,N_17548,N_17541);
or U17602 (N_17602,N_17592,N_17402);
nand U17603 (N_17603,N_17565,N_17481);
or U17604 (N_17604,N_17539,N_17409);
or U17605 (N_17605,N_17598,N_17569);
nand U17606 (N_17606,N_17554,N_17410);
nor U17607 (N_17607,N_17505,N_17599);
or U17608 (N_17608,N_17543,N_17479);
nor U17609 (N_17609,N_17401,N_17421);
xnor U17610 (N_17610,N_17491,N_17536);
nand U17611 (N_17611,N_17446,N_17485);
nand U17612 (N_17612,N_17549,N_17597);
and U17613 (N_17613,N_17494,N_17460);
nor U17614 (N_17614,N_17480,N_17468);
nor U17615 (N_17615,N_17492,N_17453);
or U17616 (N_17616,N_17438,N_17596);
nand U17617 (N_17617,N_17506,N_17507);
nor U17618 (N_17618,N_17466,N_17593);
or U17619 (N_17619,N_17447,N_17452);
nand U17620 (N_17620,N_17591,N_17576);
xor U17621 (N_17621,N_17420,N_17566);
xnor U17622 (N_17622,N_17477,N_17581);
nand U17623 (N_17623,N_17583,N_17568);
or U17624 (N_17624,N_17499,N_17572);
or U17625 (N_17625,N_17483,N_17472);
nor U17626 (N_17626,N_17462,N_17443);
nand U17627 (N_17627,N_17423,N_17442);
nor U17628 (N_17628,N_17510,N_17573);
nor U17629 (N_17629,N_17450,N_17474);
or U17630 (N_17630,N_17528,N_17445);
nand U17631 (N_17631,N_17411,N_17493);
or U17632 (N_17632,N_17535,N_17545);
nand U17633 (N_17633,N_17415,N_17590);
nand U17634 (N_17634,N_17585,N_17439);
nor U17635 (N_17635,N_17512,N_17589);
and U17636 (N_17636,N_17487,N_17521);
xor U17637 (N_17637,N_17414,N_17551);
or U17638 (N_17638,N_17555,N_17503);
or U17639 (N_17639,N_17553,N_17513);
nand U17640 (N_17640,N_17488,N_17407);
or U17641 (N_17641,N_17461,N_17449);
or U17642 (N_17642,N_17559,N_17463);
nor U17643 (N_17643,N_17594,N_17522);
and U17644 (N_17644,N_17464,N_17511);
and U17645 (N_17645,N_17455,N_17509);
nand U17646 (N_17646,N_17562,N_17556);
nand U17647 (N_17647,N_17557,N_17534);
nor U17648 (N_17648,N_17434,N_17575);
or U17649 (N_17649,N_17425,N_17588);
xnor U17650 (N_17650,N_17489,N_17437);
nor U17651 (N_17651,N_17470,N_17473);
and U17652 (N_17652,N_17564,N_17459);
nor U17653 (N_17653,N_17501,N_17523);
xnor U17654 (N_17654,N_17582,N_17570);
nand U17655 (N_17655,N_17502,N_17403);
nand U17656 (N_17656,N_17400,N_17586);
and U17657 (N_17657,N_17426,N_17563);
nand U17658 (N_17658,N_17406,N_17404);
or U17659 (N_17659,N_17515,N_17440);
nor U17660 (N_17660,N_17577,N_17433);
nand U17661 (N_17661,N_17417,N_17490);
and U17662 (N_17662,N_17432,N_17448);
or U17663 (N_17663,N_17529,N_17516);
or U17664 (N_17664,N_17544,N_17419);
nand U17665 (N_17665,N_17422,N_17475);
nor U17666 (N_17666,N_17574,N_17441);
and U17667 (N_17667,N_17495,N_17435);
or U17668 (N_17668,N_17413,N_17476);
xnor U17669 (N_17669,N_17542,N_17469);
nand U17670 (N_17670,N_17532,N_17517);
nor U17671 (N_17671,N_17436,N_17428);
or U17672 (N_17672,N_17500,N_17584);
nand U17673 (N_17673,N_17465,N_17427);
and U17674 (N_17674,N_17546,N_17524);
xnor U17675 (N_17675,N_17454,N_17537);
nor U17676 (N_17676,N_17531,N_17580);
and U17677 (N_17677,N_17408,N_17497);
xnor U17678 (N_17678,N_17571,N_17456);
nor U17679 (N_17679,N_17504,N_17405);
and U17680 (N_17680,N_17482,N_17451);
or U17681 (N_17681,N_17579,N_17486);
nor U17682 (N_17682,N_17416,N_17538);
nor U17683 (N_17683,N_17431,N_17484);
or U17684 (N_17684,N_17525,N_17508);
and U17685 (N_17685,N_17587,N_17496);
nor U17686 (N_17686,N_17444,N_17560);
xnor U17687 (N_17687,N_17561,N_17429);
nand U17688 (N_17688,N_17547,N_17578);
or U17689 (N_17689,N_17526,N_17550);
or U17690 (N_17690,N_17498,N_17527);
and U17691 (N_17691,N_17558,N_17424);
or U17692 (N_17692,N_17533,N_17595);
and U17693 (N_17693,N_17471,N_17458);
or U17694 (N_17694,N_17430,N_17478);
and U17695 (N_17695,N_17412,N_17540);
nor U17696 (N_17696,N_17418,N_17520);
and U17697 (N_17697,N_17552,N_17519);
or U17698 (N_17698,N_17518,N_17530);
and U17699 (N_17699,N_17567,N_17457);
nand U17700 (N_17700,N_17546,N_17592);
or U17701 (N_17701,N_17418,N_17442);
nor U17702 (N_17702,N_17427,N_17415);
nor U17703 (N_17703,N_17485,N_17562);
nand U17704 (N_17704,N_17525,N_17557);
and U17705 (N_17705,N_17464,N_17421);
nor U17706 (N_17706,N_17412,N_17402);
nor U17707 (N_17707,N_17477,N_17542);
nor U17708 (N_17708,N_17537,N_17405);
nand U17709 (N_17709,N_17489,N_17447);
nor U17710 (N_17710,N_17408,N_17594);
nand U17711 (N_17711,N_17436,N_17540);
or U17712 (N_17712,N_17429,N_17445);
xor U17713 (N_17713,N_17582,N_17575);
or U17714 (N_17714,N_17553,N_17455);
nor U17715 (N_17715,N_17552,N_17579);
xnor U17716 (N_17716,N_17451,N_17400);
nand U17717 (N_17717,N_17572,N_17522);
nor U17718 (N_17718,N_17527,N_17547);
and U17719 (N_17719,N_17488,N_17591);
xnor U17720 (N_17720,N_17533,N_17586);
or U17721 (N_17721,N_17485,N_17448);
nor U17722 (N_17722,N_17552,N_17561);
nand U17723 (N_17723,N_17425,N_17563);
nand U17724 (N_17724,N_17476,N_17473);
and U17725 (N_17725,N_17542,N_17559);
and U17726 (N_17726,N_17570,N_17529);
nand U17727 (N_17727,N_17546,N_17455);
nand U17728 (N_17728,N_17444,N_17515);
nand U17729 (N_17729,N_17578,N_17441);
or U17730 (N_17730,N_17563,N_17411);
or U17731 (N_17731,N_17411,N_17495);
nor U17732 (N_17732,N_17433,N_17455);
or U17733 (N_17733,N_17482,N_17431);
xor U17734 (N_17734,N_17580,N_17539);
or U17735 (N_17735,N_17416,N_17419);
nor U17736 (N_17736,N_17523,N_17563);
nor U17737 (N_17737,N_17503,N_17568);
and U17738 (N_17738,N_17471,N_17567);
and U17739 (N_17739,N_17441,N_17446);
nand U17740 (N_17740,N_17536,N_17413);
xor U17741 (N_17741,N_17432,N_17461);
or U17742 (N_17742,N_17416,N_17512);
and U17743 (N_17743,N_17545,N_17567);
nor U17744 (N_17744,N_17407,N_17403);
nand U17745 (N_17745,N_17529,N_17411);
nor U17746 (N_17746,N_17424,N_17520);
nand U17747 (N_17747,N_17436,N_17432);
nand U17748 (N_17748,N_17583,N_17446);
and U17749 (N_17749,N_17555,N_17498);
nand U17750 (N_17750,N_17438,N_17551);
or U17751 (N_17751,N_17429,N_17496);
and U17752 (N_17752,N_17536,N_17596);
nor U17753 (N_17753,N_17439,N_17580);
nor U17754 (N_17754,N_17510,N_17525);
or U17755 (N_17755,N_17537,N_17491);
nand U17756 (N_17756,N_17473,N_17554);
xor U17757 (N_17757,N_17435,N_17593);
xnor U17758 (N_17758,N_17483,N_17508);
or U17759 (N_17759,N_17592,N_17527);
and U17760 (N_17760,N_17478,N_17464);
nor U17761 (N_17761,N_17449,N_17512);
nand U17762 (N_17762,N_17416,N_17575);
and U17763 (N_17763,N_17465,N_17530);
xor U17764 (N_17764,N_17453,N_17572);
xor U17765 (N_17765,N_17483,N_17433);
nand U17766 (N_17766,N_17459,N_17512);
and U17767 (N_17767,N_17443,N_17541);
or U17768 (N_17768,N_17431,N_17487);
nor U17769 (N_17769,N_17419,N_17554);
xnor U17770 (N_17770,N_17571,N_17567);
or U17771 (N_17771,N_17562,N_17453);
nand U17772 (N_17772,N_17445,N_17550);
or U17773 (N_17773,N_17532,N_17596);
nor U17774 (N_17774,N_17513,N_17454);
nand U17775 (N_17775,N_17543,N_17473);
and U17776 (N_17776,N_17594,N_17452);
xnor U17777 (N_17777,N_17457,N_17597);
xor U17778 (N_17778,N_17526,N_17560);
xor U17779 (N_17779,N_17550,N_17452);
or U17780 (N_17780,N_17410,N_17499);
and U17781 (N_17781,N_17416,N_17443);
and U17782 (N_17782,N_17551,N_17503);
or U17783 (N_17783,N_17597,N_17494);
or U17784 (N_17784,N_17511,N_17536);
nor U17785 (N_17785,N_17584,N_17566);
nand U17786 (N_17786,N_17568,N_17426);
nand U17787 (N_17787,N_17544,N_17531);
or U17788 (N_17788,N_17403,N_17510);
nand U17789 (N_17789,N_17561,N_17482);
nor U17790 (N_17790,N_17536,N_17589);
xor U17791 (N_17791,N_17437,N_17595);
nand U17792 (N_17792,N_17477,N_17525);
nor U17793 (N_17793,N_17554,N_17411);
and U17794 (N_17794,N_17448,N_17460);
or U17795 (N_17795,N_17546,N_17525);
nor U17796 (N_17796,N_17521,N_17505);
or U17797 (N_17797,N_17546,N_17574);
nand U17798 (N_17798,N_17444,N_17429);
nand U17799 (N_17799,N_17449,N_17587);
xnor U17800 (N_17800,N_17770,N_17791);
or U17801 (N_17801,N_17600,N_17604);
and U17802 (N_17802,N_17727,N_17681);
or U17803 (N_17803,N_17665,N_17653);
nand U17804 (N_17804,N_17633,N_17629);
and U17805 (N_17805,N_17794,N_17786);
nand U17806 (N_17806,N_17729,N_17637);
or U17807 (N_17807,N_17660,N_17667);
xnor U17808 (N_17808,N_17743,N_17669);
and U17809 (N_17809,N_17776,N_17643);
and U17810 (N_17810,N_17623,N_17734);
or U17811 (N_17811,N_17671,N_17603);
and U17812 (N_17812,N_17718,N_17746);
or U17813 (N_17813,N_17764,N_17783);
or U17814 (N_17814,N_17748,N_17687);
nand U17815 (N_17815,N_17676,N_17608);
or U17816 (N_17816,N_17679,N_17750);
nor U17817 (N_17817,N_17722,N_17787);
nand U17818 (N_17818,N_17741,N_17702);
nor U17819 (N_17819,N_17630,N_17714);
nand U17820 (N_17820,N_17758,N_17773);
and U17821 (N_17821,N_17744,N_17733);
nand U17822 (N_17822,N_17663,N_17710);
nor U17823 (N_17823,N_17641,N_17767);
nand U17824 (N_17824,N_17726,N_17703);
nand U17825 (N_17825,N_17693,N_17615);
nand U17826 (N_17826,N_17697,N_17708);
nor U17827 (N_17827,N_17700,N_17793);
nor U17828 (N_17828,N_17607,N_17652);
nor U17829 (N_17829,N_17745,N_17752);
xnor U17830 (N_17830,N_17619,N_17685);
nand U17831 (N_17831,N_17605,N_17650);
xnor U17832 (N_17832,N_17659,N_17649);
nand U17833 (N_17833,N_17716,N_17784);
and U17834 (N_17834,N_17684,N_17774);
nand U17835 (N_17835,N_17728,N_17781);
nand U17836 (N_17836,N_17622,N_17709);
and U17837 (N_17837,N_17680,N_17725);
nand U17838 (N_17838,N_17740,N_17717);
nand U17839 (N_17839,N_17614,N_17631);
nor U17840 (N_17840,N_17672,N_17769);
nand U17841 (N_17841,N_17715,N_17755);
nor U17842 (N_17842,N_17624,N_17797);
and U17843 (N_17843,N_17670,N_17602);
and U17844 (N_17844,N_17747,N_17668);
and U17845 (N_17845,N_17756,N_17677);
xor U17846 (N_17846,N_17648,N_17705);
and U17847 (N_17847,N_17739,N_17768);
or U17848 (N_17848,N_17759,N_17642);
and U17849 (N_17849,N_17712,N_17606);
or U17850 (N_17850,N_17707,N_17673);
or U17851 (N_17851,N_17654,N_17790);
nand U17852 (N_17852,N_17634,N_17742);
nor U17853 (N_17853,N_17628,N_17699);
nand U17854 (N_17854,N_17620,N_17788);
nand U17855 (N_17855,N_17611,N_17675);
nor U17856 (N_17856,N_17735,N_17775);
nand U17857 (N_17857,N_17798,N_17780);
or U17858 (N_17858,N_17640,N_17662);
or U17859 (N_17859,N_17638,N_17753);
nand U17860 (N_17860,N_17706,N_17738);
nor U17861 (N_17861,N_17772,N_17632);
xnor U17862 (N_17862,N_17711,N_17760);
nor U17863 (N_17863,N_17658,N_17730);
and U17864 (N_17864,N_17757,N_17689);
and U17865 (N_17865,N_17656,N_17799);
or U17866 (N_17866,N_17701,N_17645);
nor U17867 (N_17867,N_17795,N_17779);
and U17868 (N_17868,N_17749,N_17639);
and U17869 (N_17869,N_17792,N_17616);
and U17870 (N_17870,N_17751,N_17723);
or U17871 (N_17871,N_17657,N_17736);
and U17872 (N_17872,N_17651,N_17771);
nor U17873 (N_17873,N_17683,N_17796);
xnor U17874 (N_17874,N_17610,N_17761);
xnor U17875 (N_17875,N_17635,N_17636);
nand U17876 (N_17876,N_17782,N_17789);
nand U17877 (N_17877,N_17785,N_17690);
or U17878 (N_17878,N_17762,N_17691);
nand U17879 (N_17879,N_17626,N_17704);
nand U17880 (N_17880,N_17621,N_17609);
nor U17881 (N_17881,N_17766,N_17601);
nor U17882 (N_17882,N_17666,N_17688);
nand U17883 (N_17883,N_17618,N_17724);
nor U17884 (N_17884,N_17719,N_17674);
nand U17885 (N_17885,N_17627,N_17678);
and U17886 (N_17886,N_17765,N_17754);
nor U17887 (N_17887,N_17612,N_17694);
or U17888 (N_17888,N_17720,N_17731);
and U17889 (N_17889,N_17698,N_17777);
or U17890 (N_17890,N_17613,N_17737);
nor U17891 (N_17891,N_17647,N_17695);
or U17892 (N_17892,N_17644,N_17661);
or U17893 (N_17893,N_17646,N_17778);
or U17894 (N_17894,N_17686,N_17664);
or U17895 (N_17895,N_17763,N_17625);
xor U17896 (N_17896,N_17617,N_17655);
or U17897 (N_17897,N_17696,N_17692);
nor U17898 (N_17898,N_17721,N_17682);
nand U17899 (N_17899,N_17713,N_17732);
nor U17900 (N_17900,N_17642,N_17603);
or U17901 (N_17901,N_17606,N_17611);
or U17902 (N_17902,N_17712,N_17779);
nand U17903 (N_17903,N_17694,N_17670);
or U17904 (N_17904,N_17789,N_17613);
and U17905 (N_17905,N_17615,N_17740);
and U17906 (N_17906,N_17780,N_17682);
and U17907 (N_17907,N_17708,N_17737);
nor U17908 (N_17908,N_17664,N_17774);
and U17909 (N_17909,N_17749,N_17755);
or U17910 (N_17910,N_17747,N_17611);
xor U17911 (N_17911,N_17715,N_17608);
or U17912 (N_17912,N_17776,N_17696);
nor U17913 (N_17913,N_17649,N_17687);
or U17914 (N_17914,N_17734,N_17672);
nor U17915 (N_17915,N_17743,N_17678);
nand U17916 (N_17916,N_17668,N_17738);
xor U17917 (N_17917,N_17662,N_17730);
and U17918 (N_17918,N_17793,N_17770);
and U17919 (N_17919,N_17680,N_17757);
and U17920 (N_17920,N_17644,N_17609);
or U17921 (N_17921,N_17629,N_17767);
nand U17922 (N_17922,N_17603,N_17782);
and U17923 (N_17923,N_17613,N_17670);
and U17924 (N_17924,N_17744,N_17626);
and U17925 (N_17925,N_17722,N_17752);
nor U17926 (N_17926,N_17765,N_17739);
or U17927 (N_17927,N_17759,N_17656);
or U17928 (N_17928,N_17613,N_17681);
or U17929 (N_17929,N_17784,N_17790);
and U17930 (N_17930,N_17732,N_17618);
nand U17931 (N_17931,N_17688,N_17619);
and U17932 (N_17932,N_17715,N_17721);
and U17933 (N_17933,N_17610,N_17781);
nor U17934 (N_17934,N_17698,N_17634);
or U17935 (N_17935,N_17630,N_17664);
and U17936 (N_17936,N_17796,N_17741);
or U17937 (N_17937,N_17746,N_17728);
or U17938 (N_17938,N_17627,N_17601);
or U17939 (N_17939,N_17739,N_17691);
or U17940 (N_17940,N_17636,N_17655);
nor U17941 (N_17941,N_17630,N_17767);
xor U17942 (N_17942,N_17629,N_17666);
nor U17943 (N_17943,N_17711,N_17679);
and U17944 (N_17944,N_17721,N_17798);
xnor U17945 (N_17945,N_17719,N_17662);
nor U17946 (N_17946,N_17690,N_17662);
xor U17947 (N_17947,N_17756,N_17600);
xor U17948 (N_17948,N_17781,N_17674);
and U17949 (N_17949,N_17655,N_17649);
nor U17950 (N_17950,N_17611,N_17749);
nand U17951 (N_17951,N_17664,N_17771);
nor U17952 (N_17952,N_17776,N_17634);
and U17953 (N_17953,N_17754,N_17679);
nand U17954 (N_17954,N_17732,N_17638);
nand U17955 (N_17955,N_17761,N_17797);
xor U17956 (N_17956,N_17632,N_17748);
nor U17957 (N_17957,N_17660,N_17763);
and U17958 (N_17958,N_17791,N_17647);
and U17959 (N_17959,N_17784,N_17654);
nor U17960 (N_17960,N_17706,N_17766);
nor U17961 (N_17961,N_17719,N_17661);
nor U17962 (N_17962,N_17736,N_17681);
xnor U17963 (N_17963,N_17648,N_17775);
nand U17964 (N_17964,N_17674,N_17661);
nand U17965 (N_17965,N_17651,N_17686);
or U17966 (N_17966,N_17604,N_17749);
or U17967 (N_17967,N_17711,N_17671);
and U17968 (N_17968,N_17622,N_17640);
xor U17969 (N_17969,N_17656,N_17744);
nand U17970 (N_17970,N_17631,N_17645);
or U17971 (N_17971,N_17628,N_17622);
nand U17972 (N_17972,N_17619,N_17630);
nand U17973 (N_17973,N_17639,N_17740);
or U17974 (N_17974,N_17679,N_17656);
and U17975 (N_17975,N_17618,N_17731);
nor U17976 (N_17976,N_17795,N_17759);
and U17977 (N_17977,N_17795,N_17602);
or U17978 (N_17978,N_17623,N_17716);
nand U17979 (N_17979,N_17687,N_17608);
xnor U17980 (N_17980,N_17709,N_17727);
or U17981 (N_17981,N_17695,N_17660);
or U17982 (N_17982,N_17761,N_17738);
or U17983 (N_17983,N_17718,N_17682);
xnor U17984 (N_17984,N_17766,N_17697);
and U17985 (N_17985,N_17722,N_17768);
or U17986 (N_17986,N_17717,N_17751);
xnor U17987 (N_17987,N_17654,N_17651);
or U17988 (N_17988,N_17686,N_17786);
and U17989 (N_17989,N_17791,N_17724);
nor U17990 (N_17990,N_17737,N_17721);
nor U17991 (N_17991,N_17692,N_17742);
and U17992 (N_17992,N_17750,N_17667);
or U17993 (N_17993,N_17738,N_17760);
nand U17994 (N_17994,N_17649,N_17714);
nor U17995 (N_17995,N_17792,N_17670);
or U17996 (N_17996,N_17706,N_17747);
nand U17997 (N_17997,N_17745,N_17648);
nor U17998 (N_17998,N_17774,N_17632);
xor U17999 (N_17999,N_17681,N_17744);
and U18000 (N_18000,N_17837,N_17920);
or U18001 (N_18001,N_17852,N_17968);
or U18002 (N_18002,N_17856,N_17842);
nand U18003 (N_18003,N_17824,N_17877);
nor U18004 (N_18004,N_17857,N_17889);
nand U18005 (N_18005,N_17953,N_17850);
or U18006 (N_18006,N_17921,N_17872);
and U18007 (N_18007,N_17887,N_17975);
and U18008 (N_18008,N_17870,N_17943);
nand U18009 (N_18009,N_17977,N_17853);
nor U18010 (N_18010,N_17809,N_17838);
nor U18011 (N_18011,N_17983,N_17956);
or U18012 (N_18012,N_17976,N_17923);
nor U18013 (N_18013,N_17801,N_17884);
nand U18014 (N_18014,N_17836,N_17875);
and U18015 (N_18015,N_17833,N_17944);
or U18016 (N_18016,N_17819,N_17947);
or U18017 (N_18017,N_17807,N_17902);
nor U18018 (N_18018,N_17969,N_17961);
or U18019 (N_18019,N_17992,N_17903);
nand U18020 (N_18020,N_17967,N_17821);
and U18021 (N_18021,N_17803,N_17997);
or U18022 (N_18022,N_17922,N_17813);
nor U18023 (N_18023,N_17994,N_17957);
nand U18024 (N_18024,N_17843,N_17805);
or U18025 (N_18025,N_17892,N_17941);
or U18026 (N_18026,N_17907,N_17945);
or U18027 (N_18027,N_17908,N_17873);
nor U18028 (N_18028,N_17881,N_17904);
nand U18029 (N_18029,N_17937,N_17885);
nand U18030 (N_18030,N_17986,N_17825);
xor U18031 (N_18031,N_17935,N_17839);
nand U18032 (N_18032,N_17959,N_17864);
nand U18033 (N_18033,N_17913,N_17849);
or U18034 (N_18034,N_17980,N_17909);
nor U18035 (N_18035,N_17895,N_17826);
nand U18036 (N_18036,N_17919,N_17874);
or U18037 (N_18037,N_17954,N_17830);
and U18038 (N_18038,N_17806,N_17800);
or U18039 (N_18039,N_17886,N_17844);
and U18040 (N_18040,N_17829,N_17979);
nand U18041 (N_18041,N_17946,N_17942);
and U18042 (N_18042,N_17859,N_17905);
nand U18043 (N_18043,N_17910,N_17893);
and U18044 (N_18044,N_17900,N_17999);
nand U18045 (N_18045,N_17860,N_17912);
nor U18046 (N_18046,N_17862,N_17939);
xor U18047 (N_18047,N_17985,N_17840);
nor U18048 (N_18048,N_17869,N_17896);
nor U18049 (N_18049,N_17934,N_17820);
nor U18050 (N_18050,N_17906,N_17911);
and U18051 (N_18051,N_17822,N_17938);
and U18052 (N_18052,N_17970,N_17928);
nor U18053 (N_18053,N_17878,N_17816);
and U18054 (N_18054,N_17933,N_17998);
nor U18055 (N_18055,N_17828,N_17931);
or U18056 (N_18056,N_17880,N_17901);
nor U18057 (N_18057,N_17974,N_17841);
nor U18058 (N_18058,N_17832,N_17972);
nor U18059 (N_18059,N_17831,N_17810);
or U18060 (N_18060,N_17924,N_17846);
nand U18061 (N_18061,N_17865,N_17991);
nand U18062 (N_18062,N_17802,N_17894);
xor U18063 (N_18063,N_17882,N_17823);
nor U18064 (N_18064,N_17989,N_17918);
nand U18065 (N_18065,N_17812,N_17835);
and U18066 (N_18066,N_17995,N_17890);
or U18067 (N_18067,N_17854,N_17930);
or U18068 (N_18068,N_17964,N_17915);
nand U18069 (N_18069,N_17932,N_17811);
and U18070 (N_18070,N_17868,N_17815);
nand U18071 (N_18071,N_17888,N_17987);
xnor U18072 (N_18072,N_17982,N_17960);
and U18073 (N_18073,N_17847,N_17867);
nand U18074 (N_18074,N_17978,N_17817);
nand U18075 (N_18075,N_17827,N_17804);
and U18076 (N_18076,N_17927,N_17971);
nand U18077 (N_18077,N_17984,N_17899);
or U18078 (N_18078,N_17950,N_17808);
xor U18079 (N_18079,N_17925,N_17965);
and U18080 (N_18080,N_17973,N_17958);
nor U18081 (N_18081,N_17996,N_17990);
or U18082 (N_18082,N_17951,N_17871);
xor U18083 (N_18083,N_17858,N_17926);
and U18084 (N_18084,N_17949,N_17866);
xor U18085 (N_18085,N_17917,N_17940);
or U18086 (N_18086,N_17845,N_17834);
xor U18087 (N_18087,N_17963,N_17898);
xnor U18088 (N_18088,N_17818,N_17981);
or U18089 (N_18089,N_17851,N_17966);
and U18090 (N_18090,N_17879,N_17891);
or U18091 (N_18091,N_17883,N_17955);
nor U18092 (N_18092,N_17814,N_17936);
nand U18093 (N_18093,N_17929,N_17952);
or U18094 (N_18094,N_17861,N_17876);
nor U18095 (N_18095,N_17916,N_17897);
and U18096 (N_18096,N_17962,N_17948);
or U18097 (N_18097,N_17914,N_17863);
or U18098 (N_18098,N_17848,N_17855);
nor U18099 (N_18099,N_17988,N_17993);
nor U18100 (N_18100,N_17875,N_17819);
and U18101 (N_18101,N_17908,N_17864);
and U18102 (N_18102,N_17962,N_17802);
and U18103 (N_18103,N_17995,N_17827);
xor U18104 (N_18104,N_17967,N_17890);
and U18105 (N_18105,N_17937,N_17952);
and U18106 (N_18106,N_17893,N_17843);
and U18107 (N_18107,N_17957,N_17960);
nor U18108 (N_18108,N_17956,N_17998);
and U18109 (N_18109,N_17968,N_17982);
and U18110 (N_18110,N_17943,N_17824);
nor U18111 (N_18111,N_17977,N_17850);
or U18112 (N_18112,N_17853,N_17976);
nand U18113 (N_18113,N_17828,N_17904);
or U18114 (N_18114,N_17871,N_17814);
nor U18115 (N_18115,N_17876,N_17992);
or U18116 (N_18116,N_17915,N_17973);
nand U18117 (N_18117,N_17811,N_17983);
or U18118 (N_18118,N_17964,N_17896);
or U18119 (N_18119,N_17856,N_17968);
or U18120 (N_18120,N_17985,N_17848);
nor U18121 (N_18121,N_17822,N_17961);
nand U18122 (N_18122,N_17945,N_17852);
nand U18123 (N_18123,N_17833,N_17808);
xor U18124 (N_18124,N_17989,N_17833);
nand U18125 (N_18125,N_17898,N_17997);
nand U18126 (N_18126,N_17961,N_17949);
xor U18127 (N_18127,N_17891,N_17886);
or U18128 (N_18128,N_17801,N_17867);
xnor U18129 (N_18129,N_17996,N_17897);
and U18130 (N_18130,N_17926,N_17982);
or U18131 (N_18131,N_17883,N_17948);
and U18132 (N_18132,N_17947,N_17807);
nand U18133 (N_18133,N_17818,N_17977);
and U18134 (N_18134,N_17803,N_17976);
or U18135 (N_18135,N_17825,N_17938);
xor U18136 (N_18136,N_17852,N_17906);
and U18137 (N_18137,N_17857,N_17866);
xor U18138 (N_18138,N_17990,N_17830);
nand U18139 (N_18139,N_17966,N_17870);
or U18140 (N_18140,N_17973,N_17856);
nor U18141 (N_18141,N_17983,N_17820);
or U18142 (N_18142,N_17963,N_17863);
nand U18143 (N_18143,N_17991,N_17816);
or U18144 (N_18144,N_17961,N_17853);
nor U18145 (N_18145,N_17997,N_17902);
and U18146 (N_18146,N_17917,N_17895);
or U18147 (N_18147,N_17971,N_17843);
nor U18148 (N_18148,N_17851,N_17819);
nand U18149 (N_18149,N_17881,N_17971);
nand U18150 (N_18150,N_17852,N_17868);
or U18151 (N_18151,N_17849,N_17897);
or U18152 (N_18152,N_17824,N_17821);
and U18153 (N_18153,N_17977,N_17941);
and U18154 (N_18154,N_17807,N_17994);
and U18155 (N_18155,N_17987,N_17856);
or U18156 (N_18156,N_17937,N_17858);
xnor U18157 (N_18157,N_17818,N_17892);
nor U18158 (N_18158,N_17884,N_17823);
or U18159 (N_18159,N_17911,N_17992);
nor U18160 (N_18160,N_17833,N_17849);
or U18161 (N_18161,N_17802,N_17905);
or U18162 (N_18162,N_17921,N_17965);
or U18163 (N_18163,N_17827,N_17918);
nor U18164 (N_18164,N_17838,N_17986);
and U18165 (N_18165,N_17868,N_17966);
nor U18166 (N_18166,N_17845,N_17930);
nor U18167 (N_18167,N_17852,N_17830);
nand U18168 (N_18168,N_17836,N_17808);
nand U18169 (N_18169,N_17855,N_17915);
and U18170 (N_18170,N_17954,N_17814);
or U18171 (N_18171,N_17901,N_17932);
nand U18172 (N_18172,N_17990,N_17906);
or U18173 (N_18173,N_17941,N_17826);
nor U18174 (N_18174,N_17851,N_17950);
nand U18175 (N_18175,N_17949,N_17990);
and U18176 (N_18176,N_17985,N_17849);
nand U18177 (N_18177,N_17942,N_17884);
or U18178 (N_18178,N_17962,N_17961);
and U18179 (N_18179,N_17969,N_17963);
nand U18180 (N_18180,N_17864,N_17902);
or U18181 (N_18181,N_17847,N_17818);
nand U18182 (N_18182,N_17853,N_17941);
and U18183 (N_18183,N_17941,N_17918);
nand U18184 (N_18184,N_17870,N_17926);
nand U18185 (N_18185,N_17836,N_17850);
and U18186 (N_18186,N_17811,N_17843);
xor U18187 (N_18187,N_17820,N_17961);
and U18188 (N_18188,N_17973,N_17955);
nand U18189 (N_18189,N_17840,N_17917);
xnor U18190 (N_18190,N_17885,N_17948);
xor U18191 (N_18191,N_17947,N_17868);
nor U18192 (N_18192,N_17905,N_17897);
or U18193 (N_18193,N_17861,N_17887);
nand U18194 (N_18194,N_17918,N_17848);
or U18195 (N_18195,N_17921,N_17907);
nand U18196 (N_18196,N_17913,N_17818);
or U18197 (N_18197,N_17985,N_17838);
or U18198 (N_18198,N_17834,N_17909);
and U18199 (N_18199,N_17973,N_17940);
xor U18200 (N_18200,N_18024,N_18074);
nor U18201 (N_18201,N_18132,N_18197);
nor U18202 (N_18202,N_18118,N_18107);
nor U18203 (N_18203,N_18142,N_18198);
nor U18204 (N_18204,N_18034,N_18177);
and U18205 (N_18205,N_18092,N_18106);
or U18206 (N_18206,N_18027,N_18028);
nor U18207 (N_18207,N_18033,N_18152);
nor U18208 (N_18208,N_18113,N_18014);
and U18209 (N_18209,N_18031,N_18188);
or U18210 (N_18210,N_18063,N_18133);
nor U18211 (N_18211,N_18004,N_18109);
or U18212 (N_18212,N_18174,N_18191);
and U18213 (N_18213,N_18172,N_18017);
and U18214 (N_18214,N_18051,N_18023);
and U18215 (N_18215,N_18052,N_18158);
or U18216 (N_18216,N_18070,N_18002);
nor U18217 (N_18217,N_18125,N_18076);
xnor U18218 (N_18218,N_18093,N_18049);
nand U18219 (N_18219,N_18068,N_18189);
nor U18220 (N_18220,N_18166,N_18053);
nor U18221 (N_18221,N_18140,N_18061);
and U18222 (N_18222,N_18091,N_18194);
and U18223 (N_18223,N_18148,N_18046);
or U18224 (N_18224,N_18193,N_18071);
and U18225 (N_18225,N_18021,N_18134);
xnor U18226 (N_18226,N_18056,N_18089);
or U18227 (N_18227,N_18081,N_18110);
nor U18228 (N_18228,N_18005,N_18072);
nor U18229 (N_18229,N_18102,N_18114);
and U18230 (N_18230,N_18058,N_18159);
nand U18231 (N_18231,N_18149,N_18147);
and U18232 (N_18232,N_18138,N_18196);
and U18233 (N_18233,N_18047,N_18048);
nor U18234 (N_18234,N_18157,N_18123);
nor U18235 (N_18235,N_18131,N_18096);
nor U18236 (N_18236,N_18080,N_18000);
and U18237 (N_18237,N_18181,N_18141);
and U18238 (N_18238,N_18195,N_18120);
and U18239 (N_18239,N_18183,N_18156);
or U18240 (N_18240,N_18184,N_18153);
nand U18241 (N_18241,N_18060,N_18038);
or U18242 (N_18242,N_18016,N_18013);
nor U18243 (N_18243,N_18145,N_18054);
or U18244 (N_18244,N_18026,N_18100);
nand U18245 (N_18245,N_18040,N_18192);
nor U18246 (N_18246,N_18150,N_18055);
or U18247 (N_18247,N_18009,N_18035);
nor U18248 (N_18248,N_18154,N_18059);
or U18249 (N_18249,N_18098,N_18086);
or U18250 (N_18250,N_18042,N_18139);
or U18251 (N_18251,N_18043,N_18122);
nor U18252 (N_18252,N_18128,N_18044);
or U18253 (N_18253,N_18111,N_18176);
xor U18254 (N_18254,N_18030,N_18173);
nor U18255 (N_18255,N_18065,N_18171);
nand U18256 (N_18256,N_18101,N_18105);
or U18257 (N_18257,N_18041,N_18077);
nor U18258 (N_18258,N_18007,N_18025);
nor U18259 (N_18259,N_18087,N_18185);
nand U18260 (N_18260,N_18085,N_18079);
or U18261 (N_18261,N_18160,N_18146);
nor U18262 (N_18262,N_18199,N_18144);
nand U18263 (N_18263,N_18126,N_18083);
or U18264 (N_18264,N_18078,N_18075);
or U18265 (N_18265,N_18036,N_18155);
or U18266 (N_18266,N_18022,N_18066);
or U18267 (N_18267,N_18062,N_18019);
nand U18268 (N_18268,N_18097,N_18015);
xor U18269 (N_18269,N_18137,N_18108);
and U18270 (N_18270,N_18008,N_18127);
nor U18271 (N_18271,N_18069,N_18018);
nand U18272 (N_18272,N_18115,N_18094);
xor U18273 (N_18273,N_18190,N_18020);
nand U18274 (N_18274,N_18012,N_18124);
xor U18275 (N_18275,N_18164,N_18151);
nor U18276 (N_18276,N_18090,N_18057);
and U18277 (N_18277,N_18029,N_18084);
or U18278 (N_18278,N_18129,N_18099);
or U18279 (N_18279,N_18050,N_18135);
or U18280 (N_18280,N_18162,N_18010);
xor U18281 (N_18281,N_18119,N_18169);
nor U18282 (N_18282,N_18167,N_18039);
or U18283 (N_18283,N_18073,N_18186);
and U18284 (N_18284,N_18082,N_18011);
and U18285 (N_18285,N_18095,N_18182);
nand U18286 (N_18286,N_18170,N_18165);
nand U18287 (N_18287,N_18163,N_18006);
and U18288 (N_18288,N_18003,N_18178);
nor U18289 (N_18289,N_18103,N_18130);
xnor U18290 (N_18290,N_18136,N_18117);
or U18291 (N_18291,N_18088,N_18037);
or U18292 (N_18292,N_18187,N_18175);
nor U18293 (N_18293,N_18161,N_18001);
or U18294 (N_18294,N_18064,N_18180);
and U18295 (N_18295,N_18121,N_18104);
nor U18296 (N_18296,N_18045,N_18067);
xor U18297 (N_18297,N_18143,N_18179);
and U18298 (N_18298,N_18168,N_18116);
and U18299 (N_18299,N_18032,N_18112);
xor U18300 (N_18300,N_18162,N_18170);
and U18301 (N_18301,N_18147,N_18023);
and U18302 (N_18302,N_18160,N_18127);
nand U18303 (N_18303,N_18199,N_18135);
and U18304 (N_18304,N_18141,N_18061);
nand U18305 (N_18305,N_18155,N_18095);
xnor U18306 (N_18306,N_18052,N_18165);
and U18307 (N_18307,N_18050,N_18044);
nor U18308 (N_18308,N_18003,N_18110);
and U18309 (N_18309,N_18173,N_18112);
or U18310 (N_18310,N_18173,N_18123);
nor U18311 (N_18311,N_18001,N_18083);
and U18312 (N_18312,N_18017,N_18142);
or U18313 (N_18313,N_18172,N_18028);
and U18314 (N_18314,N_18197,N_18160);
nand U18315 (N_18315,N_18199,N_18189);
and U18316 (N_18316,N_18189,N_18094);
and U18317 (N_18317,N_18056,N_18011);
nand U18318 (N_18318,N_18107,N_18028);
xnor U18319 (N_18319,N_18129,N_18042);
nand U18320 (N_18320,N_18002,N_18054);
or U18321 (N_18321,N_18168,N_18156);
nand U18322 (N_18322,N_18080,N_18146);
nand U18323 (N_18323,N_18161,N_18081);
and U18324 (N_18324,N_18104,N_18164);
xnor U18325 (N_18325,N_18004,N_18195);
or U18326 (N_18326,N_18030,N_18117);
nor U18327 (N_18327,N_18026,N_18191);
or U18328 (N_18328,N_18076,N_18150);
nor U18329 (N_18329,N_18098,N_18006);
nor U18330 (N_18330,N_18181,N_18176);
or U18331 (N_18331,N_18166,N_18068);
nor U18332 (N_18332,N_18181,N_18192);
nor U18333 (N_18333,N_18147,N_18082);
nand U18334 (N_18334,N_18115,N_18185);
nor U18335 (N_18335,N_18095,N_18172);
nand U18336 (N_18336,N_18047,N_18115);
and U18337 (N_18337,N_18164,N_18130);
and U18338 (N_18338,N_18006,N_18161);
nor U18339 (N_18339,N_18167,N_18003);
nand U18340 (N_18340,N_18174,N_18077);
and U18341 (N_18341,N_18169,N_18036);
nand U18342 (N_18342,N_18170,N_18024);
and U18343 (N_18343,N_18161,N_18178);
nand U18344 (N_18344,N_18139,N_18010);
or U18345 (N_18345,N_18087,N_18025);
nand U18346 (N_18346,N_18073,N_18065);
or U18347 (N_18347,N_18047,N_18038);
or U18348 (N_18348,N_18115,N_18086);
or U18349 (N_18349,N_18128,N_18191);
and U18350 (N_18350,N_18157,N_18145);
and U18351 (N_18351,N_18023,N_18079);
or U18352 (N_18352,N_18127,N_18043);
and U18353 (N_18353,N_18039,N_18033);
and U18354 (N_18354,N_18113,N_18138);
and U18355 (N_18355,N_18144,N_18171);
nand U18356 (N_18356,N_18055,N_18028);
nand U18357 (N_18357,N_18128,N_18152);
nor U18358 (N_18358,N_18089,N_18024);
or U18359 (N_18359,N_18169,N_18012);
and U18360 (N_18360,N_18158,N_18033);
nand U18361 (N_18361,N_18063,N_18182);
nand U18362 (N_18362,N_18179,N_18116);
and U18363 (N_18363,N_18150,N_18086);
and U18364 (N_18364,N_18132,N_18176);
nand U18365 (N_18365,N_18008,N_18113);
or U18366 (N_18366,N_18173,N_18010);
or U18367 (N_18367,N_18187,N_18199);
xor U18368 (N_18368,N_18141,N_18011);
and U18369 (N_18369,N_18140,N_18130);
and U18370 (N_18370,N_18003,N_18180);
or U18371 (N_18371,N_18135,N_18120);
and U18372 (N_18372,N_18187,N_18186);
nor U18373 (N_18373,N_18003,N_18045);
nor U18374 (N_18374,N_18187,N_18032);
nor U18375 (N_18375,N_18029,N_18198);
nand U18376 (N_18376,N_18074,N_18055);
nand U18377 (N_18377,N_18071,N_18141);
nand U18378 (N_18378,N_18033,N_18116);
and U18379 (N_18379,N_18166,N_18025);
nand U18380 (N_18380,N_18175,N_18064);
nor U18381 (N_18381,N_18117,N_18097);
and U18382 (N_18382,N_18108,N_18070);
or U18383 (N_18383,N_18183,N_18126);
xnor U18384 (N_18384,N_18199,N_18115);
and U18385 (N_18385,N_18031,N_18038);
nand U18386 (N_18386,N_18037,N_18185);
and U18387 (N_18387,N_18121,N_18035);
nand U18388 (N_18388,N_18057,N_18163);
nand U18389 (N_18389,N_18190,N_18122);
nand U18390 (N_18390,N_18157,N_18094);
xor U18391 (N_18391,N_18018,N_18092);
xnor U18392 (N_18392,N_18139,N_18032);
or U18393 (N_18393,N_18101,N_18023);
xnor U18394 (N_18394,N_18180,N_18043);
nor U18395 (N_18395,N_18053,N_18179);
nand U18396 (N_18396,N_18113,N_18048);
nand U18397 (N_18397,N_18010,N_18136);
nand U18398 (N_18398,N_18197,N_18140);
xnor U18399 (N_18399,N_18007,N_18052);
xnor U18400 (N_18400,N_18294,N_18355);
and U18401 (N_18401,N_18350,N_18363);
and U18402 (N_18402,N_18227,N_18390);
and U18403 (N_18403,N_18348,N_18342);
xor U18404 (N_18404,N_18232,N_18394);
or U18405 (N_18405,N_18284,N_18386);
nand U18406 (N_18406,N_18255,N_18236);
or U18407 (N_18407,N_18203,N_18301);
xor U18408 (N_18408,N_18217,N_18392);
nor U18409 (N_18409,N_18242,N_18366);
or U18410 (N_18410,N_18319,N_18321);
nand U18411 (N_18411,N_18207,N_18211);
nand U18412 (N_18412,N_18323,N_18279);
xnor U18413 (N_18413,N_18273,N_18311);
nor U18414 (N_18414,N_18380,N_18327);
or U18415 (N_18415,N_18317,N_18361);
nand U18416 (N_18416,N_18326,N_18341);
nor U18417 (N_18417,N_18228,N_18346);
and U18418 (N_18418,N_18270,N_18241);
xor U18419 (N_18419,N_18280,N_18286);
nor U18420 (N_18420,N_18237,N_18267);
and U18421 (N_18421,N_18378,N_18303);
nand U18422 (N_18422,N_18365,N_18262);
and U18423 (N_18423,N_18252,N_18291);
nand U18424 (N_18424,N_18292,N_18324);
or U18425 (N_18425,N_18336,N_18297);
nor U18426 (N_18426,N_18261,N_18330);
and U18427 (N_18427,N_18351,N_18360);
or U18428 (N_18428,N_18298,N_18204);
and U18429 (N_18429,N_18274,N_18256);
or U18430 (N_18430,N_18266,N_18353);
or U18431 (N_18431,N_18331,N_18362);
nand U18432 (N_18432,N_18314,N_18375);
and U18433 (N_18433,N_18238,N_18325);
and U18434 (N_18434,N_18308,N_18293);
nand U18435 (N_18435,N_18215,N_18397);
xnor U18436 (N_18436,N_18288,N_18368);
nor U18437 (N_18437,N_18285,N_18304);
nand U18438 (N_18438,N_18334,N_18318);
nor U18439 (N_18439,N_18202,N_18258);
or U18440 (N_18440,N_18271,N_18328);
or U18441 (N_18441,N_18214,N_18276);
or U18442 (N_18442,N_18302,N_18359);
nand U18443 (N_18443,N_18264,N_18315);
nor U18444 (N_18444,N_18344,N_18277);
and U18445 (N_18445,N_18372,N_18339);
or U18446 (N_18446,N_18384,N_18282);
nor U18447 (N_18447,N_18235,N_18260);
and U18448 (N_18448,N_18212,N_18295);
and U18449 (N_18449,N_18349,N_18310);
or U18450 (N_18450,N_18379,N_18387);
xnor U18451 (N_18451,N_18254,N_18358);
and U18452 (N_18452,N_18305,N_18381);
and U18453 (N_18453,N_18206,N_18231);
nor U18454 (N_18454,N_18354,N_18389);
or U18455 (N_18455,N_18220,N_18347);
nand U18456 (N_18456,N_18352,N_18225);
and U18457 (N_18457,N_18287,N_18257);
or U18458 (N_18458,N_18399,N_18364);
or U18459 (N_18459,N_18223,N_18306);
and U18460 (N_18460,N_18219,N_18320);
nand U18461 (N_18461,N_18356,N_18251);
nand U18462 (N_18462,N_18249,N_18200);
nand U18463 (N_18463,N_18289,N_18296);
xor U18464 (N_18464,N_18313,N_18391);
nand U18465 (N_18465,N_18322,N_18385);
nor U18466 (N_18466,N_18393,N_18374);
nor U18467 (N_18467,N_18234,N_18395);
nand U18468 (N_18468,N_18244,N_18201);
nand U18469 (N_18469,N_18224,N_18367);
and U18470 (N_18470,N_18309,N_18343);
xor U18471 (N_18471,N_18222,N_18335);
and U18472 (N_18472,N_18272,N_18259);
nand U18473 (N_18473,N_18248,N_18253);
nand U18474 (N_18474,N_18316,N_18369);
or U18475 (N_18475,N_18218,N_18240);
and U18476 (N_18476,N_18268,N_18245);
xor U18477 (N_18477,N_18265,N_18329);
and U18478 (N_18478,N_18208,N_18210);
or U18479 (N_18479,N_18383,N_18373);
and U18480 (N_18480,N_18345,N_18281);
or U18481 (N_18481,N_18398,N_18230);
or U18482 (N_18482,N_18290,N_18396);
or U18483 (N_18483,N_18209,N_18246);
and U18484 (N_18484,N_18205,N_18307);
and U18485 (N_18485,N_18338,N_18377);
nand U18486 (N_18486,N_18239,N_18250);
nor U18487 (N_18487,N_18333,N_18263);
or U18488 (N_18488,N_18213,N_18216);
nand U18489 (N_18489,N_18332,N_18376);
nand U18490 (N_18490,N_18278,N_18221);
xor U18491 (N_18491,N_18388,N_18269);
or U18492 (N_18492,N_18243,N_18300);
nor U18493 (N_18493,N_18299,N_18247);
nor U18494 (N_18494,N_18312,N_18382);
and U18495 (N_18495,N_18371,N_18370);
or U18496 (N_18496,N_18337,N_18283);
and U18497 (N_18497,N_18233,N_18275);
or U18498 (N_18498,N_18340,N_18229);
or U18499 (N_18499,N_18357,N_18226);
or U18500 (N_18500,N_18347,N_18253);
nand U18501 (N_18501,N_18320,N_18340);
nor U18502 (N_18502,N_18346,N_18375);
nand U18503 (N_18503,N_18261,N_18365);
xnor U18504 (N_18504,N_18386,N_18397);
and U18505 (N_18505,N_18399,N_18390);
and U18506 (N_18506,N_18382,N_18240);
and U18507 (N_18507,N_18386,N_18304);
and U18508 (N_18508,N_18325,N_18247);
and U18509 (N_18509,N_18333,N_18288);
and U18510 (N_18510,N_18373,N_18323);
or U18511 (N_18511,N_18349,N_18278);
xnor U18512 (N_18512,N_18216,N_18220);
xnor U18513 (N_18513,N_18374,N_18388);
or U18514 (N_18514,N_18299,N_18365);
or U18515 (N_18515,N_18312,N_18347);
nor U18516 (N_18516,N_18229,N_18357);
or U18517 (N_18517,N_18295,N_18379);
nor U18518 (N_18518,N_18348,N_18299);
or U18519 (N_18519,N_18289,N_18379);
or U18520 (N_18520,N_18362,N_18340);
and U18521 (N_18521,N_18386,N_18260);
nand U18522 (N_18522,N_18266,N_18397);
xnor U18523 (N_18523,N_18208,N_18370);
nor U18524 (N_18524,N_18258,N_18255);
and U18525 (N_18525,N_18391,N_18258);
nor U18526 (N_18526,N_18261,N_18296);
and U18527 (N_18527,N_18232,N_18230);
nor U18528 (N_18528,N_18249,N_18240);
and U18529 (N_18529,N_18289,N_18250);
or U18530 (N_18530,N_18224,N_18230);
and U18531 (N_18531,N_18372,N_18393);
or U18532 (N_18532,N_18377,N_18386);
nor U18533 (N_18533,N_18330,N_18393);
and U18534 (N_18534,N_18205,N_18282);
and U18535 (N_18535,N_18304,N_18292);
or U18536 (N_18536,N_18308,N_18239);
and U18537 (N_18537,N_18298,N_18259);
nor U18538 (N_18538,N_18230,N_18298);
and U18539 (N_18539,N_18342,N_18379);
nand U18540 (N_18540,N_18216,N_18354);
and U18541 (N_18541,N_18242,N_18396);
and U18542 (N_18542,N_18264,N_18306);
xor U18543 (N_18543,N_18211,N_18387);
nand U18544 (N_18544,N_18279,N_18312);
nor U18545 (N_18545,N_18345,N_18291);
nand U18546 (N_18546,N_18238,N_18297);
xnor U18547 (N_18547,N_18392,N_18395);
and U18548 (N_18548,N_18325,N_18313);
xnor U18549 (N_18549,N_18212,N_18371);
nor U18550 (N_18550,N_18347,N_18316);
nor U18551 (N_18551,N_18319,N_18261);
nor U18552 (N_18552,N_18238,N_18383);
and U18553 (N_18553,N_18274,N_18293);
or U18554 (N_18554,N_18323,N_18229);
and U18555 (N_18555,N_18281,N_18202);
nor U18556 (N_18556,N_18398,N_18251);
nand U18557 (N_18557,N_18381,N_18242);
nand U18558 (N_18558,N_18344,N_18291);
xor U18559 (N_18559,N_18219,N_18339);
nor U18560 (N_18560,N_18304,N_18322);
or U18561 (N_18561,N_18211,N_18309);
nor U18562 (N_18562,N_18242,N_18213);
nor U18563 (N_18563,N_18396,N_18276);
xnor U18564 (N_18564,N_18398,N_18212);
and U18565 (N_18565,N_18274,N_18325);
xor U18566 (N_18566,N_18395,N_18360);
or U18567 (N_18567,N_18298,N_18389);
nand U18568 (N_18568,N_18322,N_18387);
xnor U18569 (N_18569,N_18274,N_18310);
nand U18570 (N_18570,N_18213,N_18315);
and U18571 (N_18571,N_18307,N_18247);
nand U18572 (N_18572,N_18241,N_18396);
nand U18573 (N_18573,N_18244,N_18203);
nand U18574 (N_18574,N_18386,N_18259);
or U18575 (N_18575,N_18358,N_18250);
and U18576 (N_18576,N_18246,N_18380);
and U18577 (N_18577,N_18375,N_18210);
or U18578 (N_18578,N_18202,N_18314);
and U18579 (N_18579,N_18302,N_18326);
nor U18580 (N_18580,N_18298,N_18272);
nor U18581 (N_18581,N_18214,N_18393);
nor U18582 (N_18582,N_18207,N_18367);
nor U18583 (N_18583,N_18353,N_18316);
nand U18584 (N_18584,N_18393,N_18287);
or U18585 (N_18585,N_18246,N_18357);
xor U18586 (N_18586,N_18245,N_18213);
xnor U18587 (N_18587,N_18222,N_18368);
and U18588 (N_18588,N_18261,N_18241);
nand U18589 (N_18589,N_18264,N_18294);
and U18590 (N_18590,N_18331,N_18239);
and U18591 (N_18591,N_18301,N_18318);
or U18592 (N_18592,N_18268,N_18251);
nor U18593 (N_18593,N_18243,N_18377);
xnor U18594 (N_18594,N_18215,N_18250);
or U18595 (N_18595,N_18347,N_18368);
or U18596 (N_18596,N_18218,N_18251);
nand U18597 (N_18597,N_18291,N_18336);
and U18598 (N_18598,N_18258,N_18378);
nand U18599 (N_18599,N_18328,N_18296);
and U18600 (N_18600,N_18499,N_18409);
and U18601 (N_18601,N_18428,N_18537);
or U18602 (N_18602,N_18495,N_18400);
or U18603 (N_18603,N_18417,N_18547);
xor U18604 (N_18604,N_18559,N_18434);
or U18605 (N_18605,N_18440,N_18454);
nor U18606 (N_18606,N_18572,N_18493);
nand U18607 (N_18607,N_18561,N_18595);
nand U18608 (N_18608,N_18574,N_18597);
xor U18609 (N_18609,N_18411,N_18462);
nand U18610 (N_18610,N_18510,N_18532);
and U18611 (N_18611,N_18433,N_18435);
nor U18612 (N_18612,N_18451,N_18422);
nand U18613 (N_18613,N_18550,N_18589);
nor U18614 (N_18614,N_18580,N_18503);
or U18615 (N_18615,N_18587,N_18447);
and U18616 (N_18616,N_18402,N_18483);
and U18617 (N_18617,N_18401,N_18449);
nor U18618 (N_18618,N_18517,N_18519);
or U18619 (N_18619,N_18575,N_18554);
nor U18620 (N_18620,N_18484,N_18430);
or U18621 (N_18621,N_18522,N_18592);
or U18622 (N_18622,N_18505,N_18596);
and U18623 (N_18623,N_18413,N_18556);
nand U18624 (N_18624,N_18583,N_18406);
or U18625 (N_18625,N_18553,N_18540);
or U18626 (N_18626,N_18541,N_18506);
xor U18627 (N_18627,N_18481,N_18427);
xor U18628 (N_18628,N_18560,N_18557);
nor U18629 (N_18629,N_18446,N_18585);
nor U18630 (N_18630,N_18460,N_18415);
xor U18631 (N_18631,N_18423,N_18542);
nor U18632 (N_18632,N_18485,N_18593);
xnor U18633 (N_18633,N_18512,N_18591);
nor U18634 (N_18634,N_18568,N_18544);
xnor U18635 (N_18635,N_18420,N_18562);
nor U18636 (N_18636,N_18476,N_18528);
nor U18637 (N_18637,N_18576,N_18477);
xnor U18638 (N_18638,N_18453,N_18436);
or U18639 (N_18639,N_18588,N_18577);
or U18640 (N_18640,N_18416,N_18457);
and U18641 (N_18641,N_18598,N_18501);
nand U18642 (N_18642,N_18509,N_18590);
xnor U18643 (N_18643,N_18530,N_18514);
nand U18644 (N_18644,N_18408,N_18511);
and U18645 (N_18645,N_18478,N_18450);
nor U18646 (N_18646,N_18502,N_18431);
nand U18647 (N_18647,N_18570,N_18452);
nand U18648 (N_18648,N_18581,N_18468);
xor U18649 (N_18649,N_18520,N_18521);
or U18650 (N_18650,N_18407,N_18443);
nand U18651 (N_18651,N_18491,N_18578);
xnor U18652 (N_18652,N_18444,N_18529);
and U18653 (N_18653,N_18490,N_18421);
or U18654 (N_18654,N_18459,N_18463);
or U18655 (N_18655,N_18599,N_18455);
nor U18656 (N_18656,N_18563,N_18497);
xor U18657 (N_18657,N_18412,N_18573);
or U18658 (N_18658,N_18404,N_18492);
nor U18659 (N_18659,N_18475,N_18565);
or U18660 (N_18660,N_18548,N_18448);
nand U18661 (N_18661,N_18479,N_18486);
nor U18662 (N_18662,N_18425,N_18546);
xnor U18663 (N_18663,N_18571,N_18579);
and U18664 (N_18664,N_18545,N_18441);
or U18665 (N_18665,N_18539,N_18508);
or U18666 (N_18666,N_18586,N_18555);
and U18667 (N_18667,N_18531,N_18584);
and U18668 (N_18668,N_18496,N_18552);
and U18669 (N_18669,N_18480,N_18487);
and U18670 (N_18670,N_18549,N_18467);
or U18671 (N_18671,N_18465,N_18518);
or U18672 (N_18672,N_18474,N_18515);
and U18673 (N_18673,N_18533,N_18405);
nor U18674 (N_18674,N_18471,N_18524);
or U18675 (N_18675,N_18567,N_18456);
or U18676 (N_18676,N_18472,N_18458);
and U18677 (N_18677,N_18498,N_18536);
or U18678 (N_18678,N_18469,N_18418);
or U18679 (N_18679,N_18523,N_18403);
or U18680 (N_18680,N_18566,N_18569);
nand U18681 (N_18681,N_18525,N_18543);
xnor U18682 (N_18682,N_18489,N_18527);
or U18683 (N_18683,N_18414,N_18538);
or U18684 (N_18684,N_18564,N_18558);
nor U18685 (N_18685,N_18470,N_18594);
and U18686 (N_18686,N_18513,N_18488);
nand U18687 (N_18687,N_18507,N_18445);
nor U18688 (N_18688,N_18504,N_18438);
nand U18689 (N_18689,N_18494,N_18410);
nand U18690 (N_18690,N_18534,N_18464);
nand U18691 (N_18691,N_18473,N_18516);
nor U18692 (N_18692,N_18419,N_18526);
or U18693 (N_18693,N_18437,N_18442);
nor U18694 (N_18694,N_18429,N_18424);
nor U18695 (N_18695,N_18500,N_18426);
or U18696 (N_18696,N_18461,N_18551);
and U18697 (N_18697,N_18432,N_18439);
nor U18698 (N_18698,N_18482,N_18582);
and U18699 (N_18699,N_18535,N_18466);
nand U18700 (N_18700,N_18489,N_18424);
xnor U18701 (N_18701,N_18501,N_18482);
nand U18702 (N_18702,N_18413,N_18572);
and U18703 (N_18703,N_18589,N_18419);
nor U18704 (N_18704,N_18541,N_18452);
nor U18705 (N_18705,N_18484,N_18478);
nor U18706 (N_18706,N_18493,N_18561);
or U18707 (N_18707,N_18467,N_18428);
and U18708 (N_18708,N_18477,N_18580);
xnor U18709 (N_18709,N_18454,N_18495);
xor U18710 (N_18710,N_18431,N_18504);
and U18711 (N_18711,N_18527,N_18434);
xnor U18712 (N_18712,N_18473,N_18446);
nor U18713 (N_18713,N_18428,N_18576);
and U18714 (N_18714,N_18518,N_18503);
nand U18715 (N_18715,N_18487,N_18461);
and U18716 (N_18716,N_18504,N_18422);
xnor U18717 (N_18717,N_18482,N_18491);
nor U18718 (N_18718,N_18488,N_18443);
nor U18719 (N_18719,N_18488,N_18567);
and U18720 (N_18720,N_18522,N_18420);
and U18721 (N_18721,N_18443,N_18427);
nand U18722 (N_18722,N_18507,N_18518);
nand U18723 (N_18723,N_18404,N_18493);
xor U18724 (N_18724,N_18511,N_18451);
and U18725 (N_18725,N_18426,N_18404);
xnor U18726 (N_18726,N_18555,N_18553);
or U18727 (N_18727,N_18468,N_18515);
or U18728 (N_18728,N_18424,N_18450);
or U18729 (N_18729,N_18525,N_18439);
and U18730 (N_18730,N_18496,N_18586);
nand U18731 (N_18731,N_18430,N_18569);
and U18732 (N_18732,N_18439,N_18426);
nor U18733 (N_18733,N_18427,N_18534);
and U18734 (N_18734,N_18516,N_18415);
nor U18735 (N_18735,N_18500,N_18563);
and U18736 (N_18736,N_18580,N_18589);
nand U18737 (N_18737,N_18593,N_18477);
and U18738 (N_18738,N_18472,N_18437);
and U18739 (N_18739,N_18507,N_18597);
nand U18740 (N_18740,N_18545,N_18450);
nand U18741 (N_18741,N_18427,N_18429);
nor U18742 (N_18742,N_18520,N_18462);
nand U18743 (N_18743,N_18558,N_18426);
nand U18744 (N_18744,N_18446,N_18581);
or U18745 (N_18745,N_18402,N_18508);
xor U18746 (N_18746,N_18566,N_18588);
nor U18747 (N_18747,N_18557,N_18574);
or U18748 (N_18748,N_18453,N_18425);
and U18749 (N_18749,N_18555,N_18412);
or U18750 (N_18750,N_18416,N_18492);
or U18751 (N_18751,N_18470,N_18518);
or U18752 (N_18752,N_18506,N_18562);
or U18753 (N_18753,N_18422,N_18460);
nand U18754 (N_18754,N_18429,N_18415);
or U18755 (N_18755,N_18510,N_18593);
and U18756 (N_18756,N_18494,N_18521);
xnor U18757 (N_18757,N_18555,N_18576);
nor U18758 (N_18758,N_18557,N_18417);
xor U18759 (N_18759,N_18487,N_18592);
and U18760 (N_18760,N_18568,N_18421);
xor U18761 (N_18761,N_18495,N_18448);
or U18762 (N_18762,N_18407,N_18456);
nand U18763 (N_18763,N_18410,N_18548);
and U18764 (N_18764,N_18563,N_18599);
xnor U18765 (N_18765,N_18435,N_18509);
and U18766 (N_18766,N_18500,N_18504);
and U18767 (N_18767,N_18486,N_18585);
or U18768 (N_18768,N_18587,N_18592);
and U18769 (N_18769,N_18517,N_18538);
or U18770 (N_18770,N_18585,N_18534);
nand U18771 (N_18771,N_18435,N_18476);
nand U18772 (N_18772,N_18463,N_18464);
nor U18773 (N_18773,N_18547,N_18462);
and U18774 (N_18774,N_18462,N_18534);
nor U18775 (N_18775,N_18440,N_18469);
and U18776 (N_18776,N_18480,N_18551);
or U18777 (N_18777,N_18476,N_18427);
nand U18778 (N_18778,N_18475,N_18574);
and U18779 (N_18779,N_18498,N_18488);
nand U18780 (N_18780,N_18470,N_18575);
and U18781 (N_18781,N_18422,N_18438);
nor U18782 (N_18782,N_18412,N_18512);
nor U18783 (N_18783,N_18581,N_18571);
nor U18784 (N_18784,N_18414,N_18533);
nor U18785 (N_18785,N_18542,N_18535);
nand U18786 (N_18786,N_18453,N_18445);
nand U18787 (N_18787,N_18448,N_18457);
nor U18788 (N_18788,N_18487,N_18482);
nand U18789 (N_18789,N_18407,N_18562);
and U18790 (N_18790,N_18408,N_18500);
nor U18791 (N_18791,N_18486,N_18436);
nor U18792 (N_18792,N_18461,N_18592);
or U18793 (N_18793,N_18459,N_18583);
nand U18794 (N_18794,N_18464,N_18512);
nand U18795 (N_18795,N_18541,N_18464);
nor U18796 (N_18796,N_18542,N_18505);
nor U18797 (N_18797,N_18421,N_18450);
and U18798 (N_18798,N_18411,N_18433);
nor U18799 (N_18799,N_18411,N_18421);
or U18800 (N_18800,N_18640,N_18669);
nor U18801 (N_18801,N_18681,N_18623);
nor U18802 (N_18802,N_18695,N_18682);
or U18803 (N_18803,N_18724,N_18707);
or U18804 (N_18804,N_18648,N_18641);
nand U18805 (N_18805,N_18668,N_18601);
nor U18806 (N_18806,N_18606,N_18782);
or U18807 (N_18807,N_18610,N_18658);
and U18808 (N_18808,N_18717,N_18638);
nand U18809 (N_18809,N_18696,N_18665);
nor U18810 (N_18810,N_18715,N_18798);
and U18811 (N_18811,N_18667,N_18657);
nand U18812 (N_18812,N_18746,N_18709);
nor U18813 (N_18813,N_18636,N_18646);
xnor U18814 (N_18814,N_18611,N_18618);
nand U18815 (N_18815,N_18689,N_18757);
xnor U18816 (N_18816,N_18754,N_18692);
and U18817 (N_18817,N_18720,N_18699);
nor U18818 (N_18818,N_18738,N_18745);
xor U18819 (N_18819,N_18781,N_18680);
nand U18820 (N_18820,N_18613,N_18622);
nor U18821 (N_18821,N_18786,N_18647);
nor U18822 (N_18822,N_18656,N_18714);
or U18823 (N_18823,N_18766,N_18734);
nor U18824 (N_18824,N_18752,N_18755);
xor U18825 (N_18825,N_18674,N_18629);
and U18826 (N_18826,N_18687,N_18708);
or U18827 (N_18827,N_18609,N_18780);
or U18828 (N_18828,N_18761,N_18719);
nor U18829 (N_18829,N_18607,N_18770);
nand U18830 (N_18830,N_18747,N_18653);
nor U18831 (N_18831,N_18730,N_18704);
nand U18832 (N_18832,N_18790,N_18765);
nor U18833 (N_18833,N_18671,N_18652);
nand U18834 (N_18834,N_18779,N_18711);
xor U18835 (N_18835,N_18672,N_18750);
and U18836 (N_18836,N_18663,N_18799);
nand U18837 (N_18837,N_18688,N_18694);
or U18838 (N_18838,N_18649,N_18710);
nand U18839 (N_18839,N_18661,N_18650);
and U18840 (N_18840,N_18624,N_18604);
and U18841 (N_18841,N_18679,N_18660);
nand U18842 (N_18842,N_18716,N_18791);
and U18843 (N_18843,N_18787,N_18732);
or U18844 (N_18844,N_18617,N_18795);
nor U18845 (N_18845,N_18683,N_18666);
nor U18846 (N_18846,N_18684,N_18677);
nor U18847 (N_18847,N_18758,N_18691);
nand U18848 (N_18848,N_18794,N_18740);
or U18849 (N_18849,N_18741,N_18764);
xnor U18850 (N_18850,N_18792,N_18620);
xor U18851 (N_18851,N_18615,N_18706);
and U18852 (N_18852,N_18759,N_18775);
nand U18853 (N_18853,N_18701,N_18612);
nand U18854 (N_18854,N_18793,N_18602);
or U18855 (N_18855,N_18614,N_18702);
or U18856 (N_18856,N_18722,N_18703);
and U18857 (N_18857,N_18651,N_18739);
nor U18858 (N_18858,N_18769,N_18645);
nand U18859 (N_18859,N_18644,N_18797);
or U18860 (N_18860,N_18630,N_18789);
or U18861 (N_18861,N_18603,N_18698);
xor U18862 (N_18862,N_18774,N_18628);
or U18863 (N_18863,N_18718,N_18662);
nor U18864 (N_18864,N_18664,N_18639);
nand U18865 (N_18865,N_18736,N_18678);
nor U18866 (N_18866,N_18631,N_18642);
or U18867 (N_18867,N_18728,N_18686);
nand U18868 (N_18868,N_18778,N_18743);
nand U18869 (N_18869,N_18748,N_18670);
or U18870 (N_18870,N_18725,N_18762);
nor U18871 (N_18871,N_18676,N_18605);
nor U18872 (N_18872,N_18675,N_18627);
xnor U18873 (N_18873,N_18723,N_18690);
and U18874 (N_18874,N_18771,N_18749);
nor U18875 (N_18875,N_18608,N_18685);
nand U18876 (N_18876,N_18626,N_18643);
nand U18877 (N_18877,N_18776,N_18700);
and U18878 (N_18878,N_18616,N_18735);
nand U18879 (N_18879,N_18777,N_18773);
nor U18880 (N_18880,N_18729,N_18659);
or U18881 (N_18881,N_18753,N_18768);
nand U18882 (N_18882,N_18756,N_18760);
nand U18883 (N_18883,N_18655,N_18654);
nor U18884 (N_18884,N_18744,N_18772);
and U18885 (N_18885,N_18600,N_18697);
or U18886 (N_18886,N_18705,N_18712);
nor U18887 (N_18887,N_18784,N_18634);
nor U18888 (N_18888,N_18632,N_18733);
or U18889 (N_18889,N_18721,N_18625);
nand U18890 (N_18890,N_18727,N_18763);
and U18891 (N_18891,N_18742,N_18619);
nor U18892 (N_18892,N_18783,N_18693);
and U18893 (N_18893,N_18726,N_18796);
or U18894 (N_18894,N_18635,N_18751);
nand U18895 (N_18895,N_18731,N_18637);
and U18896 (N_18896,N_18785,N_18737);
and U18897 (N_18897,N_18713,N_18767);
or U18898 (N_18898,N_18633,N_18673);
or U18899 (N_18899,N_18621,N_18788);
nand U18900 (N_18900,N_18684,N_18742);
and U18901 (N_18901,N_18663,N_18746);
nand U18902 (N_18902,N_18775,N_18649);
and U18903 (N_18903,N_18642,N_18606);
or U18904 (N_18904,N_18693,N_18604);
nand U18905 (N_18905,N_18644,N_18710);
or U18906 (N_18906,N_18628,N_18785);
or U18907 (N_18907,N_18692,N_18730);
and U18908 (N_18908,N_18783,N_18695);
nand U18909 (N_18909,N_18734,N_18668);
or U18910 (N_18910,N_18761,N_18670);
nand U18911 (N_18911,N_18760,N_18641);
nand U18912 (N_18912,N_18661,N_18693);
nand U18913 (N_18913,N_18711,N_18790);
xor U18914 (N_18914,N_18766,N_18694);
nor U18915 (N_18915,N_18785,N_18795);
nand U18916 (N_18916,N_18702,N_18639);
nand U18917 (N_18917,N_18656,N_18621);
nor U18918 (N_18918,N_18798,N_18730);
nand U18919 (N_18919,N_18791,N_18703);
or U18920 (N_18920,N_18756,N_18646);
nor U18921 (N_18921,N_18748,N_18753);
and U18922 (N_18922,N_18612,N_18601);
xor U18923 (N_18923,N_18649,N_18698);
nor U18924 (N_18924,N_18771,N_18606);
nor U18925 (N_18925,N_18635,N_18700);
nand U18926 (N_18926,N_18610,N_18770);
or U18927 (N_18927,N_18665,N_18729);
or U18928 (N_18928,N_18648,N_18646);
xor U18929 (N_18929,N_18773,N_18656);
nor U18930 (N_18930,N_18796,N_18620);
nand U18931 (N_18931,N_18699,N_18714);
or U18932 (N_18932,N_18701,N_18696);
nor U18933 (N_18933,N_18661,N_18624);
nor U18934 (N_18934,N_18653,N_18656);
or U18935 (N_18935,N_18616,N_18751);
nor U18936 (N_18936,N_18782,N_18728);
or U18937 (N_18937,N_18727,N_18667);
nand U18938 (N_18938,N_18602,N_18630);
nand U18939 (N_18939,N_18740,N_18610);
nand U18940 (N_18940,N_18739,N_18646);
or U18941 (N_18941,N_18613,N_18736);
or U18942 (N_18942,N_18711,N_18774);
and U18943 (N_18943,N_18691,N_18618);
and U18944 (N_18944,N_18798,N_18698);
xor U18945 (N_18945,N_18601,N_18780);
or U18946 (N_18946,N_18662,N_18630);
and U18947 (N_18947,N_18724,N_18622);
nand U18948 (N_18948,N_18610,N_18735);
xnor U18949 (N_18949,N_18757,N_18629);
or U18950 (N_18950,N_18683,N_18625);
nor U18951 (N_18951,N_18686,N_18630);
xnor U18952 (N_18952,N_18779,N_18712);
nand U18953 (N_18953,N_18770,N_18698);
or U18954 (N_18954,N_18714,N_18784);
nor U18955 (N_18955,N_18693,N_18744);
nor U18956 (N_18956,N_18686,N_18793);
nor U18957 (N_18957,N_18693,N_18780);
and U18958 (N_18958,N_18774,N_18652);
nor U18959 (N_18959,N_18676,N_18673);
xor U18960 (N_18960,N_18669,N_18619);
or U18961 (N_18961,N_18769,N_18675);
and U18962 (N_18962,N_18696,N_18626);
or U18963 (N_18963,N_18623,N_18647);
nand U18964 (N_18964,N_18649,N_18749);
nand U18965 (N_18965,N_18767,N_18727);
and U18966 (N_18966,N_18627,N_18679);
nor U18967 (N_18967,N_18740,N_18765);
xnor U18968 (N_18968,N_18757,N_18703);
nor U18969 (N_18969,N_18788,N_18695);
or U18970 (N_18970,N_18765,N_18608);
nand U18971 (N_18971,N_18782,N_18613);
nor U18972 (N_18972,N_18684,N_18662);
or U18973 (N_18973,N_18695,N_18781);
nor U18974 (N_18974,N_18677,N_18617);
and U18975 (N_18975,N_18740,N_18783);
nand U18976 (N_18976,N_18604,N_18750);
xor U18977 (N_18977,N_18688,N_18771);
or U18978 (N_18978,N_18728,N_18760);
xor U18979 (N_18979,N_18781,N_18666);
nand U18980 (N_18980,N_18703,N_18620);
xor U18981 (N_18981,N_18797,N_18773);
nor U18982 (N_18982,N_18738,N_18683);
and U18983 (N_18983,N_18646,N_18634);
nor U18984 (N_18984,N_18780,N_18680);
nor U18985 (N_18985,N_18602,N_18740);
xnor U18986 (N_18986,N_18756,N_18610);
and U18987 (N_18987,N_18733,N_18691);
nand U18988 (N_18988,N_18635,N_18723);
xnor U18989 (N_18989,N_18717,N_18669);
nor U18990 (N_18990,N_18788,N_18647);
and U18991 (N_18991,N_18660,N_18779);
nand U18992 (N_18992,N_18647,N_18760);
or U18993 (N_18993,N_18626,N_18629);
nand U18994 (N_18994,N_18609,N_18662);
nand U18995 (N_18995,N_18762,N_18754);
or U18996 (N_18996,N_18768,N_18662);
nor U18997 (N_18997,N_18749,N_18763);
and U18998 (N_18998,N_18664,N_18776);
xor U18999 (N_18999,N_18786,N_18743);
nor U19000 (N_19000,N_18861,N_18878);
nor U19001 (N_19001,N_18966,N_18994);
nand U19002 (N_19002,N_18937,N_18823);
xor U19003 (N_19003,N_18940,N_18986);
and U19004 (N_19004,N_18929,N_18913);
xnor U19005 (N_19005,N_18997,N_18809);
and U19006 (N_19006,N_18962,N_18876);
or U19007 (N_19007,N_18891,N_18895);
or U19008 (N_19008,N_18867,N_18934);
nand U19009 (N_19009,N_18993,N_18910);
and U19010 (N_19010,N_18965,N_18859);
and U19011 (N_19011,N_18970,N_18889);
nor U19012 (N_19012,N_18902,N_18810);
nor U19013 (N_19013,N_18816,N_18874);
xor U19014 (N_19014,N_18989,N_18808);
xnor U19015 (N_19015,N_18953,N_18905);
or U19016 (N_19016,N_18836,N_18857);
nand U19017 (N_19017,N_18872,N_18945);
xor U19018 (N_19018,N_18866,N_18975);
nand U19019 (N_19019,N_18916,N_18885);
nor U19020 (N_19020,N_18906,N_18964);
nand U19021 (N_19021,N_18958,N_18898);
nand U19022 (N_19022,N_18921,N_18842);
xor U19023 (N_19023,N_18848,N_18979);
or U19024 (N_19024,N_18930,N_18985);
nor U19025 (N_19025,N_18984,N_18835);
nor U19026 (N_19026,N_18936,N_18896);
or U19027 (N_19027,N_18923,N_18963);
nor U19028 (N_19028,N_18819,N_18814);
nand U19029 (N_19029,N_18884,N_18893);
and U19030 (N_19030,N_18933,N_18988);
or U19031 (N_19031,N_18822,N_18900);
xor U19032 (N_19032,N_18862,N_18943);
or U19033 (N_19033,N_18915,N_18955);
and U19034 (N_19034,N_18846,N_18883);
or U19035 (N_19035,N_18879,N_18804);
nand U19036 (N_19036,N_18826,N_18897);
nand U19037 (N_19037,N_18805,N_18991);
or U19038 (N_19038,N_18870,N_18865);
xor U19039 (N_19039,N_18841,N_18815);
nand U19040 (N_19040,N_18869,N_18852);
nor U19041 (N_19041,N_18925,N_18947);
or U19042 (N_19042,N_18961,N_18967);
or U19043 (N_19043,N_18853,N_18840);
nor U19044 (N_19044,N_18802,N_18946);
nand U19045 (N_19045,N_18959,N_18871);
and U19046 (N_19046,N_18854,N_18911);
and U19047 (N_19047,N_18969,N_18942);
nor U19048 (N_19048,N_18980,N_18833);
and U19049 (N_19049,N_18952,N_18939);
nand U19050 (N_19050,N_18981,N_18950);
nand U19051 (N_19051,N_18894,N_18818);
nand U19052 (N_19052,N_18830,N_18817);
nor U19053 (N_19053,N_18998,N_18813);
or U19054 (N_19054,N_18899,N_18935);
nor U19055 (N_19055,N_18888,N_18907);
nand U19056 (N_19056,N_18931,N_18954);
and U19057 (N_19057,N_18995,N_18996);
or U19058 (N_19058,N_18838,N_18827);
nor U19059 (N_19059,N_18886,N_18803);
nand U19060 (N_19060,N_18858,N_18957);
and U19061 (N_19061,N_18892,N_18992);
nor U19062 (N_19062,N_18978,N_18917);
and U19063 (N_19063,N_18927,N_18831);
nand U19064 (N_19064,N_18976,N_18825);
nand U19065 (N_19065,N_18999,N_18877);
nor U19066 (N_19066,N_18922,N_18977);
or U19067 (N_19067,N_18800,N_18956);
or U19068 (N_19068,N_18828,N_18924);
nor U19069 (N_19069,N_18856,N_18812);
or U19070 (N_19070,N_18882,N_18839);
nand U19071 (N_19071,N_18941,N_18837);
and U19072 (N_19072,N_18972,N_18960);
nand U19073 (N_19073,N_18843,N_18909);
nor U19074 (N_19074,N_18845,N_18887);
nand U19075 (N_19075,N_18864,N_18912);
and U19076 (N_19076,N_18851,N_18982);
nand U19077 (N_19077,N_18949,N_18971);
xnor U19078 (N_19078,N_18820,N_18920);
and U19079 (N_19079,N_18926,N_18983);
or U19080 (N_19080,N_18844,N_18928);
and U19081 (N_19081,N_18855,N_18821);
nor U19082 (N_19082,N_18832,N_18807);
or U19083 (N_19083,N_18968,N_18987);
nand U19084 (N_19084,N_18901,N_18873);
nor U19085 (N_19085,N_18806,N_18875);
nand U19086 (N_19086,N_18824,N_18863);
nor U19087 (N_19087,N_18918,N_18801);
xnor U19088 (N_19088,N_18860,N_18880);
and U19089 (N_19089,N_18890,N_18948);
nand U19090 (N_19090,N_18908,N_18974);
nand U19091 (N_19091,N_18850,N_18829);
nor U19092 (N_19092,N_18914,N_18868);
nor U19093 (N_19093,N_18834,N_18990);
xor U19094 (N_19094,N_18973,N_18919);
nand U19095 (N_19095,N_18904,N_18849);
nor U19096 (N_19096,N_18938,N_18944);
or U19097 (N_19097,N_18811,N_18951);
nand U19098 (N_19098,N_18932,N_18881);
nand U19099 (N_19099,N_18847,N_18903);
and U19100 (N_19100,N_18870,N_18840);
nand U19101 (N_19101,N_18955,N_18977);
or U19102 (N_19102,N_18969,N_18876);
nor U19103 (N_19103,N_18949,N_18945);
nor U19104 (N_19104,N_18800,N_18859);
xnor U19105 (N_19105,N_18937,N_18940);
nand U19106 (N_19106,N_18846,N_18939);
xnor U19107 (N_19107,N_18884,N_18875);
nand U19108 (N_19108,N_18869,N_18895);
or U19109 (N_19109,N_18944,N_18914);
or U19110 (N_19110,N_18906,N_18950);
xnor U19111 (N_19111,N_18845,N_18853);
nor U19112 (N_19112,N_18807,N_18980);
and U19113 (N_19113,N_18874,N_18918);
nand U19114 (N_19114,N_18804,N_18988);
and U19115 (N_19115,N_18836,N_18947);
xor U19116 (N_19116,N_18919,N_18890);
nor U19117 (N_19117,N_18941,N_18832);
and U19118 (N_19118,N_18975,N_18854);
and U19119 (N_19119,N_18807,N_18922);
nand U19120 (N_19120,N_18822,N_18916);
and U19121 (N_19121,N_18845,N_18840);
nor U19122 (N_19122,N_18977,N_18965);
or U19123 (N_19123,N_18989,N_18863);
or U19124 (N_19124,N_18927,N_18930);
and U19125 (N_19125,N_18825,N_18910);
xnor U19126 (N_19126,N_18830,N_18953);
nand U19127 (N_19127,N_18890,N_18818);
or U19128 (N_19128,N_18921,N_18800);
nor U19129 (N_19129,N_18984,N_18931);
nor U19130 (N_19130,N_18939,N_18886);
nand U19131 (N_19131,N_18854,N_18945);
nor U19132 (N_19132,N_18838,N_18825);
nand U19133 (N_19133,N_18882,N_18929);
nand U19134 (N_19134,N_18877,N_18837);
nor U19135 (N_19135,N_18822,N_18889);
or U19136 (N_19136,N_18971,N_18855);
nor U19137 (N_19137,N_18876,N_18848);
xnor U19138 (N_19138,N_18819,N_18968);
and U19139 (N_19139,N_18942,N_18909);
nand U19140 (N_19140,N_18942,N_18830);
nor U19141 (N_19141,N_18886,N_18849);
or U19142 (N_19142,N_18935,N_18868);
or U19143 (N_19143,N_18820,N_18865);
and U19144 (N_19144,N_18839,N_18924);
nor U19145 (N_19145,N_18814,N_18984);
nor U19146 (N_19146,N_18990,N_18929);
nor U19147 (N_19147,N_18989,N_18909);
and U19148 (N_19148,N_18819,N_18924);
and U19149 (N_19149,N_18964,N_18864);
nor U19150 (N_19150,N_18930,N_18901);
nor U19151 (N_19151,N_18977,N_18944);
nand U19152 (N_19152,N_18962,N_18973);
nor U19153 (N_19153,N_18901,N_18883);
nor U19154 (N_19154,N_18863,N_18965);
xnor U19155 (N_19155,N_18900,N_18852);
or U19156 (N_19156,N_18881,N_18972);
and U19157 (N_19157,N_18813,N_18838);
or U19158 (N_19158,N_18868,N_18996);
nand U19159 (N_19159,N_18943,N_18968);
and U19160 (N_19160,N_18894,N_18999);
nand U19161 (N_19161,N_18954,N_18875);
nor U19162 (N_19162,N_18844,N_18830);
nand U19163 (N_19163,N_18972,N_18803);
and U19164 (N_19164,N_18807,N_18830);
nor U19165 (N_19165,N_18829,N_18958);
nand U19166 (N_19166,N_18850,N_18880);
and U19167 (N_19167,N_18850,N_18862);
or U19168 (N_19168,N_18963,N_18909);
nand U19169 (N_19169,N_18950,N_18885);
xnor U19170 (N_19170,N_18947,N_18851);
or U19171 (N_19171,N_18944,N_18993);
and U19172 (N_19172,N_18878,N_18913);
or U19173 (N_19173,N_18971,N_18903);
xnor U19174 (N_19174,N_18968,N_18875);
nand U19175 (N_19175,N_18894,N_18812);
nor U19176 (N_19176,N_18879,N_18941);
nor U19177 (N_19177,N_18877,N_18899);
nand U19178 (N_19178,N_18866,N_18832);
and U19179 (N_19179,N_18877,N_18984);
nor U19180 (N_19180,N_18994,N_18903);
or U19181 (N_19181,N_18957,N_18807);
nor U19182 (N_19182,N_18892,N_18943);
nand U19183 (N_19183,N_18928,N_18999);
nor U19184 (N_19184,N_18996,N_18946);
or U19185 (N_19185,N_18891,N_18914);
nor U19186 (N_19186,N_18825,N_18974);
or U19187 (N_19187,N_18971,N_18991);
nor U19188 (N_19188,N_18902,N_18974);
xor U19189 (N_19189,N_18925,N_18974);
xnor U19190 (N_19190,N_18919,N_18907);
or U19191 (N_19191,N_18977,N_18942);
xor U19192 (N_19192,N_18990,N_18973);
nand U19193 (N_19193,N_18846,N_18877);
nor U19194 (N_19194,N_18965,N_18905);
and U19195 (N_19195,N_18916,N_18874);
nand U19196 (N_19196,N_18844,N_18976);
and U19197 (N_19197,N_18891,N_18827);
and U19198 (N_19198,N_18930,N_18879);
nand U19199 (N_19199,N_18845,N_18899);
nor U19200 (N_19200,N_19113,N_19022);
and U19201 (N_19201,N_19147,N_19074);
or U19202 (N_19202,N_19060,N_19011);
nor U19203 (N_19203,N_19144,N_19170);
nand U19204 (N_19204,N_19134,N_19059);
or U19205 (N_19205,N_19108,N_19065);
or U19206 (N_19206,N_19000,N_19056);
and U19207 (N_19207,N_19177,N_19067);
and U19208 (N_19208,N_19194,N_19143);
nand U19209 (N_19209,N_19031,N_19127);
nor U19210 (N_19210,N_19032,N_19027);
and U19211 (N_19211,N_19186,N_19048);
and U19212 (N_19212,N_19198,N_19173);
nor U19213 (N_19213,N_19165,N_19136);
and U19214 (N_19214,N_19039,N_19007);
nor U19215 (N_19215,N_19171,N_19077);
and U19216 (N_19216,N_19174,N_19179);
nand U19217 (N_19217,N_19195,N_19149);
nand U19218 (N_19218,N_19097,N_19141);
xnor U19219 (N_19219,N_19068,N_19138);
xnor U19220 (N_19220,N_19193,N_19129);
nand U19221 (N_19221,N_19093,N_19047);
nand U19222 (N_19222,N_19043,N_19044);
nor U19223 (N_19223,N_19063,N_19159);
and U19224 (N_19224,N_19050,N_19101);
and U19225 (N_19225,N_19025,N_19166);
nor U19226 (N_19226,N_19040,N_19098);
nand U19227 (N_19227,N_19055,N_19158);
and U19228 (N_19228,N_19153,N_19045);
nor U19229 (N_19229,N_19066,N_19169);
or U19230 (N_19230,N_19140,N_19085);
or U19231 (N_19231,N_19006,N_19100);
or U19232 (N_19232,N_19124,N_19145);
nor U19233 (N_19233,N_19054,N_19035);
and U19234 (N_19234,N_19062,N_19163);
xnor U19235 (N_19235,N_19151,N_19041);
xor U19236 (N_19236,N_19162,N_19038);
or U19237 (N_19237,N_19087,N_19185);
nand U19238 (N_19238,N_19105,N_19137);
nand U19239 (N_19239,N_19103,N_19155);
and U19240 (N_19240,N_19191,N_19086);
or U19241 (N_19241,N_19160,N_19181);
nor U19242 (N_19242,N_19003,N_19088);
nand U19243 (N_19243,N_19182,N_19073);
xnor U19244 (N_19244,N_19161,N_19197);
nand U19245 (N_19245,N_19072,N_19018);
or U19246 (N_19246,N_19010,N_19164);
or U19247 (N_19247,N_19116,N_19172);
and U19248 (N_19248,N_19064,N_19090);
and U19249 (N_19249,N_19157,N_19148);
or U19250 (N_19250,N_19167,N_19115);
nor U19251 (N_19251,N_19046,N_19114);
nor U19252 (N_19252,N_19037,N_19019);
and U19253 (N_19253,N_19049,N_19069);
or U19254 (N_19254,N_19092,N_19130);
or U19255 (N_19255,N_19080,N_19107);
and U19256 (N_19256,N_19152,N_19094);
xor U19257 (N_19257,N_19014,N_19030);
or U19258 (N_19258,N_19075,N_19057);
or U19259 (N_19259,N_19199,N_19109);
nand U19260 (N_19260,N_19146,N_19112);
or U19261 (N_19261,N_19023,N_19175);
xnor U19262 (N_19262,N_19081,N_19099);
or U19263 (N_19263,N_19036,N_19089);
nand U19264 (N_19264,N_19096,N_19102);
nand U19265 (N_19265,N_19071,N_19029);
nor U19266 (N_19266,N_19015,N_19128);
nand U19267 (N_19267,N_19133,N_19188);
or U19268 (N_19268,N_19021,N_19189);
nand U19269 (N_19269,N_19156,N_19119);
and U19270 (N_19270,N_19013,N_19123);
nor U19271 (N_19271,N_19034,N_19016);
nand U19272 (N_19272,N_19070,N_19192);
or U19273 (N_19273,N_19196,N_19001);
nand U19274 (N_19274,N_19076,N_19122);
nand U19275 (N_19275,N_19178,N_19111);
nand U19276 (N_19276,N_19168,N_19083);
nor U19277 (N_19277,N_19079,N_19190);
and U19278 (N_19278,N_19142,N_19012);
nor U19279 (N_19279,N_19117,N_19154);
or U19280 (N_19280,N_19187,N_19051);
and U19281 (N_19281,N_19042,N_19118);
nand U19282 (N_19282,N_19028,N_19005);
or U19283 (N_19283,N_19058,N_19082);
nand U19284 (N_19284,N_19126,N_19008);
nand U19285 (N_19285,N_19104,N_19184);
nand U19286 (N_19286,N_19002,N_19091);
nand U19287 (N_19287,N_19020,N_19132);
nand U19288 (N_19288,N_19183,N_19106);
nand U19289 (N_19289,N_19033,N_19061);
nand U19290 (N_19290,N_19095,N_19131);
and U19291 (N_19291,N_19017,N_19150);
xor U19292 (N_19292,N_19110,N_19139);
and U19293 (N_19293,N_19125,N_19135);
or U19294 (N_19294,N_19084,N_19052);
nor U19295 (N_19295,N_19026,N_19078);
and U19296 (N_19296,N_19009,N_19176);
and U19297 (N_19297,N_19024,N_19053);
nand U19298 (N_19298,N_19004,N_19180);
nand U19299 (N_19299,N_19121,N_19120);
or U19300 (N_19300,N_19150,N_19004);
nand U19301 (N_19301,N_19177,N_19049);
nor U19302 (N_19302,N_19069,N_19041);
or U19303 (N_19303,N_19111,N_19099);
nor U19304 (N_19304,N_19070,N_19106);
or U19305 (N_19305,N_19133,N_19123);
or U19306 (N_19306,N_19001,N_19031);
nand U19307 (N_19307,N_19041,N_19137);
and U19308 (N_19308,N_19103,N_19096);
or U19309 (N_19309,N_19053,N_19076);
or U19310 (N_19310,N_19035,N_19140);
and U19311 (N_19311,N_19083,N_19166);
or U19312 (N_19312,N_19178,N_19153);
and U19313 (N_19313,N_19187,N_19116);
nor U19314 (N_19314,N_19115,N_19051);
and U19315 (N_19315,N_19193,N_19113);
nor U19316 (N_19316,N_19082,N_19076);
nor U19317 (N_19317,N_19164,N_19197);
and U19318 (N_19318,N_19093,N_19120);
nor U19319 (N_19319,N_19049,N_19184);
and U19320 (N_19320,N_19135,N_19009);
and U19321 (N_19321,N_19024,N_19078);
and U19322 (N_19322,N_19046,N_19033);
nor U19323 (N_19323,N_19152,N_19013);
or U19324 (N_19324,N_19180,N_19041);
nor U19325 (N_19325,N_19097,N_19046);
or U19326 (N_19326,N_19011,N_19028);
xnor U19327 (N_19327,N_19157,N_19194);
and U19328 (N_19328,N_19024,N_19064);
and U19329 (N_19329,N_19110,N_19159);
nand U19330 (N_19330,N_19185,N_19079);
nand U19331 (N_19331,N_19069,N_19062);
or U19332 (N_19332,N_19197,N_19168);
or U19333 (N_19333,N_19130,N_19149);
xnor U19334 (N_19334,N_19036,N_19081);
or U19335 (N_19335,N_19113,N_19061);
xor U19336 (N_19336,N_19081,N_19065);
nor U19337 (N_19337,N_19062,N_19035);
xor U19338 (N_19338,N_19130,N_19185);
nor U19339 (N_19339,N_19043,N_19183);
and U19340 (N_19340,N_19191,N_19111);
xnor U19341 (N_19341,N_19158,N_19125);
or U19342 (N_19342,N_19006,N_19120);
or U19343 (N_19343,N_19157,N_19095);
nand U19344 (N_19344,N_19103,N_19025);
or U19345 (N_19345,N_19023,N_19155);
nor U19346 (N_19346,N_19096,N_19004);
or U19347 (N_19347,N_19012,N_19135);
xnor U19348 (N_19348,N_19032,N_19058);
nor U19349 (N_19349,N_19176,N_19114);
nand U19350 (N_19350,N_19122,N_19012);
and U19351 (N_19351,N_19092,N_19066);
nand U19352 (N_19352,N_19042,N_19051);
nor U19353 (N_19353,N_19088,N_19118);
xor U19354 (N_19354,N_19085,N_19008);
or U19355 (N_19355,N_19183,N_19186);
and U19356 (N_19356,N_19102,N_19063);
or U19357 (N_19357,N_19078,N_19004);
nor U19358 (N_19358,N_19003,N_19166);
or U19359 (N_19359,N_19113,N_19166);
nand U19360 (N_19360,N_19108,N_19160);
nor U19361 (N_19361,N_19035,N_19198);
and U19362 (N_19362,N_19165,N_19029);
nor U19363 (N_19363,N_19169,N_19124);
and U19364 (N_19364,N_19177,N_19111);
nor U19365 (N_19365,N_19149,N_19180);
xnor U19366 (N_19366,N_19021,N_19038);
xnor U19367 (N_19367,N_19049,N_19189);
and U19368 (N_19368,N_19030,N_19182);
nand U19369 (N_19369,N_19150,N_19058);
or U19370 (N_19370,N_19032,N_19166);
nand U19371 (N_19371,N_19028,N_19072);
nor U19372 (N_19372,N_19125,N_19116);
nor U19373 (N_19373,N_19143,N_19131);
and U19374 (N_19374,N_19185,N_19077);
and U19375 (N_19375,N_19123,N_19082);
or U19376 (N_19376,N_19153,N_19199);
nor U19377 (N_19377,N_19089,N_19127);
or U19378 (N_19378,N_19135,N_19019);
and U19379 (N_19379,N_19017,N_19170);
xnor U19380 (N_19380,N_19023,N_19118);
nor U19381 (N_19381,N_19020,N_19072);
or U19382 (N_19382,N_19064,N_19167);
nor U19383 (N_19383,N_19184,N_19107);
and U19384 (N_19384,N_19034,N_19189);
and U19385 (N_19385,N_19192,N_19098);
nand U19386 (N_19386,N_19074,N_19174);
nand U19387 (N_19387,N_19072,N_19071);
or U19388 (N_19388,N_19061,N_19104);
nor U19389 (N_19389,N_19039,N_19194);
nor U19390 (N_19390,N_19029,N_19012);
nand U19391 (N_19391,N_19030,N_19068);
or U19392 (N_19392,N_19007,N_19041);
nor U19393 (N_19393,N_19188,N_19128);
nor U19394 (N_19394,N_19154,N_19157);
and U19395 (N_19395,N_19159,N_19001);
or U19396 (N_19396,N_19173,N_19029);
and U19397 (N_19397,N_19117,N_19062);
nor U19398 (N_19398,N_19193,N_19110);
and U19399 (N_19399,N_19105,N_19051);
nand U19400 (N_19400,N_19279,N_19295);
nor U19401 (N_19401,N_19271,N_19316);
nand U19402 (N_19402,N_19353,N_19255);
nor U19403 (N_19403,N_19370,N_19208);
and U19404 (N_19404,N_19352,N_19260);
nand U19405 (N_19405,N_19224,N_19345);
or U19406 (N_19406,N_19376,N_19235);
nand U19407 (N_19407,N_19354,N_19356);
and U19408 (N_19408,N_19315,N_19296);
and U19409 (N_19409,N_19344,N_19283);
nor U19410 (N_19410,N_19321,N_19364);
nand U19411 (N_19411,N_19351,N_19268);
xor U19412 (N_19412,N_19237,N_19392);
xnor U19413 (N_19413,N_19302,N_19294);
nor U19414 (N_19414,N_19385,N_19336);
xor U19415 (N_19415,N_19250,N_19375);
or U19416 (N_19416,N_19209,N_19361);
or U19417 (N_19417,N_19387,N_19388);
and U19418 (N_19418,N_19310,N_19277);
or U19419 (N_19419,N_19319,N_19257);
or U19420 (N_19420,N_19382,N_19236);
or U19421 (N_19421,N_19244,N_19234);
or U19422 (N_19422,N_19258,N_19333);
nand U19423 (N_19423,N_19281,N_19301);
nor U19424 (N_19424,N_19280,N_19332);
nand U19425 (N_19425,N_19396,N_19338);
or U19426 (N_19426,N_19335,N_19327);
and U19427 (N_19427,N_19232,N_19222);
xor U19428 (N_19428,N_19263,N_19306);
and U19429 (N_19429,N_19223,N_19313);
nand U19430 (N_19430,N_19233,N_19220);
or U19431 (N_19431,N_19297,N_19307);
xor U19432 (N_19432,N_19329,N_19308);
xnor U19433 (N_19433,N_19290,N_19379);
xnor U19434 (N_19434,N_19241,N_19239);
nor U19435 (N_19435,N_19386,N_19289);
and U19436 (N_19436,N_19265,N_19398);
xnor U19437 (N_19437,N_19276,N_19347);
and U19438 (N_19438,N_19215,N_19285);
nand U19439 (N_19439,N_19346,N_19328);
or U19440 (N_19440,N_19348,N_19372);
and U19441 (N_19441,N_19355,N_19324);
or U19442 (N_19442,N_19331,N_19202);
nand U19443 (N_19443,N_19286,N_19261);
and U19444 (N_19444,N_19391,N_19300);
or U19445 (N_19445,N_19221,N_19311);
nor U19446 (N_19446,N_19211,N_19217);
nand U19447 (N_19447,N_19225,N_19323);
xor U19448 (N_19448,N_19360,N_19359);
and U19449 (N_19449,N_19251,N_19274);
and U19450 (N_19450,N_19287,N_19216);
nor U19451 (N_19451,N_19342,N_19341);
or U19452 (N_19452,N_19358,N_19349);
nor U19453 (N_19453,N_19243,N_19309);
and U19454 (N_19454,N_19380,N_19254);
nand U19455 (N_19455,N_19339,N_19377);
nand U19456 (N_19456,N_19288,N_19325);
and U19457 (N_19457,N_19262,N_19245);
and U19458 (N_19458,N_19206,N_19374);
or U19459 (N_19459,N_19397,N_19350);
or U19460 (N_19460,N_19298,N_19264);
nor U19461 (N_19461,N_19210,N_19334);
or U19462 (N_19462,N_19267,N_19282);
nor U19463 (N_19463,N_19242,N_19205);
or U19464 (N_19464,N_19259,N_19240);
nor U19465 (N_19465,N_19228,N_19278);
or U19466 (N_19466,N_19213,N_19365);
or U19467 (N_19467,N_19390,N_19273);
nand U19468 (N_19468,N_19337,N_19395);
and U19469 (N_19469,N_19389,N_19291);
nor U19470 (N_19470,N_19203,N_19266);
nor U19471 (N_19471,N_19381,N_19330);
nand U19472 (N_19472,N_19284,N_19368);
and U19473 (N_19473,N_19305,N_19292);
nand U19474 (N_19474,N_19343,N_19394);
and U19475 (N_19475,N_19214,N_19312);
nor U19476 (N_19476,N_19246,N_19229);
and U19477 (N_19477,N_19357,N_19303);
nand U19478 (N_19478,N_19275,N_19304);
nand U19479 (N_19479,N_19201,N_19366);
nand U19480 (N_19480,N_19318,N_19367);
xor U19481 (N_19481,N_19218,N_19320);
and U19482 (N_19482,N_19231,N_19369);
nor U19483 (N_19483,N_19371,N_19227);
or U19484 (N_19484,N_19299,N_19362);
or U19485 (N_19485,N_19238,N_19200);
nand U19486 (N_19486,N_19322,N_19212);
nand U19487 (N_19487,N_19207,N_19384);
nand U19488 (N_19488,N_19256,N_19204);
nand U19489 (N_19489,N_19248,N_19226);
or U19490 (N_19490,N_19314,N_19317);
nand U19491 (N_19491,N_19247,N_19269);
nand U19492 (N_19492,N_19230,N_19399);
and U19493 (N_19493,N_19363,N_19393);
or U19494 (N_19494,N_19270,N_19378);
or U19495 (N_19495,N_19219,N_19373);
and U19496 (N_19496,N_19383,N_19249);
xnor U19497 (N_19497,N_19340,N_19326);
and U19498 (N_19498,N_19252,N_19272);
or U19499 (N_19499,N_19293,N_19253);
nand U19500 (N_19500,N_19393,N_19318);
or U19501 (N_19501,N_19262,N_19321);
nor U19502 (N_19502,N_19365,N_19335);
xor U19503 (N_19503,N_19204,N_19306);
nand U19504 (N_19504,N_19272,N_19346);
nand U19505 (N_19505,N_19238,N_19313);
or U19506 (N_19506,N_19319,N_19381);
xor U19507 (N_19507,N_19291,N_19320);
nor U19508 (N_19508,N_19258,N_19209);
or U19509 (N_19509,N_19270,N_19336);
nand U19510 (N_19510,N_19200,N_19261);
nand U19511 (N_19511,N_19306,N_19347);
nand U19512 (N_19512,N_19211,N_19259);
nor U19513 (N_19513,N_19384,N_19354);
xnor U19514 (N_19514,N_19316,N_19273);
or U19515 (N_19515,N_19342,N_19270);
or U19516 (N_19516,N_19360,N_19234);
nand U19517 (N_19517,N_19396,N_19235);
and U19518 (N_19518,N_19247,N_19284);
nor U19519 (N_19519,N_19228,N_19323);
nand U19520 (N_19520,N_19354,N_19323);
nor U19521 (N_19521,N_19216,N_19283);
nor U19522 (N_19522,N_19378,N_19233);
nor U19523 (N_19523,N_19385,N_19296);
xor U19524 (N_19524,N_19310,N_19221);
nand U19525 (N_19525,N_19305,N_19282);
nor U19526 (N_19526,N_19274,N_19372);
nor U19527 (N_19527,N_19216,N_19278);
or U19528 (N_19528,N_19373,N_19346);
xnor U19529 (N_19529,N_19313,N_19397);
nand U19530 (N_19530,N_19283,N_19320);
or U19531 (N_19531,N_19262,N_19241);
and U19532 (N_19532,N_19213,N_19343);
nor U19533 (N_19533,N_19322,N_19337);
and U19534 (N_19534,N_19367,N_19265);
nor U19535 (N_19535,N_19234,N_19379);
or U19536 (N_19536,N_19200,N_19327);
nand U19537 (N_19537,N_19245,N_19326);
and U19538 (N_19538,N_19238,N_19342);
nand U19539 (N_19539,N_19222,N_19294);
or U19540 (N_19540,N_19294,N_19279);
nand U19541 (N_19541,N_19352,N_19332);
nor U19542 (N_19542,N_19370,N_19345);
or U19543 (N_19543,N_19372,N_19324);
nand U19544 (N_19544,N_19256,N_19314);
and U19545 (N_19545,N_19247,N_19271);
xor U19546 (N_19546,N_19399,N_19209);
nor U19547 (N_19547,N_19333,N_19286);
nand U19548 (N_19548,N_19342,N_19387);
or U19549 (N_19549,N_19217,N_19322);
nor U19550 (N_19550,N_19361,N_19349);
xor U19551 (N_19551,N_19293,N_19265);
and U19552 (N_19552,N_19265,N_19222);
and U19553 (N_19553,N_19208,N_19274);
or U19554 (N_19554,N_19368,N_19201);
nor U19555 (N_19555,N_19311,N_19369);
nand U19556 (N_19556,N_19375,N_19268);
nor U19557 (N_19557,N_19238,N_19223);
or U19558 (N_19558,N_19310,N_19359);
or U19559 (N_19559,N_19289,N_19320);
nand U19560 (N_19560,N_19215,N_19263);
or U19561 (N_19561,N_19227,N_19248);
nor U19562 (N_19562,N_19315,N_19216);
xnor U19563 (N_19563,N_19290,N_19303);
or U19564 (N_19564,N_19339,N_19288);
or U19565 (N_19565,N_19258,N_19310);
and U19566 (N_19566,N_19241,N_19200);
or U19567 (N_19567,N_19310,N_19252);
and U19568 (N_19568,N_19200,N_19349);
and U19569 (N_19569,N_19361,N_19249);
or U19570 (N_19570,N_19266,N_19209);
xor U19571 (N_19571,N_19344,N_19298);
nor U19572 (N_19572,N_19250,N_19331);
or U19573 (N_19573,N_19323,N_19293);
nor U19574 (N_19574,N_19235,N_19273);
and U19575 (N_19575,N_19338,N_19359);
or U19576 (N_19576,N_19214,N_19341);
and U19577 (N_19577,N_19245,N_19294);
xor U19578 (N_19578,N_19365,N_19278);
nand U19579 (N_19579,N_19233,N_19201);
and U19580 (N_19580,N_19265,N_19395);
or U19581 (N_19581,N_19228,N_19269);
and U19582 (N_19582,N_19231,N_19280);
nor U19583 (N_19583,N_19364,N_19319);
nand U19584 (N_19584,N_19333,N_19380);
xnor U19585 (N_19585,N_19202,N_19264);
nor U19586 (N_19586,N_19361,N_19296);
nor U19587 (N_19587,N_19210,N_19264);
or U19588 (N_19588,N_19314,N_19372);
or U19589 (N_19589,N_19300,N_19368);
nand U19590 (N_19590,N_19327,N_19271);
and U19591 (N_19591,N_19231,N_19304);
or U19592 (N_19592,N_19218,N_19373);
and U19593 (N_19593,N_19217,N_19234);
nor U19594 (N_19594,N_19373,N_19280);
or U19595 (N_19595,N_19353,N_19206);
xnor U19596 (N_19596,N_19395,N_19282);
or U19597 (N_19597,N_19302,N_19299);
and U19598 (N_19598,N_19281,N_19283);
and U19599 (N_19599,N_19354,N_19269);
and U19600 (N_19600,N_19425,N_19502);
or U19601 (N_19601,N_19436,N_19478);
or U19602 (N_19602,N_19530,N_19486);
nor U19603 (N_19603,N_19414,N_19444);
nor U19604 (N_19604,N_19552,N_19514);
or U19605 (N_19605,N_19406,N_19430);
or U19606 (N_19606,N_19469,N_19472);
or U19607 (N_19607,N_19553,N_19400);
nor U19608 (N_19608,N_19494,N_19488);
nor U19609 (N_19609,N_19519,N_19590);
xnor U19610 (N_19610,N_19540,N_19550);
or U19611 (N_19611,N_19575,N_19578);
or U19612 (N_19612,N_19477,N_19547);
nor U19613 (N_19613,N_19588,N_19489);
and U19614 (N_19614,N_19545,N_19504);
or U19615 (N_19615,N_19466,N_19429);
nor U19616 (N_19616,N_19498,N_19420);
nand U19617 (N_19617,N_19585,N_19431);
xor U19618 (N_19618,N_19404,N_19490);
and U19619 (N_19619,N_19598,N_19450);
xnor U19620 (N_19620,N_19487,N_19546);
and U19621 (N_19621,N_19568,N_19559);
nor U19622 (N_19622,N_19426,N_19518);
nor U19623 (N_19623,N_19505,N_19438);
nor U19624 (N_19624,N_19543,N_19493);
nand U19625 (N_19625,N_19447,N_19491);
nor U19626 (N_19626,N_19577,N_19538);
or U19627 (N_19627,N_19599,N_19422);
xnor U19628 (N_19628,N_19419,N_19508);
nor U19629 (N_19629,N_19587,N_19462);
or U19630 (N_19630,N_19536,N_19537);
or U19631 (N_19631,N_19511,N_19448);
or U19632 (N_19632,N_19564,N_19573);
xor U19633 (N_19633,N_19432,N_19461);
xor U19634 (N_19634,N_19418,N_19459);
or U19635 (N_19635,N_19467,N_19566);
xnor U19636 (N_19636,N_19557,N_19596);
nor U19637 (N_19637,N_19421,N_19458);
and U19638 (N_19638,N_19501,N_19574);
or U19639 (N_19639,N_19417,N_19569);
or U19640 (N_19640,N_19463,N_19582);
nor U19641 (N_19641,N_19539,N_19453);
nor U19642 (N_19642,N_19509,N_19482);
and U19643 (N_19643,N_19401,N_19558);
nand U19644 (N_19644,N_19591,N_19551);
nor U19645 (N_19645,N_19423,N_19446);
and U19646 (N_19646,N_19480,N_19476);
nand U19647 (N_19647,N_19570,N_19521);
or U19648 (N_19648,N_19442,N_19500);
or U19649 (N_19649,N_19416,N_19524);
or U19650 (N_19650,N_19481,N_19441);
xor U19651 (N_19651,N_19464,N_19456);
and U19652 (N_19652,N_19457,N_19593);
nor U19653 (N_19653,N_19506,N_19405);
nand U19654 (N_19654,N_19556,N_19433);
nor U19655 (N_19655,N_19584,N_19497);
or U19656 (N_19656,N_19492,N_19445);
xnor U19657 (N_19657,N_19532,N_19529);
and U19658 (N_19658,N_19411,N_19548);
nor U19659 (N_19659,N_19403,N_19443);
nor U19660 (N_19660,N_19522,N_19424);
or U19661 (N_19661,N_19542,N_19499);
nand U19662 (N_19662,N_19525,N_19526);
nand U19663 (N_19663,N_19510,N_19579);
and U19664 (N_19664,N_19485,N_19562);
or U19665 (N_19665,N_19428,N_19580);
nand U19666 (N_19666,N_19440,N_19589);
and U19667 (N_19667,N_19449,N_19455);
and U19668 (N_19668,N_19474,N_19452);
nor U19669 (N_19669,N_19427,N_19495);
and U19670 (N_19670,N_19567,N_19512);
nand U19671 (N_19671,N_19435,N_19594);
nand U19672 (N_19672,N_19408,N_19451);
and U19673 (N_19673,N_19473,N_19415);
nand U19674 (N_19674,N_19533,N_19434);
nand U19675 (N_19675,N_19528,N_19439);
nand U19676 (N_19676,N_19527,N_19563);
and U19677 (N_19677,N_19483,N_19479);
nor U19678 (N_19678,N_19595,N_19412);
and U19679 (N_19679,N_19454,N_19592);
xor U19680 (N_19680,N_19507,N_19535);
and U19681 (N_19681,N_19496,N_19471);
nand U19682 (N_19682,N_19465,N_19581);
nor U19683 (N_19683,N_19583,N_19413);
and U19684 (N_19684,N_19407,N_19437);
nor U19685 (N_19685,N_19523,N_19410);
xor U19686 (N_19686,N_19571,N_19513);
or U19687 (N_19687,N_19555,N_19586);
and U19688 (N_19688,N_19576,N_19531);
nor U19689 (N_19689,N_19534,N_19409);
and U19690 (N_19690,N_19515,N_19541);
or U19691 (N_19691,N_19597,N_19565);
or U19692 (N_19692,N_19549,N_19460);
nand U19693 (N_19693,N_19402,N_19516);
or U19694 (N_19694,N_19517,N_19544);
or U19695 (N_19695,N_19554,N_19560);
and U19696 (N_19696,N_19484,N_19572);
and U19697 (N_19697,N_19520,N_19468);
nand U19698 (N_19698,N_19561,N_19470);
nand U19699 (N_19699,N_19475,N_19503);
nand U19700 (N_19700,N_19497,N_19585);
and U19701 (N_19701,N_19477,N_19590);
or U19702 (N_19702,N_19514,N_19481);
nor U19703 (N_19703,N_19437,N_19485);
nand U19704 (N_19704,N_19518,N_19590);
nand U19705 (N_19705,N_19416,N_19429);
nor U19706 (N_19706,N_19578,N_19460);
nor U19707 (N_19707,N_19439,N_19501);
xor U19708 (N_19708,N_19527,N_19561);
nor U19709 (N_19709,N_19518,N_19584);
and U19710 (N_19710,N_19493,N_19476);
nand U19711 (N_19711,N_19471,N_19525);
xor U19712 (N_19712,N_19572,N_19494);
and U19713 (N_19713,N_19560,N_19485);
xor U19714 (N_19714,N_19410,N_19571);
xor U19715 (N_19715,N_19427,N_19459);
nor U19716 (N_19716,N_19559,N_19428);
nand U19717 (N_19717,N_19484,N_19468);
or U19718 (N_19718,N_19559,N_19455);
or U19719 (N_19719,N_19532,N_19490);
or U19720 (N_19720,N_19561,N_19583);
xor U19721 (N_19721,N_19503,N_19526);
and U19722 (N_19722,N_19414,N_19500);
and U19723 (N_19723,N_19548,N_19570);
and U19724 (N_19724,N_19442,N_19594);
nand U19725 (N_19725,N_19512,N_19414);
nand U19726 (N_19726,N_19482,N_19456);
or U19727 (N_19727,N_19428,N_19485);
and U19728 (N_19728,N_19418,N_19435);
xor U19729 (N_19729,N_19559,N_19427);
nand U19730 (N_19730,N_19558,N_19525);
nand U19731 (N_19731,N_19541,N_19445);
nor U19732 (N_19732,N_19459,N_19400);
and U19733 (N_19733,N_19493,N_19508);
and U19734 (N_19734,N_19488,N_19460);
nand U19735 (N_19735,N_19525,N_19456);
nor U19736 (N_19736,N_19429,N_19437);
nor U19737 (N_19737,N_19576,N_19450);
or U19738 (N_19738,N_19504,N_19400);
or U19739 (N_19739,N_19428,N_19482);
nand U19740 (N_19740,N_19482,N_19540);
and U19741 (N_19741,N_19430,N_19512);
nand U19742 (N_19742,N_19532,N_19458);
nor U19743 (N_19743,N_19403,N_19462);
nand U19744 (N_19744,N_19500,N_19561);
nor U19745 (N_19745,N_19530,N_19542);
and U19746 (N_19746,N_19485,N_19411);
and U19747 (N_19747,N_19466,N_19518);
xnor U19748 (N_19748,N_19538,N_19597);
nor U19749 (N_19749,N_19430,N_19526);
nand U19750 (N_19750,N_19508,N_19560);
or U19751 (N_19751,N_19575,N_19588);
or U19752 (N_19752,N_19535,N_19466);
nor U19753 (N_19753,N_19451,N_19546);
and U19754 (N_19754,N_19442,N_19586);
and U19755 (N_19755,N_19442,N_19495);
or U19756 (N_19756,N_19500,N_19518);
and U19757 (N_19757,N_19466,N_19431);
and U19758 (N_19758,N_19530,N_19535);
nor U19759 (N_19759,N_19429,N_19419);
nand U19760 (N_19760,N_19437,N_19472);
nor U19761 (N_19761,N_19501,N_19565);
nand U19762 (N_19762,N_19584,N_19414);
nand U19763 (N_19763,N_19413,N_19469);
nand U19764 (N_19764,N_19499,N_19457);
or U19765 (N_19765,N_19552,N_19430);
nand U19766 (N_19766,N_19564,N_19468);
and U19767 (N_19767,N_19465,N_19413);
or U19768 (N_19768,N_19497,N_19457);
nand U19769 (N_19769,N_19545,N_19431);
nor U19770 (N_19770,N_19597,N_19427);
nor U19771 (N_19771,N_19566,N_19531);
nor U19772 (N_19772,N_19444,N_19549);
nand U19773 (N_19773,N_19454,N_19565);
nand U19774 (N_19774,N_19423,N_19533);
nor U19775 (N_19775,N_19561,N_19590);
and U19776 (N_19776,N_19545,N_19411);
nand U19777 (N_19777,N_19586,N_19597);
and U19778 (N_19778,N_19589,N_19577);
nor U19779 (N_19779,N_19415,N_19519);
nor U19780 (N_19780,N_19454,N_19550);
and U19781 (N_19781,N_19477,N_19569);
nor U19782 (N_19782,N_19565,N_19517);
and U19783 (N_19783,N_19511,N_19498);
and U19784 (N_19784,N_19460,N_19504);
and U19785 (N_19785,N_19543,N_19472);
or U19786 (N_19786,N_19538,N_19441);
or U19787 (N_19787,N_19426,N_19598);
nand U19788 (N_19788,N_19504,N_19483);
nor U19789 (N_19789,N_19500,N_19582);
nand U19790 (N_19790,N_19546,N_19437);
and U19791 (N_19791,N_19576,N_19520);
and U19792 (N_19792,N_19447,N_19507);
xnor U19793 (N_19793,N_19566,N_19580);
nor U19794 (N_19794,N_19526,N_19587);
and U19795 (N_19795,N_19454,N_19494);
nand U19796 (N_19796,N_19458,N_19474);
or U19797 (N_19797,N_19515,N_19497);
and U19798 (N_19798,N_19418,N_19579);
or U19799 (N_19799,N_19467,N_19418);
or U19800 (N_19800,N_19645,N_19698);
nand U19801 (N_19801,N_19697,N_19653);
and U19802 (N_19802,N_19690,N_19723);
nor U19803 (N_19803,N_19746,N_19620);
or U19804 (N_19804,N_19774,N_19617);
xor U19805 (N_19805,N_19739,N_19694);
or U19806 (N_19806,N_19753,N_19606);
nor U19807 (N_19807,N_19662,N_19627);
nand U19808 (N_19808,N_19670,N_19796);
nor U19809 (N_19809,N_19658,N_19671);
or U19810 (N_19810,N_19752,N_19794);
nand U19811 (N_19811,N_19637,N_19769);
and U19812 (N_19812,N_19649,N_19646);
nand U19813 (N_19813,N_19777,N_19675);
nor U19814 (N_19814,N_19695,N_19615);
or U19815 (N_19815,N_19710,N_19651);
or U19816 (N_19816,N_19773,N_19634);
or U19817 (N_19817,N_19795,N_19619);
xor U19818 (N_19818,N_19605,N_19727);
nand U19819 (N_19819,N_19785,N_19745);
and U19820 (N_19820,N_19603,N_19660);
and U19821 (N_19821,N_19701,N_19713);
nor U19822 (N_19822,N_19642,N_19706);
nor U19823 (N_19823,N_19728,N_19733);
and U19824 (N_19824,N_19643,N_19692);
nor U19825 (N_19825,N_19766,N_19640);
nor U19826 (N_19826,N_19784,N_19636);
nor U19827 (N_19827,N_19799,N_19737);
or U19828 (N_19828,N_19711,N_19780);
or U19829 (N_19829,N_19689,N_19602);
xnor U19830 (N_19830,N_19622,N_19715);
xor U19831 (N_19831,N_19741,N_19731);
xor U19832 (N_19832,N_19702,N_19758);
nand U19833 (N_19833,N_19765,N_19783);
and U19834 (N_19834,N_19750,N_19680);
nand U19835 (N_19835,N_19718,N_19779);
and U19836 (N_19836,N_19631,N_19629);
or U19837 (N_19837,N_19704,N_19687);
nand U19838 (N_19838,N_19663,N_19604);
nand U19839 (N_19839,N_19621,N_19635);
and U19840 (N_19840,N_19760,N_19664);
nor U19841 (N_19841,N_19612,N_19650);
nor U19842 (N_19842,N_19781,N_19652);
or U19843 (N_19843,N_19686,N_19764);
and U19844 (N_19844,N_19696,N_19744);
and U19845 (N_19845,N_19736,N_19788);
and U19846 (N_19846,N_19668,N_19786);
nor U19847 (N_19847,N_19759,N_19628);
and U19848 (N_19848,N_19638,N_19705);
nand U19849 (N_19849,N_19679,N_19756);
nor U19850 (N_19850,N_19755,N_19730);
nand U19851 (N_19851,N_19648,N_19610);
nand U19852 (N_19852,N_19655,N_19790);
nand U19853 (N_19853,N_19724,N_19616);
xnor U19854 (N_19854,N_19714,N_19797);
or U19855 (N_19855,N_19747,N_19729);
or U19856 (N_19856,N_19654,N_19632);
nor U19857 (N_19857,N_19682,N_19742);
nand U19858 (N_19858,N_19709,N_19613);
nor U19859 (N_19859,N_19776,N_19688);
nor U19860 (N_19860,N_19775,N_19630);
nor U19861 (N_19861,N_19661,N_19639);
or U19862 (N_19862,N_19707,N_19735);
nand U19863 (N_19863,N_19625,N_19789);
nor U19864 (N_19864,N_19666,N_19738);
nor U19865 (N_19865,N_19725,N_19683);
and U19866 (N_19866,N_19712,N_19600);
xor U19867 (N_19867,N_19677,N_19749);
nand U19868 (N_19868,N_19665,N_19626);
nor U19869 (N_19869,N_19607,N_19618);
nand U19870 (N_19870,N_19772,N_19601);
and U19871 (N_19871,N_19647,N_19726);
nand U19872 (N_19872,N_19757,N_19787);
or U19873 (N_19873,N_19624,N_19754);
or U19874 (N_19874,N_19768,N_19700);
nand U19875 (N_19875,N_19761,N_19762);
or U19876 (N_19876,N_19743,N_19608);
xor U19877 (N_19877,N_19732,N_19748);
or U19878 (N_19878,N_19657,N_19609);
nor U19879 (N_19879,N_19798,N_19678);
xnor U19880 (N_19880,N_19672,N_19722);
nor U19881 (N_19881,N_19767,N_19641);
xor U19882 (N_19882,N_19659,N_19720);
and U19883 (N_19883,N_19751,N_19667);
nor U19884 (N_19884,N_19770,N_19791);
and U19885 (N_19885,N_19674,N_19703);
and U19886 (N_19886,N_19669,N_19644);
nand U19887 (N_19887,N_19782,N_19771);
and U19888 (N_19888,N_19681,N_19691);
nor U19889 (N_19889,N_19716,N_19673);
and U19890 (N_19890,N_19676,N_19721);
and U19891 (N_19891,N_19614,N_19699);
nand U19892 (N_19892,N_19685,N_19740);
nand U19893 (N_19893,N_19611,N_19717);
and U19894 (N_19894,N_19708,N_19623);
nor U19895 (N_19895,N_19684,N_19693);
or U19896 (N_19896,N_19792,N_19734);
and U19897 (N_19897,N_19763,N_19793);
xnor U19898 (N_19898,N_19778,N_19719);
nor U19899 (N_19899,N_19633,N_19656);
nor U19900 (N_19900,N_19686,N_19743);
nand U19901 (N_19901,N_19663,N_19786);
nand U19902 (N_19902,N_19647,N_19666);
nor U19903 (N_19903,N_19618,N_19728);
or U19904 (N_19904,N_19620,N_19773);
and U19905 (N_19905,N_19674,N_19728);
or U19906 (N_19906,N_19637,N_19712);
or U19907 (N_19907,N_19676,N_19663);
and U19908 (N_19908,N_19662,N_19639);
or U19909 (N_19909,N_19686,N_19608);
nor U19910 (N_19910,N_19603,N_19615);
or U19911 (N_19911,N_19700,N_19601);
nor U19912 (N_19912,N_19766,N_19613);
nand U19913 (N_19913,N_19640,N_19688);
nor U19914 (N_19914,N_19677,N_19723);
and U19915 (N_19915,N_19601,N_19656);
nor U19916 (N_19916,N_19790,N_19639);
and U19917 (N_19917,N_19780,N_19666);
and U19918 (N_19918,N_19684,N_19688);
and U19919 (N_19919,N_19731,N_19627);
nand U19920 (N_19920,N_19663,N_19714);
nand U19921 (N_19921,N_19654,N_19732);
nand U19922 (N_19922,N_19785,N_19601);
and U19923 (N_19923,N_19734,N_19645);
and U19924 (N_19924,N_19706,N_19699);
or U19925 (N_19925,N_19686,N_19679);
nor U19926 (N_19926,N_19611,N_19718);
nor U19927 (N_19927,N_19688,N_19740);
nand U19928 (N_19928,N_19661,N_19622);
or U19929 (N_19929,N_19654,N_19776);
or U19930 (N_19930,N_19737,N_19661);
nor U19931 (N_19931,N_19662,N_19605);
and U19932 (N_19932,N_19771,N_19727);
and U19933 (N_19933,N_19698,N_19676);
or U19934 (N_19934,N_19793,N_19723);
xnor U19935 (N_19935,N_19688,N_19754);
nor U19936 (N_19936,N_19638,N_19725);
and U19937 (N_19937,N_19630,N_19755);
nand U19938 (N_19938,N_19697,N_19684);
nor U19939 (N_19939,N_19641,N_19797);
or U19940 (N_19940,N_19617,N_19780);
or U19941 (N_19941,N_19724,N_19606);
nor U19942 (N_19942,N_19602,N_19715);
xor U19943 (N_19943,N_19741,N_19740);
and U19944 (N_19944,N_19610,N_19638);
and U19945 (N_19945,N_19799,N_19701);
and U19946 (N_19946,N_19775,N_19642);
nand U19947 (N_19947,N_19742,N_19626);
or U19948 (N_19948,N_19692,N_19605);
nand U19949 (N_19949,N_19764,N_19601);
and U19950 (N_19950,N_19618,N_19620);
or U19951 (N_19951,N_19646,N_19615);
xnor U19952 (N_19952,N_19794,N_19683);
nor U19953 (N_19953,N_19613,N_19642);
xnor U19954 (N_19954,N_19795,N_19680);
xor U19955 (N_19955,N_19728,N_19672);
nor U19956 (N_19956,N_19662,N_19781);
and U19957 (N_19957,N_19771,N_19601);
or U19958 (N_19958,N_19691,N_19708);
and U19959 (N_19959,N_19733,N_19614);
and U19960 (N_19960,N_19711,N_19661);
or U19961 (N_19961,N_19759,N_19638);
or U19962 (N_19962,N_19736,N_19607);
nand U19963 (N_19963,N_19674,N_19654);
nand U19964 (N_19964,N_19613,N_19739);
and U19965 (N_19965,N_19651,N_19648);
or U19966 (N_19966,N_19631,N_19620);
xor U19967 (N_19967,N_19662,N_19614);
and U19968 (N_19968,N_19699,N_19719);
and U19969 (N_19969,N_19656,N_19698);
xor U19970 (N_19970,N_19701,N_19748);
xnor U19971 (N_19971,N_19694,N_19674);
nor U19972 (N_19972,N_19600,N_19663);
or U19973 (N_19973,N_19640,N_19617);
or U19974 (N_19974,N_19718,N_19692);
nand U19975 (N_19975,N_19622,N_19759);
nor U19976 (N_19976,N_19797,N_19617);
or U19977 (N_19977,N_19798,N_19723);
nor U19978 (N_19978,N_19718,N_19691);
or U19979 (N_19979,N_19650,N_19669);
nor U19980 (N_19980,N_19783,N_19640);
nand U19981 (N_19981,N_19670,N_19781);
or U19982 (N_19982,N_19776,N_19644);
xor U19983 (N_19983,N_19640,N_19661);
and U19984 (N_19984,N_19765,N_19607);
and U19985 (N_19985,N_19629,N_19700);
nand U19986 (N_19986,N_19710,N_19668);
nor U19987 (N_19987,N_19666,N_19674);
nand U19988 (N_19988,N_19764,N_19724);
xnor U19989 (N_19989,N_19674,N_19797);
xnor U19990 (N_19990,N_19754,N_19638);
nand U19991 (N_19991,N_19710,N_19754);
or U19992 (N_19992,N_19627,N_19691);
or U19993 (N_19993,N_19689,N_19690);
or U19994 (N_19994,N_19784,N_19680);
nor U19995 (N_19995,N_19758,N_19728);
nand U19996 (N_19996,N_19765,N_19782);
or U19997 (N_19997,N_19774,N_19694);
or U19998 (N_19998,N_19607,N_19785);
and U19999 (N_19999,N_19725,N_19694);
and U20000 (N_20000,N_19872,N_19866);
and U20001 (N_20001,N_19834,N_19888);
nand U20002 (N_20002,N_19826,N_19938);
or U20003 (N_20003,N_19835,N_19932);
nor U20004 (N_20004,N_19810,N_19953);
and U20005 (N_20005,N_19863,N_19919);
nor U20006 (N_20006,N_19928,N_19930);
and U20007 (N_20007,N_19956,N_19849);
and U20008 (N_20008,N_19947,N_19804);
nand U20009 (N_20009,N_19942,N_19975);
nand U20010 (N_20010,N_19952,N_19870);
nor U20011 (N_20011,N_19830,N_19802);
nand U20012 (N_20012,N_19861,N_19855);
xnor U20013 (N_20013,N_19901,N_19908);
or U20014 (N_20014,N_19865,N_19967);
or U20015 (N_20015,N_19836,N_19875);
nand U20016 (N_20016,N_19807,N_19937);
nand U20017 (N_20017,N_19976,N_19891);
and U20018 (N_20018,N_19852,N_19980);
and U20019 (N_20019,N_19824,N_19851);
or U20020 (N_20020,N_19904,N_19964);
and U20021 (N_20021,N_19945,N_19894);
and U20022 (N_20022,N_19931,N_19903);
nand U20023 (N_20023,N_19853,N_19998);
xor U20024 (N_20024,N_19969,N_19913);
and U20025 (N_20025,N_19800,N_19993);
or U20026 (N_20026,N_19848,N_19957);
or U20027 (N_20027,N_19858,N_19939);
and U20028 (N_20028,N_19944,N_19963);
and U20029 (N_20029,N_19959,N_19921);
and U20030 (N_20030,N_19879,N_19880);
nor U20031 (N_20031,N_19911,N_19902);
and U20032 (N_20032,N_19845,N_19914);
or U20033 (N_20033,N_19950,N_19847);
or U20034 (N_20034,N_19907,N_19869);
nand U20035 (N_20035,N_19949,N_19811);
nand U20036 (N_20036,N_19946,N_19996);
nand U20037 (N_20037,N_19815,N_19962);
or U20038 (N_20038,N_19829,N_19883);
nor U20039 (N_20039,N_19823,N_19805);
xor U20040 (N_20040,N_19933,N_19817);
nor U20041 (N_20041,N_19906,N_19862);
and U20042 (N_20042,N_19828,N_19889);
nand U20043 (N_20043,N_19974,N_19965);
nor U20044 (N_20044,N_19825,N_19896);
or U20045 (N_20045,N_19958,N_19832);
and U20046 (N_20046,N_19813,N_19920);
and U20047 (N_20047,N_19961,N_19886);
and U20048 (N_20048,N_19841,N_19857);
xor U20049 (N_20049,N_19842,N_19917);
nor U20050 (N_20050,N_19924,N_19999);
and U20051 (N_20051,N_19856,N_19812);
and U20052 (N_20052,N_19971,N_19951);
or U20053 (N_20053,N_19987,N_19981);
nor U20054 (N_20054,N_19882,N_19801);
nand U20055 (N_20055,N_19892,N_19833);
nor U20056 (N_20056,N_19838,N_19809);
or U20057 (N_20057,N_19927,N_19822);
xnor U20058 (N_20058,N_19867,N_19995);
xnor U20059 (N_20059,N_19955,N_19986);
nand U20060 (N_20060,N_19874,N_19816);
or U20061 (N_20061,N_19994,N_19827);
nand U20062 (N_20062,N_19923,N_19893);
nor U20063 (N_20063,N_19900,N_19873);
nor U20064 (N_20064,N_19990,N_19806);
or U20065 (N_20065,N_19820,N_19814);
and U20066 (N_20066,N_19915,N_19984);
or U20067 (N_20067,N_19941,N_19983);
nor U20068 (N_20068,N_19854,N_19899);
xor U20069 (N_20069,N_19885,N_19878);
xor U20070 (N_20070,N_19918,N_19982);
xnor U20071 (N_20071,N_19934,N_19881);
nand U20072 (N_20072,N_19843,N_19985);
nor U20073 (N_20073,N_19979,N_19940);
nor U20074 (N_20074,N_19803,N_19871);
nand U20075 (N_20075,N_19890,N_19978);
xor U20076 (N_20076,N_19808,N_19876);
or U20077 (N_20077,N_19821,N_19992);
nand U20078 (N_20078,N_19989,N_19831);
or U20079 (N_20079,N_19837,N_19910);
nor U20080 (N_20080,N_19898,N_19966);
nand U20081 (N_20081,N_19840,N_19970);
or U20082 (N_20082,N_19839,N_19948);
or U20083 (N_20083,N_19991,N_19895);
nor U20084 (N_20084,N_19972,N_19977);
nor U20085 (N_20085,N_19954,N_19909);
or U20086 (N_20086,N_19887,N_19988);
nor U20087 (N_20087,N_19868,N_19864);
nor U20088 (N_20088,N_19968,N_19960);
or U20089 (N_20089,N_19973,N_19818);
or U20090 (N_20090,N_19925,N_19844);
nand U20091 (N_20091,N_19922,N_19936);
nand U20092 (N_20092,N_19897,N_19929);
nor U20093 (N_20093,N_19877,N_19850);
nand U20094 (N_20094,N_19912,N_19860);
nand U20095 (N_20095,N_19916,N_19819);
or U20096 (N_20096,N_19997,N_19935);
nand U20097 (N_20097,N_19943,N_19846);
and U20098 (N_20098,N_19884,N_19926);
or U20099 (N_20099,N_19905,N_19859);
or U20100 (N_20100,N_19996,N_19909);
or U20101 (N_20101,N_19959,N_19800);
nor U20102 (N_20102,N_19952,N_19998);
and U20103 (N_20103,N_19873,N_19939);
xnor U20104 (N_20104,N_19840,N_19988);
or U20105 (N_20105,N_19959,N_19885);
nor U20106 (N_20106,N_19930,N_19926);
xnor U20107 (N_20107,N_19954,N_19861);
or U20108 (N_20108,N_19998,N_19844);
nand U20109 (N_20109,N_19837,N_19935);
nand U20110 (N_20110,N_19942,N_19950);
xnor U20111 (N_20111,N_19994,N_19940);
xor U20112 (N_20112,N_19976,N_19867);
and U20113 (N_20113,N_19809,N_19955);
xnor U20114 (N_20114,N_19990,N_19834);
and U20115 (N_20115,N_19901,N_19879);
nand U20116 (N_20116,N_19876,N_19908);
and U20117 (N_20117,N_19983,N_19800);
and U20118 (N_20118,N_19924,N_19917);
xnor U20119 (N_20119,N_19987,N_19863);
nand U20120 (N_20120,N_19922,N_19947);
and U20121 (N_20121,N_19940,N_19821);
nand U20122 (N_20122,N_19800,N_19844);
nor U20123 (N_20123,N_19932,N_19931);
nor U20124 (N_20124,N_19817,N_19961);
and U20125 (N_20125,N_19803,N_19950);
xnor U20126 (N_20126,N_19968,N_19823);
or U20127 (N_20127,N_19844,N_19973);
or U20128 (N_20128,N_19956,N_19808);
and U20129 (N_20129,N_19977,N_19987);
or U20130 (N_20130,N_19815,N_19835);
nor U20131 (N_20131,N_19984,N_19997);
nand U20132 (N_20132,N_19968,N_19898);
or U20133 (N_20133,N_19804,N_19848);
and U20134 (N_20134,N_19975,N_19887);
and U20135 (N_20135,N_19891,N_19871);
nand U20136 (N_20136,N_19983,N_19831);
and U20137 (N_20137,N_19944,N_19959);
or U20138 (N_20138,N_19844,N_19858);
nand U20139 (N_20139,N_19842,N_19961);
nand U20140 (N_20140,N_19959,N_19967);
and U20141 (N_20141,N_19969,N_19986);
nand U20142 (N_20142,N_19872,N_19966);
or U20143 (N_20143,N_19854,N_19879);
nand U20144 (N_20144,N_19938,N_19801);
nand U20145 (N_20145,N_19833,N_19920);
and U20146 (N_20146,N_19844,N_19954);
nand U20147 (N_20147,N_19845,N_19858);
or U20148 (N_20148,N_19969,N_19838);
or U20149 (N_20149,N_19828,N_19914);
nor U20150 (N_20150,N_19858,N_19974);
nand U20151 (N_20151,N_19814,N_19945);
and U20152 (N_20152,N_19984,N_19918);
or U20153 (N_20153,N_19891,N_19903);
or U20154 (N_20154,N_19971,N_19956);
nor U20155 (N_20155,N_19803,N_19855);
or U20156 (N_20156,N_19924,N_19945);
nand U20157 (N_20157,N_19864,N_19811);
nor U20158 (N_20158,N_19990,N_19999);
nor U20159 (N_20159,N_19849,N_19948);
and U20160 (N_20160,N_19837,N_19839);
nand U20161 (N_20161,N_19928,N_19999);
nor U20162 (N_20162,N_19922,N_19869);
xor U20163 (N_20163,N_19944,N_19992);
nor U20164 (N_20164,N_19849,N_19830);
or U20165 (N_20165,N_19884,N_19993);
and U20166 (N_20166,N_19916,N_19852);
xor U20167 (N_20167,N_19867,N_19833);
nor U20168 (N_20168,N_19867,N_19809);
nand U20169 (N_20169,N_19917,N_19944);
nand U20170 (N_20170,N_19805,N_19879);
or U20171 (N_20171,N_19855,N_19868);
or U20172 (N_20172,N_19838,N_19841);
nor U20173 (N_20173,N_19851,N_19926);
or U20174 (N_20174,N_19972,N_19843);
nor U20175 (N_20175,N_19993,N_19970);
or U20176 (N_20176,N_19965,N_19929);
and U20177 (N_20177,N_19932,N_19849);
or U20178 (N_20178,N_19902,N_19935);
and U20179 (N_20179,N_19890,N_19898);
nor U20180 (N_20180,N_19885,N_19837);
xnor U20181 (N_20181,N_19893,N_19907);
xnor U20182 (N_20182,N_19895,N_19857);
nand U20183 (N_20183,N_19847,N_19839);
and U20184 (N_20184,N_19999,N_19866);
nor U20185 (N_20185,N_19856,N_19938);
nor U20186 (N_20186,N_19810,N_19956);
or U20187 (N_20187,N_19991,N_19809);
and U20188 (N_20188,N_19854,N_19921);
xnor U20189 (N_20189,N_19879,N_19945);
or U20190 (N_20190,N_19963,N_19884);
nor U20191 (N_20191,N_19952,N_19999);
or U20192 (N_20192,N_19865,N_19839);
or U20193 (N_20193,N_19958,N_19884);
or U20194 (N_20194,N_19909,N_19893);
and U20195 (N_20195,N_19998,N_19989);
nor U20196 (N_20196,N_19923,N_19987);
nand U20197 (N_20197,N_19916,N_19888);
xnor U20198 (N_20198,N_19913,N_19919);
xnor U20199 (N_20199,N_19924,N_19822);
nand U20200 (N_20200,N_20163,N_20085);
or U20201 (N_20201,N_20195,N_20142);
or U20202 (N_20202,N_20102,N_20004);
or U20203 (N_20203,N_20106,N_20017);
nor U20204 (N_20204,N_20076,N_20104);
nor U20205 (N_20205,N_20198,N_20062);
and U20206 (N_20206,N_20147,N_20082);
xnor U20207 (N_20207,N_20118,N_20083);
nand U20208 (N_20208,N_20029,N_20024);
and U20209 (N_20209,N_20159,N_20068);
xor U20210 (N_20210,N_20079,N_20196);
or U20211 (N_20211,N_20047,N_20067);
nor U20212 (N_20212,N_20122,N_20049);
and U20213 (N_20213,N_20114,N_20141);
and U20214 (N_20214,N_20188,N_20095);
nand U20215 (N_20215,N_20026,N_20182);
xor U20216 (N_20216,N_20148,N_20116);
nand U20217 (N_20217,N_20077,N_20042);
nand U20218 (N_20218,N_20063,N_20121);
xnor U20219 (N_20219,N_20050,N_20112);
nor U20220 (N_20220,N_20000,N_20009);
nand U20221 (N_20221,N_20041,N_20027);
or U20222 (N_20222,N_20157,N_20130);
and U20223 (N_20223,N_20132,N_20185);
or U20224 (N_20224,N_20057,N_20133);
or U20225 (N_20225,N_20138,N_20107);
nand U20226 (N_20226,N_20014,N_20075);
nor U20227 (N_20227,N_20007,N_20015);
xor U20228 (N_20228,N_20018,N_20168);
nor U20229 (N_20229,N_20105,N_20080);
and U20230 (N_20230,N_20183,N_20139);
or U20231 (N_20231,N_20161,N_20137);
nand U20232 (N_20232,N_20061,N_20064);
and U20233 (N_20233,N_20180,N_20078);
nand U20234 (N_20234,N_20054,N_20113);
nand U20235 (N_20235,N_20028,N_20171);
xor U20236 (N_20236,N_20140,N_20094);
or U20237 (N_20237,N_20155,N_20020);
nor U20238 (N_20238,N_20001,N_20022);
xor U20239 (N_20239,N_20092,N_20103);
or U20240 (N_20240,N_20190,N_20158);
nor U20241 (N_20241,N_20143,N_20123);
nand U20242 (N_20242,N_20129,N_20101);
and U20243 (N_20243,N_20184,N_20152);
or U20244 (N_20244,N_20012,N_20175);
and U20245 (N_20245,N_20043,N_20053);
and U20246 (N_20246,N_20045,N_20179);
nand U20247 (N_20247,N_20099,N_20131);
or U20248 (N_20248,N_20164,N_20069);
and U20249 (N_20249,N_20034,N_20019);
nand U20250 (N_20250,N_20166,N_20192);
and U20251 (N_20251,N_20178,N_20193);
nor U20252 (N_20252,N_20070,N_20127);
and U20253 (N_20253,N_20153,N_20117);
nor U20254 (N_20254,N_20066,N_20109);
or U20255 (N_20255,N_20011,N_20181);
nand U20256 (N_20256,N_20073,N_20033);
and U20257 (N_20257,N_20037,N_20170);
and U20258 (N_20258,N_20174,N_20165);
or U20259 (N_20259,N_20032,N_20031);
xnor U20260 (N_20260,N_20016,N_20144);
nor U20261 (N_20261,N_20194,N_20097);
nand U20262 (N_20262,N_20044,N_20134);
and U20263 (N_20263,N_20046,N_20058);
and U20264 (N_20264,N_20167,N_20115);
nor U20265 (N_20265,N_20074,N_20065);
or U20266 (N_20266,N_20189,N_20021);
nor U20267 (N_20267,N_20187,N_20128);
xor U20268 (N_20268,N_20151,N_20119);
nor U20269 (N_20269,N_20197,N_20110);
nand U20270 (N_20270,N_20002,N_20060);
nand U20271 (N_20271,N_20172,N_20010);
or U20272 (N_20272,N_20048,N_20059);
nor U20273 (N_20273,N_20091,N_20149);
xor U20274 (N_20274,N_20088,N_20186);
and U20275 (N_20275,N_20154,N_20013);
or U20276 (N_20276,N_20005,N_20150);
nor U20277 (N_20277,N_20191,N_20036);
xor U20278 (N_20278,N_20156,N_20081);
nor U20279 (N_20279,N_20177,N_20030);
and U20280 (N_20280,N_20093,N_20145);
and U20281 (N_20281,N_20086,N_20176);
nor U20282 (N_20282,N_20100,N_20173);
and U20283 (N_20283,N_20035,N_20111);
nor U20284 (N_20284,N_20056,N_20124);
nand U20285 (N_20285,N_20136,N_20090);
or U20286 (N_20286,N_20162,N_20052);
nand U20287 (N_20287,N_20098,N_20084);
nand U20288 (N_20288,N_20146,N_20025);
nor U20289 (N_20289,N_20135,N_20039);
nor U20290 (N_20290,N_20126,N_20087);
nand U20291 (N_20291,N_20023,N_20120);
and U20292 (N_20292,N_20006,N_20072);
nand U20293 (N_20293,N_20040,N_20038);
xor U20294 (N_20294,N_20108,N_20199);
nand U20295 (N_20295,N_20051,N_20008);
or U20296 (N_20296,N_20003,N_20125);
or U20297 (N_20297,N_20169,N_20055);
and U20298 (N_20298,N_20089,N_20160);
nand U20299 (N_20299,N_20071,N_20096);
and U20300 (N_20300,N_20152,N_20172);
nor U20301 (N_20301,N_20163,N_20054);
or U20302 (N_20302,N_20016,N_20149);
nor U20303 (N_20303,N_20095,N_20149);
nand U20304 (N_20304,N_20057,N_20153);
nand U20305 (N_20305,N_20075,N_20008);
or U20306 (N_20306,N_20131,N_20020);
nand U20307 (N_20307,N_20113,N_20186);
and U20308 (N_20308,N_20098,N_20087);
and U20309 (N_20309,N_20040,N_20041);
or U20310 (N_20310,N_20162,N_20177);
and U20311 (N_20311,N_20076,N_20117);
nor U20312 (N_20312,N_20092,N_20105);
nor U20313 (N_20313,N_20178,N_20005);
or U20314 (N_20314,N_20197,N_20030);
nand U20315 (N_20315,N_20123,N_20046);
nand U20316 (N_20316,N_20092,N_20066);
nand U20317 (N_20317,N_20002,N_20056);
and U20318 (N_20318,N_20095,N_20160);
nor U20319 (N_20319,N_20166,N_20017);
nand U20320 (N_20320,N_20051,N_20190);
nor U20321 (N_20321,N_20173,N_20139);
and U20322 (N_20322,N_20194,N_20060);
xnor U20323 (N_20323,N_20083,N_20000);
and U20324 (N_20324,N_20043,N_20091);
or U20325 (N_20325,N_20046,N_20146);
and U20326 (N_20326,N_20168,N_20109);
nor U20327 (N_20327,N_20049,N_20178);
and U20328 (N_20328,N_20001,N_20065);
or U20329 (N_20329,N_20152,N_20079);
and U20330 (N_20330,N_20095,N_20124);
or U20331 (N_20331,N_20149,N_20045);
nand U20332 (N_20332,N_20073,N_20021);
nor U20333 (N_20333,N_20043,N_20039);
xnor U20334 (N_20334,N_20010,N_20042);
nor U20335 (N_20335,N_20078,N_20190);
nor U20336 (N_20336,N_20057,N_20149);
and U20337 (N_20337,N_20177,N_20007);
xor U20338 (N_20338,N_20148,N_20112);
nor U20339 (N_20339,N_20097,N_20185);
or U20340 (N_20340,N_20164,N_20098);
nor U20341 (N_20341,N_20124,N_20178);
nand U20342 (N_20342,N_20171,N_20056);
or U20343 (N_20343,N_20111,N_20097);
and U20344 (N_20344,N_20001,N_20111);
nand U20345 (N_20345,N_20112,N_20185);
and U20346 (N_20346,N_20188,N_20048);
xnor U20347 (N_20347,N_20184,N_20021);
nand U20348 (N_20348,N_20015,N_20076);
nor U20349 (N_20349,N_20196,N_20063);
nand U20350 (N_20350,N_20092,N_20111);
and U20351 (N_20351,N_20055,N_20014);
xor U20352 (N_20352,N_20109,N_20191);
and U20353 (N_20353,N_20135,N_20025);
xnor U20354 (N_20354,N_20119,N_20194);
nand U20355 (N_20355,N_20154,N_20189);
or U20356 (N_20356,N_20025,N_20102);
nor U20357 (N_20357,N_20076,N_20133);
nor U20358 (N_20358,N_20144,N_20012);
and U20359 (N_20359,N_20171,N_20196);
or U20360 (N_20360,N_20110,N_20065);
and U20361 (N_20361,N_20026,N_20142);
nand U20362 (N_20362,N_20002,N_20070);
nor U20363 (N_20363,N_20001,N_20003);
xor U20364 (N_20364,N_20020,N_20167);
nand U20365 (N_20365,N_20027,N_20030);
xor U20366 (N_20366,N_20085,N_20024);
and U20367 (N_20367,N_20141,N_20178);
and U20368 (N_20368,N_20004,N_20157);
and U20369 (N_20369,N_20095,N_20114);
and U20370 (N_20370,N_20021,N_20070);
and U20371 (N_20371,N_20025,N_20165);
and U20372 (N_20372,N_20055,N_20181);
nand U20373 (N_20373,N_20108,N_20131);
nor U20374 (N_20374,N_20188,N_20060);
and U20375 (N_20375,N_20179,N_20077);
or U20376 (N_20376,N_20083,N_20042);
nor U20377 (N_20377,N_20054,N_20075);
xor U20378 (N_20378,N_20046,N_20188);
or U20379 (N_20379,N_20163,N_20017);
or U20380 (N_20380,N_20037,N_20189);
nor U20381 (N_20381,N_20030,N_20194);
nand U20382 (N_20382,N_20104,N_20015);
nor U20383 (N_20383,N_20068,N_20092);
nand U20384 (N_20384,N_20154,N_20038);
or U20385 (N_20385,N_20127,N_20084);
and U20386 (N_20386,N_20106,N_20120);
or U20387 (N_20387,N_20142,N_20018);
nand U20388 (N_20388,N_20184,N_20197);
and U20389 (N_20389,N_20081,N_20130);
nor U20390 (N_20390,N_20183,N_20047);
nand U20391 (N_20391,N_20034,N_20052);
or U20392 (N_20392,N_20137,N_20065);
and U20393 (N_20393,N_20004,N_20160);
or U20394 (N_20394,N_20162,N_20040);
nor U20395 (N_20395,N_20078,N_20089);
nand U20396 (N_20396,N_20110,N_20134);
xor U20397 (N_20397,N_20115,N_20111);
and U20398 (N_20398,N_20128,N_20164);
and U20399 (N_20399,N_20101,N_20026);
and U20400 (N_20400,N_20370,N_20343);
nor U20401 (N_20401,N_20310,N_20315);
xor U20402 (N_20402,N_20201,N_20252);
nor U20403 (N_20403,N_20361,N_20278);
xnor U20404 (N_20404,N_20210,N_20214);
nor U20405 (N_20405,N_20247,N_20399);
and U20406 (N_20406,N_20307,N_20233);
nor U20407 (N_20407,N_20264,N_20240);
or U20408 (N_20408,N_20355,N_20276);
and U20409 (N_20409,N_20372,N_20313);
xnor U20410 (N_20410,N_20292,N_20272);
nor U20411 (N_20411,N_20288,N_20204);
nor U20412 (N_20412,N_20318,N_20294);
and U20413 (N_20413,N_20266,N_20270);
xor U20414 (N_20414,N_20291,N_20348);
and U20415 (N_20415,N_20301,N_20384);
or U20416 (N_20416,N_20212,N_20353);
or U20417 (N_20417,N_20256,N_20216);
and U20418 (N_20418,N_20223,N_20312);
nand U20419 (N_20419,N_20302,N_20297);
nand U20420 (N_20420,N_20218,N_20320);
and U20421 (N_20421,N_20251,N_20394);
and U20422 (N_20422,N_20308,N_20235);
nor U20423 (N_20423,N_20365,N_20236);
or U20424 (N_20424,N_20351,N_20249);
nand U20425 (N_20425,N_20362,N_20349);
and U20426 (N_20426,N_20222,N_20350);
or U20427 (N_20427,N_20385,N_20300);
and U20428 (N_20428,N_20289,N_20395);
and U20429 (N_20429,N_20225,N_20209);
nand U20430 (N_20430,N_20255,N_20335);
nand U20431 (N_20431,N_20284,N_20230);
xor U20432 (N_20432,N_20227,N_20366);
and U20433 (N_20433,N_20298,N_20281);
nand U20434 (N_20434,N_20244,N_20333);
nor U20435 (N_20435,N_20234,N_20316);
or U20436 (N_20436,N_20379,N_20293);
or U20437 (N_20437,N_20285,N_20322);
or U20438 (N_20438,N_20324,N_20306);
or U20439 (N_20439,N_20246,N_20398);
and U20440 (N_20440,N_20381,N_20211);
nand U20441 (N_20441,N_20220,N_20269);
xor U20442 (N_20442,N_20273,N_20331);
xor U20443 (N_20443,N_20241,N_20368);
nand U20444 (N_20444,N_20275,N_20397);
and U20445 (N_20445,N_20347,N_20338);
and U20446 (N_20446,N_20346,N_20257);
nor U20447 (N_20447,N_20279,N_20304);
nand U20448 (N_20448,N_20377,N_20260);
and U20449 (N_20449,N_20369,N_20382);
nand U20450 (N_20450,N_20376,N_20364);
xor U20451 (N_20451,N_20207,N_20339);
xor U20452 (N_20452,N_20245,N_20287);
nor U20453 (N_20453,N_20213,N_20259);
or U20454 (N_20454,N_20295,N_20277);
nor U20455 (N_20455,N_20340,N_20248);
nand U20456 (N_20456,N_20303,N_20224);
or U20457 (N_20457,N_20267,N_20296);
or U20458 (N_20458,N_20342,N_20392);
nand U20459 (N_20459,N_20387,N_20283);
and U20460 (N_20460,N_20268,N_20232);
and U20461 (N_20461,N_20299,N_20282);
xnor U20462 (N_20462,N_20373,N_20389);
and U20463 (N_20463,N_20242,N_20258);
nor U20464 (N_20464,N_20325,N_20286);
and U20465 (N_20465,N_20229,N_20357);
or U20466 (N_20466,N_20311,N_20206);
nor U20467 (N_20467,N_20396,N_20321);
and U20468 (N_20468,N_20202,N_20332);
or U20469 (N_20469,N_20323,N_20327);
and U20470 (N_20470,N_20388,N_20205);
xnor U20471 (N_20471,N_20203,N_20326);
nor U20472 (N_20472,N_20243,N_20334);
nor U20473 (N_20473,N_20378,N_20367);
xnor U20474 (N_20474,N_20330,N_20352);
or U20475 (N_20475,N_20386,N_20254);
or U20476 (N_20476,N_20261,N_20221);
xor U20477 (N_20477,N_20356,N_20341);
and U20478 (N_20478,N_20309,N_20380);
nand U20479 (N_20479,N_20290,N_20263);
or U20480 (N_20480,N_20317,N_20239);
or U20481 (N_20481,N_20358,N_20371);
nand U20482 (N_20482,N_20265,N_20226);
or U20483 (N_20483,N_20208,N_20271);
xor U20484 (N_20484,N_20305,N_20391);
and U20485 (N_20485,N_20383,N_20337);
nor U20486 (N_20486,N_20336,N_20344);
nand U20487 (N_20487,N_20262,N_20219);
xor U20488 (N_20488,N_20237,N_20314);
nand U20489 (N_20489,N_20390,N_20253);
nand U20490 (N_20490,N_20319,N_20375);
xnor U20491 (N_20491,N_20231,N_20274);
nor U20492 (N_20492,N_20215,N_20359);
nand U20493 (N_20493,N_20354,N_20345);
or U20494 (N_20494,N_20250,N_20200);
nand U20495 (N_20495,N_20238,N_20360);
and U20496 (N_20496,N_20374,N_20228);
nand U20497 (N_20497,N_20217,N_20329);
nor U20498 (N_20498,N_20328,N_20393);
or U20499 (N_20499,N_20363,N_20280);
nand U20500 (N_20500,N_20296,N_20383);
nor U20501 (N_20501,N_20383,N_20276);
or U20502 (N_20502,N_20214,N_20366);
nor U20503 (N_20503,N_20206,N_20315);
xor U20504 (N_20504,N_20217,N_20255);
nor U20505 (N_20505,N_20302,N_20260);
nor U20506 (N_20506,N_20325,N_20206);
nor U20507 (N_20507,N_20243,N_20279);
or U20508 (N_20508,N_20364,N_20236);
and U20509 (N_20509,N_20224,N_20241);
nand U20510 (N_20510,N_20310,N_20332);
or U20511 (N_20511,N_20314,N_20272);
nor U20512 (N_20512,N_20279,N_20335);
and U20513 (N_20513,N_20339,N_20367);
and U20514 (N_20514,N_20225,N_20203);
nor U20515 (N_20515,N_20391,N_20208);
nor U20516 (N_20516,N_20329,N_20378);
nand U20517 (N_20517,N_20398,N_20207);
or U20518 (N_20518,N_20255,N_20275);
nor U20519 (N_20519,N_20350,N_20323);
nor U20520 (N_20520,N_20267,N_20390);
xor U20521 (N_20521,N_20268,N_20360);
and U20522 (N_20522,N_20321,N_20240);
and U20523 (N_20523,N_20386,N_20290);
nand U20524 (N_20524,N_20397,N_20391);
nor U20525 (N_20525,N_20341,N_20377);
nor U20526 (N_20526,N_20305,N_20326);
nand U20527 (N_20527,N_20231,N_20305);
or U20528 (N_20528,N_20287,N_20330);
or U20529 (N_20529,N_20276,N_20261);
nor U20530 (N_20530,N_20337,N_20305);
nand U20531 (N_20531,N_20207,N_20235);
or U20532 (N_20532,N_20297,N_20390);
or U20533 (N_20533,N_20322,N_20397);
nand U20534 (N_20534,N_20274,N_20292);
or U20535 (N_20535,N_20305,N_20370);
and U20536 (N_20536,N_20232,N_20309);
or U20537 (N_20537,N_20369,N_20232);
and U20538 (N_20538,N_20304,N_20353);
and U20539 (N_20539,N_20209,N_20270);
nand U20540 (N_20540,N_20310,N_20384);
xor U20541 (N_20541,N_20371,N_20334);
xnor U20542 (N_20542,N_20265,N_20317);
xnor U20543 (N_20543,N_20338,N_20326);
nor U20544 (N_20544,N_20275,N_20243);
and U20545 (N_20545,N_20320,N_20342);
nor U20546 (N_20546,N_20290,N_20399);
nand U20547 (N_20547,N_20240,N_20245);
nand U20548 (N_20548,N_20260,N_20385);
nor U20549 (N_20549,N_20281,N_20275);
and U20550 (N_20550,N_20361,N_20272);
nand U20551 (N_20551,N_20378,N_20276);
or U20552 (N_20552,N_20232,N_20267);
xnor U20553 (N_20553,N_20337,N_20381);
nor U20554 (N_20554,N_20371,N_20315);
xnor U20555 (N_20555,N_20273,N_20286);
nand U20556 (N_20556,N_20259,N_20250);
or U20557 (N_20557,N_20310,N_20297);
nand U20558 (N_20558,N_20322,N_20241);
nand U20559 (N_20559,N_20270,N_20360);
nand U20560 (N_20560,N_20318,N_20374);
and U20561 (N_20561,N_20293,N_20214);
and U20562 (N_20562,N_20365,N_20261);
and U20563 (N_20563,N_20210,N_20387);
nand U20564 (N_20564,N_20229,N_20264);
xor U20565 (N_20565,N_20269,N_20294);
nand U20566 (N_20566,N_20397,N_20305);
nand U20567 (N_20567,N_20331,N_20352);
and U20568 (N_20568,N_20295,N_20301);
nand U20569 (N_20569,N_20211,N_20215);
nor U20570 (N_20570,N_20244,N_20256);
nand U20571 (N_20571,N_20225,N_20224);
nor U20572 (N_20572,N_20215,N_20331);
nand U20573 (N_20573,N_20369,N_20208);
nor U20574 (N_20574,N_20364,N_20328);
xnor U20575 (N_20575,N_20230,N_20258);
or U20576 (N_20576,N_20355,N_20328);
xor U20577 (N_20577,N_20386,N_20394);
or U20578 (N_20578,N_20319,N_20339);
nor U20579 (N_20579,N_20360,N_20247);
nor U20580 (N_20580,N_20357,N_20340);
or U20581 (N_20581,N_20234,N_20272);
nor U20582 (N_20582,N_20295,N_20303);
nand U20583 (N_20583,N_20261,N_20227);
nand U20584 (N_20584,N_20354,N_20388);
xor U20585 (N_20585,N_20263,N_20236);
or U20586 (N_20586,N_20258,N_20211);
and U20587 (N_20587,N_20268,N_20317);
xor U20588 (N_20588,N_20345,N_20289);
or U20589 (N_20589,N_20280,N_20376);
xnor U20590 (N_20590,N_20389,N_20353);
and U20591 (N_20591,N_20298,N_20211);
nand U20592 (N_20592,N_20368,N_20386);
and U20593 (N_20593,N_20254,N_20202);
nand U20594 (N_20594,N_20298,N_20383);
or U20595 (N_20595,N_20353,N_20397);
and U20596 (N_20596,N_20353,N_20379);
nor U20597 (N_20597,N_20329,N_20385);
nand U20598 (N_20598,N_20358,N_20257);
nand U20599 (N_20599,N_20390,N_20355);
nor U20600 (N_20600,N_20420,N_20467);
and U20601 (N_20601,N_20563,N_20528);
or U20602 (N_20602,N_20509,N_20573);
nor U20603 (N_20603,N_20434,N_20463);
or U20604 (N_20604,N_20400,N_20537);
or U20605 (N_20605,N_20476,N_20564);
or U20606 (N_20606,N_20550,N_20429);
nand U20607 (N_20607,N_20438,N_20462);
xor U20608 (N_20608,N_20512,N_20483);
nor U20609 (N_20609,N_20524,N_20422);
or U20610 (N_20610,N_20486,N_20406);
nand U20611 (N_20611,N_20530,N_20562);
nand U20612 (N_20612,N_20430,N_20408);
or U20613 (N_20613,N_20594,N_20587);
and U20614 (N_20614,N_20580,N_20506);
or U20615 (N_20615,N_20599,N_20591);
nand U20616 (N_20616,N_20470,N_20495);
and U20617 (N_20617,N_20458,N_20551);
nand U20618 (N_20618,N_20487,N_20445);
and U20619 (N_20619,N_20477,N_20541);
and U20620 (N_20620,N_20582,N_20540);
nor U20621 (N_20621,N_20576,N_20440);
nor U20622 (N_20622,N_20427,N_20584);
and U20623 (N_20623,N_20543,N_20535);
nor U20624 (N_20624,N_20407,N_20572);
nand U20625 (N_20625,N_20496,N_20553);
and U20626 (N_20626,N_20507,N_20414);
nor U20627 (N_20627,N_20560,N_20479);
and U20628 (N_20628,N_20539,N_20527);
nand U20629 (N_20629,N_20574,N_20416);
nand U20630 (N_20630,N_20525,N_20598);
nor U20631 (N_20631,N_20519,N_20471);
and U20632 (N_20632,N_20466,N_20450);
xor U20633 (N_20633,N_20554,N_20425);
or U20634 (N_20634,N_20451,N_20446);
nand U20635 (N_20635,N_20556,N_20449);
xor U20636 (N_20636,N_20474,N_20411);
or U20637 (N_20637,N_20452,N_20590);
nor U20638 (N_20638,N_20518,N_20510);
nand U20639 (N_20639,N_20546,N_20549);
nand U20640 (N_20640,N_20529,N_20577);
nor U20641 (N_20641,N_20557,N_20532);
nand U20642 (N_20642,N_20558,N_20480);
and U20643 (N_20643,N_20514,N_20475);
nor U20644 (N_20644,N_20405,N_20439);
and U20645 (N_20645,N_20473,N_20459);
or U20646 (N_20646,N_20404,N_20547);
nand U20647 (N_20647,N_20433,N_20538);
xor U20648 (N_20648,N_20578,N_20436);
nor U20649 (N_20649,N_20403,N_20453);
xnor U20650 (N_20650,N_20418,N_20465);
nor U20651 (N_20651,N_20575,N_20424);
and U20652 (N_20652,N_20454,N_20432);
nor U20653 (N_20653,N_20402,N_20423);
or U20654 (N_20654,N_20513,N_20570);
and U20655 (N_20655,N_20468,N_20501);
nand U20656 (N_20656,N_20502,N_20461);
and U20657 (N_20657,N_20504,N_20409);
and U20658 (N_20658,N_20516,N_20478);
and U20659 (N_20659,N_20567,N_20464);
and U20660 (N_20660,N_20484,N_20566);
and U20661 (N_20661,N_20413,N_20526);
and U20662 (N_20662,N_20508,N_20401);
nor U20663 (N_20663,N_20579,N_20491);
nor U20664 (N_20664,N_20428,N_20515);
xnor U20665 (N_20665,N_20583,N_20410);
nor U20666 (N_20666,N_20597,N_20531);
nand U20667 (N_20667,N_20426,N_20447);
nor U20668 (N_20668,N_20442,N_20585);
nor U20669 (N_20669,N_20421,N_20523);
or U20670 (N_20670,N_20494,N_20482);
xnor U20671 (N_20671,N_20457,N_20460);
nand U20672 (N_20672,N_20581,N_20561);
nor U20673 (N_20673,N_20492,N_20586);
and U20674 (N_20674,N_20493,N_20443);
nor U20675 (N_20675,N_20593,N_20521);
xnor U20676 (N_20676,N_20498,N_20559);
xnor U20677 (N_20677,N_20485,N_20488);
nor U20678 (N_20678,N_20522,N_20456);
or U20679 (N_20679,N_20444,N_20469);
nor U20680 (N_20680,N_20481,N_20500);
nand U20681 (N_20681,N_20588,N_20412);
and U20682 (N_20682,N_20441,N_20503);
and U20683 (N_20683,N_20415,N_20490);
and U20684 (N_20684,N_20555,N_20542);
nand U20685 (N_20685,N_20419,N_20448);
or U20686 (N_20686,N_20548,N_20505);
or U20687 (N_20687,N_20417,N_20534);
or U20688 (N_20688,N_20565,N_20595);
nand U20689 (N_20689,N_20511,N_20520);
and U20690 (N_20690,N_20431,N_20544);
nor U20691 (N_20691,N_20455,N_20489);
nor U20692 (N_20692,N_20596,N_20571);
nor U20693 (N_20693,N_20499,N_20552);
nor U20694 (N_20694,N_20533,N_20497);
and U20695 (N_20695,N_20589,N_20435);
and U20696 (N_20696,N_20536,N_20545);
and U20697 (N_20697,N_20472,N_20437);
xor U20698 (N_20698,N_20592,N_20568);
or U20699 (N_20699,N_20569,N_20517);
or U20700 (N_20700,N_20430,N_20543);
and U20701 (N_20701,N_20552,N_20419);
nor U20702 (N_20702,N_20408,N_20448);
or U20703 (N_20703,N_20486,N_20599);
and U20704 (N_20704,N_20496,N_20472);
nor U20705 (N_20705,N_20404,N_20587);
nand U20706 (N_20706,N_20571,N_20423);
nand U20707 (N_20707,N_20570,N_20548);
nor U20708 (N_20708,N_20503,N_20559);
and U20709 (N_20709,N_20565,N_20466);
nor U20710 (N_20710,N_20578,N_20575);
xnor U20711 (N_20711,N_20418,N_20425);
nand U20712 (N_20712,N_20515,N_20424);
and U20713 (N_20713,N_20486,N_20480);
nand U20714 (N_20714,N_20575,N_20471);
and U20715 (N_20715,N_20416,N_20573);
nor U20716 (N_20716,N_20578,N_20550);
or U20717 (N_20717,N_20439,N_20599);
or U20718 (N_20718,N_20508,N_20558);
or U20719 (N_20719,N_20566,N_20504);
or U20720 (N_20720,N_20557,N_20583);
or U20721 (N_20721,N_20502,N_20448);
or U20722 (N_20722,N_20566,N_20583);
or U20723 (N_20723,N_20454,N_20472);
and U20724 (N_20724,N_20471,N_20454);
xor U20725 (N_20725,N_20458,N_20544);
and U20726 (N_20726,N_20494,N_20510);
and U20727 (N_20727,N_20463,N_20432);
xnor U20728 (N_20728,N_20450,N_20593);
or U20729 (N_20729,N_20450,N_20402);
nor U20730 (N_20730,N_20563,N_20494);
nand U20731 (N_20731,N_20426,N_20534);
nand U20732 (N_20732,N_20485,N_20594);
nor U20733 (N_20733,N_20530,N_20513);
nand U20734 (N_20734,N_20409,N_20563);
or U20735 (N_20735,N_20539,N_20557);
or U20736 (N_20736,N_20535,N_20568);
or U20737 (N_20737,N_20549,N_20460);
xnor U20738 (N_20738,N_20439,N_20510);
and U20739 (N_20739,N_20558,N_20406);
nor U20740 (N_20740,N_20582,N_20529);
nor U20741 (N_20741,N_20427,N_20551);
xnor U20742 (N_20742,N_20544,N_20437);
and U20743 (N_20743,N_20531,N_20559);
nand U20744 (N_20744,N_20529,N_20478);
or U20745 (N_20745,N_20408,N_20512);
and U20746 (N_20746,N_20582,N_20579);
nand U20747 (N_20747,N_20485,N_20512);
nor U20748 (N_20748,N_20474,N_20461);
and U20749 (N_20749,N_20559,N_20572);
nand U20750 (N_20750,N_20472,N_20474);
nand U20751 (N_20751,N_20443,N_20415);
nand U20752 (N_20752,N_20482,N_20413);
nand U20753 (N_20753,N_20414,N_20592);
nand U20754 (N_20754,N_20561,N_20427);
or U20755 (N_20755,N_20581,N_20473);
or U20756 (N_20756,N_20552,N_20437);
nand U20757 (N_20757,N_20505,N_20460);
nor U20758 (N_20758,N_20532,N_20400);
nor U20759 (N_20759,N_20467,N_20459);
and U20760 (N_20760,N_20539,N_20556);
or U20761 (N_20761,N_20526,N_20425);
nor U20762 (N_20762,N_20545,N_20435);
or U20763 (N_20763,N_20471,N_20558);
nor U20764 (N_20764,N_20405,N_20452);
nand U20765 (N_20765,N_20433,N_20443);
and U20766 (N_20766,N_20514,N_20470);
nor U20767 (N_20767,N_20573,N_20536);
nor U20768 (N_20768,N_20532,N_20423);
nor U20769 (N_20769,N_20573,N_20524);
nor U20770 (N_20770,N_20488,N_20403);
nand U20771 (N_20771,N_20453,N_20406);
and U20772 (N_20772,N_20542,N_20549);
or U20773 (N_20773,N_20558,N_20556);
and U20774 (N_20774,N_20447,N_20456);
nor U20775 (N_20775,N_20564,N_20473);
nor U20776 (N_20776,N_20408,N_20545);
and U20777 (N_20777,N_20527,N_20471);
and U20778 (N_20778,N_20538,N_20483);
nor U20779 (N_20779,N_20436,N_20496);
and U20780 (N_20780,N_20503,N_20548);
and U20781 (N_20781,N_20594,N_20428);
and U20782 (N_20782,N_20561,N_20538);
nand U20783 (N_20783,N_20524,N_20489);
nor U20784 (N_20784,N_20563,N_20493);
xnor U20785 (N_20785,N_20557,N_20568);
nor U20786 (N_20786,N_20432,N_20577);
and U20787 (N_20787,N_20406,N_20438);
or U20788 (N_20788,N_20482,N_20502);
and U20789 (N_20789,N_20414,N_20585);
or U20790 (N_20790,N_20441,N_20414);
and U20791 (N_20791,N_20530,N_20508);
nand U20792 (N_20792,N_20436,N_20536);
nand U20793 (N_20793,N_20416,N_20499);
and U20794 (N_20794,N_20517,N_20448);
nand U20795 (N_20795,N_20479,N_20459);
or U20796 (N_20796,N_20493,N_20479);
nor U20797 (N_20797,N_20460,N_20419);
xnor U20798 (N_20798,N_20464,N_20435);
and U20799 (N_20799,N_20490,N_20578);
nand U20800 (N_20800,N_20623,N_20794);
and U20801 (N_20801,N_20672,N_20726);
nor U20802 (N_20802,N_20636,N_20729);
nand U20803 (N_20803,N_20741,N_20717);
nand U20804 (N_20804,N_20724,N_20638);
nor U20805 (N_20805,N_20632,N_20604);
nor U20806 (N_20806,N_20670,N_20754);
nand U20807 (N_20807,N_20669,N_20748);
nor U20808 (N_20808,N_20785,N_20613);
and U20809 (N_20809,N_20781,N_20706);
xnor U20810 (N_20810,N_20647,N_20736);
or U20811 (N_20811,N_20648,N_20772);
or U20812 (N_20812,N_20753,N_20642);
and U20813 (N_20813,N_20611,N_20789);
nand U20814 (N_20814,N_20628,N_20619);
nand U20815 (N_20815,N_20610,N_20652);
and U20816 (N_20816,N_20650,N_20627);
nor U20817 (N_20817,N_20682,N_20693);
and U20818 (N_20818,N_20764,N_20665);
and U20819 (N_20819,N_20637,N_20783);
xor U20820 (N_20820,N_20631,N_20600);
or U20821 (N_20821,N_20723,N_20713);
or U20822 (N_20822,N_20784,N_20630);
nand U20823 (N_20823,N_20714,N_20700);
nor U20824 (N_20824,N_20734,N_20721);
nor U20825 (N_20825,N_20653,N_20733);
nand U20826 (N_20826,N_20707,N_20779);
xnor U20827 (N_20827,N_20656,N_20678);
xnor U20828 (N_20828,N_20601,N_20743);
or U20829 (N_20829,N_20758,N_20715);
nand U20830 (N_20830,N_20688,N_20645);
and U20831 (N_20831,N_20719,N_20657);
or U20832 (N_20832,N_20641,N_20718);
and U20833 (N_20833,N_20649,N_20658);
nand U20834 (N_20834,N_20716,N_20740);
nand U20835 (N_20835,N_20643,N_20692);
or U20836 (N_20836,N_20676,N_20771);
and U20837 (N_20837,N_20798,N_20680);
nor U20838 (N_20838,N_20755,N_20703);
and U20839 (N_20839,N_20756,N_20775);
or U20840 (N_20840,N_20752,N_20727);
and U20841 (N_20841,N_20691,N_20728);
and U20842 (N_20842,N_20732,N_20749);
nand U20843 (N_20843,N_20773,N_20762);
xnor U20844 (N_20844,N_20739,N_20710);
nor U20845 (N_20845,N_20757,N_20704);
nand U20846 (N_20846,N_20639,N_20709);
or U20847 (N_20847,N_20626,N_20770);
and U20848 (N_20848,N_20694,N_20644);
or U20849 (N_20849,N_20763,N_20602);
nor U20850 (N_20850,N_20786,N_20609);
and U20851 (N_20851,N_20792,N_20659);
nor U20852 (N_20852,N_20702,N_20618);
xnor U20853 (N_20853,N_20685,N_20765);
nor U20854 (N_20854,N_20747,N_20606);
xnor U20855 (N_20855,N_20769,N_20625);
nand U20856 (N_20856,N_20614,N_20663);
or U20857 (N_20857,N_20788,N_20684);
or U20858 (N_20858,N_20696,N_20689);
nand U20859 (N_20859,N_20686,N_20687);
and U20860 (N_20860,N_20745,N_20651);
nor U20861 (N_20861,N_20607,N_20738);
xor U20862 (N_20862,N_20760,N_20620);
or U20863 (N_20863,N_20712,N_20622);
nor U20864 (N_20864,N_20675,N_20612);
and U20865 (N_20865,N_20624,N_20795);
nand U20866 (N_20866,N_20660,N_20793);
or U20867 (N_20867,N_20616,N_20671);
xnor U20868 (N_20868,N_20698,N_20635);
and U20869 (N_20869,N_20662,N_20797);
or U20870 (N_20870,N_20668,N_20667);
or U20871 (N_20871,N_20787,N_20750);
and U20872 (N_20872,N_20778,N_20646);
or U20873 (N_20873,N_20796,N_20681);
and U20874 (N_20874,N_20776,N_20720);
nand U20875 (N_20875,N_20655,N_20701);
or U20876 (N_20876,N_20791,N_20799);
nand U20877 (N_20877,N_20677,N_20654);
xor U20878 (N_20878,N_20708,N_20780);
nand U20879 (N_20879,N_20633,N_20705);
xnor U20880 (N_20880,N_20767,N_20777);
or U20881 (N_20881,N_20766,N_20774);
and U20882 (N_20882,N_20615,N_20751);
nand U20883 (N_20883,N_20666,N_20674);
or U20884 (N_20884,N_20768,N_20759);
or U20885 (N_20885,N_20725,N_20731);
nand U20886 (N_20886,N_20679,N_20735);
xnor U20887 (N_20887,N_20617,N_20640);
nor U20888 (N_20888,N_20664,N_20690);
xor U20889 (N_20889,N_20730,N_20742);
nor U20890 (N_20890,N_20673,N_20761);
nor U20891 (N_20891,N_20629,N_20790);
nor U20892 (N_20892,N_20695,N_20683);
nand U20893 (N_20893,N_20697,N_20737);
and U20894 (N_20894,N_20722,N_20608);
and U20895 (N_20895,N_20744,N_20782);
and U20896 (N_20896,N_20661,N_20634);
xor U20897 (N_20897,N_20621,N_20711);
and U20898 (N_20898,N_20699,N_20603);
nand U20899 (N_20899,N_20746,N_20605);
nor U20900 (N_20900,N_20739,N_20676);
xnor U20901 (N_20901,N_20624,N_20619);
nor U20902 (N_20902,N_20629,N_20613);
or U20903 (N_20903,N_20607,N_20625);
xnor U20904 (N_20904,N_20619,N_20643);
and U20905 (N_20905,N_20708,N_20701);
or U20906 (N_20906,N_20697,N_20676);
and U20907 (N_20907,N_20759,N_20683);
and U20908 (N_20908,N_20643,N_20730);
nor U20909 (N_20909,N_20694,N_20756);
nor U20910 (N_20910,N_20629,N_20795);
and U20911 (N_20911,N_20661,N_20648);
nand U20912 (N_20912,N_20691,N_20649);
or U20913 (N_20913,N_20641,N_20673);
nor U20914 (N_20914,N_20741,N_20650);
or U20915 (N_20915,N_20717,N_20663);
xnor U20916 (N_20916,N_20717,N_20615);
nand U20917 (N_20917,N_20732,N_20639);
and U20918 (N_20918,N_20624,N_20647);
and U20919 (N_20919,N_20621,N_20721);
or U20920 (N_20920,N_20662,N_20728);
nor U20921 (N_20921,N_20727,N_20610);
nand U20922 (N_20922,N_20646,N_20754);
and U20923 (N_20923,N_20725,N_20713);
nor U20924 (N_20924,N_20617,N_20719);
and U20925 (N_20925,N_20616,N_20614);
and U20926 (N_20926,N_20707,N_20700);
or U20927 (N_20927,N_20733,N_20641);
nand U20928 (N_20928,N_20674,N_20729);
nor U20929 (N_20929,N_20600,N_20736);
and U20930 (N_20930,N_20723,N_20761);
or U20931 (N_20931,N_20735,N_20777);
nor U20932 (N_20932,N_20615,N_20732);
nor U20933 (N_20933,N_20744,N_20778);
and U20934 (N_20934,N_20667,N_20729);
and U20935 (N_20935,N_20639,N_20608);
or U20936 (N_20936,N_20661,N_20785);
and U20937 (N_20937,N_20729,N_20615);
nand U20938 (N_20938,N_20787,N_20700);
and U20939 (N_20939,N_20695,N_20770);
and U20940 (N_20940,N_20752,N_20707);
nor U20941 (N_20941,N_20747,N_20685);
or U20942 (N_20942,N_20666,N_20750);
xnor U20943 (N_20943,N_20621,N_20708);
nand U20944 (N_20944,N_20652,N_20721);
nor U20945 (N_20945,N_20745,N_20627);
and U20946 (N_20946,N_20765,N_20669);
nor U20947 (N_20947,N_20764,N_20615);
nor U20948 (N_20948,N_20719,N_20668);
or U20949 (N_20949,N_20723,N_20687);
xor U20950 (N_20950,N_20767,N_20782);
xnor U20951 (N_20951,N_20653,N_20784);
or U20952 (N_20952,N_20783,N_20676);
xor U20953 (N_20953,N_20756,N_20674);
and U20954 (N_20954,N_20737,N_20752);
or U20955 (N_20955,N_20734,N_20733);
and U20956 (N_20956,N_20730,N_20662);
and U20957 (N_20957,N_20665,N_20796);
or U20958 (N_20958,N_20792,N_20764);
or U20959 (N_20959,N_20601,N_20798);
nand U20960 (N_20960,N_20621,N_20736);
or U20961 (N_20961,N_20754,N_20600);
nor U20962 (N_20962,N_20670,N_20764);
and U20963 (N_20963,N_20614,N_20783);
nor U20964 (N_20964,N_20690,N_20760);
nand U20965 (N_20965,N_20741,N_20633);
xnor U20966 (N_20966,N_20633,N_20711);
or U20967 (N_20967,N_20755,N_20796);
nand U20968 (N_20968,N_20677,N_20611);
or U20969 (N_20969,N_20619,N_20720);
nand U20970 (N_20970,N_20797,N_20666);
and U20971 (N_20971,N_20764,N_20647);
nor U20972 (N_20972,N_20739,N_20701);
nand U20973 (N_20973,N_20768,N_20719);
nor U20974 (N_20974,N_20774,N_20671);
or U20975 (N_20975,N_20729,N_20785);
nor U20976 (N_20976,N_20646,N_20725);
xnor U20977 (N_20977,N_20683,N_20622);
or U20978 (N_20978,N_20675,N_20611);
and U20979 (N_20979,N_20601,N_20707);
or U20980 (N_20980,N_20714,N_20602);
nand U20981 (N_20981,N_20652,N_20702);
nor U20982 (N_20982,N_20726,N_20723);
nor U20983 (N_20983,N_20760,N_20636);
nor U20984 (N_20984,N_20798,N_20725);
xnor U20985 (N_20985,N_20624,N_20699);
or U20986 (N_20986,N_20706,N_20626);
or U20987 (N_20987,N_20757,N_20660);
and U20988 (N_20988,N_20705,N_20700);
nand U20989 (N_20989,N_20721,N_20641);
nor U20990 (N_20990,N_20646,N_20724);
nor U20991 (N_20991,N_20773,N_20638);
nand U20992 (N_20992,N_20775,N_20728);
nand U20993 (N_20993,N_20657,N_20611);
nand U20994 (N_20994,N_20786,N_20682);
or U20995 (N_20995,N_20619,N_20609);
nor U20996 (N_20996,N_20751,N_20734);
or U20997 (N_20997,N_20726,N_20757);
nor U20998 (N_20998,N_20759,N_20716);
nand U20999 (N_20999,N_20668,N_20695);
and U21000 (N_21000,N_20935,N_20907);
and U21001 (N_21001,N_20848,N_20997);
nor U21002 (N_21002,N_20849,N_20931);
or U21003 (N_21003,N_20853,N_20828);
and U21004 (N_21004,N_20917,N_20948);
nor U21005 (N_21005,N_20830,N_20898);
or U21006 (N_21006,N_20987,N_20862);
nor U21007 (N_21007,N_20805,N_20906);
nor U21008 (N_21008,N_20964,N_20866);
nand U21009 (N_21009,N_20899,N_20944);
xnor U21010 (N_21010,N_20963,N_20863);
nand U21011 (N_21011,N_20980,N_20909);
nor U21012 (N_21012,N_20842,N_20843);
nor U21013 (N_21013,N_20834,N_20873);
or U21014 (N_21014,N_20816,N_20946);
nor U21015 (N_21015,N_20810,N_20923);
or U21016 (N_21016,N_20954,N_20823);
nand U21017 (N_21017,N_20820,N_20845);
xor U21018 (N_21018,N_20975,N_20856);
nand U21019 (N_21019,N_20970,N_20983);
nor U21020 (N_21020,N_20950,N_20832);
xor U21021 (N_21021,N_20920,N_20939);
or U21022 (N_21022,N_20959,N_20851);
or U21023 (N_21023,N_20807,N_20951);
nor U21024 (N_21024,N_20955,N_20903);
and U21025 (N_21025,N_20883,N_20837);
nand U21026 (N_21026,N_20850,N_20818);
and U21027 (N_21027,N_20982,N_20870);
nor U21028 (N_21028,N_20803,N_20952);
nor U21029 (N_21029,N_20960,N_20932);
or U21030 (N_21030,N_20990,N_20804);
nor U21031 (N_21031,N_20992,N_20840);
xor U21032 (N_21032,N_20922,N_20918);
and U21033 (N_21033,N_20874,N_20938);
nor U21034 (N_21034,N_20864,N_20949);
and U21035 (N_21035,N_20976,N_20839);
and U21036 (N_21036,N_20915,N_20854);
or U21037 (N_21037,N_20936,N_20912);
xnor U21038 (N_21038,N_20927,N_20968);
or U21039 (N_21039,N_20835,N_20809);
nand U21040 (N_21040,N_20994,N_20928);
nand U21041 (N_21041,N_20973,N_20985);
and U21042 (N_21042,N_20967,N_20806);
or U21043 (N_21043,N_20800,N_20861);
nor U21044 (N_21044,N_20897,N_20913);
or U21045 (N_21045,N_20888,N_20978);
or U21046 (N_21046,N_20865,N_20890);
xnor U21047 (N_21047,N_20930,N_20858);
and U21048 (N_21048,N_20958,N_20855);
or U21049 (N_21049,N_20872,N_20817);
xnor U21050 (N_21050,N_20965,N_20943);
nand U21051 (N_21051,N_20884,N_20940);
nor U21052 (N_21052,N_20847,N_20894);
and U21053 (N_21053,N_20891,N_20801);
and U21054 (N_21054,N_20981,N_20972);
or U21055 (N_21055,N_20900,N_20838);
and U21056 (N_21056,N_20814,N_20867);
or U21057 (N_21057,N_20869,N_20896);
or U21058 (N_21058,N_20941,N_20986);
xnor U21059 (N_21059,N_20825,N_20821);
or U21060 (N_21060,N_20945,N_20878);
xnor U21061 (N_21061,N_20886,N_20859);
and U21062 (N_21062,N_20905,N_20881);
nand U21063 (N_21063,N_20984,N_20880);
and U21064 (N_21064,N_20877,N_20902);
or U21065 (N_21065,N_20876,N_20813);
and U21066 (N_21066,N_20947,N_20824);
and U21067 (N_21067,N_20827,N_20901);
and U21068 (N_21068,N_20921,N_20819);
and U21069 (N_21069,N_20996,N_20860);
nand U21070 (N_21070,N_20889,N_20893);
and U21071 (N_21071,N_20942,N_20882);
and U21072 (N_21072,N_20826,N_20841);
nor U21073 (N_21073,N_20995,N_20892);
or U21074 (N_21074,N_20887,N_20929);
or U21075 (N_21075,N_20904,N_20993);
or U21076 (N_21076,N_20811,N_20979);
nand U21077 (N_21077,N_20871,N_20895);
or U21078 (N_21078,N_20991,N_20971);
xnor U21079 (N_21079,N_20808,N_20988);
nand U21080 (N_21080,N_20914,N_20961);
nand U21081 (N_21081,N_20911,N_20836);
and U21082 (N_21082,N_20933,N_20974);
or U21083 (N_21083,N_20857,N_20868);
nand U21084 (N_21084,N_20962,N_20956);
nand U21085 (N_21085,N_20846,N_20926);
and U21086 (N_21086,N_20916,N_20812);
nor U21087 (N_21087,N_20802,N_20885);
or U21088 (N_21088,N_20815,N_20833);
and U21089 (N_21089,N_20875,N_20822);
or U21090 (N_21090,N_20989,N_20844);
and U21091 (N_21091,N_20831,N_20953);
and U21092 (N_21092,N_20879,N_20998);
nor U21093 (N_21093,N_20934,N_20829);
or U21094 (N_21094,N_20966,N_20924);
or U21095 (N_21095,N_20908,N_20969);
nor U21096 (N_21096,N_20937,N_20925);
and U21097 (N_21097,N_20957,N_20999);
or U21098 (N_21098,N_20919,N_20910);
or U21099 (N_21099,N_20852,N_20977);
xnor U21100 (N_21100,N_20868,N_20903);
nand U21101 (N_21101,N_20866,N_20863);
nand U21102 (N_21102,N_20824,N_20800);
nand U21103 (N_21103,N_20861,N_20915);
and U21104 (N_21104,N_20830,N_20905);
and U21105 (N_21105,N_20803,N_20846);
nor U21106 (N_21106,N_20863,N_20937);
nor U21107 (N_21107,N_20957,N_20841);
nand U21108 (N_21108,N_20882,N_20895);
nand U21109 (N_21109,N_20832,N_20817);
nand U21110 (N_21110,N_20919,N_20893);
xnor U21111 (N_21111,N_20942,N_20834);
nand U21112 (N_21112,N_20916,N_20800);
and U21113 (N_21113,N_20901,N_20824);
nand U21114 (N_21114,N_20926,N_20858);
or U21115 (N_21115,N_20841,N_20807);
or U21116 (N_21116,N_20989,N_20923);
nor U21117 (N_21117,N_20849,N_20884);
nand U21118 (N_21118,N_20874,N_20800);
nand U21119 (N_21119,N_20889,N_20861);
xnor U21120 (N_21120,N_20836,N_20818);
and U21121 (N_21121,N_20962,N_20805);
nor U21122 (N_21122,N_20804,N_20981);
xnor U21123 (N_21123,N_20968,N_20978);
or U21124 (N_21124,N_20947,N_20861);
nand U21125 (N_21125,N_20963,N_20966);
xor U21126 (N_21126,N_20976,N_20881);
or U21127 (N_21127,N_20948,N_20806);
or U21128 (N_21128,N_20970,N_20977);
or U21129 (N_21129,N_20965,N_20994);
nor U21130 (N_21130,N_20968,N_20848);
or U21131 (N_21131,N_20871,N_20993);
and U21132 (N_21132,N_20801,N_20809);
nand U21133 (N_21133,N_20847,N_20987);
nor U21134 (N_21134,N_20925,N_20919);
nand U21135 (N_21135,N_20907,N_20941);
nand U21136 (N_21136,N_20855,N_20847);
and U21137 (N_21137,N_20990,N_20855);
or U21138 (N_21138,N_20998,N_20852);
nor U21139 (N_21139,N_20858,N_20933);
nand U21140 (N_21140,N_20840,N_20847);
nor U21141 (N_21141,N_20903,N_20960);
and U21142 (N_21142,N_20941,N_20817);
and U21143 (N_21143,N_20873,N_20800);
nand U21144 (N_21144,N_20806,N_20950);
nand U21145 (N_21145,N_20997,N_20801);
nand U21146 (N_21146,N_20802,N_20954);
and U21147 (N_21147,N_20807,N_20849);
nor U21148 (N_21148,N_20860,N_20849);
or U21149 (N_21149,N_20823,N_20904);
or U21150 (N_21150,N_20818,N_20960);
or U21151 (N_21151,N_20878,N_20857);
nand U21152 (N_21152,N_20907,N_20804);
nand U21153 (N_21153,N_20839,N_20822);
or U21154 (N_21154,N_20900,N_20877);
or U21155 (N_21155,N_20882,N_20957);
and U21156 (N_21156,N_20901,N_20971);
nor U21157 (N_21157,N_20859,N_20942);
and U21158 (N_21158,N_20981,N_20848);
or U21159 (N_21159,N_20800,N_20950);
nand U21160 (N_21160,N_20935,N_20908);
and U21161 (N_21161,N_20909,N_20845);
nor U21162 (N_21162,N_20934,N_20835);
nor U21163 (N_21163,N_20976,N_20865);
nor U21164 (N_21164,N_20933,N_20948);
or U21165 (N_21165,N_20817,N_20873);
nand U21166 (N_21166,N_20864,N_20931);
and U21167 (N_21167,N_20870,N_20979);
or U21168 (N_21168,N_20953,N_20978);
xnor U21169 (N_21169,N_20910,N_20982);
and U21170 (N_21170,N_20990,N_20828);
nor U21171 (N_21171,N_20851,N_20876);
nor U21172 (N_21172,N_20909,N_20916);
nand U21173 (N_21173,N_20887,N_20840);
xor U21174 (N_21174,N_20979,N_20938);
nand U21175 (N_21175,N_20935,N_20970);
xor U21176 (N_21176,N_20873,N_20908);
nor U21177 (N_21177,N_20940,N_20919);
xnor U21178 (N_21178,N_20930,N_20908);
and U21179 (N_21179,N_20902,N_20907);
nand U21180 (N_21180,N_20956,N_20990);
nor U21181 (N_21181,N_20835,N_20961);
nor U21182 (N_21182,N_20890,N_20926);
nand U21183 (N_21183,N_20876,N_20814);
or U21184 (N_21184,N_20831,N_20922);
or U21185 (N_21185,N_20814,N_20941);
nand U21186 (N_21186,N_20939,N_20942);
or U21187 (N_21187,N_20875,N_20884);
or U21188 (N_21188,N_20833,N_20827);
nand U21189 (N_21189,N_20833,N_20957);
or U21190 (N_21190,N_20942,N_20853);
nor U21191 (N_21191,N_20936,N_20851);
nor U21192 (N_21192,N_20805,N_20839);
nand U21193 (N_21193,N_20933,N_20819);
nand U21194 (N_21194,N_20823,N_20955);
or U21195 (N_21195,N_20811,N_20986);
or U21196 (N_21196,N_20907,N_20985);
and U21197 (N_21197,N_20836,N_20889);
xor U21198 (N_21198,N_20972,N_20857);
xnor U21199 (N_21199,N_20983,N_20989);
and U21200 (N_21200,N_21166,N_21144);
nand U21201 (N_21201,N_21161,N_21014);
or U21202 (N_21202,N_21185,N_21124);
or U21203 (N_21203,N_21069,N_21138);
nand U21204 (N_21204,N_21007,N_21061);
and U21205 (N_21205,N_21075,N_21157);
and U21206 (N_21206,N_21164,N_21184);
nor U21207 (N_21207,N_21002,N_21199);
nand U21208 (N_21208,N_21143,N_21165);
nand U21209 (N_21209,N_21171,N_21162);
and U21210 (N_21210,N_21085,N_21175);
or U21211 (N_21211,N_21054,N_21105);
or U21212 (N_21212,N_21088,N_21020);
or U21213 (N_21213,N_21029,N_21056);
and U21214 (N_21214,N_21120,N_21083);
or U21215 (N_21215,N_21090,N_21052);
nand U21216 (N_21216,N_21129,N_21047);
or U21217 (N_21217,N_21084,N_21167);
nand U21218 (N_21218,N_21113,N_21177);
nand U21219 (N_21219,N_21114,N_21180);
nand U21220 (N_21220,N_21102,N_21022);
nand U21221 (N_21221,N_21132,N_21033);
or U21222 (N_21222,N_21041,N_21034);
nand U21223 (N_21223,N_21019,N_21096);
nand U21224 (N_21224,N_21195,N_21013);
and U21225 (N_21225,N_21178,N_21038);
nor U21226 (N_21226,N_21112,N_21080);
nand U21227 (N_21227,N_21156,N_21035);
and U21228 (N_21228,N_21150,N_21118);
nor U21229 (N_21229,N_21133,N_21123);
or U21230 (N_21230,N_21160,N_21037);
nand U21231 (N_21231,N_21082,N_21070);
nor U21232 (N_21232,N_21072,N_21107);
nand U21233 (N_21233,N_21023,N_21091);
or U21234 (N_21234,N_21001,N_21170);
and U21235 (N_21235,N_21187,N_21101);
nand U21236 (N_21236,N_21174,N_21018);
or U21237 (N_21237,N_21191,N_21000);
nand U21238 (N_21238,N_21030,N_21087);
or U21239 (N_21239,N_21057,N_21098);
xnor U21240 (N_21240,N_21094,N_21086);
and U21241 (N_21241,N_21004,N_21006);
or U21242 (N_21242,N_21142,N_21039);
xnor U21243 (N_21243,N_21042,N_21134);
nand U21244 (N_21244,N_21103,N_21027);
nor U21245 (N_21245,N_21089,N_21078);
or U21246 (N_21246,N_21032,N_21139);
or U21247 (N_21247,N_21140,N_21062);
or U21248 (N_21248,N_21067,N_21108);
nor U21249 (N_21249,N_21110,N_21192);
or U21250 (N_21250,N_21106,N_21193);
nand U21251 (N_21251,N_21076,N_21026);
xor U21252 (N_21252,N_21116,N_21189);
nand U21253 (N_21253,N_21126,N_21117);
or U21254 (N_21254,N_21173,N_21043);
nor U21255 (N_21255,N_21121,N_21073);
nor U21256 (N_21256,N_21127,N_21050);
nand U21257 (N_21257,N_21168,N_21115);
or U21258 (N_21258,N_21131,N_21016);
or U21259 (N_21259,N_21136,N_21148);
nor U21260 (N_21260,N_21053,N_21151);
nor U21261 (N_21261,N_21104,N_21141);
nand U21262 (N_21262,N_21152,N_21181);
or U21263 (N_21263,N_21111,N_21172);
or U21264 (N_21264,N_21074,N_21119);
nor U21265 (N_21265,N_21099,N_21068);
nand U21266 (N_21266,N_21147,N_21017);
nand U21267 (N_21267,N_21010,N_21066);
nand U21268 (N_21268,N_21065,N_21155);
and U21269 (N_21269,N_21122,N_21182);
or U21270 (N_21270,N_21130,N_21146);
nor U21271 (N_21271,N_21100,N_21028);
or U21272 (N_21272,N_21186,N_21158);
nand U21273 (N_21273,N_21021,N_21009);
nand U21274 (N_21274,N_21079,N_21071);
nand U21275 (N_21275,N_21059,N_21149);
xor U21276 (N_21276,N_21025,N_21163);
and U21277 (N_21277,N_21024,N_21109);
nand U21278 (N_21278,N_21188,N_21169);
nor U21279 (N_21279,N_21049,N_21092);
nor U21280 (N_21280,N_21055,N_21183);
nand U21281 (N_21281,N_21011,N_21058);
and U21282 (N_21282,N_21077,N_21051);
nand U21283 (N_21283,N_21125,N_21179);
nand U21284 (N_21284,N_21154,N_21003);
and U21285 (N_21285,N_21012,N_21008);
nand U21286 (N_21286,N_21093,N_21045);
nand U21287 (N_21287,N_21194,N_21031);
nor U21288 (N_21288,N_21081,N_21005);
xor U21289 (N_21289,N_21060,N_21159);
nor U21290 (N_21290,N_21196,N_21048);
nand U21291 (N_21291,N_21097,N_21197);
nand U21292 (N_21292,N_21046,N_21198);
or U21293 (N_21293,N_21145,N_21015);
nor U21294 (N_21294,N_21153,N_21040);
xnor U21295 (N_21295,N_21063,N_21064);
xnor U21296 (N_21296,N_21135,N_21044);
or U21297 (N_21297,N_21095,N_21176);
nor U21298 (N_21298,N_21128,N_21137);
or U21299 (N_21299,N_21190,N_21036);
or U21300 (N_21300,N_21011,N_21192);
nand U21301 (N_21301,N_21047,N_21083);
or U21302 (N_21302,N_21040,N_21038);
or U21303 (N_21303,N_21042,N_21044);
and U21304 (N_21304,N_21162,N_21137);
xor U21305 (N_21305,N_21053,N_21069);
and U21306 (N_21306,N_21166,N_21123);
xnor U21307 (N_21307,N_21086,N_21095);
xnor U21308 (N_21308,N_21125,N_21191);
xor U21309 (N_21309,N_21047,N_21169);
nand U21310 (N_21310,N_21110,N_21141);
nand U21311 (N_21311,N_21101,N_21004);
or U21312 (N_21312,N_21187,N_21048);
nor U21313 (N_21313,N_21075,N_21058);
and U21314 (N_21314,N_21192,N_21102);
nand U21315 (N_21315,N_21193,N_21111);
nand U21316 (N_21316,N_21073,N_21042);
xor U21317 (N_21317,N_21113,N_21135);
nand U21318 (N_21318,N_21141,N_21151);
and U21319 (N_21319,N_21086,N_21124);
nor U21320 (N_21320,N_21124,N_21013);
and U21321 (N_21321,N_21072,N_21059);
and U21322 (N_21322,N_21096,N_21181);
xor U21323 (N_21323,N_21042,N_21103);
xnor U21324 (N_21324,N_21134,N_21081);
nor U21325 (N_21325,N_21069,N_21159);
nor U21326 (N_21326,N_21155,N_21041);
nand U21327 (N_21327,N_21150,N_21037);
xor U21328 (N_21328,N_21000,N_21018);
nand U21329 (N_21329,N_21166,N_21161);
nor U21330 (N_21330,N_21043,N_21070);
or U21331 (N_21331,N_21066,N_21031);
nand U21332 (N_21332,N_21050,N_21054);
and U21333 (N_21333,N_21176,N_21087);
or U21334 (N_21334,N_21189,N_21161);
xor U21335 (N_21335,N_21073,N_21017);
nor U21336 (N_21336,N_21173,N_21015);
and U21337 (N_21337,N_21081,N_21186);
nand U21338 (N_21338,N_21073,N_21144);
nor U21339 (N_21339,N_21181,N_21061);
and U21340 (N_21340,N_21058,N_21112);
or U21341 (N_21341,N_21054,N_21009);
xnor U21342 (N_21342,N_21044,N_21148);
or U21343 (N_21343,N_21041,N_21016);
nand U21344 (N_21344,N_21087,N_21174);
or U21345 (N_21345,N_21004,N_21091);
and U21346 (N_21346,N_21098,N_21190);
or U21347 (N_21347,N_21103,N_21193);
and U21348 (N_21348,N_21030,N_21192);
nor U21349 (N_21349,N_21096,N_21156);
nor U21350 (N_21350,N_21124,N_21171);
nand U21351 (N_21351,N_21039,N_21170);
and U21352 (N_21352,N_21060,N_21122);
and U21353 (N_21353,N_21051,N_21012);
and U21354 (N_21354,N_21064,N_21145);
nand U21355 (N_21355,N_21133,N_21187);
nand U21356 (N_21356,N_21143,N_21112);
and U21357 (N_21357,N_21141,N_21094);
nor U21358 (N_21358,N_21168,N_21017);
nor U21359 (N_21359,N_21087,N_21120);
nand U21360 (N_21360,N_21068,N_21065);
or U21361 (N_21361,N_21044,N_21131);
or U21362 (N_21362,N_21129,N_21161);
and U21363 (N_21363,N_21096,N_21058);
nand U21364 (N_21364,N_21140,N_21141);
nor U21365 (N_21365,N_21103,N_21107);
nand U21366 (N_21366,N_21002,N_21192);
or U21367 (N_21367,N_21059,N_21028);
nand U21368 (N_21368,N_21073,N_21160);
nor U21369 (N_21369,N_21135,N_21007);
xnor U21370 (N_21370,N_21152,N_21189);
nand U21371 (N_21371,N_21001,N_21046);
or U21372 (N_21372,N_21116,N_21070);
nand U21373 (N_21373,N_21041,N_21015);
or U21374 (N_21374,N_21044,N_21030);
or U21375 (N_21375,N_21100,N_21043);
xor U21376 (N_21376,N_21040,N_21072);
and U21377 (N_21377,N_21028,N_21020);
nand U21378 (N_21378,N_21053,N_21188);
xnor U21379 (N_21379,N_21165,N_21172);
or U21380 (N_21380,N_21048,N_21092);
nor U21381 (N_21381,N_21184,N_21091);
xor U21382 (N_21382,N_21088,N_21193);
or U21383 (N_21383,N_21191,N_21031);
or U21384 (N_21384,N_21144,N_21023);
nor U21385 (N_21385,N_21185,N_21140);
nand U21386 (N_21386,N_21155,N_21195);
or U21387 (N_21387,N_21047,N_21027);
and U21388 (N_21388,N_21019,N_21121);
xor U21389 (N_21389,N_21074,N_21149);
or U21390 (N_21390,N_21132,N_21171);
or U21391 (N_21391,N_21099,N_21155);
and U21392 (N_21392,N_21143,N_21188);
nor U21393 (N_21393,N_21191,N_21024);
or U21394 (N_21394,N_21082,N_21170);
nor U21395 (N_21395,N_21029,N_21168);
and U21396 (N_21396,N_21095,N_21045);
nand U21397 (N_21397,N_21158,N_21004);
xor U21398 (N_21398,N_21129,N_21144);
and U21399 (N_21399,N_21006,N_21137);
and U21400 (N_21400,N_21254,N_21268);
and U21401 (N_21401,N_21322,N_21262);
and U21402 (N_21402,N_21349,N_21247);
or U21403 (N_21403,N_21396,N_21320);
or U21404 (N_21404,N_21200,N_21248);
nor U21405 (N_21405,N_21227,N_21390);
nor U21406 (N_21406,N_21252,N_21359);
xnor U21407 (N_21407,N_21272,N_21371);
and U21408 (N_21408,N_21339,N_21365);
nand U21409 (N_21409,N_21281,N_21380);
and U21410 (N_21410,N_21259,N_21377);
nor U21411 (N_21411,N_21341,N_21274);
or U21412 (N_21412,N_21256,N_21271);
xor U21413 (N_21413,N_21354,N_21295);
nand U21414 (N_21414,N_21340,N_21279);
or U21415 (N_21415,N_21245,N_21324);
nor U21416 (N_21416,N_21361,N_21214);
nand U21417 (N_21417,N_21310,N_21229);
or U21418 (N_21418,N_21282,N_21211);
nor U21419 (N_21419,N_21373,N_21260);
nor U21420 (N_21420,N_21303,N_21216);
xor U21421 (N_21421,N_21238,N_21331);
nor U21422 (N_21422,N_21270,N_21207);
or U21423 (N_21423,N_21264,N_21394);
xnor U21424 (N_21424,N_21283,N_21358);
and U21425 (N_21425,N_21203,N_21383);
or U21426 (N_21426,N_21253,N_21378);
nor U21427 (N_21427,N_21315,N_21273);
nand U21428 (N_21428,N_21355,N_21343);
nand U21429 (N_21429,N_21250,N_21258);
nor U21430 (N_21430,N_21317,N_21255);
and U21431 (N_21431,N_21239,N_21392);
nand U21432 (N_21432,N_21266,N_21220);
nand U21433 (N_21433,N_21374,N_21219);
nand U21434 (N_21434,N_21313,N_21225);
nor U21435 (N_21435,N_21240,N_21232);
and U21436 (N_21436,N_21381,N_21399);
nor U21437 (N_21437,N_21210,N_21212);
nand U21438 (N_21438,N_21202,N_21265);
xnor U21439 (N_21439,N_21329,N_21337);
or U21440 (N_21440,N_21294,N_21382);
nand U21441 (N_21441,N_21209,N_21292);
xor U21442 (N_21442,N_21261,N_21226);
or U21443 (N_21443,N_21251,N_21336);
and U21444 (N_21444,N_21357,N_21328);
and U21445 (N_21445,N_21384,N_21376);
nand U21446 (N_21446,N_21241,N_21333);
and U21447 (N_21447,N_21368,N_21342);
nor U21448 (N_21448,N_21244,N_21284);
nand U21449 (N_21449,N_21301,N_21334);
and U21450 (N_21450,N_21335,N_21305);
and U21451 (N_21451,N_21224,N_21300);
and U21452 (N_21452,N_21293,N_21332);
and U21453 (N_21453,N_21298,N_21319);
nand U21454 (N_21454,N_21222,N_21296);
and U21455 (N_21455,N_21351,N_21348);
or U21456 (N_21456,N_21237,N_21280);
nand U21457 (N_21457,N_21326,N_21321);
or U21458 (N_21458,N_21364,N_21323);
nand U21459 (N_21459,N_21276,N_21217);
nor U21460 (N_21460,N_21388,N_21309);
and U21461 (N_21461,N_21263,N_21387);
and U21462 (N_21462,N_21314,N_21228);
xor U21463 (N_21463,N_21243,N_21330);
nor U21464 (N_21464,N_21308,N_21346);
or U21465 (N_21465,N_21291,N_21325);
and U21466 (N_21466,N_21230,N_21391);
or U21467 (N_21467,N_21393,N_21208);
nand U21468 (N_21468,N_21242,N_21246);
nand U21469 (N_21469,N_21362,N_21350);
and U21470 (N_21470,N_21356,N_21257);
xnor U21471 (N_21471,N_21277,N_21221);
nand U21472 (N_21472,N_21234,N_21344);
nor U21473 (N_21473,N_21318,N_21386);
or U21474 (N_21474,N_21345,N_21375);
xnor U21475 (N_21475,N_21360,N_21286);
or U21476 (N_21476,N_21206,N_21397);
or U21477 (N_21477,N_21347,N_21389);
xor U21478 (N_21478,N_21353,N_21299);
nand U21479 (N_21479,N_21288,N_21306);
nand U21480 (N_21480,N_21398,N_21352);
or U21481 (N_21481,N_21218,N_21302);
nand U21482 (N_21482,N_21312,N_21233);
nor U21483 (N_21483,N_21275,N_21213);
nor U21484 (N_21484,N_21297,N_21311);
xor U21485 (N_21485,N_21215,N_21304);
and U21486 (N_21486,N_21379,N_21223);
or U21487 (N_21487,N_21278,N_21363);
xnor U21488 (N_21488,N_21205,N_21269);
or U21489 (N_21489,N_21231,N_21372);
or U21490 (N_21490,N_21290,N_21204);
or U21491 (N_21491,N_21366,N_21338);
or U21492 (N_21492,N_21327,N_21267);
nor U21493 (N_21493,N_21236,N_21235);
nand U21494 (N_21494,N_21285,N_21385);
or U21495 (N_21495,N_21370,N_21289);
nor U21496 (N_21496,N_21307,N_21316);
or U21497 (N_21497,N_21249,N_21201);
and U21498 (N_21498,N_21395,N_21287);
nor U21499 (N_21499,N_21367,N_21369);
nor U21500 (N_21500,N_21272,N_21205);
or U21501 (N_21501,N_21255,N_21301);
nor U21502 (N_21502,N_21271,N_21269);
and U21503 (N_21503,N_21240,N_21236);
xor U21504 (N_21504,N_21224,N_21258);
or U21505 (N_21505,N_21330,N_21377);
and U21506 (N_21506,N_21236,N_21286);
or U21507 (N_21507,N_21387,N_21211);
xnor U21508 (N_21508,N_21387,N_21235);
or U21509 (N_21509,N_21301,N_21287);
nor U21510 (N_21510,N_21258,N_21237);
and U21511 (N_21511,N_21389,N_21309);
nand U21512 (N_21512,N_21292,N_21381);
or U21513 (N_21513,N_21308,N_21215);
nor U21514 (N_21514,N_21288,N_21256);
nor U21515 (N_21515,N_21321,N_21226);
or U21516 (N_21516,N_21395,N_21373);
or U21517 (N_21517,N_21203,N_21242);
and U21518 (N_21518,N_21259,N_21294);
nor U21519 (N_21519,N_21265,N_21393);
xnor U21520 (N_21520,N_21388,N_21297);
or U21521 (N_21521,N_21388,N_21281);
nor U21522 (N_21522,N_21225,N_21290);
nor U21523 (N_21523,N_21210,N_21292);
nand U21524 (N_21524,N_21274,N_21256);
nand U21525 (N_21525,N_21331,N_21317);
nor U21526 (N_21526,N_21230,N_21229);
or U21527 (N_21527,N_21253,N_21284);
xnor U21528 (N_21528,N_21308,N_21210);
and U21529 (N_21529,N_21334,N_21206);
or U21530 (N_21530,N_21276,N_21340);
and U21531 (N_21531,N_21291,N_21317);
and U21532 (N_21532,N_21319,N_21234);
nor U21533 (N_21533,N_21246,N_21315);
nand U21534 (N_21534,N_21326,N_21299);
and U21535 (N_21535,N_21244,N_21394);
and U21536 (N_21536,N_21318,N_21297);
and U21537 (N_21537,N_21321,N_21211);
nand U21538 (N_21538,N_21367,N_21378);
and U21539 (N_21539,N_21340,N_21270);
nand U21540 (N_21540,N_21301,N_21335);
nor U21541 (N_21541,N_21395,N_21378);
nand U21542 (N_21542,N_21343,N_21210);
and U21543 (N_21543,N_21304,N_21352);
or U21544 (N_21544,N_21323,N_21200);
or U21545 (N_21545,N_21212,N_21328);
or U21546 (N_21546,N_21366,N_21271);
and U21547 (N_21547,N_21376,N_21339);
nor U21548 (N_21548,N_21326,N_21314);
or U21549 (N_21549,N_21263,N_21228);
nand U21550 (N_21550,N_21272,N_21293);
or U21551 (N_21551,N_21283,N_21254);
nand U21552 (N_21552,N_21246,N_21342);
nand U21553 (N_21553,N_21204,N_21322);
xnor U21554 (N_21554,N_21273,N_21217);
nand U21555 (N_21555,N_21248,N_21271);
nand U21556 (N_21556,N_21300,N_21225);
and U21557 (N_21557,N_21276,N_21374);
and U21558 (N_21558,N_21316,N_21273);
nand U21559 (N_21559,N_21331,N_21209);
nor U21560 (N_21560,N_21362,N_21325);
and U21561 (N_21561,N_21280,N_21225);
nor U21562 (N_21562,N_21347,N_21317);
or U21563 (N_21563,N_21211,N_21317);
nor U21564 (N_21564,N_21366,N_21233);
nand U21565 (N_21565,N_21377,N_21394);
nor U21566 (N_21566,N_21323,N_21307);
and U21567 (N_21567,N_21386,N_21252);
or U21568 (N_21568,N_21230,N_21286);
and U21569 (N_21569,N_21306,N_21353);
and U21570 (N_21570,N_21387,N_21370);
nand U21571 (N_21571,N_21333,N_21342);
or U21572 (N_21572,N_21332,N_21259);
or U21573 (N_21573,N_21272,N_21260);
or U21574 (N_21574,N_21266,N_21231);
and U21575 (N_21575,N_21289,N_21245);
nand U21576 (N_21576,N_21231,N_21236);
or U21577 (N_21577,N_21277,N_21286);
nor U21578 (N_21578,N_21246,N_21376);
nor U21579 (N_21579,N_21373,N_21226);
nor U21580 (N_21580,N_21391,N_21238);
and U21581 (N_21581,N_21338,N_21342);
or U21582 (N_21582,N_21228,N_21243);
nor U21583 (N_21583,N_21320,N_21218);
nor U21584 (N_21584,N_21389,N_21284);
and U21585 (N_21585,N_21207,N_21268);
nor U21586 (N_21586,N_21271,N_21224);
and U21587 (N_21587,N_21276,N_21345);
nand U21588 (N_21588,N_21227,N_21367);
or U21589 (N_21589,N_21359,N_21248);
nor U21590 (N_21590,N_21351,N_21352);
nand U21591 (N_21591,N_21212,N_21381);
nand U21592 (N_21592,N_21283,N_21340);
nor U21593 (N_21593,N_21297,N_21368);
nand U21594 (N_21594,N_21326,N_21284);
nor U21595 (N_21595,N_21392,N_21292);
or U21596 (N_21596,N_21286,N_21338);
or U21597 (N_21597,N_21291,N_21367);
and U21598 (N_21598,N_21267,N_21362);
or U21599 (N_21599,N_21308,N_21258);
and U21600 (N_21600,N_21568,N_21540);
nor U21601 (N_21601,N_21422,N_21483);
and U21602 (N_21602,N_21508,N_21526);
or U21603 (N_21603,N_21432,N_21567);
or U21604 (N_21604,N_21489,N_21465);
or U21605 (N_21605,N_21573,N_21589);
nand U21606 (N_21606,N_21518,N_21463);
nor U21607 (N_21607,N_21495,N_21597);
or U21608 (N_21608,N_21452,N_21494);
or U21609 (N_21609,N_21481,N_21453);
or U21610 (N_21610,N_21598,N_21493);
nand U21611 (N_21611,N_21516,N_21504);
or U21612 (N_21612,N_21549,N_21466);
nand U21613 (N_21613,N_21513,N_21414);
nor U21614 (N_21614,N_21557,N_21442);
nor U21615 (N_21615,N_21469,N_21460);
and U21616 (N_21616,N_21500,N_21529);
nor U21617 (N_21617,N_21541,N_21417);
nand U21618 (N_21618,N_21401,N_21487);
or U21619 (N_21619,N_21461,N_21402);
nor U21620 (N_21620,N_21475,N_21509);
nand U21621 (N_21621,N_21534,N_21559);
or U21622 (N_21622,N_21588,N_21521);
nor U21623 (N_21623,N_21490,N_21431);
nand U21624 (N_21624,N_21595,N_21464);
xnor U21625 (N_21625,N_21480,N_21554);
or U21626 (N_21626,N_21507,N_21524);
and U21627 (N_21627,N_21551,N_21581);
and U21628 (N_21628,N_21436,N_21553);
nand U21629 (N_21629,N_21499,N_21425);
nor U21630 (N_21630,N_21497,N_21435);
or U21631 (N_21631,N_21515,N_21514);
or U21632 (N_21632,N_21531,N_21512);
nor U21633 (N_21633,N_21583,N_21582);
nand U21634 (N_21634,N_21471,N_21522);
nand U21635 (N_21635,N_21438,N_21478);
nand U21636 (N_21636,N_21506,N_21415);
xnor U21637 (N_21637,N_21510,N_21537);
nand U21638 (N_21638,N_21468,N_21416);
nor U21639 (N_21639,N_21586,N_21538);
nor U21640 (N_21640,N_21574,N_21420);
and U21641 (N_21641,N_21457,N_21410);
or U21642 (N_21642,N_21548,N_21407);
or U21643 (N_21643,N_21484,N_21532);
xnor U21644 (N_21644,N_21547,N_21450);
nand U21645 (N_21645,N_21569,N_21498);
and U21646 (N_21646,N_21587,N_21520);
or U21647 (N_21647,N_21545,N_21562);
and U21648 (N_21648,N_21561,N_21578);
and U21649 (N_21649,N_21428,N_21426);
nand U21650 (N_21650,N_21555,N_21570);
nor U21651 (N_21651,N_21488,N_21444);
nand U21652 (N_21652,N_21527,N_21405);
nand U21653 (N_21653,N_21473,N_21590);
or U21654 (N_21654,N_21519,N_21523);
nand U21655 (N_21655,N_21451,N_21421);
nand U21656 (N_21656,N_21593,N_21544);
nand U21657 (N_21657,N_21543,N_21528);
nand U21658 (N_21658,N_21418,N_21400);
nor U21659 (N_21659,N_21479,N_21413);
or U21660 (N_21660,N_21448,N_21445);
or U21661 (N_21661,N_21446,N_21434);
nand U21662 (N_21662,N_21533,N_21579);
nor U21663 (N_21663,N_21505,N_21572);
and U21664 (N_21664,N_21501,N_21535);
nor U21665 (N_21665,N_21552,N_21409);
nand U21666 (N_21666,N_21580,N_21467);
nand U21667 (N_21667,N_21486,N_21536);
nor U21668 (N_21668,N_21454,N_21511);
xor U21669 (N_21669,N_21575,N_21403);
and U21670 (N_21670,N_21591,N_21455);
or U21671 (N_21671,N_21556,N_21530);
xnor U21672 (N_21672,N_21462,N_21577);
or U21673 (N_21673,N_21408,N_21423);
and U21674 (N_21674,N_21419,N_21566);
nand U21675 (N_21675,N_21592,N_21485);
nor U21676 (N_21676,N_21599,N_21492);
nor U21677 (N_21677,N_21449,N_21576);
nand U21678 (N_21678,N_21433,N_21558);
nand U21679 (N_21679,N_21571,N_21458);
nand U21680 (N_21680,N_21565,N_21470);
nand U21681 (N_21681,N_21482,N_21447);
or U21682 (N_21682,N_21546,N_21472);
and U21683 (N_21683,N_21542,N_21503);
and U21684 (N_21684,N_21459,N_21476);
and U21685 (N_21685,N_21594,N_21517);
or U21686 (N_21686,N_21424,N_21525);
and U21687 (N_21687,N_21443,N_21560);
nand U21688 (N_21688,N_21584,N_21539);
nor U21689 (N_21689,N_21596,N_21429);
xnor U21690 (N_21690,N_21491,N_21585);
or U21691 (N_21691,N_21412,N_21474);
nor U21692 (N_21692,N_21496,N_21441);
nand U21693 (N_21693,N_21427,N_21502);
or U21694 (N_21694,N_21550,N_21430);
nand U21695 (N_21695,N_21563,N_21440);
nor U21696 (N_21696,N_21404,N_21456);
and U21697 (N_21697,N_21477,N_21564);
nor U21698 (N_21698,N_21406,N_21437);
and U21699 (N_21699,N_21439,N_21411);
or U21700 (N_21700,N_21591,N_21510);
nand U21701 (N_21701,N_21449,N_21466);
nand U21702 (N_21702,N_21471,N_21577);
and U21703 (N_21703,N_21592,N_21479);
nand U21704 (N_21704,N_21572,N_21514);
nor U21705 (N_21705,N_21459,N_21533);
and U21706 (N_21706,N_21534,N_21408);
and U21707 (N_21707,N_21585,N_21475);
nand U21708 (N_21708,N_21474,N_21518);
or U21709 (N_21709,N_21417,N_21454);
xor U21710 (N_21710,N_21551,N_21594);
and U21711 (N_21711,N_21401,N_21461);
xor U21712 (N_21712,N_21553,N_21497);
nand U21713 (N_21713,N_21560,N_21415);
and U21714 (N_21714,N_21464,N_21583);
nor U21715 (N_21715,N_21458,N_21474);
nand U21716 (N_21716,N_21580,N_21560);
nor U21717 (N_21717,N_21512,N_21414);
and U21718 (N_21718,N_21568,N_21460);
and U21719 (N_21719,N_21403,N_21441);
nor U21720 (N_21720,N_21543,N_21545);
and U21721 (N_21721,N_21446,N_21423);
nand U21722 (N_21722,N_21516,N_21570);
nor U21723 (N_21723,N_21449,N_21480);
nor U21724 (N_21724,N_21509,N_21555);
or U21725 (N_21725,N_21577,N_21431);
and U21726 (N_21726,N_21596,N_21497);
nor U21727 (N_21727,N_21516,N_21532);
or U21728 (N_21728,N_21594,N_21400);
and U21729 (N_21729,N_21443,N_21433);
and U21730 (N_21730,N_21505,N_21519);
nand U21731 (N_21731,N_21530,N_21492);
nand U21732 (N_21732,N_21484,N_21453);
or U21733 (N_21733,N_21407,N_21591);
xor U21734 (N_21734,N_21567,N_21598);
and U21735 (N_21735,N_21444,N_21555);
nor U21736 (N_21736,N_21451,N_21580);
and U21737 (N_21737,N_21550,N_21455);
nand U21738 (N_21738,N_21458,N_21545);
or U21739 (N_21739,N_21517,N_21543);
and U21740 (N_21740,N_21426,N_21579);
and U21741 (N_21741,N_21492,N_21462);
and U21742 (N_21742,N_21501,N_21507);
nand U21743 (N_21743,N_21482,N_21502);
or U21744 (N_21744,N_21442,N_21461);
or U21745 (N_21745,N_21509,N_21461);
nor U21746 (N_21746,N_21570,N_21524);
and U21747 (N_21747,N_21425,N_21540);
nor U21748 (N_21748,N_21402,N_21530);
nand U21749 (N_21749,N_21425,N_21525);
or U21750 (N_21750,N_21536,N_21591);
and U21751 (N_21751,N_21563,N_21445);
or U21752 (N_21752,N_21406,N_21441);
and U21753 (N_21753,N_21485,N_21400);
nand U21754 (N_21754,N_21580,N_21445);
nand U21755 (N_21755,N_21473,N_21461);
xnor U21756 (N_21756,N_21430,N_21437);
nor U21757 (N_21757,N_21515,N_21588);
and U21758 (N_21758,N_21400,N_21450);
and U21759 (N_21759,N_21514,N_21432);
or U21760 (N_21760,N_21484,N_21425);
nor U21761 (N_21761,N_21415,N_21465);
nor U21762 (N_21762,N_21489,N_21575);
and U21763 (N_21763,N_21413,N_21507);
nand U21764 (N_21764,N_21403,N_21456);
nand U21765 (N_21765,N_21416,N_21555);
xnor U21766 (N_21766,N_21482,N_21457);
nand U21767 (N_21767,N_21412,N_21516);
xnor U21768 (N_21768,N_21594,N_21534);
and U21769 (N_21769,N_21463,N_21504);
or U21770 (N_21770,N_21551,N_21536);
nand U21771 (N_21771,N_21427,N_21586);
or U21772 (N_21772,N_21440,N_21473);
nand U21773 (N_21773,N_21543,N_21403);
nand U21774 (N_21774,N_21421,N_21490);
nand U21775 (N_21775,N_21558,N_21410);
or U21776 (N_21776,N_21599,N_21486);
nand U21777 (N_21777,N_21513,N_21527);
nor U21778 (N_21778,N_21520,N_21566);
or U21779 (N_21779,N_21414,N_21576);
or U21780 (N_21780,N_21553,N_21519);
nand U21781 (N_21781,N_21551,N_21532);
nor U21782 (N_21782,N_21571,N_21594);
or U21783 (N_21783,N_21414,N_21440);
nand U21784 (N_21784,N_21547,N_21445);
xor U21785 (N_21785,N_21414,N_21567);
or U21786 (N_21786,N_21528,N_21568);
nand U21787 (N_21787,N_21494,N_21553);
or U21788 (N_21788,N_21580,N_21438);
nand U21789 (N_21789,N_21428,N_21422);
nor U21790 (N_21790,N_21450,N_21535);
and U21791 (N_21791,N_21427,N_21461);
nor U21792 (N_21792,N_21538,N_21587);
and U21793 (N_21793,N_21445,N_21451);
nand U21794 (N_21794,N_21529,N_21598);
xnor U21795 (N_21795,N_21550,N_21453);
nand U21796 (N_21796,N_21474,N_21551);
nor U21797 (N_21797,N_21468,N_21438);
and U21798 (N_21798,N_21461,N_21464);
nand U21799 (N_21799,N_21552,N_21469);
nor U21800 (N_21800,N_21677,N_21674);
nand U21801 (N_21801,N_21765,N_21726);
or U21802 (N_21802,N_21712,N_21609);
nor U21803 (N_21803,N_21752,N_21699);
nor U21804 (N_21804,N_21620,N_21692);
nor U21805 (N_21805,N_21644,N_21707);
and U21806 (N_21806,N_21708,N_21642);
nor U21807 (N_21807,N_21612,N_21600);
nor U21808 (N_21808,N_21788,N_21728);
and U21809 (N_21809,N_21755,N_21686);
and U21810 (N_21810,N_21790,N_21774);
or U21811 (N_21811,N_21624,N_21610);
nand U21812 (N_21812,N_21616,N_21649);
xnor U21813 (N_21813,N_21710,N_21757);
xor U21814 (N_21814,N_21756,N_21682);
and U21815 (N_21815,N_21743,N_21727);
or U21816 (N_21816,N_21732,N_21725);
nand U21817 (N_21817,N_21664,N_21691);
and U21818 (N_21818,N_21604,N_21643);
nand U21819 (N_21819,N_21781,N_21722);
nand U21820 (N_21820,N_21621,N_21602);
and U21821 (N_21821,N_21775,N_21650);
nor U21822 (N_21822,N_21676,N_21611);
nor U21823 (N_21823,N_21723,N_21639);
and U21824 (N_21824,N_21760,N_21690);
or U21825 (N_21825,N_21766,N_21715);
nor U21826 (N_21826,N_21720,N_21635);
or U21827 (N_21827,N_21764,N_21736);
or U21828 (N_21828,N_21769,N_21648);
or U21829 (N_21829,N_21672,N_21670);
and U21830 (N_21830,N_21794,N_21799);
or U21831 (N_21831,N_21660,N_21749);
nand U21832 (N_21832,N_21713,N_21633);
nor U21833 (N_21833,N_21661,N_21787);
or U21834 (N_21834,N_21714,N_21745);
or U21835 (N_21835,N_21748,N_21773);
or U21836 (N_21836,N_21750,N_21735);
or U21837 (N_21837,N_21758,N_21739);
nand U21838 (N_21838,N_21771,N_21717);
nor U21839 (N_21839,N_21785,N_21729);
or U21840 (N_21840,N_21606,N_21646);
xnor U21841 (N_21841,N_21683,N_21669);
and U21842 (N_21842,N_21614,N_21663);
nand U21843 (N_21843,N_21605,N_21716);
nand U21844 (N_21844,N_21637,N_21731);
xor U21845 (N_21845,N_21623,N_21629);
xor U21846 (N_21846,N_21608,N_21619);
nand U21847 (N_21847,N_21741,N_21615);
nand U21848 (N_21848,N_21656,N_21657);
nor U21849 (N_21849,N_21627,N_21640);
or U21850 (N_21850,N_21667,N_21742);
nand U21851 (N_21851,N_21747,N_21770);
xnor U21852 (N_21852,N_21701,N_21703);
nor U21853 (N_21853,N_21733,N_21671);
nor U21854 (N_21854,N_21645,N_21798);
or U21855 (N_21855,N_21777,N_21696);
nand U21856 (N_21856,N_21655,N_21719);
nor U21857 (N_21857,N_21704,N_21636);
and U21858 (N_21858,N_21630,N_21622);
and U21859 (N_21859,N_21776,N_21680);
xnor U21860 (N_21860,N_21617,N_21734);
or U21861 (N_21861,N_21698,N_21638);
xor U21862 (N_21862,N_21767,N_21652);
and U21863 (N_21863,N_21753,N_21763);
nand U21864 (N_21864,N_21628,N_21618);
or U21865 (N_21865,N_21675,N_21689);
or U21866 (N_21866,N_21778,N_21706);
and U21867 (N_21867,N_21631,N_21738);
and U21868 (N_21868,N_21795,N_21694);
nand U21869 (N_21869,N_21705,N_21641);
nor U21870 (N_21870,N_21786,N_21784);
xnor U21871 (N_21871,N_21768,N_21603);
xor U21872 (N_21872,N_21737,N_21601);
or U21873 (N_21873,N_21721,N_21679);
xnor U21874 (N_21874,N_21700,N_21744);
nand U21875 (N_21875,N_21796,N_21792);
and U21876 (N_21876,N_21746,N_21779);
nand U21877 (N_21877,N_21695,N_21780);
nor U21878 (N_21878,N_21626,N_21709);
or U21879 (N_21879,N_21632,N_21791);
nor U21880 (N_21880,N_21697,N_21678);
or U21881 (N_21881,N_21668,N_21625);
and U21882 (N_21882,N_21711,N_21688);
and U21883 (N_21883,N_21673,N_21797);
or U21884 (N_21884,N_21613,N_21702);
nand U21885 (N_21885,N_21685,N_21665);
nor U21886 (N_21886,N_21693,N_21782);
and U21887 (N_21887,N_21761,N_21740);
xor U21888 (N_21888,N_21651,N_21659);
or U21889 (N_21889,N_21653,N_21793);
nand U21890 (N_21890,N_21718,N_21634);
and U21891 (N_21891,N_21783,N_21730);
nor U21892 (N_21892,N_21724,N_21789);
or U21893 (N_21893,N_21647,N_21666);
and U21894 (N_21894,N_21772,N_21662);
nor U21895 (N_21895,N_21759,N_21681);
nand U21896 (N_21896,N_21687,N_21762);
nand U21897 (N_21897,N_21607,N_21658);
or U21898 (N_21898,N_21654,N_21754);
or U21899 (N_21899,N_21684,N_21751);
and U21900 (N_21900,N_21681,N_21772);
and U21901 (N_21901,N_21687,N_21780);
or U21902 (N_21902,N_21640,N_21655);
or U21903 (N_21903,N_21759,N_21713);
nor U21904 (N_21904,N_21677,N_21711);
nor U21905 (N_21905,N_21773,N_21696);
nand U21906 (N_21906,N_21799,N_21765);
nand U21907 (N_21907,N_21652,N_21690);
and U21908 (N_21908,N_21609,N_21768);
nand U21909 (N_21909,N_21756,N_21760);
or U21910 (N_21910,N_21727,N_21720);
xnor U21911 (N_21911,N_21774,N_21747);
or U21912 (N_21912,N_21642,N_21755);
nor U21913 (N_21913,N_21660,N_21676);
and U21914 (N_21914,N_21612,N_21764);
xnor U21915 (N_21915,N_21628,N_21785);
or U21916 (N_21916,N_21709,N_21785);
xor U21917 (N_21917,N_21728,N_21754);
xor U21918 (N_21918,N_21626,N_21685);
or U21919 (N_21919,N_21777,N_21751);
or U21920 (N_21920,N_21650,N_21621);
and U21921 (N_21921,N_21629,N_21674);
nand U21922 (N_21922,N_21607,N_21688);
xnor U21923 (N_21923,N_21775,N_21613);
nand U21924 (N_21924,N_21780,N_21773);
and U21925 (N_21925,N_21710,N_21675);
nor U21926 (N_21926,N_21605,N_21708);
nor U21927 (N_21927,N_21643,N_21788);
nand U21928 (N_21928,N_21604,N_21669);
or U21929 (N_21929,N_21685,N_21624);
and U21930 (N_21930,N_21612,N_21601);
and U21931 (N_21931,N_21647,N_21796);
and U21932 (N_21932,N_21673,N_21623);
nor U21933 (N_21933,N_21796,N_21687);
and U21934 (N_21934,N_21611,N_21712);
or U21935 (N_21935,N_21797,N_21619);
and U21936 (N_21936,N_21774,N_21609);
nor U21937 (N_21937,N_21603,N_21711);
nor U21938 (N_21938,N_21604,N_21701);
nand U21939 (N_21939,N_21666,N_21731);
xnor U21940 (N_21940,N_21713,N_21741);
nor U21941 (N_21941,N_21740,N_21714);
and U21942 (N_21942,N_21773,N_21635);
nor U21943 (N_21943,N_21676,N_21627);
nand U21944 (N_21944,N_21748,N_21694);
and U21945 (N_21945,N_21771,N_21612);
and U21946 (N_21946,N_21606,N_21758);
nor U21947 (N_21947,N_21746,N_21688);
nor U21948 (N_21948,N_21741,N_21674);
and U21949 (N_21949,N_21790,N_21725);
nor U21950 (N_21950,N_21721,N_21658);
and U21951 (N_21951,N_21731,N_21674);
and U21952 (N_21952,N_21730,N_21646);
xor U21953 (N_21953,N_21752,N_21697);
and U21954 (N_21954,N_21619,N_21600);
or U21955 (N_21955,N_21684,N_21779);
nand U21956 (N_21956,N_21652,N_21758);
nor U21957 (N_21957,N_21670,N_21647);
nor U21958 (N_21958,N_21796,N_21754);
xnor U21959 (N_21959,N_21729,N_21734);
and U21960 (N_21960,N_21680,N_21683);
nand U21961 (N_21961,N_21634,N_21794);
or U21962 (N_21962,N_21702,N_21733);
or U21963 (N_21963,N_21762,N_21713);
and U21964 (N_21964,N_21739,N_21612);
or U21965 (N_21965,N_21634,N_21643);
or U21966 (N_21966,N_21737,N_21715);
nor U21967 (N_21967,N_21672,N_21778);
nor U21968 (N_21968,N_21640,N_21799);
nor U21969 (N_21969,N_21631,N_21774);
and U21970 (N_21970,N_21668,N_21772);
nand U21971 (N_21971,N_21673,N_21735);
or U21972 (N_21972,N_21793,N_21608);
xnor U21973 (N_21973,N_21675,N_21663);
nor U21974 (N_21974,N_21626,N_21641);
nor U21975 (N_21975,N_21739,N_21766);
or U21976 (N_21976,N_21659,N_21602);
nand U21977 (N_21977,N_21741,N_21605);
or U21978 (N_21978,N_21693,N_21743);
xor U21979 (N_21979,N_21657,N_21714);
nor U21980 (N_21980,N_21615,N_21711);
and U21981 (N_21981,N_21606,N_21792);
nor U21982 (N_21982,N_21667,N_21748);
or U21983 (N_21983,N_21751,N_21631);
nor U21984 (N_21984,N_21644,N_21700);
or U21985 (N_21985,N_21654,N_21750);
or U21986 (N_21986,N_21746,N_21708);
or U21987 (N_21987,N_21754,N_21687);
nand U21988 (N_21988,N_21659,N_21600);
and U21989 (N_21989,N_21741,N_21705);
nand U21990 (N_21990,N_21678,N_21782);
or U21991 (N_21991,N_21763,N_21769);
nor U21992 (N_21992,N_21734,N_21615);
and U21993 (N_21993,N_21643,N_21731);
nor U21994 (N_21994,N_21647,N_21668);
nor U21995 (N_21995,N_21686,N_21641);
xnor U21996 (N_21996,N_21734,N_21784);
nand U21997 (N_21997,N_21641,N_21770);
or U21998 (N_21998,N_21763,N_21793);
nor U21999 (N_21999,N_21798,N_21799);
and U22000 (N_22000,N_21817,N_21891);
nor U22001 (N_22001,N_21845,N_21888);
xnor U22002 (N_22002,N_21965,N_21851);
and U22003 (N_22003,N_21880,N_21983);
nor U22004 (N_22004,N_21940,N_21867);
nand U22005 (N_22005,N_21958,N_21863);
or U22006 (N_22006,N_21873,N_21875);
nand U22007 (N_22007,N_21827,N_21991);
xor U22008 (N_22008,N_21869,N_21828);
or U22009 (N_22009,N_21897,N_21979);
nor U22010 (N_22010,N_21802,N_21947);
or U22011 (N_22011,N_21930,N_21945);
nand U22012 (N_22012,N_21987,N_21859);
or U22013 (N_22013,N_21901,N_21878);
nand U22014 (N_22014,N_21813,N_21829);
and U22015 (N_22015,N_21824,N_21865);
nand U22016 (N_22016,N_21938,N_21884);
and U22017 (N_22017,N_21975,N_21808);
or U22018 (N_22018,N_21962,N_21924);
nand U22019 (N_22019,N_21830,N_21870);
nor U22020 (N_22020,N_21803,N_21956);
and U22021 (N_22021,N_21852,N_21821);
xor U22022 (N_22022,N_21915,N_21892);
nand U22023 (N_22023,N_21853,N_21810);
nor U22024 (N_22024,N_21960,N_21942);
and U22025 (N_22025,N_21970,N_21804);
nor U22026 (N_22026,N_21847,N_21874);
or U22027 (N_22027,N_21887,N_21883);
nor U22028 (N_22028,N_21978,N_21946);
or U22029 (N_22029,N_21860,N_21834);
and U22030 (N_22030,N_21997,N_21848);
or U22031 (N_22031,N_21876,N_21909);
and U22032 (N_22032,N_21833,N_21996);
xor U22033 (N_22033,N_21855,N_21879);
and U22034 (N_22034,N_21966,N_21949);
and U22035 (N_22035,N_21919,N_21937);
nand U22036 (N_22036,N_21925,N_21910);
nand U22037 (N_22037,N_21964,N_21886);
nand U22038 (N_22038,N_21927,N_21928);
or U22039 (N_22039,N_21895,N_21844);
or U22040 (N_22040,N_21904,N_21843);
and U22041 (N_22041,N_21974,N_21872);
or U22042 (N_22042,N_21973,N_21850);
xnor U22043 (N_22043,N_21939,N_21906);
nor U22044 (N_22044,N_21814,N_21818);
nand U22045 (N_22045,N_21862,N_21842);
nor U22046 (N_22046,N_21838,N_21999);
and U22047 (N_22047,N_21941,N_21809);
and U22048 (N_22048,N_21963,N_21986);
or U22049 (N_22049,N_21846,N_21861);
nand U22050 (N_22050,N_21837,N_21898);
xnor U22051 (N_22051,N_21820,N_21957);
and U22052 (N_22052,N_21835,N_21980);
nand U22053 (N_22053,N_21936,N_21926);
nand U22054 (N_22054,N_21993,N_21900);
nand U22055 (N_22055,N_21836,N_21972);
and U22056 (N_22056,N_21841,N_21893);
nor U22057 (N_22057,N_21806,N_21932);
nand U22058 (N_22058,N_21988,N_21995);
nor U22059 (N_22059,N_21931,N_21922);
nor U22060 (N_22060,N_21882,N_21961);
nand U22061 (N_22061,N_21934,N_21994);
and U22062 (N_22062,N_21856,N_21984);
and U22063 (N_22063,N_21826,N_21959);
and U22064 (N_22064,N_21952,N_21969);
nor U22065 (N_22065,N_21933,N_21816);
or U22066 (N_22066,N_21890,N_21825);
xnor U22067 (N_22067,N_21977,N_21968);
or U22068 (N_22068,N_21839,N_21811);
and U22069 (N_22069,N_21823,N_21967);
nor U22070 (N_22070,N_21920,N_21881);
and U22071 (N_22071,N_21868,N_21871);
nand U22072 (N_22072,N_21894,N_21899);
or U22073 (N_22073,N_21857,N_21921);
nand U22074 (N_22074,N_21992,N_21864);
and U22075 (N_22075,N_21923,N_21812);
xnor U22076 (N_22076,N_21889,N_21918);
nor U22077 (N_22077,N_21914,N_21807);
and U22078 (N_22078,N_21998,N_21976);
nor U22079 (N_22079,N_21908,N_21911);
or U22080 (N_22080,N_21805,N_21943);
and U22081 (N_22081,N_21953,N_21955);
nor U22082 (N_22082,N_21819,N_21929);
or U22083 (N_22083,N_21831,N_21854);
and U22084 (N_22084,N_21885,N_21913);
or U22085 (N_22085,N_21877,N_21982);
xnor U22086 (N_22086,N_21935,N_21902);
nand U22087 (N_22087,N_21971,N_21985);
and U22088 (N_22088,N_21917,N_21832);
and U22089 (N_22089,N_21858,N_21903);
or U22090 (N_22090,N_21907,N_21950);
or U22091 (N_22091,N_21800,N_21912);
nor U22092 (N_22092,N_21801,N_21822);
or U22093 (N_22093,N_21948,N_21896);
and U22094 (N_22094,N_21866,N_21990);
or U22095 (N_22095,N_21916,N_21849);
or U22096 (N_22096,N_21944,N_21989);
or U22097 (N_22097,N_21951,N_21954);
xor U22098 (N_22098,N_21840,N_21815);
or U22099 (N_22099,N_21981,N_21905);
nor U22100 (N_22100,N_21951,N_21989);
nand U22101 (N_22101,N_21988,N_21906);
nor U22102 (N_22102,N_21824,N_21942);
or U22103 (N_22103,N_21823,N_21934);
nor U22104 (N_22104,N_21945,N_21873);
nand U22105 (N_22105,N_21966,N_21853);
nand U22106 (N_22106,N_21960,N_21804);
and U22107 (N_22107,N_21966,N_21854);
xor U22108 (N_22108,N_21921,N_21979);
or U22109 (N_22109,N_21882,N_21884);
nand U22110 (N_22110,N_21957,N_21890);
xnor U22111 (N_22111,N_21952,N_21943);
and U22112 (N_22112,N_21994,N_21959);
nand U22113 (N_22113,N_21936,N_21990);
or U22114 (N_22114,N_21931,N_21932);
nand U22115 (N_22115,N_21808,N_21933);
nor U22116 (N_22116,N_21930,N_21925);
or U22117 (N_22117,N_21969,N_21975);
and U22118 (N_22118,N_21990,N_21916);
and U22119 (N_22119,N_21826,N_21811);
nor U22120 (N_22120,N_21818,N_21918);
and U22121 (N_22121,N_21893,N_21926);
and U22122 (N_22122,N_21958,N_21941);
nor U22123 (N_22123,N_21934,N_21856);
nand U22124 (N_22124,N_21901,N_21833);
nand U22125 (N_22125,N_21962,N_21943);
nor U22126 (N_22126,N_21978,N_21994);
nor U22127 (N_22127,N_21866,N_21917);
nor U22128 (N_22128,N_21819,N_21848);
or U22129 (N_22129,N_21809,N_21951);
or U22130 (N_22130,N_21995,N_21878);
nand U22131 (N_22131,N_21803,N_21870);
nand U22132 (N_22132,N_21831,N_21855);
and U22133 (N_22133,N_21880,N_21804);
nor U22134 (N_22134,N_21910,N_21854);
and U22135 (N_22135,N_21875,N_21825);
xnor U22136 (N_22136,N_21801,N_21839);
nor U22137 (N_22137,N_21849,N_21956);
and U22138 (N_22138,N_21855,N_21966);
nand U22139 (N_22139,N_21931,N_21824);
nor U22140 (N_22140,N_21888,N_21990);
nand U22141 (N_22141,N_21979,N_21988);
nor U22142 (N_22142,N_21924,N_21823);
and U22143 (N_22143,N_21899,N_21812);
or U22144 (N_22144,N_21840,N_21828);
or U22145 (N_22145,N_21857,N_21814);
and U22146 (N_22146,N_21804,N_21852);
and U22147 (N_22147,N_21923,N_21988);
or U22148 (N_22148,N_21866,N_21801);
nand U22149 (N_22149,N_21966,N_21938);
nand U22150 (N_22150,N_21809,N_21859);
nor U22151 (N_22151,N_21929,N_21907);
nand U22152 (N_22152,N_21886,N_21838);
or U22153 (N_22153,N_21914,N_21983);
nand U22154 (N_22154,N_21817,N_21933);
nor U22155 (N_22155,N_21962,N_21904);
or U22156 (N_22156,N_21946,N_21871);
or U22157 (N_22157,N_21954,N_21860);
nor U22158 (N_22158,N_21991,N_21865);
nor U22159 (N_22159,N_21908,N_21959);
or U22160 (N_22160,N_21925,N_21929);
nand U22161 (N_22161,N_21924,N_21889);
nand U22162 (N_22162,N_21984,N_21830);
and U22163 (N_22163,N_21854,N_21924);
nor U22164 (N_22164,N_21800,N_21867);
and U22165 (N_22165,N_21920,N_21912);
and U22166 (N_22166,N_21933,N_21944);
or U22167 (N_22167,N_21934,N_21839);
or U22168 (N_22168,N_21857,N_21967);
nor U22169 (N_22169,N_21830,N_21929);
or U22170 (N_22170,N_21884,N_21896);
or U22171 (N_22171,N_21805,N_21832);
nor U22172 (N_22172,N_21993,N_21882);
nor U22173 (N_22173,N_21929,N_21845);
nand U22174 (N_22174,N_21827,N_21823);
and U22175 (N_22175,N_21951,N_21802);
and U22176 (N_22176,N_21863,N_21807);
nor U22177 (N_22177,N_21924,N_21951);
xor U22178 (N_22178,N_21919,N_21830);
or U22179 (N_22179,N_21926,N_21915);
nor U22180 (N_22180,N_21928,N_21891);
and U22181 (N_22181,N_21889,N_21922);
nor U22182 (N_22182,N_21949,N_21951);
and U22183 (N_22183,N_21804,N_21848);
and U22184 (N_22184,N_21928,N_21945);
nand U22185 (N_22185,N_21802,N_21940);
and U22186 (N_22186,N_21983,N_21960);
and U22187 (N_22187,N_21976,N_21996);
or U22188 (N_22188,N_21862,N_21846);
or U22189 (N_22189,N_21813,N_21891);
nor U22190 (N_22190,N_21918,N_21869);
xor U22191 (N_22191,N_21838,N_21969);
or U22192 (N_22192,N_21829,N_21973);
and U22193 (N_22193,N_21854,N_21946);
nand U22194 (N_22194,N_21914,N_21933);
nor U22195 (N_22195,N_21920,N_21990);
nand U22196 (N_22196,N_21835,N_21952);
nor U22197 (N_22197,N_21813,N_21921);
xnor U22198 (N_22198,N_21949,N_21959);
nand U22199 (N_22199,N_21810,N_21895);
xor U22200 (N_22200,N_22128,N_22019);
nand U22201 (N_22201,N_22078,N_22015);
nor U22202 (N_22202,N_22046,N_22088);
nand U22203 (N_22203,N_22156,N_22186);
or U22204 (N_22204,N_22005,N_22179);
nor U22205 (N_22205,N_22153,N_22080);
and U22206 (N_22206,N_22126,N_22065);
nor U22207 (N_22207,N_22119,N_22079);
nand U22208 (N_22208,N_22137,N_22073);
or U22209 (N_22209,N_22150,N_22011);
and U22210 (N_22210,N_22169,N_22028);
and U22211 (N_22211,N_22081,N_22101);
or U22212 (N_22212,N_22180,N_22068);
or U22213 (N_22213,N_22050,N_22157);
and U22214 (N_22214,N_22199,N_22087);
and U22215 (N_22215,N_22004,N_22163);
xnor U22216 (N_22216,N_22021,N_22172);
nor U22217 (N_22217,N_22164,N_22109);
nor U22218 (N_22218,N_22012,N_22111);
and U22219 (N_22219,N_22095,N_22192);
or U22220 (N_22220,N_22056,N_22125);
nand U22221 (N_22221,N_22132,N_22002);
or U22222 (N_22222,N_22149,N_22194);
and U22223 (N_22223,N_22069,N_22123);
or U22224 (N_22224,N_22084,N_22178);
nand U22225 (N_22225,N_22110,N_22060);
or U22226 (N_22226,N_22189,N_22176);
nand U22227 (N_22227,N_22035,N_22092);
xnor U22228 (N_22228,N_22130,N_22097);
and U22229 (N_22229,N_22170,N_22196);
or U22230 (N_22230,N_22049,N_22001);
and U22231 (N_22231,N_22122,N_22010);
nand U22232 (N_22232,N_22051,N_22098);
nor U22233 (N_22233,N_22053,N_22096);
and U22234 (N_22234,N_22070,N_22127);
and U22235 (N_22235,N_22031,N_22131);
and U22236 (N_22236,N_22147,N_22198);
and U22237 (N_22237,N_22102,N_22168);
xor U22238 (N_22238,N_22134,N_22182);
and U22239 (N_22239,N_22171,N_22190);
or U22240 (N_22240,N_22066,N_22183);
nand U22241 (N_22241,N_22055,N_22036);
and U22242 (N_22242,N_22181,N_22144);
and U22243 (N_22243,N_22043,N_22191);
nor U22244 (N_22244,N_22121,N_22072);
nor U22245 (N_22245,N_22136,N_22006);
nand U22246 (N_22246,N_22003,N_22082);
nor U22247 (N_22247,N_22117,N_22175);
nand U22248 (N_22248,N_22029,N_22041);
nand U22249 (N_22249,N_22146,N_22140);
or U22250 (N_22250,N_22113,N_22047);
nor U22251 (N_22251,N_22090,N_22103);
nor U22252 (N_22252,N_22104,N_22009);
or U22253 (N_22253,N_22173,N_22148);
nand U22254 (N_22254,N_22177,N_22052);
or U22255 (N_22255,N_22094,N_22106);
and U22256 (N_22256,N_22145,N_22187);
or U22257 (N_22257,N_22120,N_22040);
nand U22258 (N_22258,N_22034,N_22016);
nand U22259 (N_22259,N_22032,N_22185);
and U22260 (N_22260,N_22100,N_22155);
and U22261 (N_22261,N_22159,N_22118);
and U22262 (N_22262,N_22024,N_22057);
and U22263 (N_22263,N_22048,N_22165);
nor U22264 (N_22264,N_22115,N_22152);
nand U22265 (N_22265,N_22017,N_22184);
or U22266 (N_22266,N_22174,N_22074);
nand U22267 (N_22267,N_22161,N_22030);
or U22268 (N_22268,N_22162,N_22129);
and U22269 (N_22269,N_22023,N_22022);
and U22270 (N_22270,N_22105,N_22124);
xnor U22271 (N_22271,N_22142,N_22154);
xor U22272 (N_22272,N_22099,N_22013);
and U22273 (N_22273,N_22085,N_22167);
and U22274 (N_22274,N_22045,N_22062);
nand U22275 (N_22275,N_22000,N_22018);
and U22276 (N_22276,N_22026,N_22114);
and U22277 (N_22277,N_22058,N_22139);
nor U22278 (N_22278,N_22197,N_22195);
nand U22279 (N_22279,N_22188,N_22025);
nor U22280 (N_22280,N_22020,N_22071);
and U22281 (N_22281,N_22014,N_22083);
nand U22282 (N_22282,N_22067,N_22112);
or U22283 (N_22283,N_22160,N_22138);
nor U22284 (N_22284,N_22151,N_22061);
and U22285 (N_22285,N_22027,N_22108);
xor U22286 (N_22286,N_22044,N_22059);
and U22287 (N_22287,N_22033,N_22039);
or U22288 (N_22288,N_22037,N_22193);
xor U22289 (N_22289,N_22076,N_22077);
nor U22290 (N_22290,N_22008,N_22086);
nor U22291 (N_22291,N_22141,N_22007);
xnor U22292 (N_22292,N_22063,N_22042);
nand U22293 (N_22293,N_22107,N_22093);
or U22294 (N_22294,N_22038,N_22158);
nand U22295 (N_22295,N_22116,N_22089);
xnor U22296 (N_22296,N_22091,N_22075);
and U22297 (N_22297,N_22064,N_22135);
or U22298 (N_22298,N_22166,N_22133);
xor U22299 (N_22299,N_22054,N_22143);
xnor U22300 (N_22300,N_22159,N_22069);
nor U22301 (N_22301,N_22166,N_22149);
or U22302 (N_22302,N_22098,N_22157);
or U22303 (N_22303,N_22098,N_22010);
and U22304 (N_22304,N_22107,N_22082);
and U22305 (N_22305,N_22165,N_22034);
or U22306 (N_22306,N_22012,N_22134);
xor U22307 (N_22307,N_22092,N_22020);
or U22308 (N_22308,N_22013,N_22125);
or U22309 (N_22309,N_22035,N_22165);
nand U22310 (N_22310,N_22093,N_22064);
and U22311 (N_22311,N_22051,N_22018);
or U22312 (N_22312,N_22000,N_22150);
nand U22313 (N_22313,N_22197,N_22046);
nor U22314 (N_22314,N_22189,N_22079);
and U22315 (N_22315,N_22087,N_22080);
nand U22316 (N_22316,N_22098,N_22064);
xnor U22317 (N_22317,N_22188,N_22139);
nor U22318 (N_22318,N_22039,N_22083);
xor U22319 (N_22319,N_22132,N_22054);
nand U22320 (N_22320,N_22081,N_22009);
nand U22321 (N_22321,N_22198,N_22104);
nand U22322 (N_22322,N_22064,N_22033);
and U22323 (N_22323,N_22138,N_22170);
and U22324 (N_22324,N_22078,N_22150);
and U22325 (N_22325,N_22028,N_22082);
nand U22326 (N_22326,N_22021,N_22025);
or U22327 (N_22327,N_22073,N_22086);
or U22328 (N_22328,N_22047,N_22087);
and U22329 (N_22329,N_22174,N_22195);
nand U22330 (N_22330,N_22124,N_22151);
nand U22331 (N_22331,N_22153,N_22114);
nand U22332 (N_22332,N_22191,N_22188);
nand U22333 (N_22333,N_22098,N_22111);
xor U22334 (N_22334,N_22093,N_22180);
nor U22335 (N_22335,N_22114,N_22084);
or U22336 (N_22336,N_22182,N_22059);
and U22337 (N_22337,N_22125,N_22112);
or U22338 (N_22338,N_22019,N_22073);
and U22339 (N_22339,N_22023,N_22104);
or U22340 (N_22340,N_22001,N_22056);
nand U22341 (N_22341,N_22040,N_22112);
or U22342 (N_22342,N_22127,N_22145);
nand U22343 (N_22343,N_22121,N_22196);
xor U22344 (N_22344,N_22014,N_22013);
nand U22345 (N_22345,N_22198,N_22000);
and U22346 (N_22346,N_22098,N_22092);
nand U22347 (N_22347,N_22163,N_22090);
nand U22348 (N_22348,N_22152,N_22071);
or U22349 (N_22349,N_22001,N_22071);
and U22350 (N_22350,N_22145,N_22078);
or U22351 (N_22351,N_22103,N_22081);
nand U22352 (N_22352,N_22175,N_22185);
or U22353 (N_22353,N_22178,N_22018);
nor U22354 (N_22354,N_22186,N_22184);
and U22355 (N_22355,N_22195,N_22125);
and U22356 (N_22356,N_22091,N_22171);
and U22357 (N_22357,N_22057,N_22184);
nand U22358 (N_22358,N_22173,N_22055);
nor U22359 (N_22359,N_22093,N_22099);
and U22360 (N_22360,N_22126,N_22085);
or U22361 (N_22361,N_22009,N_22027);
nand U22362 (N_22362,N_22145,N_22132);
or U22363 (N_22363,N_22021,N_22130);
xnor U22364 (N_22364,N_22020,N_22032);
nor U22365 (N_22365,N_22137,N_22128);
nor U22366 (N_22366,N_22156,N_22123);
nand U22367 (N_22367,N_22049,N_22020);
xnor U22368 (N_22368,N_22195,N_22062);
nand U22369 (N_22369,N_22136,N_22150);
nor U22370 (N_22370,N_22009,N_22052);
xor U22371 (N_22371,N_22033,N_22035);
and U22372 (N_22372,N_22151,N_22079);
or U22373 (N_22373,N_22006,N_22153);
and U22374 (N_22374,N_22130,N_22139);
xor U22375 (N_22375,N_22017,N_22174);
nand U22376 (N_22376,N_22058,N_22006);
nor U22377 (N_22377,N_22180,N_22187);
nand U22378 (N_22378,N_22006,N_22079);
and U22379 (N_22379,N_22068,N_22017);
nand U22380 (N_22380,N_22194,N_22109);
nand U22381 (N_22381,N_22041,N_22091);
and U22382 (N_22382,N_22136,N_22124);
and U22383 (N_22383,N_22123,N_22050);
nor U22384 (N_22384,N_22117,N_22082);
xor U22385 (N_22385,N_22026,N_22067);
nor U22386 (N_22386,N_22159,N_22157);
and U22387 (N_22387,N_22003,N_22150);
xor U22388 (N_22388,N_22090,N_22190);
nand U22389 (N_22389,N_22072,N_22053);
or U22390 (N_22390,N_22069,N_22070);
nor U22391 (N_22391,N_22174,N_22057);
nor U22392 (N_22392,N_22132,N_22161);
or U22393 (N_22393,N_22091,N_22162);
xor U22394 (N_22394,N_22084,N_22095);
and U22395 (N_22395,N_22164,N_22036);
or U22396 (N_22396,N_22002,N_22146);
and U22397 (N_22397,N_22054,N_22124);
nand U22398 (N_22398,N_22025,N_22148);
xor U22399 (N_22399,N_22099,N_22081);
and U22400 (N_22400,N_22262,N_22249);
or U22401 (N_22401,N_22264,N_22288);
nor U22402 (N_22402,N_22320,N_22278);
and U22403 (N_22403,N_22398,N_22318);
nand U22404 (N_22404,N_22270,N_22238);
and U22405 (N_22405,N_22258,N_22212);
nor U22406 (N_22406,N_22390,N_22204);
xor U22407 (N_22407,N_22384,N_22216);
or U22408 (N_22408,N_22241,N_22272);
or U22409 (N_22409,N_22225,N_22344);
nand U22410 (N_22410,N_22309,N_22302);
xor U22411 (N_22411,N_22381,N_22339);
or U22412 (N_22412,N_22224,N_22229);
nand U22413 (N_22413,N_22341,N_22222);
nand U22414 (N_22414,N_22243,N_22275);
nand U22415 (N_22415,N_22266,N_22325);
xor U22416 (N_22416,N_22315,N_22327);
xnor U22417 (N_22417,N_22338,N_22373);
xnor U22418 (N_22418,N_22230,N_22392);
and U22419 (N_22419,N_22372,N_22271);
nor U22420 (N_22420,N_22324,N_22274);
or U22421 (N_22421,N_22268,N_22367);
nand U22422 (N_22422,N_22323,N_22334);
nor U22423 (N_22423,N_22218,N_22387);
nor U22424 (N_22424,N_22291,N_22350);
xnor U22425 (N_22425,N_22215,N_22364);
nor U22426 (N_22426,N_22379,N_22386);
nor U22427 (N_22427,N_22371,N_22317);
or U22428 (N_22428,N_22214,N_22296);
xor U22429 (N_22429,N_22231,N_22254);
nand U22430 (N_22430,N_22360,N_22233);
and U22431 (N_22431,N_22248,N_22399);
and U22432 (N_22432,N_22376,N_22365);
and U22433 (N_22433,N_22281,N_22245);
and U22434 (N_22434,N_22242,N_22312);
xnor U22435 (N_22435,N_22255,N_22203);
and U22436 (N_22436,N_22273,N_22206);
nor U22437 (N_22437,N_22213,N_22368);
or U22438 (N_22438,N_22321,N_22232);
nand U22439 (N_22439,N_22363,N_22347);
nand U22440 (N_22440,N_22211,N_22370);
nand U22441 (N_22441,N_22369,N_22263);
nor U22442 (N_22442,N_22202,N_22253);
nor U22443 (N_22443,N_22205,N_22329);
nor U22444 (N_22444,N_22340,N_22345);
or U22445 (N_22445,N_22269,N_22362);
nor U22446 (N_22446,N_22343,N_22303);
nand U22447 (N_22447,N_22280,N_22285);
nor U22448 (N_22448,N_22374,N_22335);
nand U22449 (N_22449,N_22261,N_22375);
xnor U22450 (N_22450,N_22236,N_22353);
and U22451 (N_22451,N_22337,N_22286);
nor U22452 (N_22452,N_22397,N_22385);
nor U22453 (N_22453,N_22277,N_22348);
and U22454 (N_22454,N_22294,N_22319);
nand U22455 (N_22455,N_22391,N_22295);
xnor U22456 (N_22456,N_22265,N_22395);
xor U22457 (N_22457,N_22293,N_22259);
nand U22458 (N_22458,N_22342,N_22276);
nand U22459 (N_22459,N_22396,N_22200);
nand U22460 (N_22460,N_22352,N_22246);
xor U22461 (N_22461,N_22217,N_22207);
nand U22462 (N_22462,N_22223,N_22358);
or U22463 (N_22463,N_22331,N_22287);
or U22464 (N_22464,N_22292,N_22378);
or U22465 (N_22465,N_22284,N_22351);
or U22466 (N_22466,N_22210,N_22235);
and U22467 (N_22467,N_22308,N_22228);
nand U22468 (N_22468,N_22322,N_22393);
or U22469 (N_22469,N_22247,N_22377);
and U22470 (N_22470,N_22221,N_22356);
nor U22471 (N_22471,N_22279,N_22208);
xnor U22472 (N_22472,N_22251,N_22366);
or U22473 (N_22473,N_22306,N_22382);
or U22474 (N_22474,N_22310,N_22305);
xor U22475 (N_22475,N_22332,N_22257);
and U22476 (N_22476,N_22227,N_22244);
xor U22477 (N_22477,N_22389,N_22240);
nand U22478 (N_22478,N_22209,N_22283);
nand U22479 (N_22479,N_22326,N_22354);
xor U22480 (N_22480,N_22234,N_22383);
and U22481 (N_22481,N_22388,N_22226);
nor U22482 (N_22482,N_22219,N_22333);
or U22483 (N_22483,N_22355,N_22252);
xnor U22484 (N_22484,N_22256,N_22289);
and U22485 (N_22485,N_22349,N_22267);
and U22486 (N_22486,N_22300,N_22307);
or U22487 (N_22487,N_22361,N_22201);
nor U22488 (N_22488,N_22316,N_22313);
or U22489 (N_22489,N_22260,N_22314);
and U22490 (N_22490,N_22290,N_22220);
nand U22491 (N_22491,N_22346,N_22250);
and U22492 (N_22492,N_22311,N_22328);
and U22493 (N_22493,N_22282,N_22380);
nor U22494 (N_22494,N_22301,N_22237);
or U22495 (N_22495,N_22336,N_22239);
nand U22496 (N_22496,N_22330,N_22394);
nand U22497 (N_22497,N_22297,N_22304);
nand U22498 (N_22498,N_22359,N_22357);
nand U22499 (N_22499,N_22298,N_22299);
nor U22500 (N_22500,N_22249,N_22396);
nor U22501 (N_22501,N_22300,N_22381);
and U22502 (N_22502,N_22392,N_22250);
nand U22503 (N_22503,N_22346,N_22245);
nand U22504 (N_22504,N_22309,N_22212);
or U22505 (N_22505,N_22344,N_22284);
or U22506 (N_22506,N_22356,N_22267);
xnor U22507 (N_22507,N_22249,N_22311);
nand U22508 (N_22508,N_22254,N_22232);
nand U22509 (N_22509,N_22371,N_22244);
xnor U22510 (N_22510,N_22326,N_22213);
nor U22511 (N_22511,N_22285,N_22398);
and U22512 (N_22512,N_22323,N_22388);
and U22513 (N_22513,N_22391,N_22383);
and U22514 (N_22514,N_22277,N_22236);
nor U22515 (N_22515,N_22376,N_22382);
nand U22516 (N_22516,N_22306,N_22357);
nor U22517 (N_22517,N_22274,N_22224);
or U22518 (N_22518,N_22284,N_22377);
and U22519 (N_22519,N_22246,N_22278);
nor U22520 (N_22520,N_22283,N_22286);
nor U22521 (N_22521,N_22324,N_22359);
nor U22522 (N_22522,N_22238,N_22244);
nor U22523 (N_22523,N_22324,N_22312);
or U22524 (N_22524,N_22330,N_22253);
or U22525 (N_22525,N_22381,N_22390);
nor U22526 (N_22526,N_22334,N_22216);
and U22527 (N_22527,N_22284,N_22215);
nor U22528 (N_22528,N_22377,N_22399);
nor U22529 (N_22529,N_22278,N_22368);
nand U22530 (N_22530,N_22281,N_22293);
nand U22531 (N_22531,N_22346,N_22200);
and U22532 (N_22532,N_22276,N_22389);
xor U22533 (N_22533,N_22266,N_22200);
and U22534 (N_22534,N_22377,N_22391);
nand U22535 (N_22535,N_22305,N_22323);
nor U22536 (N_22536,N_22305,N_22300);
nand U22537 (N_22537,N_22201,N_22294);
nor U22538 (N_22538,N_22220,N_22219);
nor U22539 (N_22539,N_22380,N_22225);
nor U22540 (N_22540,N_22383,N_22315);
or U22541 (N_22541,N_22334,N_22256);
or U22542 (N_22542,N_22238,N_22396);
or U22543 (N_22543,N_22299,N_22375);
or U22544 (N_22544,N_22291,N_22333);
nand U22545 (N_22545,N_22236,N_22338);
nor U22546 (N_22546,N_22225,N_22306);
and U22547 (N_22547,N_22340,N_22222);
nor U22548 (N_22548,N_22348,N_22247);
xnor U22549 (N_22549,N_22368,N_22337);
and U22550 (N_22550,N_22332,N_22206);
nor U22551 (N_22551,N_22367,N_22358);
nor U22552 (N_22552,N_22228,N_22273);
nand U22553 (N_22553,N_22257,N_22396);
nor U22554 (N_22554,N_22379,N_22295);
or U22555 (N_22555,N_22372,N_22223);
nand U22556 (N_22556,N_22320,N_22304);
nand U22557 (N_22557,N_22262,N_22391);
or U22558 (N_22558,N_22315,N_22295);
nand U22559 (N_22559,N_22361,N_22245);
or U22560 (N_22560,N_22322,N_22345);
or U22561 (N_22561,N_22231,N_22377);
nand U22562 (N_22562,N_22244,N_22209);
nor U22563 (N_22563,N_22290,N_22356);
nand U22564 (N_22564,N_22323,N_22223);
or U22565 (N_22565,N_22366,N_22353);
and U22566 (N_22566,N_22348,N_22262);
nor U22567 (N_22567,N_22213,N_22236);
or U22568 (N_22568,N_22230,N_22235);
or U22569 (N_22569,N_22218,N_22263);
nand U22570 (N_22570,N_22301,N_22349);
xnor U22571 (N_22571,N_22248,N_22287);
nor U22572 (N_22572,N_22250,N_22357);
nand U22573 (N_22573,N_22220,N_22314);
and U22574 (N_22574,N_22346,N_22330);
nand U22575 (N_22575,N_22320,N_22200);
or U22576 (N_22576,N_22366,N_22295);
or U22577 (N_22577,N_22335,N_22291);
and U22578 (N_22578,N_22373,N_22301);
nand U22579 (N_22579,N_22368,N_22333);
nor U22580 (N_22580,N_22381,N_22222);
or U22581 (N_22581,N_22214,N_22383);
nand U22582 (N_22582,N_22392,N_22385);
or U22583 (N_22583,N_22257,N_22282);
and U22584 (N_22584,N_22273,N_22258);
nand U22585 (N_22585,N_22383,N_22278);
nand U22586 (N_22586,N_22368,N_22302);
or U22587 (N_22587,N_22201,N_22281);
nor U22588 (N_22588,N_22311,N_22230);
nor U22589 (N_22589,N_22349,N_22218);
nand U22590 (N_22590,N_22394,N_22327);
nor U22591 (N_22591,N_22202,N_22210);
or U22592 (N_22592,N_22325,N_22384);
and U22593 (N_22593,N_22289,N_22354);
nor U22594 (N_22594,N_22244,N_22323);
or U22595 (N_22595,N_22395,N_22384);
or U22596 (N_22596,N_22231,N_22272);
xor U22597 (N_22597,N_22325,N_22250);
and U22598 (N_22598,N_22307,N_22266);
nor U22599 (N_22599,N_22249,N_22336);
or U22600 (N_22600,N_22530,N_22599);
nor U22601 (N_22601,N_22513,N_22514);
or U22602 (N_22602,N_22416,N_22587);
or U22603 (N_22603,N_22459,N_22449);
nand U22604 (N_22604,N_22420,N_22524);
nand U22605 (N_22605,N_22438,N_22575);
xor U22606 (N_22606,N_22447,N_22490);
nor U22607 (N_22607,N_22407,N_22572);
or U22608 (N_22608,N_22552,N_22410);
xor U22609 (N_22609,N_22532,N_22501);
nand U22610 (N_22610,N_22432,N_22468);
nand U22611 (N_22611,N_22480,N_22492);
nor U22612 (N_22612,N_22458,N_22488);
and U22613 (N_22613,N_22537,N_22426);
or U22614 (N_22614,N_22486,N_22479);
xor U22615 (N_22615,N_22521,N_22429);
nor U22616 (N_22616,N_22476,N_22585);
and U22617 (N_22617,N_22564,N_22577);
nor U22618 (N_22618,N_22554,N_22460);
nor U22619 (N_22619,N_22515,N_22457);
nor U22620 (N_22620,N_22406,N_22408);
nand U22621 (N_22621,N_22519,N_22582);
or U22622 (N_22622,N_22456,N_22596);
and U22623 (N_22623,N_22547,N_22409);
nand U22624 (N_22624,N_22425,N_22414);
nor U22625 (N_22625,N_22452,N_22527);
nor U22626 (N_22626,N_22422,N_22510);
xnor U22627 (N_22627,N_22453,N_22469);
or U22628 (N_22628,N_22494,N_22566);
xnor U22629 (N_22629,N_22487,N_22463);
or U22630 (N_22630,N_22451,N_22549);
or U22631 (N_22631,N_22512,N_22499);
and U22632 (N_22632,N_22538,N_22477);
or U22633 (N_22633,N_22442,N_22567);
or U22634 (N_22634,N_22484,N_22402);
and U22635 (N_22635,N_22419,N_22470);
nand U22636 (N_22636,N_22590,N_22483);
nand U22637 (N_22637,N_22413,N_22445);
nand U22638 (N_22638,N_22466,N_22462);
and U22639 (N_22639,N_22583,N_22465);
and U22640 (N_22640,N_22529,N_22541);
nand U22641 (N_22641,N_22424,N_22544);
and U22642 (N_22642,N_22560,N_22472);
xor U22643 (N_22643,N_22412,N_22454);
and U22644 (N_22644,N_22516,N_22533);
nand U22645 (N_22645,N_22525,N_22588);
and U22646 (N_22646,N_22435,N_22534);
xnor U22647 (N_22647,N_22592,N_22471);
or U22648 (N_22648,N_22594,N_22573);
or U22649 (N_22649,N_22511,N_22474);
and U22650 (N_22650,N_22591,N_22539);
and U22651 (N_22651,N_22568,N_22440);
or U22652 (N_22652,N_22418,N_22520);
nand U22653 (N_22653,N_22598,N_22431);
nand U22654 (N_22654,N_22593,N_22423);
or U22655 (N_22655,N_22497,N_22580);
nor U22656 (N_22656,N_22421,N_22405);
xnor U22657 (N_22657,N_22411,N_22509);
and U22658 (N_22658,N_22478,N_22441);
or U22659 (N_22659,N_22565,N_22545);
and U22660 (N_22660,N_22400,N_22506);
and U22661 (N_22661,N_22546,N_22563);
and U22662 (N_22662,N_22427,N_22500);
nor U22663 (N_22663,N_22502,N_22526);
or U22664 (N_22664,N_22489,N_22428);
nor U22665 (N_22665,N_22446,N_22505);
or U22666 (N_22666,N_22455,N_22464);
nor U22667 (N_22667,N_22569,N_22576);
nor U22668 (N_22668,N_22550,N_22461);
or U22669 (N_22669,N_22473,N_22571);
nand U22670 (N_22670,N_22551,N_22548);
nand U22671 (N_22671,N_22553,N_22528);
nand U22672 (N_22672,N_22417,N_22493);
and U22673 (N_22673,N_22481,N_22584);
nor U22674 (N_22674,N_22507,N_22508);
or U22675 (N_22675,N_22491,N_22485);
nand U22676 (N_22676,N_22581,N_22522);
nand U22677 (N_22677,N_22401,N_22439);
nor U22678 (N_22678,N_22433,N_22558);
nor U22679 (N_22679,N_22403,N_22517);
nor U22680 (N_22680,N_22448,N_22574);
or U22681 (N_22681,N_22495,N_22559);
or U22682 (N_22682,N_22543,N_22415);
and U22683 (N_22683,N_22578,N_22536);
xnor U22684 (N_22684,N_22504,N_22404);
and U22685 (N_22685,N_22523,N_22434);
and U22686 (N_22686,N_22586,N_22535);
nor U22687 (N_22687,N_22444,N_22540);
and U22688 (N_22688,N_22503,N_22498);
or U22689 (N_22689,N_22467,N_22555);
nand U22690 (N_22690,N_22597,N_22589);
xnor U22691 (N_22691,N_22450,N_22518);
and U22692 (N_22692,N_22542,N_22496);
xor U22693 (N_22693,N_22475,N_22437);
nand U22694 (N_22694,N_22570,N_22561);
nand U22695 (N_22695,N_22557,N_22556);
and U22696 (N_22696,N_22443,N_22562);
nor U22697 (N_22697,N_22430,N_22482);
xor U22698 (N_22698,N_22595,N_22436);
nand U22699 (N_22699,N_22579,N_22531);
nand U22700 (N_22700,N_22434,N_22400);
or U22701 (N_22701,N_22421,N_22553);
or U22702 (N_22702,N_22552,N_22493);
nand U22703 (N_22703,N_22480,N_22406);
nand U22704 (N_22704,N_22502,N_22548);
nor U22705 (N_22705,N_22570,N_22550);
nor U22706 (N_22706,N_22490,N_22522);
nand U22707 (N_22707,N_22516,N_22508);
nand U22708 (N_22708,N_22481,N_22519);
and U22709 (N_22709,N_22569,N_22518);
or U22710 (N_22710,N_22510,N_22558);
nor U22711 (N_22711,N_22462,N_22423);
or U22712 (N_22712,N_22499,N_22457);
or U22713 (N_22713,N_22479,N_22551);
nor U22714 (N_22714,N_22584,N_22514);
nand U22715 (N_22715,N_22480,N_22573);
or U22716 (N_22716,N_22497,N_22407);
nand U22717 (N_22717,N_22413,N_22428);
and U22718 (N_22718,N_22420,N_22506);
nand U22719 (N_22719,N_22549,N_22470);
or U22720 (N_22720,N_22440,N_22557);
and U22721 (N_22721,N_22437,N_22499);
and U22722 (N_22722,N_22470,N_22445);
or U22723 (N_22723,N_22442,N_22527);
nor U22724 (N_22724,N_22530,N_22574);
nor U22725 (N_22725,N_22443,N_22439);
nand U22726 (N_22726,N_22453,N_22534);
or U22727 (N_22727,N_22526,N_22530);
xnor U22728 (N_22728,N_22587,N_22530);
nand U22729 (N_22729,N_22496,N_22474);
nand U22730 (N_22730,N_22401,N_22418);
or U22731 (N_22731,N_22429,N_22583);
nor U22732 (N_22732,N_22412,N_22455);
xor U22733 (N_22733,N_22595,N_22540);
xnor U22734 (N_22734,N_22530,N_22557);
and U22735 (N_22735,N_22597,N_22446);
xor U22736 (N_22736,N_22540,N_22422);
or U22737 (N_22737,N_22468,N_22451);
nor U22738 (N_22738,N_22425,N_22401);
nor U22739 (N_22739,N_22597,N_22568);
and U22740 (N_22740,N_22408,N_22523);
nand U22741 (N_22741,N_22468,N_22475);
or U22742 (N_22742,N_22415,N_22560);
or U22743 (N_22743,N_22509,N_22406);
nor U22744 (N_22744,N_22589,N_22593);
and U22745 (N_22745,N_22580,N_22463);
and U22746 (N_22746,N_22558,N_22496);
xnor U22747 (N_22747,N_22599,N_22593);
nand U22748 (N_22748,N_22567,N_22598);
and U22749 (N_22749,N_22536,N_22549);
or U22750 (N_22750,N_22419,N_22444);
or U22751 (N_22751,N_22494,N_22513);
and U22752 (N_22752,N_22478,N_22492);
nor U22753 (N_22753,N_22510,N_22552);
or U22754 (N_22754,N_22424,N_22459);
xor U22755 (N_22755,N_22491,N_22596);
xnor U22756 (N_22756,N_22445,N_22492);
nand U22757 (N_22757,N_22507,N_22429);
nand U22758 (N_22758,N_22485,N_22537);
or U22759 (N_22759,N_22521,N_22456);
or U22760 (N_22760,N_22419,N_22589);
or U22761 (N_22761,N_22503,N_22418);
nand U22762 (N_22762,N_22504,N_22555);
and U22763 (N_22763,N_22559,N_22422);
or U22764 (N_22764,N_22490,N_22501);
nor U22765 (N_22765,N_22546,N_22501);
and U22766 (N_22766,N_22468,N_22513);
nand U22767 (N_22767,N_22440,N_22549);
nand U22768 (N_22768,N_22533,N_22437);
or U22769 (N_22769,N_22599,N_22408);
nor U22770 (N_22770,N_22505,N_22478);
and U22771 (N_22771,N_22530,N_22467);
xnor U22772 (N_22772,N_22591,N_22522);
xor U22773 (N_22773,N_22481,N_22478);
and U22774 (N_22774,N_22471,N_22430);
or U22775 (N_22775,N_22575,N_22462);
nor U22776 (N_22776,N_22543,N_22573);
nor U22777 (N_22777,N_22563,N_22482);
nor U22778 (N_22778,N_22537,N_22464);
and U22779 (N_22779,N_22478,N_22408);
or U22780 (N_22780,N_22513,N_22543);
nand U22781 (N_22781,N_22464,N_22559);
nor U22782 (N_22782,N_22544,N_22431);
and U22783 (N_22783,N_22489,N_22426);
nand U22784 (N_22784,N_22512,N_22592);
or U22785 (N_22785,N_22416,N_22465);
nor U22786 (N_22786,N_22505,N_22406);
or U22787 (N_22787,N_22412,N_22415);
and U22788 (N_22788,N_22566,N_22578);
nand U22789 (N_22789,N_22599,N_22401);
or U22790 (N_22790,N_22479,N_22448);
and U22791 (N_22791,N_22553,N_22591);
nor U22792 (N_22792,N_22511,N_22464);
nor U22793 (N_22793,N_22413,N_22530);
xor U22794 (N_22794,N_22545,N_22516);
and U22795 (N_22795,N_22524,N_22451);
nand U22796 (N_22796,N_22586,N_22577);
nor U22797 (N_22797,N_22545,N_22561);
and U22798 (N_22798,N_22472,N_22551);
nor U22799 (N_22799,N_22503,N_22407);
or U22800 (N_22800,N_22690,N_22675);
or U22801 (N_22801,N_22662,N_22686);
nor U22802 (N_22802,N_22723,N_22617);
xor U22803 (N_22803,N_22705,N_22742);
xnor U22804 (N_22804,N_22676,N_22674);
and U22805 (N_22805,N_22740,N_22678);
nor U22806 (N_22806,N_22636,N_22658);
and U22807 (N_22807,N_22683,N_22655);
nand U22808 (N_22808,N_22672,N_22763);
or U22809 (N_22809,N_22761,N_22748);
and U22810 (N_22810,N_22665,N_22608);
nand U22811 (N_22811,N_22741,N_22651);
nand U22812 (N_22812,N_22647,N_22778);
or U22813 (N_22813,N_22762,N_22795);
or U22814 (N_22814,N_22768,N_22728);
nor U22815 (N_22815,N_22620,N_22770);
nand U22816 (N_22816,N_22746,N_22792);
or U22817 (N_22817,N_22616,N_22789);
nand U22818 (N_22818,N_22663,N_22775);
nand U22819 (N_22819,N_22718,N_22630);
and U22820 (N_22820,N_22777,N_22657);
nand U22821 (N_22821,N_22753,N_22656);
and U22822 (N_22822,N_22633,N_22760);
and U22823 (N_22823,N_22708,N_22606);
nor U22824 (N_22824,N_22769,N_22738);
nor U22825 (N_22825,N_22650,N_22684);
xor U22826 (N_22826,N_22643,N_22735);
or U22827 (N_22827,N_22783,N_22755);
xnor U22828 (N_22828,N_22612,N_22779);
or U22829 (N_22829,N_22786,N_22619);
nor U22830 (N_22830,N_22790,N_22625);
nor U22831 (N_22831,N_22693,N_22635);
and U22832 (N_22832,N_22689,N_22600);
nor U22833 (N_22833,N_22654,N_22764);
or U22834 (N_22834,N_22704,N_22745);
or U22835 (N_22835,N_22711,N_22734);
nor U22836 (N_22836,N_22751,N_22695);
and U22837 (N_22837,N_22621,N_22774);
and U22838 (N_22838,N_22709,N_22668);
nor U22839 (N_22839,N_22720,N_22759);
nand U22840 (N_22840,N_22677,N_22796);
nor U22841 (N_22841,N_22671,N_22703);
nor U22842 (N_22842,N_22785,N_22688);
nor U22843 (N_22843,N_22640,N_22702);
nor U22844 (N_22844,N_22714,N_22788);
and U22845 (N_22845,N_22696,N_22604);
nor U22846 (N_22846,N_22700,N_22772);
and U22847 (N_22847,N_22781,N_22629);
nor U22848 (N_22848,N_22730,N_22639);
or U22849 (N_22849,N_22767,N_22793);
nand U22850 (N_22850,N_22727,N_22797);
nand U22851 (N_22851,N_22729,N_22610);
nand U22852 (N_22852,N_22687,N_22713);
nand U22853 (N_22853,N_22725,N_22794);
and U22854 (N_22854,N_22724,N_22609);
and U22855 (N_22855,N_22691,N_22660);
or U22856 (N_22856,N_22638,N_22765);
and U22857 (N_22857,N_22707,N_22771);
nand U22858 (N_22858,N_22747,N_22780);
or U22859 (N_22859,N_22721,N_22782);
nand U22860 (N_22860,N_22787,N_22679);
nand U22861 (N_22861,N_22627,N_22634);
or U22862 (N_22862,N_22652,N_22737);
nand U22863 (N_22863,N_22682,N_22669);
or U22864 (N_22864,N_22766,N_22685);
nand U22865 (N_22865,N_22628,N_22692);
nor U22866 (N_22866,N_22623,N_22661);
nor U22867 (N_22867,N_22699,N_22739);
and U22868 (N_22868,N_22757,N_22642);
and U22869 (N_22869,N_22659,N_22605);
or U22870 (N_22870,N_22649,N_22618);
nand U22871 (N_22871,N_22602,N_22736);
nand U22872 (N_22872,N_22750,N_22667);
and U22873 (N_22873,N_22799,N_22613);
and U22874 (N_22874,N_22731,N_22798);
nand U22875 (N_22875,N_22615,N_22601);
nand U22876 (N_22876,N_22710,N_22743);
nand U22877 (N_22877,N_22719,N_22701);
xor U22878 (N_22878,N_22614,N_22645);
or U22879 (N_22879,N_22752,N_22744);
nor U22880 (N_22880,N_22726,N_22758);
nand U22881 (N_22881,N_22697,N_22680);
or U22882 (N_22882,N_22622,N_22784);
and U22883 (N_22883,N_22717,N_22607);
xnor U22884 (N_22884,N_22754,N_22626);
nand U22885 (N_22885,N_22732,N_22648);
nor U22886 (N_22886,N_22712,N_22715);
and U22887 (N_22887,N_22694,N_22631);
and U22888 (N_22888,N_22611,N_22733);
nand U22889 (N_22889,N_22722,N_22603);
or U22890 (N_22890,N_22653,N_22641);
nor U22891 (N_22891,N_22670,N_22664);
xor U22892 (N_22892,N_22749,N_22773);
xnor U22893 (N_22893,N_22776,N_22756);
nand U22894 (N_22894,N_22624,N_22698);
nand U22895 (N_22895,N_22637,N_22644);
nand U22896 (N_22896,N_22681,N_22673);
nor U22897 (N_22897,N_22646,N_22791);
or U22898 (N_22898,N_22706,N_22666);
and U22899 (N_22899,N_22632,N_22716);
xnor U22900 (N_22900,N_22739,N_22639);
or U22901 (N_22901,N_22787,N_22704);
nor U22902 (N_22902,N_22613,N_22687);
and U22903 (N_22903,N_22769,N_22675);
and U22904 (N_22904,N_22709,N_22779);
and U22905 (N_22905,N_22669,N_22698);
nor U22906 (N_22906,N_22656,N_22606);
and U22907 (N_22907,N_22796,N_22734);
nor U22908 (N_22908,N_22670,N_22600);
or U22909 (N_22909,N_22727,N_22757);
xnor U22910 (N_22910,N_22617,N_22774);
nor U22911 (N_22911,N_22643,N_22672);
nand U22912 (N_22912,N_22743,N_22639);
and U22913 (N_22913,N_22704,N_22772);
nand U22914 (N_22914,N_22796,N_22740);
or U22915 (N_22915,N_22692,N_22754);
nand U22916 (N_22916,N_22672,N_22789);
and U22917 (N_22917,N_22783,N_22724);
nand U22918 (N_22918,N_22649,N_22753);
or U22919 (N_22919,N_22614,N_22724);
and U22920 (N_22920,N_22656,N_22614);
or U22921 (N_22921,N_22651,N_22754);
nor U22922 (N_22922,N_22624,N_22601);
nor U22923 (N_22923,N_22712,N_22623);
nand U22924 (N_22924,N_22781,N_22636);
xor U22925 (N_22925,N_22611,N_22752);
xor U22926 (N_22926,N_22690,N_22732);
and U22927 (N_22927,N_22627,N_22749);
nor U22928 (N_22928,N_22608,N_22741);
xor U22929 (N_22929,N_22776,N_22748);
xnor U22930 (N_22930,N_22754,N_22706);
or U22931 (N_22931,N_22627,N_22678);
or U22932 (N_22932,N_22789,N_22724);
nand U22933 (N_22933,N_22614,N_22658);
nand U22934 (N_22934,N_22735,N_22668);
or U22935 (N_22935,N_22698,N_22742);
xor U22936 (N_22936,N_22792,N_22610);
nor U22937 (N_22937,N_22757,N_22734);
nand U22938 (N_22938,N_22683,N_22764);
or U22939 (N_22939,N_22668,N_22611);
nor U22940 (N_22940,N_22730,N_22718);
or U22941 (N_22941,N_22677,N_22779);
xnor U22942 (N_22942,N_22646,N_22651);
nor U22943 (N_22943,N_22676,N_22658);
nand U22944 (N_22944,N_22613,N_22733);
and U22945 (N_22945,N_22755,N_22764);
xor U22946 (N_22946,N_22755,N_22778);
nand U22947 (N_22947,N_22681,N_22601);
xor U22948 (N_22948,N_22651,N_22780);
nor U22949 (N_22949,N_22615,N_22619);
nand U22950 (N_22950,N_22651,N_22687);
or U22951 (N_22951,N_22776,N_22644);
nand U22952 (N_22952,N_22655,N_22738);
nand U22953 (N_22953,N_22733,N_22742);
or U22954 (N_22954,N_22703,N_22738);
nor U22955 (N_22955,N_22655,N_22765);
nor U22956 (N_22956,N_22715,N_22673);
nor U22957 (N_22957,N_22698,N_22797);
nand U22958 (N_22958,N_22617,N_22724);
xor U22959 (N_22959,N_22645,N_22651);
nand U22960 (N_22960,N_22769,N_22753);
nand U22961 (N_22961,N_22722,N_22623);
or U22962 (N_22962,N_22727,N_22608);
or U22963 (N_22963,N_22748,N_22740);
and U22964 (N_22964,N_22637,N_22611);
and U22965 (N_22965,N_22600,N_22765);
nor U22966 (N_22966,N_22705,N_22677);
nor U22967 (N_22967,N_22631,N_22748);
and U22968 (N_22968,N_22728,N_22712);
xor U22969 (N_22969,N_22705,N_22694);
or U22970 (N_22970,N_22646,N_22624);
xor U22971 (N_22971,N_22780,N_22717);
and U22972 (N_22972,N_22631,N_22726);
and U22973 (N_22973,N_22774,N_22752);
and U22974 (N_22974,N_22704,N_22759);
and U22975 (N_22975,N_22686,N_22776);
nand U22976 (N_22976,N_22751,N_22667);
xor U22977 (N_22977,N_22683,N_22624);
nand U22978 (N_22978,N_22797,N_22607);
nand U22979 (N_22979,N_22620,N_22778);
nor U22980 (N_22980,N_22604,N_22655);
nor U22981 (N_22981,N_22780,N_22616);
nor U22982 (N_22982,N_22686,N_22756);
nor U22983 (N_22983,N_22793,N_22649);
or U22984 (N_22984,N_22700,N_22793);
nand U22985 (N_22985,N_22757,N_22677);
or U22986 (N_22986,N_22798,N_22756);
or U22987 (N_22987,N_22729,N_22742);
and U22988 (N_22988,N_22653,N_22707);
nand U22989 (N_22989,N_22795,N_22768);
xnor U22990 (N_22990,N_22605,N_22669);
nand U22991 (N_22991,N_22691,N_22673);
and U22992 (N_22992,N_22762,N_22779);
nor U22993 (N_22993,N_22797,N_22786);
and U22994 (N_22994,N_22725,N_22602);
and U22995 (N_22995,N_22783,N_22688);
and U22996 (N_22996,N_22701,N_22752);
and U22997 (N_22997,N_22631,N_22790);
nand U22998 (N_22998,N_22771,N_22792);
nand U22999 (N_22999,N_22691,N_22633);
nand U23000 (N_23000,N_22940,N_22875);
or U23001 (N_23001,N_22840,N_22843);
nor U23002 (N_23002,N_22876,N_22932);
xnor U23003 (N_23003,N_22899,N_22996);
or U23004 (N_23004,N_22862,N_22968);
and U23005 (N_23005,N_22980,N_22837);
and U23006 (N_23006,N_22866,N_22820);
and U23007 (N_23007,N_22846,N_22823);
and U23008 (N_23008,N_22908,N_22916);
nand U23009 (N_23009,N_22879,N_22985);
and U23010 (N_23010,N_22805,N_22995);
and U23011 (N_23011,N_22841,N_22989);
nand U23012 (N_23012,N_22966,N_22835);
nand U23013 (N_23013,N_22921,N_22913);
nor U23014 (N_23014,N_22975,N_22931);
or U23015 (N_23015,N_22824,N_22850);
nand U23016 (N_23016,N_22864,N_22818);
nor U23017 (N_23017,N_22886,N_22883);
nor U23018 (N_23018,N_22830,N_22842);
nand U23019 (N_23019,N_22953,N_22873);
nand U23020 (N_23020,N_22826,N_22811);
nor U23021 (N_23021,N_22858,N_22892);
and U23022 (N_23022,N_22874,N_22915);
and U23023 (N_23023,N_22827,N_22860);
nand U23024 (N_23024,N_22926,N_22861);
and U23025 (N_23025,N_22834,N_22859);
nor U23026 (N_23026,N_22971,N_22807);
nand U23027 (N_23027,N_22952,N_22954);
nor U23028 (N_23028,N_22964,N_22895);
or U23029 (N_23029,N_22800,N_22911);
nor U23030 (N_23030,N_22813,N_22901);
xor U23031 (N_23031,N_22885,N_22918);
nor U23032 (N_23032,N_22933,N_22851);
and U23033 (N_23033,N_22986,N_22935);
or U23034 (N_23034,N_22997,N_22865);
xnor U23035 (N_23035,N_22863,N_22959);
nor U23036 (N_23036,N_22869,N_22893);
or U23037 (N_23037,N_22982,N_22888);
xnor U23038 (N_23038,N_22852,N_22829);
or U23039 (N_23039,N_22801,N_22803);
nand U23040 (N_23040,N_22853,N_22970);
and U23041 (N_23041,N_22808,N_22956);
nand U23042 (N_23042,N_22965,N_22961);
nor U23043 (N_23043,N_22878,N_22810);
or U23044 (N_23044,N_22962,N_22833);
xnor U23045 (N_23045,N_22900,N_22884);
nand U23046 (N_23046,N_22816,N_22838);
nor U23047 (N_23047,N_22922,N_22839);
or U23048 (N_23048,N_22809,N_22917);
nor U23049 (N_23049,N_22825,N_22868);
or U23050 (N_23050,N_22993,N_22806);
xnor U23051 (N_23051,N_22815,N_22944);
nor U23052 (N_23052,N_22976,N_22802);
or U23053 (N_23053,N_22949,N_22960);
nor U23054 (N_23054,N_22969,N_22974);
or U23055 (N_23055,N_22914,N_22854);
or U23056 (N_23056,N_22929,N_22882);
and U23057 (N_23057,N_22967,N_22939);
nor U23058 (N_23058,N_22828,N_22957);
nand U23059 (N_23059,N_22946,N_22924);
nor U23060 (N_23060,N_22981,N_22844);
nor U23061 (N_23061,N_22831,N_22896);
xnor U23062 (N_23062,N_22979,N_22943);
and U23063 (N_23063,N_22832,N_22906);
nand U23064 (N_23064,N_22988,N_22912);
nor U23065 (N_23065,N_22951,N_22947);
nor U23066 (N_23066,N_22978,N_22909);
nand U23067 (N_23067,N_22990,N_22910);
and U23068 (N_23068,N_22928,N_22992);
nor U23069 (N_23069,N_22905,N_22821);
xor U23070 (N_23070,N_22887,N_22867);
and U23071 (N_23071,N_22907,N_22855);
xor U23072 (N_23072,N_22856,N_22920);
and U23073 (N_23073,N_22941,N_22897);
xnor U23074 (N_23074,N_22890,N_22889);
xor U23075 (N_23075,N_22991,N_22880);
nand U23076 (N_23076,N_22958,N_22955);
nand U23077 (N_23077,N_22925,N_22881);
and U23078 (N_23078,N_22898,N_22857);
nor U23079 (N_23079,N_22973,N_22848);
or U23080 (N_23080,N_22817,N_22963);
and U23081 (N_23081,N_22923,N_22984);
nand U23082 (N_23082,N_22836,N_22819);
and U23083 (N_23083,N_22945,N_22845);
and U23084 (N_23084,N_22999,N_22927);
or U23085 (N_23085,N_22998,N_22814);
nor U23086 (N_23086,N_22894,N_22919);
and U23087 (N_23087,N_22948,N_22904);
xnor U23088 (N_23088,N_22930,N_22937);
nor U23089 (N_23089,N_22849,N_22942);
xnor U23090 (N_23090,N_22934,N_22804);
xnor U23091 (N_23091,N_22871,N_22938);
nand U23092 (N_23092,N_22877,N_22903);
nor U23093 (N_23093,N_22950,N_22812);
or U23094 (N_23094,N_22870,N_22822);
nand U23095 (N_23095,N_22994,N_22872);
nand U23096 (N_23096,N_22972,N_22902);
nor U23097 (N_23097,N_22891,N_22987);
or U23098 (N_23098,N_22977,N_22983);
and U23099 (N_23099,N_22847,N_22936);
nor U23100 (N_23100,N_22978,N_22902);
or U23101 (N_23101,N_22920,N_22874);
and U23102 (N_23102,N_22894,N_22941);
nand U23103 (N_23103,N_22921,N_22938);
nor U23104 (N_23104,N_22841,N_22801);
xnor U23105 (N_23105,N_22831,N_22858);
and U23106 (N_23106,N_22873,N_22895);
and U23107 (N_23107,N_22910,N_22875);
nor U23108 (N_23108,N_22911,N_22971);
and U23109 (N_23109,N_22810,N_22952);
and U23110 (N_23110,N_22865,N_22844);
nor U23111 (N_23111,N_22899,N_22924);
and U23112 (N_23112,N_22974,N_22991);
nor U23113 (N_23113,N_22884,N_22989);
nand U23114 (N_23114,N_22836,N_22840);
or U23115 (N_23115,N_22935,N_22872);
xnor U23116 (N_23116,N_22948,N_22906);
or U23117 (N_23117,N_22972,N_22910);
or U23118 (N_23118,N_22852,N_22928);
nand U23119 (N_23119,N_22844,N_22963);
nand U23120 (N_23120,N_22907,N_22875);
nand U23121 (N_23121,N_22892,N_22814);
and U23122 (N_23122,N_22968,N_22939);
nand U23123 (N_23123,N_22828,N_22930);
nor U23124 (N_23124,N_22822,N_22976);
nor U23125 (N_23125,N_22908,N_22867);
or U23126 (N_23126,N_22924,N_22937);
nor U23127 (N_23127,N_22964,N_22940);
or U23128 (N_23128,N_22830,N_22912);
nand U23129 (N_23129,N_22860,N_22818);
nand U23130 (N_23130,N_22945,N_22880);
and U23131 (N_23131,N_22950,N_22913);
nand U23132 (N_23132,N_22988,N_22924);
and U23133 (N_23133,N_22900,N_22955);
and U23134 (N_23134,N_22920,N_22830);
or U23135 (N_23135,N_22859,N_22944);
and U23136 (N_23136,N_22969,N_22878);
nand U23137 (N_23137,N_22994,N_22819);
nand U23138 (N_23138,N_22856,N_22868);
or U23139 (N_23139,N_22911,N_22864);
xor U23140 (N_23140,N_22916,N_22884);
and U23141 (N_23141,N_22829,N_22888);
nor U23142 (N_23142,N_22811,N_22895);
nor U23143 (N_23143,N_22955,N_22918);
xor U23144 (N_23144,N_22903,N_22824);
xnor U23145 (N_23145,N_22986,N_22888);
nor U23146 (N_23146,N_22905,N_22808);
nand U23147 (N_23147,N_22841,N_22914);
nor U23148 (N_23148,N_22927,N_22923);
nor U23149 (N_23149,N_22932,N_22904);
nor U23150 (N_23150,N_22987,N_22807);
nor U23151 (N_23151,N_22975,N_22843);
nand U23152 (N_23152,N_22847,N_22825);
xor U23153 (N_23153,N_22989,N_22887);
nand U23154 (N_23154,N_22822,N_22927);
nand U23155 (N_23155,N_22921,N_22861);
and U23156 (N_23156,N_22807,N_22965);
or U23157 (N_23157,N_22905,N_22859);
xnor U23158 (N_23158,N_22854,N_22943);
or U23159 (N_23159,N_22918,N_22812);
or U23160 (N_23160,N_22952,N_22936);
or U23161 (N_23161,N_22961,N_22924);
and U23162 (N_23162,N_22821,N_22878);
nand U23163 (N_23163,N_22892,N_22891);
nand U23164 (N_23164,N_22980,N_22855);
or U23165 (N_23165,N_22982,N_22829);
nand U23166 (N_23166,N_22819,N_22965);
or U23167 (N_23167,N_22930,N_22910);
and U23168 (N_23168,N_22948,N_22848);
nor U23169 (N_23169,N_22926,N_22903);
or U23170 (N_23170,N_22881,N_22970);
and U23171 (N_23171,N_22834,N_22892);
nor U23172 (N_23172,N_22862,N_22942);
or U23173 (N_23173,N_22800,N_22865);
nor U23174 (N_23174,N_22809,N_22971);
nand U23175 (N_23175,N_22811,N_22969);
xor U23176 (N_23176,N_22880,N_22850);
or U23177 (N_23177,N_22985,N_22996);
or U23178 (N_23178,N_22927,N_22917);
nor U23179 (N_23179,N_22875,N_22900);
nor U23180 (N_23180,N_22948,N_22974);
nand U23181 (N_23181,N_22842,N_22942);
nand U23182 (N_23182,N_22816,N_22961);
or U23183 (N_23183,N_22909,N_22986);
nor U23184 (N_23184,N_22915,N_22996);
nor U23185 (N_23185,N_22884,N_22990);
xnor U23186 (N_23186,N_22953,N_22843);
or U23187 (N_23187,N_22966,N_22869);
nor U23188 (N_23188,N_22992,N_22850);
and U23189 (N_23189,N_22957,N_22857);
nor U23190 (N_23190,N_22932,N_22901);
nor U23191 (N_23191,N_22877,N_22931);
nand U23192 (N_23192,N_22861,N_22830);
or U23193 (N_23193,N_22943,N_22830);
nor U23194 (N_23194,N_22811,N_22878);
nor U23195 (N_23195,N_22803,N_22829);
and U23196 (N_23196,N_22867,N_22968);
or U23197 (N_23197,N_22815,N_22866);
and U23198 (N_23198,N_22991,N_22894);
nand U23199 (N_23199,N_22916,N_22981);
and U23200 (N_23200,N_23129,N_23181);
and U23201 (N_23201,N_23184,N_23143);
and U23202 (N_23202,N_23060,N_23078);
nand U23203 (N_23203,N_23095,N_23100);
nand U23204 (N_23204,N_23097,N_23120);
and U23205 (N_23205,N_23160,N_23132);
xnor U23206 (N_23206,N_23191,N_23170);
nand U23207 (N_23207,N_23071,N_23063);
or U23208 (N_23208,N_23001,N_23152);
nand U23209 (N_23209,N_23192,N_23065);
nor U23210 (N_23210,N_23026,N_23146);
and U23211 (N_23211,N_23131,N_23049);
nand U23212 (N_23212,N_23188,N_23115);
nand U23213 (N_23213,N_23122,N_23157);
nor U23214 (N_23214,N_23003,N_23090);
or U23215 (N_23215,N_23150,N_23123);
and U23216 (N_23216,N_23045,N_23105);
nand U23217 (N_23217,N_23187,N_23064);
xnor U23218 (N_23218,N_23000,N_23077);
xor U23219 (N_23219,N_23037,N_23052);
and U23220 (N_23220,N_23135,N_23020);
or U23221 (N_23221,N_23008,N_23177);
and U23222 (N_23222,N_23139,N_23074);
xor U23223 (N_23223,N_23108,N_23125);
or U23224 (N_23224,N_23031,N_23007);
and U23225 (N_23225,N_23002,N_23009);
and U23226 (N_23226,N_23185,N_23173);
and U23227 (N_23227,N_23076,N_23018);
and U23228 (N_23228,N_23155,N_23094);
nor U23229 (N_23229,N_23016,N_23085);
or U23230 (N_23230,N_23089,N_23101);
and U23231 (N_23231,N_23021,N_23156);
nand U23232 (N_23232,N_23196,N_23011);
and U23233 (N_23233,N_23199,N_23015);
nor U23234 (N_23234,N_23180,N_23172);
and U23235 (N_23235,N_23004,N_23092);
nor U23236 (N_23236,N_23036,N_23055);
nand U23237 (N_23237,N_23186,N_23151);
nand U23238 (N_23238,N_23083,N_23112);
nor U23239 (N_23239,N_23145,N_23117);
or U23240 (N_23240,N_23033,N_23168);
and U23241 (N_23241,N_23161,N_23118);
or U23242 (N_23242,N_23107,N_23133);
and U23243 (N_23243,N_23058,N_23111);
nand U23244 (N_23244,N_23126,N_23017);
nor U23245 (N_23245,N_23134,N_23179);
xnor U23246 (N_23246,N_23121,N_23022);
or U23247 (N_23247,N_23029,N_23127);
and U23248 (N_23248,N_23164,N_23153);
nand U23249 (N_23249,N_23110,N_23194);
nor U23250 (N_23250,N_23091,N_23013);
or U23251 (N_23251,N_23030,N_23119);
xor U23252 (N_23252,N_23096,N_23072);
or U23253 (N_23253,N_23136,N_23023);
and U23254 (N_23254,N_23159,N_23104);
and U23255 (N_23255,N_23070,N_23027);
and U23256 (N_23256,N_23178,N_23182);
or U23257 (N_23257,N_23174,N_23098);
nor U23258 (N_23258,N_23106,N_23005);
nor U23259 (N_23259,N_23050,N_23189);
and U23260 (N_23260,N_23066,N_23041);
nand U23261 (N_23261,N_23048,N_23056);
xor U23262 (N_23262,N_23025,N_23038);
and U23263 (N_23263,N_23044,N_23138);
and U23264 (N_23264,N_23158,N_23099);
xnor U23265 (N_23265,N_23062,N_23024);
or U23266 (N_23266,N_23079,N_23040);
nand U23267 (N_23267,N_23197,N_23102);
or U23268 (N_23268,N_23046,N_23190);
and U23269 (N_23269,N_23080,N_23103);
or U23270 (N_23270,N_23147,N_23148);
nand U23271 (N_23271,N_23128,N_23019);
xor U23272 (N_23272,N_23034,N_23176);
xnor U23273 (N_23273,N_23028,N_23198);
or U23274 (N_23274,N_23081,N_23175);
and U23275 (N_23275,N_23053,N_23061);
xnor U23276 (N_23276,N_23142,N_23043);
nand U23277 (N_23277,N_23012,N_23082);
nor U23278 (N_23278,N_23059,N_23109);
nor U23279 (N_23279,N_23141,N_23116);
nor U23280 (N_23280,N_23165,N_23069);
or U23281 (N_23281,N_23163,N_23039);
or U23282 (N_23282,N_23162,N_23195);
or U23283 (N_23283,N_23047,N_23073);
nor U23284 (N_23284,N_23154,N_23051);
and U23285 (N_23285,N_23171,N_23010);
nand U23286 (N_23286,N_23114,N_23093);
nor U23287 (N_23287,N_23113,N_23068);
xor U23288 (N_23288,N_23032,N_23035);
nor U23289 (N_23289,N_23087,N_23006);
nor U23290 (N_23290,N_23193,N_23167);
nor U23291 (N_23291,N_23067,N_23075);
nor U23292 (N_23292,N_23014,N_23140);
nand U23293 (N_23293,N_23169,N_23144);
nand U23294 (N_23294,N_23137,N_23084);
xor U23295 (N_23295,N_23166,N_23086);
and U23296 (N_23296,N_23057,N_23183);
nand U23297 (N_23297,N_23054,N_23088);
and U23298 (N_23298,N_23124,N_23149);
or U23299 (N_23299,N_23042,N_23130);
nor U23300 (N_23300,N_23020,N_23084);
or U23301 (N_23301,N_23138,N_23186);
nor U23302 (N_23302,N_23077,N_23032);
or U23303 (N_23303,N_23089,N_23087);
nand U23304 (N_23304,N_23185,N_23071);
nand U23305 (N_23305,N_23090,N_23080);
and U23306 (N_23306,N_23109,N_23018);
or U23307 (N_23307,N_23139,N_23157);
nand U23308 (N_23308,N_23187,N_23093);
and U23309 (N_23309,N_23035,N_23159);
nand U23310 (N_23310,N_23135,N_23189);
or U23311 (N_23311,N_23172,N_23112);
or U23312 (N_23312,N_23127,N_23040);
and U23313 (N_23313,N_23155,N_23008);
nand U23314 (N_23314,N_23046,N_23042);
and U23315 (N_23315,N_23021,N_23117);
or U23316 (N_23316,N_23147,N_23078);
xor U23317 (N_23317,N_23139,N_23090);
nand U23318 (N_23318,N_23062,N_23187);
or U23319 (N_23319,N_23060,N_23187);
or U23320 (N_23320,N_23051,N_23023);
or U23321 (N_23321,N_23002,N_23187);
and U23322 (N_23322,N_23173,N_23086);
nor U23323 (N_23323,N_23176,N_23187);
nand U23324 (N_23324,N_23138,N_23191);
or U23325 (N_23325,N_23127,N_23188);
xnor U23326 (N_23326,N_23169,N_23115);
nor U23327 (N_23327,N_23171,N_23040);
nand U23328 (N_23328,N_23038,N_23171);
nand U23329 (N_23329,N_23120,N_23075);
or U23330 (N_23330,N_23145,N_23134);
nor U23331 (N_23331,N_23019,N_23161);
or U23332 (N_23332,N_23050,N_23169);
nand U23333 (N_23333,N_23164,N_23092);
nand U23334 (N_23334,N_23048,N_23131);
nor U23335 (N_23335,N_23131,N_23091);
nand U23336 (N_23336,N_23024,N_23139);
or U23337 (N_23337,N_23049,N_23065);
nor U23338 (N_23338,N_23034,N_23175);
or U23339 (N_23339,N_23168,N_23006);
and U23340 (N_23340,N_23112,N_23084);
xor U23341 (N_23341,N_23039,N_23016);
nand U23342 (N_23342,N_23107,N_23153);
nor U23343 (N_23343,N_23126,N_23091);
nand U23344 (N_23344,N_23061,N_23035);
nand U23345 (N_23345,N_23080,N_23146);
nor U23346 (N_23346,N_23074,N_23094);
or U23347 (N_23347,N_23056,N_23003);
nor U23348 (N_23348,N_23137,N_23070);
nor U23349 (N_23349,N_23013,N_23098);
or U23350 (N_23350,N_23182,N_23107);
nor U23351 (N_23351,N_23147,N_23045);
nor U23352 (N_23352,N_23193,N_23062);
and U23353 (N_23353,N_23114,N_23083);
or U23354 (N_23354,N_23134,N_23036);
nor U23355 (N_23355,N_23158,N_23184);
and U23356 (N_23356,N_23114,N_23033);
nor U23357 (N_23357,N_23192,N_23171);
nor U23358 (N_23358,N_23024,N_23023);
or U23359 (N_23359,N_23154,N_23183);
or U23360 (N_23360,N_23082,N_23033);
xnor U23361 (N_23361,N_23026,N_23121);
and U23362 (N_23362,N_23072,N_23049);
and U23363 (N_23363,N_23009,N_23168);
and U23364 (N_23364,N_23140,N_23034);
nand U23365 (N_23365,N_23051,N_23167);
xnor U23366 (N_23366,N_23101,N_23115);
or U23367 (N_23367,N_23052,N_23171);
nor U23368 (N_23368,N_23029,N_23110);
nand U23369 (N_23369,N_23196,N_23075);
or U23370 (N_23370,N_23072,N_23087);
or U23371 (N_23371,N_23194,N_23021);
nand U23372 (N_23372,N_23132,N_23085);
or U23373 (N_23373,N_23001,N_23141);
nand U23374 (N_23374,N_23084,N_23073);
nand U23375 (N_23375,N_23034,N_23151);
xor U23376 (N_23376,N_23033,N_23000);
nor U23377 (N_23377,N_23195,N_23146);
or U23378 (N_23378,N_23006,N_23042);
or U23379 (N_23379,N_23054,N_23000);
nor U23380 (N_23380,N_23024,N_23001);
or U23381 (N_23381,N_23159,N_23069);
nand U23382 (N_23382,N_23076,N_23149);
and U23383 (N_23383,N_23004,N_23150);
or U23384 (N_23384,N_23109,N_23160);
and U23385 (N_23385,N_23195,N_23066);
nor U23386 (N_23386,N_23198,N_23068);
nor U23387 (N_23387,N_23044,N_23131);
nand U23388 (N_23388,N_23048,N_23190);
or U23389 (N_23389,N_23019,N_23028);
nor U23390 (N_23390,N_23061,N_23065);
nand U23391 (N_23391,N_23040,N_23047);
and U23392 (N_23392,N_23164,N_23029);
nand U23393 (N_23393,N_23147,N_23019);
and U23394 (N_23394,N_23129,N_23027);
nor U23395 (N_23395,N_23119,N_23161);
nor U23396 (N_23396,N_23101,N_23199);
nor U23397 (N_23397,N_23185,N_23003);
nor U23398 (N_23398,N_23107,N_23108);
and U23399 (N_23399,N_23044,N_23029);
nand U23400 (N_23400,N_23204,N_23350);
nor U23401 (N_23401,N_23359,N_23277);
nand U23402 (N_23402,N_23239,N_23345);
nand U23403 (N_23403,N_23255,N_23298);
or U23404 (N_23404,N_23327,N_23253);
and U23405 (N_23405,N_23348,N_23258);
or U23406 (N_23406,N_23302,N_23280);
nand U23407 (N_23407,N_23294,N_23281);
nand U23408 (N_23408,N_23392,N_23343);
and U23409 (N_23409,N_23355,N_23293);
xnor U23410 (N_23410,N_23214,N_23238);
nand U23411 (N_23411,N_23310,N_23220);
and U23412 (N_23412,N_23358,N_23396);
and U23413 (N_23413,N_23289,N_23334);
xnor U23414 (N_23414,N_23306,N_23329);
or U23415 (N_23415,N_23330,N_23398);
nor U23416 (N_23416,N_23221,N_23228);
and U23417 (N_23417,N_23248,N_23372);
or U23418 (N_23418,N_23260,N_23278);
nor U23419 (N_23419,N_23378,N_23215);
and U23420 (N_23420,N_23271,N_23200);
nand U23421 (N_23421,N_23257,N_23326);
and U23422 (N_23422,N_23344,N_23320);
and U23423 (N_23423,N_23380,N_23244);
or U23424 (N_23424,N_23219,N_23242);
and U23425 (N_23425,N_23365,N_23331);
or U23426 (N_23426,N_23216,N_23399);
or U23427 (N_23427,N_23357,N_23384);
nor U23428 (N_23428,N_23207,N_23375);
and U23429 (N_23429,N_23367,N_23395);
nand U23430 (N_23430,N_23376,N_23362);
nor U23431 (N_23431,N_23314,N_23337);
xor U23432 (N_23432,N_23287,N_23387);
nor U23433 (N_23433,N_23394,N_23364);
nand U23434 (N_23434,N_23341,N_23299);
or U23435 (N_23435,N_23373,N_23241);
or U23436 (N_23436,N_23285,N_23232);
nand U23437 (N_23437,N_23203,N_23231);
nor U23438 (N_23438,N_23324,N_23304);
and U23439 (N_23439,N_23249,N_23284);
nand U23440 (N_23440,N_23230,N_23332);
nor U23441 (N_23441,N_23206,N_23300);
xor U23442 (N_23442,N_23322,N_23247);
nor U23443 (N_23443,N_23295,N_23223);
and U23444 (N_23444,N_23208,N_23256);
nand U23445 (N_23445,N_23340,N_23273);
nand U23446 (N_23446,N_23233,N_23316);
or U23447 (N_23447,N_23390,N_23272);
nor U23448 (N_23448,N_23202,N_23279);
nand U23449 (N_23449,N_23290,N_23296);
or U23450 (N_23450,N_23303,N_23276);
and U23451 (N_23451,N_23269,N_23356);
nand U23452 (N_23452,N_23381,N_23385);
or U23453 (N_23453,N_23313,N_23268);
and U23454 (N_23454,N_23319,N_23307);
and U23455 (N_23455,N_23318,N_23379);
or U23456 (N_23456,N_23226,N_23229);
xor U23457 (N_23457,N_23351,N_23235);
nor U23458 (N_23458,N_23267,N_23224);
nor U23459 (N_23459,N_23274,N_23368);
nor U23460 (N_23460,N_23270,N_23251);
or U23461 (N_23461,N_23371,N_23265);
and U23462 (N_23462,N_23237,N_23377);
and U23463 (N_23463,N_23245,N_23336);
and U23464 (N_23464,N_23338,N_23339);
and U23465 (N_23465,N_23225,N_23397);
nor U23466 (N_23466,N_23212,N_23353);
nor U23467 (N_23467,N_23393,N_23315);
and U23468 (N_23468,N_23209,N_23370);
nand U23469 (N_23469,N_23236,N_23361);
nor U23470 (N_23470,N_23264,N_23389);
nor U23471 (N_23471,N_23325,N_23266);
or U23472 (N_23472,N_23386,N_23227);
and U23473 (N_23473,N_23282,N_23305);
or U23474 (N_23474,N_23342,N_23309);
nor U23475 (N_23475,N_23301,N_23391);
or U23476 (N_23476,N_23354,N_23311);
nor U23477 (N_23477,N_23288,N_23323);
or U23478 (N_23478,N_23308,N_23328);
nor U23479 (N_23479,N_23211,N_23360);
nand U23480 (N_23480,N_23259,N_23297);
and U23481 (N_23481,N_23383,N_23275);
nand U23482 (N_23482,N_23374,N_23250);
nand U23483 (N_23483,N_23222,N_23218);
or U23484 (N_23484,N_23292,N_23261);
xor U23485 (N_23485,N_23217,N_23201);
nand U23486 (N_23486,N_23317,N_23254);
nand U23487 (N_23487,N_23349,N_23333);
and U23488 (N_23488,N_23240,N_23286);
xor U23489 (N_23489,N_23388,N_23246);
or U23490 (N_23490,N_23263,N_23346);
and U23491 (N_23491,N_23213,N_23252);
nand U23492 (N_23492,N_23234,N_23366);
nor U23493 (N_23493,N_23262,N_23352);
nor U23494 (N_23494,N_23243,N_23283);
or U23495 (N_23495,N_23291,N_23321);
nor U23496 (N_23496,N_23312,N_23335);
nand U23497 (N_23497,N_23347,N_23363);
or U23498 (N_23498,N_23369,N_23210);
and U23499 (N_23499,N_23205,N_23382);
nand U23500 (N_23500,N_23346,N_23371);
and U23501 (N_23501,N_23218,N_23368);
nor U23502 (N_23502,N_23244,N_23362);
and U23503 (N_23503,N_23238,N_23228);
or U23504 (N_23504,N_23397,N_23395);
or U23505 (N_23505,N_23329,N_23327);
nand U23506 (N_23506,N_23274,N_23212);
nor U23507 (N_23507,N_23343,N_23209);
nor U23508 (N_23508,N_23383,N_23247);
nand U23509 (N_23509,N_23297,N_23232);
and U23510 (N_23510,N_23305,N_23313);
nor U23511 (N_23511,N_23339,N_23299);
and U23512 (N_23512,N_23208,N_23358);
and U23513 (N_23513,N_23263,N_23259);
or U23514 (N_23514,N_23216,N_23317);
nand U23515 (N_23515,N_23350,N_23206);
and U23516 (N_23516,N_23313,N_23392);
nor U23517 (N_23517,N_23336,N_23212);
or U23518 (N_23518,N_23352,N_23333);
nand U23519 (N_23519,N_23398,N_23373);
nor U23520 (N_23520,N_23241,N_23392);
nand U23521 (N_23521,N_23286,N_23283);
or U23522 (N_23522,N_23305,N_23343);
and U23523 (N_23523,N_23290,N_23354);
and U23524 (N_23524,N_23272,N_23332);
and U23525 (N_23525,N_23395,N_23244);
nor U23526 (N_23526,N_23340,N_23265);
or U23527 (N_23527,N_23343,N_23246);
nand U23528 (N_23528,N_23213,N_23362);
nor U23529 (N_23529,N_23200,N_23335);
and U23530 (N_23530,N_23295,N_23336);
nand U23531 (N_23531,N_23257,N_23244);
and U23532 (N_23532,N_23238,N_23325);
or U23533 (N_23533,N_23249,N_23377);
nor U23534 (N_23534,N_23205,N_23288);
and U23535 (N_23535,N_23353,N_23330);
nor U23536 (N_23536,N_23234,N_23264);
nand U23537 (N_23537,N_23332,N_23334);
or U23538 (N_23538,N_23234,N_23227);
or U23539 (N_23539,N_23230,N_23386);
and U23540 (N_23540,N_23212,N_23397);
nand U23541 (N_23541,N_23218,N_23286);
nor U23542 (N_23542,N_23259,N_23336);
or U23543 (N_23543,N_23326,N_23253);
or U23544 (N_23544,N_23360,N_23324);
nand U23545 (N_23545,N_23223,N_23319);
or U23546 (N_23546,N_23357,N_23205);
and U23547 (N_23547,N_23217,N_23292);
nand U23548 (N_23548,N_23335,N_23234);
xnor U23549 (N_23549,N_23363,N_23292);
and U23550 (N_23550,N_23249,N_23209);
or U23551 (N_23551,N_23343,N_23336);
and U23552 (N_23552,N_23397,N_23256);
or U23553 (N_23553,N_23361,N_23387);
and U23554 (N_23554,N_23261,N_23267);
nor U23555 (N_23555,N_23369,N_23209);
nor U23556 (N_23556,N_23352,N_23322);
nand U23557 (N_23557,N_23392,N_23257);
or U23558 (N_23558,N_23208,N_23291);
or U23559 (N_23559,N_23313,N_23251);
xor U23560 (N_23560,N_23243,N_23236);
nor U23561 (N_23561,N_23244,N_23304);
xor U23562 (N_23562,N_23389,N_23212);
or U23563 (N_23563,N_23352,N_23381);
or U23564 (N_23564,N_23356,N_23298);
nand U23565 (N_23565,N_23378,N_23261);
and U23566 (N_23566,N_23367,N_23281);
or U23567 (N_23567,N_23262,N_23321);
xnor U23568 (N_23568,N_23277,N_23341);
nand U23569 (N_23569,N_23291,N_23214);
and U23570 (N_23570,N_23229,N_23248);
xor U23571 (N_23571,N_23318,N_23369);
or U23572 (N_23572,N_23333,N_23232);
nand U23573 (N_23573,N_23208,N_23382);
or U23574 (N_23574,N_23339,N_23253);
or U23575 (N_23575,N_23327,N_23225);
or U23576 (N_23576,N_23371,N_23279);
nand U23577 (N_23577,N_23331,N_23363);
and U23578 (N_23578,N_23219,N_23201);
nand U23579 (N_23579,N_23300,N_23363);
xnor U23580 (N_23580,N_23349,N_23286);
nor U23581 (N_23581,N_23200,N_23395);
or U23582 (N_23582,N_23370,N_23202);
nand U23583 (N_23583,N_23339,N_23238);
and U23584 (N_23584,N_23397,N_23220);
xnor U23585 (N_23585,N_23334,N_23331);
nor U23586 (N_23586,N_23321,N_23251);
nand U23587 (N_23587,N_23288,N_23322);
nand U23588 (N_23588,N_23369,N_23277);
xnor U23589 (N_23589,N_23325,N_23349);
xnor U23590 (N_23590,N_23304,N_23243);
xor U23591 (N_23591,N_23287,N_23297);
nand U23592 (N_23592,N_23378,N_23394);
xor U23593 (N_23593,N_23216,N_23210);
xnor U23594 (N_23594,N_23388,N_23247);
nand U23595 (N_23595,N_23221,N_23277);
nand U23596 (N_23596,N_23370,N_23283);
or U23597 (N_23597,N_23237,N_23258);
nor U23598 (N_23598,N_23334,N_23306);
nor U23599 (N_23599,N_23231,N_23296);
nor U23600 (N_23600,N_23511,N_23512);
and U23601 (N_23601,N_23552,N_23565);
and U23602 (N_23602,N_23592,N_23524);
nand U23603 (N_23603,N_23556,N_23437);
nand U23604 (N_23604,N_23443,N_23466);
or U23605 (N_23605,N_23589,N_23498);
and U23606 (N_23606,N_23561,N_23471);
nand U23607 (N_23607,N_23584,N_23518);
nand U23608 (N_23608,N_23405,N_23583);
or U23609 (N_23609,N_23539,N_23429);
and U23610 (N_23610,N_23529,N_23541);
xor U23611 (N_23611,N_23425,N_23407);
nand U23612 (N_23612,N_23523,N_23450);
nor U23613 (N_23613,N_23540,N_23567);
or U23614 (N_23614,N_23557,N_23482);
and U23615 (N_23615,N_23416,N_23554);
nor U23616 (N_23616,N_23560,N_23453);
or U23617 (N_23617,N_23445,N_23456);
xor U23618 (N_23618,N_23480,N_23506);
nor U23619 (N_23619,N_23486,N_23496);
or U23620 (N_23620,N_23444,N_23481);
nor U23621 (N_23621,N_23545,N_23479);
nand U23622 (N_23622,N_23517,N_23454);
nand U23623 (N_23623,N_23535,N_23546);
or U23624 (N_23624,N_23504,N_23412);
nor U23625 (N_23625,N_23566,N_23497);
and U23626 (N_23626,N_23510,N_23598);
and U23627 (N_23627,N_23428,N_23577);
nor U23628 (N_23628,N_23503,N_23528);
and U23629 (N_23629,N_23418,N_23562);
nand U23630 (N_23630,N_23489,N_23502);
xnor U23631 (N_23631,N_23469,N_23483);
nor U23632 (N_23632,N_23433,N_23575);
xor U23633 (N_23633,N_23423,N_23551);
or U23634 (N_23634,N_23446,N_23475);
nor U23635 (N_23635,N_23586,N_23599);
xor U23636 (N_23636,N_23465,N_23495);
nand U23637 (N_23637,N_23572,N_23432);
or U23638 (N_23638,N_23464,N_23521);
xor U23639 (N_23639,N_23441,N_23404);
or U23640 (N_23640,N_23564,N_23537);
nand U23641 (N_23641,N_23544,N_23526);
nor U23642 (N_23642,N_23403,N_23547);
or U23643 (N_23643,N_23595,N_23485);
nand U23644 (N_23644,N_23500,N_23542);
nor U23645 (N_23645,N_23491,N_23580);
or U23646 (N_23646,N_23415,N_23513);
nor U23647 (N_23647,N_23499,N_23520);
or U23648 (N_23648,N_23474,N_23417);
and U23649 (N_23649,N_23484,N_23531);
nor U23650 (N_23650,N_23477,N_23525);
xor U23651 (N_23651,N_23587,N_23514);
nor U23652 (N_23652,N_23509,N_23596);
nor U23653 (N_23653,N_23409,N_23530);
nor U23654 (N_23654,N_23436,N_23558);
or U23655 (N_23655,N_23424,N_23550);
xnor U23656 (N_23656,N_23588,N_23494);
nand U23657 (N_23657,N_23440,N_23515);
nor U23658 (N_23658,N_23508,N_23419);
nand U23659 (N_23659,N_23597,N_23411);
nor U23660 (N_23660,N_23548,N_23533);
nor U23661 (N_23661,N_23473,N_23420);
or U23662 (N_23662,N_23408,N_23488);
and U23663 (N_23663,N_23459,N_23449);
or U23664 (N_23664,N_23532,N_23461);
and U23665 (N_23665,N_23538,N_23573);
xnor U23666 (N_23666,N_23413,N_23468);
or U23667 (N_23667,N_23593,N_23406);
nor U23668 (N_23668,N_23568,N_23549);
nand U23669 (N_23669,N_23578,N_23579);
and U23670 (N_23670,N_23435,N_23426);
nor U23671 (N_23671,N_23458,N_23431);
xnor U23672 (N_23672,N_23569,N_23448);
nor U23673 (N_23673,N_23576,N_23492);
or U23674 (N_23674,N_23559,N_23421);
xor U23675 (N_23675,N_23427,N_23455);
and U23676 (N_23676,N_23400,N_23527);
xor U23677 (N_23677,N_23505,N_23478);
and U23678 (N_23678,N_23594,N_23463);
nand U23679 (N_23679,N_23472,N_23581);
nor U23680 (N_23680,N_23470,N_23574);
or U23681 (N_23681,N_23536,N_23414);
nor U23682 (N_23682,N_23507,N_23534);
nor U23683 (N_23683,N_23582,N_23563);
nor U23684 (N_23684,N_23516,N_23410);
nor U23685 (N_23685,N_23501,N_23490);
nor U23686 (N_23686,N_23571,N_23438);
nand U23687 (N_23687,N_23434,N_23439);
or U23688 (N_23688,N_23555,N_23457);
nor U23689 (N_23689,N_23585,N_23570);
and U23690 (N_23690,N_23590,N_23493);
or U23691 (N_23691,N_23543,N_23447);
nand U23692 (N_23692,N_23519,N_23553);
nor U23693 (N_23693,N_23467,N_23522);
nand U23694 (N_23694,N_23422,N_23401);
xor U23695 (N_23695,N_23451,N_23402);
or U23696 (N_23696,N_23476,N_23442);
nand U23697 (N_23697,N_23591,N_23487);
nor U23698 (N_23698,N_23462,N_23452);
nor U23699 (N_23699,N_23430,N_23460);
nor U23700 (N_23700,N_23561,N_23450);
nor U23701 (N_23701,N_23482,N_23416);
or U23702 (N_23702,N_23419,N_23433);
or U23703 (N_23703,N_23400,N_23426);
or U23704 (N_23704,N_23572,N_23588);
nand U23705 (N_23705,N_23479,N_23445);
nand U23706 (N_23706,N_23585,N_23454);
and U23707 (N_23707,N_23489,N_23548);
nand U23708 (N_23708,N_23561,N_23483);
xor U23709 (N_23709,N_23438,N_23466);
and U23710 (N_23710,N_23450,N_23559);
and U23711 (N_23711,N_23481,N_23533);
nor U23712 (N_23712,N_23487,N_23526);
or U23713 (N_23713,N_23596,N_23511);
nor U23714 (N_23714,N_23422,N_23468);
and U23715 (N_23715,N_23512,N_23508);
or U23716 (N_23716,N_23432,N_23486);
and U23717 (N_23717,N_23521,N_23458);
and U23718 (N_23718,N_23462,N_23494);
nand U23719 (N_23719,N_23556,N_23515);
nor U23720 (N_23720,N_23596,N_23537);
nor U23721 (N_23721,N_23499,N_23429);
nand U23722 (N_23722,N_23511,N_23416);
xor U23723 (N_23723,N_23457,N_23479);
nand U23724 (N_23724,N_23527,N_23519);
nand U23725 (N_23725,N_23408,N_23503);
or U23726 (N_23726,N_23555,N_23416);
nand U23727 (N_23727,N_23572,N_23404);
nand U23728 (N_23728,N_23494,N_23497);
nor U23729 (N_23729,N_23484,N_23585);
or U23730 (N_23730,N_23596,N_23559);
and U23731 (N_23731,N_23487,N_23438);
nor U23732 (N_23732,N_23593,N_23425);
nand U23733 (N_23733,N_23497,N_23455);
nor U23734 (N_23734,N_23435,N_23405);
nand U23735 (N_23735,N_23541,N_23502);
xnor U23736 (N_23736,N_23534,N_23563);
or U23737 (N_23737,N_23596,N_23470);
or U23738 (N_23738,N_23438,N_23589);
nor U23739 (N_23739,N_23504,N_23402);
or U23740 (N_23740,N_23504,N_23564);
and U23741 (N_23741,N_23471,N_23580);
and U23742 (N_23742,N_23440,N_23494);
nor U23743 (N_23743,N_23465,N_23587);
nand U23744 (N_23744,N_23427,N_23410);
nand U23745 (N_23745,N_23427,N_23544);
nand U23746 (N_23746,N_23524,N_23508);
xnor U23747 (N_23747,N_23581,N_23582);
nor U23748 (N_23748,N_23415,N_23521);
and U23749 (N_23749,N_23590,N_23492);
or U23750 (N_23750,N_23560,N_23401);
or U23751 (N_23751,N_23416,N_23409);
or U23752 (N_23752,N_23487,N_23402);
or U23753 (N_23753,N_23540,N_23466);
or U23754 (N_23754,N_23550,N_23572);
and U23755 (N_23755,N_23435,N_23551);
nand U23756 (N_23756,N_23486,N_23540);
and U23757 (N_23757,N_23437,N_23446);
nor U23758 (N_23758,N_23436,N_23528);
or U23759 (N_23759,N_23565,N_23419);
or U23760 (N_23760,N_23406,N_23491);
or U23761 (N_23761,N_23552,N_23523);
nor U23762 (N_23762,N_23471,N_23530);
nor U23763 (N_23763,N_23456,N_23400);
and U23764 (N_23764,N_23521,N_23547);
nor U23765 (N_23765,N_23416,N_23521);
nand U23766 (N_23766,N_23586,N_23512);
and U23767 (N_23767,N_23556,N_23567);
xnor U23768 (N_23768,N_23515,N_23571);
or U23769 (N_23769,N_23468,N_23571);
and U23770 (N_23770,N_23525,N_23403);
xor U23771 (N_23771,N_23463,N_23417);
xor U23772 (N_23772,N_23446,N_23401);
or U23773 (N_23773,N_23586,N_23571);
or U23774 (N_23774,N_23577,N_23422);
or U23775 (N_23775,N_23414,N_23418);
nand U23776 (N_23776,N_23428,N_23475);
or U23777 (N_23777,N_23520,N_23522);
or U23778 (N_23778,N_23473,N_23495);
and U23779 (N_23779,N_23574,N_23450);
or U23780 (N_23780,N_23422,N_23412);
or U23781 (N_23781,N_23417,N_23521);
and U23782 (N_23782,N_23563,N_23445);
nor U23783 (N_23783,N_23529,N_23555);
nand U23784 (N_23784,N_23537,N_23474);
nor U23785 (N_23785,N_23496,N_23470);
nand U23786 (N_23786,N_23596,N_23417);
and U23787 (N_23787,N_23427,N_23489);
nand U23788 (N_23788,N_23562,N_23499);
and U23789 (N_23789,N_23541,N_23442);
xnor U23790 (N_23790,N_23421,N_23552);
and U23791 (N_23791,N_23456,N_23543);
nor U23792 (N_23792,N_23454,N_23453);
nor U23793 (N_23793,N_23530,N_23540);
nand U23794 (N_23794,N_23453,N_23504);
nand U23795 (N_23795,N_23421,N_23476);
nor U23796 (N_23796,N_23451,N_23518);
nor U23797 (N_23797,N_23489,N_23584);
nor U23798 (N_23798,N_23581,N_23425);
or U23799 (N_23799,N_23414,N_23463);
nand U23800 (N_23800,N_23631,N_23684);
and U23801 (N_23801,N_23715,N_23620);
nor U23802 (N_23802,N_23651,N_23769);
nand U23803 (N_23803,N_23674,N_23604);
or U23804 (N_23804,N_23713,N_23709);
nand U23805 (N_23805,N_23721,N_23602);
nand U23806 (N_23806,N_23729,N_23704);
nor U23807 (N_23807,N_23641,N_23761);
nor U23808 (N_23808,N_23686,N_23758);
and U23809 (N_23809,N_23662,N_23740);
and U23810 (N_23810,N_23689,N_23690);
xor U23811 (N_23811,N_23666,N_23673);
or U23812 (N_23812,N_23730,N_23613);
and U23813 (N_23813,N_23731,N_23759);
nor U23814 (N_23814,N_23675,N_23617);
nor U23815 (N_23815,N_23782,N_23714);
nand U23816 (N_23816,N_23653,N_23677);
nor U23817 (N_23817,N_23647,N_23603);
nor U23818 (N_23818,N_23642,N_23752);
or U23819 (N_23819,N_23670,N_23632);
nand U23820 (N_23820,N_23744,N_23616);
xor U23821 (N_23821,N_23705,N_23696);
nor U23822 (N_23822,N_23747,N_23655);
and U23823 (N_23823,N_23716,N_23692);
and U23824 (N_23824,N_23676,N_23796);
and U23825 (N_23825,N_23718,N_23646);
or U23826 (N_23826,N_23777,N_23739);
nand U23827 (N_23827,N_23678,N_23726);
or U23828 (N_23828,N_23764,N_23753);
or U23829 (N_23829,N_23656,N_23628);
nand U23830 (N_23830,N_23717,N_23772);
nand U23831 (N_23831,N_23627,N_23630);
nor U23832 (N_23832,N_23732,N_23614);
or U23833 (N_23833,N_23600,N_23609);
xnor U23834 (N_23834,N_23738,N_23756);
nor U23835 (N_23835,N_23762,N_23601);
or U23836 (N_23836,N_23707,N_23664);
nor U23837 (N_23837,N_23697,N_23773);
or U23838 (N_23838,N_23748,N_23790);
and U23839 (N_23839,N_23785,N_23799);
nand U23840 (N_23840,N_23625,N_23734);
or U23841 (N_23841,N_23650,N_23710);
nor U23842 (N_23842,N_23755,N_23742);
xor U23843 (N_23843,N_23698,N_23669);
or U23844 (N_23844,N_23766,N_23702);
nand U23845 (N_23845,N_23671,N_23737);
nor U23846 (N_23846,N_23611,N_23683);
nand U23847 (N_23847,N_23741,N_23733);
nand U23848 (N_23848,N_23608,N_23658);
and U23849 (N_23849,N_23636,N_23645);
nor U23850 (N_23850,N_23638,N_23722);
nand U23851 (N_23851,N_23765,N_23661);
and U23852 (N_23852,N_23607,N_23667);
nor U23853 (N_23853,N_23606,N_23660);
nor U23854 (N_23854,N_23640,N_23746);
nor U23855 (N_23855,N_23712,N_23680);
nand U23856 (N_23856,N_23725,N_23685);
and U23857 (N_23857,N_23679,N_23792);
or U23858 (N_23858,N_23623,N_23688);
or U23859 (N_23859,N_23605,N_23788);
and U23860 (N_23860,N_23711,N_23724);
nand U23861 (N_23861,N_23723,N_23771);
xor U23862 (N_23862,N_23644,N_23767);
nor U23863 (N_23863,N_23778,N_23798);
xnor U23864 (N_23864,N_23615,N_23635);
or U23865 (N_23865,N_23633,N_23720);
or U23866 (N_23866,N_23701,N_23629);
or U23867 (N_23867,N_23706,N_23637);
and U23868 (N_23868,N_23797,N_23774);
nor U23869 (N_23869,N_23654,N_23657);
or U23870 (N_23870,N_23789,N_23735);
or U23871 (N_23871,N_23694,N_23776);
or U23872 (N_23872,N_23750,N_23784);
or U23873 (N_23873,N_23719,N_23708);
nor U23874 (N_23874,N_23626,N_23668);
nor U23875 (N_23875,N_23639,N_23621);
or U23876 (N_23876,N_23693,N_23682);
nor U23877 (N_23877,N_23754,N_23648);
or U23878 (N_23878,N_23699,N_23745);
nand U23879 (N_23879,N_23622,N_23787);
nand U23880 (N_23880,N_23768,N_23751);
and U23881 (N_23881,N_23780,N_23663);
nor U23882 (N_23882,N_23736,N_23760);
nor U23883 (N_23883,N_23781,N_23728);
or U23884 (N_23884,N_23791,N_23786);
nand U23885 (N_23885,N_23681,N_23610);
or U23886 (N_23886,N_23749,N_23672);
and U23887 (N_23887,N_23691,N_23763);
xnor U23888 (N_23888,N_23612,N_23783);
nor U23889 (N_23889,N_23634,N_23703);
and U23890 (N_23890,N_23779,N_23687);
or U23891 (N_23891,N_23775,N_23652);
nand U23892 (N_23892,N_23619,N_23665);
nor U23893 (N_23893,N_23770,N_23649);
nor U23894 (N_23894,N_23793,N_23700);
xnor U23895 (N_23895,N_23757,N_23659);
xor U23896 (N_23896,N_23743,N_23794);
nor U23897 (N_23897,N_23618,N_23624);
or U23898 (N_23898,N_23643,N_23795);
nor U23899 (N_23899,N_23727,N_23695);
nor U23900 (N_23900,N_23637,N_23742);
and U23901 (N_23901,N_23635,N_23634);
nor U23902 (N_23902,N_23745,N_23736);
xnor U23903 (N_23903,N_23722,N_23781);
or U23904 (N_23904,N_23682,N_23740);
and U23905 (N_23905,N_23695,N_23668);
and U23906 (N_23906,N_23613,N_23641);
and U23907 (N_23907,N_23632,N_23789);
nor U23908 (N_23908,N_23706,N_23722);
or U23909 (N_23909,N_23713,N_23701);
and U23910 (N_23910,N_23705,N_23611);
nand U23911 (N_23911,N_23791,N_23633);
or U23912 (N_23912,N_23645,N_23730);
xnor U23913 (N_23913,N_23726,N_23689);
nand U23914 (N_23914,N_23609,N_23619);
and U23915 (N_23915,N_23649,N_23709);
and U23916 (N_23916,N_23633,N_23693);
nor U23917 (N_23917,N_23733,N_23753);
nand U23918 (N_23918,N_23697,N_23612);
and U23919 (N_23919,N_23604,N_23719);
and U23920 (N_23920,N_23743,N_23656);
nor U23921 (N_23921,N_23722,N_23768);
and U23922 (N_23922,N_23753,N_23695);
or U23923 (N_23923,N_23694,N_23754);
or U23924 (N_23924,N_23721,N_23601);
nand U23925 (N_23925,N_23733,N_23634);
or U23926 (N_23926,N_23734,N_23789);
xor U23927 (N_23927,N_23670,N_23798);
nand U23928 (N_23928,N_23730,N_23777);
or U23929 (N_23929,N_23654,N_23637);
and U23930 (N_23930,N_23662,N_23778);
nand U23931 (N_23931,N_23701,N_23655);
and U23932 (N_23932,N_23653,N_23604);
nand U23933 (N_23933,N_23761,N_23618);
nand U23934 (N_23934,N_23617,N_23757);
nor U23935 (N_23935,N_23732,N_23626);
and U23936 (N_23936,N_23725,N_23664);
xor U23937 (N_23937,N_23747,N_23766);
or U23938 (N_23938,N_23797,N_23744);
nor U23939 (N_23939,N_23780,N_23793);
nor U23940 (N_23940,N_23657,N_23745);
and U23941 (N_23941,N_23776,N_23607);
or U23942 (N_23942,N_23704,N_23620);
nor U23943 (N_23943,N_23696,N_23691);
or U23944 (N_23944,N_23648,N_23738);
xnor U23945 (N_23945,N_23765,N_23735);
or U23946 (N_23946,N_23645,N_23711);
nor U23947 (N_23947,N_23607,N_23731);
and U23948 (N_23948,N_23761,N_23706);
nand U23949 (N_23949,N_23621,N_23764);
or U23950 (N_23950,N_23638,N_23647);
nand U23951 (N_23951,N_23651,N_23615);
xor U23952 (N_23952,N_23604,N_23703);
or U23953 (N_23953,N_23780,N_23654);
nand U23954 (N_23954,N_23603,N_23646);
xnor U23955 (N_23955,N_23741,N_23620);
nand U23956 (N_23956,N_23602,N_23607);
or U23957 (N_23957,N_23610,N_23713);
and U23958 (N_23958,N_23639,N_23787);
and U23959 (N_23959,N_23751,N_23679);
nor U23960 (N_23960,N_23676,N_23686);
xnor U23961 (N_23961,N_23720,N_23738);
or U23962 (N_23962,N_23629,N_23605);
nor U23963 (N_23963,N_23668,N_23667);
nand U23964 (N_23964,N_23703,N_23747);
nand U23965 (N_23965,N_23749,N_23609);
nand U23966 (N_23966,N_23672,N_23698);
and U23967 (N_23967,N_23674,N_23793);
nand U23968 (N_23968,N_23612,N_23645);
nor U23969 (N_23969,N_23669,N_23618);
xor U23970 (N_23970,N_23675,N_23701);
xnor U23971 (N_23971,N_23638,N_23754);
nor U23972 (N_23972,N_23622,N_23777);
nor U23973 (N_23973,N_23740,N_23792);
and U23974 (N_23974,N_23781,N_23616);
nand U23975 (N_23975,N_23775,N_23650);
nor U23976 (N_23976,N_23621,N_23691);
nor U23977 (N_23977,N_23641,N_23741);
nor U23978 (N_23978,N_23742,N_23667);
and U23979 (N_23979,N_23747,N_23684);
or U23980 (N_23980,N_23634,N_23623);
or U23981 (N_23981,N_23710,N_23661);
and U23982 (N_23982,N_23624,N_23626);
or U23983 (N_23983,N_23798,N_23687);
nand U23984 (N_23984,N_23796,N_23746);
or U23985 (N_23985,N_23790,N_23717);
nor U23986 (N_23986,N_23738,N_23672);
and U23987 (N_23987,N_23738,N_23778);
and U23988 (N_23988,N_23622,N_23700);
nand U23989 (N_23989,N_23775,N_23615);
xnor U23990 (N_23990,N_23684,N_23628);
nor U23991 (N_23991,N_23690,N_23668);
nor U23992 (N_23992,N_23673,N_23618);
nor U23993 (N_23993,N_23624,N_23628);
nor U23994 (N_23994,N_23632,N_23640);
and U23995 (N_23995,N_23775,N_23618);
and U23996 (N_23996,N_23665,N_23726);
nand U23997 (N_23997,N_23611,N_23749);
or U23998 (N_23998,N_23685,N_23662);
nor U23999 (N_23999,N_23633,N_23746);
and U24000 (N_24000,N_23939,N_23844);
or U24001 (N_24001,N_23807,N_23912);
nor U24002 (N_24002,N_23822,N_23969);
and U24003 (N_24003,N_23983,N_23812);
and U24004 (N_24004,N_23881,N_23940);
nand U24005 (N_24005,N_23854,N_23831);
or U24006 (N_24006,N_23941,N_23865);
xor U24007 (N_24007,N_23832,N_23900);
nor U24008 (N_24008,N_23801,N_23943);
and U24009 (N_24009,N_23907,N_23905);
nor U24010 (N_24010,N_23989,N_23921);
nor U24011 (N_24011,N_23990,N_23910);
nand U24012 (N_24012,N_23877,N_23987);
or U24013 (N_24013,N_23986,N_23984);
and U24014 (N_24014,N_23938,N_23962);
and U24015 (N_24015,N_23827,N_23849);
nor U24016 (N_24016,N_23888,N_23955);
and U24017 (N_24017,N_23897,N_23818);
nand U24018 (N_24018,N_23842,N_23851);
and U24019 (N_24019,N_23985,N_23963);
xor U24020 (N_24020,N_23883,N_23954);
nor U24021 (N_24021,N_23988,N_23874);
xnor U24022 (N_24022,N_23893,N_23889);
or U24023 (N_24023,N_23840,N_23852);
nor U24024 (N_24024,N_23913,N_23808);
xor U24025 (N_24025,N_23846,N_23861);
nand U24026 (N_24026,N_23982,N_23873);
xor U24027 (N_24027,N_23970,N_23823);
nand U24028 (N_24028,N_23876,N_23804);
xnor U24029 (N_24029,N_23820,N_23813);
and U24030 (N_24030,N_23869,N_23930);
nor U24031 (N_24031,N_23917,N_23850);
nor U24032 (N_24032,N_23980,N_23960);
or U24033 (N_24033,N_23834,N_23802);
nand U24034 (N_24034,N_23995,N_23856);
nand U24035 (N_24035,N_23973,N_23957);
nor U24036 (N_24036,N_23992,N_23862);
nor U24037 (N_24037,N_23964,N_23800);
and U24038 (N_24038,N_23872,N_23934);
or U24039 (N_24039,N_23945,N_23927);
or U24040 (N_24040,N_23965,N_23867);
nand U24041 (N_24041,N_23997,N_23841);
and U24042 (N_24042,N_23847,N_23891);
and U24043 (N_24043,N_23976,N_23811);
nor U24044 (N_24044,N_23979,N_23896);
and U24045 (N_24045,N_23809,N_23908);
and U24046 (N_24046,N_23871,N_23952);
nand U24047 (N_24047,N_23884,N_23899);
nor U24048 (N_24048,N_23879,N_23882);
nand U24049 (N_24049,N_23926,N_23966);
or U24050 (N_24050,N_23868,N_23830);
and U24051 (N_24051,N_23836,N_23931);
xor U24052 (N_24052,N_23833,N_23857);
nor U24053 (N_24053,N_23835,N_23961);
and U24054 (N_24054,N_23999,N_23914);
or U24055 (N_24055,N_23972,N_23918);
nor U24056 (N_24056,N_23919,N_23829);
or U24057 (N_24057,N_23929,N_23971);
and U24058 (N_24058,N_23991,N_23967);
and U24059 (N_24059,N_23996,N_23920);
or U24060 (N_24060,N_23895,N_23932);
nand U24061 (N_24061,N_23815,N_23859);
nand U24062 (N_24062,N_23848,N_23916);
or U24063 (N_24063,N_23816,N_23885);
and U24064 (N_24064,N_23950,N_23942);
xnor U24065 (N_24065,N_23951,N_23860);
xnor U24066 (N_24066,N_23821,N_23806);
nand U24067 (N_24067,N_23855,N_23838);
and U24068 (N_24068,N_23902,N_23948);
nand U24069 (N_24069,N_23928,N_23968);
and U24070 (N_24070,N_23892,N_23878);
or U24071 (N_24071,N_23875,N_23819);
nor U24072 (N_24072,N_23901,N_23898);
or U24073 (N_24073,N_23956,N_23894);
or U24074 (N_24074,N_23810,N_23998);
or U24075 (N_24075,N_23974,N_23946);
and U24076 (N_24076,N_23904,N_23949);
or U24077 (N_24077,N_23870,N_23977);
and U24078 (N_24078,N_23853,N_23817);
xnor U24079 (N_24079,N_23936,N_23825);
or U24080 (N_24080,N_23958,N_23906);
and U24081 (N_24081,N_23925,N_23886);
nor U24082 (N_24082,N_23922,N_23935);
and U24083 (N_24083,N_23909,N_23903);
nand U24084 (N_24084,N_23845,N_23837);
and U24085 (N_24085,N_23944,N_23824);
nand U24086 (N_24086,N_23915,N_23978);
and U24087 (N_24087,N_23828,N_23803);
or U24088 (N_24088,N_23887,N_23923);
nor U24089 (N_24089,N_23947,N_23933);
nor U24090 (N_24090,N_23866,N_23975);
and U24091 (N_24091,N_23839,N_23924);
nor U24092 (N_24092,N_23805,N_23953);
xor U24093 (N_24093,N_23814,N_23959);
and U24094 (N_24094,N_23863,N_23937);
xor U24095 (N_24095,N_23890,N_23880);
nor U24096 (N_24096,N_23981,N_23994);
nand U24097 (N_24097,N_23826,N_23858);
or U24098 (N_24098,N_23993,N_23864);
or U24099 (N_24099,N_23843,N_23911);
nand U24100 (N_24100,N_23822,N_23804);
and U24101 (N_24101,N_23820,N_23873);
and U24102 (N_24102,N_23805,N_23879);
and U24103 (N_24103,N_23892,N_23829);
nor U24104 (N_24104,N_23849,N_23968);
or U24105 (N_24105,N_23956,N_23811);
or U24106 (N_24106,N_23807,N_23892);
nand U24107 (N_24107,N_23894,N_23996);
and U24108 (N_24108,N_23870,N_23954);
and U24109 (N_24109,N_23916,N_23945);
and U24110 (N_24110,N_23891,N_23803);
or U24111 (N_24111,N_23971,N_23911);
and U24112 (N_24112,N_23939,N_23848);
nand U24113 (N_24113,N_23915,N_23882);
nor U24114 (N_24114,N_23834,N_23883);
and U24115 (N_24115,N_23849,N_23922);
nand U24116 (N_24116,N_23875,N_23843);
nor U24117 (N_24117,N_23839,N_23916);
and U24118 (N_24118,N_23963,N_23971);
nor U24119 (N_24119,N_23809,N_23962);
and U24120 (N_24120,N_23834,N_23902);
nand U24121 (N_24121,N_23873,N_23830);
nor U24122 (N_24122,N_23846,N_23802);
and U24123 (N_24123,N_23802,N_23972);
nor U24124 (N_24124,N_23849,N_23845);
nand U24125 (N_24125,N_23884,N_23953);
nand U24126 (N_24126,N_23812,N_23802);
and U24127 (N_24127,N_23944,N_23868);
nor U24128 (N_24128,N_23964,N_23878);
or U24129 (N_24129,N_23986,N_23977);
and U24130 (N_24130,N_23812,N_23973);
and U24131 (N_24131,N_23931,N_23947);
or U24132 (N_24132,N_23945,N_23868);
nor U24133 (N_24133,N_23937,N_23903);
nand U24134 (N_24134,N_23911,N_23825);
xnor U24135 (N_24135,N_23840,N_23809);
and U24136 (N_24136,N_23956,N_23814);
and U24137 (N_24137,N_23812,N_23898);
and U24138 (N_24138,N_23998,N_23912);
nor U24139 (N_24139,N_23882,N_23880);
or U24140 (N_24140,N_23807,N_23880);
or U24141 (N_24141,N_23976,N_23810);
or U24142 (N_24142,N_23978,N_23893);
and U24143 (N_24143,N_23840,N_23882);
or U24144 (N_24144,N_23884,N_23969);
and U24145 (N_24145,N_23850,N_23810);
xnor U24146 (N_24146,N_23977,N_23992);
and U24147 (N_24147,N_23850,N_23907);
and U24148 (N_24148,N_23948,N_23951);
and U24149 (N_24149,N_23861,N_23987);
nor U24150 (N_24150,N_23927,N_23991);
nor U24151 (N_24151,N_23949,N_23850);
and U24152 (N_24152,N_23930,N_23837);
nand U24153 (N_24153,N_23900,N_23838);
and U24154 (N_24154,N_23901,N_23854);
and U24155 (N_24155,N_23906,N_23872);
nand U24156 (N_24156,N_23849,N_23921);
or U24157 (N_24157,N_23877,N_23902);
and U24158 (N_24158,N_23912,N_23930);
nor U24159 (N_24159,N_23977,N_23837);
nand U24160 (N_24160,N_23981,N_23855);
nor U24161 (N_24161,N_23884,N_23902);
and U24162 (N_24162,N_23904,N_23857);
or U24163 (N_24163,N_23816,N_23800);
nor U24164 (N_24164,N_23818,N_23928);
nand U24165 (N_24165,N_23976,N_23867);
nor U24166 (N_24166,N_23844,N_23980);
or U24167 (N_24167,N_23982,N_23909);
or U24168 (N_24168,N_23897,N_23968);
or U24169 (N_24169,N_23964,N_23834);
or U24170 (N_24170,N_23829,N_23824);
nor U24171 (N_24171,N_23819,N_23860);
or U24172 (N_24172,N_23888,N_23989);
nand U24173 (N_24173,N_23871,N_23866);
nand U24174 (N_24174,N_23885,N_23979);
nor U24175 (N_24175,N_23880,N_23819);
nand U24176 (N_24176,N_23937,N_23926);
and U24177 (N_24177,N_23903,N_23892);
nor U24178 (N_24178,N_23859,N_23917);
nand U24179 (N_24179,N_23834,N_23890);
nand U24180 (N_24180,N_23924,N_23919);
nor U24181 (N_24181,N_23858,N_23844);
nor U24182 (N_24182,N_23866,N_23956);
nand U24183 (N_24183,N_23817,N_23869);
and U24184 (N_24184,N_23845,N_23994);
nand U24185 (N_24185,N_23840,N_23990);
xor U24186 (N_24186,N_23892,N_23943);
nor U24187 (N_24187,N_23800,N_23961);
xnor U24188 (N_24188,N_23849,N_23989);
or U24189 (N_24189,N_23864,N_23964);
nand U24190 (N_24190,N_23955,N_23963);
xnor U24191 (N_24191,N_23862,N_23845);
nand U24192 (N_24192,N_23875,N_23852);
or U24193 (N_24193,N_23802,N_23907);
nor U24194 (N_24194,N_23884,N_23986);
nand U24195 (N_24195,N_23985,N_23801);
nor U24196 (N_24196,N_23994,N_23967);
nand U24197 (N_24197,N_23976,N_23804);
xor U24198 (N_24198,N_23815,N_23885);
and U24199 (N_24199,N_23985,N_23915);
or U24200 (N_24200,N_24155,N_24052);
nand U24201 (N_24201,N_24139,N_24065);
nor U24202 (N_24202,N_24063,N_24059);
or U24203 (N_24203,N_24190,N_24070);
nor U24204 (N_24204,N_24008,N_24050);
and U24205 (N_24205,N_24133,N_24141);
and U24206 (N_24206,N_24157,N_24027);
nor U24207 (N_24207,N_24134,N_24098);
or U24208 (N_24208,N_24080,N_24140);
or U24209 (N_24209,N_24086,N_24111);
nand U24210 (N_24210,N_24137,N_24183);
and U24211 (N_24211,N_24069,N_24024);
nand U24212 (N_24212,N_24004,N_24022);
and U24213 (N_24213,N_24031,N_24104);
nor U24214 (N_24214,N_24192,N_24002);
and U24215 (N_24215,N_24093,N_24084);
or U24216 (N_24216,N_24081,N_24005);
or U24217 (N_24217,N_24078,N_24072);
nand U24218 (N_24218,N_24017,N_24087);
nand U24219 (N_24219,N_24107,N_24130);
nor U24220 (N_24220,N_24073,N_24125);
and U24221 (N_24221,N_24077,N_24082);
and U24222 (N_24222,N_24096,N_24193);
or U24223 (N_24223,N_24144,N_24006);
nor U24224 (N_24224,N_24102,N_24138);
xnor U24225 (N_24225,N_24172,N_24108);
nor U24226 (N_24226,N_24013,N_24101);
and U24227 (N_24227,N_24146,N_24003);
and U24228 (N_24228,N_24035,N_24051);
or U24229 (N_24229,N_24189,N_24151);
and U24230 (N_24230,N_24195,N_24043);
xor U24231 (N_24231,N_24166,N_24176);
or U24232 (N_24232,N_24023,N_24015);
and U24233 (N_24233,N_24109,N_24135);
nor U24234 (N_24234,N_24152,N_24180);
or U24235 (N_24235,N_24106,N_24030);
nor U24236 (N_24236,N_24115,N_24012);
nand U24237 (N_24237,N_24067,N_24198);
xor U24238 (N_24238,N_24041,N_24196);
nor U24239 (N_24239,N_24037,N_24154);
or U24240 (N_24240,N_24010,N_24194);
or U24241 (N_24241,N_24129,N_24150);
nand U24242 (N_24242,N_24036,N_24047);
xnor U24243 (N_24243,N_24057,N_24169);
nand U24244 (N_24244,N_24016,N_24123);
and U24245 (N_24245,N_24126,N_24145);
nand U24246 (N_24246,N_24161,N_24117);
and U24247 (N_24247,N_24042,N_24177);
nand U24248 (N_24248,N_24040,N_24097);
nand U24249 (N_24249,N_24079,N_24044);
nor U24250 (N_24250,N_24175,N_24049);
nor U24251 (N_24251,N_24018,N_24110);
or U24252 (N_24252,N_24038,N_24029);
nor U24253 (N_24253,N_24119,N_24179);
nor U24254 (N_24254,N_24120,N_24142);
nand U24255 (N_24255,N_24056,N_24088);
or U24256 (N_24256,N_24127,N_24100);
or U24257 (N_24257,N_24089,N_24091);
and U24258 (N_24258,N_24163,N_24075);
nor U24259 (N_24259,N_24185,N_24178);
nor U24260 (N_24260,N_24034,N_24020);
xor U24261 (N_24261,N_24009,N_24053);
and U24262 (N_24262,N_24164,N_24147);
nor U24263 (N_24263,N_24148,N_24054);
nor U24264 (N_24264,N_24085,N_24103);
or U24265 (N_24265,N_24039,N_24055);
and U24266 (N_24266,N_24182,N_24026);
xnor U24267 (N_24267,N_24113,N_24191);
or U24268 (N_24268,N_24092,N_24158);
nand U24269 (N_24269,N_24048,N_24045);
nor U24270 (N_24270,N_24019,N_24032);
xnor U24271 (N_24271,N_24136,N_24066);
xnor U24272 (N_24272,N_24094,N_24173);
nor U24273 (N_24273,N_24068,N_24074);
nand U24274 (N_24274,N_24011,N_24046);
or U24275 (N_24275,N_24143,N_24186);
nor U24276 (N_24276,N_24132,N_24116);
and U24277 (N_24277,N_24124,N_24099);
nand U24278 (N_24278,N_24162,N_24170);
nor U24279 (N_24279,N_24168,N_24058);
or U24280 (N_24280,N_24060,N_24064);
or U24281 (N_24281,N_24033,N_24014);
or U24282 (N_24282,N_24090,N_24105);
or U24283 (N_24283,N_24174,N_24118);
and U24284 (N_24284,N_24071,N_24028);
nand U24285 (N_24285,N_24121,N_24076);
nor U24286 (N_24286,N_24083,N_24181);
or U24287 (N_24287,N_24112,N_24153);
and U24288 (N_24288,N_24007,N_24160);
or U24289 (N_24289,N_24000,N_24095);
and U24290 (N_24290,N_24021,N_24149);
nor U24291 (N_24291,N_24159,N_24122);
nand U24292 (N_24292,N_24197,N_24199);
nor U24293 (N_24293,N_24188,N_24156);
nand U24294 (N_24294,N_24171,N_24184);
and U24295 (N_24295,N_24128,N_24165);
and U24296 (N_24296,N_24167,N_24001);
or U24297 (N_24297,N_24131,N_24025);
or U24298 (N_24298,N_24187,N_24114);
or U24299 (N_24299,N_24062,N_24061);
and U24300 (N_24300,N_24065,N_24130);
and U24301 (N_24301,N_24199,N_24021);
nor U24302 (N_24302,N_24083,N_24017);
xor U24303 (N_24303,N_24130,N_24051);
nand U24304 (N_24304,N_24161,N_24041);
nor U24305 (N_24305,N_24051,N_24049);
nand U24306 (N_24306,N_24091,N_24008);
nor U24307 (N_24307,N_24051,N_24004);
and U24308 (N_24308,N_24109,N_24141);
or U24309 (N_24309,N_24021,N_24157);
and U24310 (N_24310,N_24150,N_24186);
nor U24311 (N_24311,N_24115,N_24198);
nor U24312 (N_24312,N_24197,N_24105);
and U24313 (N_24313,N_24096,N_24081);
nand U24314 (N_24314,N_24009,N_24086);
nand U24315 (N_24315,N_24100,N_24179);
and U24316 (N_24316,N_24064,N_24078);
or U24317 (N_24317,N_24087,N_24099);
nand U24318 (N_24318,N_24141,N_24125);
xor U24319 (N_24319,N_24161,N_24018);
and U24320 (N_24320,N_24124,N_24188);
and U24321 (N_24321,N_24020,N_24102);
xnor U24322 (N_24322,N_24175,N_24082);
nor U24323 (N_24323,N_24197,N_24145);
nand U24324 (N_24324,N_24093,N_24073);
xor U24325 (N_24325,N_24136,N_24004);
nand U24326 (N_24326,N_24025,N_24173);
nand U24327 (N_24327,N_24181,N_24092);
xnor U24328 (N_24328,N_24173,N_24189);
xnor U24329 (N_24329,N_24059,N_24052);
nand U24330 (N_24330,N_24061,N_24100);
and U24331 (N_24331,N_24023,N_24039);
nand U24332 (N_24332,N_24174,N_24045);
and U24333 (N_24333,N_24091,N_24078);
or U24334 (N_24334,N_24146,N_24033);
nor U24335 (N_24335,N_24010,N_24052);
nor U24336 (N_24336,N_24171,N_24071);
or U24337 (N_24337,N_24176,N_24081);
xnor U24338 (N_24338,N_24090,N_24110);
nor U24339 (N_24339,N_24136,N_24014);
xor U24340 (N_24340,N_24178,N_24164);
nor U24341 (N_24341,N_24114,N_24185);
or U24342 (N_24342,N_24146,N_24067);
or U24343 (N_24343,N_24123,N_24080);
nor U24344 (N_24344,N_24031,N_24149);
nand U24345 (N_24345,N_24126,N_24136);
and U24346 (N_24346,N_24027,N_24142);
nand U24347 (N_24347,N_24160,N_24125);
and U24348 (N_24348,N_24122,N_24146);
xnor U24349 (N_24349,N_24175,N_24041);
and U24350 (N_24350,N_24082,N_24193);
or U24351 (N_24351,N_24108,N_24156);
nand U24352 (N_24352,N_24068,N_24122);
xnor U24353 (N_24353,N_24195,N_24125);
nand U24354 (N_24354,N_24157,N_24070);
nand U24355 (N_24355,N_24025,N_24139);
and U24356 (N_24356,N_24097,N_24061);
and U24357 (N_24357,N_24148,N_24029);
or U24358 (N_24358,N_24198,N_24142);
xor U24359 (N_24359,N_24006,N_24005);
nor U24360 (N_24360,N_24084,N_24137);
or U24361 (N_24361,N_24123,N_24084);
nand U24362 (N_24362,N_24035,N_24079);
or U24363 (N_24363,N_24179,N_24030);
and U24364 (N_24364,N_24009,N_24160);
or U24365 (N_24365,N_24180,N_24065);
nor U24366 (N_24366,N_24100,N_24105);
or U24367 (N_24367,N_24091,N_24053);
nand U24368 (N_24368,N_24040,N_24145);
and U24369 (N_24369,N_24115,N_24040);
or U24370 (N_24370,N_24005,N_24067);
or U24371 (N_24371,N_24006,N_24048);
nor U24372 (N_24372,N_24100,N_24096);
nor U24373 (N_24373,N_24114,N_24082);
and U24374 (N_24374,N_24123,N_24052);
and U24375 (N_24375,N_24010,N_24078);
or U24376 (N_24376,N_24051,N_24190);
nor U24377 (N_24377,N_24014,N_24199);
nand U24378 (N_24378,N_24010,N_24175);
nand U24379 (N_24379,N_24067,N_24019);
nand U24380 (N_24380,N_24130,N_24085);
nor U24381 (N_24381,N_24086,N_24107);
nor U24382 (N_24382,N_24167,N_24078);
and U24383 (N_24383,N_24106,N_24078);
or U24384 (N_24384,N_24116,N_24005);
nand U24385 (N_24385,N_24183,N_24142);
or U24386 (N_24386,N_24146,N_24144);
or U24387 (N_24387,N_24169,N_24114);
nor U24388 (N_24388,N_24140,N_24004);
nor U24389 (N_24389,N_24087,N_24073);
xor U24390 (N_24390,N_24115,N_24025);
or U24391 (N_24391,N_24165,N_24019);
nand U24392 (N_24392,N_24135,N_24176);
nand U24393 (N_24393,N_24123,N_24074);
nor U24394 (N_24394,N_24073,N_24058);
nand U24395 (N_24395,N_24077,N_24118);
xor U24396 (N_24396,N_24177,N_24004);
xnor U24397 (N_24397,N_24022,N_24135);
or U24398 (N_24398,N_24006,N_24070);
and U24399 (N_24399,N_24174,N_24178);
or U24400 (N_24400,N_24365,N_24362);
and U24401 (N_24401,N_24316,N_24322);
nand U24402 (N_24402,N_24346,N_24245);
nor U24403 (N_24403,N_24249,N_24260);
or U24404 (N_24404,N_24219,N_24207);
nor U24405 (N_24405,N_24339,N_24215);
xnor U24406 (N_24406,N_24330,N_24258);
nor U24407 (N_24407,N_24327,N_24369);
and U24408 (N_24408,N_24384,N_24298);
or U24409 (N_24409,N_24206,N_24284);
xnor U24410 (N_24410,N_24210,N_24268);
xor U24411 (N_24411,N_24276,N_24397);
nor U24412 (N_24412,N_24396,N_24269);
or U24413 (N_24413,N_24264,N_24263);
or U24414 (N_24414,N_24317,N_24209);
nor U24415 (N_24415,N_24234,N_24237);
and U24416 (N_24416,N_24286,N_24229);
nor U24417 (N_24417,N_24357,N_24204);
nor U24418 (N_24418,N_24377,N_24311);
nor U24419 (N_24419,N_24279,N_24341);
nor U24420 (N_24420,N_24220,N_24200);
or U24421 (N_24421,N_24364,N_24309);
nor U24422 (N_24422,N_24390,N_24315);
or U24423 (N_24423,N_24386,N_24214);
or U24424 (N_24424,N_24259,N_24270);
and U24425 (N_24425,N_24310,N_24308);
nor U24426 (N_24426,N_24300,N_24366);
nand U24427 (N_24427,N_24302,N_24367);
and U24428 (N_24428,N_24333,N_24332);
or U24429 (N_24429,N_24304,N_24319);
nor U24430 (N_24430,N_24251,N_24391);
or U24431 (N_24431,N_24278,N_24299);
or U24432 (N_24432,N_24227,N_24274);
or U24433 (N_24433,N_24208,N_24297);
or U24434 (N_24434,N_24267,N_24370);
and U24435 (N_24435,N_24340,N_24216);
nand U24436 (N_24436,N_24325,N_24290);
nor U24437 (N_24437,N_24233,N_24383);
nor U24438 (N_24438,N_24225,N_24307);
nand U24439 (N_24439,N_24349,N_24277);
and U24440 (N_24440,N_24352,N_24373);
nand U24441 (N_24441,N_24353,N_24261);
nor U24442 (N_24442,N_24372,N_24385);
xnor U24443 (N_24443,N_24241,N_24360);
and U24444 (N_24444,N_24231,N_24217);
nor U24445 (N_24445,N_24399,N_24271);
nor U24446 (N_24446,N_24288,N_24296);
xnor U24447 (N_24447,N_24238,N_24345);
and U24448 (N_24448,N_24374,N_24354);
and U24449 (N_24449,N_24376,N_24336);
and U24450 (N_24450,N_24289,N_24328);
xnor U24451 (N_24451,N_24313,N_24244);
xor U24452 (N_24452,N_24337,N_24283);
nand U24453 (N_24453,N_24203,N_24240);
and U24454 (N_24454,N_24398,N_24342);
or U24455 (N_24455,N_24343,N_24212);
nand U24456 (N_24456,N_24228,N_24235);
nor U24457 (N_24457,N_24246,N_24255);
and U24458 (N_24458,N_24201,N_24224);
and U24459 (N_24459,N_24252,N_24293);
nand U24460 (N_24460,N_24379,N_24226);
nand U24461 (N_24461,N_24223,N_24382);
nand U24462 (N_24462,N_24329,N_24254);
xnor U24463 (N_24463,N_24301,N_24221);
nand U24464 (N_24464,N_24287,N_24242);
xnor U24465 (N_24465,N_24266,N_24348);
or U24466 (N_24466,N_24292,N_24371);
nand U24467 (N_24467,N_24256,N_24232);
nor U24468 (N_24468,N_24230,N_24211);
or U24469 (N_24469,N_24368,N_24387);
or U24470 (N_24470,N_24222,N_24375);
nand U24471 (N_24471,N_24321,N_24282);
xor U24472 (N_24472,N_24247,N_24305);
nor U24473 (N_24473,N_24213,N_24388);
or U24474 (N_24474,N_24389,N_24294);
nor U24475 (N_24475,N_24306,N_24395);
and U24476 (N_24476,N_24303,N_24239);
xnor U24477 (N_24477,N_24323,N_24334);
nor U24478 (N_24478,N_24265,N_24318);
or U24479 (N_24479,N_24324,N_24262);
xnor U24480 (N_24480,N_24331,N_24359);
xnor U24481 (N_24481,N_24218,N_24326);
and U24482 (N_24482,N_24280,N_24295);
or U24483 (N_24483,N_24273,N_24312);
nand U24484 (N_24484,N_24335,N_24250);
or U24485 (N_24485,N_24363,N_24380);
or U24486 (N_24486,N_24381,N_24253);
nor U24487 (N_24487,N_24338,N_24243);
nor U24488 (N_24488,N_24285,N_24202);
and U24489 (N_24489,N_24344,N_24361);
or U24490 (N_24490,N_24356,N_24275);
and U24491 (N_24491,N_24205,N_24378);
nor U24492 (N_24492,N_24350,N_24257);
or U24493 (N_24493,N_24358,N_24291);
and U24494 (N_24494,N_24236,N_24281);
nor U24495 (N_24495,N_24347,N_24355);
and U24496 (N_24496,N_24272,N_24248);
nand U24497 (N_24497,N_24320,N_24314);
nand U24498 (N_24498,N_24351,N_24393);
nand U24499 (N_24499,N_24394,N_24392);
nor U24500 (N_24500,N_24295,N_24322);
nor U24501 (N_24501,N_24349,N_24276);
and U24502 (N_24502,N_24338,N_24213);
or U24503 (N_24503,N_24382,N_24210);
and U24504 (N_24504,N_24330,N_24261);
nand U24505 (N_24505,N_24210,N_24235);
xnor U24506 (N_24506,N_24272,N_24336);
or U24507 (N_24507,N_24224,N_24301);
and U24508 (N_24508,N_24336,N_24223);
or U24509 (N_24509,N_24299,N_24310);
nand U24510 (N_24510,N_24383,N_24275);
nand U24511 (N_24511,N_24253,N_24304);
nand U24512 (N_24512,N_24288,N_24252);
nor U24513 (N_24513,N_24264,N_24235);
xor U24514 (N_24514,N_24218,N_24205);
and U24515 (N_24515,N_24226,N_24351);
and U24516 (N_24516,N_24358,N_24348);
nand U24517 (N_24517,N_24389,N_24262);
nand U24518 (N_24518,N_24246,N_24342);
nor U24519 (N_24519,N_24376,N_24345);
and U24520 (N_24520,N_24261,N_24378);
nand U24521 (N_24521,N_24365,N_24293);
nor U24522 (N_24522,N_24298,N_24244);
and U24523 (N_24523,N_24237,N_24371);
nor U24524 (N_24524,N_24297,N_24345);
xnor U24525 (N_24525,N_24212,N_24316);
nand U24526 (N_24526,N_24397,N_24320);
and U24527 (N_24527,N_24309,N_24262);
xnor U24528 (N_24528,N_24223,N_24237);
or U24529 (N_24529,N_24310,N_24372);
and U24530 (N_24530,N_24201,N_24358);
nor U24531 (N_24531,N_24382,N_24350);
nor U24532 (N_24532,N_24220,N_24289);
or U24533 (N_24533,N_24278,N_24367);
xor U24534 (N_24534,N_24378,N_24326);
nand U24535 (N_24535,N_24389,N_24248);
nand U24536 (N_24536,N_24270,N_24266);
nor U24537 (N_24537,N_24396,N_24300);
nand U24538 (N_24538,N_24369,N_24379);
and U24539 (N_24539,N_24277,N_24312);
nor U24540 (N_24540,N_24273,N_24231);
and U24541 (N_24541,N_24374,N_24236);
nand U24542 (N_24542,N_24233,N_24335);
and U24543 (N_24543,N_24281,N_24270);
xor U24544 (N_24544,N_24389,N_24361);
nand U24545 (N_24545,N_24312,N_24391);
nor U24546 (N_24546,N_24276,N_24300);
xor U24547 (N_24547,N_24298,N_24320);
and U24548 (N_24548,N_24322,N_24378);
nor U24549 (N_24549,N_24312,N_24289);
nand U24550 (N_24550,N_24296,N_24333);
nand U24551 (N_24551,N_24213,N_24257);
xor U24552 (N_24552,N_24319,N_24211);
nand U24553 (N_24553,N_24223,N_24381);
xor U24554 (N_24554,N_24368,N_24315);
or U24555 (N_24555,N_24395,N_24228);
or U24556 (N_24556,N_24352,N_24299);
nor U24557 (N_24557,N_24296,N_24378);
or U24558 (N_24558,N_24305,N_24368);
and U24559 (N_24559,N_24229,N_24263);
nand U24560 (N_24560,N_24270,N_24277);
nor U24561 (N_24561,N_24205,N_24227);
and U24562 (N_24562,N_24302,N_24368);
nand U24563 (N_24563,N_24319,N_24325);
nor U24564 (N_24564,N_24220,N_24216);
xor U24565 (N_24565,N_24342,N_24399);
nor U24566 (N_24566,N_24222,N_24256);
or U24567 (N_24567,N_24345,N_24344);
nand U24568 (N_24568,N_24234,N_24236);
nand U24569 (N_24569,N_24227,N_24329);
nor U24570 (N_24570,N_24303,N_24202);
nor U24571 (N_24571,N_24234,N_24344);
nor U24572 (N_24572,N_24398,N_24318);
or U24573 (N_24573,N_24374,N_24232);
nor U24574 (N_24574,N_24224,N_24229);
and U24575 (N_24575,N_24203,N_24267);
nor U24576 (N_24576,N_24334,N_24273);
and U24577 (N_24577,N_24377,N_24200);
and U24578 (N_24578,N_24291,N_24258);
and U24579 (N_24579,N_24327,N_24212);
nand U24580 (N_24580,N_24384,N_24378);
or U24581 (N_24581,N_24208,N_24267);
xnor U24582 (N_24582,N_24256,N_24285);
xnor U24583 (N_24583,N_24233,N_24227);
or U24584 (N_24584,N_24235,N_24320);
and U24585 (N_24585,N_24215,N_24208);
nand U24586 (N_24586,N_24385,N_24345);
nand U24587 (N_24587,N_24230,N_24310);
nor U24588 (N_24588,N_24310,N_24399);
or U24589 (N_24589,N_24243,N_24218);
and U24590 (N_24590,N_24268,N_24290);
xnor U24591 (N_24591,N_24354,N_24304);
nor U24592 (N_24592,N_24310,N_24315);
and U24593 (N_24593,N_24349,N_24233);
xor U24594 (N_24594,N_24243,N_24380);
nor U24595 (N_24595,N_24360,N_24271);
nor U24596 (N_24596,N_24200,N_24356);
nand U24597 (N_24597,N_24327,N_24257);
and U24598 (N_24598,N_24392,N_24367);
nand U24599 (N_24599,N_24331,N_24360);
or U24600 (N_24600,N_24452,N_24520);
nand U24601 (N_24601,N_24597,N_24523);
or U24602 (N_24602,N_24504,N_24587);
and U24603 (N_24603,N_24422,N_24434);
nand U24604 (N_24604,N_24525,N_24496);
nor U24605 (N_24605,N_24599,N_24448);
xnor U24606 (N_24606,N_24487,N_24494);
xnor U24607 (N_24607,N_24536,N_24440);
or U24608 (N_24608,N_24539,N_24438);
nor U24609 (N_24609,N_24591,N_24421);
or U24610 (N_24610,N_24436,N_24509);
nand U24611 (N_24611,N_24480,N_24537);
nand U24612 (N_24612,N_24511,N_24561);
and U24613 (N_24613,N_24566,N_24428);
nor U24614 (N_24614,N_24588,N_24555);
nand U24615 (N_24615,N_24470,N_24472);
and U24616 (N_24616,N_24559,N_24481);
xnor U24617 (N_24617,N_24571,N_24489);
and U24618 (N_24618,N_24426,N_24420);
xnor U24619 (N_24619,N_24402,N_24579);
or U24620 (N_24620,N_24431,N_24497);
or U24621 (N_24621,N_24593,N_24408);
nand U24622 (N_24622,N_24486,N_24545);
nor U24623 (N_24623,N_24595,N_24473);
or U24624 (N_24624,N_24488,N_24590);
nand U24625 (N_24625,N_24584,N_24517);
or U24626 (N_24626,N_24544,N_24450);
nand U24627 (N_24627,N_24449,N_24560);
and U24628 (N_24628,N_24543,N_24585);
nand U24629 (N_24629,N_24457,N_24530);
or U24630 (N_24630,N_24503,N_24581);
nor U24631 (N_24631,N_24534,N_24578);
or U24632 (N_24632,N_24549,N_24557);
or U24633 (N_24633,N_24541,N_24437);
nand U24634 (N_24634,N_24563,N_24477);
nand U24635 (N_24635,N_24576,N_24479);
nand U24636 (N_24636,N_24492,N_24458);
nor U24637 (N_24637,N_24466,N_24499);
xnor U24638 (N_24638,N_24594,N_24418);
nand U24639 (N_24639,N_24569,N_24455);
xnor U24640 (N_24640,N_24592,N_24506);
nor U24641 (N_24641,N_24582,N_24412);
or U24642 (N_24642,N_24409,N_24467);
nand U24643 (N_24643,N_24567,N_24427);
or U24644 (N_24644,N_24589,N_24586);
or U24645 (N_24645,N_24540,N_24446);
nand U24646 (N_24646,N_24469,N_24514);
and U24647 (N_24647,N_24460,N_24495);
nand U24648 (N_24648,N_24414,N_24462);
xor U24649 (N_24649,N_24573,N_24505);
and U24650 (N_24650,N_24538,N_24507);
nor U24651 (N_24651,N_24528,N_24454);
and U24652 (N_24652,N_24419,N_24413);
nor U24653 (N_24653,N_24456,N_24501);
and U24654 (N_24654,N_24407,N_24429);
and U24655 (N_24655,N_24512,N_24531);
and U24656 (N_24656,N_24404,N_24475);
nand U24657 (N_24657,N_24476,N_24403);
or U24658 (N_24658,N_24568,N_24513);
and U24659 (N_24659,N_24529,N_24551);
nand U24660 (N_24660,N_24583,N_24405);
xor U24661 (N_24661,N_24527,N_24498);
or U24662 (N_24662,N_24532,N_24482);
nor U24663 (N_24663,N_24424,N_24401);
nand U24664 (N_24664,N_24553,N_24464);
nand U24665 (N_24665,N_24432,N_24400);
nor U24666 (N_24666,N_24548,N_24411);
and U24667 (N_24667,N_24441,N_24562);
nor U24668 (N_24668,N_24552,N_24515);
or U24669 (N_24669,N_24522,N_24471);
and U24670 (N_24670,N_24516,N_24575);
or U24671 (N_24671,N_24564,N_24519);
nand U24672 (N_24672,N_24474,N_24459);
or U24673 (N_24673,N_24478,N_24433);
and U24674 (N_24674,N_24439,N_24500);
or U24675 (N_24675,N_24447,N_24485);
nand U24676 (N_24676,N_24542,N_24574);
nand U24677 (N_24677,N_24577,N_24435);
or U24678 (N_24678,N_24468,N_24453);
and U24679 (N_24679,N_24535,N_24554);
nor U24680 (N_24680,N_24445,N_24415);
nand U24681 (N_24681,N_24558,N_24491);
nor U24682 (N_24682,N_24461,N_24490);
xnor U24683 (N_24683,N_24580,N_24526);
nor U24684 (N_24684,N_24484,N_24533);
nor U24685 (N_24685,N_24596,N_24546);
nor U24686 (N_24686,N_24416,N_24570);
nand U24687 (N_24687,N_24550,N_24443);
and U24688 (N_24688,N_24423,N_24442);
and U24689 (N_24689,N_24463,N_24565);
or U24690 (N_24690,N_24410,N_24425);
or U24691 (N_24691,N_24572,N_24547);
and U24692 (N_24692,N_24510,N_24502);
or U24693 (N_24693,N_24444,N_24524);
nand U24694 (N_24694,N_24518,N_24451);
nand U24695 (N_24695,N_24406,N_24556);
or U24696 (N_24696,N_24521,N_24483);
and U24697 (N_24697,N_24598,N_24417);
and U24698 (N_24698,N_24508,N_24430);
nor U24699 (N_24699,N_24493,N_24465);
or U24700 (N_24700,N_24520,N_24465);
nor U24701 (N_24701,N_24517,N_24486);
nor U24702 (N_24702,N_24474,N_24569);
and U24703 (N_24703,N_24462,N_24545);
and U24704 (N_24704,N_24472,N_24549);
nor U24705 (N_24705,N_24528,N_24550);
or U24706 (N_24706,N_24521,N_24569);
or U24707 (N_24707,N_24462,N_24485);
and U24708 (N_24708,N_24492,N_24432);
xor U24709 (N_24709,N_24426,N_24506);
nor U24710 (N_24710,N_24584,N_24598);
xnor U24711 (N_24711,N_24470,N_24486);
nand U24712 (N_24712,N_24496,N_24576);
and U24713 (N_24713,N_24557,N_24470);
nor U24714 (N_24714,N_24528,N_24428);
nor U24715 (N_24715,N_24481,N_24460);
and U24716 (N_24716,N_24545,N_24470);
and U24717 (N_24717,N_24565,N_24595);
nor U24718 (N_24718,N_24546,N_24441);
nor U24719 (N_24719,N_24433,N_24414);
nand U24720 (N_24720,N_24451,N_24506);
xor U24721 (N_24721,N_24537,N_24473);
nand U24722 (N_24722,N_24507,N_24599);
nand U24723 (N_24723,N_24517,N_24467);
nor U24724 (N_24724,N_24467,N_24429);
or U24725 (N_24725,N_24523,N_24430);
nand U24726 (N_24726,N_24505,N_24565);
or U24727 (N_24727,N_24585,N_24561);
and U24728 (N_24728,N_24581,N_24418);
nand U24729 (N_24729,N_24401,N_24558);
nand U24730 (N_24730,N_24512,N_24597);
nor U24731 (N_24731,N_24457,N_24543);
nand U24732 (N_24732,N_24542,N_24548);
and U24733 (N_24733,N_24469,N_24516);
or U24734 (N_24734,N_24514,N_24425);
xnor U24735 (N_24735,N_24410,N_24582);
nand U24736 (N_24736,N_24412,N_24592);
and U24737 (N_24737,N_24451,N_24497);
or U24738 (N_24738,N_24422,N_24421);
or U24739 (N_24739,N_24484,N_24458);
or U24740 (N_24740,N_24483,N_24416);
and U24741 (N_24741,N_24412,N_24407);
nand U24742 (N_24742,N_24427,N_24437);
nor U24743 (N_24743,N_24409,N_24482);
and U24744 (N_24744,N_24526,N_24571);
or U24745 (N_24745,N_24582,N_24544);
or U24746 (N_24746,N_24437,N_24441);
and U24747 (N_24747,N_24425,N_24566);
nor U24748 (N_24748,N_24437,N_24408);
xor U24749 (N_24749,N_24468,N_24429);
nand U24750 (N_24750,N_24402,N_24590);
nand U24751 (N_24751,N_24422,N_24488);
or U24752 (N_24752,N_24407,N_24446);
and U24753 (N_24753,N_24524,N_24434);
and U24754 (N_24754,N_24573,N_24565);
nand U24755 (N_24755,N_24517,N_24478);
nor U24756 (N_24756,N_24535,N_24539);
nor U24757 (N_24757,N_24528,N_24437);
nor U24758 (N_24758,N_24497,N_24560);
or U24759 (N_24759,N_24479,N_24476);
nor U24760 (N_24760,N_24439,N_24546);
nor U24761 (N_24761,N_24549,N_24583);
nor U24762 (N_24762,N_24402,N_24512);
nand U24763 (N_24763,N_24478,N_24570);
nor U24764 (N_24764,N_24544,N_24430);
and U24765 (N_24765,N_24555,N_24502);
or U24766 (N_24766,N_24540,N_24596);
nand U24767 (N_24767,N_24584,N_24523);
and U24768 (N_24768,N_24537,N_24527);
nand U24769 (N_24769,N_24444,N_24501);
or U24770 (N_24770,N_24471,N_24505);
nor U24771 (N_24771,N_24486,N_24583);
nand U24772 (N_24772,N_24452,N_24412);
nand U24773 (N_24773,N_24418,N_24442);
and U24774 (N_24774,N_24415,N_24569);
nor U24775 (N_24775,N_24447,N_24527);
or U24776 (N_24776,N_24497,N_24522);
nand U24777 (N_24777,N_24530,N_24407);
and U24778 (N_24778,N_24599,N_24500);
nor U24779 (N_24779,N_24420,N_24452);
nor U24780 (N_24780,N_24417,N_24503);
nor U24781 (N_24781,N_24575,N_24465);
nor U24782 (N_24782,N_24465,N_24510);
or U24783 (N_24783,N_24581,N_24494);
nand U24784 (N_24784,N_24567,N_24524);
nor U24785 (N_24785,N_24478,N_24465);
or U24786 (N_24786,N_24420,N_24559);
or U24787 (N_24787,N_24476,N_24426);
or U24788 (N_24788,N_24474,N_24573);
xnor U24789 (N_24789,N_24475,N_24428);
or U24790 (N_24790,N_24450,N_24535);
nor U24791 (N_24791,N_24526,N_24473);
nand U24792 (N_24792,N_24425,N_24549);
nor U24793 (N_24793,N_24491,N_24571);
nand U24794 (N_24794,N_24495,N_24400);
xnor U24795 (N_24795,N_24513,N_24594);
and U24796 (N_24796,N_24583,N_24422);
or U24797 (N_24797,N_24479,N_24449);
nand U24798 (N_24798,N_24523,N_24543);
or U24799 (N_24799,N_24505,N_24402);
nand U24800 (N_24800,N_24733,N_24681);
and U24801 (N_24801,N_24743,N_24729);
and U24802 (N_24802,N_24708,N_24712);
xor U24803 (N_24803,N_24638,N_24784);
xnor U24804 (N_24804,N_24780,N_24782);
nand U24805 (N_24805,N_24707,N_24693);
nor U24806 (N_24806,N_24793,N_24674);
nor U24807 (N_24807,N_24767,N_24749);
and U24808 (N_24808,N_24702,N_24673);
nor U24809 (N_24809,N_24646,N_24652);
nor U24810 (N_24810,N_24713,N_24601);
and U24811 (N_24811,N_24742,N_24647);
and U24812 (N_24812,N_24658,N_24687);
or U24813 (N_24813,N_24755,N_24617);
nand U24814 (N_24814,N_24694,N_24703);
nor U24815 (N_24815,N_24626,N_24683);
nor U24816 (N_24816,N_24611,N_24657);
or U24817 (N_24817,N_24671,N_24636);
nor U24818 (N_24818,N_24668,N_24631);
and U24819 (N_24819,N_24774,N_24635);
and U24820 (N_24820,N_24685,N_24698);
nor U24821 (N_24821,N_24630,N_24692);
nor U24822 (N_24822,N_24754,N_24672);
nand U24823 (N_24823,N_24699,N_24794);
xnor U24824 (N_24824,N_24763,N_24637);
or U24825 (N_24825,N_24797,N_24644);
nand U24826 (N_24826,N_24704,N_24615);
nand U24827 (N_24827,N_24609,N_24696);
nor U24828 (N_24828,N_24798,N_24779);
nor U24829 (N_24829,N_24776,N_24641);
or U24830 (N_24830,N_24608,N_24614);
nand U24831 (N_24831,N_24628,N_24706);
xor U24832 (N_24832,N_24639,N_24732);
nor U24833 (N_24833,N_24781,N_24736);
or U24834 (N_24834,N_24783,N_24610);
nand U24835 (N_24835,N_24669,N_24649);
nor U24836 (N_24836,N_24758,N_24747);
nand U24837 (N_24837,N_24745,N_24719);
and U24838 (N_24838,N_24680,N_24709);
or U24839 (N_24839,N_24607,N_24790);
and U24840 (N_24840,N_24632,N_24714);
or U24841 (N_24841,N_24697,N_24622);
and U24842 (N_24842,N_24720,N_24788);
and U24843 (N_24843,N_24748,N_24640);
nor U24844 (N_24844,N_24651,N_24665);
nor U24845 (N_24845,N_24752,N_24744);
or U24846 (N_24846,N_24756,N_24751);
xnor U24847 (N_24847,N_24603,N_24686);
nand U24848 (N_24848,N_24765,N_24656);
or U24849 (N_24849,N_24710,N_24761);
or U24850 (N_24850,N_24791,N_24633);
and U24851 (N_24851,N_24730,N_24722);
nor U24852 (N_24852,N_24796,N_24773);
and U24853 (N_24853,N_24660,N_24724);
and U24854 (N_24854,N_24735,N_24664);
or U24855 (N_24855,N_24634,N_24663);
or U24856 (N_24856,N_24625,N_24750);
nor U24857 (N_24857,N_24726,N_24764);
or U24858 (N_24858,N_24792,N_24734);
nand U24859 (N_24859,N_24604,N_24716);
or U24860 (N_24860,N_24740,N_24760);
or U24861 (N_24861,N_24653,N_24619);
and U24862 (N_24862,N_24645,N_24688);
and U24863 (N_24863,N_24701,N_24769);
nor U24864 (N_24864,N_24731,N_24621);
and U24865 (N_24865,N_24772,N_24602);
and U24866 (N_24866,N_24741,N_24777);
xor U24867 (N_24867,N_24655,N_24670);
nand U24868 (N_24868,N_24725,N_24661);
and U24869 (N_24869,N_24623,N_24715);
nor U24870 (N_24870,N_24606,N_24762);
xor U24871 (N_24871,N_24667,N_24675);
and U24872 (N_24872,N_24717,N_24659);
nand U24873 (N_24873,N_24795,N_24705);
and U24874 (N_24874,N_24746,N_24739);
nor U24875 (N_24875,N_24700,N_24648);
nor U24876 (N_24876,N_24654,N_24786);
nor U24877 (N_24877,N_24771,N_24662);
nor U24878 (N_24878,N_24738,N_24616);
and U24879 (N_24879,N_24690,N_24605);
or U24880 (N_24880,N_24775,N_24676);
xor U24881 (N_24881,N_24770,N_24627);
and U24882 (N_24882,N_24768,N_24689);
and U24883 (N_24883,N_24643,N_24718);
or U24884 (N_24884,N_24613,N_24789);
nand U24885 (N_24885,N_24721,N_24759);
or U24886 (N_24886,N_24642,N_24753);
or U24887 (N_24887,N_24629,N_24620);
nand U24888 (N_24888,N_24737,N_24679);
nand U24889 (N_24889,N_24682,N_24691);
or U24890 (N_24890,N_24624,N_24666);
or U24891 (N_24891,N_24684,N_24695);
or U24892 (N_24892,N_24757,N_24723);
nand U24893 (N_24893,N_24678,N_24799);
or U24894 (N_24894,N_24711,N_24618);
and U24895 (N_24895,N_24766,N_24677);
and U24896 (N_24896,N_24778,N_24650);
nor U24897 (N_24897,N_24600,N_24728);
and U24898 (N_24898,N_24727,N_24612);
or U24899 (N_24899,N_24785,N_24787);
or U24900 (N_24900,N_24689,N_24601);
nor U24901 (N_24901,N_24608,N_24718);
xor U24902 (N_24902,N_24761,N_24768);
nand U24903 (N_24903,N_24725,N_24683);
nand U24904 (N_24904,N_24670,N_24779);
and U24905 (N_24905,N_24751,N_24645);
nor U24906 (N_24906,N_24713,N_24799);
or U24907 (N_24907,N_24716,N_24705);
nor U24908 (N_24908,N_24770,N_24680);
or U24909 (N_24909,N_24610,N_24665);
and U24910 (N_24910,N_24771,N_24610);
nor U24911 (N_24911,N_24707,N_24625);
xor U24912 (N_24912,N_24659,N_24751);
nor U24913 (N_24913,N_24626,N_24696);
or U24914 (N_24914,N_24797,N_24791);
nand U24915 (N_24915,N_24698,N_24657);
or U24916 (N_24916,N_24730,N_24645);
nand U24917 (N_24917,N_24635,N_24664);
nand U24918 (N_24918,N_24743,N_24648);
or U24919 (N_24919,N_24766,N_24723);
and U24920 (N_24920,N_24783,N_24647);
nand U24921 (N_24921,N_24778,N_24630);
or U24922 (N_24922,N_24603,N_24664);
nand U24923 (N_24923,N_24683,N_24716);
and U24924 (N_24924,N_24646,N_24775);
and U24925 (N_24925,N_24707,N_24757);
and U24926 (N_24926,N_24713,N_24779);
or U24927 (N_24927,N_24648,N_24605);
nand U24928 (N_24928,N_24652,N_24729);
and U24929 (N_24929,N_24708,N_24646);
or U24930 (N_24930,N_24767,N_24678);
nand U24931 (N_24931,N_24713,N_24664);
nand U24932 (N_24932,N_24656,N_24604);
or U24933 (N_24933,N_24610,N_24689);
nand U24934 (N_24934,N_24758,N_24643);
and U24935 (N_24935,N_24685,N_24602);
nand U24936 (N_24936,N_24623,N_24738);
or U24937 (N_24937,N_24798,N_24781);
and U24938 (N_24938,N_24678,N_24715);
xnor U24939 (N_24939,N_24643,N_24607);
and U24940 (N_24940,N_24757,N_24724);
nor U24941 (N_24941,N_24623,N_24700);
nand U24942 (N_24942,N_24723,N_24636);
nor U24943 (N_24943,N_24602,N_24601);
nor U24944 (N_24944,N_24617,N_24609);
nand U24945 (N_24945,N_24787,N_24644);
nor U24946 (N_24946,N_24602,N_24668);
nand U24947 (N_24947,N_24757,N_24685);
and U24948 (N_24948,N_24689,N_24770);
nand U24949 (N_24949,N_24798,N_24645);
or U24950 (N_24950,N_24601,N_24691);
nand U24951 (N_24951,N_24600,N_24691);
xnor U24952 (N_24952,N_24612,N_24709);
nor U24953 (N_24953,N_24799,N_24607);
and U24954 (N_24954,N_24686,N_24743);
or U24955 (N_24955,N_24797,N_24630);
nand U24956 (N_24956,N_24789,N_24643);
or U24957 (N_24957,N_24657,N_24655);
or U24958 (N_24958,N_24795,N_24644);
nand U24959 (N_24959,N_24654,N_24728);
or U24960 (N_24960,N_24761,N_24735);
nor U24961 (N_24961,N_24721,N_24753);
or U24962 (N_24962,N_24716,N_24798);
and U24963 (N_24963,N_24706,N_24659);
or U24964 (N_24964,N_24696,N_24724);
nor U24965 (N_24965,N_24693,N_24724);
nor U24966 (N_24966,N_24786,N_24788);
nor U24967 (N_24967,N_24652,N_24669);
or U24968 (N_24968,N_24781,N_24797);
nand U24969 (N_24969,N_24697,N_24645);
nor U24970 (N_24970,N_24729,N_24649);
or U24971 (N_24971,N_24647,N_24673);
and U24972 (N_24972,N_24759,N_24628);
or U24973 (N_24973,N_24764,N_24714);
nand U24974 (N_24974,N_24626,N_24790);
or U24975 (N_24975,N_24635,N_24706);
and U24976 (N_24976,N_24747,N_24741);
and U24977 (N_24977,N_24632,N_24617);
nand U24978 (N_24978,N_24657,N_24769);
and U24979 (N_24979,N_24758,N_24689);
and U24980 (N_24980,N_24629,N_24639);
nor U24981 (N_24981,N_24716,N_24647);
or U24982 (N_24982,N_24728,N_24739);
xor U24983 (N_24983,N_24622,N_24793);
or U24984 (N_24984,N_24682,N_24749);
and U24985 (N_24985,N_24699,N_24635);
nor U24986 (N_24986,N_24627,N_24743);
or U24987 (N_24987,N_24635,N_24721);
nand U24988 (N_24988,N_24662,N_24688);
xor U24989 (N_24989,N_24798,N_24662);
and U24990 (N_24990,N_24692,N_24742);
xnor U24991 (N_24991,N_24778,N_24643);
nand U24992 (N_24992,N_24714,N_24611);
or U24993 (N_24993,N_24663,N_24702);
nand U24994 (N_24994,N_24616,N_24635);
nor U24995 (N_24995,N_24726,N_24750);
or U24996 (N_24996,N_24617,N_24691);
nor U24997 (N_24997,N_24663,N_24678);
xor U24998 (N_24998,N_24602,N_24748);
or U24999 (N_24999,N_24606,N_24619);
nand UO_0 (O_0,N_24857,N_24940);
or UO_1 (O_1,N_24835,N_24921);
or UO_2 (O_2,N_24991,N_24825);
and UO_3 (O_3,N_24826,N_24862);
nand UO_4 (O_4,N_24845,N_24929);
nand UO_5 (O_5,N_24902,N_24830);
nor UO_6 (O_6,N_24985,N_24922);
xor UO_7 (O_7,N_24873,N_24858);
nor UO_8 (O_8,N_24927,N_24980);
or UO_9 (O_9,N_24861,N_24990);
nand UO_10 (O_10,N_24901,N_24923);
or UO_11 (O_11,N_24920,N_24821);
or UO_12 (O_12,N_24935,N_24957);
nand UO_13 (O_13,N_24892,N_24854);
nand UO_14 (O_14,N_24905,N_24952);
xnor UO_15 (O_15,N_24885,N_24950);
or UO_16 (O_16,N_24938,N_24973);
or UO_17 (O_17,N_24919,N_24823);
nand UO_18 (O_18,N_24876,N_24846);
xnor UO_19 (O_19,N_24908,N_24998);
nor UO_20 (O_20,N_24891,N_24877);
or UO_21 (O_21,N_24833,N_24910);
nand UO_22 (O_22,N_24997,N_24931);
nand UO_23 (O_23,N_24936,N_24996);
nor UO_24 (O_24,N_24983,N_24893);
or UO_25 (O_25,N_24993,N_24813);
nand UO_26 (O_26,N_24971,N_24800);
or UO_27 (O_27,N_24970,N_24817);
or UO_28 (O_28,N_24956,N_24868);
nor UO_29 (O_29,N_24987,N_24949);
nand UO_30 (O_30,N_24803,N_24900);
nand UO_31 (O_31,N_24838,N_24889);
nor UO_32 (O_32,N_24874,N_24865);
nor UO_33 (O_33,N_24934,N_24839);
nand UO_34 (O_34,N_24962,N_24969);
and UO_35 (O_35,N_24866,N_24974);
or UO_36 (O_36,N_24943,N_24979);
nand UO_37 (O_37,N_24831,N_24939);
nand UO_38 (O_38,N_24975,N_24872);
nand UO_39 (O_39,N_24942,N_24882);
nand UO_40 (O_40,N_24994,N_24802);
or UO_41 (O_41,N_24828,N_24977);
nand UO_42 (O_42,N_24945,N_24960);
or UO_43 (O_43,N_24853,N_24859);
or UO_44 (O_44,N_24961,N_24941);
and UO_45 (O_45,N_24804,N_24888);
or UO_46 (O_46,N_24811,N_24847);
nand UO_47 (O_47,N_24903,N_24818);
nand UO_48 (O_48,N_24808,N_24850);
and UO_49 (O_49,N_24896,N_24815);
or UO_50 (O_50,N_24932,N_24926);
nor UO_51 (O_51,N_24937,N_24879);
nor UO_52 (O_52,N_24863,N_24984);
or UO_53 (O_53,N_24899,N_24871);
nand UO_54 (O_54,N_24955,N_24959);
nand UO_55 (O_55,N_24914,N_24992);
or UO_56 (O_56,N_24898,N_24849);
xor UO_57 (O_57,N_24807,N_24965);
and UO_58 (O_58,N_24933,N_24805);
nor UO_59 (O_59,N_24886,N_24967);
and UO_60 (O_60,N_24834,N_24887);
nand UO_61 (O_61,N_24806,N_24814);
nand UO_62 (O_62,N_24946,N_24809);
or UO_63 (O_63,N_24958,N_24912);
nor UO_64 (O_64,N_24966,N_24963);
nor UO_65 (O_65,N_24995,N_24913);
or UO_66 (O_66,N_24829,N_24856);
xnor UO_67 (O_67,N_24982,N_24988);
or UO_68 (O_68,N_24953,N_24822);
and UO_69 (O_69,N_24827,N_24848);
xnor UO_70 (O_70,N_24832,N_24841);
or UO_71 (O_71,N_24916,N_24928);
nand UO_72 (O_72,N_24864,N_24890);
nand UO_73 (O_73,N_24884,N_24816);
nand UO_74 (O_74,N_24948,N_24918);
xnor UO_75 (O_75,N_24843,N_24925);
xor UO_76 (O_76,N_24924,N_24819);
nor UO_77 (O_77,N_24875,N_24867);
and UO_78 (O_78,N_24836,N_24909);
or UO_79 (O_79,N_24860,N_24812);
or UO_80 (O_80,N_24981,N_24907);
nor UO_81 (O_81,N_24930,N_24954);
nor UO_82 (O_82,N_24911,N_24894);
or UO_83 (O_83,N_24904,N_24917);
nand UO_84 (O_84,N_24989,N_24976);
nor UO_85 (O_85,N_24820,N_24999);
nor UO_86 (O_86,N_24951,N_24944);
or UO_87 (O_87,N_24801,N_24842);
xnor UO_88 (O_88,N_24840,N_24968);
or UO_89 (O_89,N_24986,N_24915);
or UO_90 (O_90,N_24947,N_24824);
nand UO_91 (O_91,N_24881,N_24906);
and UO_92 (O_92,N_24810,N_24855);
nand UO_93 (O_93,N_24880,N_24978);
nand UO_94 (O_94,N_24878,N_24852);
and UO_95 (O_95,N_24870,N_24883);
xnor UO_96 (O_96,N_24964,N_24897);
xor UO_97 (O_97,N_24844,N_24972);
nor UO_98 (O_98,N_24895,N_24837);
nand UO_99 (O_99,N_24869,N_24851);
xnor UO_100 (O_100,N_24808,N_24887);
nor UO_101 (O_101,N_24981,N_24994);
nand UO_102 (O_102,N_24962,N_24964);
or UO_103 (O_103,N_24995,N_24908);
or UO_104 (O_104,N_24906,N_24926);
and UO_105 (O_105,N_24837,N_24816);
nor UO_106 (O_106,N_24961,N_24837);
xor UO_107 (O_107,N_24851,N_24954);
nand UO_108 (O_108,N_24876,N_24815);
nor UO_109 (O_109,N_24961,N_24926);
and UO_110 (O_110,N_24953,N_24865);
and UO_111 (O_111,N_24913,N_24912);
xor UO_112 (O_112,N_24895,N_24936);
nor UO_113 (O_113,N_24988,N_24864);
or UO_114 (O_114,N_24803,N_24996);
nand UO_115 (O_115,N_24993,N_24815);
xnor UO_116 (O_116,N_24871,N_24996);
or UO_117 (O_117,N_24864,N_24957);
xnor UO_118 (O_118,N_24894,N_24954);
nand UO_119 (O_119,N_24812,N_24867);
nand UO_120 (O_120,N_24959,N_24899);
and UO_121 (O_121,N_24966,N_24973);
or UO_122 (O_122,N_24817,N_24837);
or UO_123 (O_123,N_24926,N_24918);
nand UO_124 (O_124,N_24868,N_24840);
or UO_125 (O_125,N_24906,N_24876);
nor UO_126 (O_126,N_24902,N_24967);
nor UO_127 (O_127,N_24850,N_24991);
nand UO_128 (O_128,N_24977,N_24923);
nand UO_129 (O_129,N_24954,N_24899);
xor UO_130 (O_130,N_24936,N_24864);
nand UO_131 (O_131,N_24999,N_24943);
or UO_132 (O_132,N_24971,N_24833);
and UO_133 (O_133,N_24809,N_24801);
or UO_134 (O_134,N_24873,N_24826);
or UO_135 (O_135,N_24985,N_24855);
nor UO_136 (O_136,N_24858,N_24863);
xnor UO_137 (O_137,N_24938,N_24801);
and UO_138 (O_138,N_24822,N_24915);
or UO_139 (O_139,N_24921,N_24829);
nand UO_140 (O_140,N_24930,N_24810);
nor UO_141 (O_141,N_24881,N_24891);
or UO_142 (O_142,N_24901,N_24914);
nand UO_143 (O_143,N_24993,N_24940);
xnor UO_144 (O_144,N_24998,N_24900);
or UO_145 (O_145,N_24930,N_24922);
nand UO_146 (O_146,N_24830,N_24951);
and UO_147 (O_147,N_24894,N_24937);
nand UO_148 (O_148,N_24986,N_24848);
nand UO_149 (O_149,N_24806,N_24848);
and UO_150 (O_150,N_24914,N_24982);
or UO_151 (O_151,N_24971,N_24986);
or UO_152 (O_152,N_24906,N_24962);
nand UO_153 (O_153,N_24979,N_24905);
xnor UO_154 (O_154,N_24865,N_24952);
nor UO_155 (O_155,N_24954,N_24941);
nand UO_156 (O_156,N_24847,N_24980);
and UO_157 (O_157,N_24990,N_24877);
nand UO_158 (O_158,N_24900,N_24914);
xnor UO_159 (O_159,N_24883,N_24861);
and UO_160 (O_160,N_24879,N_24857);
nor UO_161 (O_161,N_24947,N_24805);
nor UO_162 (O_162,N_24948,N_24860);
and UO_163 (O_163,N_24965,N_24919);
or UO_164 (O_164,N_24843,N_24929);
or UO_165 (O_165,N_24837,N_24927);
or UO_166 (O_166,N_24850,N_24972);
nor UO_167 (O_167,N_24953,N_24836);
xnor UO_168 (O_168,N_24913,N_24804);
or UO_169 (O_169,N_24993,N_24876);
nand UO_170 (O_170,N_24838,N_24880);
and UO_171 (O_171,N_24887,N_24954);
and UO_172 (O_172,N_24835,N_24895);
or UO_173 (O_173,N_24914,N_24860);
nand UO_174 (O_174,N_24941,N_24992);
nand UO_175 (O_175,N_24837,N_24990);
nand UO_176 (O_176,N_24885,N_24959);
and UO_177 (O_177,N_24853,N_24850);
nand UO_178 (O_178,N_24887,N_24934);
and UO_179 (O_179,N_24931,N_24915);
nor UO_180 (O_180,N_24967,N_24915);
nand UO_181 (O_181,N_24912,N_24889);
nand UO_182 (O_182,N_24996,N_24883);
or UO_183 (O_183,N_24864,N_24863);
and UO_184 (O_184,N_24967,N_24979);
or UO_185 (O_185,N_24977,N_24837);
nand UO_186 (O_186,N_24898,N_24998);
nor UO_187 (O_187,N_24923,N_24810);
nor UO_188 (O_188,N_24813,N_24977);
and UO_189 (O_189,N_24914,N_24890);
and UO_190 (O_190,N_24971,N_24903);
or UO_191 (O_191,N_24830,N_24818);
or UO_192 (O_192,N_24977,N_24997);
and UO_193 (O_193,N_24823,N_24848);
nand UO_194 (O_194,N_24989,N_24883);
xor UO_195 (O_195,N_24882,N_24869);
nor UO_196 (O_196,N_24981,N_24908);
or UO_197 (O_197,N_24826,N_24950);
xnor UO_198 (O_198,N_24982,N_24845);
nor UO_199 (O_199,N_24956,N_24965);
or UO_200 (O_200,N_24819,N_24872);
nor UO_201 (O_201,N_24891,N_24942);
and UO_202 (O_202,N_24868,N_24990);
and UO_203 (O_203,N_24986,N_24954);
nor UO_204 (O_204,N_24863,N_24936);
nor UO_205 (O_205,N_24901,N_24896);
and UO_206 (O_206,N_24974,N_24945);
and UO_207 (O_207,N_24911,N_24845);
nand UO_208 (O_208,N_24808,N_24904);
xor UO_209 (O_209,N_24919,N_24830);
nand UO_210 (O_210,N_24852,N_24904);
or UO_211 (O_211,N_24962,N_24849);
nand UO_212 (O_212,N_24974,N_24992);
and UO_213 (O_213,N_24894,N_24902);
nand UO_214 (O_214,N_24993,N_24801);
or UO_215 (O_215,N_24939,N_24970);
nor UO_216 (O_216,N_24924,N_24822);
and UO_217 (O_217,N_24813,N_24941);
xor UO_218 (O_218,N_24914,N_24847);
and UO_219 (O_219,N_24897,N_24882);
or UO_220 (O_220,N_24920,N_24884);
and UO_221 (O_221,N_24973,N_24937);
or UO_222 (O_222,N_24892,N_24887);
nor UO_223 (O_223,N_24857,N_24883);
nand UO_224 (O_224,N_24912,N_24860);
and UO_225 (O_225,N_24843,N_24811);
xor UO_226 (O_226,N_24983,N_24837);
or UO_227 (O_227,N_24988,N_24968);
nor UO_228 (O_228,N_24971,N_24962);
nand UO_229 (O_229,N_24987,N_24880);
and UO_230 (O_230,N_24935,N_24965);
xor UO_231 (O_231,N_24936,N_24812);
nor UO_232 (O_232,N_24822,N_24800);
or UO_233 (O_233,N_24893,N_24906);
or UO_234 (O_234,N_24952,N_24900);
and UO_235 (O_235,N_24878,N_24805);
nor UO_236 (O_236,N_24942,N_24862);
or UO_237 (O_237,N_24833,N_24940);
and UO_238 (O_238,N_24808,N_24948);
nor UO_239 (O_239,N_24819,N_24840);
xnor UO_240 (O_240,N_24974,N_24888);
nand UO_241 (O_241,N_24964,N_24887);
or UO_242 (O_242,N_24859,N_24900);
nand UO_243 (O_243,N_24818,N_24815);
or UO_244 (O_244,N_24825,N_24839);
nand UO_245 (O_245,N_24904,N_24996);
nand UO_246 (O_246,N_24929,N_24958);
nor UO_247 (O_247,N_24854,N_24902);
nor UO_248 (O_248,N_24821,N_24991);
nor UO_249 (O_249,N_24882,N_24916);
or UO_250 (O_250,N_24955,N_24990);
and UO_251 (O_251,N_24930,N_24800);
nand UO_252 (O_252,N_24913,N_24865);
nand UO_253 (O_253,N_24895,N_24832);
nor UO_254 (O_254,N_24866,N_24857);
or UO_255 (O_255,N_24863,N_24906);
nor UO_256 (O_256,N_24999,N_24834);
nor UO_257 (O_257,N_24808,N_24991);
or UO_258 (O_258,N_24891,N_24924);
or UO_259 (O_259,N_24961,N_24959);
nor UO_260 (O_260,N_24876,N_24832);
nand UO_261 (O_261,N_24951,N_24880);
nand UO_262 (O_262,N_24945,N_24944);
or UO_263 (O_263,N_24876,N_24991);
nand UO_264 (O_264,N_24856,N_24843);
nand UO_265 (O_265,N_24894,N_24809);
xor UO_266 (O_266,N_24892,N_24970);
nor UO_267 (O_267,N_24853,N_24841);
and UO_268 (O_268,N_24900,N_24854);
and UO_269 (O_269,N_24834,N_24801);
nand UO_270 (O_270,N_24893,N_24951);
nand UO_271 (O_271,N_24945,N_24831);
and UO_272 (O_272,N_24835,N_24968);
or UO_273 (O_273,N_24903,N_24941);
or UO_274 (O_274,N_24909,N_24974);
nand UO_275 (O_275,N_24908,N_24844);
nor UO_276 (O_276,N_24817,N_24871);
nand UO_277 (O_277,N_24910,N_24996);
and UO_278 (O_278,N_24898,N_24824);
or UO_279 (O_279,N_24936,N_24816);
and UO_280 (O_280,N_24951,N_24982);
xor UO_281 (O_281,N_24925,N_24857);
nor UO_282 (O_282,N_24865,N_24930);
and UO_283 (O_283,N_24927,N_24809);
nand UO_284 (O_284,N_24942,N_24883);
nand UO_285 (O_285,N_24823,N_24832);
nor UO_286 (O_286,N_24826,N_24816);
nand UO_287 (O_287,N_24983,N_24995);
or UO_288 (O_288,N_24889,N_24849);
or UO_289 (O_289,N_24850,N_24863);
or UO_290 (O_290,N_24878,N_24942);
and UO_291 (O_291,N_24875,N_24954);
and UO_292 (O_292,N_24833,N_24929);
nor UO_293 (O_293,N_24874,N_24979);
nor UO_294 (O_294,N_24986,N_24967);
or UO_295 (O_295,N_24883,N_24912);
nor UO_296 (O_296,N_24814,N_24963);
nor UO_297 (O_297,N_24804,N_24951);
nand UO_298 (O_298,N_24855,N_24938);
or UO_299 (O_299,N_24989,N_24889);
nor UO_300 (O_300,N_24892,N_24930);
and UO_301 (O_301,N_24867,N_24873);
or UO_302 (O_302,N_24826,N_24898);
nand UO_303 (O_303,N_24907,N_24840);
nor UO_304 (O_304,N_24956,N_24989);
or UO_305 (O_305,N_24997,N_24934);
and UO_306 (O_306,N_24913,N_24822);
nor UO_307 (O_307,N_24962,N_24859);
and UO_308 (O_308,N_24825,N_24863);
and UO_309 (O_309,N_24859,N_24850);
or UO_310 (O_310,N_24959,N_24933);
nor UO_311 (O_311,N_24828,N_24844);
and UO_312 (O_312,N_24924,N_24854);
and UO_313 (O_313,N_24853,N_24883);
or UO_314 (O_314,N_24926,N_24903);
nor UO_315 (O_315,N_24988,N_24989);
or UO_316 (O_316,N_24985,N_24935);
nor UO_317 (O_317,N_24997,N_24845);
and UO_318 (O_318,N_24810,N_24991);
nand UO_319 (O_319,N_24936,N_24892);
or UO_320 (O_320,N_24948,N_24830);
or UO_321 (O_321,N_24905,N_24885);
and UO_322 (O_322,N_24870,N_24836);
and UO_323 (O_323,N_24968,N_24962);
or UO_324 (O_324,N_24823,N_24830);
or UO_325 (O_325,N_24993,N_24937);
xnor UO_326 (O_326,N_24855,N_24909);
nand UO_327 (O_327,N_24942,N_24838);
and UO_328 (O_328,N_24866,N_24812);
or UO_329 (O_329,N_24834,N_24917);
or UO_330 (O_330,N_24821,N_24846);
and UO_331 (O_331,N_24857,N_24890);
nor UO_332 (O_332,N_24818,N_24894);
or UO_333 (O_333,N_24903,N_24952);
nor UO_334 (O_334,N_24864,N_24977);
or UO_335 (O_335,N_24888,N_24953);
xnor UO_336 (O_336,N_24832,N_24988);
or UO_337 (O_337,N_24849,N_24852);
nand UO_338 (O_338,N_24937,N_24814);
xor UO_339 (O_339,N_24821,N_24831);
and UO_340 (O_340,N_24882,N_24941);
and UO_341 (O_341,N_24835,N_24881);
xor UO_342 (O_342,N_24887,N_24987);
nor UO_343 (O_343,N_24907,N_24950);
nand UO_344 (O_344,N_24833,N_24960);
or UO_345 (O_345,N_24955,N_24903);
nor UO_346 (O_346,N_24824,N_24955);
nand UO_347 (O_347,N_24996,N_24833);
and UO_348 (O_348,N_24937,N_24825);
and UO_349 (O_349,N_24820,N_24847);
and UO_350 (O_350,N_24907,N_24913);
nor UO_351 (O_351,N_24862,N_24856);
xor UO_352 (O_352,N_24817,N_24991);
nor UO_353 (O_353,N_24858,N_24977);
and UO_354 (O_354,N_24912,N_24996);
xor UO_355 (O_355,N_24987,N_24996);
and UO_356 (O_356,N_24882,N_24952);
or UO_357 (O_357,N_24923,N_24883);
xor UO_358 (O_358,N_24955,N_24997);
nand UO_359 (O_359,N_24874,N_24836);
nor UO_360 (O_360,N_24808,N_24803);
and UO_361 (O_361,N_24840,N_24953);
nand UO_362 (O_362,N_24942,N_24887);
nor UO_363 (O_363,N_24855,N_24917);
nand UO_364 (O_364,N_24870,N_24881);
and UO_365 (O_365,N_24955,N_24994);
nor UO_366 (O_366,N_24961,N_24962);
nand UO_367 (O_367,N_24861,N_24892);
and UO_368 (O_368,N_24921,N_24995);
nor UO_369 (O_369,N_24882,N_24954);
nand UO_370 (O_370,N_24898,N_24814);
or UO_371 (O_371,N_24943,N_24818);
xnor UO_372 (O_372,N_24971,N_24871);
or UO_373 (O_373,N_24937,N_24885);
nor UO_374 (O_374,N_24874,N_24923);
nand UO_375 (O_375,N_24971,N_24842);
and UO_376 (O_376,N_24877,N_24836);
or UO_377 (O_377,N_24919,N_24944);
and UO_378 (O_378,N_24823,N_24981);
nor UO_379 (O_379,N_24960,N_24882);
nor UO_380 (O_380,N_24947,N_24898);
nand UO_381 (O_381,N_24802,N_24953);
nor UO_382 (O_382,N_24971,N_24827);
nor UO_383 (O_383,N_24803,N_24921);
and UO_384 (O_384,N_24857,N_24828);
nand UO_385 (O_385,N_24946,N_24845);
nand UO_386 (O_386,N_24901,N_24983);
and UO_387 (O_387,N_24932,N_24963);
xor UO_388 (O_388,N_24828,N_24820);
xor UO_389 (O_389,N_24841,N_24989);
nand UO_390 (O_390,N_24821,N_24939);
nor UO_391 (O_391,N_24955,N_24966);
and UO_392 (O_392,N_24854,N_24843);
nor UO_393 (O_393,N_24881,N_24915);
xor UO_394 (O_394,N_24967,N_24911);
nand UO_395 (O_395,N_24881,N_24955);
nand UO_396 (O_396,N_24981,N_24800);
nand UO_397 (O_397,N_24815,N_24870);
nand UO_398 (O_398,N_24882,N_24910);
xnor UO_399 (O_399,N_24856,N_24980);
nor UO_400 (O_400,N_24898,N_24823);
xor UO_401 (O_401,N_24895,N_24966);
nor UO_402 (O_402,N_24861,N_24839);
or UO_403 (O_403,N_24995,N_24874);
nand UO_404 (O_404,N_24805,N_24981);
nor UO_405 (O_405,N_24924,N_24903);
xor UO_406 (O_406,N_24966,N_24866);
and UO_407 (O_407,N_24865,N_24835);
and UO_408 (O_408,N_24825,N_24906);
nand UO_409 (O_409,N_24921,N_24827);
or UO_410 (O_410,N_24862,N_24881);
nor UO_411 (O_411,N_24922,N_24911);
nor UO_412 (O_412,N_24971,N_24889);
or UO_413 (O_413,N_24906,N_24960);
nor UO_414 (O_414,N_24854,N_24829);
nand UO_415 (O_415,N_24887,N_24893);
nor UO_416 (O_416,N_24978,N_24953);
nand UO_417 (O_417,N_24917,N_24878);
or UO_418 (O_418,N_24941,N_24847);
and UO_419 (O_419,N_24818,N_24826);
or UO_420 (O_420,N_24973,N_24801);
nand UO_421 (O_421,N_24901,N_24807);
nand UO_422 (O_422,N_24861,N_24938);
and UO_423 (O_423,N_24990,N_24863);
nor UO_424 (O_424,N_24856,N_24914);
xor UO_425 (O_425,N_24980,N_24971);
or UO_426 (O_426,N_24840,N_24926);
nor UO_427 (O_427,N_24834,N_24874);
nor UO_428 (O_428,N_24818,N_24882);
and UO_429 (O_429,N_24882,N_24949);
nand UO_430 (O_430,N_24853,N_24888);
nand UO_431 (O_431,N_24905,N_24962);
or UO_432 (O_432,N_24892,N_24906);
or UO_433 (O_433,N_24905,N_24975);
nand UO_434 (O_434,N_24836,N_24820);
nand UO_435 (O_435,N_24968,N_24985);
nor UO_436 (O_436,N_24938,N_24967);
xor UO_437 (O_437,N_24993,N_24932);
nor UO_438 (O_438,N_24802,N_24937);
and UO_439 (O_439,N_24847,N_24870);
and UO_440 (O_440,N_24867,N_24914);
nor UO_441 (O_441,N_24981,N_24804);
nor UO_442 (O_442,N_24952,N_24985);
xnor UO_443 (O_443,N_24993,N_24910);
nand UO_444 (O_444,N_24975,N_24994);
and UO_445 (O_445,N_24846,N_24906);
nor UO_446 (O_446,N_24882,N_24810);
and UO_447 (O_447,N_24945,N_24985);
or UO_448 (O_448,N_24862,N_24959);
or UO_449 (O_449,N_24843,N_24829);
nand UO_450 (O_450,N_24998,N_24971);
or UO_451 (O_451,N_24936,N_24937);
nand UO_452 (O_452,N_24828,N_24957);
nor UO_453 (O_453,N_24982,N_24892);
nand UO_454 (O_454,N_24949,N_24945);
and UO_455 (O_455,N_24875,N_24896);
nor UO_456 (O_456,N_24990,N_24946);
nor UO_457 (O_457,N_24922,N_24874);
and UO_458 (O_458,N_24907,N_24848);
nor UO_459 (O_459,N_24936,N_24838);
xnor UO_460 (O_460,N_24953,N_24967);
and UO_461 (O_461,N_24980,N_24846);
and UO_462 (O_462,N_24831,N_24805);
or UO_463 (O_463,N_24939,N_24842);
or UO_464 (O_464,N_24993,N_24810);
nand UO_465 (O_465,N_24891,N_24991);
xnor UO_466 (O_466,N_24992,N_24811);
and UO_467 (O_467,N_24930,N_24924);
or UO_468 (O_468,N_24814,N_24938);
or UO_469 (O_469,N_24832,N_24972);
xnor UO_470 (O_470,N_24886,N_24904);
nor UO_471 (O_471,N_24917,N_24978);
nor UO_472 (O_472,N_24867,N_24883);
or UO_473 (O_473,N_24934,N_24912);
nor UO_474 (O_474,N_24911,N_24910);
nand UO_475 (O_475,N_24886,N_24950);
and UO_476 (O_476,N_24807,N_24830);
xnor UO_477 (O_477,N_24824,N_24837);
nand UO_478 (O_478,N_24999,N_24853);
nor UO_479 (O_479,N_24993,N_24896);
xor UO_480 (O_480,N_24927,N_24885);
and UO_481 (O_481,N_24903,N_24932);
and UO_482 (O_482,N_24908,N_24818);
nand UO_483 (O_483,N_24889,N_24809);
or UO_484 (O_484,N_24822,N_24888);
nor UO_485 (O_485,N_24936,N_24989);
nand UO_486 (O_486,N_24873,N_24972);
nor UO_487 (O_487,N_24913,N_24852);
nand UO_488 (O_488,N_24836,N_24892);
or UO_489 (O_489,N_24811,N_24812);
nand UO_490 (O_490,N_24984,N_24867);
and UO_491 (O_491,N_24951,N_24828);
and UO_492 (O_492,N_24902,N_24939);
and UO_493 (O_493,N_24947,N_24849);
or UO_494 (O_494,N_24843,N_24923);
nor UO_495 (O_495,N_24840,N_24870);
or UO_496 (O_496,N_24951,N_24824);
and UO_497 (O_497,N_24824,N_24807);
and UO_498 (O_498,N_24950,N_24860);
nand UO_499 (O_499,N_24844,N_24950);
or UO_500 (O_500,N_24841,N_24900);
and UO_501 (O_501,N_24908,N_24895);
nand UO_502 (O_502,N_24935,N_24862);
and UO_503 (O_503,N_24956,N_24973);
nor UO_504 (O_504,N_24949,N_24930);
and UO_505 (O_505,N_24849,N_24989);
xor UO_506 (O_506,N_24890,N_24931);
nand UO_507 (O_507,N_24956,N_24841);
nand UO_508 (O_508,N_24965,N_24983);
and UO_509 (O_509,N_24831,N_24977);
nor UO_510 (O_510,N_24889,N_24902);
nor UO_511 (O_511,N_24961,N_24852);
nor UO_512 (O_512,N_24836,N_24839);
nor UO_513 (O_513,N_24935,N_24827);
nor UO_514 (O_514,N_24803,N_24896);
nor UO_515 (O_515,N_24827,N_24970);
and UO_516 (O_516,N_24999,N_24920);
nor UO_517 (O_517,N_24867,N_24965);
nor UO_518 (O_518,N_24806,N_24932);
or UO_519 (O_519,N_24806,N_24822);
or UO_520 (O_520,N_24880,N_24897);
or UO_521 (O_521,N_24952,N_24825);
and UO_522 (O_522,N_24961,N_24997);
and UO_523 (O_523,N_24833,N_24943);
xnor UO_524 (O_524,N_24991,N_24863);
nor UO_525 (O_525,N_24937,N_24853);
nor UO_526 (O_526,N_24832,N_24849);
and UO_527 (O_527,N_24929,N_24887);
or UO_528 (O_528,N_24959,N_24909);
or UO_529 (O_529,N_24989,N_24813);
nand UO_530 (O_530,N_24846,N_24898);
or UO_531 (O_531,N_24918,N_24939);
or UO_532 (O_532,N_24938,N_24971);
nor UO_533 (O_533,N_24933,N_24847);
and UO_534 (O_534,N_24909,N_24941);
or UO_535 (O_535,N_24883,N_24858);
nand UO_536 (O_536,N_24882,N_24980);
and UO_537 (O_537,N_24807,N_24985);
xor UO_538 (O_538,N_24866,N_24997);
nor UO_539 (O_539,N_24942,N_24911);
nand UO_540 (O_540,N_24832,N_24947);
or UO_541 (O_541,N_24986,N_24831);
xnor UO_542 (O_542,N_24812,N_24851);
xor UO_543 (O_543,N_24866,N_24891);
nand UO_544 (O_544,N_24927,N_24801);
nand UO_545 (O_545,N_24850,N_24882);
or UO_546 (O_546,N_24989,N_24912);
nand UO_547 (O_547,N_24852,N_24992);
nand UO_548 (O_548,N_24950,N_24887);
nor UO_549 (O_549,N_24981,N_24827);
nor UO_550 (O_550,N_24979,N_24829);
or UO_551 (O_551,N_24810,N_24829);
nand UO_552 (O_552,N_24948,N_24986);
and UO_553 (O_553,N_24854,N_24857);
and UO_554 (O_554,N_24909,N_24966);
nand UO_555 (O_555,N_24880,N_24969);
nand UO_556 (O_556,N_24816,N_24991);
or UO_557 (O_557,N_24912,N_24843);
nor UO_558 (O_558,N_24941,N_24900);
and UO_559 (O_559,N_24971,N_24911);
nand UO_560 (O_560,N_24906,N_24901);
nand UO_561 (O_561,N_24861,N_24988);
or UO_562 (O_562,N_24839,N_24806);
or UO_563 (O_563,N_24905,N_24828);
and UO_564 (O_564,N_24946,N_24834);
nor UO_565 (O_565,N_24917,N_24850);
or UO_566 (O_566,N_24896,N_24930);
xnor UO_567 (O_567,N_24993,N_24807);
nand UO_568 (O_568,N_24888,N_24947);
nand UO_569 (O_569,N_24927,N_24939);
nor UO_570 (O_570,N_24976,N_24850);
nand UO_571 (O_571,N_24955,N_24979);
nand UO_572 (O_572,N_24892,N_24983);
and UO_573 (O_573,N_24896,N_24970);
nand UO_574 (O_574,N_24902,N_24878);
xor UO_575 (O_575,N_24927,N_24830);
nor UO_576 (O_576,N_24921,N_24926);
and UO_577 (O_577,N_24931,N_24965);
xnor UO_578 (O_578,N_24971,N_24952);
nand UO_579 (O_579,N_24857,N_24984);
or UO_580 (O_580,N_24957,N_24919);
or UO_581 (O_581,N_24897,N_24873);
and UO_582 (O_582,N_24969,N_24935);
or UO_583 (O_583,N_24940,N_24982);
nor UO_584 (O_584,N_24994,N_24954);
and UO_585 (O_585,N_24848,N_24951);
and UO_586 (O_586,N_24961,N_24856);
or UO_587 (O_587,N_24873,N_24957);
and UO_588 (O_588,N_24963,N_24803);
nand UO_589 (O_589,N_24914,N_24839);
nor UO_590 (O_590,N_24860,N_24853);
or UO_591 (O_591,N_24925,N_24987);
and UO_592 (O_592,N_24994,N_24959);
nand UO_593 (O_593,N_24897,N_24966);
nor UO_594 (O_594,N_24969,N_24848);
and UO_595 (O_595,N_24900,N_24902);
nand UO_596 (O_596,N_24983,N_24835);
nor UO_597 (O_597,N_24820,N_24920);
nor UO_598 (O_598,N_24910,N_24800);
and UO_599 (O_599,N_24861,N_24827);
nand UO_600 (O_600,N_24855,N_24823);
nor UO_601 (O_601,N_24941,N_24947);
or UO_602 (O_602,N_24984,N_24829);
xor UO_603 (O_603,N_24843,N_24921);
or UO_604 (O_604,N_24803,N_24822);
nand UO_605 (O_605,N_24834,N_24823);
xnor UO_606 (O_606,N_24989,N_24902);
or UO_607 (O_607,N_24857,N_24920);
nor UO_608 (O_608,N_24989,N_24863);
and UO_609 (O_609,N_24880,N_24882);
and UO_610 (O_610,N_24925,N_24905);
or UO_611 (O_611,N_24934,N_24929);
xor UO_612 (O_612,N_24942,N_24902);
and UO_613 (O_613,N_24842,N_24831);
nand UO_614 (O_614,N_24823,N_24877);
or UO_615 (O_615,N_24823,N_24946);
or UO_616 (O_616,N_24952,N_24997);
nor UO_617 (O_617,N_24828,N_24908);
nand UO_618 (O_618,N_24886,N_24965);
or UO_619 (O_619,N_24896,N_24880);
nand UO_620 (O_620,N_24890,N_24845);
nand UO_621 (O_621,N_24898,N_24907);
and UO_622 (O_622,N_24817,N_24850);
or UO_623 (O_623,N_24962,N_24826);
nand UO_624 (O_624,N_24866,N_24803);
nand UO_625 (O_625,N_24991,N_24968);
and UO_626 (O_626,N_24933,N_24872);
xnor UO_627 (O_627,N_24948,N_24846);
or UO_628 (O_628,N_24898,N_24881);
nor UO_629 (O_629,N_24967,N_24932);
and UO_630 (O_630,N_24887,N_24870);
nand UO_631 (O_631,N_24958,N_24836);
nand UO_632 (O_632,N_24903,N_24886);
and UO_633 (O_633,N_24949,N_24879);
or UO_634 (O_634,N_24821,N_24950);
nor UO_635 (O_635,N_24838,N_24851);
nor UO_636 (O_636,N_24987,N_24946);
nor UO_637 (O_637,N_24938,N_24999);
and UO_638 (O_638,N_24885,N_24825);
nand UO_639 (O_639,N_24859,N_24992);
nor UO_640 (O_640,N_24888,N_24884);
nand UO_641 (O_641,N_24952,N_24891);
nand UO_642 (O_642,N_24851,N_24915);
nand UO_643 (O_643,N_24882,N_24913);
or UO_644 (O_644,N_24944,N_24825);
nand UO_645 (O_645,N_24940,N_24828);
or UO_646 (O_646,N_24932,N_24832);
nand UO_647 (O_647,N_24939,N_24995);
nand UO_648 (O_648,N_24844,N_24825);
or UO_649 (O_649,N_24893,N_24868);
or UO_650 (O_650,N_24895,N_24819);
nand UO_651 (O_651,N_24847,N_24961);
nor UO_652 (O_652,N_24902,N_24874);
nand UO_653 (O_653,N_24967,N_24989);
xnor UO_654 (O_654,N_24877,N_24894);
nor UO_655 (O_655,N_24937,N_24922);
and UO_656 (O_656,N_24958,N_24903);
nor UO_657 (O_657,N_24874,N_24868);
nand UO_658 (O_658,N_24801,N_24886);
and UO_659 (O_659,N_24921,N_24939);
nor UO_660 (O_660,N_24812,N_24890);
or UO_661 (O_661,N_24894,N_24803);
nand UO_662 (O_662,N_24834,N_24911);
nand UO_663 (O_663,N_24838,N_24800);
nor UO_664 (O_664,N_24953,N_24858);
and UO_665 (O_665,N_24933,N_24938);
xor UO_666 (O_666,N_24959,N_24837);
nor UO_667 (O_667,N_24846,N_24848);
or UO_668 (O_668,N_24831,N_24834);
xor UO_669 (O_669,N_24823,N_24999);
xnor UO_670 (O_670,N_24930,N_24999);
nor UO_671 (O_671,N_24859,N_24932);
nand UO_672 (O_672,N_24898,N_24980);
and UO_673 (O_673,N_24815,N_24877);
and UO_674 (O_674,N_24807,N_24864);
and UO_675 (O_675,N_24979,N_24858);
and UO_676 (O_676,N_24908,N_24961);
xor UO_677 (O_677,N_24935,N_24974);
or UO_678 (O_678,N_24911,N_24866);
or UO_679 (O_679,N_24848,N_24861);
nor UO_680 (O_680,N_24979,N_24984);
nor UO_681 (O_681,N_24842,N_24904);
nand UO_682 (O_682,N_24839,N_24850);
nand UO_683 (O_683,N_24921,N_24851);
and UO_684 (O_684,N_24808,N_24824);
and UO_685 (O_685,N_24822,N_24894);
nor UO_686 (O_686,N_24839,N_24987);
nor UO_687 (O_687,N_24879,N_24888);
nand UO_688 (O_688,N_24907,N_24836);
or UO_689 (O_689,N_24802,N_24863);
nand UO_690 (O_690,N_24971,N_24894);
or UO_691 (O_691,N_24865,N_24851);
nand UO_692 (O_692,N_24952,N_24940);
or UO_693 (O_693,N_24870,N_24960);
or UO_694 (O_694,N_24815,N_24849);
or UO_695 (O_695,N_24893,N_24896);
and UO_696 (O_696,N_24973,N_24942);
or UO_697 (O_697,N_24946,N_24885);
and UO_698 (O_698,N_24924,N_24864);
or UO_699 (O_699,N_24933,N_24802);
xnor UO_700 (O_700,N_24971,N_24972);
xnor UO_701 (O_701,N_24809,N_24937);
nand UO_702 (O_702,N_24837,N_24839);
nor UO_703 (O_703,N_24947,N_24801);
or UO_704 (O_704,N_24804,N_24921);
nand UO_705 (O_705,N_24847,N_24855);
and UO_706 (O_706,N_24956,N_24976);
nor UO_707 (O_707,N_24937,N_24986);
nor UO_708 (O_708,N_24942,N_24804);
nand UO_709 (O_709,N_24907,N_24941);
or UO_710 (O_710,N_24890,N_24971);
nor UO_711 (O_711,N_24995,N_24916);
nor UO_712 (O_712,N_24991,N_24946);
nor UO_713 (O_713,N_24855,N_24903);
xor UO_714 (O_714,N_24815,N_24922);
nand UO_715 (O_715,N_24829,N_24909);
or UO_716 (O_716,N_24938,N_24850);
or UO_717 (O_717,N_24838,N_24945);
and UO_718 (O_718,N_24883,N_24839);
nor UO_719 (O_719,N_24929,N_24947);
nor UO_720 (O_720,N_24970,N_24997);
nor UO_721 (O_721,N_24819,N_24836);
nor UO_722 (O_722,N_24995,N_24824);
and UO_723 (O_723,N_24973,N_24852);
nand UO_724 (O_724,N_24922,N_24876);
nand UO_725 (O_725,N_24832,N_24907);
xor UO_726 (O_726,N_24924,N_24858);
and UO_727 (O_727,N_24872,N_24998);
nand UO_728 (O_728,N_24935,N_24837);
xor UO_729 (O_729,N_24998,N_24947);
nand UO_730 (O_730,N_24819,N_24964);
nor UO_731 (O_731,N_24813,N_24860);
nor UO_732 (O_732,N_24916,N_24973);
and UO_733 (O_733,N_24832,N_24801);
nor UO_734 (O_734,N_24827,N_24977);
nand UO_735 (O_735,N_24855,N_24978);
or UO_736 (O_736,N_24930,N_24926);
nor UO_737 (O_737,N_24826,N_24949);
or UO_738 (O_738,N_24972,N_24843);
and UO_739 (O_739,N_24841,N_24890);
or UO_740 (O_740,N_24880,N_24985);
nand UO_741 (O_741,N_24832,N_24934);
nor UO_742 (O_742,N_24942,N_24975);
xnor UO_743 (O_743,N_24815,N_24953);
or UO_744 (O_744,N_24820,N_24910);
or UO_745 (O_745,N_24969,N_24940);
and UO_746 (O_746,N_24911,N_24948);
or UO_747 (O_747,N_24840,N_24892);
and UO_748 (O_748,N_24894,N_24960);
nand UO_749 (O_749,N_24940,N_24851);
nor UO_750 (O_750,N_24845,N_24972);
and UO_751 (O_751,N_24922,N_24998);
and UO_752 (O_752,N_24825,N_24881);
nand UO_753 (O_753,N_24911,N_24950);
and UO_754 (O_754,N_24918,N_24895);
or UO_755 (O_755,N_24899,N_24874);
nand UO_756 (O_756,N_24945,N_24837);
or UO_757 (O_757,N_24999,N_24871);
xor UO_758 (O_758,N_24903,N_24891);
and UO_759 (O_759,N_24979,N_24959);
nand UO_760 (O_760,N_24915,N_24925);
or UO_761 (O_761,N_24877,N_24930);
nor UO_762 (O_762,N_24888,N_24915);
and UO_763 (O_763,N_24815,N_24940);
nor UO_764 (O_764,N_24940,N_24955);
nor UO_765 (O_765,N_24834,N_24979);
or UO_766 (O_766,N_24960,N_24841);
nor UO_767 (O_767,N_24821,N_24892);
or UO_768 (O_768,N_24820,N_24886);
nand UO_769 (O_769,N_24841,N_24851);
and UO_770 (O_770,N_24934,N_24881);
or UO_771 (O_771,N_24979,N_24972);
and UO_772 (O_772,N_24925,N_24963);
xor UO_773 (O_773,N_24820,N_24851);
nand UO_774 (O_774,N_24978,N_24998);
xor UO_775 (O_775,N_24943,N_24908);
nand UO_776 (O_776,N_24817,N_24833);
xor UO_777 (O_777,N_24949,N_24849);
and UO_778 (O_778,N_24894,N_24882);
xnor UO_779 (O_779,N_24889,N_24828);
or UO_780 (O_780,N_24916,N_24989);
and UO_781 (O_781,N_24980,N_24852);
xor UO_782 (O_782,N_24880,N_24918);
nor UO_783 (O_783,N_24891,N_24801);
or UO_784 (O_784,N_24926,N_24883);
nand UO_785 (O_785,N_24966,N_24820);
or UO_786 (O_786,N_24995,N_24937);
and UO_787 (O_787,N_24854,N_24890);
nor UO_788 (O_788,N_24881,N_24932);
nand UO_789 (O_789,N_24927,N_24874);
and UO_790 (O_790,N_24958,N_24995);
nor UO_791 (O_791,N_24980,N_24924);
nor UO_792 (O_792,N_24992,N_24913);
nor UO_793 (O_793,N_24979,N_24854);
and UO_794 (O_794,N_24977,N_24871);
nor UO_795 (O_795,N_24917,N_24940);
nor UO_796 (O_796,N_24802,N_24998);
or UO_797 (O_797,N_24878,N_24874);
and UO_798 (O_798,N_24960,N_24903);
xor UO_799 (O_799,N_24865,N_24898);
nor UO_800 (O_800,N_24967,N_24855);
and UO_801 (O_801,N_24947,N_24950);
nand UO_802 (O_802,N_24838,N_24884);
nand UO_803 (O_803,N_24962,N_24955);
or UO_804 (O_804,N_24949,N_24855);
nand UO_805 (O_805,N_24964,N_24938);
nor UO_806 (O_806,N_24982,N_24886);
and UO_807 (O_807,N_24819,N_24870);
xnor UO_808 (O_808,N_24987,N_24952);
and UO_809 (O_809,N_24923,N_24909);
and UO_810 (O_810,N_24877,N_24967);
and UO_811 (O_811,N_24986,N_24844);
or UO_812 (O_812,N_24860,N_24800);
nand UO_813 (O_813,N_24883,N_24881);
or UO_814 (O_814,N_24823,N_24801);
nor UO_815 (O_815,N_24908,N_24970);
nand UO_816 (O_816,N_24947,N_24901);
or UO_817 (O_817,N_24867,N_24943);
nand UO_818 (O_818,N_24921,N_24903);
nand UO_819 (O_819,N_24826,N_24975);
nand UO_820 (O_820,N_24904,N_24963);
nand UO_821 (O_821,N_24812,N_24949);
nor UO_822 (O_822,N_24816,N_24828);
xnor UO_823 (O_823,N_24937,N_24921);
or UO_824 (O_824,N_24855,N_24801);
and UO_825 (O_825,N_24956,N_24886);
or UO_826 (O_826,N_24900,N_24937);
and UO_827 (O_827,N_24836,N_24896);
nor UO_828 (O_828,N_24879,N_24828);
nor UO_829 (O_829,N_24823,N_24954);
or UO_830 (O_830,N_24979,N_24921);
nand UO_831 (O_831,N_24983,N_24975);
and UO_832 (O_832,N_24975,N_24917);
nand UO_833 (O_833,N_24871,N_24959);
nand UO_834 (O_834,N_24903,N_24969);
nand UO_835 (O_835,N_24924,N_24945);
nand UO_836 (O_836,N_24981,N_24811);
nand UO_837 (O_837,N_24905,N_24982);
or UO_838 (O_838,N_24914,N_24980);
nor UO_839 (O_839,N_24856,N_24941);
nand UO_840 (O_840,N_24882,N_24867);
xor UO_841 (O_841,N_24903,N_24947);
and UO_842 (O_842,N_24815,N_24905);
nand UO_843 (O_843,N_24939,N_24904);
and UO_844 (O_844,N_24887,N_24948);
nor UO_845 (O_845,N_24841,N_24857);
or UO_846 (O_846,N_24979,N_24932);
nand UO_847 (O_847,N_24937,N_24924);
nor UO_848 (O_848,N_24980,N_24813);
nand UO_849 (O_849,N_24814,N_24893);
and UO_850 (O_850,N_24818,N_24982);
and UO_851 (O_851,N_24850,N_24875);
and UO_852 (O_852,N_24837,N_24864);
or UO_853 (O_853,N_24864,N_24819);
nand UO_854 (O_854,N_24836,N_24824);
and UO_855 (O_855,N_24811,N_24922);
xor UO_856 (O_856,N_24996,N_24957);
xor UO_857 (O_857,N_24986,N_24807);
or UO_858 (O_858,N_24994,N_24896);
or UO_859 (O_859,N_24944,N_24839);
nor UO_860 (O_860,N_24952,N_24992);
xor UO_861 (O_861,N_24856,N_24921);
and UO_862 (O_862,N_24986,N_24916);
or UO_863 (O_863,N_24847,N_24825);
nand UO_864 (O_864,N_24953,N_24916);
nor UO_865 (O_865,N_24910,N_24946);
or UO_866 (O_866,N_24882,N_24829);
nor UO_867 (O_867,N_24869,N_24953);
xnor UO_868 (O_868,N_24844,N_24955);
nor UO_869 (O_869,N_24860,N_24807);
xor UO_870 (O_870,N_24819,N_24971);
nor UO_871 (O_871,N_24832,N_24880);
or UO_872 (O_872,N_24972,N_24862);
and UO_873 (O_873,N_24962,N_24876);
nand UO_874 (O_874,N_24877,N_24903);
nand UO_875 (O_875,N_24961,N_24855);
nor UO_876 (O_876,N_24855,N_24963);
and UO_877 (O_877,N_24842,N_24950);
and UO_878 (O_878,N_24884,N_24853);
nor UO_879 (O_879,N_24911,N_24980);
nand UO_880 (O_880,N_24941,N_24843);
xor UO_881 (O_881,N_24949,N_24863);
nand UO_882 (O_882,N_24920,N_24990);
nand UO_883 (O_883,N_24815,N_24950);
xnor UO_884 (O_884,N_24879,N_24951);
or UO_885 (O_885,N_24820,N_24849);
nand UO_886 (O_886,N_24811,N_24908);
or UO_887 (O_887,N_24969,N_24876);
and UO_888 (O_888,N_24975,N_24865);
nand UO_889 (O_889,N_24864,N_24952);
nand UO_890 (O_890,N_24911,N_24886);
nor UO_891 (O_891,N_24816,N_24971);
or UO_892 (O_892,N_24854,N_24870);
or UO_893 (O_893,N_24888,N_24845);
xor UO_894 (O_894,N_24846,N_24911);
and UO_895 (O_895,N_24875,N_24964);
nand UO_896 (O_896,N_24964,N_24950);
and UO_897 (O_897,N_24904,N_24877);
nand UO_898 (O_898,N_24936,N_24848);
and UO_899 (O_899,N_24880,N_24937);
or UO_900 (O_900,N_24956,N_24818);
nand UO_901 (O_901,N_24874,N_24994);
nand UO_902 (O_902,N_24954,N_24824);
nand UO_903 (O_903,N_24842,N_24965);
xnor UO_904 (O_904,N_24822,N_24863);
or UO_905 (O_905,N_24934,N_24804);
and UO_906 (O_906,N_24953,N_24996);
nand UO_907 (O_907,N_24861,N_24953);
and UO_908 (O_908,N_24870,N_24827);
and UO_909 (O_909,N_24907,N_24888);
nand UO_910 (O_910,N_24868,N_24892);
and UO_911 (O_911,N_24884,N_24818);
nand UO_912 (O_912,N_24938,N_24808);
and UO_913 (O_913,N_24964,N_24811);
nor UO_914 (O_914,N_24962,N_24843);
nor UO_915 (O_915,N_24874,N_24945);
or UO_916 (O_916,N_24872,N_24813);
nand UO_917 (O_917,N_24994,N_24870);
or UO_918 (O_918,N_24931,N_24843);
or UO_919 (O_919,N_24923,N_24995);
or UO_920 (O_920,N_24855,N_24970);
nor UO_921 (O_921,N_24951,N_24872);
nor UO_922 (O_922,N_24978,N_24913);
xor UO_923 (O_923,N_24884,N_24937);
xor UO_924 (O_924,N_24938,N_24915);
or UO_925 (O_925,N_24992,N_24892);
nand UO_926 (O_926,N_24963,N_24805);
or UO_927 (O_927,N_24842,N_24827);
and UO_928 (O_928,N_24856,N_24952);
and UO_929 (O_929,N_24820,N_24941);
xor UO_930 (O_930,N_24849,N_24891);
and UO_931 (O_931,N_24981,N_24914);
nor UO_932 (O_932,N_24865,N_24877);
xor UO_933 (O_933,N_24812,N_24887);
and UO_934 (O_934,N_24920,N_24827);
nand UO_935 (O_935,N_24806,N_24861);
or UO_936 (O_936,N_24890,N_24904);
xnor UO_937 (O_937,N_24810,N_24843);
nor UO_938 (O_938,N_24848,N_24855);
or UO_939 (O_939,N_24988,N_24969);
and UO_940 (O_940,N_24943,N_24803);
nand UO_941 (O_941,N_24816,N_24872);
or UO_942 (O_942,N_24928,N_24926);
nor UO_943 (O_943,N_24942,N_24892);
and UO_944 (O_944,N_24822,N_24864);
or UO_945 (O_945,N_24993,N_24880);
nor UO_946 (O_946,N_24922,N_24829);
or UO_947 (O_947,N_24998,N_24919);
or UO_948 (O_948,N_24972,N_24821);
and UO_949 (O_949,N_24948,N_24897);
nor UO_950 (O_950,N_24881,N_24801);
xnor UO_951 (O_951,N_24852,N_24949);
and UO_952 (O_952,N_24967,N_24890);
or UO_953 (O_953,N_24811,N_24888);
nand UO_954 (O_954,N_24973,N_24947);
nor UO_955 (O_955,N_24863,N_24820);
xor UO_956 (O_956,N_24827,N_24896);
or UO_957 (O_957,N_24863,N_24962);
or UO_958 (O_958,N_24902,N_24907);
and UO_959 (O_959,N_24845,N_24958);
nor UO_960 (O_960,N_24928,N_24925);
xnor UO_961 (O_961,N_24845,N_24962);
nor UO_962 (O_962,N_24987,N_24993);
or UO_963 (O_963,N_24811,N_24834);
nand UO_964 (O_964,N_24837,N_24955);
nor UO_965 (O_965,N_24802,N_24985);
or UO_966 (O_966,N_24959,N_24939);
nand UO_967 (O_967,N_24819,N_24903);
nand UO_968 (O_968,N_24931,N_24998);
xor UO_969 (O_969,N_24928,N_24905);
and UO_970 (O_970,N_24801,N_24827);
nor UO_971 (O_971,N_24966,N_24860);
nor UO_972 (O_972,N_24923,N_24832);
nor UO_973 (O_973,N_24894,N_24842);
nor UO_974 (O_974,N_24821,N_24891);
or UO_975 (O_975,N_24993,N_24846);
nand UO_976 (O_976,N_24839,N_24979);
nor UO_977 (O_977,N_24995,N_24904);
nand UO_978 (O_978,N_24906,N_24992);
nand UO_979 (O_979,N_24950,N_24946);
xor UO_980 (O_980,N_24817,N_24875);
nor UO_981 (O_981,N_24813,N_24957);
xnor UO_982 (O_982,N_24886,N_24979);
nor UO_983 (O_983,N_24993,N_24912);
nand UO_984 (O_984,N_24874,N_24889);
or UO_985 (O_985,N_24944,N_24854);
and UO_986 (O_986,N_24976,N_24931);
xnor UO_987 (O_987,N_24889,N_24993);
and UO_988 (O_988,N_24803,N_24856);
and UO_989 (O_989,N_24887,N_24904);
nor UO_990 (O_990,N_24859,N_24917);
or UO_991 (O_991,N_24955,N_24915);
and UO_992 (O_992,N_24961,N_24983);
or UO_993 (O_993,N_24891,N_24861);
and UO_994 (O_994,N_24830,N_24971);
and UO_995 (O_995,N_24877,N_24926);
xnor UO_996 (O_996,N_24887,N_24924);
and UO_997 (O_997,N_24897,N_24822);
nor UO_998 (O_998,N_24905,N_24930);
nor UO_999 (O_999,N_24997,N_24942);
and UO_1000 (O_1000,N_24942,N_24935);
nand UO_1001 (O_1001,N_24848,N_24860);
or UO_1002 (O_1002,N_24998,N_24942);
nor UO_1003 (O_1003,N_24869,N_24928);
nand UO_1004 (O_1004,N_24997,N_24853);
and UO_1005 (O_1005,N_24936,N_24955);
or UO_1006 (O_1006,N_24862,N_24934);
nor UO_1007 (O_1007,N_24899,N_24849);
and UO_1008 (O_1008,N_24816,N_24906);
or UO_1009 (O_1009,N_24813,N_24952);
nand UO_1010 (O_1010,N_24960,N_24815);
and UO_1011 (O_1011,N_24997,N_24926);
nand UO_1012 (O_1012,N_24975,N_24848);
nand UO_1013 (O_1013,N_24866,N_24805);
and UO_1014 (O_1014,N_24841,N_24905);
nand UO_1015 (O_1015,N_24911,N_24992);
nand UO_1016 (O_1016,N_24841,N_24941);
nand UO_1017 (O_1017,N_24865,N_24946);
or UO_1018 (O_1018,N_24922,N_24893);
nor UO_1019 (O_1019,N_24863,N_24993);
nand UO_1020 (O_1020,N_24954,N_24950);
nor UO_1021 (O_1021,N_24875,N_24877);
nor UO_1022 (O_1022,N_24952,N_24954);
and UO_1023 (O_1023,N_24829,N_24998);
or UO_1024 (O_1024,N_24818,N_24889);
or UO_1025 (O_1025,N_24857,N_24872);
nor UO_1026 (O_1026,N_24804,N_24825);
nor UO_1027 (O_1027,N_24994,N_24853);
nor UO_1028 (O_1028,N_24815,N_24851);
nand UO_1029 (O_1029,N_24963,N_24965);
nand UO_1030 (O_1030,N_24805,N_24889);
and UO_1031 (O_1031,N_24893,N_24946);
nand UO_1032 (O_1032,N_24878,N_24922);
nand UO_1033 (O_1033,N_24813,N_24892);
nand UO_1034 (O_1034,N_24958,N_24813);
and UO_1035 (O_1035,N_24875,N_24854);
and UO_1036 (O_1036,N_24909,N_24935);
and UO_1037 (O_1037,N_24853,N_24965);
xnor UO_1038 (O_1038,N_24959,N_24942);
nand UO_1039 (O_1039,N_24875,N_24893);
nand UO_1040 (O_1040,N_24861,N_24996);
and UO_1041 (O_1041,N_24953,N_24842);
nor UO_1042 (O_1042,N_24896,N_24969);
nand UO_1043 (O_1043,N_24853,N_24927);
and UO_1044 (O_1044,N_24987,N_24874);
nor UO_1045 (O_1045,N_24809,N_24998);
and UO_1046 (O_1046,N_24868,N_24823);
nor UO_1047 (O_1047,N_24877,N_24813);
xor UO_1048 (O_1048,N_24834,N_24929);
nor UO_1049 (O_1049,N_24844,N_24902);
or UO_1050 (O_1050,N_24872,N_24806);
and UO_1051 (O_1051,N_24814,N_24840);
nor UO_1052 (O_1052,N_24992,N_24813);
nor UO_1053 (O_1053,N_24908,N_24894);
or UO_1054 (O_1054,N_24806,N_24999);
xnor UO_1055 (O_1055,N_24938,N_24974);
nand UO_1056 (O_1056,N_24865,N_24847);
or UO_1057 (O_1057,N_24958,N_24893);
nand UO_1058 (O_1058,N_24827,N_24832);
or UO_1059 (O_1059,N_24989,N_24866);
and UO_1060 (O_1060,N_24869,N_24850);
or UO_1061 (O_1061,N_24970,N_24821);
or UO_1062 (O_1062,N_24994,N_24889);
and UO_1063 (O_1063,N_24947,N_24852);
nand UO_1064 (O_1064,N_24832,N_24965);
and UO_1065 (O_1065,N_24805,N_24965);
nor UO_1066 (O_1066,N_24892,N_24873);
or UO_1067 (O_1067,N_24943,N_24905);
or UO_1068 (O_1068,N_24929,N_24856);
nor UO_1069 (O_1069,N_24968,N_24811);
or UO_1070 (O_1070,N_24903,N_24862);
nor UO_1071 (O_1071,N_24884,N_24972);
or UO_1072 (O_1072,N_24844,N_24808);
nor UO_1073 (O_1073,N_24909,N_24980);
nor UO_1074 (O_1074,N_24921,N_24836);
nor UO_1075 (O_1075,N_24934,N_24977);
and UO_1076 (O_1076,N_24993,N_24984);
and UO_1077 (O_1077,N_24805,N_24880);
nor UO_1078 (O_1078,N_24977,N_24816);
nand UO_1079 (O_1079,N_24861,N_24928);
xnor UO_1080 (O_1080,N_24869,N_24899);
or UO_1081 (O_1081,N_24829,N_24802);
xnor UO_1082 (O_1082,N_24900,N_24942);
and UO_1083 (O_1083,N_24860,N_24957);
nor UO_1084 (O_1084,N_24946,N_24864);
xnor UO_1085 (O_1085,N_24880,N_24995);
and UO_1086 (O_1086,N_24867,N_24901);
nand UO_1087 (O_1087,N_24930,N_24858);
and UO_1088 (O_1088,N_24973,N_24936);
or UO_1089 (O_1089,N_24903,N_24849);
xor UO_1090 (O_1090,N_24830,N_24988);
nand UO_1091 (O_1091,N_24991,N_24903);
or UO_1092 (O_1092,N_24911,N_24977);
or UO_1093 (O_1093,N_24874,N_24844);
and UO_1094 (O_1094,N_24920,N_24804);
or UO_1095 (O_1095,N_24941,N_24842);
nand UO_1096 (O_1096,N_24976,N_24875);
nand UO_1097 (O_1097,N_24864,N_24885);
nand UO_1098 (O_1098,N_24811,N_24813);
xor UO_1099 (O_1099,N_24930,N_24955);
xor UO_1100 (O_1100,N_24915,N_24906);
nand UO_1101 (O_1101,N_24828,N_24853);
and UO_1102 (O_1102,N_24965,N_24976);
or UO_1103 (O_1103,N_24965,N_24972);
nor UO_1104 (O_1104,N_24970,N_24918);
nand UO_1105 (O_1105,N_24949,N_24864);
and UO_1106 (O_1106,N_24900,N_24825);
or UO_1107 (O_1107,N_24853,N_24861);
or UO_1108 (O_1108,N_24925,N_24819);
and UO_1109 (O_1109,N_24910,N_24890);
nand UO_1110 (O_1110,N_24880,N_24802);
nor UO_1111 (O_1111,N_24939,N_24983);
nor UO_1112 (O_1112,N_24995,N_24837);
nand UO_1113 (O_1113,N_24914,N_24998);
nand UO_1114 (O_1114,N_24918,N_24930);
nor UO_1115 (O_1115,N_24830,N_24994);
xnor UO_1116 (O_1116,N_24807,N_24827);
or UO_1117 (O_1117,N_24851,N_24823);
and UO_1118 (O_1118,N_24810,N_24808);
nor UO_1119 (O_1119,N_24897,N_24951);
or UO_1120 (O_1120,N_24806,N_24888);
nand UO_1121 (O_1121,N_24996,N_24804);
nand UO_1122 (O_1122,N_24973,N_24815);
xor UO_1123 (O_1123,N_24886,N_24855);
or UO_1124 (O_1124,N_24862,N_24836);
and UO_1125 (O_1125,N_24913,N_24884);
nor UO_1126 (O_1126,N_24856,N_24801);
nor UO_1127 (O_1127,N_24814,N_24944);
and UO_1128 (O_1128,N_24985,N_24948);
nor UO_1129 (O_1129,N_24928,N_24814);
nand UO_1130 (O_1130,N_24812,N_24964);
and UO_1131 (O_1131,N_24954,N_24820);
and UO_1132 (O_1132,N_24844,N_24823);
or UO_1133 (O_1133,N_24824,N_24804);
nand UO_1134 (O_1134,N_24936,N_24846);
nand UO_1135 (O_1135,N_24815,N_24958);
or UO_1136 (O_1136,N_24985,N_24940);
or UO_1137 (O_1137,N_24946,N_24839);
or UO_1138 (O_1138,N_24809,N_24854);
and UO_1139 (O_1139,N_24847,N_24903);
or UO_1140 (O_1140,N_24999,N_24804);
nor UO_1141 (O_1141,N_24804,N_24889);
nor UO_1142 (O_1142,N_24936,N_24805);
nor UO_1143 (O_1143,N_24852,N_24805);
xnor UO_1144 (O_1144,N_24994,N_24851);
nand UO_1145 (O_1145,N_24808,N_24857);
xnor UO_1146 (O_1146,N_24977,N_24861);
and UO_1147 (O_1147,N_24871,N_24832);
or UO_1148 (O_1148,N_24982,N_24939);
nor UO_1149 (O_1149,N_24988,N_24997);
or UO_1150 (O_1150,N_24848,N_24813);
and UO_1151 (O_1151,N_24949,N_24932);
nand UO_1152 (O_1152,N_24867,N_24833);
and UO_1153 (O_1153,N_24950,N_24902);
nand UO_1154 (O_1154,N_24857,N_24952);
nor UO_1155 (O_1155,N_24829,N_24900);
and UO_1156 (O_1156,N_24931,N_24853);
nand UO_1157 (O_1157,N_24960,N_24952);
or UO_1158 (O_1158,N_24913,N_24854);
nor UO_1159 (O_1159,N_24914,N_24942);
and UO_1160 (O_1160,N_24868,N_24833);
and UO_1161 (O_1161,N_24886,N_24895);
or UO_1162 (O_1162,N_24988,N_24913);
nand UO_1163 (O_1163,N_24984,N_24908);
nor UO_1164 (O_1164,N_24940,N_24992);
or UO_1165 (O_1165,N_24925,N_24875);
nand UO_1166 (O_1166,N_24944,N_24985);
nor UO_1167 (O_1167,N_24911,N_24812);
and UO_1168 (O_1168,N_24883,N_24955);
xnor UO_1169 (O_1169,N_24867,N_24818);
and UO_1170 (O_1170,N_24972,N_24910);
nor UO_1171 (O_1171,N_24841,N_24884);
nand UO_1172 (O_1172,N_24975,N_24901);
nand UO_1173 (O_1173,N_24962,N_24999);
nor UO_1174 (O_1174,N_24935,N_24914);
and UO_1175 (O_1175,N_24804,N_24967);
and UO_1176 (O_1176,N_24858,N_24919);
nor UO_1177 (O_1177,N_24888,N_24991);
and UO_1178 (O_1178,N_24808,N_24915);
or UO_1179 (O_1179,N_24916,N_24896);
and UO_1180 (O_1180,N_24926,N_24809);
or UO_1181 (O_1181,N_24993,N_24873);
and UO_1182 (O_1182,N_24850,N_24876);
nand UO_1183 (O_1183,N_24807,N_24922);
xor UO_1184 (O_1184,N_24811,N_24941);
nand UO_1185 (O_1185,N_24879,N_24869);
nor UO_1186 (O_1186,N_24817,N_24908);
nand UO_1187 (O_1187,N_24941,N_24904);
and UO_1188 (O_1188,N_24991,N_24878);
or UO_1189 (O_1189,N_24976,N_24821);
nor UO_1190 (O_1190,N_24971,N_24880);
nor UO_1191 (O_1191,N_24939,N_24891);
and UO_1192 (O_1192,N_24912,N_24829);
nand UO_1193 (O_1193,N_24864,N_24801);
nand UO_1194 (O_1194,N_24836,N_24935);
and UO_1195 (O_1195,N_24827,N_24821);
nand UO_1196 (O_1196,N_24905,N_24921);
or UO_1197 (O_1197,N_24954,N_24831);
and UO_1198 (O_1198,N_24903,N_24801);
and UO_1199 (O_1199,N_24998,N_24962);
or UO_1200 (O_1200,N_24896,N_24869);
nor UO_1201 (O_1201,N_24933,N_24941);
and UO_1202 (O_1202,N_24955,N_24818);
and UO_1203 (O_1203,N_24949,N_24831);
nor UO_1204 (O_1204,N_24800,N_24836);
nand UO_1205 (O_1205,N_24884,N_24911);
and UO_1206 (O_1206,N_24803,N_24888);
nand UO_1207 (O_1207,N_24854,N_24899);
or UO_1208 (O_1208,N_24846,N_24972);
and UO_1209 (O_1209,N_24994,N_24902);
nor UO_1210 (O_1210,N_24883,N_24944);
nand UO_1211 (O_1211,N_24882,N_24876);
nor UO_1212 (O_1212,N_24861,N_24831);
or UO_1213 (O_1213,N_24981,N_24986);
nor UO_1214 (O_1214,N_24820,N_24980);
nor UO_1215 (O_1215,N_24896,N_24863);
or UO_1216 (O_1216,N_24814,N_24841);
xor UO_1217 (O_1217,N_24936,N_24896);
nand UO_1218 (O_1218,N_24844,N_24968);
xnor UO_1219 (O_1219,N_24853,N_24907);
nand UO_1220 (O_1220,N_24956,N_24970);
nand UO_1221 (O_1221,N_24888,N_24941);
nand UO_1222 (O_1222,N_24913,N_24870);
nand UO_1223 (O_1223,N_24875,N_24868);
and UO_1224 (O_1224,N_24883,N_24972);
xor UO_1225 (O_1225,N_24919,N_24868);
or UO_1226 (O_1226,N_24888,N_24905);
or UO_1227 (O_1227,N_24911,N_24912);
or UO_1228 (O_1228,N_24806,N_24952);
nand UO_1229 (O_1229,N_24914,N_24919);
nand UO_1230 (O_1230,N_24879,N_24870);
nand UO_1231 (O_1231,N_24915,N_24811);
and UO_1232 (O_1232,N_24997,N_24885);
and UO_1233 (O_1233,N_24900,N_24965);
nor UO_1234 (O_1234,N_24831,N_24870);
nand UO_1235 (O_1235,N_24888,N_24942);
nand UO_1236 (O_1236,N_24912,N_24808);
nand UO_1237 (O_1237,N_24885,N_24909);
or UO_1238 (O_1238,N_24965,N_24989);
xor UO_1239 (O_1239,N_24905,N_24896);
or UO_1240 (O_1240,N_24953,N_24962);
nand UO_1241 (O_1241,N_24885,N_24816);
and UO_1242 (O_1242,N_24975,N_24907);
and UO_1243 (O_1243,N_24888,N_24944);
nor UO_1244 (O_1244,N_24896,N_24947);
or UO_1245 (O_1245,N_24932,N_24862);
nand UO_1246 (O_1246,N_24816,N_24934);
nor UO_1247 (O_1247,N_24832,N_24973);
nand UO_1248 (O_1248,N_24999,N_24856);
nand UO_1249 (O_1249,N_24868,N_24930);
and UO_1250 (O_1250,N_24932,N_24804);
nor UO_1251 (O_1251,N_24848,N_24864);
nor UO_1252 (O_1252,N_24801,N_24982);
nand UO_1253 (O_1253,N_24873,N_24998);
and UO_1254 (O_1254,N_24859,N_24870);
and UO_1255 (O_1255,N_24982,N_24902);
and UO_1256 (O_1256,N_24902,N_24949);
or UO_1257 (O_1257,N_24964,N_24914);
and UO_1258 (O_1258,N_24984,N_24962);
or UO_1259 (O_1259,N_24846,N_24908);
nor UO_1260 (O_1260,N_24816,N_24806);
or UO_1261 (O_1261,N_24875,N_24866);
nor UO_1262 (O_1262,N_24926,N_24839);
nand UO_1263 (O_1263,N_24856,N_24869);
xnor UO_1264 (O_1264,N_24958,N_24967);
or UO_1265 (O_1265,N_24919,N_24888);
and UO_1266 (O_1266,N_24904,N_24901);
or UO_1267 (O_1267,N_24842,N_24923);
nand UO_1268 (O_1268,N_24829,N_24850);
or UO_1269 (O_1269,N_24864,N_24953);
and UO_1270 (O_1270,N_24956,N_24987);
and UO_1271 (O_1271,N_24808,N_24957);
or UO_1272 (O_1272,N_24836,N_24915);
and UO_1273 (O_1273,N_24882,N_24931);
and UO_1274 (O_1274,N_24994,N_24815);
nand UO_1275 (O_1275,N_24934,N_24818);
nor UO_1276 (O_1276,N_24934,N_24998);
nand UO_1277 (O_1277,N_24959,N_24993);
and UO_1278 (O_1278,N_24833,N_24990);
nor UO_1279 (O_1279,N_24890,N_24901);
and UO_1280 (O_1280,N_24910,N_24915);
or UO_1281 (O_1281,N_24811,N_24855);
and UO_1282 (O_1282,N_24858,N_24932);
xor UO_1283 (O_1283,N_24956,N_24981);
and UO_1284 (O_1284,N_24901,N_24940);
nor UO_1285 (O_1285,N_24824,N_24829);
nor UO_1286 (O_1286,N_24801,N_24846);
nand UO_1287 (O_1287,N_24830,N_24820);
nor UO_1288 (O_1288,N_24804,N_24963);
xnor UO_1289 (O_1289,N_24843,N_24907);
nand UO_1290 (O_1290,N_24928,N_24846);
xnor UO_1291 (O_1291,N_24942,N_24979);
or UO_1292 (O_1292,N_24948,N_24904);
or UO_1293 (O_1293,N_24988,N_24971);
or UO_1294 (O_1294,N_24979,N_24946);
nand UO_1295 (O_1295,N_24994,N_24842);
nand UO_1296 (O_1296,N_24857,N_24914);
or UO_1297 (O_1297,N_24962,N_24841);
nand UO_1298 (O_1298,N_24969,N_24839);
nand UO_1299 (O_1299,N_24989,N_24949);
and UO_1300 (O_1300,N_24971,N_24828);
xnor UO_1301 (O_1301,N_24974,N_24980);
nand UO_1302 (O_1302,N_24862,N_24914);
nor UO_1303 (O_1303,N_24980,N_24848);
nand UO_1304 (O_1304,N_24850,N_24804);
or UO_1305 (O_1305,N_24935,N_24885);
xor UO_1306 (O_1306,N_24804,N_24917);
xnor UO_1307 (O_1307,N_24853,N_24824);
xnor UO_1308 (O_1308,N_24999,N_24928);
and UO_1309 (O_1309,N_24953,N_24876);
and UO_1310 (O_1310,N_24878,N_24962);
xor UO_1311 (O_1311,N_24966,N_24928);
nand UO_1312 (O_1312,N_24951,N_24891);
nand UO_1313 (O_1313,N_24911,N_24951);
or UO_1314 (O_1314,N_24919,N_24971);
and UO_1315 (O_1315,N_24921,N_24977);
nand UO_1316 (O_1316,N_24977,N_24887);
or UO_1317 (O_1317,N_24920,N_24956);
nor UO_1318 (O_1318,N_24877,N_24921);
xnor UO_1319 (O_1319,N_24889,N_24965);
and UO_1320 (O_1320,N_24857,N_24942);
nand UO_1321 (O_1321,N_24937,N_24941);
or UO_1322 (O_1322,N_24969,N_24826);
or UO_1323 (O_1323,N_24932,N_24810);
or UO_1324 (O_1324,N_24825,N_24961);
xnor UO_1325 (O_1325,N_24944,N_24871);
nor UO_1326 (O_1326,N_24972,N_24966);
or UO_1327 (O_1327,N_24864,N_24999);
xnor UO_1328 (O_1328,N_24968,N_24993);
or UO_1329 (O_1329,N_24948,N_24970);
and UO_1330 (O_1330,N_24963,N_24846);
and UO_1331 (O_1331,N_24893,N_24902);
xor UO_1332 (O_1332,N_24802,N_24836);
or UO_1333 (O_1333,N_24956,N_24986);
and UO_1334 (O_1334,N_24977,N_24845);
nor UO_1335 (O_1335,N_24948,N_24876);
xnor UO_1336 (O_1336,N_24903,N_24815);
nor UO_1337 (O_1337,N_24915,N_24846);
or UO_1338 (O_1338,N_24964,N_24919);
and UO_1339 (O_1339,N_24846,N_24953);
xor UO_1340 (O_1340,N_24978,N_24926);
nand UO_1341 (O_1341,N_24862,N_24889);
and UO_1342 (O_1342,N_24821,N_24802);
or UO_1343 (O_1343,N_24843,N_24840);
or UO_1344 (O_1344,N_24917,N_24911);
nand UO_1345 (O_1345,N_24866,N_24893);
nor UO_1346 (O_1346,N_24863,N_24883);
xnor UO_1347 (O_1347,N_24868,N_24992);
or UO_1348 (O_1348,N_24893,N_24890);
nand UO_1349 (O_1349,N_24807,N_24811);
or UO_1350 (O_1350,N_24836,N_24969);
nand UO_1351 (O_1351,N_24972,N_24847);
nor UO_1352 (O_1352,N_24872,N_24853);
nor UO_1353 (O_1353,N_24800,N_24966);
nand UO_1354 (O_1354,N_24844,N_24971);
and UO_1355 (O_1355,N_24934,N_24992);
nand UO_1356 (O_1356,N_24937,N_24923);
and UO_1357 (O_1357,N_24863,N_24998);
or UO_1358 (O_1358,N_24976,N_24979);
and UO_1359 (O_1359,N_24824,N_24993);
nand UO_1360 (O_1360,N_24865,N_24940);
nand UO_1361 (O_1361,N_24952,N_24966);
nor UO_1362 (O_1362,N_24989,N_24843);
and UO_1363 (O_1363,N_24869,N_24913);
and UO_1364 (O_1364,N_24823,N_24978);
and UO_1365 (O_1365,N_24851,N_24860);
or UO_1366 (O_1366,N_24919,N_24805);
nand UO_1367 (O_1367,N_24940,N_24981);
and UO_1368 (O_1368,N_24835,N_24914);
xnor UO_1369 (O_1369,N_24891,N_24957);
and UO_1370 (O_1370,N_24836,N_24840);
or UO_1371 (O_1371,N_24859,N_24851);
xnor UO_1372 (O_1372,N_24885,N_24803);
and UO_1373 (O_1373,N_24888,N_24945);
xnor UO_1374 (O_1374,N_24810,N_24807);
or UO_1375 (O_1375,N_24826,N_24828);
and UO_1376 (O_1376,N_24937,N_24829);
and UO_1377 (O_1377,N_24805,N_24875);
nand UO_1378 (O_1378,N_24967,N_24978);
or UO_1379 (O_1379,N_24899,N_24866);
nor UO_1380 (O_1380,N_24990,N_24815);
and UO_1381 (O_1381,N_24933,N_24838);
nand UO_1382 (O_1382,N_24816,N_24970);
nor UO_1383 (O_1383,N_24855,N_24958);
xnor UO_1384 (O_1384,N_24869,N_24883);
nor UO_1385 (O_1385,N_24819,N_24907);
nand UO_1386 (O_1386,N_24865,N_24806);
nor UO_1387 (O_1387,N_24895,N_24962);
and UO_1388 (O_1388,N_24970,N_24875);
nand UO_1389 (O_1389,N_24955,N_24807);
nor UO_1390 (O_1390,N_24942,N_24818);
nor UO_1391 (O_1391,N_24890,N_24811);
nand UO_1392 (O_1392,N_24849,N_24895);
nor UO_1393 (O_1393,N_24963,N_24897);
or UO_1394 (O_1394,N_24941,N_24964);
and UO_1395 (O_1395,N_24868,N_24881);
nor UO_1396 (O_1396,N_24801,N_24867);
nand UO_1397 (O_1397,N_24907,N_24820);
or UO_1398 (O_1398,N_24876,N_24944);
nor UO_1399 (O_1399,N_24926,N_24838);
or UO_1400 (O_1400,N_24984,N_24897);
nand UO_1401 (O_1401,N_24934,N_24953);
nor UO_1402 (O_1402,N_24982,N_24884);
nor UO_1403 (O_1403,N_24891,N_24967);
and UO_1404 (O_1404,N_24971,N_24817);
nand UO_1405 (O_1405,N_24866,N_24840);
or UO_1406 (O_1406,N_24808,N_24932);
or UO_1407 (O_1407,N_24987,N_24932);
xor UO_1408 (O_1408,N_24821,N_24903);
nor UO_1409 (O_1409,N_24934,N_24984);
or UO_1410 (O_1410,N_24904,N_24923);
xor UO_1411 (O_1411,N_24933,N_24825);
and UO_1412 (O_1412,N_24811,N_24884);
xor UO_1413 (O_1413,N_24964,N_24974);
and UO_1414 (O_1414,N_24928,N_24969);
nand UO_1415 (O_1415,N_24825,N_24829);
or UO_1416 (O_1416,N_24983,N_24890);
and UO_1417 (O_1417,N_24944,N_24915);
or UO_1418 (O_1418,N_24949,N_24845);
nand UO_1419 (O_1419,N_24813,N_24911);
nor UO_1420 (O_1420,N_24802,N_24955);
xnor UO_1421 (O_1421,N_24867,N_24956);
nand UO_1422 (O_1422,N_24926,N_24963);
and UO_1423 (O_1423,N_24937,N_24980);
nand UO_1424 (O_1424,N_24953,N_24986);
xnor UO_1425 (O_1425,N_24816,N_24990);
and UO_1426 (O_1426,N_24853,N_24908);
nor UO_1427 (O_1427,N_24959,N_24931);
and UO_1428 (O_1428,N_24958,N_24804);
xor UO_1429 (O_1429,N_24885,N_24919);
nor UO_1430 (O_1430,N_24903,N_24851);
xnor UO_1431 (O_1431,N_24928,N_24954);
nand UO_1432 (O_1432,N_24849,N_24930);
nand UO_1433 (O_1433,N_24839,N_24994);
nand UO_1434 (O_1434,N_24874,N_24992);
nand UO_1435 (O_1435,N_24942,N_24931);
or UO_1436 (O_1436,N_24918,N_24890);
nand UO_1437 (O_1437,N_24812,N_24969);
and UO_1438 (O_1438,N_24909,N_24972);
or UO_1439 (O_1439,N_24989,N_24922);
or UO_1440 (O_1440,N_24828,N_24825);
nand UO_1441 (O_1441,N_24956,N_24808);
nand UO_1442 (O_1442,N_24837,N_24891);
and UO_1443 (O_1443,N_24942,N_24814);
or UO_1444 (O_1444,N_24811,N_24817);
and UO_1445 (O_1445,N_24949,N_24870);
nor UO_1446 (O_1446,N_24881,N_24962);
and UO_1447 (O_1447,N_24985,N_24971);
nand UO_1448 (O_1448,N_24978,N_24977);
nor UO_1449 (O_1449,N_24929,N_24994);
and UO_1450 (O_1450,N_24997,N_24986);
or UO_1451 (O_1451,N_24994,N_24940);
and UO_1452 (O_1452,N_24832,N_24861);
or UO_1453 (O_1453,N_24829,N_24916);
nor UO_1454 (O_1454,N_24981,N_24854);
nand UO_1455 (O_1455,N_24986,N_24889);
or UO_1456 (O_1456,N_24999,N_24959);
or UO_1457 (O_1457,N_24826,N_24945);
nor UO_1458 (O_1458,N_24971,N_24994);
and UO_1459 (O_1459,N_24962,N_24910);
and UO_1460 (O_1460,N_24899,N_24801);
and UO_1461 (O_1461,N_24834,N_24835);
nor UO_1462 (O_1462,N_24932,N_24844);
or UO_1463 (O_1463,N_24910,N_24877);
nor UO_1464 (O_1464,N_24881,N_24913);
nand UO_1465 (O_1465,N_24935,N_24889);
and UO_1466 (O_1466,N_24871,N_24813);
nor UO_1467 (O_1467,N_24811,N_24887);
and UO_1468 (O_1468,N_24928,N_24919);
and UO_1469 (O_1469,N_24955,N_24953);
nor UO_1470 (O_1470,N_24893,N_24825);
and UO_1471 (O_1471,N_24925,N_24828);
and UO_1472 (O_1472,N_24993,N_24909);
and UO_1473 (O_1473,N_24913,N_24929);
or UO_1474 (O_1474,N_24871,N_24851);
and UO_1475 (O_1475,N_24970,N_24813);
and UO_1476 (O_1476,N_24902,N_24941);
and UO_1477 (O_1477,N_24991,N_24985);
nor UO_1478 (O_1478,N_24970,N_24929);
xnor UO_1479 (O_1479,N_24847,N_24845);
nor UO_1480 (O_1480,N_24896,N_24955);
and UO_1481 (O_1481,N_24841,N_24917);
nand UO_1482 (O_1482,N_24859,N_24978);
or UO_1483 (O_1483,N_24944,N_24890);
or UO_1484 (O_1484,N_24985,N_24915);
or UO_1485 (O_1485,N_24941,N_24855);
and UO_1486 (O_1486,N_24810,N_24927);
or UO_1487 (O_1487,N_24869,N_24923);
nand UO_1488 (O_1488,N_24833,N_24906);
nor UO_1489 (O_1489,N_24877,N_24802);
nand UO_1490 (O_1490,N_24847,N_24975);
and UO_1491 (O_1491,N_24904,N_24967);
nand UO_1492 (O_1492,N_24954,N_24978);
nand UO_1493 (O_1493,N_24972,N_24893);
nand UO_1494 (O_1494,N_24868,N_24812);
xor UO_1495 (O_1495,N_24925,N_24893);
xor UO_1496 (O_1496,N_24896,N_24805);
nor UO_1497 (O_1497,N_24823,N_24856);
nor UO_1498 (O_1498,N_24975,N_24996);
and UO_1499 (O_1499,N_24929,N_24871);
or UO_1500 (O_1500,N_24840,N_24934);
and UO_1501 (O_1501,N_24892,N_24978);
or UO_1502 (O_1502,N_24827,N_24915);
or UO_1503 (O_1503,N_24829,N_24981);
nor UO_1504 (O_1504,N_24818,N_24953);
or UO_1505 (O_1505,N_24822,N_24929);
xor UO_1506 (O_1506,N_24880,N_24873);
nor UO_1507 (O_1507,N_24855,N_24808);
nand UO_1508 (O_1508,N_24897,N_24925);
and UO_1509 (O_1509,N_24836,N_24865);
and UO_1510 (O_1510,N_24966,N_24890);
nand UO_1511 (O_1511,N_24974,N_24884);
or UO_1512 (O_1512,N_24937,N_24914);
nor UO_1513 (O_1513,N_24961,N_24991);
nor UO_1514 (O_1514,N_24894,N_24949);
nor UO_1515 (O_1515,N_24910,N_24922);
nor UO_1516 (O_1516,N_24816,N_24843);
and UO_1517 (O_1517,N_24950,N_24830);
nor UO_1518 (O_1518,N_24806,N_24956);
or UO_1519 (O_1519,N_24828,N_24822);
nor UO_1520 (O_1520,N_24975,N_24935);
or UO_1521 (O_1521,N_24850,N_24803);
or UO_1522 (O_1522,N_24998,N_24979);
nand UO_1523 (O_1523,N_24827,N_24826);
nand UO_1524 (O_1524,N_24896,N_24850);
nand UO_1525 (O_1525,N_24879,N_24823);
nand UO_1526 (O_1526,N_24873,N_24818);
or UO_1527 (O_1527,N_24916,N_24900);
nand UO_1528 (O_1528,N_24940,N_24966);
nand UO_1529 (O_1529,N_24870,N_24977);
and UO_1530 (O_1530,N_24850,N_24834);
nor UO_1531 (O_1531,N_24959,N_24884);
nor UO_1532 (O_1532,N_24955,N_24987);
nor UO_1533 (O_1533,N_24994,N_24908);
and UO_1534 (O_1534,N_24808,N_24964);
nor UO_1535 (O_1535,N_24985,N_24907);
nand UO_1536 (O_1536,N_24895,N_24903);
xnor UO_1537 (O_1537,N_24846,N_24914);
nor UO_1538 (O_1538,N_24982,N_24865);
nor UO_1539 (O_1539,N_24898,N_24949);
nand UO_1540 (O_1540,N_24930,N_24945);
nor UO_1541 (O_1541,N_24927,N_24890);
nor UO_1542 (O_1542,N_24883,N_24873);
xnor UO_1543 (O_1543,N_24845,N_24959);
nand UO_1544 (O_1544,N_24916,N_24831);
nand UO_1545 (O_1545,N_24902,N_24869);
and UO_1546 (O_1546,N_24956,N_24949);
nor UO_1547 (O_1547,N_24844,N_24803);
nand UO_1548 (O_1548,N_24901,N_24873);
and UO_1549 (O_1549,N_24899,N_24851);
nor UO_1550 (O_1550,N_24805,N_24808);
or UO_1551 (O_1551,N_24836,N_24867);
xor UO_1552 (O_1552,N_24922,N_24872);
or UO_1553 (O_1553,N_24936,N_24960);
nor UO_1554 (O_1554,N_24933,N_24857);
and UO_1555 (O_1555,N_24928,N_24806);
nor UO_1556 (O_1556,N_24912,N_24863);
and UO_1557 (O_1557,N_24843,N_24909);
or UO_1558 (O_1558,N_24832,N_24976);
nand UO_1559 (O_1559,N_24827,N_24860);
nor UO_1560 (O_1560,N_24965,N_24986);
nand UO_1561 (O_1561,N_24905,N_24964);
and UO_1562 (O_1562,N_24802,N_24890);
and UO_1563 (O_1563,N_24999,N_24802);
and UO_1564 (O_1564,N_24975,N_24881);
nor UO_1565 (O_1565,N_24960,N_24992);
nand UO_1566 (O_1566,N_24998,N_24930);
or UO_1567 (O_1567,N_24899,N_24808);
or UO_1568 (O_1568,N_24975,N_24887);
nand UO_1569 (O_1569,N_24995,N_24990);
nor UO_1570 (O_1570,N_24993,N_24826);
xnor UO_1571 (O_1571,N_24855,N_24881);
or UO_1572 (O_1572,N_24824,N_24814);
and UO_1573 (O_1573,N_24923,N_24847);
nor UO_1574 (O_1574,N_24885,N_24801);
and UO_1575 (O_1575,N_24994,N_24979);
and UO_1576 (O_1576,N_24940,N_24801);
and UO_1577 (O_1577,N_24941,N_24827);
or UO_1578 (O_1578,N_24857,N_24851);
nor UO_1579 (O_1579,N_24866,N_24941);
nor UO_1580 (O_1580,N_24853,N_24929);
or UO_1581 (O_1581,N_24910,N_24992);
nor UO_1582 (O_1582,N_24857,N_24935);
nand UO_1583 (O_1583,N_24867,N_24846);
or UO_1584 (O_1584,N_24835,N_24851);
xor UO_1585 (O_1585,N_24910,N_24822);
and UO_1586 (O_1586,N_24950,N_24998);
and UO_1587 (O_1587,N_24877,N_24899);
nand UO_1588 (O_1588,N_24812,N_24816);
nor UO_1589 (O_1589,N_24800,N_24906);
xor UO_1590 (O_1590,N_24930,N_24829);
or UO_1591 (O_1591,N_24942,N_24993);
and UO_1592 (O_1592,N_24829,N_24951);
nor UO_1593 (O_1593,N_24904,N_24946);
nor UO_1594 (O_1594,N_24828,N_24975);
or UO_1595 (O_1595,N_24866,N_24825);
nand UO_1596 (O_1596,N_24975,N_24879);
nor UO_1597 (O_1597,N_24899,N_24936);
nand UO_1598 (O_1598,N_24962,N_24877);
nor UO_1599 (O_1599,N_24837,N_24992);
nand UO_1600 (O_1600,N_24984,N_24848);
nor UO_1601 (O_1601,N_24997,N_24817);
and UO_1602 (O_1602,N_24812,N_24914);
nand UO_1603 (O_1603,N_24932,N_24888);
nor UO_1604 (O_1604,N_24854,N_24820);
nand UO_1605 (O_1605,N_24920,N_24815);
or UO_1606 (O_1606,N_24953,N_24897);
nor UO_1607 (O_1607,N_24946,N_24828);
xnor UO_1608 (O_1608,N_24894,N_24884);
nor UO_1609 (O_1609,N_24977,N_24834);
nor UO_1610 (O_1610,N_24951,N_24993);
and UO_1611 (O_1611,N_24941,N_24833);
or UO_1612 (O_1612,N_24850,N_24821);
nor UO_1613 (O_1613,N_24940,N_24960);
nand UO_1614 (O_1614,N_24824,N_24937);
nand UO_1615 (O_1615,N_24803,N_24810);
and UO_1616 (O_1616,N_24808,N_24907);
nand UO_1617 (O_1617,N_24887,N_24956);
or UO_1618 (O_1618,N_24854,N_24822);
or UO_1619 (O_1619,N_24942,N_24858);
or UO_1620 (O_1620,N_24838,N_24950);
nor UO_1621 (O_1621,N_24921,N_24817);
xnor UO_1622 (O_1622,N_24895,N_24885);
nand UO_1623 (O_1623,N_24955,N_24806);
and UO_1624 (O_1624,N_24928,N_24997);
xnor UO_1625 (O_1625,N_24894,N_24930);
nor UO_1626 (O_1626,N_24814,N_24816);
xor UO_1627 (O_1627,N_24886,N_24823);
nand UO_1628 (O_1628,N_24987,N_24870);
nor UO_1629 (O_1629,N_24812,N_24943);
nor UO_1630 (O_1630,N_24821,N_24811);
nor UO_1631 (O_1631,N_24918,N_24822);
or UO_1632 (O_1632,N_24939,N_24805);
or UO_1633 (O_1633,N_24823,N_24869);
nand UO_1634 (O_1634,N_24826,N_24984);
xor UO_1635 (O_1635,N_24806,N_24880);
xor UO_1636 (O_1636,N_24909,N_24812);
xnor UO_1637 (O_1637,N_24872,N_24849);
nor UO_1638 (O_1638,N_24916,N_24832);
or UO_1639 (O_1639,N_24933,N_24822);
nand UO_1640 (O_1640,N_24877,N_24829);
nor UO_1641 (O_1641,N_24946,N_24920);
nor UO_1642 (O_1642,N_24994,N_24945);
nor UO_1643 (O_1643,N_24889,N_24857);
or UO_1644 (O_1644,N_24848,N_24807);
nor UO_1645 (O_1645,N_24845,N_24965);
or UO_1646 (O_1646,N_24891,N_24993);
and UO_1647 (O_1647,N_24953,N_24928);
xor UO_1648 (O_1648,N_24800,N_24997);
or UO_1649 (O_1649,N_24823,N_24958);
nor UO_1650 (O_1650,N_24868,N_24894);
nand UO_1651 (O_1651,N_24878,N_24929);
and UO_1652 (O_1652,N_24933,N_24815);
or UO_1653 (O_1653,N_24804,N_24811);
nand UO_1654 (O_1654,N_24857,N_24896);
and UO_1655 (O_1655,N_24828,N_24805);
nand UO_1656 (O_1656,N_24815,N_24800);
and UO_1657 (O_1657,N_24802,N_24813);
nand UO_1658 (O_1658,N_24972,N_24806);
or UO_1659 (O_1659,N_24851,N_24980);
and UO_1660 (O_1660,N_24943,N_24903);
nor UO_1661 (O_1661,N_24902,N_24843);
and UO_1662 (O_1662,N_24873,N_24872);
nor UO_1663 (O_1663,N_24809,N_24890);
and UO_1664 (O_1664,N_24928,N_24911);
or UO_1665 (O_1665,N_24834,N_24940);
or UO_1666 (O_1666,N_24831,N_24806);
nor UO_1667 (O_1667,N_24992,N_24844);
nor UO_1668 (O_1668,N_24959,N_24928);
or UO_1669 (O_1669,N_24867,N_24811);
nor UO_1670 (O_1670,N_24910,N_24987);
nor UO_1671 (O_1671,N_24970,N_24851);
and UO_1672 (O_1672,N_24915,N_24992);
or UO_1673 (O_1673,N_24878,N_24982);
and UO_1674 (O_1674,N_24803,N_24895);
or UO_1675 (O_1675,N_24901,N_24910);
or UO_1676 (O_1676,N_24881,N_24890);
or UO_1677 (O_1677,N_24961,N_24976);
nand UO_1678 (O_1678,N_24866,N_24937);
nand UO_1679 (O_1679,N_24983,N_24989);
nor UO_1680 (O_1680,N_24948,N_24925);
nor UO_1681 (O_1681,N_24822,N_24970);
nand UO_1682 (O_1682,N_24948,N_24827);
and UO_1683 (O_1683,N_24975,N_24855);
nor UO_1684 (O_1684,N_24828,N_24923);
nor UO_1685 (O_1685,N_24938,N_24946);
and UO_1686 (O_1686,N_24962,N_24902);
and UO_1687 (O_1687,N_24848,N_24978);
nand UO_1688 (O_1688,N_24974,N_24969);
and UO_1689 (O_1689,N_24944,N_24897);
and UO_1690 (O_1690,N_24946,N_24863);
and UO_1691 (O_1691,N_24896,N_24831);
nor UO_1692 (O_1692,N_24975,N_24836);
xnor UO_1693 (O_1693,N_24804,N_24928);
nor UO_1694 (O_1694,N_24889,N_24983);
or UO_1695 (O_1695,N_24847,N_24834);
nand UO_1696 (O_1696,N_24834,N_24857);
or UO_1697 (O_1697,N_24866,N_24946);
and UO_1698 (O_1698,N_24829,N_24865);
nor UO_1699 (O_1699,N_24841,N_24922);
and UO_1700 (O_1700,N_24903,N_24942);
or UO_1701 (O_1701,N_24896,N_24929);
and UO_1702 (O_1702,N_24919,N_24980);
nor UO_1703 (O_1703,N_24994,N_24933);
nor UO_1704 (O_1704,N_24901,N_24825);
nor UO_1705 (O_1705,N_24971,N_24979);
nand UO_1706 (O_1706,N_24838,N_24847);
or UO_1707 (O_1707,N_24996,N_24862);
and UO_1708 (O_1708,N_24987,N_24953);
nand UO_1709 (O_1709,N_24823,N_24861);
and UO_1710 (O_1710,N_24890,N_24908);
nand UO_1711 (O_1711,N_24972,N_24985);
nand UO_1712 (O_1712,N_24974,N_24910);
or UO_1713 (O_1713,N_24800,N_24851);
nor UO_1714 (O_1714,N_24929,N_24905);
or UO_1715 (O_1715,N_24904,N_24894);
nand UO_1716 (O_1716,N_24813,N_24930);
and UO_1717 (O_1717,N_24968,N_24898);
and UO_1718 (O_1718,N_24971,N_24809);
and UO_1719 (O_1719,N_24808,N_24927);
or UO_1720 (O_1720,N_24864,N_24986);
or UO_1721 (O_1721,N_24970,N_24988);
nand UO_1722 (O_1722,N_24801,N_24879);
or UO_1723 (O_1723,N_24871,N_24907);
and UO_1724 (O_1724,N_24916,N_24915);
nand UO_1725 (O_1725,N_24831,N_24812);
nor UO_1726 (O_1726,N_24943,N_24843);
nor UO_1727 (O_1727,N_24865,N_24883);
nor UO_1728 (O_1728,N_24817,N_24944);
nand UO_1729 (O_1729,N_24810,N_24948);
and UO_1730 (O_1730,N_24939,N_24867);
nand UO_1731 (O_1731,N_24946,N_24872);
and UO_1732 (O_1732,N_24928,N_24924);
xnor UO_1733 (O_1733,N_24852,N_24946);
or UO_1734 (O_1734,N_24914,N_24948);
nand UO_1735 (O_1735,N_24928,N_24818);
nor UO_1736 (O_1736,N_24976,N_24934);
xor UO_1737 (O_1737,N_24948,N_24995);
and UO_1738 (O_1738,N_24958,N_24838);
xor UO_1739 (O_1739,N_24917,N_24808);
or UO_1740 (O_1740,N_24807,N_24833);
nand UO_1741 (O_1741,N_24882,N_24994);
nand UO_1742 (O_1742,N_24955,N_24856);
nor UO_1743 (O_1743,N_24935,N_24999);
and UO_1744 (O_1744,N_24962,N_24909);
or UO_1745 (O_1745,N_24953,N_24957);
and UO_1746 (O_1746,N_24813,N_24915);
nor UO_1747 (O_1747,N_24835,N_24846);
and UO_1748 (O_1748,N_24861,N_24835);
or UO_1749 (O_1749,N_24827,N_24991);
or UO_1750 (O_1750,N_24991,N_24875);
nand UO_1751 (O_1751,N_24865,N_24931);
or UO_1752 (O_1752,N_24895,N_24975);
nand UO_1753 (O_1753,N_24851,N_24909);
or UO_1754 (O_1754,N_24819,N_24941);
nand UO_1755 (O_1755,N_24838,N_24898);
or UO_1756 (O_1756,N_24862,N_24827);
and UO_1757 (O_1757,N_24824,N_24883);
and UO_1758 (O_1758,N_24929,N_24982);
and UO_1759 (O_1759,N_24865,N_24934);
nor UO_1760 (O_1760,N_24963,N_24889);
and UO_1761 (O_1761,N_24907,N_24939);
xnor UO_1762 (O_1762,N_24923,N_24866);
and UO_1763 (O_1763,N_24917,N_24988);
and UO_1764 (O_1764,N_24880,N_24996);
and UO_1765 (O_1765,N_24861,N_24888);
nand UO_1766 (O_1766,N_24914,N_24905);
nor UO_1767 (O_1767,N_24924,N_24913);
nand UO_1768 (O_1768,N_24830,N_24833);
or UO_1769 (O_1769,N_24900,N_24912);
and UO_1770 (O_1770,N_24964,N_24988);
nand UO_1771 (O_1771,N_24999,N_24868);
or UO_1772 (O_1772,N_24998,N_24981);
nand UO_1773 (O_1773,N_24986,N_24840);
and UO_1774 (O_1774,N_24824,N_24991);
and UO_1775 (O_1775,N_24825,N_24998);
and UO_1776 (O_1776,N_24908,N_24866);
nand UO_1777 (O_1777,N_24818,N_24876);
xnor UO_1778 (O_1778,N_24852,N_24887);
xnor UO_1779 (O_1779,N_24861,N_24871);
xnor UO_1780 (O_1780,N_24823,N_24876);
nand UO_1781 (O_1781,N_24833,N_24865);
and UO_1782 (O_1782,N_24833,N_24958);
nor UO_1783 (O_1783,N_24902,N_24837);
nor UO_1784 (O_1784,N_24915,N_24893);
xor UO_1785 (O_1785,N_24959,N_24966);
or UO_1786 (O_1786,N_24803,N_24859);
or UO_1787 (O_1787,N_24885,N_24805);
or UO_1788 (O_1788,N_24868,N_24899);
nand UO_1789 (O_1789,N_24931,N_24909);
nand UO_1790 (O_1790,N_24883,N_24807);
and UO_1791 (O_1791,N_24828,N_24881);
or UO_1792 (O_1792,N_24985,N_24883);
or UO_1793 (O_1793,N_24947,N_24893);
or UO_1794 (O_1794,N_24846,N_24916);
or UO_1795 (O_1795,N_24902,N_24825);
nand UO_1796 (O_1796,N_24959,N_24957);
nand UO_1797 (O_1797,N_24852,N_24808);
nand UO_1798 (O_1798,N_24871,N_24917);
and UO_1799 (O_1799,N_24980,N_24866);
nand UO_1800 (O_1800,N_24859,N_24943);
and UO_1801 (O_1801,N_24963,N_24911);
xnor UO_1802 (O_1802,N_24999,N_24878);
xnor UO_1803 (O_1803,N_24809,N_24984);
and UO_1804 (O_1804,N_24995,N_24903);
or UO_1805 (O_1805,N_24816,N_24813);
or UO_1806 (O_1806,N_24926,N_24816);
nor UO_1807 (O_1807,N_24975,N_24883);
or UO_1808 (O_1808,N_24894,N_24861);
and UO_1809 (O_1809,N_24829,N_24863);
or UO_1810 (O_1810,N_24916,N_24840);
or UO_1811 (O_1811,N_24899,N_24940);
nor UO_1812 (O_1812,N_24978,N_24918);
and UO_1813 (O_1813,N_24815,N_24959);
and UO_1814 (O_1814,N_24871,N_24987);
nand UO_1815 (O_1815,N_24925,N_24979);
nand UO_1816 (O_1816,N_24968,N_24862);
nor UO_1817 (O_1817,N_24960,N_24877);
and UO_1818 (O_1818,N_24989,N_24918);
or UO_1819 (O_1819,N_24811,N_24978);
and UO_1820 (O_1820,N_24911,N_24819);
nand UO_1821 (O_1821,N_24896,N_24963);
or UO_1822 (O_1822,N_24900,N_24923);
or UO_1823 (O_1823,N_24985,N_24874);
and UO_1824 (O_1824,N_24964,N_24997);
and UO_1825 (O_1825,N_24930,N_24933);
nor UO_1826 (O_1826,N_24907,N_24895);
and UO_1827 (O_1827,N_24975,N_24889);
and UO_1828 (O_1828,N_24836,N_24913);
and UO_1829 (O_1829,N_24908,N_24878);
nand UO_1830 (O_1830,N_24840,N_24817);
nand UO_1831 (O_1831,N_24809,N_24931);
nor UO_1832 (O_1832,N_24972,N_24961);
or UO_1833 (O_1833,N_24973,N_24839);
and UO_1834 (O_1834,N_24891,N_24838);
or UO_1835 (O_1835,N_24948,N_24920);
and UO_1836 (O_1836,N_24895,N_24833);
or UO_1837 (O_1837,N_24824,N_24983);
or UO_1838 (O_1838,N_24966,N_24945);
nor UO_1839 (O_1839,N_24927,N_24978);
and UO_1840 (O_1840,N_24949,N_24995);
and UO_1841 (O_1841,N_24803,N_24987);
or UO_1842 (O_1842,N_24971,N_24929);
nand UO_1843 (O_1843,N_24887,N_24869);
and UO_1844 (O_1844,N_24896,N_24941);
nor UO_1845 (O_1845,N_24975,N_24813);
xnor UO_1846 (O_1846,N_24811,N_24826);
nor UO_1847 (O_1847,N_24910,N_24969);
or UO_1848 (O_1848,N_24818,N_24979);
nor UO_1849 (O_1849,N_24880,N_24861);
and UO_1850 (O_1850,N_24996,N_24937);
or UO_1851 (O_1851,N_24848,N_24972);
nand UO_1852 (O_1852,N_24863,N_24973);
nand UO_1853 (O_1853,N_24999,N_24821);
nand UO_1854 (O_1854,N_24947,N_24874);
nand UO_1855 (O_1855,N_24834,N_24805);
or UO_1856 (O_1856,N_24890,N_24952);
or UO_1857 (O_1857,N_24989,N_24984);
xnor UO_1858 (O_1858,N_24914,N_24989);
nand UO_1859 (O_1859,N_24929,N_24902);
or UO_1860 (O_1860,N_24963,N_24981);
and UO_1861 (O_1861,N_24972,N_24878);
nand UO_1862 (O_1862,N_24930,N_24962);
xnor UO_1863 (O_1863,N_24956,N_24964);
nor UO_1864 (O_1864,N_24911,N_24956);
or UO_1865 (O_1865,N_24976,N_24841);
nor UO_1866 (O_1866,N_24954,N_24860);
nor UO_1867 (O_1867,N_24810,N_24917);
nor UO_1868 (O_1868,N_24862,N_24933);
and UO_1869 (O_1869,N_24830,N_24963);
xnor UO_1870 (O_1870,N_24895,N_24860);
and UO_1871 (O_1871,N_24981,N_24833);
and UO_1872 (O_1872,N_24975,N_24923);
xor UO_1873 (O_1873,N_24845,N_24988);
nand UO_1874 (O_1874,N_24985,N_24916);
nand UO_1875 (O_1875,N_24950,N_24992);
and UO_1876 (O_1876,N_24857,N_24825);
and UO_1877 (O_1877,N_24952,N_24899);
or UO_1878 (O_1878,N_24816,N_24951);
nand UO_1879 (O_1879,N_24933,N_24889);
and UO_1880 (O_1880,N_24990,N_24848);
or UO_1881 (O_1881,N_24902,N_24812);
or UO_1882 (O_1882,N_24881,N_24991);
nor UO_1883 (O_1883,N_24985,N_24953);
nor UO_1884 (O_1884,N_24892,N_24972);
and UO_1885 (O_1885,N_24881,N_24902);
nand UO_1886 (O_1886,N_24981,N_24958);
and UO_1887 (O_1887,N_24977,N_24994);
and UO_1888 (O_1888,N_24865,N_24813);
nand UO_1889 (O_1889,N_24842,N_24802);
nor UO_1890 (O_1890,N_24950,N_24808);
nand UO_1891 (O_1891,N_24897,N_24891);
or UO_1892 (O_1892,N_24919,N_24838);
nor UO_1893 (O_1893,N_24989,N_24892);
nor UO_1894 (O_1894,N_24862,N_24831);
or UO_1895 (O_1895,N_24999,N_24974);
nand UO_1896 (O_1896,N_24993,N_24965);
nand UO_1897 (O_1897,N_24948,N_24943);
nand UO_1898 (O_1898,N_24954,N_24959);
nand UO_1899 (O_1899,N_24861,N_24914);
and UO_1900 (O_1900,N_24918,N_24868);
nor UO_1901 (O_1901,N_24838,N_24823);
nor UO_1902 (O_1902,N_24925,N_24924);
nor UO_1903 (O_1903,N_24958,N_24930);
or UO_1904 (O_1904,N_24829,N_24956);
or UO_1905 (O_1905,N_24917,N_24933);
and UO_1906 (O_1906,N_24919,N_24845);
nor UO_1907 (O_1907,N_24801,N_24812);
nand UO_1908 (O_1908,N_24931,N_24841);
and UO_1909 (O_1909,N_24869,N_24832);
nand UO_1910 (O_1910,N_24954,N_24968);
or UO_1911 (O_1911,N_24850,N_24868);
or UO_1912 (O_1912,N_24990,N_24916);
nand UO_1913 (O_1913,N_24991,N_24947);
xnor UO_1914 (O_1914,N_24840,N_24896);
or UO_1915 (O_1915,N_24835,N_24814);
nand UO_1916 (O_1916,N_24841,N_24969);
or UO_1917 (O_1917,N_24842,N_24809);
nand UO_1918 (O_1918,N_24956,N_24823);
or UO_1919 (O_1919,N_24863,N_24848);
or UO_1920 (O_1920,N_24879,N_24962);
nand UO_1921 (O_1921,N_24990,N_24967);
nand UO_1922 (O_1922,N_24968,N_24809);
or UO_1923 (O_1923,N_24910,N_24920);
nor UO_1924 (O_1924,N_24890,N_24882);
and UO_1925 (O_1925,N_24928,N_24816);
and UO_1926 (O_1926,N_24869,N_24995);
nand UO_1927 (O_1927,N_24875,N_24872);
and UO_1928 (O_1928,N_24880,N_24935);
nor UO_1929 (O_1929,N_24940,N_24937);
and UO_1930 (O_1930,N_24955,N_24998);
or UO_1931 (O_1931,N_24868,N_24819);
or UO_1932 (O_1932,N_24865,N_24846);
nand UO_1933 (O_1933,N_24868,N_24926);
nor UO_1934 (O_1934,N_24946,N_24880);
and UO_1935 (O_1935,N_24901,N_24831);
and UO_1936 (O_1936,N_24914,N_24910);
nand UO_1937 (O_1937,N_24995,N_24996);
nor UO_1938 (O_1938,N_24918,N_24965);
xor UO_1939 (O_1939,N_24862,N_24989);
nand UO_1940 (O_1940,N_24902,N_24842);
nand UO_1941 (O_1941,N_24911,N_24840);
nor UO_1942 (O_1942,N_24946,N_24860);
or UO_1943 (O_1943,N_24877,N_24978);
nand UO_1944 (O_1944,N_24943,N_24917);
nor UO_1945 (O_1945,N_24849,N_24956);
or UO_1946 (O_1946,N_24957,N_24936);
or UO_1947 (O_1947,N_24872,N_24956);
nand UO_1948 (O_1948,N_24843,N_24848);
nand UO_1949 (O_1949,N_24962,N_24815);
or UO_1950 (O_1950,N_24953,N_24863);
nand UO_1951 (O_1951,N_24931,N_24939);
nor UO_1952 (O_1952,N_24920,N_24945);
nor UO_1953 (O_1953,N_24854,N_24801);
xor UO_1954 (O_1954,N_24894,N_24994);
and UO_1955 (O_1955,N_24960,N_24813);
nor UO_1956 (O_1956,N_24818,N_24973);
nor UO_1957 (O_1957,N_24905,N_24983);
and UO_1958 (O_1958,N_24949,N_24834);
and UO_1959 (O_1959,N_24853,N_24939);
and UO_1960 (O_1960,N_24878,N_24869);
or UO_1961 (O_1961,N_24888,N_24917);
nor UO_1962 (O_1962,N_24890,N_24816);
nor UO_1963 (O_1963,N_24999,N_24850);
nand UO_1964 (O_1964,N_24959,N_24892);
nor UO_1965 (O_1965,N_24967,N_24936);
nor UO_1966 (O_1966,N_24884,N_24877);
and UO_1967 (O_1967,N_24853,N_24886);
xnor UO_1968 (O_1968,N_24930,N_24831);
nor UO_1969 (O_1969,N_24830,N_24966);
and UO_1970 (O_1970,N_24957,N_24882);
or UO_1971 (O_1971,N_24860,N_24828);
nand UO_1972 (O_1972,N_24815,N_24839);
or UO_1973 (O_1973,N_24883,N_24843);
or UO_1974 (O_1974,N_24881,N_24997);
and UO_1975 (O_1975,N_24844,N_24895);
or UO_1976 (O_1976,N_24928,N_24994);
and UO_1977 (O_1977,N_24929,N_24908);
xnor UO_1978 (O_1978,N_24844,N_24993);
nand UO_1979 (O_1979,N_24926,N_24916);
nor UO_1980 (O_1980,N_24987,N_24895);
nand UO_1981 (O_1981,N_24830,N_24992);
and UO_1982 (O_1982,N_24887,N_24983);
or UO_1983 (O_1983,N_24934,N_24802);
nor UO_1984 (O_1984,N_24882,N_24926);
xnor UO_1985 (O_1985,N_24992,N_24848);
nand UO_1986 (O_1986,N_24865,N_24929);
or UO_1987 (O_1987,N_24941,N_24846);
or UO_1988 (O_1988,N_24916,N_24866);
and UO_1989 (O_1989,N_24985,N_24886);
nor UO_1990 (O_1990,N_24923,N_24933);
and UO_1991 (O_1991,N_24846,N_24956);
nand UO_1992 (O_1992,N_24817,N_24928);
nor UO_1993 (O_1993,N_24908,N_24967);
nor UO_1994 (O_1994,N_24824,N_24960);
xor UO_1995 (O_1995,N_24866,N_24996);
and UO_1996 (O_1996,N_24858,N_24808);
nor UO_1997 (O_1997,N_24907,N_24953);
nand UO_1998 (O_1998,N_24865,N_24939);
and UO_1999 (O_1999,N_24888,N_24970);
nor UO_2000 (O_2000,N_24822,N_24905);
nand UO_2001 (O_2001,N_24930,N_24882);
nor UO_2002 (O_2002,N_24804,N_24877);
nand UO_2003 (O_2003,N_24925,N_24835);
nor UO_2004 (O_2004,N_24830,N_24921);
or UO_2005 (O_2005,N_24817,N_24976);
and UO_2006 (O_2006,N_24837,N_24850);
nor UO_2007 (O_2007,N_24866,N_24820);
and UO_2008 (O_2008,N_24837,N_24879);
nand UO_2009 (O_2009,N_24991,N_24941);
xnor UO_2010 (O_2010,N_24828,N_24919);
xor UO_2011 (O_2011,N_24972,N_24902);
or UO_2012 (O_2012,N_24848,N_24819);
nor UO_2013 (O_2013,N_24815,N_24806);
nand UO_2014 (O_2014,N_24960,N_24997);
nand UO_2015 (O_2015,N_24947,N_24814);
or UO_2016 (O_2016,N_24885,N_24891);
nand UO_2017 (O_2017,N_24815,N_24840);
nand UO_2018 (O_2018,N_24811,N_24895);
nor UO_2019 (O_2019,N_24987,N_24864);
and UO_2020 (O_2020,N_24917,N_24836);
or UO_2021 (O_2021,N_24802,N_24866);
nor UO_2022 (O_2022,N_24891,N_24817);
or UO_2023 (O_2023,N_24861,N_24901);
nand UO_2024 (O_2024,N_24866,N_24978);
nor UO_2025 (O_2025,N_24804,N_24803);
nand UO_2026 (O_2026,N_24846,N_24950);
nand UO_2027 (O_2027,N_24900,N_24936);
and UO_2028 (O_2028,N_24881,N_24805);
or UO_2029 (O_2029,N_24934,N_24812);
xor UO_2030 (O_2030,N_24947,N_24808);
nand UO_2031 (O_2031,N_24902,N_24986);
nand UO_2032 (O_2032,N_24884,N_24882);
or UO_2033 (O_2033,N_24923,N_24840);
nand UO_2034 (O_2034,N_24912,N_24873);
xnor UO_2035 (O_2035,N_24817,N_24892);
nand UO_2036 (O_2036,N_24952,N_24963);
and UO_2037 (O_2037,N_24884,N_24829);
nand UO_2038 (O_2038,N_24808,N_24839);
or UO_2039 (O_2039,N_24872,N_24807);
nand UO_2040 (O_2040,N_24952,N_24826);
xor UO_2041 (O_2041,N_24981,N_24906);
nand UO_2042 (O_2042,N_24899,N_24892);
nor UO_2043 (O_2043,N_24888,N_24819);
xnor UO_2044 (O_2044,N_24897,N_24818);
and UO_2045 (O_2045,N_24928,N_24839);
and UO_2046 (O_2046,N_24949,N_24883);
and UO_2047 (O_2047,N_24922,N_24857);
nand UO_2048 (O_2048,N_24993,N_24943);
nand UO_2049 (O_2049,N_24941,N_24835);
nor UO_2050 (O_2050,N_24951,N_24997);
xor UO_2051 (O_2051,N_24837,N_24814);
nand UO_2052 (O_2052,N_24876,N_24810);
or UO_2053 (O_2053,N_24835,N_24932);
or UO_2054 (O_2054,N_24830,N_24947);
nand UO_2055 (O_2055,N_24941,N_24927);
xnor UO_2056 (O_2056,N_24968,N_24951);
nand UO_2057 (O_2057,N_24887,N_24863);
or UO_2058 (O_2058,N_24813,N_24933);
nor UO_2059 (O_2059,N_24805,N_24850);
and UO_2060 (O_2060,N_24827,N_24901);
or UO_2061 (O_2061,N_24989,N_24858);
nor UO_2062 (O_2062,N_24900,N_24915);
nand UO_2063 (O_2063,N_24907,N_24869);
nor UO_2064 (O_2064,N_24884,N_24930);
and UO_2065 (O_2065,N_24907,N_24830);
and UO_2066 (O_2066,N_24816,N_24913);
and UO_2067 (O_2067,N_24848,N_24803);
and UO_2068 (O_2068,N_24820,N_24986);
and UO_2069 (O_2069,N_24848,N_24958);
or UO_2070 (O_2070,N_24954,N_24815);
nor UO_2071 (O_2071,N_24893,N_24844);
xnor UO_2072 (O_2072,N_24934,N_24864);
xnor UO_2073 (O_2073,N_24928,N_24983);
and UO_2074 (O_2074,N_24967,N_24887);
nor UO_2075 (O_2075,N_24906,N_24912);
nand UO_2076 (O_2076,N_24810,N_24847);
and UO_2077 (O_2077,N_24963,N_24938);
or UO_2078 (O_2078,N_24803,N_24853);
nor UO_2079 (O_2079,N_24921,N_24908);
nor UO_2080 (O_2080,N_24810,N_24944);
and UO_2081 (O_2081,N_24989,N_24856);
nand UO_2082 (O_2082,N_24906,N_24807);
nor UO_2083 (O_2083,N_24903,N_24917);
nor UO_2084 (O_2084,N_24852,N_24830);
or UO_2085 (O_2085,N_24979,N_24899);
nor UO_2086 (O_2086,N_24906,N_24964);
or UO_2087 (O_2087,N_24821,N_24893);
and UO_2088 (O_2088,N_24912,N_24853);
and UO_2089 (O_2089,N_24813,N_24849);
nand UO_2090 (O_2090,N_24934,N_24950);
nor UO_2091 (O_2091,N_24977,N_24896);
nor UO_2092 (O_2092,N_24883,N_24945);
nor UO_2093 (O_2093,N_24892,N_24961);
xnor UO_2094 (O_2094,N_24876,N_24855);
or UO_2095 (O_2095,N_24951,N_24843);
and UO_2096 (O_2096,N_24927,N_24993);
nand UO_2097 (O_2097,N_24990,N_24819);
nand UO_2098 (O_2098,N_24877,N_24989);
and UO_2099 (O_2099,N_24854,N_24878);
and UO_2100 (O_2100,N_24863,N_24915);
nand UO_2101 (O_2101,N_24929,N_24955);
or UO_2102 (O_2102,N_24889,N_24860);
xnor UO_2103 (O_2103,N_24930,N_24860);
nand UO_2104 (O_2104,N_24929,N_24810);
nor UO_2105 (O_2105,N_24931,N_24922);
or UO_2106 (O_2106,N_24865,N_24972);
nand UO_2107 (O_2107,N_24876,N_24861);
and UO_2108 (O_2108,N_24838,N_24850);
or UO_2109 (O_2109,N_24955,N_24914);
and UO_2110 (O_2110,N_24896,N_24965);
xor UO_2111 (O_2111,N_24903,N_24918);
and UO_2112 (O_2112,N_24956,N_24842);
or UO_2113 (O_2113,N_24855,N_24950);
or UO_2114 (O_2114,N_24873,N_24959);
and UO_2115 (O_2115,N_24923,N_24804);
nor UO_2116 (O_2116,N_24833,N_24962);
or UO_2117 (O_2117,N_24872,N_24991);
or UO_2118 (O_2118,N_24845,N_24968);
and UO_2119 (O_2119,N_24858,N_24931);
and UO_2120 (O_2120,N_24874,N_24888);
or UO_2121 (O_2121,N_24948,N_24877);
and UO_2122 (O_2122,N_24985,N_24998);
and UO_2123 (O_2123,N_24961,N_24923);
xor UO_2124 (O_2124,N_24847,N_24849);
or UO_2125 (O_2125,N_24990,N_24915);
nor UO_2126 (O_2126,N_24879,N_24970);
nand UO_2127 (O_2127,N_24884,N_24996);
or UO_2128 (O_2128,N_24967,N_24941);
nand UO_2129 (O_2129,N_24813,N_24825);
nor UO_2130 (O_2130,N_24844,N_24865);
or UO_2131 (O_2131,N_24964,N_24953);
or UO_2132 (O_2132,N_24849,N_24997);
nor UO_2133 (O_2133,N_24978,N_24857);
xnor UO_2134 (O_2134,N_24961,N_24914);
and UO_2135 (O_2135,N_24977,N_24909);
nor UO_2136 (O_2136,N_24980,N_24944);
and UO_2137 (O_2137,N_24925,N_24992);
nand UO_2138 (O_2138,N_24808,N_24827);
or UO_2139 (O_2139,N_24848,N_24998);
nand UO_2140 (O_2140,N_24889,N_24915);
nand UO_2141 (O_2141,N_24834,N_24918);
and UO_2142 (O_2142,N_24894,N_24950);
nand UO_2143 (O_2143,N_24930,N_24838);
or UO_2144 (O_2144,N_24897,N_24848);
nor UO_2145 (O_2145,N_24994,N_24909);
or UO_2146 (O_2146,N_24830,N_24930);
nand UO_2147 (O_2147,N_24876,N_24997);
nor UO_2148 (O_2148,N_24853,N_24813);
nand UO_2149 (O_2149,N_24808,N_24982);
nand UO_2150 (O_2150,N_24968,N_24952);
and UO_2151 (O_2151,N_24812,N_24846);
and UO_2152 (O_2152,N_24830,N_24997);
and UO_2153 (O_2153,N_24990,N_24822);
and UO_2154 (O_2154,N_24983,N_24988);
nand UO_2155 (O_2155,N_24807,N_24856);
nand UO_2156 (O_2156,N_24802,N_24906);
nor UO_2157 (O_2157,N_24849,N_24944);
nand UO_2158 (O_2158,N_24964,N_24881);
or UO_2159 (O_2159,N_24845,N_24952);
nor UO_2160 (O_2160,N_24822,N_24984);
or UO_2161 (O_2161,N_24802,N_24967);
or UO_2162 (O_2162,N_24832,N_24967);
and UO_2163 (O_2163,N_24818,N_24852);
and UO_2164 (O_2164,N_24839,N_24886);
nand UO_2165 (O_2165,N_24896,N_24838);
or UO_2166 (O_2166,N_24947,N_24999);
nor UO_2167 (O_2167,N_24949,N_24872);
nand UO_2168 (O_2168,N_24839,N_24858);
xnor UO_2169 (O_2169,N_24930,N_24900);
and UO_2170 (O_2170,N_24822,N_24960);
and UO_2171 (O_2171,N_24872,N_24923);
nand UO_2172 (O_2172,N_24999,N_24854);
or UO_2173 (O_2173,N_24801,N_24915);
and UO_2174 (O_2174,N_24982,N_24827);
nand UO_2175 (O_2175,N_24954,N_24937);
nor UO_2176 (O_2176,N_24836,N_24858);
and UO_2177 (O_2177,N_24975,N_24845);
or UO_2178 (O_2178,N_24820,N_24857);
xor UO_2179 (O_2179,N_24861,N_24866);
and UO_2180 (O_2180,N_24834,N_24820);
nand UO_2181 (O_2181,N_24921,N_24901);
or UO_2182 (O_2182,N_24899,N_24821);
or UO_2183 (O_2183,N_24823,N_24916);
xor UO_2184 (O_2184,N_24974,N_24873);
nand UO_2185 (O_2185,N_24906,N_24988);
nand UO_2186 (O_2186,N_24855,N_24835);
or UO_2187 (O_2187,N_24994,N_24867);
and UO_2188 (O_2188,N_24909,N_24879);
and UO_2189 (O_2189,N_24966,N_24998);
or UO_2190 (O_2190,N_24817,N_24920);
and UO_2191 (O_2191,N_24838,N_24984);
nand UO_2192 (O_2192,N_24912,N_24950);
nor UO_2193 (O_2193,N_24978,N_24816);
nand UO_2194 (O_2194,N_24969,N_24850);
nor UO_2195 (O_2195,N_24800,N_24870);
nand UO_2196 (O_2196,N_24862,N_24987);
or UO_2197 (O_2197,N_24851,N_24971);
nand UO_2198 (O_2198,N_24892,N_24847);
and UO_2199 (O_2199,N_24838,N_24864);
or UO_2200 (O_2200,N_24927,N_24896);
and UO_2201 (O_2201,N_24932,N_24941);
nor UO_2202 (O_2202,N_24936,N_24815);
nand UO_2203 (O_2203,N_24981,N_24935);
xnor UO_2204 (O_2204,N_24871,N_24822);
nand UO_2205 (O_2205,N_24879,N_24896);
and UO_2206 (O_2206,N_24803,N_24864);
nand UO_2207 (O_2207,N_24825,N_24927);
nand UO_2208 (O_2208,N_24877,N_24838);
nand UO_2209 (O_2209,N_24861,N_24864);
nor UO_2210 (O_2210,N_24881,N_24864);
or UO_2211 (O_2211,N_24975,N_24853);
or UO_2212 (O_2212,N_24819,N_24812);
and UO_2213 (O_2213,N_24839,N_24968);
and UO_2214 (O_2214,N_24825,N_24823);
and UO_2215 (O_2215,N_24943,N_24895);
or UO_2216 (O_2216,N_24801,N_24803);
nand UO_2217 (O_2217,N_24972,N_24995);
or UO_2218 (O_2218,N_24854,N_24871);
nand UO_2219 (O_2219,N_24812,N_24824);
nand UO_2220 (O_2220,N_24827,N_24909);
nand UO_2221 (O_2221,N_24943,N_24998);
and UO_2222 (O_2222,N_24987,N_24894);
or UO_2223 (O_2223,N_24828,N_24877);
and UO_2224 (O_2224,N_24954,N_24924);
xnor UO_2225 (O_2225,N_24886,N_24884);
nor UO_2226 (O_2226,N_24845,N_24961);
and UO_2227 (O_2227,N_24939,N_24987);
and UO_2228 (O_2228,N_24915,N_24970);
or UO_2229 (O_2229,N_24828,N_24831);
nor UO_2230 (O_2230,N_24876,N_24819);
nand UO_2231 (O_2231,N_24835,N_24860);
and UO_2232 (O_2232,N_24816,N_24966);
or UO_2233 (O_2233,N_24869,N_24881);
nor UO_2234 (O_2234,N_24899,N_24844);
xnor UO_2235 (O_2235,N_24871,N_24951);
and UO_2236 (O_2236,N_24960,N_24885);
nand UO_2237 (O_2237,N_24870,N_24845);
and UO_2238 (O_2238,N_24963,N_24906);
nand UO_2239 (O_2239,N_24899,N_24833);
nand UO_2240 (O_2240,N_24892,N_24990);
nor UO_2241 (O_2241,N_24912,N_24918);
nor UO_2242 (O_2242,N_24904,N_24978);
nand UO_2243 (O_2243,N_24909,N_24821);
and UO_2244 (O_2244,N_24940,N_24844);
or UO_2245 (O_2245,N_24917,N_24950);
or UO_2246 (O_2246,N_24987,N_24852);
and UO_2247 (O_2247,N_24870,N_24920);
nand UO_2248 (O_2248,N_24820,N_24950);
xnor UO_2249 (O_2249,N_24920,N_24835);
or UO_2250 (O_2250,N_24844,N_24939);
or UO_2251 (O_2251,N_24995,N_24963);
nand UO_2252 (O_2252,N_24874,N_24910);
or UO_2253 (O_2253,N_24839,N_24859);
or UO_2254 (O_2254,N_24851,N_24826);
nand UO_2255 (O_2255,N_24830,N_24895);
and UO_2256 (O_2256,N_24989,N_24971);
nor UO_2257 (O_2257,N_24856,N_24904);
nand UO_2258 (O_2258,N_24911,N_24859);
and UO_2259 (O_2259,N_24845,N_24803);
nor UO_2260 (O_2260,N_24993,N_24850);
nand UO_2261 (O_2261,N_24905,N_24892);
xor UO_2262 (O_2262,N_24976,N_24844);
and UO_2263 (O_2263,N_24801,N_24869);
and UO_2264 (O_2264,N_24909,N_24946);
and UO_2265 (O_2265,N_24981,N_24868);
nand UO_2266 (O_2266,N_24998,N_24878);
and UO_2267 (O_2267,N_24825,N_24936);
nor UO_2268 (O_2268,N_24925,N_24988);
nand UO_2269 (O_2269,N_24965,N_24818);
nor UO_2270 (O_2270,N_24812,N_24959);
nor UO_2271 (O_2271,N_24879,N_24840);
and UO_2272 (O_2272,N_24833,N_24925);
nand UO_2273 (O_2273,N_24816,N_24933);
nor UO_2274 (O_2274,N_24800,N_24916);
nor UO_2275 (O_2275,N_24825,N_24834);
nand UO_2276 (O_2276,N_24948,N_24837);
nor UO_2277 (O_2277,N_24921,N_24809);
nor UO_2278 (O_2278,N_24998,N_24995);
and UO_2279 (O_2279,N_24884,N_24977);
or UO_2280 (O_2280,N_24936,N_24953);
nand UO_2281 (O_2281,N_24871,N_24978);
xor UO_2282 (O_2282,N_24917,N_24814);
nor UO_2283 (O_2283,N_24815,N_24868);
or UO_2284 (O_2284,N_24965,N_24998);
or UO_2285 (O_2285,N_24856,N_24871);
nor UO_2286 (O_2286,N_24943,N_24891);
or UO_2287 (O_2287,N_24983,N_24801);
nor UO_2288 (O_2288,N_24964,N_24824);
xor UO_2289 (O_2289,N_24818,N_24969);
nor UO_2290 (O_2290,N_24845,N_24966);
nand UO_2291 (O_2291,N_24824,N_24943);
nor UO_2292 (O_2292,N_24903,N_24985);
xnor UO_2293 (O_2293,N_24884,N_24994);
nand UO_2294 (O_2294,N_24826,N_24885);
nor UO_2295 (O_2295,N_24970,N_24807);
nor UO_2296 (O_2296,N_24886,N_24984);
and UO_2297 (O_2297,N_24869,N_24839);
and UO_2298 (O_2298,N_24874,N_24929);
and UO_2299 (O_2299,N_24861,N_24817);
xor UO_2300 (O_2300,N_24837,N_24872);
xnor UO_2301 (O_2301,N_24817,N_24938);
and UO_2302 (O_2302,N_24998,N_24977);
and UO_2303 (O_2303,N_24888,N_24982);
and UO_2304 (O_2304,N_24804,N_24827);
nor UO_2305 (O_2305,N_24802,N_24958);
nand UO_2306 (O_2306,N_24806,N_24986);
nand UO_2307 (O_2307,N_24931,N_24954);
and UO_2308 (O_2308,N_24959,N_24951);
nor UO_2309 (O_2309,N_24809,N_24932);
and UO_2310 (O_2310,N_24839,N_24949);
or UO_2311 (O_2311,N_24967,N_24829);
nand UO_2312 (O_2312,N_24812,N_24823);
nand UO_2313 (O_2313,N_24871,N_24963);
nand UO_2314 (O_2314,N_24938,N_24866);
xor UO_2315 (O_2315,N_24933,N_24971);
nor UO_2316 (O_2316,N_24920,N_24932);
nor UO_2317 (O_2317,N_24973,N_24850);
or UO_2318 (O_2318,N_24897,N_24802);
xnor UO_2319 (O_2319,N_24971,N_24877);
nand UO_2320 (O_2320,N_24818,N_24861);
and UO_2321 (O_2321,N_24836,N_24829);
nand UO_2322 (O_2322,N_24801,N_24861);
or UO_2323 (O_2323,N_24817,N_24854);
nor UO_2324 (O_2324,N_24806,N_24841);
or UO_2325 (O_2325,N_24940,N_24971);
nor UO_2326 (O_2326,N_24852,N_24827);
xor UO_2327 (O_2327,N_24850,N_24964);
nor UO_2328 (O_2328,N_24840,N_24984);
nand UO_2329 (O_2329,N_24973,N_24827);
and UO_2330 (O_2330,N_24845,N_24932);
nor UO_2331 (O_2331,N_24813,N_24827);
xnor UO_2332 (O_2332,N_24815,N_24972);
and UO_2333 (O_2333,N_24969,N_24807);
and UO_2334 (O_2334,N_24873,N_24813);
and UO_2335 (O_2335,N_24999,N_24932);
nand UO_2336 (O_2336,N_24967,N_24933);
nand UO_2337 (O_2337,N_24871,N_24810);
nor UO_2338 (O_2338,N_24985,N_24853);
or UO_2339 (O_2339,N_24823,N_24922);
nand UO_2340 (O_2340,N_24865,N_24979);
or UO_2341 (O_2341,N_24917,N_24995);
and UO_2342 (O_2342,N_24989,N_24901);
and UO_2343 (O_2343,N_24953,N_24850);
or UO_2344 (O_2344,N_24891,N_24803);
nand UO_2345 (O_2345,N_24897,N_24900);
or UO_2346 (O_2346,N_24805,N_24918);
nor UO_2347 (O_2347,N_24954,N_24843);
xnor UO_2348 (O_2348,N_24907,N_24968);
and UO_2349 (O_2349,N_24846,N_24851);
xor UO_2350 (O_2350,N_24877,N_24825);
or UO_2351 (O_2351,N_24937,N_24959);
and UO_2352 (O_2352,N_24882,N_24917);
and UO_2353 (O_2353,N_24833,N_24826);
nor UO_2354 (O_2354,N_24924,N_24866);
nand UO_2355 (O_2355,N_24872,N_24916);
or UO_2356 (O_2356,N_24918,N_24872);
or UO_2357 (O_2357,N_24967,N_24900);
nor UO_2358 (O_2358,N_24820,N_24918);
nor UO_2359 (O_2359,N_24996,N_24879);
nand UO_2360 (O_2360,N_24897,N_24806);
xor UO_2361 (O_2361,N_24869,N_24982);
or UO_2362 (O_2362,N_24964,N_24835);
nor UO_2363 (O_2363,N_24882,N_24830);
nand UO_2364 (O_2364,N_24858,N_24856);
xor UO_2365 (O_2365,N_24801,N_24943);
xor UO_2366 (O_2366,N_24937,N_24967);
xnor UO_2367 (O_2367,N_24923,N_24815);
nor UO_2368 (O_2368,N_24996,N_24847);
nor UO_2369 (O_2369,N_24963,N_24821);
or UO_2370 (O_2370,N_24862,N_24875);
xor UO_2371 (O_2371,N_24898,N_24886);
nand UO_2372 (O_2372,N_24973,N_24894);
or UO_2373 (O_2373,N_24954,N_24953);
nand UO_2374 (O_2374,N_24829,N_24948);
xor UO_2375 (O_2375,N_24864,N_24929);
and UO_2376 (O_2376,N_24978,N_24832);
and UO_2377 (O_2377,N_24992,N_24957);
or UO_2378 (O_2378,N_24885,N_24933);
nand UO_2379 (O_2379,N_24890,N_24969);
nand UO_2380 (O_2380,N_24939,N_24911);
nand UO_2381 (O_2381,N_24868,N_24997);
nor UO_2382 (O_2382,N_24965,N_24938);
nor UO_2383 (O_2383,N_24958,N_24853);
or UO_2384 (O_2384,N_24853,N_24920);
xnor UO_2385 (O_2385,N_24985,N_24967);
nor UO_2386 (O_2386,N_24862,N_24877);
or UO_2387 (O_2387,N_24998,N_24905);
or UO_2388 (O_2388,N_24913,N_24931);
or UO_2389 (O_2389,N_24847,N_24886);
or UO_2390 (O_2390,N_24860,N_24978);
nand UO_2391 (O_2391,N_24814,N_24994);
or UO_2392 (O_2392,N_24817,N_24855);
nor UO_2393 (O_2393,N_24853,N_24866);
and UO_2394 (O_2394,N_24940,N_24991);
xor UO_2395 (O_2395,N_24965,N_24914);
nand UO_2396 (O_2396,N_24974,N_24912);
xor UO_2397 (O_2397,N_24864,N_24868);
or UO_2398 (O_2398,N_24905,N_24872);
or UO_2399 (O_2399,N_24952,N_24824);
or UO_2400 (O_2400,N_24999,N_24898);
nand UO_2401 (O_2401,N_24908,N_24972);
or UO_2402 (O_2402,N_24969,N_24802);
or UO_2403 (O_2403,N_24854,N_24867);
and UO_2404 (O_2404,N_24882,N_24929);
and UO_2405 (O_2405,N_24940,N_24903);
or UO_2406 (O_2406,N_24825,N_24975);
nand UO_2407 (O_2407,N_24997,N_24906);
and UO_2408 (O_2408,N_24916,N_24806);
or UO_2409 (O_2409,N_24847,N_24880);
nand UO_2410 (O_2410,N_24907,N_24931);
nand UO_2411 (O_2411,N_24844,N_24973);
and UO_2412 (O_2412,N_24838,N_24920);
nor UO_2413 (O_2413,N_24902,N_24883);
nand UO_2414 (O_2414,N_24809,N_24911);
xnor UO_2415 (O_2415,N_24981,N_24932);
nand UO_2416 (O_2416,N_24891,N_24810);
nand UO_2417 (O_2417,N_24868,N_24882);
or UO_2418 (O_2418,N_24972,N_24999);
and UO_2419 (O_2419,N_24961,N_24863);
xor UO_2420 (O_2420,N_24907,N_24828);
nand UO_2421 (O_2421,N_24837,N_24875);
or UO_2422 (O_2422,N_24922,N_24933);
and UO_2423 (O_2423,N_24877,N_24895);
and UO_2424 (O_2424,N_24834,N_24992);
nand UO_2425 (O_2425,N_24865,N_24991);
nand UO_2426 (O_2426,N_24902,N_24814);
nor UO_2427 (O_2427,N_24923,N_24823);
nand UO_2428 (O_2428,N_24839,N_24971);
and UO_2429 (O_2429,N_24993,N_24885);
xnor UO_2430 (O_2430,N_24808,N_24930);
or UO_2431 (O_2431,N_24847,N_24804);
or UO_2432 (O_2432,N_24990,N_24856);
nand UO_2433 (O_2433,N_24950,N_24893);
and UO_2434 (O_2434,N_24943,N_24842);
xor UO_2435 (O_2435,N_24819,N_24975);
and UO_2436 (O_2436,N_24901,N_24812);
or UO_2437 (O_2437,N_24881,N_24815);
nand UO_2438 (O_2438,N_24859,N_24884);
and UO_2439 (O_2439,N_24976,N_24848);
or UO_2440 (O_2440,N_24924,N_24966);
and UO_2441 (O_2441,N_24844,N_24833);
nand UO_2442 (O_2442,N_24873,N_24940);
nor UO_2443 (O_2443,N_24938,N_24825);
nand UO_2444 (O_2444,N_24894,N_24991);
xnor UO_2445 (O_2445,N_24904,N_24944);
nand UO_2446 (O_2446,N_24920,N_24986);
and UO_2447 (O_2447,N_24928,N_24871);
and UO_2448 (O_2448,N_24857,N_24956);
nor UO_2449 (O_2449,N_24826,N_24934);
nand UO_2450 (O_2450,N_24844,N_24980);
and UO_2451 (O_2451,N_24813,N_24994);
and UO_2452 (O_2452,N_24816,N_24950);
nor UO_2453 (O_2453,N_24934,N_24908);
and UO_2454 (O_2454,N_24943,N_24930);
and UO_2455 (O_2455,N_24988,N_24962);
or UO_2456 (O_2456,N_24919,N_24844);
xnor UO_2457 (O_2457,N_24986,N_24989);
or UO_2458 (O_2458,N_24877,N_24824);
or UO_2459 (O_2459,N_24918,N_24983);
xnor UO_2460 (O_2460,N_24931,N_24861);
and UO_2461 (O_2461,N_24827,N_24966);
xnor UO_2462 (O_2462,N_24919,N_24897);
nor UO_2463 (O_2463,N_24908,N_24851);
nand UO_2464 (O_2464,N_24884,N_24997);
nor UO_2465 (O_2465,N_24890,N_24981);
nor UO_2466 (O_2466,N_24848,N_24896);
and UO_2467 (O_2467,N_24959,N_24893);
nand UO_2468 (O_2468,N_24917,N_24907);
nand UO_2469 (O_2469,N_24846,N_24805);
xnor UO_2470 (O_2470,N_24950,N_24967);
nand UO_2471 (O_2471,N_24820,N_24879);
xor UO_2472 (O_2472,N_24843,N_24877);
nand UO_2473 (O_2473,N_24948,N_24882);
nor UO_2474 (O_2474,N_24814,N_24866);
or UO_2475 (O_2475,N_24996,N_24890);
and UO_2476 (O_2476,N_24984,N_24910);
and UO_2477 (O_2477,N_24887,N_24817);
and UO_2478 (O_2478,N_24847,N_24995);
nand UO_2479 (O_2479,N_24845,N_24933);
and UO_2480 (O_2480,N_24929,N_24825);
or UO_2481 (O_2481,N_24930,N_24941);
nor UO_2482 (O_2482,N_24968,N_24850);
or UO_2483 (O_2483,N_24957,N_24841);
and UO_2484 (O_2484,N_24806,N_24998);
xor UO_2485 (O_2485,N_24888,N_24935);
or UO_2486 (O_2486,N_24938,N_24961);
nor UO_2487 (O_2487,N_24815,N_24988);
and UO_2488 (O_2488,N_24953,N_24835);
and UO_2489 (O_2489,N_24836,N_24904);
or UO_2490 (O_2490,N_24958,N_24904);
nor UO_2491 (O_2491,N_24830,N_24849);
or UO_2492 (O_2492,N_24854,N_24980);
and UO_2493 (O_2493,N_24972,N_24836);
nor UO_2494 (O_2494,N_24930,N_24857);
nand UO_2495 (O_2495,N_24875,N_24926);
nor UO_2496 (O_2496,N_24837,N_24993);
or UO_2497 (O_2497,N_24811,N_24891);
and UO_2498 (O_2498,N_24820,N_24967);
nand UO_2499 (O_2499,N_24988,N_24941);
xor UO_2500 (O_2500,N_24872,N_24841);
nor UO_2501 (O_2501,N_24867,N_24872);
xor UO_2502 (O_2502,N_24842,N_24882);
and UO_2503 (O_2503,N_24800,N_24965);
nand UO_2504 (O_2504,N_24921,N_24972);
nand UO_2505 (O_2505,N_24802,N_24886);
or UO_2506 (O_2506,N_24897,N_24816);
xnor UO_2507 (O_2507,N_24956,N_24936);
or UO_2508 (O_2508,N_24824,N_24881);
and UO_2509 (O_2509,N_24881,N_24861);
nand UO_2510 (O_2510,N_24856,N_24824);
and UO_2511 (O_2511,N_24831,N_24912);
nor UO_2512 (O_2512,N_24818,N_24865);
and UO_2513 (O_2513,N_24876,N_24946);
and UO_2514 (O_2514,N_24880,N_24975);
nand UO_2515 (O_2515,N_24849,N_24910);
and UO_2516 (O_2516,N_24857,N_24964);
or UO_2517 (O_2517,N_24970,N_24814);
nand UO_2518 (O_2518,N_24867,N_24832);
nor UO_2519 (O_2519,N_24950,N_24935);
nand UO_2520 (O_2520,N_24973,N_24877);
nor UO_2521 (O_2521,N_24931,N_24994);
nor UO_2522 (O_2522,N_24989,N_24802);
nor UO_2523 (O_2523,N_24826,N_24991);
and UO_2524 (O_2524,N_24840,N_24993);
or UO_2525 (O_2525,N_24856,N_24879);
and UO_2526 (O_2526,N_24855,N_24820);
and UO_2527 (O_2527,N_24916,N_24975);
nor UO_2528 (O_2528,N_24820,N_24971);
nand UO_2529 (O_2529,N_24868,N_24910);
nor UO_2530 (O_2530,N_24978,N_24991);
or UO_2531 (O_2531,N_24955,N_24941);
nor UO_2532 (O_2532,N_24959,N_24853);
xor UO_2533 (O_2533,N_24852,N_24955);
nor UO_2534 (O_2534,N_24816,N_24899);
nor UO_2535 (O_2535,N_24828,N_24872);
xnor UO_2536 (O_2536,N_24821,N_24974);
and UO_2537 (O_2537,N_24922,N_24943);
or UO_2538 (O_2538,N_24967,N_24878);
nand UO_2539 (O_2539,N_24819,N_24980);
and UO_2540 (O_2540,N_24847,N_24827);
nand UO_2541 (O_2541,N_24889,N_24877);
nand UO_2542 (O_2542,N_24893,N_24940);
nand UO_2543 (O_2543,N_24969,N_24905);
or UO_2544 (O_2544,N_24939,N_24928);
or UO_2545 (O_2545,N_24913,N_24976);
nand UO_2546 (O_2546,N_24949,N_24909);
nand UO_2547 (O_2547,N_24900,N_24874);
and UO_2548 (O_2548,N_24922,N_24839);
nand UO_2549 (O_2549,N_24998,N_24877);
xnor UO_2550 (O_2550,N_24832,N_24937);
and UO_2551 (O_2551,N_24835,N_24839);
xor UO_2552 (O_2552,N_24871,N_24890);
nor UO_2553 (O_2553,N_24940,N_24880);
and UO_2554 (O_2554,N_24865,N_24886);
nand UO_2555 (O_2555,N_24951,N_24896);
or UO_2556 (O_2556,N_24843,N_24922);
nor UO_2557 (O_2557,N_24809,N_24817);
or UO_2558 (O_2558,N_24838,N_24863);
xnor UO_2559 (O_2559,N_24883,N_24908);
or UO_2560 (O_2560,N_24841,N_24990);
nor UO_2561 (O_2561,N_24921,N_24898);
or UO_2562 (O_2562,N_24834,N_24944);
nor UO_2563 (O_2563,N_24955,N_24984);
nand UO_2564 (O_2564,N_24862,N_24976);
nand UO_2565 (O_2565,N_24858,N_24920);
nor UO_2566 (O_2566,N_24916,N_24938);
xnor UO_2567 (O_2567,N_24987,N_24859);
or UO_2568 (O_2568,N_24929,N_24841);
nor UO_2569 (O_2569,N_24818,N_24823);
xor UO_2570 (O_2570,N_24999,N_24945);
or UO_2571 (O_2571,N_24955,N_24822);
nand UO_2572 (O_2572,N_24930,N_24915);
and UO_2573 (O_2573,N_24824,N_24891);
or UO_2574 (O_2574,N_24869,N_24855);
and UO_2575 (O_2575,N_24922,N_24952);
or UO_2576 (O_2576,N_24880,N_24803);
xor UO_2577 (O_2577,N_24814,N_24861);
or UO_2578 (O_2578,N_24889,N_24982);
nor UO_2579 (O_2579,N_24884,N_24928);
or UO_2580 (O_2580,N_24966,N_24964);
and UO_2581 (O_2581,N_24989,N_24888);
nand UO_2582 (O_2582,N_24912,N_24847);
nor UO_2583 (O_2583,N_24929,N_24826);
xnor UO_2584 (O_2584,N_24854,N_24873);
nor UO_2585 (O_2585,N_24985,N_24828);
nor UO_2586 (O_2586,N_24871,N_24916);
nand UO_2587 (O_2587,N_24890,N_24925);
nor UO_2588 (O_2588,N_24826,N_24869);
and UO_2589 (O_2589,N_24928,N_24882);
and UO_2590 (O_2590,N_24918,N_24878);
xor UO_2591 (O_2591,N_24940,N_24875);
and UO_2592 (O_2592,N_24801,N_24850);
nand UO_2593 (O_2593,N_24864,N_24919);
or UO_2594 (O_2594,N_24909,N_24913);
or UO_2595 (O_2595,N_24816,N_24874);
nor UO_2596 (O_2596,N_24911,N_24821);
nor UO_2597 (O_2597,N_24942,N_24822);
and UO_2598 (O_2598,N_24919,N_24882);
and UO_2599 (O_2599,N_24978,N_24951);
nand UO_2600 (O_2600,N_24951,N_24966);
nor UO_2601 (O_2601,N_24998,N_24896);
nand UO_2602 (O_2602,N_24982,N_24909);
and UO_2603 (O_2603,N_24964,N_24886);
or UO_2604 (O_2604,N_24847,N_24867);
and UO_2605 (O_2605,N_24869,N_24842);
nand UO_2606 (O_2606,N_24842,N_24868);
nor UO_2607 (O_2607,N_24813,N_24917);
xor UO_2608 (O_2608,N_24929,N_24915);
or UO_2609 (O_2609,N_24833,N_24890);
nand UO_2610 (O_2610,N_24809,N_24985);
or UO_2611 (O_2611,N_24991,N_24938);
nor UO_2612 (O_2612,N_24880,N_24994);
nor UO_2613 (O_2613,N_24969,N_24842);
and UO_2614 (O_2614,N_24863,N_24938);
or UO_2615 (O_2615,N_24857,N_24910);
nand UO_2616 (O_2616,N_24916,N_24959);
or UO_2617 (O_2617,N_24912,N_24859);
xor UO_2618 (O_2618,N_24894,N_24917);
nor UO_2619 (O_2619,N_24959,N_24867);
xor UO_2620 (O_2620,N_24906,N_24948);
and UO_2621 (O_2621,N_24933,N_24897);
and UO_2622 (O_2622,N_24807,N_24873);
or UO_2623 (O_2623,N_24998,N_24812);
nor UO_2624 (O_2624,N_24864,N_24922);
or UO_2625 (O_2625,N_24985,N_24961);
and UO_2626 (O_2626,N_24915,N_24914);
nand UO_2627 (O_2627,N_24915,N_24954);
and UO_2628 (O_2628,N_24815,N_24845);
nand UO_2629 (O_2629,N_24802,N_24978);
and UO_2630 (O_2630,N_24963,N_24922);
or UO_2631 (O_2631,N_24890,N_24940);
nor UO_2632 (O_2632,N_24875,N_24901);
and UO_2633 (O_2633,N_24983,N_24800);
nor UO_2634 (O_2634,N_24826,N_24977);
or UO_2635 (O_2635,N_24919,N_24854);
nor UO_2636 (O_2636,N_24825,N_24949);
or UO_2637 (O_2637,N_24933,N_24888);
nor UO_2638 (O_2638,N_24822,N_24943);
or UO_2639 (O_2639,N_24847,N_24813);
and UO_2640 (O_2640,N_24886,N_24916);
nand UO_2641 (O_2641,N_24847,N_24920);
nand UO_2642 (O_2642,N_24815,N_24904);
or UO_2643 (O_2643,N_24963,N_24837);
nor UO_2644 (O_2644,N_24994,N_24864);
or UO_2645 (O_2645,N_24864,N_24954);
or UO_2646 (O_2646,N_24856,N_24893);
nor UO_2647 (O_2647,N_24837,N_24956);
and UO_2648 (O_2648,N_24948,N_24852);
and UO_2649 (O_2649,N_24851,N_24966);
or UO_2650 (O_2650,N_24883,N_24901);
nor UO_2651 (O_2651,N_24834,N_24804);
nand UO_2652 (O_2652,N_24944,N_24962);
or UO_2653 (O_2653,N_24902,N_24997);
nand UO_2654 (O_2654,N_24832,N_24825);
xnor UO_2655 (O_2655,N_24879,N_24919);
nand UO_2656 (O_2656,N_24845,N_24813);
and UO_2657 (O_2657,N_24962,N_24800);
nor UO_2658 (O_2658,N_24981,N_24853);
or UO_2659 (O_2659,N_24812,N_24912);
or UO_2660 (O_2660,N_24990,N_24989);
xnor UO_2661 (O_2661,N_24810,N_24959);
nor UO_2662 (O_2662,N_24807,N_24938);
and UO_2663 (O_2663,N_24960,N_24929);
nand UO_2664 (O_2664,N_24884,N_24822);
nand UO_2665 (O_2665,N_24889,N_24924);
nor UO_2666 (O_2666,N_24957,N_24805);
nand UO_2667 (O_2667,N_24912,N_24896);
xnor UO_2668 (O_2668,N_24823,N_24945);
or UO_2669 (O_2669,N_24858,N_24997);
and UO_2670 (O_2670,N_24886,N_24988);
or UO_2671 (O_2671,N_24935,N_24822);
xnor UO_2672 (O_2672,N_24946,N_24911);
nor UO_2673 (O_2673,N_24894,N_24995);
nand UO_2674 (O_2674,N_24953,N_24872);
nand UO_2675 (O_2675,N_24806,N_24901);
nand UO_2676 (O_2676,N_24830,N_24867);
nand UO_2677 (O_2677,N_24861,N_24812);
and UO_2678 (O_2678,N_24853,N_24954);
and UO_2679 (O_2679,N_24809,N_24964);
or UO_2680 (O_2680,N_24911,N_24954);
xnor UO_2681 (O_2681,N_24960,N_24875);
or UO_2682 (O_2682,N_24948,N_24899);
nor UO_2683 (O_2683,N_24990,N_24898);
or UO_2684 (O_2684,N_24864,N_24867);
and UO_2685 (O_2685,N_24960,N_24857);
or UO_2686 (O_2686,N_24999,N_24966);
xnor UO_2687 (O_2687,N_24932,N_24807);
and UO_2688 (O_2688,N_24893,N_24849);
or UO_2689 (O_2689,N_24919,N_24826);
nor UO_2690 (O_2690,N_24833,N_24858);
xnor UO_2691 (O_2691,N_24917,N_24860);
xnor UO_2692 (O_2692,N_24862,N_24820);
or UO_2693 (O_2693,N_24868,N_24855);
and UO_2694 (O_2694,N_24937,N_24907);
or UO_2695 (O_2695,N_24853,N_24898);
and UO_2696 (O_2696,N_24877,N_24949);
nand UO_2697 (O_2697,N_24906,N_24885);
and UO_2698 (O_2698,N_24833,N_24836);
or UO_2699 (O_2699,N_24961,N_24886);
and UO_2700 (O_2700,N_24889,N_24985);
and UO_2701 (O_2701,N_24833,N_24886);
and UO_2702 (O_2702,N_24965,N_24928);
xor UO_2703 (O_2703,N_24975,N_24959);
xnor UO_2704 (O_2704,N_24881,N_24917);
nand UO_2705 (O_2705,N_24824,N_24945);
or UO_2706 (O_2706,N_24959,N_24973);
or UO_2707 (O_2707,N_24813,N_24973);
nor UO_2708 (O_2708,N_24990,N_24821);
nand UO_2709 (O_2709,N_24964,N_24846);
and UO_2710 (O_2710,N_24951,N_24907);
nor UO_2711 (O_2711,N_24997,N_24819);
xnor UO_2712 (O_2712,N_24914,N_24870);
nor UO_2713 (O_2713,N_24961,N_24988);
or UO_2714 (O_2714,N_24830,N_24926);
and UO_2715 (O_2715,N_24873,N_24819);
nand UO_2716 (O_2716,N_24984,N_24922);
and UO_2717 (O_2717,N_24992,N_24964);
xnor UO_2718 (O_2718,N_24883,N_24957);
and UO_2719 (O_2719,N_24950,N_24997);
and UO_2720 (O_2720,N_24894,N_24804);
and UO_2721 (O_2721,N_24818,N_24992);
nand UO_2722 (O_2722,N_24904,N_24826);
nand UO_2723 (O_2723,N_24960,N_24840);
nand UO_2724 (O_2724,N_24913,N_24904);
or UO_2725 (O_2725,N_24900,N_24805);
and UO_2726 (O_2726,N_24980,N_24900);
and UO_2727 (O_2727,N_24940,N_24907);
nand UO_2728 (O_2728,N_24938,N_24805);
nand UO_2729 (O_2729,N_24832,N_24953);
xor UO_2730 (O_2730,N_24925,N_24829);
xor UO_2731 (O_2731,N_24848,N_24963);
and UO_2732 (O_2732,N_24959,N_24838);
nor UO_2733 (O_2733,N_24935,N_24830);
nand UO_2734 (O_2734,N_24831,N_24860);
xnor UO_2735 (O_2735,N_24930,N_24919);
nand UO_2736 (O_2736,N_24852,N_24909);
or UO_2737 (O_2737,N_24981,N_24968);
nand UO_2738 (O_2738,N_24985,N_24854);
or UO_2739 (O_2739,N_24916,N_24932);
and UO_2740 (O_2740,N_24903,N_24962);
xnor UO_2741 (O_2741,N_24942,N_24962);
and UO_2742 (O_2742,N_24895,N_24863);
or UO_2743 (O_2743,N_24947,N_24853);
nor UO_2744 (O_2744,N_24992,N_24961);
or UO_2745 (O_2745,N_24899,N_24985);
nor UO_2746 (O_2746,N_24896,N_24968);
and UO_2747 (O_2747,N_24995,N_24914);
nor UO_2748 (O_2748,N_24969,N_24955);
nor UO_2749 (O_2749,N_24972,N_24842);
and UO_2750 (O_2750,N_24915,N_24896);
nor UO_2751 (O_2751,N_24927,N_24952);
nand UO_2752 (O_2752,N_24873,N_24865);
or UO_2753 (O_2753,N_24871,N_24975);
nand UO_2754 (O_2754,N_24964,N_24879);
or UO_2755 (O_2755,N_24914,N_24823);
nand UO_2756 (O_2756,N_24983,N_24846);
or UO_2757 (O_2757,N_24836,N_24977);
nor UO_2758 (O_2758,N_24835,N_24841);
or UO_2759 (O_2759,N_24837,N_24876);
nor UO_2760 (O_2760,N_24925,N_24879);
nor UO_2761 (O_2761,N_24889,N_24801);
nor UO_2762 (O_2762,N_24908,N_24876);
xor UO_2763 (O_2763,N_24930,N_24901);
xnor UO_2764 (O_2764,N_24936,N_24952);
nand UO_2765 (O_2765,N_24883,N_24995);
or UO_2766 (O_2766,N_24937,N_24985);
or UO_2767 (O_2767,N_24897,N_24988);
nor UO_2768 (O_2768,N_24903,N_24870);
nand UO_2769 (O_2769,N_24962,N_24888);
nand UO_2770 (O_2770,N_24959,N_24941);
nor UO_2771 (O_2771,N_24984,N_24976);
and UO_2772 (O_2772,N_24807,N_24806);
or UO_2773 (O_2773,N_24967,N_24858);
nor UO_2774 (O_2774,N_24857,N_24931);
nor UO_2775 (O_2775,N_24944,N_24813);
and UO_2776 (O_2776,N_24983,N_24847);
nor UO_2777 (O_2777,N_24990,N_24886);
nand UO_2778 (O_2778,N_24871,N_24879);
or UO_2779 (O_2779,N_24877,N_24997);
or UO_2780 (O_2780,N_24815,N_24801);
nor UO_2781 (O_2781,N_24868,N_24923);
xor UO_2782 (O_2782,N_24941,N_24812);
and UO_2783 (O_2783,N_24847,N_24812);
xor UO_2784 (O_2784,N_24853,N_24816);
xnor UO_2785 (O_2785,N_24843,N_24809);
and UO_2786 (O_2786,N_24987,N_24826);
nand UO_2787 (O_2787,N_24809,N_24835);
nand UO_2788 (O_2788,N_24880,N_24964);
nand UO_2789 (O_2789,N_24861,N_24954);
nand UO_2790 (O_2790,N_24986,N_24906);
or UO_2791 (O_2791,N_24995,N_24811);
nand UO_2792 (O_2792,N_24916,N_24980);
or UO_2793 (O_2793,N_24844,N_24802);
xor UO_2794 (O_2794,N_24882,N_24969);
nand UO_2795 (O_2795,N_24962,N_24929);
nor UO_2796 (O_2796,N_24872,N_24829);
nand UO_2797 (O_2797,N_24846,N_24996);
nand UO_2798 (O_2798,N_24821,N_24856);
nor UO_2799 (O_2799,N_24841,N_24828);
nor UO_2800 (O_2800,N_24939,N_24974);
or UO_2801 (O_2801,N_24952,N_24842);
or UO_2802 (O_2802,N_24818,N_24878);
nor UO_2803 (O_2803,N_24902,N_24826);
nand UO_2804 (O_2804,N_24981,N_24843);
nor UO_2805 (O_2805,N_24884,N_24866);
xnor UO_2806 (O_2806,N_24810,N_24859);
nand UO_2807 (O_2807,N_24873,N_24899);
nand UO_2808 (O_2808,N_24938,N_24939);
nor UO_2809 (O_2809,N_24904,N_24921);
nor UO_2810 (O_2810,N_24965,N_24929);
or UO_2811 (O_2811,N_24948,N_24885);
nand UO_2812 (O_2812,N_24921,N_24944);
and UO_2813 (O_2813,N_24855,N_24989);
nand UO_2814 (O_2814,N_24882,N_24922);
and UO_2815 (O_2815,N_24959,N_24818);
and UO_2816 (O_2816,N_24878,N_24961);
or UO_2817 (O_2817,N_24848,N_24857);
xnor UO_2818 (O_2818,N_24951,N_24903);
nor UO_2819 (O_2819,N_24992,N_24816);
nand UO_2820 (O_2820,N_24840,N_24813);
and UO_2821 (O_2821,N_24868,N_24973);
or UO_2822 (O_2822,N_24983,N_24830);
nand UO_2823 (O_2823,N_24997,N_24807);
nor UO_2824 (O_2824,N_24885,N_24985);
and UO_2825 (O_2825,N_24937,N_24817);
nor UO_2826 (O_2826,N_24807,N_24911);
nor UO_2827 (O_2827,N_24825,N_24878);
nand UO_2828 (O_2828,N_24974,N_24820);
or UO_2829 (O_2829,N_24915,N_24841);
and UO_2830 (O_2830,N_24806,N_24929);
nand UO_2831 (O_2831,N_24851,N_24965);
and UO_2832 (O_2832,N_24937,N_24890);
and UO_2833 (O_2833,N_24930,N_24863);
and UO_2834 (O_2834,N_24951,N_24855);
nor UO_2835 (O_2835,N_24841,N_24907);
and UO_2836 (O_2836,N_24991,N_24969);
xor UO_2837 (O_2837,N_24960,N_24819);
nor UO_2838 (O_2838,N_24927,N_24858);
and UO_2839 (O_2839,N_24930,N_24867);
and UO_2840 (O_2840,N_24819,N_24926);
or UO_2841 (O_2841,N_24809,N_24941);
xor UO_2842 (O_2842,N_24800,N_24900);
and UO_2843 (O_2843,N_24802,N_24850);
nand UO_2844 (O_2844,N_24876,N_24829);
and UO_2845 (O_2845,N_24996,N_24917);
nand UO_2846 (O_2846,N_24823,N_24935);
nor UO_2847 (O_2847,N_24833,N_24882);
nor UO_2848 (O_2848,N_24939,N_24863);
xor UO_2849 (O_2849,N_24936,N_24977);
or UO_2850 (O_2850,N_24876,N_24938);
nand UO_2851 (O_2851,N_24945,N_24911);
or UO_2852 (O_2852,N_24869,N_24952);
or UO_2853 (O_2853,N_24979,N_24802);
xnor UO_2854 (O_2854,N_24929,N_24986);
nor UO_2855 (O_2855,N_24812,N_24938);
and UO_2856 (O_2856,N_24924,N_24934);
or UO_2857 (O_2857,N_24903,N_24923);
or UO_2858 (O_2858,N_24947,N_24835);
xnor UO_2859 (O_2859,N_24964,N_24854);
nand UO_2860 (O_2860,N_24903,N_24846);
nor UO_2861 (O_2861,N_24877,N_24985);
nor UO_2862 (O_2862,N_24884,N_24897);
nand UO_2863 (O_2863,N_24980,N_24965);
or UO_2864 (O_2864,N_24852,N_24894);
xnor UO_2865 (O_2865,N_24888,N_24849);
and UO_2866 (O_2866,N_24977,N_24860);
nand UO_2867 (O_2867,N_24822,N_24836);
and UO_2868 (O_2868,N_24925,N_24937);
nor UO_2869 (O_2869,N_24806,N_24843);
nor UO_2870 (O_2870,N_24830,N_24810);
or UO_2871 (O_2871,N_24895,N_24916);
or UO_2872 (O_2872,N_24964,N_24918);
nor UO_2873 (O_2873,N_24969,N_24808);
nand UO_2874 (O_2874,N_24989,N_24800);
nor UO_2875 (O_2875,N_24806,N_24941);
nand UO_2876 (O_2876,N_24865,N_24999);
or UO_2877 (O_2877,N_24982,N_24840);
or UO_2878 (O_2878,N_24861,N_24994);
xor UO_2879 (O_2879,N_24873,N_24980);
nor UO_2880 (O_2880,N_24825,N_24959);
nand UO_2881 (O_2881,N_24804,N_24910);
nand UO_2882 (O_2882,N_24819,N_24882);
or UO_2883 (O_2883,N_24939,N_24971);
or UO_2884 (O_2884,N_24905,N_24954);
and UO_2885 (O_2885,N_24851,N_24938);
nor UO_2886 (O_2886,N_24911,N_24970);
and UO_2887 (O_2887,N_24849,N_24861);
and UO_2888 (O_2888,N_24826,N_24855);
and UO_2889 (O_2889,N_24811,N_24830);
or UO_2890 (O_2890,N_24962,N_24980);
nand UO_2891 (O_2891,N_24869,N_24893);
nor UO_2892 (O_2892,N_24846,N_24818);
nand UO_2893 (O_2893,N_24852,N_24879);
nor UO_2894 (O_2894,N_24933,N_24934);
xor UO_2895 (O_2895,N_24843,N_24863);
nand UO_2896 (O_2896,N_24973,N_24931);
nand UO_2897 (O_2897,N_24911,N_24851);
nand UO_2898 (O_2898,N_24843,N_24969);
xor UO_2899 (O_2899,N_24978,N_24815);
and UO_2900 (O_2900,N_24810,N_24838);
nor UO_2901 (O_2901,N_24836,N_24815);
nor UO_2902 (O_2902,N_24807,N_24919);
nand UO_2903 (O_2903,N_24846,N_24998);
and UO_2904 (O_2904,N_24943,N_24850);
nand UO_2905 (O_2905,N_24846,N_24918);
or UO_2906 (O_2906,N_24994,N_24987);
and UO_2907 (O_2907,N_24929,N_24808);
and UO_2908 (O_2908,N_24906,N_24937);
or UO_2909 (O_2909,N_24899,N_24981);
nor UO_2910 (O_2910,N_24820,N_24919);
nand UO_2911 (O_2911,N_24909,N_24867);
and UO_2912 (O_2912,N_24887,N_24810);
and UO_2913 (O_2913,N_24951,N_24913);
or UO_2914 (O_2914,N_24815,N_24872);
and UO_2915 (O_2915,N_24878,N_24947);
xor UO_2916 (O_2916,N_24848,N_24899);
nand UO_2917 (O_2917,N_24875,N_24955);
nand UO_2918 (O_2918,N_24823,N_24863);
and UO_2919 (O_2919,N_24818,N_24869);
nor UO_2920 (O_2920,N_24895,N_24954);
nor UO_2921 (O_2921,N_24878,N_24802);
nand UO_2922 (O_2922,N_24999,N_24968);
nor UO_2923 (O_2923,N_24932,N_24874);
xor UO_2924 (O_2924,N_24848,N_24939);
nand UO_2925 (O_2925,N_24888,N_24847);
and UO_2926 (O_2926,N_24837,N_24886);
nand UO_2927 (O_2927,N_24885,N_24866);
and UO_2928 (O_2928,N_24906,N_24880);
or UO_2929 (O_2929,N_24821,N_24876);
nand UO_2930 (O_2930,N_24925,N_24839);
or UO_2931 (O_2931,N_24897,N_24991);
or UO_2932 (O_2932,N_24913,N_24942);
or UO_2933 (O_2933,N_24991,N_24867);
nor UO_2934 (O_2934,N_24972,N_24956);
xnor UO_2935 (O_2935,N_24972,N_24906);
nor UO_2936 (O_2936,N_24852,N_24839);
and UO_2937 (O_2937,N_24973,N_24915);
nand UO_2938 (O_2938,N_24846,N_24904);
nand UO_2939 (O_2939,N_24816,N_24976);
and UO_2940 (O_2940,N_24907,N_24956);
xor UO_2941 (O_2941,N_24917,N_24935);
and UO_2942 (O_2942,N_24948,N_24981);
and UO_2943 (O_2943,N_24928,N_24860);
and UO_2944 (O_2944,N_24898,N_24834);
nand UO_2945 (O_2945,N_24901,N_24813);
or UO_2946 (O_2946,N_24811,N_24935);
xnor UO_2947 (O_2947,N_24990,N_24860);
nor UO_2948 (O_2948,N_24970,N_24862);
or UO_2949 (O_2949,N_24813,N_24869);
and UO_2950 (O_2950,N_24976,N_24904);
nand UO_2951 (O_2951,N_24953,N_24979);
nor UO_2952 (O_2952,N_24931,N_24916);
and UO_2953 (O_2953,N_24886,N_24858);
or UO_2954 (O_2954,N_24958,N_24954);
and UO_2955 (O_2955,N_24830,N_24892);
nand UO_2956 (O_2956,N_24881,N_24886);
and UO_2957 (O_2957,N_24936,N_24883);
and UO_2958 (O_2958,N_24976,N_24954);
nor UO_2959 (O_2959,N_24966,N_24902);
nor UO_2960 (O_2960,N_24919,N_24910);
or UO_2961 (O_2961,N_24932,N_24976);
nor UO_2962 (O_2962,N_24847,N_24851);
or UO_2963 (O_2963,N_24844,N_24928);
and UO_2964 (O_2964,N_24888,N_24830);
nor UO_2965 (O_2965,N_24996,N_24814);
nand UO_2966 (O_2966,N_24885,N_24836);
or UO_2967 (O_2967,N_24916,N_24856);
nor UO_2968 (O_2968,N_24910,N_24941);
nor UO_2969 (O_2969,N_24895,N_24847);
or UO_2970 (O_2970,N_24960,N_24999);
or UO_2971 (O_2971,N_24943,N_24906);
nor UO_2972 (O_2972,N_24820,N_24800);
xnor UO_2973 (O_2973,N_24910,N_24903);
or UO_2974 (O_2974,N_24902,N_24838);
nor UO_2975 (O_2975,N_24817,N_24818);
and UO_2976 (O_2976,N_24877,N_24864);
or UO_2977 (O_2977,N_24957,N_24876);
nor UO_2978 (O_2978,N_24902,N_24868);
xnor UO_2979 (O_2979,N_24979,N_24993);
nand UO_2980 (O_2980,N_24807,N_24927);
nor UO_2981 (O_2981,N_24989,N_24887);
nor UO_2982 (O_2982,N_24846,N_24960);
and UO_2983 (O_2983,N_24827,N_24960);
or UO_2984 (O_2984,N_24939,N_24905);
or UO_2985 (O_2985,N_24902,N_24839);
xnor UO_2986 (O_2986,N_24851,N_24852);
and UO_2987 (O_2987,N_24938,N_24836);
and UO_2988 (O_2988,N_24965,N_24961);
or UO_2989 (O_2989,N_24990,N_24809);
nand UO_2990 (O_2990,N_24954,N_24961);
and UO_2991 (O_2991,N_24801,N_24958);
xor UO_2992 (O_2992,N_24859,N_24804);
nand UO_2993 (O_2993,N_24996,N_24973);
and UO_2994 (O_2994,N_24943,N_24997);
nand UO_2995 (O_2995,N_24863,N_24977);
and UO_2996 (O_2996,N_24874,N_24971);
nor UO_2997 (O_2997,N_24888,N_24875);
and UO_2998 (O_2998,N_24800,N_24855);
or UO_2999 (O_2999,N_24893,N_24895);
endmodule