module basic_500_3000_500_30_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_312,In_100);
nor U1 (N_1,In_466,In_402);
nand U2 (N_2,In_181,In_288);
nand U3 (N_3,In_279,In_172);
or U4 (N_4,In_206,In_482);
nor U5 (N_5,In_218,In_56);
and U6 (N_6,In_316,In_342);
nor U7 (N_7,In_48,In_258);
and U8 (N_8,In_45,In_368);
nand U9 (N_9,In_201,In_203);
xnor U10 (N_10,In_371,In_391);
nand U11 (N_11,In_324,In_365);
nor U12 (N_12,In_269,In_23);
nor U13 (N_13,In_35,In_427);
or U14 (N_14,In_164,In_110);
nand U15 (N_15,In_426,In_90);
or U16 (N_16,In_451,In_198);
or U17 (N_17,In_327,In_8);
nor U18 (N_18,In_242,In_386);
nor U19 (N_19,In_339,In_27);
and U20 (N_20,In_433,In_65);
and U21 (N_21,In_244,In_464);
nand U22 (N_22,In_447,In_334);
and U23 (N_23,In_61,In_184);
and U24 (N_24,In_262,In_470);
or U25 (N_25,In_131,In_193);
nor U26 (N_26,In_301,In_360);
nor U27 (N_27,In_467,In_335);
nor U28 (N_28,In_353,In_204);
nand U29 (N_29,In_122,In_369);
or U30 (N_30,In_485,In_21);
nand U31 (N_31,In_69,In_424);
nand U32 (N_32,In_320,In_498);
and U33 (N_33,In_257,In_125);
or U34 (N_34,In_412,In_41);
or U35 (N_35,In_51,In_345);
nor U36 (N_36,In_382,In_421);
nand U37 (N_37,In_175,In_118);
or U38 (N_38,In_144,In_154);
nand U39 (N_39,In_180,In_2);
or U40 (N_40,In_230,In_481);
nand U41 (N_41,In_457,In_147);
or U42 (N_42,In_162,In_101);
or U43 (N_43,In_153,In_7);
or U44 (N_44,In_190,In_285);
and U45 (N_45,In_121,In_410);
nor U46 (N_46,In_50,In_474);
or U47 (N_47,In_140,In_418);
and U48 (N_48,In_489,In_394);
or U49 (N_49,In_321,In_333);
and U50 (N_50,In_444,In_483);
nand U51 (N_51,In_170,In_212);
nand U52 (N_52,In_194,In_17);
or U53 (N_53,In_337,In_476);
nand U54 (N_54,In_52,In_416);
xor U55 (N_55,In_494,In_77);
nand U56 (N_56,In_362,In_272);
nand U57 (N_57,In_74,In_208);
xnor U58 (N_58,In_340,In_16);
or U59 (N_59,In_59,In_216);
nor U60 (N_60,In_254,In_165);
or U61 (N_61,In_273,In_471);
and U62 (N_62,In_88,In_192);
xor U63 (N_63,In_430,In_449);
or U64 (N_64,In_383,In_231);
nand U65 (N_65,In_207,In_409);
and U66 (N_66,In_209,In_239);
xor U67 (N_67,In_63,In_249);
nand U68 (N_68,In_159,In_443);
or U69 (N_69,In_156,In_176);
xor U70 (N_70,In_267,In_404);
or U71 (N_71,In_114,In_91);
or U72 (N_72,In_160,In_343);
and U73 (N_73,In_103,In_112);
nor U74 (N_74,In_469,In_350);
nand U75 (N_75,In_119,In_33);
nand U76 (N_76,In_490,In_492);
or U77 (N_77,In_86,In_168);
nor U78 (N_78,In_438,In_349);
or U79 (N_79,In_256,In_484);
nor U80 (N_80,In_352,In_326);
nand U81 (N_81,In_178,In_379);
nand U82 (N_82,In_96,In_22);
xor U83 (N_83,In_57,In_472);
nand U84 (N_84,In_274,In_32);
nand U85 (N_85,In_313,In_167);
xnor U86 (N_86,In_75,In_82);
and U87 (N_87,In_437,In_486);
nand U88 (N_88,In_309,In_297);
nand U89 (N_89,In_259,In_452);
or U90 (N_90,In_431,In_221);
nand U91 (N_91,In_60,In_432);
and U92 (N_92,In_113,In_133);
nor U93 (N_93,In_338,In_93);
xnor U94 (N_94,In_227,In_264);
nor U95 (N_95,In_141,In_381);
nand U96 (N_96,In_450,In_473);
nand U97 (N_97,In_278,In_106);
and U98 (N_98,In_135,In_46);
or U99 (N_99,In_459,In_169);
nor U100 (N_100,N_16,N_79);
xor U101 (N_101,In_346,N_99);
or U102 (N_102,In_357,N_55);
xor U103 (N_103,N_83,In_54);
xor U104 (N_104,N_21,N_23);
or U105 (N_105,In_58,N_86);
or U106 (N_106,N_76,In_329);
or U107 (N_107,N_71,In_129);
or U108 (N_108,In_290,N_15);
nor U109 (N_109,In_456,In_434);
nand U110 (N_110,N_73,In_270);
and U111 (N_111,In_191,In_105);
and U112 (N_112,In_255,N_89);
or U113 (N_113,In_62,In_370);
nor U114 (N_114,In_89,In_398);
and U115 (N_115,N_48,In_390);
xnor U116 (N_116,N_6,In_148);
nand U117 (N_117,In_67,In_493);
and U118 (N_118,In_328,In_419);
nand U119 (N_119,N_84,In_13);
nand U120 (N_120,N_96,N_13);
or U121 (N_121,In_29,N_36);
nor U122 (N_122,In_263,In_94);
and U123 (N_123,N_44,N_91);
nand U124 (N_124,N_8,N_60);
nor U125 (N_125,In_445,N_38);
and U126 (N_126,In_425,N_3);
nand U127 (N_127,In_4,N_4);
nand U128 (N_128,In_377,In_496);
nor U129 (N_129,In_210,In_189);
or U130 (N_130,N_78,N_2);
xor U131 (N_131,In_187,In_199);
and U132 (N_132,In_39,In_414);
or U133 (N_133,In_38,In_411);
nor U134 (N_134,In_238,In_202);
and U135 (N_135,In_401,In_436);
xor U136 (N_136,In_364,In_130);
nor U137 (N_137,In_115,In_405);
or U138 (N_138,In_378,N_52);
xor U139 (N_139,In_149,In_146);
nand U140 (N_140,N_58,In_475);
xor U141 (N_141,In_384,In_214);
nor U142 (N_142,In_143,In_3);
xor U143 (N_143,In_454,In_463);
and U144 (N_144,In_79,In_399);
and U145 (N_145,In_217,N_95);
and U146 (N_146,In_289,In_186);
nand U147 (N_147,In_196,N_28);
or U148 (N_148,In_299,In_80);
xor U149 (N_149,N_14,N_37);
or U150 (N_150,In_302,In_158);
and U151 (N_151,In_64,N_70);
nor U152 (N_152,N_61,In_376);
nor U153 (N_153,N_18,In_407);
and U154 (N_154,N_92,In_173);
or U155 (N_155,In_387,In_36);
nor U156 (N_156,In_12,N_41);
nand U157 (N_157,In_223,N_54);
nor U158 (N_158,In_277,In_47);
nand U159 (N_159,In_11,In_499);
and U160 (N_160,In_348,In_136);
or U161 (N_161,In_31,In_422);
nor U162 (N_162,In_367,N_1);
nor U163 (N_163,In_71,In_373);
nor U164 (N_164,In_462,In_374);
nor U165 (N_165,In_363,In_83);
nor U166 (N_166,N_11,N_67);
or U167 (N_167,In_322,N_59);
or U168 (N_168,In_446,In_247);
nand U169 (N_169,N_94,In_250);
nand U170 (N_170,In_219,In_372);
and U171 (N_171,In_479,In_229);
nand U172 (N_172,N_75,In_314);
and U173 (N_173,In_318,In_157);
or U174 (N_174,In_14,In_171);
nand U175 (N_175,In_1,In_491);
and U176 (N_176,In_226,In_355);
and U177 (N_177,In_179,In_81);
and U178 (N_178,In_0,In_102);
or U179 (N_179,N_69,In_319);
nand U180 (N_180,In_265,In_403);
and U181 (N_181,In_304,In_420);
and U182 (N_182,In_417,In_25);
nand U183 (N_183,In_253,In_161);
nor U184 (N_184,In_366,In_232);
nor U185 (N_185,In_497,In_97);
nor U186 (N_186,N_20,In_468);
and U187 (N_187,N_33,In_174);
and U188 (N_188,In_281,In_18);
nand U189 (N_189,In_336,In_392);
nand U190 (N_190,In_236,In_183);
and U191 (N_191,In_116,N_9);
nor U192 (N_192,In_477,In_271);
nor U193 (N_193,In_20,N_25);
and U194 (N_194,N_49,In_315);
nor U195 (N_195,N_82,In_408);
nor U196 (N_196,N_63,In_220);
nand U197 (N_197,In_235,N_40);
and U198 (N_198,In_155,In_243);
or U199 (N_199,In_282,In_276);
or U200 (N_200,N_109,N_103);
nor U201 (N_201,In_423,N_178);
or U202 (N_202,In_361,In_344);
nor U203 (N_203,In_85,In_240);
nand U204 (N_204,N_57,N_117);
or U205 (N_205,In_460,In_9);
xor U206 (N_206,N_199,N_68);
nand U207 (N_207,N_0,In_480);
nor U208 (N_208,N_65,In_305);
or U209 (N_209,In_99,In_351);
or U210 (N_210,In_448,In_461);
or U211 (N_211,N_45,N_170);
nand U212 (N_212,N_93,N_185);
nor U213 (N_213,N_128,N_7);
nor U214 (N_214,In_225,In_311);
and U215 (N_215,N_149,In_395);
nor U216 (N_216,N_163,N_24);
nor U217 (N_217,In_78,N_124);
xnor U218 (N_218,In_117,In_123);
and U219 (N_219,N_35,In_87);
or U220 (N_220,N_22,In_44);
xor U221 (N_221,In_294,In_246);
nor U222 (N_222,In_295,N_160);
or U223 (N_223,In_134,In_185);
nand U224 (N_224,N_136,In_42);
and U225 (N_225,N_166,N_100);
nor U226 (N_226,In_92,N_111);
and U227 (N_227,In_393,In_248);
or U228 (N_228,N_191,N_196);
or U229 (N_229,N_171,N_150);
and U230 (N_230,N_62,N_141);
nand U231 (N_231,N_139,N_133);
nor U232 (N_232,In_465,In_435);
or U233 (N_233,In_150,N_74);
nand U234 (N_234,N_119,In_128);
nor U235 (N_235,N_143,N_107);
and U236 (N_236,In_177,In_126);
nand U237 (N_237,N_26,N_114);
or U238 (N_238,In_300,In_275);
nand U239 (N_239,In_317,In_73);
or U240 (N_240,In_195,N_168);
nor U241 (N_241,N_157,N_179);
and U242 (N_242,N_123,In_109);
nor U243 (N_243,In_323,N_10);
nor U244 (N_244,N_108,In_111);
nand U245 (N_245,In_211,In_237);
xnor U246 (N_246,N_131,In_388);
and U247 (N_247,In_213,N_156);
and U248 (N_248,In_380,In_389);
and U249 (N_249,N_72,N_151);
or U250 (N_250,In_453,In_287);
nor U251 (N_251,N_145,In_331);
or U252 (N_252,N_32,In_188);
xor U253 (N_253,In_413,N_101);
or U254 (N_254,N_43,N_46);
nor U255 (N_255,N_97,N_120);
and U256 (N_256,N_187,In_325);
or U257 (N_257,In_95,N_190);
or U258 (N_258,N_152,N_34);
and U259 (N_259,In_152,In_332);
and U260 (N_260,In_127,N_104);
nand U261 (N_261,N_116,N_153);
and U262 (N_262,N_146,N_195);
nor U263 (N_263,In_347,In_132);
nand U264 (N_264,N_167,In_293);
and U265 (N_265,N_88,N_126);
nor U266 (N_266,In_163,N_176);
and U267 (N_267,In_241,In_428);
or U268 (N_268,N_137,In_458);
nand U269 (N_269,N_125,N_19);
nor U270 (N_270,In_358,N_132);
and U271 (N_271,N_173,N_147);
and U272 (N_272,In_268,N_47);
and U273 (N_273,In_222,N_184);
nand U274 (N_274,In_205,N_66);
nor U275 (N_275,In_139,N_106);
and U276 (N_276,In_280,N_113);
nor U277 (N_277,N_129,In_30);
and U278 (N_278,N_189,In_234);
or U279 (N_279,In_495,N_138);
xnor U280 (N_280,In_37,N_192);
nor U281 (N_281,In_266,In_406);
and U282 (N_282,In_26,In_76);
or U283 (N_283,In_487,N_42);
nand U284 (N_284,N_56,In_120);
xnor U285 (N_285,In_303,In_107);
and U286 (N_286,N_154,N_77);
and U287 (N_287,In_15,N_87);
nand U288 (N_288,N_174,N_27);
or U289 (N_289,N_135,N_110);
and U290 (N_290,N_127,In_306);
nand U291 (N_291,N_162,N_155);
xnor U292 (N_292,In_251,N_98);
and U293 (N_293,N_161,In_224);
nand U294 (N_294,N_17,N_181);
nand U295 (N_295,In_151,In_298);
and U296 (N_296,N_30,N_90);
and U297 (N_297,In_108,In_34);
xnor U298 (N_298,N_182,In_98);
xor U299 (N_299,N_31,N_112);
and U300 (N_300,N_208,N_248);
and U301 (N_301,In_70,In_397);
xnor U302 (N_302,In_138,In_145);
or U303 (N_303,N_277,N_12);
or U304 (N_304,N_246,In_261);
nand U305 (N_305,N_286,In_28);
nor U306 (N_306,N_215,N_297);
xnor U307 (N_307,N_265,N_232);
nand U308 (N_308,In_359,N_198);
xor U309 (N_309,N_194,In_415);
nor U310 (N_310,N_225,N_188);
or U311 (N_311,In_245,In_68);
or U312 (N_312,In_233,N_293);
and U313 (N_313,N_296,N_214);
or U314 (N_314,N_241,N_287);
nor U315 (N_315,In_66,N_223);
or U316 (N_316,N_266,In_488);
and U317 (N_317,N_219,N_252);
nor U318 (N_318,N_81,N_222);
nand U319 (N_319,In_72,N_276);
xnor U320 (N_320,N_235,N_285);
or U321 (N_321,N_39,N_236);
nor U322 (N_322,In_354,N_228);
and U323 (N_323,In_286,In_330);
and U324 (N_324,N_294,N_250);
nand U325 (N_325,N_279,In_252);
xnor U326 (N_326,N_262,N_165);
or U327 (N_327,N_234,N_224);
or U328 (N_328,N_205,N_227);
or U329 (N_329,N_118,N_238);
nand U330 (N_330,N_269,N_233);
or U331 (N_331,In_400,N_142);
or U332 (N_332,N_230,In_441);
and U333 (N_333,N_254,N_50);
xor U334 (N_334,N_284,N_212);
nor U335 (N_335,N_245,In_137);
xor U336 (N_336,N_272,N_211);
nor U337 (N_337,N_283,N_217);
nor U338 (N_338,In_5,In_40);
and U339 (N_339,N_175,In_375);
or U340 (N_340,N_244,In_341);
nand U341 (N_341,In_455,N_260);
or U342 (N_342,In_292,In_10);
nand U343 (N_343,N_259,N_207);
and U344 (N_344,N_264,N_202);
nor U345 (N_345,In_49,In_215);
xnor U346 (N_346,In_55,N_158);
or U347 (N_347,N_140,N_172);
or U348 (N_348,N_209,In_442);
and U349 (N_349,N_249,N_213);
nand U350 (N_350,N_295,N_148);
nor U351 (N_351,N_164,In_200);
nand U352 (N_352,N_51,In_84);
nand U353 (N_353,N_289,N_102);
nor U354 (N_354,N_203,N_299);
nand U355 (N_355,N_5,N_240);
nor U356 (N_356,N_255,N_159);
and U357 (N_357,N_183,In_291);
nand U358 (N_358,N_257,In_478);
nand U359 (N_359,N_239,N_231);
or U360 (N_360,N_247,In_182);
nand U361 (N_361,N_242,N_201);
and U362 (N_362,N_29,In_296);
nand U363 (N_363,In_396,N_274);
and U364 (N_364,N_271,N_221);
nor U365 (N_365,In_142,N_115);
and U366 (N_366,N_251,In_43);
nand U367 (N_367,N_292,N_243);
or U368 (N_368,In_53,In_104);
nand U369 (N_369,In_197,N_134);
or U370 (N_370,N_229,N_180);
xnor U371 (N_371,N_261,N_85);
or U372 (N_372,In_166,N_282);
or U373 (N_373,N_273,In_385);
nand U374 (N_374,In_284,N_144);
and U375 (N_375,In_439,N_64);
or U376 (N_376,In_308,In_6);
nor U377 (N_377,N_218,N_291);
or U378 (N_378,In_24,N_268);
nor U379 (N_379,N_258,In_429);
nand U380 (N_380,N_263,N_177);
nand U381 (N_381,N_204,In_228);
nor U382 (N_382,In_260,N_290);
and U383 (N_383,N_270,N_281);
nand U384 (N_384,N_193,N_280);
xnor U385 (N_385,N_275,N_53);
nand U386 (N_386,N_197,N_169);
and U387 (N_387,N_206,In_310);
or U388 (N_388,In_440,In_283);
and U389 (N_389,N_267,N_220);
nor U390 (N_390,N_216,N_278);
nand U391 (N_391,N_200,In_19);
nor U392 (N_392,N_226,N_186);
xor U393 (N_393,N_298,In_356);
xnor U394 (N_394,N_121,N_256);
nand U395 (N_395,In_307,N_130);
and U396 (N_396,N_80,N_237);
nand U397 (N_397,N_288,In_124);
and U398 (N_398,N_253,N_105);
nor U399 (N_399,N_210,N_122);
and U400 (N_400,N_378,N_382);
nand U401 (N_401,N_328,N_391);
and U402 (N_402,N_332,N_380);
nor U403 (N_403,N_393,N_357);
or U404 (N_404,N_385,N_358);
nand U405 (N_405,N_356,N_364);
xor U406 (N_406,N_388,N_306);
nand U407 (N_407,N_383,N_390);
and U408 (N_408,N_327,N_348);
and U409 (N_409,N_374,N_384);
nor U410 (N_410,N_347,N_373);
xor U411 (N_411,N_366,N_363);
xnor U412 (N_412,N_344,N_341);
and U413 (N_413,N_389,N_340);
or U414 (N_414,N_314,N_338);
or U415 (N_415,N_333,N_326);
nor U416 (N_416,N_323,N_320);
and U417 (N_417,N_312,N_361);
nand U418 (N_418,N_330,N_334);
nand U419 (N_419,N_369,N_302);
and U420 (N_420,N_370,N_317);
or U421 (N_421,N_387,N_376);
nor U422 (N_422,N_324,N_396);
or U423 (N_423,N_355,N_325);
xnor U424 (N_424,N_398,N_365);
and U425 (N_425,N_350,N_329);
nand U426 (N_426,N_381,N_372);
and U427 (N_427,N_392,N_321);
nor U428 (N_428,N_346,N_351);
and U429 (N_429,N_395,N_315);
and U430 (N_430,N_318,N_311);
or U431 (N_431,N_319,N_301);
or U432 (N_432,N_310,N_379);
nand U433 (N_433,N_308,N_375);
nor U434 (N_434,N_397,N_322);
nand U435 (N_435,N_399,N_359);
nor U436 (N_436,N_353,N_368);
and U437 (N_437,N_386,N_345);
or U438 (N_438,N_313,N_360);
and U439 (N_439,N_339,N_367);
or U440 (N_440,N_305,N_307);
xnor U441 (N_441,N_354,N_304);
and U442 (N_442,N_337,N_336);
and U443 (N_443,N_342,N_309);
nand U444 (N_444,N_349,N_303);
or U445 (N_445,N_343,N_362);
or U446 (N_446,N_331,N_335);
and U447 (N_447,N_394,N_352);
nand U448 (N_448,N_300,N_371);
nor U449 (N_449,N_316,N_377);
nand U450 (N_450,N_340,N_367);
and U451 (N_451,N_369,N_326);
and U452 (N_452,N_353,N_393);
xor U453 (N_453,N_302,N_391);
nand U454 (N_454,N_324,N_369);
nand U455 (N_455,N_318,N_361);
or U456 (N_456,N_308,N_306);
nor U457 (N_457,N_327,N_321);
or U458 (N_458,N_311,N_334);
or U459 (N_459,N_321,N_329);
and U460 (N_460,N_374,N_335);
nand U461 (N_461,N_309,N_336);
or U462 (N_462,N_398,N_357);
nand U463 (N_463,N_344,N_396);
nand U464 (N_464,N_324,N_309);
and U465 (N_465,N_358,N_396);
nor U466 (N_466,N_376,N_371);
or U467 (N_467,N_374,N_316);
nor U468 (N_468,N_323,N_325);
nor U469 (N_469,N_349,N_366);
or U470 (N_470,N_387,N_325);
nor U471 (N_471,N_379,N_307);
or U472 (N_472,N_364,N_320);
and U473 (N_473,N_335,N_339);
nand U474 (N_474,N_371,N_322);
or U475 (N_475,N_348,N_384);
or U476 (N_476,N_383,N_367);
or U477 (N_477,N_330,N_329);
xnor U478 (N_478,N_314,N_393);
nor U479 (N_479,N_353,N_381);
nor U480 (N_480,N_360,N_319);
nand U481 (N_481,N_301,N_348);
or U482 (N_482,N_353,N_305);
or U483 (N_483,N_347,N_317);
or U484 (N_484,N_340,N_354);
nand U485 (N_485,N_349,N_350);
and U486 (N_486,N_333,N_389);
and U487 (N_487,N_321,N_371);
or U488 (N_488,N_321,N_345);
and U489 (N_489,N_316,N_329);
or U490 (N_490,N_364,N_353);
nor U491 (N_491,N_378,N_364);
or U492 (N_492,N_371,N_346);
nor U493 (N_493,N_370,N_395);
xor U494 (N_494,N_363,N_334);
nand U495 (N_495,N_351,N_359);
xor U496 (N_496,N_387,N_319);
nor U497 (N_497,N_392,N_363);
nand U498 (N_498,N_320,N_308);
nor U499 (N_499,N_348,N_365);
nand U500 (N_500,N_426,N_441);
and U501 (N_501,N_469,N_434);
or U502 (N_502,N_465,N_499);
and U503 (N_503,N_460,N_440);
nor U504 (N_504,N_450,N_480);
and U505 (N_505,N_461,N_430);
nand U506 (N_506,N_463,N_448);
nor U507 (N_507,N_452,N_400);
xor U508 (N_508,N_418,N_408);
nand U509 (N_509,N_457,N_409);
nor U510 (N_510,N_402,N_427);
and U511 (N_511,N_429,N_494);
nand U512 (N_512,N_436,N_417);
or U513 (N_513,N_486,N_459);
or U514 (N_514,N_456,N_423);
and U515 (N_515,N_445,N_449);
and U516 (N_516,N_488,N_416);
and U517 (N_517,N_483,N_458);
nand U518 (N_518,N_411,N_432);
nand U519 (N_519,N_497,N_472);
nand U520 (N_520,N_451,N_481);
and U521 (N_521,N_419,N_495);
or U522 (N_522,N_476,N_428);
and U523 (N_523,N_438,N_482);
nand U524 (N_524,N_407,N_493);
or U525 (N_525,N_453,N_471);
nor U526 (N_526,N_415,N_464);
xnor U527 (N_527,N_422,N_467);
and U528 (N_528,N_439,N_466);
and U529 (N_529,N_442,N_403);
or U530 (N_530,N_478,N_412);
and U531 (N_531,N_498,N_477);
and U532 (N_532,N_470,N_444);
nor U533 (N_533,N_405,N_468);
and U534 (N_534,N_433,N_446);
and U535 (N_535,N_462,N_491);
nor U536 (N_536,N_443,N_437);
and U537 (N_537,N_496,N_485);
nand U538 (N_538,N_492,N_404);
or U539 (N_539,N_420,N_425);
or U540 (N_540,N_454,N_406);
nand U541 (N_541,N_475,N_401);
and U542 (N_542,N_414,N_489);
nor U543 (N_543,N_421,N_435);
xor U544 (N_544,N_487,N_410);
nand U545 (N_545,N_424,N_490);
and U546 (N_546,N_473,N_479);
or U547 (N_547,N_431,N_474);
xor U548 (N_548,N_455,N_413);
nand U549 (N_549,N_447,N_484);
nand U550 (N_550,N_455,N_459);
nor U551 (N_551,N_499,N_448);
nor U552 (N_552,N_415,N_474);
and U553 (N_553,N_444,N_435);
nor U554 (N_554,N_487,N_400);
and U555 (N_555,N_430,N_442);
nand U556 (N_556,N_486,N_448);
or U557 (N_557,N_422,N_448);
or U558 (N_558,N_476,N_461);
and U559 (N_559,N_415,N_493);
or U560 (N_560,N_496,N_473);
nor U561 (N_561,N_406,N_451);
nand U562 (N_562,N_456,N_463);
nand U563 (N_563,N_416,N_408);
nor U564 (N_564,N_479,N_403);
xnor U565 (N_565,N_415,N_498);
nor U566 (N_566,N_489,N_470);
or U567 (N_567,N_482,N_464);
nor U568 (N_568,N_457,N_430);
nor U569 (N_569,N_456,N_443);
or U570 (N_570,N_487,N_440);
nor U571 (N_571,N_488,N_465);
xor U572 (N_572,N_448,N_466);
or U573 (N_573,N_467,N_456);
nand U574 (N_574,N_464,N_427);
or U575 (N_575,N_412,N_471);
nor U576 (N_576,N_465,N_471);
nor U577 (N_577,N_478,N_456);
or U578 (N_578,N_462,N_494);
and U579 (N_579,N_459,N_482);
or U580 (N_580,N_481,N_473);
nor U581 (N_581,N_469,N_494);
nor U582 (N_582,N_412,N_485);
and U583 (N_583,N_421,N_481);
xnor U584 (N_584,N_450,N_409);
nor U585 (N_585,N_482,N_476);
and U586 (N_586,N_497,N_402);
and U587 (N_587,N_485,N_451);
xor U588 (N_588,N_424,N_455);
or U589 (N_589,N_434,N_493);
and U590 (N_590,N_498,N_401);
or U591 (N_591,N_424,N_461);
or U592 (N_592,N_455,N_408);
nand U593 (N_593,N_425,N_480);
and U594 (N_594,N_446,N_413);
nand U595 (N_595,N_490,N_438);
and U596 (N_596,N_429,N_462);
nand U597 (N_597,N_471,N_473);
nand U598 (N_598,N_481,N_418);
and U599 (N_599,N_453,N_403);
and U600 (N_600,N_532,N_577);
and U601 (N_601,N_592,N_528);
or U602 (N_602,N_593,N_512);
or U603 (N_603,N_522,N_527);
or U604 (N_604,N_547,N_579);
nand U605 (N_605,N_531,N_511);
nand U606 (N_606,N_545,N_541);
and U607 (N_607,N_580,N_564);
nand U608 (N_608,N_516,N_568);
and U609 (N_609,N_566,N_536);
nor U610 (N_610,N_598,N_521);
nand U611 (N_611,N_524,N_506);
nor U612 (N_612,N_576,N_507);
nand U613 (N_613,N_518,N_504);
nand U614 (N_614,N_581,N_559);
nand U615 (N_615,N_591,N_571);
nand U616 (N_616,N_570,N_597);
and U617 (N_617,N_588,N_501);
xor U618 (N_618,N_584,N_519);
or U619 (N_619,N_589,N_537);
nand U620 (N_620,N_590,N_529);
nor U621 (N_621,N_557,N_500);
and U622 (N_622,N_517,N_523);
or U623 (N_623,N_520,N_544);
xnor U624 (N_624,N_556,N_586);
nor U625 (N_625,N_554,N_572);
xnor U626 (N_626,N_546,N_569);
nor U627 (N_627,N_509,N_540);
or U628 (N_628,N_582,N_563);
nor U629 (N_629,N_560,N_533);
xnor U630 (N_630,N_567,N_508);
nor U631 (N_631,N_555,N_549);
nor U632 (N_632,N_565,N_539);
and U633 (N_633,N_550,N_548);
nand U634 (N_634,N_543,N_551);
and U635 (N_635,N_595,N_583);
nor U636 (N_636,N_530,N_526);
or U637 (N_637,N_585,N_510);
nor U638 (N_638,N_502,N_538);
or U639 (N_639,N_513,N_578);
and U640 (N_640,N_525,N_515);
and U641 (N_641,N_573,N_575);
and U642 (N_642,N_534,N_558);
and U643 (N_643,N_553,N_514);
nand U644 (N_644,N_574,N_505);
or U645 (N_645,N_535,N_561);
nand U646 (N_646,N_596,N_587);
or U647 (N_647,N_542,N_594);
nand U648 (N_648,N_503,N_552);
nor U649 (N_649,N_562,N_599);
xnor U650 (N_650,N_560,N_525);
nor U651 (N_651,N_531,N_577);
nor U652 (N_652,N_553,N_558);
and U653 (N_653,N_541,N_593);
nor U654 (N_654,N_556,N_506);
or U655 (N_655,N_583,N_505);
or U656 (N_656,N_544,N_542);
or U657 (N_657,N_508,N_537);
xnor U658 (N_658,N_520,N_552);
nand U659 (N_659,N_506,N_576);
nor U660 (N_660,N_570,N_590);
nand U661 (N_661,N_566,N_550);
and U662 (N_662,N_546,N_577);
and U663 (N_663,N_510,N_546);
xnor U664 (N_664,N_564,N_569);
and U665 (N_665,N_561,N_530);
or U666 (N_666,N_513,N_564);
and U667 (N_667,N_536,N_586);
and U668 (N_668,N_569,N_532);
and U669 (N_669,N_504,N_512);
or U670 (N_670,N_585,N_597);
and U671 (N_671,N_505,N_551);
or U672 (N_672,N_516,N_547);
nor U673 (N_673,N_563,N_588);
and U674 (N_674,N_550,N_574);
or U675 (N_675,N_551,N_564);
nor U676 (N_676,N_506,N_555);
nor U677 (N_677,N_599,N_557);
and U678 (N_678,N_597,N_579);
and U679 (N_679,N_599,N_566);
nand U680 (N_680,N_575,N_586);
or U681 (N_681,N_582,N_523);
nand U682 (N_682,N_590,N_554);
and U683 (N_683,N_570,N_553);
and U684 (N_684,N_579,N_521);
nor U685 (N_685,N_563,N_590);
xor U686 (N_686,N_583,N_525);
nor U687 (N_687,N_559,N_569);
nor U688 (N_688,N_539,N_513);
nand U689 (N_689,N_517,N_533);
nand U690 (N_690,N_578,N_512);
nand U691 (N_691,N_561,N_565);
nand U692 (N_692,N_591,N_596);
or U693 (N_693,N_514,N_583);
or U694 (N_694,N_517,N_594);
and U695 (N_695,N_565,N_540);
nand U696 (N_696,N_538,N_528);
nor U697 (N_697,N_597,N_593);
nand U698 (N_698,N_517,N_548);
nand U699 (N_699,N_524,N_528);
xor U700 (N_700,N_601,N_622);
nor U701 (N_701,N_690,N_647);
or U702 (N_702,N_648,N_632);
xor U703 (N_703,N_666,N_697);
nor U704 (N_704,N_659,N_677);
nor U705 (N_705,N_682,N_696);
or U706 (N_706,N_652,N_645);
or U707 (N_707,N_615,N_699);
and U708 (N_708,N_605,N_630);
and U709 (N_709,N_614,N_687);
nand U710 (N_710,N_635,N_619);
or U711 (N_711,N_670,N_617);
nand U712 (N_712,N_662,N_685);
nor U713 (N_713,N_644,N_608);
and U714 (N_714,N_640,N_698);
nor U715 (N_715,N_669,N_692);
and U716 (N_716,N_602,N_660);
nor U717 (N_717,N_600,N_642);
nand U718 (N_718,N_671,N_655);
and U719 (N_719,N_634,N_643);
nor U720 (N_720,N_681,N_627);
or U721 (N_721,N_695,N_689);
or U722 (N_722,N_618,N_667);
nor U723 (N_723,N_633,N_675);
and U724 (N_724,N_673,N_637);
nand U725 (N_725,N_649,N_688);
nand U726 (N_726,N_672,N_680);
xor U727 (N_727,N_631,N_621);
or U728 (N_728,N_651,N_678);
and U729 (N_729,N_656,N_603);
and U730 (N_730,N_674,N_606);
nor U731 (N_731,N_638,N_658);
or U732 (N_732,N_661,N_607);
or U733 (N_733,N_624,N_611);
or U734 (N_734,N_641,N_693);
or U735 (N_735,N_663,N_616);
nor U736 (N_736,N_626,N_664);
nand U737 (N_737,N_636,N_613);
and U738 (N_738,N_625,N_657);
nor U739 (N_739,N_604,N_679);
nand U740 (N_740,N_668,N_609);
and U741 (N_741,N_686,N_639);
nor U742 (N_742,N_628,N_646);
nand U743 (N_743,N_684,N_694);
and U744 (N_744,N_612,N_653);
or U745 (N_745,N_665,N_620);
nand U746 (N_746,N_683,N_691);
and U747 (N_747,N_654,N_610);
nand U748 (N_748,N_676,N_623);
nand U749 (N_749,N_650,N_629);
or U750 (N_750,N_683,N_696);
nand U751 (N_751,N_699,N_606);
nand U752 (N_752,N_689,N_659);
and U753 (N_753,N_678,N_626);
nand U754 (N_754,N_674,N_653);
nand U755 (N_755,N_667,N_675);
or U756 (N_756,N_630,N_645);
and U757 (N_757,N_699,N_643);
xnor U758 (N_758,N_647,N_659);
xnor U759 (N_759,N_666,N_696);
xor U760 (N_760,N_633,N_699);
or U761 (N_761,N_651,N_603);
or U762 (N_762,N_653,N_623);
nor U763 (N_763,N_661,N_664);
nor U764 (N_764,N_657,N_624);
nor U765 (N_765,N_698,N_600);
or U766 (N_766,N_628,N_632);
or U767 (N_767,N_682,N_628);
nand U768 (N_768,N_692,N_670);
nand U769 (N_769,N_622,N_602);
and U770 (N_770,N_634,N_696);
xor U771 (N_771,N_657,N_633);
nand U772 (N_772,N_650,N_633);
and U773 (N_773,N_678,N_611);
nand U774 (N_774,N_629,N_603);
or U775 (N_775,N_671,N_668);
nor U776 (N_776,N_657,N_691);
nor U777 (N_777,N_694,N_605);
xor U778 (N_778,N_621,N_660);
and U779 (N_779,N_609,N_618);
xnor U780 (N_780,N_695,N_637);
nor U781 (N_781,N_647,N_694);
xnor U782 (N_782,N_625,N_633);
nand U783 (N_783,N_663,N_617);
nor U784 (N_784,N_699,N_627);
nand U785 (N_785,N_679,N_666);
nand U786 (N_786,N_600,N_658);
nand U787 (N_787,N_615,N_641);
nand U788 (N_788,N_614,N_628);
or U789 (N_789,N_622,N_645);
nand U790 (N_790,N_640,N_675);
xnor U791 (N_791,N_662,N_699);
and U792 (N_792,N_657,N_680);
nor U793 (N_793,N_694,N_650);
nor U794 (N_794,N_680,N_606);
nor U795 (N_795,N_673,N_622);
or U796 (N_796,N_636,N_654);
and U797 (N_797,N_659,N_670);
or U798 (N_798,N_639,N_681);
and U799 (N_799,N_659,N_684);
and U800 (N_800,N_725,N_742);
and U801 (N_801,N_765,N_783);
and U802 (N_802,N_782,N_768);
and U803 (N_803,N_775,N_795);
nor U804 (N_804,N_796,N_702);
xor U805 (N_805,N_716,N_762);
or U806 (N_806,N_776,N_755);
nor U807 (N_807,N_797,N_780);
and U808 (N_808,N_781,N_772);
xor U809 (N_809,N_794,N_791);
xnor U810 (N_810,N_759,N_752);
and U811 (N_811,N_751,N_711);
and U812 (N_812,N_756,N_761);
or U813 (N_813,N_779,N_732);
xnor U814 (N_814,N_763,N_712);
xor U815 (N_815,N_731,N_786);
nor U816 (N_816,N_790,N_757);
xnor U817 (N_817,N_700,N_724);
and U818 (N_818,N_708,N_701);
and U819 (N_819,N_793,N_717);
nand U820 (N_820,N_706,N_736);
or U821 (N_821,N_789,N_746);
and U822 (N_822,N_785,N_764);
or U823 (N_823,N_720,N_713);
xnor U824 (N_824,N_715,N_743);
and U825 (N_825,N_778,N_739);
or U826 (N_826,N_766,N_745);
or U827 (N_827,N_741,N_705);
and U828 (N_828,N_728,N_758);
or U829 (N_829,N_798,N_721);
nand U830 (N_830,N_787,N_730);
and U831 (N_831,N_788,N_770);
or U832 (N_832,N_774,N_710);
nand U833 (N_833,N_723,N_773);
or U834 (N_834,N_792,N_722);
nand U835 (N_835,N_703,N_784);
nor U836 (N_836,N_734,N_718);
nor U837 (N_837,N_714,N_737);
or U838 (N_838,N_749,N_738);
nand U839 (N_839,N_748,N_733);
nand U840 (N_840,N_719,N_767);
xnor U841 (N_841,N_704,N_799);
and U842 (N_842,N_750,N_771);
and U843 (N_843,N_747,N_709);
nand U844 (N_844,N_735,N_769);
and U845 (N_845,N_740,N_727);
and U846 (N_846,N_760,N_744);
or U847 (N_847,N_777,N_754);
nor U848 (N_848,N_707,N_726);
and U849 (N_849,N_729,N_753);
and U850 (N_850,N_708,N_749);
and U851 (N_851,N_733,N_764);
and U852 (N_852,N_702,N_799);
and U853 (N_853,N_769,N_744);
and U854 (N_854,N_773,N_792);
nand U855 (N_855,N_725,N_773);
nor U856 (N_856,N_787,N_791);
nor U857 (N_857,N_710,N_789);
or U858 (N_858,N_739,N_789);
nor U859 (N_859,N_711,N_754);
nand U860 (N_860,N_798,N_795);
or U861 (N_861,N_782,N_708);
nand U862 (N_862,N_746,N_797);
nor U863 (N_863,N_709,N_799);
nor U864 (N_864,N_730,N_746);
nor U865 (N_865,N_783,N_714);
nand U866 (N_866,N_709,N_768);
or U867 (N_867,N_796,N_760);
nor U868 (N_868,N_744,N_703);
xor U869 (N_869,N_770,N_717);
and U870 (N_870,N_799,N_712);
and U871 (N_871,N_730,N_765);
and U872 (N_872,N_725,N_796);
nand U873 (N_873,N_715,N_745);
and U874 (N_874,N_775,N_733);
and U875 (N_875,N_716,N_752);
and U876 (N_876,N_760,N_700);
and U877 (N_877,N_729,N_721);
or U878 (N_878,N_754,N_700);
xnor U879 (N_879,N_734,N_727);
nand U880 (N_880,N_775,N_729);
nand U881 (N_881,N_765,N_777);
and U882 (N_882,N_758,N_789);
nor U883 (N_883,N_700,N_769);
or U884 (N_884,N_770,N_777);
or U885 (N_885,N_752,N_720);
and U886 (N_886,N_777,N_728);
and U887 (N_887,N_754,N_714);
and U888 (N_888,N_767,N_726);
and U889 (N_889,N_738,N_763);
or U890 (N_890,N_745,N_785);
and U891 (N_891,N_707,N_750);
and U892 (N_892,N_794,N_721);
nor U893 (N_893,N_762,N_704);
and U894 (N_894,N_795,N_727);
nand U895 (N_895,N_732,N_704);
or U896 (N_896,N_796,N_778);
nor U897 (N_897,N_754,N_763);
and U898 (N_898,N_711,N_730);
or U899 (N_899,N_723,N_796);
and U900 (N_900,N_843,N_897);
or U901 (N_901,N_832,N_800);
xor U902 (N_902,N_837,N_808);
nand U903 (N_903,N_831,N_867);
nand U904 (N_904,N_840,N_873);
xor U905 (N_905,N_845,N_878);
or U906 (N_906,N_821,N_883);
and U907 (N_907,N_847,N_846);
nor U908 (N_908,N_869,N_893);
nor U909 (N_909,N_899,N_852);
or U910 (N_910,N_805,N_810);
or U911 (N_911,N_851,N_857);
or U912 (N_912,N_884,N_815);
and U913 (N_913,N_894,N_870);
nand U914 (N_914,N_885,N_818);
and U915 (N_915,N_898,N_841);
nor U916 (N_916,N_813,N_892);
and U917 (N_917,N_835,N_876);
and U918 (N_918,N_887,N_820);
xor U919 (N_919,N_868,N_830);
and U920 (N_920,N_875,N_880);
xnor U921 (N_921,N_825,N_881);
nand U922 (N_922,N_838,N_849);
nor U923 (N_923,N_827,N_803);
nand U924 (N_924,N_826,N_882);
or U925 (N_925,N_824,N_864);
and U926 (N_926,N_854,N_819);
and U927 (N_927,N_848,N_823);
nand U928 (N_928,N_850,N_859);
nor U929 (N_929,N_888,N_862);
nand U930 (N_930,N_833,N_863);
or U931 (N_931,N_866,N_896);
or U932 (N_932,N_829,N_895);
and U933 (N_933,N_860,N_817);
nor U934 (N_934,N_807,N_889);
nand U935 (N_935,N_865,N_812);
nand U936 (N_936,N_855,N_836);
nand U937 (N_937,N_872,N_816);
xor U938 (N_938,N_828,N_804);
and U939 (N_939,N_886,N_839);
nand U940 (N_940,N_891,N_853);
nand U941 (N_941,N_856,N_861);
nor U942 (N_942,N_844,N_879);
nand U943 (N_943,N_811,N_822);
nor U944 (N_944,N_842,N_858);
nand U945 (N_945,N_814,N_801);
and U946 (N_946,N_890,N_802);
nand U947 (N_947,N_877,N_806);
or U948 (N_948,N_834,N_874);
xnor U949 (N_949,N_809,N_871);
nand U950 (N_950,N_827,N_895);
nor U951 (N_951,N_897,N_838);
or U952 (N_952,N_897,N_829);
nor U953 (N_953,N_837,N_821);
or U954 (N_954,N_898,N_840);
and U955 (N_955,N_881,N_807);
nor U956 (N_956,N_852,N_832);
nor U957 (N_957,N_810,N_820);
nand U958 (N_958,N_883,N_860);
and U959 (N_959,N_854,N_855);
nor U960 (N_960,N_810,N_858);
and U961 (N_961,N_874,N_864);
or U962 (N_962,N_824,N_867);
nand U963 (N_963,N_894,N_852);
nand U964 (N_964,N_870,N_812);
and U965 (N_965,N_842,N_803);
xnor U966 (N_966,N_815,N_895);
nand U967 (N_967,N_830,N_864);
and U968 (N_968,N_818,N_899);
or U969 (N_969,N_855,N_848);
nor U970 (N_970,N_804,N_856);
or U971 (N_971,N_820,N_859);
xor U972 (N_972,N_827,N_829);
nand U973 (N_973,N_806,N_887);
xnor U974 (N_974,N_861,N_807);
nor U975 (N_975,N_813,N_831);
nor U976 (N_976,N_835,N_885);
nand U977 (N_977,N_853,N_858);
nor U978 (N_978,N_835,N_859);
or U979 (N_979,N_892,N_811);
or U980 (N_980,N_867,N_833);
xor U981 (N_981,N_837,N_866);
nand U982 (N_982,N_871,N_819);
or U983 (N_983,N_888,N_829);
or U984 (N_984,N_878,N_880);
and U985 (N_985,N_873,N_848);
nor U986 (N_986,N_860,N_805);
or U987 (N_987,N_844,N_825);
or U988 (N_988,N_861,N_879);
or U989 (N_989,N_848,N_814);
nand U990 (N_990,N_853,N_808);
nor U991 (N_991,N_882,N_806);
nor U992 (N_992,N_887,N_852);
or U993 (N_993,N_843,N_831);
or U994 (N_994,N_845,N_866);
and U995 (N_995,N_820,N_830);
and U996 (N_996,N_870,N_889);
or U997 (N_997,N_845,N_838);
nand U998 (N_998,N_822,N_810);
xor U999 (N_999,N_829,N_863);
or U1000 (N_1000,N_952,N_948);
nand U1001 (N_1001,N_957,N_961);
nor U1002 (N_1002,N_930,N_927);
xor U1003 (N_1003,N_945,N_928);
or U1004 (N_1004,N_913,N_976);
nor U1005 (N_1005,N_934,N_997);
nor U1006 (N_1006,N_904,N_936);
nand U1007 (N_1007,N_993,N_964);
xor U1008 (N_1008,N_999,N_947);
and U1009 (N_1009,N_938,N_979);
nand U1010 (N_1010,N_985,N_974);
and U1011 (N_1011,N_968,N_920);
and U1012 (N_1012,N_910,N_984);
nor U1013 (N_1013,N_940,N_901);
or U1014 (N_1014,N_960,N_925);
nor U1015 (N_1015,N_944,N_983);
xnor U1016 (N_1016,N_923,N_932);
or U1017 (N_1017,N_969,N_981);
nand U1018 (N_1018,N_989,N_941);
and U1019 (N_1019,N_953,N_973);
and U1020 (N_1020,N_951,N_990);
nand U1021 (N_1021,N_905,N_980);
nor U1022 (N_1022,N_950,N_916);
and U1023 (N_1023,N_994,N_962);
nand U1024 (N_1024,N_958,N_972);
nor U1025 (N_1025,N_911,N_975);
nand U1026 (N_1026,N_986,N_917);
nor U1027 (N_1027,N_966,N_955);
and U1028 (N_1028,N_933,N_965);
and U1029 (N_1029,N_912,N_978);
nor U1030 (N_1030,N_988,N_996);
nor U1031 (N_1031,N_914,N_939);
and U1032 (N_1032,N_909,N_908);
nand U1033 (N_1033,N_924,N_942);
nand U1034 (N_1034,N_921,N_949);
or U1035 (N_1035,N_963,N_959);
or U1036 (N_1036,N_907,N_998);
and U1037 (N_1037,N_954,N_991);
nand U1038 (N_1038,N_926,N_922);
and U1039 (N_1039,N_902,N_929);
nor U1040 (N_1040,N_967,N_906);
or U1041 (N_1041,N_900,N_992);
nor U1042 (N_1042,N_956,N_995);
nand U1043 (N_1043,N_919,N_970);
nor U1044 (N_1044,N_943,N_937);
nand U1045 (N_1045,N_918,N_977);
xor U1046 (N_1046,N_946,N_903);
or U1047 (N_1047,N_931,N_987);
nand U1048 (N_1048,N_935,N_982);
and U1049 (N_1049,N_915,N_971);
and U1050 (N_1050,N_944,N_996);
nor U1051 (N_1051,N_989,N_996);
nor U1052 (N_1052,N_928,N_901);
or U1053 (N_1053,N_953,N_946);
nor U1054 (N_1054,N_936,N_927);
nor U1055 (N_1055,N_943,N_959);
nor U1056 (N_1056,N_921,N_982);
nor U1057 (N_1057,N_988,N_998);
nand U1058 (N_1058,N_998,N_983);
nand U1059 (N_1059,N_922,N_948);
and U1060 (N_1060,N_981,N_916);
nand U1061 (N_1061,N_981,N_914);
and U1062 (N_1062,N_988,N_943);
nand U1063 (N_1063,N_954,N_902);
and U1064 (N_1064,N_966,N_912);
and U1065 (N_1065,N_912,N_902);
xor U1066 (N_1066,N_900,N_966);
nand U1067 (N_1067,N_977,N_954);
nor U1068 (N_1068,N_915,N_931);
or U1069 (N_1069,N_929,N_989);
nand U1070 (N_1070,N_940,N_915);
nand U1071 (N_1071,N_985,N_960);
and U1072 (N_1072,N_970,N_978);
or U1073 (N_1073,N_939,N_965);
xnor U1074 (N_1074,N_949,N_988);
nor U1075 (N_1075,N_936,N_910);
and U1076 (N_1076,N_904,N_977);
nand U1077 (N_1077,N_973,N_931);
nand U1078 (N_1078,N_966,N_980);
and U1079 (N_1079,N_926,N_928);
nand U1080 (N_1080,N_946,N_914);
nor U1081 (N_1081,N_930,N_967);
nor U1082 (N_1082,N_980,N_937);
and U1083 (N_1083,N_985,N_970);
nand U1084 (N_1084,N_913,N_901);
xor U1085 (N_1085,N_901,N_934);
nor U1086 (N_1086,N_920,N_932);
nor U1087 (N_1087,N_938,N_942);
or U1088 (N_1088,N_964,N_980);
nor U1089 (N_1089,N_923,N_941);
nor U1090 (N_1090,N_978,N_995);
nand U1091 (N_1091,N_954,N_978);
or U1092 (N_1092,N_958,N_933);
xor U1093 (N_1093,N_970,N_931);
or U1094 (N_1094,N_907,N_968);
nor U1095 (N_1095,N_952,N_984);
nor U1096 (N_1096,N_975,N_968);
or U1097 (N_1097,N_907,N_975);
or U1098 (N_1098,N_934,N_925);
nor U1099 (N_1099,N_980,N_979);
nor U1100 (N_1100,N_1075,N_1084);
nor U1101 (N_1101,N_1078,N_1087);
and U1102 (N_1102,N_1005,N_1035);
nor U1103 (N_1103,N_1058,N_1070);
and U1104 (N_1104,N_1027,N_1095);
xnor U1105 (N_1105,N_1018,N_1000);
nand U1106 (N_1106,N_1037,N_1081);
nand U1107 (N_1107,N_1006,N_1045);
nor U1108 (N_1108,N_1029,N_1062);
and U1109 (N_1109,N_1039,N_1085);
nand U1110 (N_1110,N_1044,N_1004);
nand U1111 (N_1111,N_1022,N_1088);
nand U1112 (N_1112,N_1092,N_1046);
and U1113 (N_1113,N_1053,N_1064);
nor U1114 (N_1114,N_1051,N_1017);
nand U1115 (N_1115,N_1079,N_1003);
nor U1116 (N_1116,N_1001,N_1096);
nand U1117 (N_1117,N_1067,N_1002);
nor U1118 (N_1118,N_1089,N_1061);
and U1119 (N_1119,N_1057,N_1023);
nor U1120 (N_1120,N_1031,N_1014);
or U1121 (N_1121,N_1012,N_1050);
and U1122 (N_1122,N_1052,N_1077);
xor U1123 (N_1123,N_1097,N_1068);
or U1124 (N_1124,N_1007,N_1043);
and U1125 (N_1125,N_1069,N_1073);
and U1126 (N_1126,N_1055,N_1026);
nand U1127 (N_1127,N_1011,N_1082);
and U1128 (N_1128,N_1008,N_1091);
nand U1129 (N_1129,N_1032,N_1063);
nor U1130 (N_1130,N_1048,N_1059);
nor U1131 (N_1131,N_1083,N_1086);
and U1132 (N_1132,N_1040,N_1009);
nor U1133 (N_1133,N_1025,N_1065);
nor U1134 (N_1134,N_1080,N_1071);
or U1135 (N_1135,N_1060,N_1056);
nor U1136 (N_1136,N_1076,N_1030);
and U1137 (N_1137,N_1047,N_1024);
and U1138 (N_1138,N_1074,N_1021);
or U1139 (N_1139,N_1010,N_1072);
nor U1140 (N_1140,N_1094,N_1019);
or U1141 (N_1141,N_1098,N_1066);
xor U1142 (N_1142,N_1020,N_1016);
or U1143 (N_1143,N_1041,N_1028);
xor U1144 (N_1144,N_1038,N_1042);
or U1145 (N_1145,N_1013,N_1093);
nor U1146 (N_1146,N_1054,N_1099);
xnor U1147 (N_1147,N_1049,N_1033);
nor U1148 (N_1148,N_1036,N_1090);
nor U1149 (N_1149,N_1034,N_1015);
and U1150 (N_1150,N_1017,N_1062);
and U1151 (N_1151,N_1065,N_1004);
and U1152 (N_1152,N_1039,N_1071);
nor U1153 (N_1153,N_1020,N_1074);
or U1154 (N_1154,N_1087,N_1050);
or U1155 (N_1155,N_1074,N_1015);
and U1156 (N_1156,N_1040,N_1068);
nor U1157 (N_1157,N_1034,N_1095);
nand U1158 (N_1158,N_1092,N_1097);
nand U1159 (N_1159,N_1061,N_1054);
nor U1160 (N_1160,N_1065,N_1001);
or U1161 (N_1161,N_1048,N_1008);
and U1162 (N_1162,N_1077,N_1047);
nand U1163 (N_1163,N_1089,N_1004);
nand U1164 (N_1164,N_1011,N_1077);
xnor U1165 (N_1165,N_1052,N_1098);
or U1166 (N_1166,N_1084,N_1048);
or U1167 (N_1167,N_1029,N_1072);
and U1168 (N_1168,N_1036,N_1089);
nand U1169 (N_1169,N_1066,N_1093);
or U1170 (N_1170,N_1050,N_1042);
or U1171 (N_1171,N_1062,N_1040);
nand U1172 (N_1172,N_1038,N_1066);
nand U1173 (N_1173,N_1037,N_1096);
nand U1174 (N_1174,N_1024,N_1078);
or U1175 (N_1175,N_1088,N_1065);
nor U1176 (N_1176,N_1030,N_1054);
or U1177 (N_1177,N_1063,N_1081);
nand U1178 (N_1178,N_1026,N_1010);
nand U1179 (N_1179,N_1007,N_1058);
and U1180 (N_1180,N_1023,N_1024);
nor U1181 (N_1181,N_1040,N_1053);
or U1182 (N_1182,N_1066,N_1069);
or U1183 (N_1183,N_1027,N_1084);
or U1184 (N_1184,N_1007,N_1095);
nor U1185 (N_1185,N_1008,N_1052);
or U1186 (N_1186,N_1007,N_1098);
nand U1187 (N_1187,N_1060,N_1031);
xnor U1188 (N_1188,N_1085,N_1091);
or U1189 (N_1189,N_1035,N_1037);
or U1190 (N_1190,N_1089,N_1059);
or U1191 (N_1191,N_1049,N_1010);
nor U1192 (N_1192,N_1053,N_1006);
nor U1193 (N_1193,N_1060,N_1038);
and U1194 (N_1194,N_1045,N_1024);
nand U1195 (N_1195,N_1042,N_1029);
or U1196 (N_1196,N_1099,N_1077);
nor U1197 (N_1197,N_1014,N_1083);
nand U1198 (N_1198,N_1053,N_1044);
and U1199 (N_1199,N_1052,N_1053);
and U1200 (N_1200,N_1101,N_1196);
nand U1201 (N_1201,N_1154,N_1102);
nand U1202 (N_1202,N_1104,N_1185);
or U1203 (N_1203,N_1100,N_1126);
nand U1204 (N_1204,N_1162,N_1153);
xnor U1205 (N_1205,N_1191,N_1199);
nand U1206 (N_1206,N_1136,N_1163);
nor U1207 (N_1207,N_1134,N_1140);
or U1208 (N_1208,N_1106,N_1144);
and U1209 (N_1209,N_1143,N_1168);
and U1210 (N_1210,N_1142,N_1173);
or U1211 (N_1211,N_1108,N_1141);
nand U1212 (N_1212,N_1112,N_1186);
and U1213 (N_1213,N_1169,N_1152);
or U1214 (N_1214,N_1189,N_1149);
or U1215 (N_1215,N_1133,N_1109);
nor U1216 (N_1216,N_1182,N_1178);
nor U1217 (N_1217,N_1190,N_1113);
or U1218 (N_1218,N_1181,N_1180);
or U1219 (N_1219,N_1159,N_1161);
nand U1220 (N_1220,N_1114,N_1146);
or U1221 (N_1221,N_1179,N_1165);
or U1222 (N_1222,N_1177,N_1147);
or U1223 (N_1223,N_1117,N_1103);
nand U1224 (N_1224,N_1120,N_1145);
nor U1225 (N_1225,N_1156,N_1198);
nand U1226 (N_1226,N_1124,N_1172);
nor U1227 (N_1227,N_1166,N_1115);
nor U1228 (N_1228,N_1194,N_1192);
and U1229 (N_1229,N_1167,N_1193);
nand U1230 (N_1230,N_1131,N_1188);
or U1231 (N_1231,N_1175,N_1128);
nor U1232 (N_1232,N_1110,N_1174);
and U1233 (N_1233,N_1121,N_1127);
or U1234 (N_1234,N_1176,N_1132);
nor U1235 (N_1235,N_1118,N_1129);
nand U1236 (N_1236,N_1150,N_1105);
nor U1237 (N_1237,N_1107,N_1151);
or U1238 (N_1238,N_1187,N_1148);
and U1239 (N_1239,N_1184,N_1164);
or U1240 (N_1240,N_1155,N_1111);
and U1241 (N_1241,N_1197,N_1119);
nor U1242 (N_1242,N_1171,N_1125);
nand U1243 (N_1243,N_1135,N_1157);
nor U1244 (N_1244,N_1195,N_1160);
nor U1245 (N_1245,N_1138,N_1183);
or U1246 (N_1246,N_1139,N_1158);
nand U1247 (N_1247,N_1137,N_1123);
or U1248 (N_1248,N_1170,N_1122);
or U1249 (N_1249,N_1130,N_1116);
xor U1250 (N_1250,N_1108,N_1117);
nand U1251 (N_1251,N_1195,N_1173);
nor U1252 (N_1252,N_1122,N_1115);
nor U1253 (N_1253,N_1174,N_1152);
or U1254 (N_1254,N_1110,N_1158);
nand U1255 (N_1255,N_1162,N_1166);
and U1256 (N_1256,N_1165,N_1107);
and U1257 (N_1257,N_1134,N_1188);
and U1258 (N_1258,N_1184,N_1197);
nor U1259 (N_1259,N_1122,N_1135);
nor U1260 (N_1260,N_1168,N_1129);
nor U1261 (N_1261,N_1144,N_1195);
nor U1262 (N_1262,N_1197,N_1178);
and U1263 (N_1263,N_1193,N_1135);
and U1264 (N_1264,N_1127,N_1113);
and U1265 (N_1265,N_1129,N_1198);
xor U1266 (N_1266,N_1134,N_1110);
and U1267 (N_1267,N_1199,N_1126);
and U1268 (N_1268,N_1121,N_1164);
or U1269 (N_1269,N_1150,N_1133);
nor U1270 (N_1270,N_1125,N_1182);
nor U1271 (N_1271,N_1168,N_1184);
nor U1272 (N_1272,N_1127,N_1155);
nand U1273 (N_1273,N_1167,N_1132);
xor U1274 (N_1274,N_1167,N_1184);
nand U1275 (N_1275,N_1112,N_1145);
nand U1276 (N_1276,N_1154,N_1181);
nor U1277 (N_1277,N_1178,N_1192);
or U1278 (N_1278,N_1117,N_1159);
nor U1279 (N_1279,N_1130,N_1179);
or U1280 (N_1280,N_1122,N_1152);
xor U1281 (N_1281,N_1161,N_1166);
xnor U1282 (N_1282,N_1109,N_1103);
nor U1283 (N_1283,N_1136,N_1100);
nor U1284 (N_1284,N_1159,N_1151);
nor U1285 (N_1285,N_1160,N_1149);
or U1286 (N_1286,N_1115,N_1101);
nand U1287 (N_1287,N_1166,N_1175);
nor U1288 (N_1288,N_1137,N_1156);
or U1289 (N_1289,N_1119,N_1133);
nor U1290 (N_1290,N_1170,N_1108);
or U1291 (N_1291,N_1117,N_1140);
or U1292 (N_1292,N_1173,N_1107);
nand U1293 (N_1293,N_1138,N_1119);
nand U1294 (N_1294,N_1134,N_1113);
and U1295 (N_1295,N_1148,N_1173);
nand U1296 (N_1296,N_1193,N_1195);
nand U1297 (N_1297,N_1184,N_1130);
or U1298 (N_1298,N_1108,N_1146);
and U1299 (N_1299,N_1169,N_1121);
and U1300 (N_1300,N_1272,N_1217);
nand U1301 (N_1301,N_1255,N_1262);
xor U1302 (N_1302,N_1267,N_1282);
and U1303 (N_1303,N_1295,N_1202);
nor U1304 (N_1304,N_1248,N_1235);
nand U1305 (N_1305,N_1245,N_1208);
nor U1306 (N_1306,N_1257,N_1292);
or U1307 (N_1307,N_1274,N_1254);
or U1308 (N_1308,N_1277,N_1269);
or U1309 (N_1309,N_1243,N_1259);
nand U1310 (N_1310,N_1239,N_1279);
nor U1311 (N_1311,N_1290,N_1266);
and U1312 (N_1312,N_1224,N_1222);
and U1313 (N_1313,N_1206,N_1244);
nor U1314 (N_1314,N_1268,N_1281);
or U1315 (N_1315,N_1232,N_1297);
or U1316 (N_1316,N_1219,N_1273);
or U1317 (N_1317,N_1225,N_1241);
or U1318 (N_1318,N_1249,N_1209);
nand U1319 (N_1319,N_1201,N_1240);
nand U1320 (N_1320,N_1278,N_1253);
nor U1321 (N_1321,N_1261,N_1298);
and U1322 (N_1322,N_1215,N_1236);
and U1323 (N_1323,N_1200,N_1286);
nor U1324 (N_1324,N_1211,N_1283);
nand U1325 (N_1325,N_1263,N_1288);
nor U1326 (N_1326,N_1289,N_1284);
nor U1327 (N_1327,N_1213,N_1275);
nand U1328 (N_1328,N_1285,N_1291);
nor U1329 (N_1329,N_1231,N_1251);
nand U1330 (N_1330,N_1296,N_1246);
or U1331 (N_1331,N_1230,N_1287);
nor U1332 (N_1332,N_1205,N_1237);
xnor U1333 (N_1333,N_1229,N_1294);
nand U1334 (N_1334,N_1221,N_1260);
and U1335 (N_1335,N_1207,N_1247);
or U1336 (N_1336,N_1242,N_1218);
or U1337 (N_1337,N_1276,N_1212);
nor U1338 (N_1338,N_1252,N_1271);
nor U1339 (N_1339,N_1238,N_1293);
nand U1340 (N_1340,N_1210,N_1270);
nor U1341 (N_1341,N_1233,N_1220);
and U1342 (N_1342,N_1299,N_1226);
and U1343 (N_1343,N_1204,N_1258);
xnor U1344 (N_1344,N_1203,N_1227);
and U1345 (N_1345,N_1265,N_1223);
xnor U1346 (N_1346,N_1228,N_1280);
xor U1347 (N_1347,N_1214,N_1250);
or U1348 (N_1348,N_1234,N_1264);
or U1349 (N_1349,N_1216,N_1256);
xor U1350 (N_1350,N_1216,N_1232);
or U1351 (N_1351,N_1270,N_1231);
and U1352 (N_1352,N_1246,N_1280);
and U1353 (N_1353,N_1202,N_1225);
or U1354 (N_1354,N_1225,N_1292);
nand U1355 (N_1355,N_1293,N_1272);
nand U1356 (N_1356,N_1210,N_1220);
nor U1357 (N_1357,N_1261,N_1262);
nand U1358 (N_1358,N_1273,N_1291);
or U1359 (N_1359,N_1250,N_1288);
and U1360 (N_1360,N_1271,N_1236);
and U1361 (N_1361,N_1248,N_1270);
xor U1362 (N_1362,N_1272,N_1201);
and U1363 (N_1363,N_1252,N_1257);
nand U1364 (N_1364,N_1293,N_1224);
nor U1365 (N_1365,N_1285,N_1261);
or U1366 (N_1366,N_1248,N_1204);
nand U1367 (N_1367,N_1219,N_1214);
xnor U1368 (N_1368,N_1206,N_1274);
or U1369 (N_1369,N_1214,N_1245);
or U1370 (N_1370,N_1223,N_1229);
nand U1371 (N_1371,N_1294,N_1274);
nor U1372 (N_1372,N_1207,N_1299);
nor U1373 (N_1373,N_1291,N_1276);
or U1374 (N_1374,N_1219,N_1213);
nand U1375 (N_1375,N_1291,N_1284);
and U1376 (N_1376,N_1253,N_1205);
or U1377 (N_1377,N_1289,N_1218);
and U1378 (N_1378,N_1209,N_1288);
or U1379 (N_1379,N_1248,N_1251);
or U1380 (N_1380,N_1289,N_1226);
or U1381 (N_1381,N_1211,N_1288);
nor U1382 (N_1382,N_1243,N_1271);
and U1383 (N_1383,N_1296,N_1227);
xnor U1384 (N_1384,N_1248,N_1250);
or U1385 (N_1385,N_1249,N_1253);
nand U1386 (N_1386,N_1268,N_1236);
nor U1387 (N_1387,N_1217,N_1265);
nor U1388 (N_1388,N_1224,N_1296);
nor U1389 (N_1389,N_1203,N_1287);
and U1390 (N_1390,N_1286,N_1230);
nor U1391 (N_1391,N_1260,N_1297);
and U1392 (N_1392,N_1241,N_1291);
and U1393 (N_1393,N_1238,N_1244);
nor U1394 (N_1394,N_1200,N_1243);
nor U1395 (N_1395,N_1232,N_1264);
nor U1396 (N_1396,N_1221,N_1268);
or U1397 (N_1397,N_1254,N_1206);
nand U1398 (N_1398,N_1229,N_1299);
or U1399 (N_1399,N_1269,N_1249);
nor U1400 (N_1400,N_1349,N_1378);
xnor U1401 (N_1401,N_1352,N_1386);
nor U1402 (N_1402,N_1397,N_1337);
xor U1403 (N_1403,N_1313,N_1364);
nand U1404 (N_1404,N_1336,N_1315);
nor U1405 (N_1405,N_1310,N_1330);
nand U1406 (N_1406,N_1306,N_1318);
and U1407 (N_1407,N_1300,N_1339);
or U1408 (N_1408,N_1319,N_1320);
and U1409 (N_1409,N_1346,N_1303);
nor U1410 (N_1410,N_1371,N_1304);
and U1411 (N_1411,N_1392,N_1370);
nand U1412 (N_1412,N_1316,N_1362);
or U1413 (N_1413,N_1345,N_1343);
or U1414 (N_1414,N_1374,N_1335);
nand U1415 (N_1415,N_1368,N_1301);
xnor U1416 (N_1416,N_1327,N_1391);
or U1417 (N_1417,N_1311,N_1393);
and U1418 (N_1418,N_1317,N_1389);
nor U1419 (N_1419,N_1309,N_1353);
nor U1420 (N_1420,N_1307,N_1394);
nand U1421 (N_1421,N_1357,N_1380);
and U1422 (N_1422,N_1344,N_1385);
or U1423 (N_1423,N_1384,N_1377);
or U1424 (N_1424,N_1333,N_1338);
nand U1425 (N_1425,N_1369,N_1372);
or U1426 (N_1426,N_1373,N_1351);
nor U1427 (N_1427,N_1322,N_1350);
nor U1428 (N_1428,N_1329,N_1375);
or U1429 (N_1429,N_1324,N_1354);
nor U1430 (N_1430,N_1367,N_1321);
nand U1431 (N_1431,N_1347,N_1308);
or U1432 (N_1432,N_1331,N_1396);
or U1433 (N_1433,N_1314,N_1325);
or U1434 (N_1434,N_1382,N_1376);
nand U1435 (N_1435,N_1348,N_1388);
or U1436 (N_1436,N_1395,N_1398);
nor U1437 (N_1437,N_1399,N_1340);
and U1438 (N_1438,N_1379,N_1355);
nand U1439 (N_1439,N_1334,N_1342);
nor U1440 (N_1440,N_1383,N_1381);
nand U1441 (N_1441,N_1305,N_1323);
or U1442 (N_1442,N_1363,N_1358);
xor U1443 (N_1443,N_1390,N_1360);
and U1444 (N_1444,N_1361,N_1359);
nand U1445 (N_1445,N_1387,N_1302);
and U1446 (N_1446,N_1312,N_1328);
nand U1447 (N_1447,N_1332,N_1366);
nand U1448 (N_1448,N_1326,N_1365);
or U1449 (N_1449,N_1356,N_1341);
or U1450 (N_1450,N_1359,N_1303);
xor U1451 (N_1451,N_1300,N_1310);
nor U1452 (N_1452,N_1320,N_1337);
nand U1453 (N_1453,N_1380,N_1318);
nor U1454 (N_1454,N_1357,N_1362);
and U1455 (N_1455,N_1302,N_1345);
nand U1456 (N_1456,N_1380,N_1392);
or U1457 (N_1457,N_1395,N_1303);
nand U1458 (N_1458,N_1344,N_1373);
nor U1459 (N_1459,N_1313,N_1350);
and U1460 (N_1460,N_1376,N_1339);
nand U1461 (N_1461,N_1354,N_1383);
nand U1462 (N_1462,N_1365,N_1340);
nand U1463 (N_1463,N_1355,N_1377);
or U1464 (N_1464,N_1308,N_1341);
nor U1465 (N_1465,N_1357,N_1375);
and U1466 (N_1466,N_1336,N_1395);
and U1467 (N_1467,N_1396,N_1368);
or U1468 (N_1468,N_1350,N_1361);
nand U1469 (N_1469,N_1348,N_1381);
and U1470 (N_1470,N_1395,N_1371);
and U1471 (N_1471,N_1396,N_1336);
and U1472 (N_1472,N_1346,N_1377);
or U1473 (N_1473,N_1342,N_1362);
nand U1474 (N_1474,N_1312,N_1366);
or U1475 (N_1475,N_1324,N_1371);
xnor U1476 (N_1476,N_1303,N_1378);
or U1477 (N_1477,N_1352,N_1333);
xnor U1478 (N_1478,N_1326,N_1381);
and U1479 (N_1479,N_1336,N_1387);
and U1480 (N_1480,N_1310,N_1399);
nand U1481 (N_1481,N_1330,N_1398);
nand U1482 (N_1482,N_1363,N_1395);
and U1483 (N_1483,N_1353,N_1358);
and U1484 (N_1484,N_1312,N_1356);
xnor U1485 (N_1485,N_1359,N_1373);
nor U1486 (N_1486,N_1306,N_1391);
nor U1487 (N_1487,N_1338,N_1315);
nand U1488 (N_1488,N_1377,N_1372);
nand U1489 (N_1489,N_1306,N_1397);
nand U1490 (N_1490,N_1381,N_1363);
nand U1491 (N_1491,N_1370,N_1328);
or U1492 (N_1492,N_1345,N_1352);
nand U1493 (N_1493,N_1355,N_1373);
or U1494 (N_1494,N_1397,N_1352);
nor U1495 (N_1495,N_1322,N_1367);
or U1496 (N_1496,N_1372,N_1320);
nand U1497 (N_1497,N_1325,N_1397);
nor U1498 (N_1498,N_1380,N_1383);
or U1499 (N_1499,N_1375,N_1361);
nand U1500 (N_1500,N_1433,N_1437);
or U1501 (N_1501,N_1432,N_1489);
nand U1502 (N_1502,N_1482,N_1491);
nor U1503 (N_1503,N_1404,N_1400);
or U1504 (N_1504,N_1461,N_1454);
nor U1505 (N_1505,N_1403,N_1450);
nand U1506 (N_1506,N_1411,N_1412);
or U1507 (N_1507,N_1456,N_1441);
nor U1508 (N_1508,N_1447,N_1478);
nor U1509 (N_1509,N_1423,N_1464);
nor U1510 (N_1510,N_1414,N_1439);
nand U1511 (N_1511,N_1453,N_1446);
nand U1512 (N_1512,N_1467,N_1430);
and U1513 (N_1513,N_1420,N_1410);
and U1514 (N_1514,N_1462,N_1405);
and U1515 (N_1515,N_1497,N_1415);
xnor U1516 (N_1516,N_1426,N_1485);
and U1517 (N_1517,N_1496,N_1493);
or U1518 (N_1518,N_1477,N_1431);
and U1519 (N_1519,N_1418,N_1428);
or U1520 (N_1520,N_1492,N_1495);
and U1521 (N_1521,N_1427,N_1498);
nor U1522 (N_1522,N_1429,N_1436);
nor U1523 (N_1523,N_1448,N_1445);
nor U1524 (N_1524,N_1435,N_1480);
nand U1525 (N_1525,N_1413,N_1425);
nor U1526 (N_1526,N_1408,N_1434);
nand U1527 (N_1527,N_1468,N_1401);
nand U1528 (N_1528,N_1407,N_1490);
nand U1529 (N_1529,N_1463,N_1419);
nand U1530 (N_1530,N_1416,N_1455);
nor U1531 (N_1531,N_1488,N_1484);
and U1532 (N_1532,N_1442,N_1451);
or U1533 (N_1533,N_1470,N_1487);
xnor U1534 (N_1534,N_1460,N_1422);
or U1535 (N_1535,N_1409,N_1486);
and U1536 (N_1536,N_1402,N_1472);
or U1537 (N_1537,N_1494,N_1457);
and U1538 (N_1538,N_1465,N_1474);
and U1539 (N_1539,N_1499,N_1479);
nand U1540 (N_1540,N_1424,N_1421);
xor U1541 (N_1541,N_1469,N_1406);
or U1542 (N_1542,N_1443,N_1449);
and U1543 (N_1543,N_1475,N_1458);
nand U1544 (N_1544,N_1466,N_1440);
nand U1545 (N_1545,N_1476,N_1473);
nor U1546 (N_1546,N_1471,N_1481);
nand U1547 (N_1547,N_1452,N_1444);
nor U1548 (N_1548,N_1459,N_1438);
xnor U1549 (N_1549,N_1417,N_1483);
and U1550 (N_1550,N_1472,N_1439);
or U1551 (N_1551,N_1457,N_1439);
xnor U1552 (N_1552,N_1427,N_1453);
nor U1553 (N_1553,N_1447,N_1401);
or U1554 (N_1554,N_1412,N_1489);
nor U1555 (N_1555,N_1420,N_1426);
nand U1556 (N_1556,N_1458,N_1404);
and U1557 (N_1557,N_1485,N_1459);
xnor U1558 (N_1558,N_1438,N_1448);
or U1559 (N_1559,N_1486,N_1460);
or U1560 (N_1560,N_1496,N_1427);
and U1561 (N_1561,N_1401,N_1449);
or U1562 (N_1562,N_1447,N_1434);
nor U1563 (N_1563,N_1490,N_1444);
or U1564 (N_1564,N_1457,N_1464);
nand U1565 (N_1565,N_1425,N_1496);
and U1566 (N_1566,N_1499,N_1465);
and U1567 (N_1567,N_1431,N_1453);
and U1568 (N_1568,N_1494,N_1400);
nor U1569 (N_1569,N_1415,N_1419);
or U1570 (N_1570,N_1489,N_1410);
nand U1571 (N_1571,N_1405,N_1407);
or U1572 (N_1572,N_1454,N_1477);
xor U1573 (N_1573,N_1424,N_1447);
xor U1574 (N_1574,N_1445,N_1464);
and U1575 (N_1575,N_1451,N_1415);
and U1576 (N_1576,N_1481,N_1442);
and U1577 (N_1577,N_1496,N_1432);
nor U1578 (N_1578,N_1481,N_1429);
xor U1579 (N_1579,N_1476,N_1450);
nor U1580 (N_1580,N_1417,N_1474);
and U1581 (N_1581,N_1498,N_1438);
or U1582 (N_1582,N_1427,N_1464);
and U1583 (N_1583,N_1418,N_1437);
nor U1584 (N_1584,N_1478,N_1401);
xor U1585 (N_1585,N_1451,N_1483);
or U1586 (N_1586,N_1410,N_1424);
or U1587 (N_1587,N_1443,N_1402);
and U1588 (N_1588,N_1494,N_1469);
nor U1589 (N_1589,N_1415,N_1470);
and U1590 (N_1590,N_1478,N_1427);
nor U1591 (N_1591,N_1474,N_1435);
or U1592 (N_1592,N_1485,N_1447);
nand U1593 (N_1593,N_1486,N_1430);
or U1594 (N_1594,N_1422,N_1499);
nor U1595 (N_1595,N_1402,N_1454);
and U1596 (N_1596,N_1499,N_1497);
and U1597 (N_1597,N_1455,N_1467);
nor U1598 (N_1598,N_1411,N_1456);
nor U1599 (N_1599,N_1459,N_1489);
nand U1600 (N_1600,N_1595,N_1509);
nor U1601 (N_1601,N_1546,N_1528);
and U1602 (N_1602,N_1533,N_1559);
or U1603 (N_1603,N_1586,N_1550);
nor U1604 (N_1604,N_1554,N_1592);
nand U1605 (N_1605,N_1536,N_1585);
nand U1606 (N_1606,N_1517,N_1553);
nor U1607 (N_1607,N_1506,N_1576);
nor U1608 (N_1608,N_1565,N_1579);
and U1609 (N_1609,N_1572,N_1541);
nand U1610 (N_1610,N_1544,N_1578);
nand U1611 (N_1611,N_1501,N_1525);
xor U1612 (N_1612,N_1582,N_1551);
nor U1613 (N_1613,N_1573,N_1504);
nand U1614 (N_1614,N_1526,N_1569);
nand U1615 (N_1615,N_1512,N_1556);
nand U1616 (N_1616,N_1543,N_1558);
xnor U1617 (N_1617,N_1547,N_1584);
or U1618 (N_1618,N_1574,N_1532);
nand U1619 (N_1619,N_1599,N_1598);
xnor U1620 (N_1620,N_1587,N_1581);
and U1621 (N_1621,N_1561,N_1508);
and U1622 (N_1622,N_1571,N_1531);
and U1623 (N_1623,N_1542,N_1534);
or U1624 (N_1624,N_1557,N_1515);
nor U1625 (N_1625,N_1563,N_1514);
xnor U1626 (N_1626,N_1591,N_1503);
or U1627 (N_1627,N_1597,N_1516);
nor U1628 (N_1628,N_1540,N_1505);
nand U1629 (N_1629,N_1524,N_1596);
and U1630 (N_1630,N_1593,N_1502);
nand U1631 (N_1631,N_1535,N_1513);
xnor U1632 (N_1632,N_1538,N_1552);
and U1633 (N_1633,N_1588,N_1530);
nand U1634 (N_1634,N_1564,N_1518);
nor U1635 (N_1635,N_1583,N_1511);
or U1636 (N_1636,N_1527,N_1562);
xnor U1637 (N_1637,N_1500,N_1529);
nor U1638 (N_1638,N_1589,N_1523);
xor U1639 (N_1639,N_1580,N_1555);
nor U1640 (N_1640,N_1590,N_1539);
or U1641 (N_1641,N_1575,N_1560);
or U1642 (N_1642,N_1519,N_1521);
or U1643 (N_1643,N_1548,N_1577);
xnor U1644 (N_1644,N_1520,N_1510);
or U1645 (N_1645,N_1568,N_1567);
nor U1646 (N_1646,N_1507,N_1537);
nor U1647 (N_1647,N_1545,N_1566);
nand U1648 (N_1648,N_1522,N_1594);
or U1649 (N_1649,N_1549,N_1570);
or U1650 (N_1650,N_1546,N_1535);
and U1651 (N_1651,N_1529,N_1577);
nor U1652 (N_1652,N_1504,N_1569);
or U1653 (N_1653,N_1584,N_1546);
nand U1654 (N_1654,N_1522,N_1521);
xor U1655 (N_1655,N_1550,N_1509);
or U1656 (N_1656,N_1580,N_1527);
or U1657 (N_1657,N_1586,N_1571);
nand U1658 (N_1658,N_1553,N_1571);
nand U1659 (N_1659,N_1515,N_1565);
or U1660 (N_1660,N_1523,N_1521);
xnor U1661 (N_1661,N_1512,N_1515);
and U1662 (N_1662,N_1503,N_1527);
or U1663 (N_1663,N_1542,N_1582);
nor U1664 (N_1664,N_1515,N_1564);
xnor U1665 (N_1665,N_1591,N_1525);
and U1666 (N_1666,N_1583,N_1524);
nand U1667 (N_1667,N_1527,N_1581);
nand U1668 (N_1668,N_1553,N_1570);
or U1669 (N_1669,N_1537,N_1571);
or U1670 (N_1670,N_1528,N_1532);
nor U1671 (N_1671,N_1555,N_1546);
nand U1672 (N_1672,N_1501,N_1539);
nand U1673 (N_1673,N_1508,N_1599);
nor U1674 (N_1674,N_1591,N_1542);
or U1675 (N_1675,N_1556,N_1562);
or U1676 (N_1676,N_1567,N_1505);
or U1677 (N_1677,N_1508,N_1530);
or U1678 (N_1678,N_1553,N_1566);
nor U1679 (N_1679,N_1512,N_1551);
xnor U1680 (N_1680,N_1595,N_1598);
xor U1681 (N_1681,N_1525,N_1508);
or U1682 (N_1682,N_1596,N_1507);
and U1683 (N_1683,N_1588,N_1591);
and U1684 (N_1684,N_1500,N_1557);
nand U1685 (N_1685,N_1587,N_1528);
nand U1686 (N_1686,N_1542,N_1596);
nand U1687 (N_1687,N_1582,N_1570);
and U1688 (N_1688,N_1519,N_1574);
or U1689 (N_1689,N_1553,N_1576);
nand U1690 (N_1690,N_1536,N_1586);
nand U1691 (N_1691,N_1554,N_1501);
or U1692 (N_1692,N_1560,N_1565);
or U1693 (N_1693,N_1523,N_1581);
nand U1694 (N_1694,N_1523,N_1598);
or U1695 (N_1695,N_1563,N_1579);
and U1696 (N_1696,N_1506,N_1515);
nand U1697 (N_1697,N_1525,N_1548);
nand U1698 (N_1698,N_1597,N_1538);
nor U1699 (N_1699,N_1521,N_1589);
nor U1700 (N_1700,N_1633,N_1656);
nor U1701 (N_1701,N_1642,N_1682);
and U1702 (N_1702,N_1645,N_1665);
and U1703 (N_1703,N_1608,N_1655);
nand U1704 (N_1704,N_1688,N_1647);
xor U1705 (N_1705,N_1690,N_1664);
or U1706 (N_1706,N_1666,N_1698);
or U1707 (N_1707,N_1622,N_1681);
nand U1708 (N_1708,N_1687,N_1636);
or U1709 (N_1709,N_1610,N_1674);
nand U1710 (N_1710,N_1667,N_1683);
nor U1711 (N_1711,N_1648,N_1637);
nand U1712 (N_1712,N_1653,N_1686);
and U1713 (N_1713,N_1657,N_1654);
and U1714 (N_1714,N_1670,N_1634);
xor U1715 (N_1715,N_1615,N_1697);
nand U1716 (N_1716,N_1604,N_1617);
nor U1717 (N_1717,N_1627,N_1612);
and U1718 (N_1718,N_1659,N_1613);
xor U1719 (N_1719,N_1676,N_1631);
and U1720 (N_1720,N_1629,N_1641);
nor U1721 (N_1721,N_1603,N_1625);
nand U1722 (N_1722,N_1691,N_1621);
nand U1723 (N_1723,N_1699,N_1643);
or U1724 (N_1724,N_1669,N_1601);
nor U1725 (N_1725,N_1635,N_1600);
or U1726 (N_1726,N_1628,N_1684);
and U1727 (N_1727,N_1678,N_1668);
and U1728 (N_1728,N_1650,N_1660);
nor U1729 (N_1729,N_1694,N_1626);
or U1730 (N_1730,N_1672,N_1609);
and U1731 (N_1731,N_1618,N_1644);
nor U1732 (N_1732,N_1602,N_1677);
nand U1733 (N_1733,N_1675,N_1689);
or U1734 (N_1734,N_1692,N_1685);
or U1735 (N_1735,N_1693,N_1607);
nand U1736 (N_1736,N_1632,N_1679);
or U1737 (N_1737,N_1671,N_1646);
xor U1738 (N_1738,N_1614,N_1662);
nand U1739 (N_1739,N_1696,N_1611);
xor U1740 (N_1740,N_1658,N_1606);
or U1741 (N_1741,N_1638,N_1630);
and U1742 (N_1742,N_1640,N_1619);
and U1743 (N_1743,N_1663,N_1661);
nor U1744 (N_1744,N_1652,N_1616);
and U1745 (N_1745,N_1620,N_1605);
and U1746 (N_1746,N_1651,N_1673);
or U1747 (N_1747,N_1695,N_1680);
nor U1748 (N_1748,N_1624,N_1649);
nor U1749 (N_1749,N_1639,N_1623);
xor U1750 (N_1750,N_1618,N_1623);
or U1751 (N_1751,N_1638,N_1644);
nand U1752 (N_1752,N_1691,N_1608);
or U1753 (N_1753,N_1608,N_1601);
or U1754 (N_1754,N_1615,N_1655);
nor U1755 (N_1755,N_1673,N_1642);
and U1756 (N_1756,N_1628,N_1682);
nor U1757 (N_1757,N_1613,N_1609);
nor U1758 (N_1758,N_1601,N_1677);
or U1759 (N_1759,N_1615,N_1692);
nor U1760 (N_1760,N_1642,N_1636);
nor U1761 (N_1761,N_1638,N_1643);
nor U1762 (N_1762,N_1674,N_1642);
or U1763 (N_1763,N_1640,N_1665);
nand U1764 (N_1764,N_1675,N_1666);
nand U1765 (N_1765,N_1600,N_1684);
nor U1766 (N_1766,N_1617,N_1647);
or U1767 (N_1767,N_1660,N_1646);
xor U1768 (N_1768,N_1653,N_1623);
nand U1769 (N_1769,N_1682,N_1689);
xor U1770 (N_1770,N_1627,N_1607);
nand U1771 (N_1771,N_1638,N_1671);
or U1772 (N_1772,N_1622,N_1609);
nor U1773 (N_1773,N_1629,N_1637);
nand U1774 (N_1774,N_1652,N_1624);
nand U1775 (N_1775,N_1668,N_1632);
nand U1776 (N_1776,N_1639,N_1674);
nor U1777 (N_1777,N_1669,N_1667);
xnor U1778 (N_1778,N_1631,N_1681);
nand U1779 (N_1779,N_1683,N_1659);
and U1780 (N_1780,N_1691,N_1640);
or U1781 (N_1781,N_1634,N_1681);
and U1782 (N_1782,N_1618,N_1660);
and U1783 (N_1783,N_1693,N_1612);
nor U1784 (N_1784,N_1677,N_1664);
and U1785 (N_1785,N_1698,N_1678);
xnor U1786 (N_1786,N_1699,N_1680);
and U1787 (N_1787,N_1611,N_1668);
or U1788 (N_1788,N_1689,N_1618);
nor U1789 (N_1789,N_1627,N_1622);
nor U1790 (N_1790,N_1654,N_1651);
nor U1791 (N_1791,N_1616,N_1619);
and U1792 (N_1792,N_1606,N_1601);
or U1793 (N_1793,N_1663,N_1613);
xor U1794 (N_1794,N_1685,N_1618);
and U1795 (N_1795,N_1699,N_1605);
nor U1796 (N_1796,N_1698,N_1675);
or U1797 (N_1797,N_1624,N_1618);
and U1798 (N_1798,N_1623,N_1600);
nand U1799 (N_1799,N_1636,N_1683);
nand U1800 (N_1800,N_1726,N_1750);
and U1801 (N_1801,N_1748,N_1782);
nand U1802 (N_1802,N_1715,N_1764);
or U1803 (N_1803,N_1797,N_1701);
nand U1804 (N_1804,N_1794,N_1723);
or U1805 (N_1805,N_1777,N_1720);
nor U1806 (N_1806,N_1703,N_1725);
nand U1807 (N_1807,N_1705,N_1771);
nand U1808 (N_1808,N_1770,N_1712);
nor U1809 (N_1809,N_1758,N_1706);
nand U1810 (N_1810,N_1785,N_1742);
nand U1811 (N_1811,N_1783,N_1773);
and U1812 (N_1812,N_1713,N_1716);
and U1813 (N_1813,N_1753,N_1769);
nand U1814 (N_1814,N_1721,N_1763);
or U1815 (N_1815,N_1775,N_1700);
or U1816 (N_1816,N_1739,N_1788);
nor U1817 (N_1817,N_1728,N_1751);
nand U1818 (N_1818,N_1718,N_1732);
or U1819 (N_1819,N_1754,N_1709);
and U1820 (N_1820,N_1724,N_1734);
or U1821 (N_1821,N_1755,N_1796);
xnor U1822 (N_1822,N_1789,N_1779);
and U1823 (N_1823,N_1727,N_1743);
or U1824 (N_1824,N_1776,N_1790);
nor U1825 (N_1825,N_1799,N_1756);
or U1826 (N_1826,N_1702,N_1736);
and U1827 (N_1827,N_1745,N_1707);
or U1828 (N_1828,N_1722,N_1795);
nor U1829 (N_1829,N_1749,N_1780);
nand U1830 (N_1830,N_1738,N_1767);
nor U1831 (N_1831,N_1729,N_1778);
xnor U1832 (N_1832,N_1740,N_1744);
xnor U1833 (N_1833,N_1733,N_1747);
xor U1834 (N_1834,N_1768,N_1784);
nand U1835 (N_1835,N_1793,N_1710);
and U1836 (N_1836,N_1762,N_1792);
or U1837 (N_1837,N_1786,N_1766);
nand U1838 (N_1838,N_1772,N_1708);
and U1839 (N_1839,N_1711,N_1760);
nand U1840 (N_1840,N_1759,N_1774);
nand U1841 (N_1841,N_1730,N_1737);
or U1842 (N_1842,N_1731,N_1741);
xor U1843 (N_1843,N_1757,N_1787);
nand U1844 (N_1844,N_1735,N_1791);
nand U1845 (N_1845,N_1719,N_1752);
or U1846 (N_1846,N_1798,N_1717);
and U1847 (N_1847,N_1746,N_1714);
or U1848 (N_1848,N_1761,N_1781);
nand U1849 (N_1849,N_1765,N_1704);
and U1850 (N_1850,N_1791,N_1707);
nor U1851 (N_1851,N_1748,N_1737);
nand U1852 (N_1852,N_1742,N_1777);
nor U1853 (N_1853,N_1725,N_1772);
and U1854 (N_1854,N_1731,N_1703);
nor U1855 (N_1855,N_1749,N_1724);
nor U1856 (N_1856,N_1792,N_1735);
nor U1857 (N_1857,N_1709,N_1736);
or U1858 (N_1858,N_1739,N_1724);
nand U1859 (N_1859,N_1729,N_1728);
nor U1860 (N_1860,N_1766,N_1709);
and U1861 (N_1861,N_1704,N_1705);
or U1862 (N_1862,N_1792,N_1702);
nand U1863 (N_1863,N_1745,N_1750);
or U1864 (N_1864,N_1779,N_1718);
nand U1865 (N_1865,N_1762,N_1788);
nand U1866 (N_1866,N_1775,N_1768);
nor U1867 (N_1867,N_1724,N_1776);
nor U1868 (N_1868,N_1746,N_1752);
and U1869 (N_1869,N_1706,N_1708);
or U1870 (N_1870,N_1786,N_1704);
and U1871 (N_1871,N_1714,N_1791);
xor U1872 (N_1872,N_1761,N_1797);
nor U1873 (N_1873,N_1778,N_1763);
and U1874 (N_1874,N_1742,N_1796);
nand U1875 (N_1875,N_1703,N_1752);
nor U1876 (N_1876,N_1764,N_1755);
or U1877 (N_1877,N_1741,N_1781);
nand U1878 (N_1878,N_1714,N_1788);
and U1879 (N_1879,N_1772,N_1723);
nor U1880 (N_1880,N_1724,N_1744);
or U1881 (N_1881,N_1715,N_1787);
or U1882 (N_1882,N_1702,N_1723);
nand U1883 (N_1883,N_1780,N_1729);
nand U1884 (N_1884,N_1799,N_1782);
nand U1885 (N_1885,N_1730,N_1752);
nand U1886 (N_1886,N_1754,N_1723);
xnor U1887 (N_1887,N_1783,N_1755);
nor U1888 (N_1888,N_1797,N_1763);
nand U1889 (N_1889,N_1758,N_1713);
nor U1890 (N_1890,N_1727,N_1764);
nor U1891 (N_1891,N_1782,N_1772);
or U1892 (N_1892,N_1713,N_1717);
or U1893 (N_1893,N_1788,N_1794);
nor U1894 (N_1894,N_1708,N_1702);
nor U1895 (N_1895,N_1756,N_1786);
nand U1896 (N_1896,N_1788,N_1704);
or U1897 (N_1897,N_1748,N_1789);
or U1898 (N_1898,N_1738,N_1757);
nor U1899 (N_1899,N_1725,N_1781);
or U1900 (N_1900,N_1868,N_1815);
xor U1901 (N_1901,N_1834,N_1866);
or U1902 (N_1902,N_1895,N_1807);
nand U1903 (N_1903,N_1844,N_1862);
xnor U1904 (N_1904,N_1825,N_1829);
or U1905 (N_1905,N_1883,N_1813);
nor U1906 (N_1906,N_1877,N_1878);
nor U1907 (N_1907,N_1857,N_1850);
or U1908 (N_1908,N_1865,N_1810);
nand U1909 (N_1909,N_1809,N_1803);
nand U1910 (N_1910,N_1811,N_1884);
or U1911 (N_1911,N_1846,N_1872);
and U1912 (N_1912,N_1836,N_1882);
nor U1913 (N_1913,N_1890,N_1818);
xnor U1914 (N_1914,N_1817,N_1852);
nand U1915 (N_1915,N_1894,N_1871);
and U1916 (N_1916,N_1800,N_1860);
or U1917 (N_1917,N_1853,N_1880);
nand U1918 (N_1918,N_1845,N_1843);
or U1919 (N_1919,N_1802,N_1879);
and U1920 (N_1920,N_1864,N_1885);
nand U1921 (N_1921,N_1837,N_1826);
and U1922 (N_1922,N_1847,N_1828);
or U1923 (N_1923,N_1801,N_1840);
nand U1924 (N_1924,N_1816,N_1888);
and U1925 (N_1925,N_1806,N_1804);
nor U1926 (N_1926,N_1889,N_1869);
and U1927 (N_1927,N_1863,N_1848);
xnor U1928 (N_1928,N_1899,N_1841);
nor U1929 (N_1929,N_1896,N_1893);
and U1930 (N_1930,N_1881,N_1838);
and U1931 (N_1931,N_1856,N_1830);
or U1932 (N_1932,N_1876,N_1819);
nor U1933 (N_1933,N_1805,N_1824);
xnor U1934 (N_1934,N_1812,N_1886);
or U1935 (N_1935,N_1822,N_1842);
nand U1936 (N_1936,N_1823,N_1821);
or U1937 (N_1937,N_1898,N_1854);
and U1938 (N_1938,N_1874,N_1855);
nand U1939 (N_1939,N_1832,N_1859);
and U1940 (N_1940,N_1861,N_1858);
nor U1941 (N_1941,N_1870,N_1851);
nor U1942 (N_1942,N_1875,N_1887);
and U1943 (N_1943,N_1849,N_1808);
nand U1944 (N_1944,N_1835,N_1891);
nor U1945 (N_1945,N_1831,N_1839);
nor U1946 (N_1946,N_1814,N_1897);
nand U1947 (N_1947,N_1820,N_1867);
or U1948 (N_1948,N_1833,N_1873);
nor U1949 (N_1949,N_1892,N_1827);
and U1950 (N_1950,N_1828,N_1872);
nand U1951 (N_1951,N_1851,N_1848);
and U1952 (N_1952,N_1848,N_1833);
nand U1953 (N_1953,N_1887,N_1820);
nand U1954 (N_1954,N_1801,N_1858);
nor U1955 (N_1955,N_1839,N_1819);
or U1956 (N_1956,N_1847,N_1825);
and U1957 (N_1957,N_1833,N_1871);
nor U1958 (N_1958,N_1847,N_1812);
or U1959 (N_1959,N_1827,N_1819);
nand U1960 (N_1960,N_1816,N_1852);
nor U1961 (N_1961,N_1846,N_1869);
and U1962 (N_1962,N_1840,N_1872);
nor U1963 (N_1963,N_1842,N_1846);
nand U1964 (N_1964,N_1866,N_1867);
nand U1965 (N_1965,N_1898,N_1867);
and U1966 (N_1966,N_1824,N_1828);
or U1967 (N_1967,N_1815,N_1804);
and U1968 (N_1968,N_1899,N_1819);
and U1969 (N_1969,N_1812,N_1835);
xnor U1970 (N_1970,N_1821,N_1866);
and U1971 (N_1971,N_1894,N_1832);
and U1972 (N_1972,N_1894,N_1819);
nand U1973 (N_1973,N_1846,N_1853);
nand U1974 (N_1974,N_1897,N_1800);
nand U1975 (N_1975,N_1835,N_1832);
xnor U1976 (N_1976,N_1845,N_1893);
and U1977 (N_1977,N_1884,N_1809);
nand U1978 (N_1978,N_1840,N_1865);
and U1979 (N_1979,N_1874,N_1830);
or U1980 (N_1980,N_1877,N_1850);
nor U1981 (N_1981,N_1845,N_1873);
nand U1982 (N_1982,N_1809,N_1886);
nor U1983 (N_1983,N_1825,N_1820);
nor U1984 (N_1984,N_1836,N_1843);
nand U1985 (N_1985,N_1831,N_1871);
nor U1986 (N_1986,N_1896,N_1873);
nand U1987 (N_1987,N_1853,N_1834);
nor U1988 (N_1988,N_1844,N_1810);
and U1989 (N_1989,N_1828,N_1813);
nand U1990 (N_1990,N_1899,N_1863);
nor U1991 (N_1991,N_1873,N_1858);
nor U1992 (N_1992,N_1851,N_1895);
nor U1993 (N_1993,N_1848,N_1803);
nand U1994 (N_1994,N_1854,N_1813);
or U1995 (N_1995,N_1807,N_1812);
and U1996 (N_1996,N_1859,N_1809);
nor U1997 (N_1997,N_1878,N_1873);
nor U1998 (N_1998,N_1837,N_1817);
or U1999 (N_1999,N_1890,N_1817);
xnor U2000 (N_2000,N_1999,N_1922);
nand U2001 (N_2001,N_1988,N_1992);
nor U2002 (N_2002,N_1989,N_1972);
nor U2003 (N_2003,N_1914,N_1979);
nand U2004 (N_2004,N_1910,N_1941);
xnor U2005 (N_2005,N_1983,N_1923);
nand U2006 (N_2006,N_1926,N_1970);
and U2007 (N_2007,N_1968,N_1953);
and U2008 (N_2008,N_1948,N_1991);
or U2009 (N_2009,N_1903,N_1956);
nand U2010 (N_2010,N_1901,N_1960);
and U2011 (N_2011,N_1978,N_1977);
and U2012 (N_2012,N_1947,N_1951);
and U2013 (N_2013,N_1969,N_1950);
and U2014 (N_2014,N_1975,N_1942);
or U2015 (N_2015,N_1945,N_1974);
or U2016 (N_2016,N_1984,N_1957);
or U2017 (N_2017,N_1964,N_1936);
nor U2018 (N_2018,N_1946,N_1931);
nand U2019 (N_2019,N_1933,N_1935);
nand U2020 (N_2020,N_1996,N_1918);
nand U2021 (N_2021,N_1925,N_1963);
nand U2022 (N_2022,N_1917,N_1909);
nand U2023 (N_2023,N_1998,N_1906);
and U2024 (N_2024,N_1939,N_1920);
nor U2025 (N_2025,N_1921,N_1927);
and U2026 (N_2026,N_1961,N_1919);
and U2027 (N_2027,N_1987,N_1944);
nor U2028 (N_2028,N_1929,N_1913);
nor U2029 (N_2029,N_1905,N_1967);
nor U2030 (N_2030,N_1952,N_1932);
nand U2031 (N_2031,N_1934,N_1928);
or U2032 (N_2032,N_1966,N_1954);
nor U2033 (N_2033,N_1955,N_1980);
and U2034 (N_2034,N_1976,N_1973);
nor U2035 (N_2035,N_1908,N_1958);
xor U2036 (N_2036,N_1930,N_1962);
and U2037 (N_2037,N_1924,N_1911);
nand U2038 (N_2038,N_1915,N_1907);
or U2039 (N_2039,N_1949,N_1993);
and U2040 (N_2040,N_1943,N_1900);
nor U2041 (N_2041,N_1982,N_1995);
xor U2042 (N_2042,N_1994,N_1902);
and U2043 (N_2043,N_1959,N_1981);
nand U2044 (N_2044,N_1997,N_1912);
and U2045 (N_2045,N_1971,N_1916);
nor U2046 (N_2046,N_1965,N_1937);
nand U2047 (N_2047,N_1985,N_1940);
nor U2048 (N_2048,N_1986,N_1938);
or U2049 (N_2049,N_1990,N_1904);
nand U2050 (N_2050,N_1954,N_1978);
or U2051 (N_2051,N_1962,N_1903);
nand U2052 (N_2052,N_1998,N_1966);
and U2053 (N_2053,N_1910,N_1992);
nor U2054 (N_2054,N_1951,N_1933);
nand U2055 (N_2055,N_1936,N_1944);
and U2056 (N_2056,N_1907,N_1911);
xor U2057 (N_2057,N_1976,N_1996);
nand U2058 (N_2058,N_1934,N_1964);
or U2059 (N_2059,N_1953,N_1963);
nand U2060 (N_2060,N_1918,N_1971);
or U2061 (N_2061,N_1959,N_1960);
nor U2062 (N_2062,N_1900,N_1966);
nor U2063 (N_2063,N_1959,N_1978);
and U2064 (N_2064,N_1964,N_1922);
and U2065 (N_2065,N_1969,N_1936);
nand U2066 (N_2066,N_1902,N_1952);
nor U2067 (N_2067,N_1997,N_1951);
nand U2068 (N_2068,N_1982,N_1937);
and U2069 (N_2069,N_1994,N_1989);
nand U2070 (N_2070,N_1922,N_1921);
and U2071 (N_2071,N_1987,N_1982);
nand U2072 (N_2072,N_1948,N_1924);
or U2073 (N_2073,N_1918,N_1973);
or U2074 (N_2074,N_1957,N_1913);
nand U2075 (N_2075,N_1901,N_1970);
nor U2076 (N_2076,N_1933,N_1930);
xnor U2077 (N_2077,N_1973,N_1906);
and U2078 (N_2078,N_1963,N_1903);
or U2079 (N_2079,N_1975,N_1904);
nand U2080 (N_2080,N_1944,N_1977);
and U2081 (N_2081,N_1998,N_1928);
and U2082 (N_2082,N_1943,N_1957);
xnor U2083 (N_2083,N_1952,N_1950);
nor U2084 (N_2084,N_1964,N_1948);
or U2085 (N_2085,N_1953,N_1957);
nor U2086 (N_2086,N_1912,N_1957);
nor U2087 (N_2087,N_1919,N_1928);
nor U2088 (N_2088,N_1978,N_1917);
and U2089 (N_2089,N_1931,N_1942);
and U2090 (N_2090,N_1960,N_1904);
and U2091 (N_2091,N_1928,N_1939);
nand U2092 (N_2092,N_1926,N_1987);
xor U2093 (N_2093,N_1986,N_1902);
nand U2094 (N_2094,N_1908,N_1948);
and U2095 (N_2095,N_1922,N_1944);
nor U2096 (N_2096,N_1907,N_1925);
or U2097 (N_2097,N_1949,N_1912);
or U2098 (N_2098,N_1995,N_1911);
or U2099 (N_2099,N_1948,N_1959);
nand U2100 (N_2100,N_2021,N_2034);
or U2101 (N_2101,N_2068,N_2012);
and U2102 (N_2102,N_2072,N_2010);
xor U2103 (N_2103,N_2032,N_2038);
or U2104 (N_2104,N_2088,N_2069);
nor U2105 (N_2105,N_2023,N_2003);
nand U2106 (N_2106,N_2035,N_2043);
and U2107 (N_2107,N_2052,N_2085);
nand U2108 (N_2108,N_2095,N_2046);
nor U2109 (N_2109,N_2044,N_2029);
or U2110 (N_2110,N_2028,N_2097);
or U2111 (N_2111,N_2041,N_2013);
and U2112 (N_2112,N_2096,N_2014);
nor U2113 (N_2113,N_2080,N_2090);
nand U2114 (N_2114,N_2008,N_2048);
nor U2115 (N_2115,N_2024,N_2075);
nor U2116 (N_2116,N_2064,N_2073);
and U2117 (N_2117,N_2011,N_2063);
and U2118 (N_2118,N_2027,N_2040);
or U2119 (N_2119,N_2055,N_2066);
or U2120 (N_2120,N_2086,N_2033);
xnor U2121 (N_2121,N_2039,N_2025);
nor U2122 (N_2122,N_2049,N_2051);
or U2123 (N_2123,N_2031,N_2007);
or U2124 (N_2124,N_2001,N_2061);
or U2125 (N_2125,N_2015,N_2056);
nor U2126 (N_2126,N_2084,N_2022);
and U2127 (N_2127,N_2057,N_2037);
nor U2128 (N_2128,N_2098,N_2081);
nor U2129 (N_2129,N_2083,N_2030);
nor U2130 (N_2130,N_2006,N_2047);
and U2131 (N_2131,N_2099,N_2004);
xor U2132 (N_2132,N_2017,N_2093);
xnor U2133 (N_2133,N_2092,N_2076);
nand U2134 (N_2134,N_2070,N_2019);
or U2135 (N_2135,N_2058,N_2054);
or U2136 (N_2136,N_2005,N_2079);
nand U2137 (N_2137,N_2000,N_2078);
and U2138 (N_2138,N_2065,N_2059);
nor U2139 (N_2139,N_2091,N_2053);
nand U2140 (N_2140,N_2018,N_2089);
xnor U2141 (N_2141,N_2020,N_2077);
and U2142 (N_2142,N_2060,N_2045);
and U2143 (N_2143,N_2016,N_2050);
nand U2144 (N_2144,N_2009,N_2062);
xor U2145 (N_2145,N_2042,N_2002);
and U2146 (N_2146,N_2026,N_2074);
or U2147 (N_2147,N_2082,N_2067);
nor U2148 (N_2148,N_2087,N_2094);
nor U2149 (N_2149,N_2036,N_2071);
and U2150 (N_2150,N_2014,N_2001);
or U2151 (N_2151,N_2047,N_2091);
nand U2152 (N_2152,N_2069,N_2050);
and U2153 (N_2153,N_2073,N_2062);
nor U2154 (N_2154,N_2070,N_2089);
nand U2155 (N_2155,N_2069,N_2051);
or U2156 (N_2156,N_2045,N_2087);
xor U2157 (N_2157,N_2027,N_2028);
nor U2158 (N_2158,N_2085,N_2051);
or U2159 (N_2159,N_2023,N_2058);
and U2160 (N_2160,N_2087,N_2031);
or U2161 (N_2161,N_2006,N_2096);
and U2162 (N_2162,N_2080,N_2053);
and U2163 (N_2163,N_2085,N_2044);
xnor U2164 (N_2164,N_2077,N_2048);
or U2165 (N_2165,N_2038,N_2050);
and U2166 (N_2166,N_2060,N_2085);
and U2167 (N_2167,N_2013,N_2079);
nor U2168 (N_2168,N_2008,N_2023);
or U2169 (N_2169,N_2044,N_2063);
xor U2170 (N_2170,N_2092,N_2066);
xnor U2171 (N_2171,N_2085,N_2065);
and U2172 (N_2172,N_2059,N_2017);
nand U2173 (N_2173,N_2026,N_2053);
and U2174 (N_2174,N_2039,N_2068);
or U2175 (N_2175,N_2030,N_2063);
nor U2176 (N_2176,N_2057,N_2049);
xnor U2177 (N_2177,N_2019,N_2066);
nand U2178 (N_2178,N_2028,N_2069);
and U2179 (N_2179,N_2010,N_2031);
or U2180 (N_2180,N_2057,N_2041);
nand U2181 (N_2181,N_2000,N_2021);
and U2182 (N_2182,N_2063,N_2007);
and U2183 (N_2183,N_2001,N_2083);
xnor U2184 (N_2184,N_2086,N_2067);
nor U2185 (N_2185,N_2051,N_2010);
xor U2186 (N_2186,N_2022,N_2039);
nor U2187 (N_2187,N_2001,N_2068);
nand U2188 (N_2188,N_2067,N_2008);
and U2189 (N_2189,N_2092,N_2012);
nor U2190 (N_2190,N_2056,N_2060);
xor U2191 (N_2191,N_2098,N_2093);
and U2192 (N_2192,N_2047,N_2043);
nand U2193 (N_2193,N_2099,N_2043);
nor U2194 (N_2194,N_2059,N_2033);
and U2195 (N_2195,N_2099,N_2064);
or U2196 (N_2196,N_2029,N_2076);
or U2197 (N_2197,N_2099,N_2017);
nand U2198 (N_2198,N_2070,N_2054);
and U2199 (N_2199,N_2003,N_2024);
and U2200 (N_2200,N_2174,N_2176);
nor U2201 (N_2201,N_2157,N_2161);
nor U2202 (N_2202,N_2188,N_2185);
xor U2203 (N_2203,N_2116,N_2146);
nand U2204 (N_2204,N_2179,N_2140);
nand U2205 (N_2205,N_2149,N_2104);
nand U2206 (N_2206,N_2171,N_2180);
nand U2207 (N_2207,N_2193,N_2183);
nand U2208 (N_2208,N_2102,N_2130);
nand U2209 (N_2209,N_2173,N_2141);
or U2210 (N_2210,N_2142,N_2129);
nand U2211 (N_2211,N_2145,N_2127);
nand U2212 (N_2212,N_2167,N_2177);
xor U2213 (N_2213,N_2151,N_2162);
nand U2214 (N_2214,N_2190,N_2175);
or U2215 (N_2215,N_2160,N_2166);
or U2216 (N_2216,N_2109,N_2186);
or U2217 (N_2217,N_2100,N_2170);
nor U2218 (N_2218,N_2198,N_2103);
or U2219 (N_2219,N_2113,N_2136);
and U2220 (N_2220,N_2189,N_2119);
or U2221 (N_2221,N_2122,N_2112);
and U2222 (N_2222,N_2139,N_2137);
or U2223 (N_2223,N_2114,N_2110);
nand U2224 (N_2224,N_2111,N_2124);
nor U2225 (N_2225,N_2195,N_2148);
or U2226 (N_2226,N_2158,N_2159);
xor U2227 (N_2227,N_2164,N_2126);
nand U2228 (N_2228,N_2101,N_2165);
nor U2229 (N_2229,N_2125,N_2121);
xnor U2230 (N_2230,N_2178,N_2152);
or U2231 (N_2231,N_2144,N_2118);
or U2232 (N_2232,N_2199,N_2184);
nand U2233 (N_2233,N_2191,N_2154);
or U2234 (N_2234,N_2197,N_2172);
nor U2235 (N_2235,N_2163,N_2192);
nor U2236 (N_2236,N_2108,N_2182);
nor U2237 (N_2237,N_2168,N_2153);
or U2238 (N_2238,N_2143,N_2156);
and U2239 (N_2239,N_2107,N_2117);
or U2240 (N_2240,N_2194,N_2115);
nand U2241 (N_2241,N_2196,N_2181);
or U2242 (N_2242,N_2120,N_2105);
nand U2243 (N_2243,N_2133,N_2150);
or U2244 (N_2244,N_2138,N_2187);
and U2245 (N_2245,N_2131,N_2135);
and U2246 (N_2246,N_2106,N_2169);
xnor U2247 (N_2247,N_2123,N_2134);
nor U2248 (N_2248,N_2155,N_2128);
nor U2249 (N_2249,N_2132,N_2147);
nor U2250 (N_2250,N_2192,N_2142);
nand U2251 (N_2251,N_2111,N_2196);
or U2252 (N_2252,N_2169,N_2154);
or U2253 (N_2253,N_2101,N_2157);
or U2254 (N_2254,N_2118,N_2167);
nor U2255 (N_2255,N_2165,N_2195);
and U2256 (N_2256,N_2183,N_2135);
nor U2257 (N_2257,N_2109,N_2105);
and U2258 (N_2258,N_2166,N_2159);
or U2259 (N_2259,N_2192,N_2184);
and U2260 (N_2260,N_2107,N_2105);
nor U2261 (N_2261,N_2187,N_2146);
nand U2262 (N_2262,N_2142,N_2107);
nand U2263 (N_2263,N_2185,N_2130);
and U2264 (N_2264,N_2178,N_2136);
nand U2265 (N_2265,N_2163,N_2170);
or U2266 (N_2266,N_2100,N_2132);
nand U2267 (N_2267,N_2188,N_2191);
and U2268 (N_2268,N_2189,N_2134);
and U2269 (N_2269,N_2196,N_2112);
xor U2270 (N_2270,N_2102,N_2137);
nor U2271 (N_2271,N_2102,N_2198);
or U2272 (N_2272,N_2126,N_2177);
or U2273 (N_2273,N_2125,N_2172);
nand U2274 (N_2274,N_2155,N_2160);
xor U2275 (N_2275,N_2197,N_2104);
and U2276 (N_2276,N_2136,N_2101);
xnor U2277 (N_2277,N_2164,N_2125);
or U2278 (N_2278,N_2156,N_2103);
or U2279 (N_2279,N_2150,N_2103);
and U2280 (N_2280,N_2165,N_2188);
nor U2281 (N_2281,N_2132,N_2116);
xnor U2282 (N_2282,N_2186,N_2164);
xnor U2283 (N_2283,N_2131,N_2159);
and U2284 (N_2284,N_2105,N_2134);
nand U2285 (N_2285,N_2196,N_2141);
or U2286 (N_2286,N_2108,N_2195);
nand U2287 (N_2287,N_2153,N_2183);
nand U2288 (N_2288,N_2181,N_2151);
xor U2289 (N_2289,N_2124,N_2184);
and U2290 (N_2290,N_2157,N_2172);
or U2291 (N_2291,N_2125,N_2163);
nor U2292 (N_2292,N_2106,N_2102);
and U2293 (N_2293,N_2194,N_2111);
and U2294 (N_2294,N_2148,N_2163);
nand U2295 (N_2295,N_2135,N_2150);
and U2296 (N_2296,N_2170,N_2168);
and U2297 (N_2297,N_2183,N_2132);
nand U2298 (N_2298,N_2136,N_2169);
nand U2299 (N_2299,N_2100,N_2169);
and U2300 (N_2300,N_2274,N_2231);
nand U2301 (N_2301,N_2209,N_2288);
and U2302 (N_2302,N_2242,N_2216);
and U2303 (N_2303,N_2269,N_2237);
nor U2304 (N_2304,N_2268,N_2289);
nor U2305 (N_2305,N_2264,N_2259);
nor U2306 (N_2306,N_2282,N_2204);
nor U2307 (N_2307,N_2248,N_2260);
or U2308 (N_2308,N_2254,N_2257);
xor U2309 (N_2309,N_2244,N_2284);
and U2310 (N_2310,N_2290,N_2283);
nand U2311 (N_2311,N_2252,N_2241);
nand U2312 (N_2312,N_2281,N_2277);
nand U2313 (N_2313,N_2266,N_2263);
xor U2314 (N_2314,N_2211,N_2219);
nor U2315 (N_2315,N_2267,N_2298);
nor U2316 (N_2316,N_2234,N_2250);
and U2317 (N_2317,N_2203,N_2200);
or U2318 (N_2318,N_2224,N_2239);
xor U2319 (N_2319,N_2223,N_2275);
nor U2320 (N_2320,N_2221,N_2287);
nor U2321 (N_2321,N_2222,N_2213);
or U2322 (N_2322,N_2235,N_2273);
and U2323 (N_2323,N_2276,N_2206);
and U2324 (N_2324,N_2265,N_2225);
or U2325 (N_2325,N_2240,N_2293);
or U2326 (N_2326,N_2255,N_2279);
nor U2327 (N_2327,N_2217,N_2215);
or U2328 (N_2328,N_2280,N_2228);
or U2329 (N_2329,N_2232,N_2236);
and U2330 (N_2330,N_2262,N_2292);
or U2331 (N_2331,N_2218,N_2285);
nor U2332 (N_2332,N_2238,N_2207);
nand U2333 (N_2333,N_2261,N_2227);
nor U2334 (N_2334,N_2210,N_2296);
or U2335 (N_2335,N_2256,N_2230);
nand U2336 (N_2336,N_2251,N_2212);
and U2337 (N_2337,N_2226,N_2208);
nand U2338 (N_2338,N_2294,N_2278);
and U2339 (N_2339,N_2297,N_2214);
xor U2340 (N_2340,N_2246,N_2249);
xnor U2341 (N_2341,N_2270,N_2245);
and U2342 (N_2342,N_2299,N_2271);
or U2343 (N_2343,N_2201,N_2243);
nand U2344 (N_2344,N_2202,N_2233);
or U2345 (N_2345,N_2253,N_2286);
xor U2346 (N_2346,N_2229,N_2220);
nor U2347 (N_2347,N_2272,N_2247);
nand U2348 (N_2348,N_2205,N_2258);
nand U2349 (N_2349,N_2291,N_2295);
nor U2350 (N_2350,N_2227,N_2211);
nand U2351 (N_2351,N_2206,N_2210);
nor U2352 (N_2352,N_2280,N_2262);
or U2353 (N_2353,N_2216,N_2251);
nand U2354 (N_2354,N_2277,N_2258);
or U2355 (N_2355,N_2291,N_2242);
or U2356 (N_2356,N_2214,N_2248);
xnor U2357 (N_2357,N_2259,N_2212);
and U2358 (N_2358,N_2295,N_2210);
and U2359 (N_2359,N_2261,N_2271);
or U2360 (N_2360,N_2210,N_2230);
xnor U2361 (N_2361,N_2277,N_2230);
nor U2362 (N_2362,N_2229,N_2245);
and U2363 (N_2363,N_2282,N_2257);
nand U2364 (N_2364,N_2209,N_2240);
nor U2365 (N_2365,N_2215,N_2214);
nor U2366 (N_2366,N_2230,N_2235);
or U2367 (N_2367,N_2256,N_2284);
nor U2368 (N_2368,N_2232,N_2287);
or U2369 (N_2369,N_2281,N_2267);
and U2370 (N_2370,N_2276,N_2228);
and U2371 (N_2371,N_2285,N_2244);
and U2372 (N_2372,N_2211,N_2251);
or U2373 (N_2373,N_2218,N_2250);
or U2374 (N_2374,N_2254,N_2287);
or U2375 (N_2375,N_2286,N_2275);
xor U2376 (N_2376,N_2257,N_2278);
or U2377 (N_2377,N_2258,N_2240);
or U2378 (N_2378,N_2226,N_2203);
and U2379 (N_2379,N_2264,N_2202);
or U2380 (N_2380,N_2251,N_2238);
nand U2381 (N_2381,N_2220,N_2242);
nand U2382 (N_2382,N_2245,N_2231);
or U2383 (N_2383,N_2235,N_2269);
and U2384 (N_2384,N_2265,N_2294);
or U2385 (N_2385,N_2264,N_2223);
nand U2386 (N_2386,N_2221,N_2220);
or U2387 (N_2387,N_2262,N_2271);
nand U2388 (N_2388,N_2262,N_2252);
or U2389 (N_2389,N_2238,N_2295);
nor U2390 (N_2390,N_2281,N_2224);
or U2391 (N_2391,N_2293,N_2288);
and U2392 (N_2392,N_2213,N_2290);
and U2393 (N_2393,N_2217,N_2249);
and U2394 (N_2394,N_2288,N_2243);
or U2395 (N_2395,N_2293,N_2208);
nor U2396 (N_2396,N_2280,N_2266);
or U2397 (N_2397,N_2296,N_2281);
nor U2398 (N_2398,N_2292,N_2279);
or U2399 (N_2399,N_2260,N_2268);
xor U2400 (N_2400,N_2377,N_2334);
nor U2401 (N_2401,N_2399,N_2341);
nor U2402 (N_2402,N_2364,N_2327);
nor U2403 (N_2403,N_2389,N_2387);
and U2404 (N_2404,N_2370,N_2342);
and U2405 (N_2405,N_2324,N_2309);
or U2406 (N_2406,N_2344,N_2325);
nand U2407 (N_2407,N_2383,N_2305);
nand U2408 (N_2408,N_2393,N_2316);
or U2409 (N_2409,N_2319,N_2310);
nor U2410 (N_2410,N_2302,N_2372);
and U2411 (N_2411,N_2361,N_2363);
nor U2412 (N_2412,N_2303,N_2374);
and U2413 (N_2413,N_2378,N_2332);
nor U2414 (N_2414,N_2351,N_2340);
nand U2415 (N_2415,N_2338,N_2330);
xnor U2416 (N_2416,N_2313,N_2312);
or U2417 (N_2417,N_2376,N_2336);
and U2418 (N_2418,N_2360,N_2356);
nand U2419 (N_2419,N_2397,N_2369);
nand U2420 (N_2420,N_2354,N_2337);
and U2421 (N_2421,N_2375,N_2304);
nor U2422 (N_2422,N_2339,N_2345);
and U2423 (N_2423,N_2322,N_2315);
and U2424 (N_2424,N_2343,N_2308);
or U2425 (N_2425,N_2331,N_2385);
or U2426 (N_2426,N_2388,N_2353);
and U2427 (N_2427,N_2346,N_2366);
and U2428 (N_2428,N_2301,N_2348);
nor U2429 (N_2429,N_2384,N_2390);
nand U2430 (N_2430,N_2311,N_2371);
nand U2431 (N_2431,N_2347,N_2329);
nand U2432 (N_2432,N_2392,N_2355);
nor U2433 (N_2433,N_2395,N_2373);
or U2434 (N_2434,N_2391,N_2333);
and U2435 (N_2435,N_2359,N_2326);
and U2436 (N_2436,N_2335,N_2320);
or U2437 (N_2437,N_2367,N_2318);
nor U2438 (N_2438,N_2357,N_2380);
nand U2439 (N_2439,N_2349,N_2396);
nor U2440 (N_2440,N_2365,N_2398);
or U2441 (N_2441,N_2321,N_2368);
nand U2442 (N_2442,N_2379,N_2386);
and U2443 (N_2443,N_2323,N_2352);
nand U2444 (N_2444,N_2300,N_2317);
nand U2445 (N_2445,N_2314,N_2306);
nor U2446 (N_2446,N_2307,N_2350);
xor U2447 (N_2447,N_2358,N_2381);
nor U2448 (N_2448,N_2394,N_2362);
nand U2449 (N_2449,N_2328,N_2382);
or U2450 (N_2450,N_2396,N_2300);
xor U2451 (N_2451,N_2392,N_2380);
or U2452 (N_2452,N_2353,N_2339);
and U2453 (N_2453,N_2324,N_2369);
and U2454 (N_2454,N_2394,N_2336);
nand U2455 (N_2455,N_2319,N_2332);
nand U2456 (N_2456,N_2364,N_2332);
nand U2457 (N_2457,N_2392,N_2310);
and U2458 (N_2458,N_2315,N_2394);
and U2459 (N_2459,N_2363,N_2329);
nor U2460 (N_2460,N_2354,N_2381);
nand U2461 (N_2461,N_2363,N_2301);
nor U2462 (N_2462,N_2384,N_2341);
nand U2463 (N_2463,N_2332,N_2327);
or U2464 (N_2464,N_2310,N_2357);
xnor U2465 (N_2465,N_2372,N_2332);
and U2466 (N_2466,N_2310,N_2395);
xnor U2467 (N_2467,N_2310,N_2364);
and U2468 (N_2468,N_2399,N_2320);
nor U2469 (N_2469,N_2339,N_2337);
xor U2470 (N_2470,N_2350,N_2349);
or U2471 (N_2471,N_2394,N_2397);
or U2472 (N_2472,N_2324,N_2312);
nand U2473 (N_2473,N_2328,N_2368);
nor U2474 (N_2474,N_2338,N_2305);
nor U2475 (N_2475,N_2339,N_2348);
nand U2476 (N_2476,N_2377,N_2367);
nand U2477 (N_2477,N_2368,N_2331);
nand U2478 (N_2478,N_2318,N_2362);
and U2479 (N_2479,N_2372,N_2397);
xnor U2480 (N_2480,N_2366,N_2312);
nor U2481 (N_2481,N_2379,N_2330);
or U2482 (N_2482,N_2339,N_2364);
xnor U2483 (N_2483,N_2390,N_2321);
xnor U2484 (N_2484,N_2328,N_2313);
and U2485 (N_2485,N_2392,N_2398);
and U2486 (N_2486,N_2355,N_2380);
xnor U2487 (N_2487,N_2372,N_2304);
nand U2488 (N_2488,N_2317,N_2384);
nand U2489 (N_2489,N_2337,N_2383);
nor U2490 (N_2490,N_2304,N_2365);
or U2491 (N_2491,N_2361,N_2355);
nand U2492 (N_2492,N_2335,N_2395);
or U2493 (N_2493,N_2370,N_2396);
or U2494 (N_2494,N_2353,N_2391);
or U2495 (N_2495,N_2314,N_2362);
and U2496 (N_2496,N_2317,N_2332);
or U2497 (N_2497,N_2306,N_2302);
nor U2498 (N_2498,N_2321,N_2309);
and U2499 (N_2499,N_2386,N_2324);
xor U2500 (N_2500,N_2411,N_2483);
and U2501 (N_2501,N_2497,N_2436);
and U2502 (N_2502,N_2480,N_2410);
and U2503 (N_2503,N_2488,N_2439);
nor U2504 (N_2504,N_2407,N_2459);
xor U2505 (N_2505,N_2465,N_2491);
or U2506 (N_2506,N_2404,N_2431);
xor U2507 (N_2507,N_2433,N_2476);
nand U2508 (N_2508,N_2432,N_2425);
or U2509 (N_2509,N_2464,N_2450);
xor U2510 (N_2510,N_2468,N_2493);
nor U2511 (N_2511,N_2490,N_2400);
or U2512 (N_2512,N_2472,N_2445);
or U2513 (N_2513,N_2449,N_2451);
nor U2514 (N_2514,N_2412,N_2478);
or U2515 (N_2515,N_2440,N_2422);
and U2516 (N_2516,N_2462,N_2496);
nand U2517 (N_2517,N_2485,N_2408);
and U2518 (N_2518,N_2434,N_2437);
or U2519 (N_2519,N_2453,N_2409);
or U2520 (N_2520,N_2438,N_2481);
nor U2521 (N_2521,N_2441,N_2405);
and U2522 (N_2522,N_2401,N_2419);
or U2523 (N_2523,N_2443,N_2415);
or U2524 (N_2524,N_2423,N_2466);
nand U2525 (N_2525,N_2498,N_2428);
xnor U2526 (N_2526,N_2463,N_2458);
or U2527 (N_2527,N_2427,N_2484);
xor U2528 (N_2528,N_2435,N_2486);
nand U2529 (N_2529,N_2487,N_2489);
nand U2530 (N_2530,N_2492,N_2460);
nor U2531 (N_2531,N_2416,N_2418);
and U2532 (N_2532,N_2430,N_2421);
nor U2533 (N_2533,N_2455,N_2456);
nor U2534 (N_2534,N_2475,N_2470);
or U2535 (N_2535,N_2474,N_2426);
or U2536 (N_2536,N_2414,N_2417);
or U2537 (N_2537,N_2444,N_2403);
nor U2538 (N_2538,N_2413,N_2494);
nand U2539 (N_2539,N_2420,N_2406);
xnor U2540 (N_2540,N_2477,N_2473);
nand U2541 (N_2541,N_2479,N_2446);
or U2542 (N_2542,N_2467,N_2482);
nand U2543 (N_2543,N_2447,N_2442);
and U2544 (N_2544,N_2469,N_2424);
or U2545 (N_2545,N_2495,N_2429);
xor U2546 (N_2546,N_2499,N_2448);
and U2547 (N_2547,N_2461,N_2402);
or U2548 (N_2548,N_2452,N_2457);
or U2549 (N_2549,N_2471,N_2454);
nor U2550 (N_2550,N_2496,N_2430);
nor U2551 (N_2551,N_2472,N_2415);
xor U2552 (N_2552,N_2408,N_2483);
or U2553 (N_2553,N_2452,N_2414);
nor U2554 (N_2554,N_2445,N_2450);
xor U2555 (N_2555,N_2463,N_2437);
or U2556 (N_2556,N_2427,N_2406);
nor U2557 (N_2557,N_2491,N_2469);
xor U2558 (N_2558,N_2406,N_2405);
and U2559 (N_2559,N_2483,N_2470);
nor U2560 (N_2560,N_2405,N_2469);
and U2561 (N_2561,N_2445,N_2460);
or U2562 (N_2562,N_2408,N_2405);
and U2563 (N_2563,N_2464,N_2434);
or U2564 (N_2564,N_2468,N_2492);
and U2565 (N_2565,N_2458,N_2465);
nand U2566 (N_2566,N_2408,N_2400);
and U2567 (N_2567,N_2460,N_2444);
and U2568 (N_2568,N_2453,N_2431);
nor U2569 (N_2569,N_2486,N_2410);
and U2570 (N_2570,N_2477,N_2472);
and U2571 (N_2571,N_2484,N_2471);
nand U2572 (N_2572,N_2499,N_2401);
or U2573 (N_2573,N_2474,N_2419);
xnor U2574 (N_2574,N_2425,N_2471);
nor U2575 (N_2575,N_2481,N_2418);
and U2576 (N_2576,N_2472,N_2419);
nor U2577 (N_2577,N_2421,N_2488);
or U2578 (N_2578,N_2404,N_2474);
nand U2579 (N_2579,N_2436,N_2409);
nand U2580 (N_2580,N_2475,N_2413);
and U2581 (N_2581,N_2451,N_2431);
or U2582 (N_2582,N_2421,N_2413);
and U2583 (N_2583,N_2489,N_2474);
or U2584 (N_2584,N_2461,N_2435);
or U2585 (N_2585,N_2408,N_2498);
nor U2586 (N_2586,N_2499,N_2444);
xnor U2587 (N_2587,N_2424,N_2491);
nand U2588 (N_2588,N_2433,N_2450);
and U2589 (N_2589,N_2426,N_2465);
or U2590 (N_2590,N_2446,N_2439);
and U2591 (N_2591,N_2460,N_2413);
and U2592 (N_2592,N_2435,N_2432);
xnor U2593 (N_2593,N_2403,N_2461);
or U2594 (N_2594,N_2401,N_2415);
nand U2595 (N_2595,N_2429,N_2448);
or U2596 (N_2596,N_2408,N_2447);
nor U2597 (N_2597,N_2477,N_2496);
and U2598 (N_2598,N_2458,N_2448);
and U2599 (N_2599,N_2441,N_2453);
or U2600 (N_2600,N_2524,N_2575);
or U2601 (N_2601,N_2548,N_2580);
nor U2602 (N_2602,N_2544,N_2532);
nand U2603 (N_2603,N_2574,N_2500);
and U2604 (N_2604,N_2563,N_2516);
and U2605 (N_2605,N_2562,N_2551);
xnor U2606 (N_2606,N_2507,N_2553);
nand U2607 (N_2607,N_2505,N_2537);
nor U2608 (N_2608,N_2583,N_2528);
or U2609 (N_2609,N_2578,N_2522);
and U2610 (N_2610,N_2518,N_2565);
and U2611 (N_2611,N_2599,N_2523);
or U2612 (N_2612,N_2555,N_2536);
and U2613 (N_2613,N_2598,N_2585);
nand U2614 (N_2614,N_2590,N_2570);
or U2615 (N_2615,N_2582,N_2579);
nand U2616 (N_2616,N_2545,N_2546);
xor U2617 (N_2617,N_2514,N_2561);
or U2618 (N_2618,N_2592,N_2521);
or U2619 (N_2619,N_2557,N_2569);
and U2620 (N_2620,N_2520,N_2556);
nor U2621 (N_2621,N_2530,N_2577);
and U2622 (N_2622,N_2541,N_2510);
nand U2623 (N_2623,N_2542,N_2502);
and U2624 (N_2624,N_2572,N_2550);
nor U2625 (N_2625,N_2554,N_2534);
nand U2626 (N_2626,N_2503,N_2539);
nor U2627 (N_2627,N_2566,N_2587);
and U2628 (N_2628,N_2558,N_2581);
nand U2629 (N_2629,N_2533,N_2593);
or U2630 (N_2630,N_2538,N_2549);
and U2631 (N_2631,N_2504,N_2506);
nor U2632 (N_2632,N_2517,N_2576);
or U2633 (N_2633,N_2564,N_2595);
nand U2634 (N_2634,N_2591,N_2586);
nand U2635 (N_2635,N_2597,N_2509);
or U2636 (N_2636,N_2594,N_2535);
and U2637 (N_2637,N_2519,N_2501);
nor U2638 (N_2638,N_2552,N_2567);
and U2639 (N_2639,N_2529,N_2588);
and U2640 (N_2640,N_2508,N_2511);
nor U2641 (N_2641,N_2540,N_2515);
nand U2642 (N_2642,N_2589,N_2527);
nor U2643 (N_2643,N_2568,N_2559);
xor U2644 (N_2644,N_2525,N_2543);
nand U2645 (N_2645,N_2584,N_2596);
xor U2646 (N_2646,N_2526,N_2547);
or U2647 (N_2647,N_2512,N_2560);
or U2648 (N_2648,N_2571,N_2573);
nor U2649 (N_2649,N_2513,N_2531);
nor U2650 (N_2650,N_2563,N_2530);
nor U2651 (N_2651,N_2534,N_2581);
or U2652 (N_2652,N_2543,N_2523);
or U2653 (N_2653,N_2586,N_2508);
xor U2654 (N_2654,N_2543,N_2539);
and U2655 (N_2655,N_2521,N_2575);
nor U2656 (N_2656,N_2532,N_2586);
nor U2657 (N_2657,N_2580,N_2518);
nand U2658 (N_2658,N_2505,N_2544);
or U2659 (N_2659,N_2535,N_2530);
nand U2660 (N_2660,N_2546,N_2564);
nor U2661 (N_2661,N_2531,N_2527);
xnor U2662 (N_2662,N_2504,N_2511);
nor U2663 (N_2663,N_2550,N_2529);
and U2664 (N_2664,N_2584,N_2566);
and U2665 (N_2665,N_2530,N_2572);
nand U2666 (N_2666,N_2539,N_2554);
and U2667 (N_2667,N_2512,N_2564);
nor U2668 (N_2668,N_2537,N_2551);
nor U2669 (N_2669,N_2570,N_2569);
nor U2670 (N_2670,N_2537,N_2526);
and U2671 (N_2671,N_2586,N_2594);
or U2672 (N_2672,N_2577,N_2569);
nand U2673 (N_2673,N_2514,N_2523);
or U2674 (N_2674,N_2564,N_2539);
or U2675 (N_2675,N_2532,N_2512);
nand U2676 (N_2676,N_2551,N_2539);
xor U2677 (N_2677,N_2569,N_2560);
nand U2678 (N_2678,N_2538,N_2570);
nor U2679 (N_2679,N_2587,N_2516);
nand U2680 (N_2680,N_2526,N_2593);
and U2681 (N_2681,N_2532,N_2589);
nor U2682 (N_2682,N_2509,N_2570);
nand U2683 (N_2683,N_2578,N_2583);
nand U2684 (N_2684,N_2542,N_2579);
nand U2685 (N_2685,N_2565,N_2561);
nand U2686 (N_2686,N_2596,N_2589);
nor U2687 (N_2687,N_2569,N_2512);
nand U2688 (N_2688,N_2517,N_2531);
or U2689 (N_2689,N_2534,N_2582);
or U2690 (N_2690,N_2515,N_2577);
nor U2691 (N_2691,N_2524,N_2529);
and U2692 (N_2692,N_2590,N_2587);
xor U2693 (N_2693,N_2501,N_2566);
or U2694 (N_2694,N_2546,N_2593);
or U2695 (N_2695,N_2537,N_2506);
and U2696 (N_2696,N_2599,N_2538);
and U2697 (N_2697,N_2563,N_2550);
nor U2698 (N_2698,N_2580,N_2537);
or U2699 (N_2699,N_2584,N_2576);
or U2700 (N_2700,N_2653,N_2620);
nand U2701 (N_2701,N_2678,N_2631);
or U2702 (N_2702,N_2654,N_2696);
nand U2703 (N_2703,N_2611,N_2608);
and U2704 (N_2704,N_2605,N_2637);
nor U2705 (N_2705,N_2633,N_2616);
or U2706 (N_2706,N_2690,N_2629);
nand U2707 (N_2707,N_2622,N_2655);
nor U2708 (N_2708,N_2606,N_2679);
or U2709 (N_2709,N_2621,N_2685);
xor U2710 (N_2710,N_2649,N_2618);
or U2711 (N_2711,N_2609,N_2694);
and U2712 (N_2712,N_2610,N_2623);
nor U2713 (N_2713,N_2676,N_2689);
or U2714 (N_2714,N_2614,N_2602);
or U2715 (N_2715,N_2630,N_2645);
nand U2716 (N_2716,N_2671,N_2646);
or U2717 (N_2717,N_2699,N_2664);
and U2718 (N_2718,N_2658,N_2668);
nand U2719 (N_2719,N_2632,N_2670);
or U2720 (N_2720,N_2669,N_2652);
nand U2721 (N_2721,N_2642,N_2693);
and U2722 (N_2722,N_2661,N_2643);
nor U2723 (N_2723,N_2635,N_2682);
nor U2724 (N_2724,N_2677,N_2659);
nor U2725 (N_2725,N_2636,N_2698);
xnor U2726 (N_2726,N_2639,N_2651);
and U2727 (N_2727,N_2683,N_2684);
nor U2728 (N_2728,N_2600,N_2647);
or U2729 (N_2729,N_2673,N_2692);
nand U2730 (N_2730,N_2675,N_2624);
and U2731 (N_2731,N_2625,N_2662);
nand U2732 (N_2732,N_2648,N_2663);
and U2733 (N_2733,N_2674,N_2680);
and U2734 (N_2734,N_2681,N_2667);
nand U2735 (N_2735,N_2627,N_2672);
or U2736 (N_2736,N_2650,N_2612);
and U2737 (N_2737,N_2628,N_2656);
nand U2738 (N_2738,N_2626,N_2640);
nor U2739 (N_2739,N_2691,N_2641);
or U2740 (N_2740,N_2615,N_2603);
nor U2741 (N_2741,N_2665,N_2657);
or U2742 (N_2742,N_2686,N_2601);
or U2743 (N_2743,N_2619,N_2695);
and U2744 (N_2744,N_2697,N_2617);
nand U2745 (N_2745,N_2666,N_2687);
nor U2746 (N_2746,N_2604,N_2688);
or U2747 (N_2747,N_2607,N_2638);
xor U2748 (N_2748,N_2660,N_2634);
nand U2749 (N_2749,N_2613,N_2644);
nor U2750 (N_2750,N_2687,N_2665);
nor U2751 (N_2751,N_2690,N_2610);
or U2752 (N_2752,N_2652,N_2608);
or U2753 (N_2753,N_2605,N_2639);
nor U2754 (N_2754,N_2626,N_2647);
nand U2755 (N_2755,N_2688,N_2678);
nand U2756 (N_2756,N_2642,N_2681);
nand U2757 (N_2757,N_2638,N_2605);
and U2758 (N_2758,N_2652,N_2667);
or U2759 (N_2759,N_2698,N_2610);
nand U2760 (N_2760,N_2633,N_2672);
and U2761 (N_2761,N_2602,N_2623);
or U2762 (N_2762,N_2650,N_2655);
nor U2763 (N_2763,N_2676,N_2612);
or U2764 (N_2764,N_2647,N_2695);
or U2765 (N_2765,N_2699,N_2685);
nand U2766 (N_2766,N_2688,N_2666);
or U2767 (N_2767,N_2653,N_2664);
and U2768 (N_2768,N_2609,N_2670);
nand U2769 (N_2769,N_2633,N_2667);
and U2770 (N_2770,N_2633,N_2631);
nor U2771 (N_2771,N_2670,N_2619);
nand U2772 (N_2772,N_2689,N_2645);
nor U2773 (N_2773,N_2623,N_2656);
and U2774 (N_2774,N_2610,N_2664);
xor U2775 (N_2775,N_2634,N_2633);
nand U2776 (N_2776,N_2620,N_2683);
xnor U2777 (N_2777,N_2651,N_2672);
xnor U2778 (N_2778,N_2677,N_2636);
nand U2779 (N_2779,N_2625,N_2651);
or U2780 (N_2780,N_2636,N_2620);
nor U2781 (N_2781,N_2616,N_2672);
nor U2782 (N_2782,N_2636,N_2656);
nor U2783 (N_2783,N_2642,N_2624);
nor U2784 (N_2784,N_2604,N_2654);
nor U2785 (N_2785,N_2694,N_2686);
nor U2786 (N_2786,N_2675,N_2644);
nor U2787 (N_2787,N_2601,N_2680);
and U2788 (N_2788,N_2687,N_2652);
or U2789 (N_2789,N_2629,N_2615);
and U2790 (N_2790,N_2624,N_2647);
and U2791 (N_2791,N_2682,N_2658);
xor U2792 (N_2792,N_2648,N_2691);
nand U2793 (N_2793,N_2662,N_2692);
or U2794 (N_2794,N_2695,N_2693);
or U2795 (N_2795,N_2666,N_2644);
and U2796 (N_2796,N_2618,N_2623);
nand U2797 (N_2797,N_2602,N_2606);
or U2798 (N_2798,N_2631,N_2606);
nand U2799 (N_2799,N_2688,N_2611);
xnor U2800 (N_2800,N_2727,N_2721);
and U2801 (N_2801,N_2725,N_2761);
xor U2802 (N_2802,N_2717,N_2748);
and U2803 (N_2803,N_2787,N_2765);
xnor U2804 (N_2804,N_2710,N_2704);
and U2805 (N_2805,N_2732,N_2737);
nand U2806 (N_2806,N_2731,N_2781);
xor U2807 (N_2807,N_2712,N_2719);
or U2808 (N_2808,N_2716,N_2714);
or U2809 (N_2809,N_2715,N_2789);
nand U2810 (N_2810,N_2767,N_2792);
nor U2811 (N_2811,N_2759,N_2701);
and U2812 (N_2812,N_2744,N_2724);
or U2813 (N_2813,N_2723,N_2793);
xor U2814 (N_2814,N_2750,N_2702);
or U2815 (N_2815,N_2762,N_2764);
nand U2816 (N_2816,N_2733,N_2709);
nor U2817 (N_2817,N_2756,N_2796);
and U2818 (N_2818,N_2728,N_2747);
nor U2819 (N_2819,N_2739,N_2774);
and U2820 (N_2820,N_2779,N_2711);
nor U2821 (N_2821,N_2776,N_2726);
nor U2822 (N_2822,N_2755,N_2708);
or U2823 (N_2823,N_2768,N_2742);
or U2824 (N_2824,N_2777,N_2720);
or U2825 (N_2825,N_2770,N_2766);
nor U2826 (N_2826,N_2753,N_2741);
nor U2827 (N_2827,N_2773,N_2775);
or U2828 (N_2828,N_2740,N_2743);
and U2829 (N_2829,N_2790,N_2700);
or U2830 (N_2830,N_2706,N_2751);
and U2831 (N_2831,N_2780,N_2785);
and U2832 (N_2832,N_2799,N_2784);
nor U2833 (N_2833,N_2798,N_2795);
or U2834 (N_2834,N_2746,N_2758);
or U2835 (N_2835,N_2772,N_2749);
nor U2836 (N_2836,N_2771,N_2783);
nand U2837 (N_2837,N_2769,N_2705);
nand U2838 (N_2838,N_2797,N_2736);
or U2839 (N_2839,N_2757,N_2794);
and U2840 (N_2840,N_2734,N_2713);
xnor U2841 (N_2841,N_2778,N_2754);
and U2842 (N_2842,N_2782,N_2788);
xor U2843 (N_2843,N_2729,N_2735);
nor U2844 (N_2844,N_2763,N_2730);
or U2845 (N_2845,N_2791,N_2738);
and U2846 (N_2846,N_2760,N_2703);
or U2847 (N_2847,N_2786,N_2722);
nor U2848 (N_2848,N_2752,N_2745);
xor U2849 (N_2849,N_2707,N_2718);
or U2850 (N_2850,N_2726,N_2710);
nor U2851 (N_2851,N_2795,N_2720);
and U2852 (N_2852,N_2700,N_2769);
nor U2853 (N_2853,N_2713,N_2744);
xnor U2854 (N_2854,N_2765,N_2727);
nor U2855 (N_2855,N_2759,N_2710);
and U2856 (N_2856,N_2727,N_2717);
or U2857 (N_2857,N_2786,N_2796);
and U2858 (N_2858,N_2798,N_2727);
nand U2859 (N_2859,N_2773,N_2723);
nand U2860 (N_2860,N_2712,N_2732);
xor U2861 (N_2861,N_2777,N_2741);
nor U2862 (N_2862,N_2757,N_2732);
nor U2863 (N_2863,N_2725,N_2759);
and U2864 (N_2864,N_2771,N_2712);
or U2865 (N_2865,N_2702,N_2743);
or U2866 (N_2866,N_2785,N_2708);
or U2867 (N_2867,N_2703,N_2716);
nand U2868 (N_2868,N_2759,N_2741);
or U2869 (N_2869,N_2725,N_2775);
nor U2870 (N_2870,N_2788,N_2721);
nor U2871 (N_2871,N_2719,N_2766);
or U2872 (N_2872,N_2793,N_2709);
or U2873 (N_2873,N_2742,N_2762);
xnor U2874 (N_2874,N_2780,N_2786);
and U2875 (N_2875,N_2726,N_2730);
nor U2876 (N_2876,N_2724,N_2794);
and U2877 (N_2877,N_2707,N_2788);
xnor U2878 (N_2878,N_2723,N_2788);
nor U2879 (N_2879,N_2721,N_2780);
nor U2880 (N_2880,N_2724,N_2757);
nand U2881 (N_2881,N_2784,N_2788);
or U2882 (N_2882,N_2788,N_2798);
nor U2883 (N_2883,N_2709,N_2742);
or U2884 (N_2884,N_2711,N_2772);
or U2885 (N_2885,N_2720,N_2726);
and U2886 (N_2886,N_2729,N_2715);
xnor U2887 (N_2887,N_2705,N_2758);
and U2888 (N_2888,N_2768,N_2721);
and U2889 (N_2889,N_2710,N_2754);
and U2890 (N_2890,N_2729,N_2790);
nand U2891 (N_2891,N_2752,N_2751);
and U2892 (N_2892,N_2767,N_2785);
or U2893 (N_2893,N_2728,N_2768);
nand U2894 (N_2894,N_2775,N_2772);
nand U2895 (N_2895,N_2705,N_2763);
or U2896 (N_2896,N_2716,N_2782);
xnor U2897 (N_2897,N_2779,N_2755);
nor U2898 (N_2898,N_2773,N_2737);
and U2899 (N_2899,N_2760,N_2762);
and U2900 (N_2900,N_2883,N_2824);
nand U2901 (N_2901,N_2889,N_2815);
and U2902 (N_2902,N_2884,N_2855);
nor U2903 (N_2903,N_2891,N_2868);
nand U2904 (N_2904,N_2809,N_2801);
and U2905 (N_2905,N_2851,N_2857);
and U2906 (N_2906,N_2810,N_2817);
and U2907 (N_2907,N_2811,N_2804);
nand U2908 (N_2908,N_2877,N_2816);
and U2909 (N_2909,N_2888,N_2870);
nor U2910 (N_2910,N_2844,N_2831);
nor U2911 (N_2911,N_2875,N_2858);
nor U2912 (N_2912,N_2896,N_2886);
nor U2913 (N_2913,N_2832,N_2828);
nand U2914 (N_2914,N_2822,N_2850);
or U2915 (N_2915,N_2890,N_2820);
xnor U2916 (N_2916,N_2826,N_2893);
or U2917 (N_2917,N_2836,N_2887);
nand U2918 (N_2918,N_2814,N_2842);
nand U2919 (N_2919,N_2848,N_2846);
or U2920 (N_2920,N_2821,N_2835);
or U2921 (N_2921,N_2841,N_2833);
or U2922 (N_2922,N_2829,N_2862);
and U2923 (N_2923,N_2818,N_2894);
nand U2924 (N_2924,N_2892,N_2881);
nand U2925 (N_2925,N_2869,N_2827);
and U2926 (N_2926,N_2879,N_2880);
nor U2927 (N_2927,N_2860,N_2840);
and U2928 (N_2928,N_2839,N_2864);
xor U2929 (N_2929,N_2837,N_2806);
nor U2930 (N_2930,N_2834,N_2845);
nor U2931 (N_2931,N_2843,N_2813);
xor U2932 (N_2932,N_2853,N_2885);
and U2933 (N_2933,N_2838,N_2871);
and U2934 (N_2934,N_2866,N_2805);
or U2935 (N_2935,N_2854,N_2872);
xnor U2936 (N_2936,N_2897,N_2819);
nor U2937 (N_2937,N_2873,N_2802);
nand U2938 (N_2938,N_2859,N_2863);
or U2939 (N_2939,N_2849,N_2861);
nand U2940 (N_2940,N_2899,N_2867);
nor U2941 (N_2941,N_2878,N_2808);
or U2942 (N_2942,N_2852,N_2803);
nand U2943 (N_2943,N_2876,N_2882);
or U2944 (N_2944,N_2823,N_2856);
and U2945 (N_2945,N_2812,N_2847);
nor U2946 (N_2946,N_2898,N_2825);
nor U2947 (N_2947,N_2874,N_2865);
nor U2948 (N_2948,N_2895,N_2830);
and U2949 (N_2949,N_2800,N_2807);
and U2950 (N_2950,N_2826,N_2870);
nor U2951 (N_2951,N_2848,N_2865);
or U2952 (N_2952,N_2889,N_2829);
nor U2953 (N_2953,N_2829,N_2842);
or U2954 (N_2954,N_2838,N_2858);
nand U2955 (N_2955,N_2837,N_2823);
nand U2956 (N_2956,N_2844,N_2856);
or U2957 (N_2957,N_2836,N_2849);
or U2958 (N_2958,N_2862,N_2805);
nor U2959 (N_2959,N_2843,N_2821);
nand U2960 (N_2960,N_2859,N_2807);
and U2961 (N_2961,N_2827,N_2871);
nand U2962 (N_2962,N_2826,N_2892);
nor U2963 (N_2963,N_2870,N_2829);
and U2964 (N_2964,N_2876,N_2827);
nand U2965 (N_2965,N_2803,N_2831);
nor U2966 (N_2966,N_2807,N_2853);
nand U2967 (N_2967,N_2804,N_2842);
nor U2968 (N_2968,N_2887,N_2862);
nor U2969 (N_2969,N_2855,N_2809);
and U2970 (N_2970,N_2849,N_2880);
and U2971 (N_2971,N_2871,N_2869);
or U2972 (N_2972,N_2824,N_2891);
or U2973 (N_2973,N_2823,N_2858);
nand U2974 (N_2974,N_2817,N_2858);
and U2975 (N_2975,N_2837,N_2858);
or U2976 (N_2976,N_2855,N_2843);
nor U2977 (N_2977,N_2805,N_2895);
nand U2978 (N_2978,N_2815,N_2803);
xnor U2979 (N_2979,N_2880,N_2854);
and U2980 (N_2980,N_2883,N_2856);
or U2981 (N_2981,N_2856,N_2809);
nor U2982 (N_2982,N_2843,N_2825);
nand U2983 (N_2983,N_2819,N_2807);
or U2984 (N_2984,N_2809,N_2869);
and U2985 (N_2985,N_2837,N_2889);
nand U2986 (N_2986,N_2805,N_2887);
nor U2987 (N_2987,N_2810,N_2829);
or U2988 (N_2988,N_2873,N_2872);
nand U2989 (N_2989,N_2811,N_2861);
xor U2990 (N_2990,N_2841,N_2868);
nor U2991 (N_2991,N_2872,N_2820);
xor U2992 (N_2992,N_2845,N_2808);
nor U2993 (N_2993,N_2838,N_2872);
and U2994 (N_2994,N_2848,N_2835);
and U2995 (N_2995,N_2830,N_2816);
nand U2996 (N_2996,N_2855,N_2864);
and U2997 (N_2997,N_2879,N_2815);
nor U2998 (N_2998,N_2802,N_2814);
and U2999 (N_2999,N_2828,N_2830);
or UO_0 (O_0,N_2989,N_2977);
nand UO_1 (O_1,N_2941,N_2934);
nand UO_2 (O_2,N_2931,N_2943);
nor UO_3 (O_3,N_2998,N_2913);
nor UO_4 (O_4,N_2958,N_2927);
nand UO_5 (O_5,N_2981,N_2960);
xor UO_6 (O_6,N_2935,N_2952);
xnor UO_7 (O_7,N_2984,N_2951);
nand UO_8 (O_8,N_2922,N_2953);
and UO_9 (O_9,N_2976,N_2924);
or UO_10 (O_10,N_2962,N_2946);
or UO_11 (O_11,N_2937,N_2956);
and UO_12 (O_12,N_2972,N_2987);
nor UO_13 (O_13,N_2945,N_2965);
nand UO_14 (O_14,N_2971,N_2940);
or UO_15 (O_15,N_2993,N_2957);
xor UO_16 (O_16,N_2949,N_2904);
xnor UO_17 (O_17,N_2911,N_2955);
nand UO_18 (O_18,N_2978,N_2906);
xnor UO_19 (O_19,N_2970,N_2916);
and UO_20 (O_20,N_2933,N_2994);
or UO_21 (O_21,N_2925,N_2919);
nand UO_22 (O_22,N_2950,N_2923);
or UO_23 (O_23,N_2990,N_2918);
or UO_24 (O_24,N_2954,N_2985);
nand UO_25 (O_25,N_2920,N_2901);
or UO_26 (O_26,N_2999,N_2902);
nand UO_27 (O_27,N_2980,N_2967);
nor UO_28 (O_28,N_2926,N_2900);
or UO_29 (O_29,N_2914,N_2975);
xor UO_30 (O_30,N_2930,N_2948);
and UO_31 (O_31,N_2983,N_2974);
and UO_32 (O_32,N_2932,N_2982);
or UO_33 (O_33,N_2928,N_2905);
nor UO_34 (O_34,N_2968,N_2969);
and UO_35 (O_35,N_2907,N_2944);
nor UO_36 (O_36,N_2939,N_2979);
nand UO_37 (O_37,N_2959,N_2991);
xnor UO_38 (O_38,N_2964,N_2909);
nor UO_39 (O_39,N_2910,N_2917);
or UO_40 (O_40,N_2992,N_2961);
and UO_41 (O_41,N_2996,N_2908);
nor UO_42 (O_42,N_2915,N_2966);
and UO_43 (O_43,N_2997,N_2986);
or UO_44 (O_44,N_2912,N_2963);
and UO_45 (O_45,N_2903,N_2942);
nand UO_46 (O_46,N_2936,N_2995);
or UO_47 (O_47,N_2947,N_2929);
and UO_48 (O_48,N_2938,N_2988);
nand UO_49 (O_49,N_2973,N_2921);
nor UO_50 (O_50,N_2913,N_2958);
xnor UO_51 (O_51,N_2924,N_2953);
and UO_52 (O_52,N_2900,N_2913);
and UO_53 (O_53,N_2915,N_2985);
and UO_54 (O_54,N_2996,N_2991);
nand UO_55 (O_55,N_2919,N_2959);
nor UO_56 (O_56,N_2908,N_2918);
and UO_57 (O_57,N_2993,N_2934);
or UO_58 (O_58,N_2997,N_2995);
and UO_59 (O_59,N_2980,N_2975);
or UO_60 (O_60,N_2994,N_2901);
or UO_61 (O_61,N_2957,N_2946);
and UO_62 (O_62,N_2999,N_2935);
nor UO_63 (O_63,N_2998,N_2923);
xnor UO_64 (O_64,N_2951,N_2913);
xor UO_65 (O_65,N_2980,N_2959);
nand UO_66 (O_66,N_2927,N_2907);
or UO_67 (O_67,N_2980,N_2964);
or UO_68 (O_68,N_2937,N_2921);
and UO_69 (O_69,N_2989,N_2987);
or UO_70 (O_70,N_2968,N_2923);
and UO_71 (O_71,N_2904,N_2942);
nor UO_72 (O_72,N_2927,N_2909);
xnor UO_73 (O_73,N_2974,N_2971);
xor UO_74 (O_74,N_2977,N_2940);
and UO_75 (O_75,N_2990,N_2944);
or UO_76 (O_76,N_2941,N_2961);
and UO_77 (O_77,N_2927,N_2938);
nand UO_78 (O_78,N_2960,N_2921);
nor UO_79 (O_79,N_2920,N_2964);
nor UO_80 (O_80,N_2935,N_2994);
nand UO_81 (O_81,N_2986,N_2967);
and UO_82 (O_82,N_2993,N_2948);
xor UO_83 (O_83,N_2975,N_2990);
nor UO_84 (O_84,N_2934,N_2930);
or UO_85 (O_85,N_2977,N_2905);
and UO_86 (O_86,N_2948,N_2900);
nor UO_87 (O_87,N_2993,N_2903);
nor UO_88 (O_88,N_2959,N_2907);
nand UO_89 (O_89,N_2977,N_2986);
nand UO_90 (O_90,N_2916,N_2934);
xor UO_91 (O_91,N_2986,N_2995);
or UO_92 (O_92,N_2909,N_2902);
or UO_93 (O_93,N_2902,N_2920);
nor UO_94 (O_94,N_2988,N_2927);
or UO_95 (O_95,N_2926,N_2923);
or UO_96 (O_96,N_2919,N_2908);
and UO_97 (O_97,N_2943,N_2967);
nand UO_98 (O_98,N_2971,N_2997);
nand UO_99 (O_99,N_2949,N_2999);
nor UO_100 (O_100,N_2936,N_2973);
and UO_101 (O_101,N_2951,N_2934);
or UO_102 (O_102,N_2942,N_2962);
and UO_103 (O_103,N_2939,N_2941);
and UO_104 (O_104,N_2984,N_2986);
nor UO_105 (O_105,N_2966,N_2919);
or UO_106 (O_106,N_2937,N_2993);
and UO_107 (O_107,N_2983,N_2949);
nand UO_108 (O_108,N_2912,N_2969);
nand UO_109 (O_109,N_2931,N_2906);
nand UO_110 (O_110,N_2976,N_2965);
and UO_111 (O_111,N_2960,N_2963);
xor UO_112 (O_112,N_2945,N_2913);
nand UO_113 (O_113,N_2986,N_2947);
and UO_114 (O_114,N_2966,N_2907);
and UO_115 (O_115,N_2985,N_2959);
nand UO_116 (O_116,N_2978,N_2961);
nor UO_117 (O_117,N_2902,N_2950);
nand UO_118 (O_118,N_2929,N_2904);
or UO_119 (O_119,N_2940,N_2952);
nor UO_120 (O_120,N_2908,N_2979);
nand UO_121 (O_121,N_2960,N_2944);
nand UO_122 (O_122,N_2972,N_2990);
nor UO_123 (O_123,N_2969,N_2906);
nor UO_124 (O_124,N_2941,N_2930);
or UO_125 (O_125,N_2923,N_2904);
or UO_126 (O_126,N_2917,N_2951);
nand UO_127 (O_127,N_2979,N_2947);
xnor UO_128 (O_128,N_2934,N_2942);
or UO_129 (O_129,N_2999,N_2909);
and UO_130 (O_130,N_2917,N_2977);
xnor UO_131 (O_131,N_2941,N_2947);
and UO_132 (O_132,N_2977,N_2934);
and UO_133 (O_133,N_2936,N_2987);
nor UO_134 (O_134,N_2951,N_2963);
nor UO_135 (O_135,N_2976,N_2936);
nor UO_136 (O_136,N_2980,N_2912);
nor UO_137 (O_137,N_2997,N_2929);
nand UO_138 (O_138,N_2920,N_2995);
and UO_139 (O_139,N_2904,N_2916);
xnor UO_140 (O_140,N_2938,N_2969);
or UO_141 (O_141,N_2911,N_2942);
nand UO_142 (O_142,N_2911,N_2988);
nand UO_143 (O_143,N_2974,N_2937);
nand UO_144 (O_144,N_2999,N_2905);
nand UO_145 (O_145,N_2949,N_2909);
nor UO_146 (O_146,N_2982,N_2904);
xnor UO_147 (O_147,N_2964,N_2969);
nand UO_148 (O_148,N_2973,N_2929);
nand UO_149 (O_149,N_2996,N_2918);
and UO_150 (O_150,N_2907,N_2953);
and UO_151 (O_151,N_2903,N_2974);
and UO_152 (O_152,N_2951,N_2946);
nand UO_153 (O_153,N_2975,N_2949);
and UO_154 (O_154,N_2968,N_2921);
nor UO_155 (O_155,N_2912,N_2978);
or UO_156 (O_156,N_2980,N_2946);
nand UO_157 (O_157,N_2950,N_2916);
nor UO_158 (O_158,N_2971,N_2948);
or UO_159 (O_159,N_2900,N_2919);
and UO_160 (O_160,N_2976,N_2914);
nor UO_161 (O_161,N_2925,N_2927);
or UO_162 (O_162,N_2949,N_2925);
or UO_163 (O_163,N_2936,N_2922);
nor UO_164 (O_164,N_2943,N_2992);
xor UO_165 (O_165,N_2990,N_2966);
or UO_166 (O_166,N_2975,N_2938);
or UO_167 (O_167,N_2905,N_2945);
or UO_168 (O_168,N_2935,N_2948);
xor UO_169 (O_169,N_2965,N_2922);
nand UO_170 (O_170,N_2932,N_2974);
xor UO_171 (O_171,N_2914,N_2918);
nor UO_172 (O_172,N_2921,N_2928);
nor UO_173 (O_173,N_2994,N_2999);
xor UO_174 (O_174,N_2984,N_2918);
or UO_175 (O_175,N_2953,N_2963);
nand UO_176 (O_176,N_2995,N_2934);
nor UO_177 (O_177,N_2965,N_2990);
nor UO_178 (O_178,N_2900,N_2941);
and UO_179 (O_179,N_2934,N_2956);
and UO_180 (O_180,N_2912,N_2971);
nand UO_181 (O_181,N_2944,N_2956);
or UO_182 (O_182,N_2980,N_2987);
nand UO_183 (O_183,N_2948,N_2980);
and UO_184 (O_184,N_2903,N_2945);
xor UO_185 (O_185,N_2962,N_2969);
nor UO_186 (O_186,N_2945,N_2995);
nand UO_187 (O_187,N_2943,N_2920);
and UO_188 (O_188,N_2953,N_2935);
nand UO_189 (O_189,N_2948,N_2968);
nand UO_190 (O_190,N_2991,N_2981);
xnor UO_191 (O_191,N_2929,N_2905);
or UO_192 (O_192,N_2912,N_2923);
nor UO_193 (O_193,N_2972,N_2991);
and UO_194 (O_194,N_2914,N_2943);
xnor UO_195 (O_195,N_2905,N_2912);
nor UO_196 (O_196,N_2928,N_2951);
nor UO_197 (O_197,N_2961,N_2952);
xnor UO_198 (O_198,N_2917,N_2919);
and UO_199 (O_199,N_2957,N_2907);
or UO_200 (O_200,N_2993,N_2924);
nand UO_201 (O_201,N_2977,N_2911);
and UO_202 (O_202,N_2990,N_2931);
nor UO_203 (O_203,N_2983,N_2925);
nor UO_204 (O_204,N_2995,N_2905);
nand UO_205 (O_205,N_2987,N_2954);
and UO_206 (O_206,N_2912,N_2965);
nor UO_207 (O_207,N_2926,N_2993);
nor UO_208 (O_208,N_2935,N_2919);
xnor UO_209 (O_209,N_2959,N_2990);
nand UO_210 (O_210,N_2994,N_2981);
nand UO_211 (O_211,N_2932,N_2965);
nor UO_212 (O_212,N_2913,N_2904);
nand UO_213 (O_213,N_2972,N_2913);
nor UO_214 (O_214,N_2957,N_2948);
xnor UO_215 (O_215,N_2983,N_2912);
or UO_216 (O_216,N_2962,N_2973);
and UO_217 (O_217,N_2909,N_2956);
and UO_218 (O_218,N_2985,N_2975);
or UO_219 (O_219,N_2998,N_2994);
nor UO_220 (O_220,N_2995,N_2931);
nor UO_221 (O_221,N_2963,N_2921);
or UO_222 (O_222,N_2936,N_2946);
nor UO_223 (O_223,N_2910,N_2923);
xor UO_224 (O_224,N_2903,N_2908);
or UO_225 (O_225,N_2917,N_2950);
or UO_226 (O_226,N_2989,N_2911);
nand UO_227 (O_227,N_2991,N_2973);
nor UO_228 (O_228,N_2952,N_2991);
nor UO_229 (O_229,N_2941,N_2923);
and UO_230 (O_230,N_2939,N_2998);
or UO_231 (O_231,N_2901,N_2986);
nand UO_232 (O_232,N_2943,N_2921);
and UO_233 (O_233,N_2927,N_2999);
and UO_234 (O_234,N_2905,N_2970);
or UO_235 (O_235,N_2925,N_2909);
or UO_236 (O_236,N_2936,N_2933);
or UO_237 (O_237,N_2915,N_2998);
xor UO_238 (O_238,N_2992,N_2933);
or UO_239 (O_239,N_2908,N_2976);
or UO_240 (O_240,N_2967,N_2992);
or UO_241 (O_241,N_2990,N_2974);
and UO_242 (O_242,N_2916,N_2966);
nor UO_243 (O_243,N_2901,N_2900);
nor UO_244 (O_244,N_2928,N_2969);
nor UO_245 (O_245,N_2952,N_2969);
nand UO_246 (O_246,N_2911,N_2994);
nand UO_247 (O_247,N_2930,N_2961);
nor UO_248 (O_248,N_2942,N_2930);
and UO_249 (O_249,N_2968,N_2929);
nor UO_250 (O_250,N_2916,N_2997);
nor UO_251 (O_251,N_2931,N_2941);
nor UO_252 (O_252,N_2968,N_2930);
and UO_253 (O_253,N_2916,N_2956);
and UO_254 (O_254,N_2941,N_2987);
nor UO_255 (O_255,N_2980,N_2974);
or UO_256 (O_256,N_2965,N_2992);
xor UO_257 (O_257,N_2938,N_2913);
nor UO_258 (O_258,N_2909,N_2960);
or UO_259 (O_259,N_2980,N_2988);
nor UO_260 (O_260,N_2974,N_2967);
and UO_261 (O_261,N_2998,N_2966);
and UO_262 (O_262,N_2990,N_2980);
nor UO_263 (O_263,N_2974,N_2955);
and UO_264 (O_264,N_2940,N_2959);
nor UO_265 (O_265,N_2917,N_2966);
or UO_266 (O_266,N_2919,N_2947);
nand UO_267 (O_267,N_2973,N_2939);
and UO_268 (O_268,N_2984,N_2982);
nor UO_269 (O_269,N_2935,N_2917);
or UO_270 (O_270,N_2958,N_2986);
nor UO_271 (O_271,N_2935,N_2944);
nor UO_272 (O_272,N_2924,N_2928);
or UO_273 (O_273,N_2995,N_2942);
xor UO_274 (O_274,N_2915,N_2952);
nand UO_275 (O_275,N_2907,N_2949);
and UO_276 (O_276,N_2972,N_2984);
or UO_277 (O_277,N_2998,N_2965);
xnor UO_278 (O_278,N_2919,N_2994);
xor UO_279 (O_279,N_2991,N_2979);
nor UO_280 (O_280,N_2948,N_2982);
nand UO_281 (O_281,N_2918,N_2983);
nor UO_282 (O_282,N_2994,N_2976);
nor UO_283 (O_283,N_2974,N_2907);
or UO_284 (O_284,N_2942,N_2944);
nand UO_285 (O_285,N_2937,N_2991);
nor UO_286 (O_286,N_2948,N_2947);
and UO_287 (O_287,N_2937,N_2945);
xor UO_288 (O_288,N_2918,N_2987);
nor UO_289 (O_289,N_2937,N_2992);
and UO_290 (O_290,N_2914,N_2989);
and UO_291 (O_291,N_2933,N_2938);
nand UO_292 (O_292,N_2972,N_2932);
and UO_293 (O_293,N_2920,N_2956);
nor UO_294 (O_294,N_2973,N_2922);
or UO_295 (O_295,N_2941,N_2936);
nand UO_296 (O_296,N_2994,N_2906);
or UO_297 (O_297,N_2968,N_2943);
and UO_298 (O_298,N_2904,N_2922);
or UO_299 (O_299,N_2998,N_2927);
and UO_300 (O_300,N_2994,N_2982);
or UO_301 (O_301,N_2904,N_2992);
and UO_302 (O_302,N_2970,N_2978);
and UO_303 (O_303,N_2946,N_2955);
or UO_304 (O_304,N_2959,N_2979);
and UO_305 (O_305,N_2939,N_2981);
or UO_306 (O_306,N_2905,N_2937);
nor UO_307 (O_307,N_2902,N_2932);
or UO_308 (O_308,N_2932,N_2920);
and UO_309 (O_309,N_2978,N_2947);
xnor UO_310 (O_310,N_2915,N_2988);
xor UO_311 (O_311,N_2910,N_2938);
nor UO_312 (O_312,N_2942,N_2931);
or UO_313 (O_313,N_2987,N_2909);
nand UO_314 (O_314,N_2911,N_2954);
nor UO_315 (O_315,N_2901,N_2992);
nand UO_316 (O_316,N_2944,N_2911);
nor UO_317 (O_317,N_2903,N_2986);
nor UO_318 (O_318,N_2994,N_2918);
and UO_319 (O_319,N_2978,N_2992);
nand UO_320 (O_320,N_2943,N_2912);
xnor UO_321 (O_321,N_2975,N_2920);
xor UO_322 (O_322,N_2957,N_2970);
and UO_323 (O_323,N_2967,N_2939);
nor UO_324 (O_324,N_2932,N_2923);
xor UO_325 (O_325,N_2963,N_2979);
or UO_326 (O_326,N_2994,N_2962);
xor UO_327 (O_327,N_2931,N_2913);
nor UO_328 (O_328,N_2945,N_2979);
xnor UO_329 (O_329,N_2963,N_2967);
nand UO_330 (O_330,N_2947,N_2998);
and UO_331 (O_331,N_2990,N_2979);
nand UO_332 (O_332,N_2977,N_2954);
nand UO_333 (O_333,N_2923,N_2911);
or UO_334 (O_334,N_2992,N_2971);
and UO_335 (O_335,N_2950,N_2985);
or UO_336 (O_336,N_2927,N_2917);
and UO_337 (O_337,N_2981,N_2929);
or UO_338 (O_338,N_2916,N_2930);
and UO_339 (O_339,N_2968,N_2992);
nand UO_340 (O_340,N_2902,N_2988);
nand UO_341 (O_341,N_2912,N_2999);
and UO_342 (O_342,N_2909,N_2967);
or UO_343 (O_343,N_2937,N_2996);
and UO_344 (O_344,N_2948,N_2938);
or UO_345 (O_345,N_2935,N_2972);
nand UO_346 (O_346,N_2980,N_2982);
xor UO_347 (O_347,N_2945,N_2911);
xnor UO_348 (O_348,N_2947,N_2907);
nand UO_349 (O_349,N_2914,N_2967);
or UO_350 (O_350,N_2911,N_2919);
nand UO_351 (O_351,N_2954,N_2971);
or UO_352 (O_352,N_2998,N_2911);
nor UO_353 (O_353,N_2965,N_2970);
and UO_354 (O_354,N_2918,N_2945);
nand UO_355 (O_355,N_2981,N_2949);
nand UO_356 (O_356,N_2978,N_2972);
nand UO_357 (O_357,N_2904,N_2975);
nand UO_358 (O_358,N_2922,N_2988);
and UO_359 (O_359,N_2985,N_2986);
or UO_360 (O_360,N_2922,N_2912);
nand UO_361 (O_361,N_2996,N_2930);
nor UO_362 (O_362,N_2927,N_2937);
and UO_363 (O_363,N_2910,N_2975);
nand UO_364 (O_364,N_2940,N_2937);
nor UO_365 (O_365,N_2980,N_2924);
nand UO_366 (O_366,N_2988,N_2944);
nor UO_367 (O_367,N_2927,N_2983);
and UO_368 (O_368,N_2961,N_2940);
or UO_369 (O_369,N_2968,N_2991);
and UO_370 (O_370,N_2974,N_2961);
nor UO_371 (O_371,N_2945,N_2961);
xnor UO_372 (O_372,N_2969,N_2988);
nor UO_373 (O_373,N_2922,N_2963);
or UO_374 (O_374,N_2919,N_2906);
nor UO_375 (O_375,N_2980,N_2925);
nor UO_376 (O_376,N_2988,N_2930);
or UO_377 (O_377,N_2900,N_2966);
nand UO_378 (O_378,N_2952,N_2956);
or UO_379 (O_379,N_2972,N_2944);
xnor UO_380 (O_380,N_2950,N_2928);
and UO_381 (O_381,N_2959,N_2976);
or UO_382 (O_382,N_2936,N_2918);
or UO_383 (O_383,N_2904,N_2984);
nand UO_384 (O_384,N_2954,N_2976);
and UO_385 (O_385,N_2938,N_2957);
or UO_386 (O_386,N_2984,N_2980);
and UO_387 (O_387,N_2938,N_2992);
nor UO_388 (O_388,N_2960,N_2939);
nand UO_389 (O_389,N_2940,N_2968);
xnor UO_390 (O_390,N_2989,N_2949);
and UO_391 (O_391,N_2937,N_2987);
or UO_392 (O_392,N_2928,N_2946);
or UO_393 (O_393,N_2901,N_2937);
nor UO_394 (O_394,N_2970,N_2984);
and UO_395 (O_395,N_2998,N_2903);
nand UO_396 (O_396,N_2910,N_2914);
or UO_397 (O_397,N_2917,N_2975);
nand UO_398 (O_398,N_2908,N_2907);
nand UO_399 (O_399,N_2968,N_2946);
and UO_400 (O_400,N_2995,N_2915);
nand UO_401 (O_401,N_2919,N_2990);
and UO_402 (O_402,N_2973,N_2961);
xnor UO_403 (O_403,N_2918,N_2975);
nand UO_404 (O_404,N_2947,N_2930);
xnor UO_405 (O_405,N_2992,N_2993);
or UO_406 (O_406,N_2936,N_2942);
nor UO_407 (O_407,N_2901,N_2923);
or UO_408 (O_408,N_2904,N_2938);
nor UO_409 (O_409,N_2996,N_2913);
or UO_410 (O_410,N_2981,N_2933);
xnor UO_411 (O_411,N_2996,N_2923);
xor UO_412 (O_412,N_2902,N_2977);
nand UO_413 (O_413,N_2962,N_2911);
or UO_414 (O_414,N_2928,N_2987);
and UO_415 (O_415,N_2987,N_2935);
nand UO_416 (O_416,N_2945,N_2904);
or UO_417 (O_417,N_2969,N_2975);
xor UO_418 (O_418,N_2934,N_2963);
and UO_419 (O_419,N_2992,N_2974);
or UO_420 (O_420,N_2948,N_2966);
or UO_421 (O_421,N_2987,N_2966);
or UO_422 (O_422,N_2954,N_2916);
and UO_423 (O_423,N_2909,N_2963);
or UO_424 (O_424,N_2977,N_2981);
and UO_425 (O_425,N_2960,N_2973);
or UO_426 (O_426,N_2955,N_2934);
nand UO_427 (O_427,N_2998,N_2945);
or UO_428 (O_428,N_2961,N_2962);
or UO_429 (O_429,N_2989,N_2953);
nor UO_430 (O_430,N_2900,N_2987);
and UO_431 (O_431,N_2959,N_2987);
nand UO_432 (O_432,N_2994,N_2967);
and UO_433 (O_433,N_2991,N_2975);
and UO_434 (O_434,N_2972,N_2916);
or UO_435 (O_435,N_2929,N_2943);
nor UO_436 (O_436,N_2920,N_2906);
nor UO_437 (O_437,N_2958,N_2977);
xor UO_438 (O_438,N_2907,N_2972);
or UO_439 (O_439,N_2982,N_2945);
nor UO_440 (O_440,N_2938,N_2991);
or UO_441 (O_441,N_2951,N_2995);
and UO_442 (O_442,N_2926,N_2997);
nor UO_443 (O_443,N_2938,N_2918);
or UO_444 (O_444,N_2912,N_2934);
or UO_445 (O_445,N_2903,N_2904);
or UO_446 (O_446,N_2971,N_2962);
nand UO_447 (O_447,N_2980,N_2940);
or UO_448 (O_448,N_2921,N_2950);
nor UO_449 (O_449,N_2999,N_2944);
nor UO_450 (O_450,N_2933,N_2947);
and UO_451 (O_451,N_2941,N_2978);
nand UO_452 (O_452,N_2975,N_2966);
and UO_453 (O_453,N_2974,N_2944);
or UO_454 (O_454,N_2905,N_2908);
or UO_455 (O_455,N_2961,N_2977);
and UO_456 (O_456,N_2934,N_2978);
and UO_457 (O_457,N_2921,N_2909);
or UO_458 (O_458,N_2973,N_2975);
nand UO_459 (O_459,N_2925,N_2962);
nand UO_460 (O_460,N_2978,N_2977);
nand UO_461 (O_461,N_2912,N_2974);
or UO_462 (O_462,N_2904,N_2950);
or UO_463 (O_463,N_2937,N_2955);
nor UO_464 (O_464,N_2998,N_2980);
or UO_465 (O_465,N_2963,N_2974);
xor UO_466 (O_466,N_2910,N_2904);
nand UO_467 (O_467,N_2995,N_2947);
nand UO_468 (O_468,N_2925,N_2914);
or UO_469 (O_469,N_2922,N_2969);
nand UO_470 (O_470,N_2967,N_2997);
and UO_471 (O_471,N_2928,N_2929);
or UO_472 (O_472,N_2973,N_2932);
and UO_473 (O_473,N_2936,N_2905);
and UO_474 (O_474,N_2901,N_2967);
or UO_475 (O_475,N_2967,N_2927);
nor UO_476 (O_476,N_2913,N_2928);
or UO_477 (O_477,N_2962,N_2992);
nor UO_478 (O_478,N_2946,N_2902);
or UO_479 (O_479,N_2976,N_2972);
or UO_480 (O_480,N_2934,N_2933);
or UO_481 (O_481,N_2992,N_2905);
or UO_482 (O_482,N_2933,N_2976);
or UO_483 (O_483,N_2904,N_2967);
xnor UO_484 (O_484,N_2973,N_2926);
nand UO_485 (O_485,N_2944,N_2943);
nand UO_486 (O_486,N_2924,N_2942);
nand UO_487 (O_487,N_2970,N_2954);
nor UO_488 (O_488,N_2931,N_2932);
nand UO_489 (O_489,N_2996,N_2992);
nand UO_490 (O_490,N_2986,N_2923);
or UO_491 (O_491,N_2975,N_2905);
xor UO_492 (O_492,N_2975,N_2907);
nand UO_493 (O_493,N_2977,N_2928);
xnor UO_494 (O_494,N_2987,N_2911);
and UO_495 (O_495,N_2925,N_2907);
nor UO_496 (O_496,N_2973,N_2971);
nor UO_497 (O_497,N_2926,N_2940);
nand UO_498 (O_498,N_2987,N_2985);
nor UO_499 (O_499,N_2945,N_2957);
endmodule