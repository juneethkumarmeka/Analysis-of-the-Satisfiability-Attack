module basic_1000_10000_1500_2_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5005,N_5007,N_5011,N_5012,N_5014,N_5017,N_5018,N_5020,N_5021,N_5022,N_5023,N_5025,N_5031,N_5033,N_5036,N_5039,N_5041,N_5042,N_5043,N_5044,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5054,N_5056,N_5058,N_5059,N_5061,N_5066,N_5067,N_5069,N_5073,N_5074,N_5076,N_5077,N_5078,N_5080,N_5082,N_5083,N_5084,N_5086,N_5089,N_5090,N_5093,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5107,N_5108,N_5110,N_5112,N_5113,N_5114,N_5116,N_5117,N_5119,N_5120,N_5124,N_5125,N_5126,N_5127,N_5129,N_5133,N_5135,N_5136,N_5137,N_5139,N_5140,N_5142,N_5144,N_5146,N_5147,N_5148,N_5149,N_5150,N_5152,N_5153,N_5155,N_5157,N_5159,N_5161,N_5163,N_5166,N_5168,N_5170,N_5173,N_5175,N_5176,N_5179,N_5180,N_5181,N_5183,N_5184,N_5185,N_5188,N_5190,N_5193,N_5194,N_5196,N_5197,N_5198,N_5199,N_5203,N_5205,N_5206,N_5207,N_5210,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5219,N_5221,N_5222,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5234,N_5236,N_5237,N_5240,N_5242,N_5244,N_5248,N_5249,N_5250,N_5253,N_5254,N_5255,N_5256,N_5257,N_5260,N_5262,N_5263,N_5264,N_5265,N_5267,N_5268,N_5269,N_5270,N_5273,N_5275,N_5278,N_5279,N_5280,N_5281,N_5282,N_5284,N_5285,N_5287,N_5288,N_5289,N_5291,N_5292,N_5295,N_5296,N_5297,N_5298,N_5300,N_5301,N_5302,N_5304,N_5305,N_5306,N_5309,N_5310,N_5312,N_5313,N_5314,N_5315,N_5318,N_5321,N_5323,N_5324,N_5326,N_5327,N_5331,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5344,N_5345,N_5346,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5356,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5367,N_5369,N_5370,N_5371,N_5372,N_5373,N_5375,N_5376,N_5378,N_5381,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5393,N_5394,N_5396,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5406,N_5407,N_5409,N_5412,N_5413,N_5415,N_5416,N_5420,N_5422,N_5423,N_5424,N_5428,N_5430,N_5431,N_5432,N_5433,N_5434,N_5436,N_5439,N_5441,N_5442,N_5444,N_5445,N_5446,N_5447,N_5450,N_5451,N_5452,N_5453,N_5454,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5463,N_5464,N_5465,N_5466,N_5468,N_5469,N_5470,N_5472,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5486,N_5490,N_5491,N_5492,N_5494,N_5495,N_5496,N_5497,N_5498,N_5501,N_5502,N_5503,N_5504,N_5505,N_5507,N_5508,N_5509,N_5510,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5529,N_5530,N_5531,N_5535,N_5538,N_5539,N_5540,N_5541,N_5544,N_5546,N_5547,N_5549,N_5550,N_5551,N_5552,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5563,N_5564,N_5565,N_5567,N_5569,N_5571,N_5572,N_5576,N_5577,N_5578,N_5581,N_5582,N_5588,N_5589,N_5590,N_5592,N_5593,N_5597,N_5598,N_5600,N_5601,N_5603,N_5604,N_5605,N_5607,N_5608,N_5610,N_5611,N_5612,N_5613,N_5615,N_5616,N_5619,N_5620,N_5621,N_5624,N_5626,N_5627,N_5629,N_5630,N_5631,N_5633,N_5634,N_5635,N_5636,N_5638,N_5641,N_5642,N_5644,N_5647,N_5649,N_5650,N_5652,N_5653,N_5655,N_5657,N_5659,N_5660,N_5661,N_5663,N_5664,N_5665,N_5666,N_5667,N_5670,N_5671,N_5672,N_5676,N_5678,N_5679,N_5680,N_5681,N_5682,N_5684,N_5685,N_5686,N_5689,N_5691,N_5693,N_5697,N_5698,N_5700,N_5701,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5710,N_5715,N_5716,N_5717,N_5718,N_5719,N_5721,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5742,N_5744,N_5746,N_5749,N_5752,N_5754,N_5757,N_5759,N_5761,N_5762,N_5763,N_5764,N_5765,N_5767,N_5769,N_5772,N_5773,N_5774,N_5775,N_5776,N_5780,N_5782,N_5784,N_5785,N_5788,N_5789,N_5791,N_5792,N_5795,N_5796,N_5797,N_5798,N_5799,N_5802,N_5805,N_5808,N_5809,N_5810,N_5812,N_5813,N_5814,N_5815,N_5817,N_5818,N_5819,N_5821,N_5827,N_5829,N_5830,N_5832,N_5834,N_5837,N_5838,N_5839,N_5841,N_5843,N_5845,N_5846,N_5848,N_5849,N_5850,N_5853,N_5854,N_5856,N_5857,N_5859,N_5861,N_5862,N_5863,N_5864,N_5866,N_5867,N_5868,N_5870,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5882,N_5883,N_5884,N_5887,N_5888,N_5889,N_5890,N_5891,N_5893,N_5894,N_5895,N_5897,N_5898,N_5900,N_5901,N_5902,N_5903,N_5906,N_5909,N_5911,N_5912,N_5914,N_5915,N_5918,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5933,N_5934,N_5935,N_5938,N_5939,N_5940,N_5941,N_5943,N_5944,N_5945,N_5952,N_5953,N_5954,N_5955,N_5957,N_5960,N_5961,N_5963,N_5964,N_5965,N_5970,N_5972,N_5973,N_5974,N_5977,N_5978,N_5980,N_5982,N_5984,N_5986,N_5987,N_5990,N_5991,N_5995,N_5996,N_5998,N_6001,N_6003,N_6004,N_6005,N_6006,N_6008,N_6009,N_6010,N_6011,N_6013,N_6017,N_6018,N_6021,N_6022,N_6025,N_6026,N_6027,N_6029,N_6034,N_6036,N_6038,N_6041,N_6044,N_6047,N_6049,N_6050,N_6051,N_6053,N_6054,N_6055,N_6056,N_6059,N_6060,N_6062,N_6063,N_6065,N_6067,N_6068,N_6070,N_6071,N_6072,N_6073,N_6076,N_6080,N_6083,N_6088,N_6089,N_6091,N_6092,N_6094,N_6097,N_6098,N_6102,N_6104,N_6105,N_6106,N_6107,N_6108,N_6110,N_6111,N_6113,N_6114,N_6115,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6130,N_6131,N_6133,N_6135,N_6136,N_6137,N_6138,N_6144,N_6146,N_6147,N_6149,N_6150,N_6151,N_6153,N_6157,N_6158,N_6161,N_6163,N_6165,N_6168,N_6169,N_6170,N_6172,N_6174,N_6176,N_6177,N_6179,N_6180,N_6181,N_6184,N_6186,N_6190,N_6191,N_6193,N_6197,N_6199,N_6200,N_6201,N_6202,N_6204,N_6205,N_6206,N_6207,N_6211,N_6217,N_6219,N_6220,N_6222,N_6224,N_6225,N_6226,N_6227,N_6229,N_6231,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6243,N_6245,N_6246,N_6252,N_6253,N_6254,N_6255,N_6256,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6267,N_6271,N_6272,N_6273,N_6274,N_6276,N_6278,N_6279,N_6280,N_6281,N_6284,N_6285,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6295,N_6296,N_6297,N_6299,N_6300,N_6301,N_6302,N_6303,N_6306,N_6307,N_6308,N_6311,N_6314,N_6315,N_6316,N_6318,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6329,N_6330,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6344,N_6345,N_6348,N_6350,N_6353,N_6355,N_6356,N_6357,N_6358,N_6362,N_6363,N_6364,N_6366,N_6367,N_6368,N_6370,N_6371,N_6372,N_6374,N_6376,N_6378,N_6379,N_6382,N_6383,N_6385,N_6389,N_6390,N_6391,N_6393,N_6396,N_6398,N_6399,N_6400,N_6402,N_6403,N_6404,N_6406,N_6407,N_6408,N_6410,N_6413,N_6415,N_6419,N_6421,N_6426,N_6427,N_6428,N_6430,N_6431,N_6432,N_6434,N_6435,N_6437,N_6439,N_6440,N_6441,N_6442,N_6444,N_6445,N_6446,N_6448,N_6449,N_6450,N_6452,N_6453,N_6454,N_6456,N_6460,N_6461,N_6462,N_6468,N_6469,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6484,N_6485,N_6486,N_6487,N_6488,N_6490,N_6492,N_6493,N_6494,N_6496,N_6497,N_6499,N_6500,N_6502,N_6503,N_6504,N_6505,N_6508,N_6509,N_6511,N_6512,N_6513,N_6515,N_6516,N_6520,N_6521,N_6522,N_6525,N_6527,N_6528,N_6529,N_6531,N_6532,N_6533,N_6534,N_6536,N_6537,N_6538,N_6540,N_6541,N_6543,N_6544,N_6545,N_6548,N_6549,N_6552,N_6554,N_6555,N_6556,N_6557,N_6559,N_6562,N_6563,N_6564,N_6565,N_6566,N_6568,N_6570,N_6571,N_6572,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6581,N_6582,N_6583,N_6586,N_6588,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6599,N_6601,N_6602,N_6603,N_6605,N_6609,N_6612,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6623,N_6625,N_6626,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6637,N_6638,N_6642,N_6643,N_6645,N_6648,N_6649,N_6652,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6662,N_6663,N_6665,N_6666,N_6669,N_6670,N_6672,N_6674,N_6676,N_6677,N_6678,N_6679,N_6686,N_6687,N_6688,N_6691,N_6692,N_6694,N_6695,N_6696,N_6697,N_6698,N_6703,N_6704,N_6705,N_6706,N_6709,N_6710,N_6711,N_6712,N_6714,N_6716,N_6717,N_6719,N_6720,N_6721,N_6725,N_6726,N_6727,N_6728,N_6729,N_6734,N_6738,N_6740,N_6742,N_6745,N_6747,N_6748,N_6751,N_6753,N_6756,N_6758,N_6761,N_6766,N_6769,N_6771,N_6772,N_6773,N_6774,N_6775,N_6777,N_6780,N_6781,N_6782,N_6783,N_6785,N_6788,N_6789,N_6792,N_6796,N_6798,N_6800,N_6801,N_6802,N_6804,N_6807,N_6808,N_6809,N_6812,N_6813,N_6814,N_6817,N_6818,N_6819,N_6820,N_6822,N_6823,N_6826,N_6831,N_6832,N_6833,N_6835,N_6836,N_6837,N_6839,N_6840,N_6843,N_6844,N_6845,N_6848,N_6850,N_6851,N_6852,N_6853,N_6855,N_6856,N_6858,N_6861,N_6864,N_6865,N_6866,N_6867,N_6870,N_6871,N_6873,N_6874,N_6875,N_6877,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6890,N_6891,N_6892,N_6895,N_6897,N_6898,N_6899,N_6900,N_6902,N_6903,N_6904,N_6905,N_6906,N_6910,N_6913,N_6915,N_6917,N_6920,N_6921,N_6922,N_6923,N_6924,N_6928,N_6929,N_6930,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6941,N_6942,N_6943,N_6946,N_6950,N_6953,N_6954,N_6955,N_6961,N_6962,N_6965,N_6966,N_6967,N_6969,N_6971,N_6973,N_6976,N_6977,N_6980,N_6982,N_6983,N_6989,N_6994,N_6995,N_6996,N_6997,N_7001,N_7003,N_7004,N_7008,N_7009,N_7010,N_7012,N_7014,N_7015,N_7016,N_7017,N_7018,N_7020,N_7021,N_7022,N_7023,N_7024,N_7027,N_7028,N_7031,N_7032,N_7033,N_7034,N_7036,N_7038,N_7039,N_7040,N_7041,N_7043,N_7044,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7058,N_7059,N_7060,N_7062,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7073,N_7075,N_7076,N_7077,N_7079,N_7081,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7090,N_7091,N_7093,N_7094,N_7096,N_7097,N_7099,N_7100,N_7102,N_7105,N_7108,N_7109,N_7110,N_7111,N_7113,N_7116,N_7117,N_7120,N_7121,N_7123,N_7125,N_7130,N_7131,N_7132,N_7134,N_7136,N_7137,N_7140,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7157,N_7158,N_7159,N_7162,N_7166,N_7167,N_7168,N_7172,N_7173,N_7175,N_7176,N_7177,N_7180,N_7181,N_7182,N_7184,N_7185,N_7186,N_7190,N_7193,N_7195,N_7196,N_7197,N_7198,N_7199,N_7201,N_7202,N_7203,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7216,N_7217,N_7218,N_7219,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7237,N_7239,N_7242,N_7246,N_7247,N_7249,N_7256,N_7258,N_7259,N_7260,N_7261,N_7263,N_7264,N_7266,N_7268,N_7270,N_7271,N_7274,N_7275,N_7277,N_7279,N_7280,N_7281,N_7283,N_7284,N_7286,N_7287,N_7289,N_7290,N_7291,N_7292,N_7293,N_7295,N_7296,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7307,N_7311,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7323,N_7324,N_7325,N_7326,N_7329,N_7334,N_7336,N_7338,N_7341,N_7343,N_7344,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7355,N_7358,N_7359,N_7361,N_7363,N_7365,N_7367,N_7370,N_7371,N_7372,N_7373,N_7374,N_7377,N_7379,N_7380,N_7382,N_7383,N_7384,N_7385,N_7386,N_7390,N_7391,N_7392,N_7396,N_7397,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7408,N_7410,N_7412,N_7413,N_7416,N_7418,N_7421,N_7422,N_7426,N_7427,N_7430,N_7431,N_7432,N_7436,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7448,N_7449,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7463,N_7465,N_7468,N_7471,N_7472,N_7473,N_7474,N_7476,N_7477,N_7478,N_7482,N_7483,N_7484,N_7485,N_7486,N_7488,N_7489,N_7491,N_7492,N_7493,N_7495,N_7496,N_7499,N_7501,N_7502,N_7504,N_7505,N_7506,N_7507,N_7509,N_7512,N_7513,N_7515,N_7517,N_7518,N_7520,N_7521,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7535,N_7536,N_7537,N_7538,N_7540,N_7541,N_7542,N_7543,N_7545,N_7546,N_7548,N_7549,N_7552,N_7553,N_7554,N_7555,N_7557,N_7558,N_7560,N_7561,N_7563,N_7564,N_7566,N_7567,N_7570,N_7572,N_7573,N_7576,N_7581,N_7583,N_7584,N_7586,N_7588,N_7590,N_7591,N_7593,N_7595,N_7597,N_7600,N_7601,N_7603,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7616,N_7617,N_7619,N_7620,N_7622,N_7623,N_7624,N_7625,N_7628,N_7632,N_7634,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7645,N_7646,N_7648,N_7650,N_7651,N_7654,N_7655,N_7656,N_7659,N_7663,N_7664,N_7666,N_7668,N_7669,N_7670,N_7674,N_7675,N_7676,N_7679,N_7680,N_7681,N_7682,N_7686,N_7687,N_7688,N_7690,N_7694,N_7695,N_7696,N_7697,N_7698,N_7700,N_7701,N_7703,N_7704,N_7705,N_7706,N_7707,N_7713,N_7715,N_7717,N_7718,N_7719,N_7720,N_7724,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7735,N_7739,N_7741,N_7742,N_7743,N_7744,N_7746,N_7750,N_7751,N_7752,N_7756,N_7757,N_7758,N_7760,N_7761,N_7763,N_7764,N_7766,N_7767,N_7769,N_7770,N_7772,N_7773,N_7779,N_7781,N_7782,N_7784,N_7785,N_7787,N_7788,N_7789,N_7791,N_7796,N_7797,N_7799,N_7800,N_7801,N_7802,N_7803,N_7805,N_7806,N_7807,N_7809,N_7811,N_7814,N_7817,N_7820,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7830,N_7832,N_7833,N_7838,N_7839,N_7844,N_7845,N_7846,N_7847,N_7849,N_7853,N_7854,N_7855,N_7858,N_7859,N_7865,N_7867,N_7868,N_7869,N_7870,N_7873,N_7875,N_7878,N_7879,N_7881,N_7883,N_7888,N_7889,N_7890,N_7892,N_7895,N_7896,N_7898,N_7899,N_7903,N_7904,N_7906,N_7907,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7918,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7931,N_7932,N_7935,N_7936,N_7942,N_7943,N_7947,N_7948,N_7950,N_7952,N_7955,N_7958,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7982,N_7983,N_7984,N_7985,N_7987,N_7991,N_7992,N_7993,N_7996,N_7997,N_7998,N_8000,N_8002,N_8003,N_8006,N_8009,N_8011,N_8012,N_8016,N_8017,N_8018,N_8019,N_8021,N_8026,N_8027,N_8029,N_8030,N_8033,N_8034,N_8038,N_8039,N_8042,N_8043,N_8044,N_8046,N_8049,N_8051,N_8054,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8063,N_8065,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8078,N_8079,N_8080,N_8084,N_8086,N_8090,N_8094,N_8096,N_8097,N_8101,N_8102,N_8105,N_8106,N_8107,N_8110,N_8111,N_8114,N_8117,N_8120,N_8121,N_8122,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8132,N_8133,N_8134,N_8136,N_8137,N_8138,N_8139,N_8142,N_8144,N_8145,N_8147,N_8148,N_8149,N_8154,N_8155,N_8156,N_8157,N_8162,N_8163,N_8164,N_8167,N_8168,N_8170,N_8172,N_8174,N_8176,N_8178,N_8179,N_8180,N_8181,N_8185,N_8188,N_8190,N_8193,N_8194,N_8195,N_8196,N_8197,N_8203,N_8205,N_8206,N_8209,N_8213,N_8214,N_8217,N_8218,N_8222,N_8224,N_8225,N_8228,N_8231,N_8235,N_8236,N_8237,N_8238,N_8239,N_8241,N_8242,N_8244,N_8245,N_8246,N_8247,N_8249,N_8250,N_8252,N_8256,N_8258,N_8260,N_8263,N_8264,N_8265,N_8266,N_8268,N_8270,N_8271,N_8273,N_8274,N_8275,N_8276,N_8278,N_8279,N_8280,N_8282,N_8284,N_8285,N_8286,N_8288,N_8290,N_8293,N_8296,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8312,N_8315,N_8316,N_8318,N_8320,N_8321,N_8324,N_8325,N_8326,N_8328,N_8330,N_8332,N_8333,N_8334,N_8337,N_8340,N_8341,N_8342,N_8344,N_8346,N_8349,N_8352,N_8357,N_8359,N_8362,N_8363,N_8364,N_8365,N_8367,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8379,N_8380,N_8381,N_8382,N_8384,N_8385,N_8388,N_8390,N_8391,N_8392,N_8396,N_8397,N_8401,N_8402,N_8403,N_8405,N_8407,N_8408,N_8409,N_8410,N_8412,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8423,N_8429,N_8430,N_8433,N_8434,N_8435,N_8436,N_8437,N_8439,N_8441,N_8442,N_8443,N_8444,N_8446,N_8447,N_8450,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8460,N_8461,N_8463,N_8464,N_8466,N_8467,N_8470,N_8472,N_8473,N_8474,N_8475,N_8477,N_8478,N_8480,N_8481,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8496,N_8498,N_8500,N_8501,N_8502,N_8505,N_8506,N_8507,N_8509,N_8511,N_8513,N_8515,N_8517,N_8518,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8535,N_8539,N_8540,N_8541,N_8542,N_8544,N_8546,N_8548,N_8549,N_8552,N_8553,N_8554,N_8556,N_8559,N_8560,N_8561,N_8563,N_8565,N_8566,N_8567,N_8568,N_8569,N_8571,N_8572,N_8574,N_8576,N_8577,N_8578,N_8580,N_8582,N_8583,N_8584,N_8586,N_8587,N_8589,N_8590,N_8591,N_8592,N_8594,N_8596,N_8600,N_8601,N_8603,N_8604,N_8606,N_8607,N_8608,N_8609,N_8610,N_8612,N_8613,N_8614,N_8615,N_8616,N_8620,N_8621,N_8622,N_8624,N_8625,N_8626,N_8628,N_8629,N_8631,N_8634,N_8635,N_8636,N_8638,N_8640,N_8642,N_8643,N_8644,N_8645,N_8649,N_8650,N_8652,N_8653,N_8654,N_8655,N_8657,N_8658,N_8659,N_8660,N_8664,N_8665,N_8666,N_8669,N_8670,N_8672,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8686,N_8688,N_8692,N_8696,N_8697,N_8699,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8710,N_8711,N_8714,N_8715,N_8716,N_8718,N_8719,N_8720,N_8721,N_8723,N_8724,N_8727,N_8728,N_8731,N_8732,N_8736,N_8740,N_8741,N_8743,N_8745,N_8746,N_8748,N_8749,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8759,N_8761,N_8762,N_8764,N_8766,N_8768,N_8770,N_8772,N_8773,N_8775,N_8776,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8788,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8799,N_8803,N_8806,N_8811,N_8813,N_8814,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8824,N_8826,N_8827,N_8828,N_8832,N_8834,N_8835,N_8837,N_8838,N_8839,N_8844,N_8846,N_8847,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8856,N_8858,N_8859,N_8860,N_8864,N_8865,N_8867,N_8868,N_8870,N_8871,N_8872,N_8873,N_8874,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8896,N_8898,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8923,N_8924,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8933,N_8935,N_8936,N_8938,N_8943,N_8946,N_8947,N_8950,N_8953,N_8954,N_8957,N_8958,N_8961,N_8962,N_8965,N_8967,N_8968,N_8970,N_8971,N_8972,N_8974,N_8978,N_8980,N_8986,N_8989,N_8991,N_8993,N_8994,N_8995,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9005,N_9007,N_9008,N_9009,N_9010,N_9014,N_9015,N_9016,N_9019,N_9021,N_9022,N_9024,N_9025,N_9026,N_9027,N_9028,N_9030,N_9031,N_9035,N_9036,N_9037,N_9038,N_9039,N_9043,N_9044,N_9045,N_9046,N_9051,N_9053,N_9054,N_9056,N_9057,N_9059,N_9062,N_9065,N_9067,N_9068,N_9070,N_9071,N_9073,N_9074,N_9075,N_9076,N_9077,N_9081,N_9082,N_9083,N_9087,N_9088,N_9090,N_9092,N_9093,N_9094,N_9096,N_9100,N_9103,N_9104,N_9105,N_9107,N_9108,N_9110,N_9111,N_9114,N_9115,N_9116,N_9119,N_9120,N_9123,N_9124,N_9125,N_9126,N_9127,N_9130,N_9131,N_9133,N_9134,N_9135,N_9136,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9146,N_9150,N_9154,N_9155,N_9156,N_9157,N_9159,N_9161,N_9162,N_9163,N_9165,N_9166,N_9169,N_9172,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9182,N_9183,N_9185,N_9188,N_9190,N_9191,N_9192,N_9193,N_9195,N_9196,N_9197,N_9198,N_9203,N_9205,N_9207,N_9209,N_9211,N_9215,N_9216,N_9217,N_9219,N_9220,N_9221,N_9222,N_9224,N_9226,N_9228,N_9229,N_9230,N_9231,N_9233,N_9235,N_9238,N_9239,N_9243,N_9244,N_9245,N_9247,N_9248,N_9249,N_9250,N_9252,N_9254,N_9255,N_9256,N_9258,N_9262,N_9263,N_9266,N_9269,N_9270,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9281,N_9283,N_9291,N_9292,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9320,N_9321,N_9324,N_9326,N_9327,N_9330,N_9331,N_9332,N_9334,N_9336,N_9338,N_9341,N_9345,N_9346,N_9349,N_9350,N_9353,N_9355,N_9356,N_9357,N_9358,N_9359,N_9361,N_9362,N_9363,N_9364,N_9365,N_9369,N_9371,N_9373,N_9375,N_9377,N_9378,N_9380,N_9384,N_9387,N_9388,N_9390,N_9393,N_9394,N_9395,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9404,N_9405,N_9406,N_9407,N_9408,N_9410,N_9412,N_9413,N_9415,N_9417,N_9418,N_9420,N_9422,N_9424,N_9426,N_9427,N_9429,N_9430,N_9431,N_9433,N_9436,N_9438,N_9439,N_9440,N_9441,N_9442,N_9445,N_9446,N_9447,N_9448,N_9449,N_9452,N_9455,N_9456,N_9461,N_9462,N_9464,N_9466,N_9469,N_9471,N_9472,N_9473,N_9474,N_9475,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9484,N_9485,N_9486,N_9490,N_9491,N_9492,N_9493,N_9494,N_9498,N_9501,N_9502,N_9504,N_9506,N_9507,N_9510,N_9512,N_9513,N_9516,N_9517,N_9518,N_9523,N_9524,N_9525,N_9527,N_9528,N_9529,N_9531,N_9533,N_9535,N_9537,N_9538,N_9540,N_9542,N_9543,N_9547,N_9549,N_9550,N_9551,N_9553,N_9554,N_9556,N_9558,N_9560,N_9561,N_9562,N_9564,N_9565,N_9566,N_9568,N_9571,N_9572,N_9573,N_9574,N_9575,N_9577,N_9578,N_9580,N_9581,N_9582,N_9583,N_9584,N_9587,N_9589,N_9590,N_9592,N_9593,N_9596,N_9598,N_9600,N_9603,N_9604,N_9605,N_9610,N_9611,N_9613,N_9616,N_9617,N_9618,N_9619,N_9623,N_9624,N_9627,N_9629,N_9630,N_9634,N_9635,N_9637,N_9639,N_9641,N_9642,N_9643,N_9644,N_9645,N_9647,N_9649,N_9650,N_9651,N_9654,N_9656,N_9658,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9669,N_9671,N_9672,N_9673,N_9675,N_9676,N_9680,N_9681,N_9684,N_9688,N_9689,N_9690,N_9694,N_9695,N_9697,N_9700,N_9702,N_9704,N_9705,N_9707,N_9708,N_9709,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9718,N_9720,N_9725,N_9726,N_9727,N_9729,N_9733,N_9735,N_9736,N_9739,N_9741,N_9742,N_9743,N_9744,N_9746,N_9748,N_9749,N_9750,N_9751,N_9753,N_9754,N_9755,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9765,N_9766,N_9768,N_9770,N_9771,N_9772,N_9773,N_9774,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9786,N_9788,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9798,N_9799,N_9800,N_9801,N_9802,N_9805,N_9808,N_9809,N_9812,N_9813,N_9814,N_9818,N_9820,N_9822,N_9824,N_9827,N_9828,N_9830,N_9831,N_9833,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9845,N_9848,N_9851,N_9852,N_9853,N_9854,N_9857,N_9858,N_9859,N_9861,N_9862,N_9863,N_9866,N_9868,N_9872,N_9873,N_9875,N_9876,N_9879,N_9880,N_9881,N_9882,N_9883,N_9888,N_9889,N_9890,N_9892,N_9895,N_9896,N_9897,N_9898,N_9900,N_9901,N_9903,N_9905,N_9906,N_9908,N_9909,N_9912,N_9913,N_9914,N_9916,N_9918,N_9919,N_9920,N_9921,N_9922,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9932,N_9934,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9946,N_9950,N_9951,N_9952,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9963,N_9964,N_9969,N_9970,N_9971,N_9972,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9990,N_9991,N_9992,N_9993,N_9996,N_9997,N_9998;
and U0 (N_0,In_303,In_281);
or U1 (N_1,In_223,In_676);
nand U2 (N_2,In_960,In_235);
nor U3 (N_3,In_4,In_945);
nor U4 (N_4,In_706,In_702);
nor U5 (N_5,In_584,In_462);
xnor U6 (N_6,In_961,In_568);
and U7 (N_7,In_209,In_670);
or U8 (N_8,In_822,In_832);
and U9 (N_9,In_616,In_878);
nor U10 (N_10,In_596,In_912);
nor U11 (N_11,In_517,In_168);
and U12 (N_12,In_577,In_870);
or U13 (N_13,In_597,In_483);
and U14 (N_14,In_218,In_682);
nand U15 (N_15,In_821,In_899);
and U16 (N_16,In_889,In_307);
nor U17 (N_17,In_109,In_309);
and U18 (N_18,In_610,In_155);
nor U19 (N_19,In_190,In_54);
nor U20 (N_20,In_313,In_57);
or U21 (N_21,In_453,In_849);
and U22 (N_22,In_824,In_216);
nand U23 (N_23,In_126,In_371);
or U24 (N_24,In_70,In_872);
and U25 (N_25,In_166,In_603);
nand U26 (N_26,In_681,In_726);
nor U27 (N_27,In_51,In_384);
or U28 (N_28,In_6,In_399);
nor U29 (N_29,In_906,In_71);
nand U30 (N_30,In_599,In_703);
and U31 (N_31,In_693,In_316);
nor U32 (N_32,In_276,In_177);
and U33 (N_33,In_966,In_994);
nor U34 (N_34,In_664,In_201);
nand U35 (N_35,In_589,In_374);
or U36 (N_36,In_748,In_141);
nor U37 (N_37,In_659,In_712);
or U38 (N_38,In_540,In_488);
nor U39 (N_39,In_474,In_741);
and U40 (N_40,In_755,In_233);
nor U41 (N_41,In_524,In_154);
and U42 (N_42,In_532,In_674);
nor U43 (N_43,In_396,In_640);
or U44 (N_44,In_151,In_965);
and U45 (N_45,In_841,In_807);
nand U46 (N_46,In_632,In_447);
nor U47 (N_47,In_636,In_379);
nand U48 (N_48,In_704,In_542);
or U49 (N_49,In_534,In_690);
nor U50 (N_50,In_354,In_308);
nor U51 (N_51,In_918,In_974);
or U52 (N_52,In_811,In_314);
nor U53 (N_53,In_300,In_465);
nor U54 (N_54,In_132,In_806);
nor U55 (N_55,In_587,In_837);
or U56 (N_56,In_716,In_147);
nand U57 (N_57,In_221,In_302);
and U58 (N_58,In_948,In_880);
nand U59 (N_59,In_156,In_123);
nand U60 (N_60,In_627,In_76);
and U61 (N_61,In_56,In_251);
nor U62 (N_62,In_479,In_290);
and U63 (N_63,In_203,In_253);
nor U64 (N_64,In_503,In_521);
or U65 (N_65,In_157,In_35);
nand U66 (N_66,In_868,In_338);
nor U67 (N_67,In_434,In_691);
nand U68 (N_68,In_138,In_771);
nor U69 (N_69,In_576,In_901);
nor U70 (N_70,In_722,In_819);
nor U71 (N_71,In_264,In_367);
or U72 (N_72,In_87,In_266);
nor U73 (N_73,In_93,In_930);
and U74 (N_74,In_916,In_717);
nand U75 (N_75,In_903,In_801);
or U76 (N_76,In_747,In_433);
or U77 (N_77,In_591,In_359);
nand U78 (N_78,In_407,In_590);
nor U79 (N_79,In_514,In_200);
nand U80 (N_80,In_937,In_803);
nand U81 (N_81,In_506,In_917);
and U82 (N_82,In_954,In_508);
nor U83 (N_83,In_24,In_998);
nand U84 (N_84,In_969,In_471);
nor U85 (N_85,In_284,In_387);
nand U86 (N_86,In_970,In_864);
and U87 (N_87,In_951,In_923);
or U88 (N_88,In_713,In_9);
nor U89 (N_89,In_431,In_364);
and U90 (N_90,In_675,In_529);
and U91 (N_91,In_452,In_790);
or U92 (N_92,In_139,In_826);
nor U93 (N_93,In_861,In_75);
nor U94 (N_94,In_993,In_692);
nor U95 (N_95,In_74,In_928);
nand U96 (N_96,In_641,In_496);
nor U97 (N_97,In_796,In_426);
and U98 (N_98,In_184,In_356);
and U99 (N_99,In_740,In_617);
and U100 (N_100,In_896,In_427);
and U101 (N_101,In_813,In_259);
xnor U102 (N_102,In_891,In_193);
and U103 (N_103,In_921,In_770);
nand U104 (N_104,In_707,In_247);
nand U105 (N_105,In_77,In_622);
nand U106 (N_106,In_229,In_871);
and U107 (N_107,In_386,In_958);
or U108 (N_108,In_325,In_679);
and U109 (N_109,In_797,In_876);
or U110 (N_110,In_225,In_935);
or U111 (N_111,In_915,In_500);
or U112 (N_112,In_606,In_708);
nor U113 (N_113,In_167,In_331);
and U114 (N_114,In_360,In_963);
nor U115 (N_115,In_291,In_683);
and U116 (N_116,In_561,In_262);
or U117 (N_117,In_105,In_68);
nor U118 (N_118,In_59,In_793);
nand U119 (N_119,In_982,In_213);
or U120 (N_120,In_898,In_14);
or U121 (N_121,In_799,In_977);
nand U122 (N_122,In_794,In_420);
and U123 (N_123,In_351,In_619);
nor U124 (N_124,In_724,In_792);
nor U125 (N_125,In_454,In_329);
nand U126 (N_126,In_689,In_851);
or U127 (N_127,In_185,In_107);
and U128 (N_128,In_875,In_996);
nand U129 (N_129,In_240,In_888);
or U130 (N_130,In_538,In_642);
nand U131 (N_131,In_121,In_212);
nand U132 (N_132,In_95,In_220);
and U133 (N_133,In_782,In_457);
and U134 (N_134,In_239,In_611);
nand U135 (N_135,In_321,In_287);
and U136 (N_136,In_415,In_478);
and U137 (N_137,In_758,In_395);
and U138 (N_138,In_501,In_980);
nor U139 (N_139,In_241,In_336);
nand U140 (N_140,In_265,In_781);
nor U141 (N_141,In_710,In_491);
nor U142 (N_142,In_818,In_949);
or U143 (N_143,In_205,In_545);
nor U144 (N_144,In_455,In_440);
nor U145 (N_145,In_477,In_380);
or U146 (N_146,In_289,In_729);
nand U147 (N_147,In_983,In_40);
nand U148 (N_148,In_709,In_327);
or U149 (N_149,In_518,In_353);
nand U150 (N_150,In_110,In_637);
and U151 (N_151,In_856,In_907);
nand U152 (N_152,In_946,In_409);
xnor U153 (N_153,In_618,In_775);
nor U154 (N_154,In_340,In_823);
nand U155 (N_155,In_42,In_342);
nor U156 (N_156,In_297,In_492);
or U157 (N_157,In_173,In_389);
and U158 (N_158,In_544,In_887);
nand U159 (N_159,In_48,In_654);
and U160 (N_160,In_523,In_728);
or U161 (N_161,In_897,In_294);
and U162 (N_162,In_553,In_365);
nand U163 (N_163,In_988,In_762);
nor U164 (N_164,In_468,In_493);
nand U165 (N_165,In_429,In_292);
nor U166 (N_166,In_145,In_487);
or U167 (N_167,In_410,In_224);
nor U168 (N_168,In_680,In_131);
or U169 (N_169,In_677,In_234);
nand U170 (N_170,In_248,In_45);
and U171 (N_171,In_720,In_23);
nand U172 (N_172,In_779,In_49);
or U173 (N_173,In_29,In_179);
or U174 (N_174,In_866,In_343);
nand U175 (N_175,In_750,In_602);
nor U176 (N_176,In_564,In_261);
or U177 (N_177,In_394,In_723);
nand U178 (N_178,In_128,In_705);
or U179 (N_179,In_260,In_684);
and U180 (N_180,In_939,In_593);
nand U181 (N_181,In_435,In_743);
or U182 (N_182,In_361,In_971);
and U183 (N_183,In_438,In_215);
nand U184 (N_184,In_774,In_385);
or U185 (N_185,In_104,In_345);
nand U186 (N_186,In_867,In_183);
nor U187 (N_187,In_688,In_122);
and U188 (N_188,In_381,In_99);
and U189 (N_189,In_249,In_258);
and U190 (N_190,In_41,In_10);
or U191 (N_191,In_368,In_277);
nor U192 (N_192,In_924,In_349);
nor U193 (N_193,In_600,In_2);
and U194 (N_194,In_194,In_947);
nor U195 (N_195,In_102,In_686);
and U196 (N_196,In_973,In_464);
nand U197 (N_197,In_990,In_809);
and U198 (N_198,In_186,In_79);
and U199 (N_199,In_129,In_651);
nand U200 (N_200,In_450,In_85);
or U201 (N_201,In_579,In_714);
or U202 (N_202,In_555,In_744);
and U203 (N_203,In_817,In_445);
nand U204 (N_204,In_446,In_869);
nand U205 (N_205,In_910,In_574);
nor U206 (N_206,In_279,In_392);
nor U207 (N_207,In_181,In_113);
nor U208 (N_208,In_358,In_513);
xor U209 (N_209,In_18,In_800);
or U210 (N_210,In_376,In_256);
xor U211 (N_211,In_117,In_853);
or U212 (N_212,In_556,In_98);
xnor U213 (N_213,In_335,In_393);
nor U214 (N_214,In_400,In_526);
nand U215 (N_215,In_67,In_789);
nand U216 (N_216,In_467,In_152);
nor U217 (N_217,In_892,In_612);
and U218 (N_218,In_839,In_926);
nor U219 (N_219,In_378,In_893);
nor U220 (N_220,In_94,In_834);
nand U221 (N_221,In_495,In_598);
or U222 (N_222,In_560,In_463);
and U223 (N_223,In_655,In_169);
and U224 (N_224,In_243,In_176);
or U225 (N_225,In_83,In_607);
and U226 (N_226,In_721,In_873);
or U227 (N_227,In_62,In_835);
nor U228 (N_228,In_148,In_119);
nand U229 (N_229,In_27,In_999);
nor U230 (N_230,In_164,In_428);
nor U231 (N_231,In_69,In_348);
or U232 (N_232,In_634,In_595);
and U233 (N_233,In_699,In_268);
nand U234 (N_234,In_512,In_546);
or U235 (N_235,In_430,In_88);
nand U236 (N_236,In_337,In_795);
nor U237 (N_237,In_698,In_572);
nand U238 (N_238,In_347,In_628);
and U239 (N_239,In_456,In_350);
nor U240 (N_240,In_558,In_298);
nand U241 (N_241,In_533,In_485);
nand U242 (N_242,In_578,In_423);
and U243 (N_243,In_32,In_270);
nand U244 (N_244,In_421,In_820);
nor U245 (N_245,In_149,In_894);
nand U246 (N_246,In_170,In_238);
nand U247 (N_247,In_159,In_814);
and U248 (N_248,In_886,In_210);
or U249 (N_249,In_569,In_660);
nor U250 (N_250,In_621,In_112);
nor U251 (N_251,In_111,In_144);
or U252 (N_252,In_377,In_746);
nor U253 (N_253,In_459,In_7);
or U254 (N_254,In_53,In_672);
or U255 (N_255,In_363,In_541);
or U256 (N_256,In_908,In_669);
nand U257 (N_257,In_283,In_175);
nand U258 (N_258,In_985,In_346);
nand U259 (N_259,In_586,In_153);
and U260 (N_260,In_769,In_763);
or U261 (N_261,In_784,In_967);
nor U262 (N_262,In_65,In_383);
and U263 (N_263,In_609,In_647);
nand U264 (N_264,In_900,In_644);
or U265 (N_265,In_658,In_28);
and U266 (N_266,In_668,In_847);
nor U267 (N_267,In_520,In_120);
nand U268 (N_268,In_525,In_972);
or U269 (N_269,In_31,In_649);
nor U270 (N_270,In_940,In_15);
or U271 (N_271,In_305,In_757);
and U272 (N_272,In_648,In_494);
or U273 (N_273,In_401,In_317);
nor U274 (N_274,In_12,In_217);
and U275 (N_275,In_161,In_613);
nor U276 (N_276,In_527,In_208);
nor U277 (N_277,In_766,In_581);
nand U278 (N_278,In_976,In_780);
or U279 (N_279,In_646,In_552);
or U280 (N_280,In_461,In_719);
nor U281 (N_281,In_328,In_573);
or U282 (N_282,In_252,In_530);
nor U283 (N_283,In_135,In_171);
and U284 (N_284,In_981,In_319);
nor U285 (N_285,In_678,In_448);
and U286 (N_286,In_245,In_288);
nor U287 (N_287,In_0,In_997);
and U288 (N_288,In_275,In_226);
or U289 (N_289,In_460,In_242);
nor U290 (N_290,In_372,In_650);
or U291 (N_291,In_759,In_964);
nor U292 (N_292,In_17,In_620);
or U293 (N_293,In_333,In_267);
nor U294 (N_294,In_785,In_933);
or U295 (N_295,In_195,In_543);
nand U296 (N_296,In_286,In_810);
or U297 (N_297,In_850,In_608);
or U298 (N_298,In_808,In_968);
or U299 (N_299,In_55,In_114);
nand U300 (N_300,In_735,In_341);
xor U301 (N_301,In_80,In_751);
and U302 (N_302,In_528,In_911);
or U303 (N_303,In_855,In_696);
nor U304 (N_304,In_843,In_318);
and U305 (N_305,In_21,In_192);
nor U306 (N_306,In_274,In_777);
and U307 (N_307,In_33,In_323);
or U308 (N_308,In_922,In_936);
nand U309 (N_309,In_332,In_580);
nor U310 (N_310,In_745,In_369);
or U311 (N_311,In_842,In_643);
nor U312 (N_312,In_1,In_730);
and U313 (N_313,In_885,In_804);
nand U314 (N_314,In_941,In_100);
nor U315 (N_315,In_504,In_442);
or U316 (N_316,In_146,In_106);
or U317 (N_317,In_742,In_989);
and U318 (N_318,In_854,In_845);
and U319 (N_319,In_406,In_418);
or U320 (N_320,In_232,In_549);
and U321 (N_321,In_163,In_441);
or U322 (N_322,In_116,In_370);
nor U323 (N_323,In_66,In_484);
or U324 (N_324,In_404,In_667);
nor U325 (N_325,In_344,In_34);
or U326 (N_326,In_196,In_522);
and U327 (N_327,In_189,In_296);
nor U328 (N_328,In_604,In_391);
nand U329 (N_329,In_204,In_548);
and U330 (N_330,In_925,In_519);
nand U331 (N_331,In_82,In_825);
or U332 (N_332,In_957,In_697);
or U333 (N_333,In_43,In_26);
or U334 (N_334,In_22,In_246);
or U335 (N_335,In_78,In_874);
nand U336 (N_336,In_827,In_978);
and U337 (N_337,In_516,In_89);
and U338 (N_338,In_739,In_752);
nand U339 (N_339,In_315,In_783);
or U340 (N_340,In_46,In_206);
and U341 (N_341,In_412,In_614);
nor U342 (N_342,In_881,In_211);
and U343 (N_343,In_437,In_398);
nor U344 (N_344,In_838,In_366);
and U345 (N_345,In_840,In_987);
and U346 (N_346,In_97,In_414);
nor U347 (N_347,In_615,In_8);
nor U348 (N_348,In_230,In_539);
or U349 (N_349,In_934,In_72);
nand U350 (N_350,In_760,In_944);
nor U351 (N_351,In_39,In_382);
and U352 (N_352,In_657,In_511);
or U353 (N_353,In_671,In_373);
nor U354 (N_354,In_60,In_443);
or U355 (N_355,In_753,In_927);
nor U356 (N_356,In_405,In_64);
nor U357 (N_357,In_115,In_58);
and U358 (N_358,In_301,In_489);
nand U359 (N_359,In_626,In_73);
nand U360 (N_360,In_497,In_436);
nor U361 (N_361,In_375,In_816);
nor U362 (N_362,In_846,In_929);
nand U363 (N_363,In_734,In_694);
nand U364 (N_364,In_482,In_571);
or U365 (N_365,In_562,In_633);
or U366 (N_366,In_623,In_727);
nor U367 (N_367,In_188,In_663);
or U368 (N_368,In_432,In_879);
and U369 (N_369,In_662,In_269);
nand U370 (N_370,In_701,In_505);
nor U371 (N_371,In_828,In_877);
nand U372 (N_372,In_127,In_992);
or U373 (N_373,In_390,In_172);
or U374 (N_374,In_905,In_857);
nor U375 (N_375,In_984,In_476);
nand U376 (N_376,In_355,In_673);
nand U377 (N_377,In_84,In_575);
nor U378 (N_378,In_451,In_731);
xnor U379 (N_379,In_550,In_202);
nand U380 (N_380,In_180,In_805);
xnor U381 (N_381,In_938,In_480);
nand U382 (N_382,In_272,In_352);
or U383 (N_383,In_509,In_557);
nand U384 (N_384,In_466,In_199);
and U385 (N_385,In_890,In_165);
or U386 (N_386,In_137,In_909);
or U387 (N_387,In_310,In_919);
nand U388 (N_388,In_601,In_36);
nand U389 (N_389,In_472,In_531);
nand U390 (N_390,In_299,In_143);
nand U391 (N_391,In_187,In_588);
and U392 (N_392,In_551,In_754);
and U393 (N_393,In_942,In_334);
nor U394 (N_394,In_830,In_214);
and U395 (N_395,In_362,In_473);
xor U396 (N_396,In_37,In_162);
and U397 (N_397,In_848,In_859);
nor U398 (N_398,In_652,In_498);
and U399 (N_399,In_904,In_403);
or U400 (N_400,In_86,In_565);
and U401 (N_401,In_844,In_955);
nand U402 (N_402,In_3,In_207);
or U403 (N_403,In_812,In_458);
or U404 (N_404,In_311,In_481);
and U405 (N_405,In_656,In_786);
nor U406 (N_406,In_920,In_858);
nor U407 (N_407,In_408,In_638);
or U408 (N_408,In_732,In_425);
nand U409 (N_409,In_711,In_424);
nand U410 (N_410,In_756,In_469);
nand U411 (N_411,In_725,In_772);
and U412 (N_412,In_685,In_914);
and U413 (N_413,In_339,In_829);
or U414 (N_414,In_499,In_738);
and U415 (N_415,In_30,In_582);
or U416 (N_416,In_178,In_475);
nand U417 (N_417,In_416,In_749);
or U418 (N_418,In_665,In_236);
and U419 (N_419,In_142,In_507);
nand U420 (N_420,In_515,In_535);
nand U421 (N_421,In_537,In_592);
and U422 (N_422,In_44,In_605);
nor U423 (N_423,In_16,In_219);
nor U424 (N_424,In_263,In_836);
nand U425 (N_425,In_295,In_995);
or U426 (N_426,In_96,In_943);
nor U427 (N_427,In_422,In_773);
nor U428 (N_428,In_902,In_630);
and U429 (N_429,In_50,In_158);
and U430 (N_430,In_767,In_991);
nand U431 (N_431,In_140,In_788);
nor U432 (N_432,In_715,In_831);
nand U433 (N_433,In_413,In_397);
nor U434 (N_434,In_160,In_280);
nor U435 (N_435,In_883,In_322);
nor U436 (N_436,In_645,In_25);
or U437 (N_437,In_134,In_761);
nor U438 (N_438,In_510,In_567);
and U439 (N_439,In_863,In_490);
or U440 (N_440,In_198,In_312);
nor U441 (N_441,In_293,In_585);
or U442 (N_442,In_860,In_470);
and U443 (N_443,In_444,In_952);
nand U444 (N_444,In_250,In_191);
nand U445 (N_445,In_962,In_718);
nand U446 (N_446,In_737,In_103);
or U447 (N_447,In_52,In_227);
and U448 (N_448,In_63,In_38);
nor U449 (N_449,In_304,In_986);
and U450 (N_450,In_802,In_244);
nor U451 (N_451,In_733,In_629);
or U452 (N_452,In_559,In_953);
nand U453 (N_453,In_130,In_566);
or U454 (N_454,In_101,In_502);
and U455 (N_455,In_554,In_439);
nand U456 (N_456,In_326,In_273);
or U457 (N_457,In_932,In_583);
nor U458 (N_458,In_695,In_271);
nand U459 (N_459,In_862,In_20);
and U460 (N_460,In_547,In_419);
nand U461 (N_461,In_449,In_357);
nor U462 (N_462,In_118,In_257);
nor U463 (N_463,In_666,In_255);
or U464 (N_464,In_791,In_635);
and U465 (N_465,In_150,In_222);
nor U466 (N_466,In_931,In_956);
nor U467 (N_467,In_631,In_979);
nand U468 (N_468,In_285,In_182);
and U469 (N_469,In_768,In_254);
and U470 (N_470,In_765,In_19);
and U471 (N_471,In_687,In_563);
or U472 (N_472,In_92,In_950);
nand U473 (N_473,In_536,In_124);
nand U474 (N_474,In_625,In_798);
or U475 (N_475,In_778,In_700);
and U476 (N_476,In_895,In_913);
nand U477 (N_477,In_815,In_237);
and U478 (N_478,In_882,In_639);
or U479 (N_479,In_653,In_417);
nand U480 (N_480,In_776,In_402);
or U481 (N_481,In_278,In_228);
nand U482 (N_482,In_47,In_411);
nor U483 (N_483,In_282,In_136);
nand U484 (N_484,In_959,In_594);
or U485 (N_485,In_81,In_865);
and U486 (N_486,In_486,In_174);
nor U487 (N_487,In_13,In_852);
and U488 (N_488,In_388,In_90);
and U489 (N_489,In_61,In_787);
or U490 (N_490,In_306,In_324);
or U491 (N_491,In_11,In_197);
nand U492 (N_492,In_5,In_661);
nand U493 (N_493,In_624,In_330);
and U494 (N_494,In_570,In_108);
or U495 (N_495,In_91,In_320);
or U496 (N_496,In_975,In_764);
nor U497 (N_497,In_125,In_736);
xnor U498 (N_498,In_231,In_833);
or U499 (N_499,In_133,In_884);
or U500 (N_500,In_154,In_498);
or U501 (N_501,In_120,In_523);
or U502 (N_502,In_230,In_233);
nand U503 (N_503,In_464,In_553);
nand U504 (N_504,In_76,In_26);
nor U505 (N_505,In_313,In_533);
and U506 (N_506,In_427,In_566);
nor U507 (N_507,In_167,In_355);
nand U508 (N_508,In_766,In_781);
nor U509 (N_509,In_441,In_950);
and U510 (N_510,In_802,In_574);
and U511 (N_511,In_283,In_339);
nand U512 (N_512,In_640,In_698);
and U513 (N_513,In_527,In_556);
and U514 (N_514,In_340,In_988);
nor U515 (N_515,In_620,In_394);
xor U516 (N_516,In_519,In_993);
nor U517 (N_517,In_636,In_942);
nor U518 (N_518,In_102,In_388);
or U519 (N_519,In_53,In_711);
nor U520 (N_520,In_480,In_464);
nor U521 (N_521,In_551,In_186);
or U522 (N_522,In_869,In_942);
and U523 (N_523,In_143,In_222);
nor U524 (N_524,In_559,In_92);
nand U525 (N_525,In_144,In_82);
nor U526 (N_526,In_622,In_606);
and U527 (N_527,In_424,In_250);
and U528 (N_528,In_61,In_134);
or U529 (N_529,In_883,In_630);
nor U530 (N_530,In_925,In_302);
nand U531 (N_531,In_322,In_799);
and U532 (N_532,In_344,In_574);
or U533 (N_533,In_482,In_893);
or U534 (N_534,In_715,In_411);
nand U535 (N_535,In_218,In_683);
nand U536 (N_536,In_906,In_32);
nand U537 (N_537,In_125,In_290);
and U538 (N_538,In_968,In_214);
or U539 (N_539,In_931,In_177);
and U540 (N_540,In_851,In_488);
nand U541 (N_541,In_687,In_964);
nand U542 (N_542,In_200,In_15);
nand U543 (N_543,In_847,In_935);
or U544 (N_544,In_498,In_438);
nor U545 (N_545,In_34,In_616);
or U546 (N_546,In_45,In_637);
or U547 (N_547,In_263,In_34);
and U548 (N_548,In_952,In_214);
nand U549 (N_549,In_254,In_721);
and U550 (N_550,In_992,In_564);
and U551 (N_551,In_673,In_248);
or U552 (N_552,In_544,In_752);
nand U553 (N_553,In_773,In_828);
or U554 (N_554,In_174,In_87);
and U555 (N_555,In_991,In_813);
or U556 (N_556,In_19,In_920);
nand U557 (N_557,In_309,In_314);
or U558 (N_558,In_965,In_57);
and U559 (N_559,In_309,In_310);
nand U560 (N_560,In_517,In_177);
and U561 (N_561,In_138,In_575);
nor U562 (N_562,In_751,In_69);
xor U563 (N_563,In_287,In_788);
and U564 (N_564,In_523,In_351);
and U565 (N_565,In_84,In_647);
nor U566 (N_566,In_409,In_441);
and U567 (N_567,In_566,In_798);
and U568 (N_568,In_561,In_937);
nor U569 (N_569,In_501,In_5);
nand U570 (N_570,In_995,In_477);
nand U571 (N_571,In_372,In_358);
nand U572 (N_572,In_214,In_655);
or U573 (N_573,In_732,In_599);
nor U574 (N_574,In_224,In_44);
and U575 (N_575,In_172,In_841);
or U576 (N_576,In_911,In_8);
or U577 (N_577,In_522,In_432);
and U578 (N_578,In_373,In_186);
or U579 (N_579,In_536,In_759);
nand U580 (N_580,In_154,In_901);
or U581 (N_581,In_181,In_820);
and U582 (N_582,In_459,In_114);
nor U583 (N_583,In_840,In_370);
and U584 (N_584,In_82,In_340);
nor U585 (N_585,In_521,In_273);
or U586 (N_586,In_59,In_549);
nor U587 (N_587,In_12,In_601);
or U588 (N_588,In_237,In_306);
or U589 (N_589,In_812,In_173);
nor U590 (N_590,In_422,In_362);
nand U591 (N_591,In_371,In_85);
nor U592 (N_592,In_600,In_872);
nor U593 (N_593,In_222,In_888);
nand U594 (N_594,In_599,In_578);
or U595 (N_595,In_510,In_126);
nand U596 (N_596,In_947,In_126);
or U597 (N_597,In_112,In_663);
and U598 (N_598,In_745,In_413);
or U599 (N_599,In_615,In_571);
or U600 (N_600,In_693,In_483);
nand U601 (N_601,In_386,In_838);
and U602 (N_602,In_136,In_281);
nor U603 (N_603,In_843,In_844);
xor U604 (N_604,In_262,In_964);
and U605 (N_605,In_273,In_0);
or U606 (N_606,In_193,In_307);
or U607 (N_607,In_206,In_106);
xor U608 (N_608,In_977,In_667);
or U609 (N_609,In_973,In_414);
or U610 (N_610,In_567,In_552);
nor U611 (N_611,In_891,In_638);
nor U612 (N_612,In_143,In_513);
nor U613 (N_613,In_827,In_851);
nor U614 (N_614,In_967,In_690);
nor U615 (N_615,In_589,In_410);
and U616 (N_616,In_418,In_687);
nand U617 (N_617,In_504,In_846);
and U618 (N_618,In_239,In_237);
nor U619 (N_619,In_559,In_691);
nor U620 (N_620,In_29,In_338);
nor U621 (N_621,In_364,In_792);
and U622 (N_622,In_108,In_382);
nand U623 (N_623,In_717,In_394);
and U624 (N_624,In_158,In_212);
nand U625 (N_625,In_714,In_846);
nand U626 (N_626,In_753,In_374);
or U627 (N_627,In_357,In_444);
nand U628 (N_628,In_361,In_114);
nor U629 (N_629,In_347,In_142);
nor U630 (N_630,In_948,In_981);
and U631 (N_631,In_465,In_436);
and U632 (N_632,In_450,In_203);
or U633 (N_633,In_913,In_234);
or U634 (N_634,In_759,In_708);
nand U635 (N_635,In_906,In_184);
nand U636 (N_636,In_830,In_794);
xor U637 (N_637,In_103,In_543);
nor U638 (N_638,In_392,In_736);
and U639 (N_639,In_783,In_480);
or U640 (N_640,In_450,In_921);
nor U641 (N_641,In_284,In_47);
or U642 (N_642,In_751,In_260);
and U643 (N_643,In_384,In_64);
or U644 (N_644,In_945,In_397);
or U645 (N_645,In_306,In_95);
nand U646 (N_646,In_397,In_578);
nor U647 (N_647,In_914,In_301);
nor U648 (N_648,In_928,In_394);
or U649 (N_649,In_949,In_407);
nor U650 (N_650,In_896,In_477);
nor U651 (N_651,In_413,In_484);
nand U652 (N_652,In_320,In_424);
and U653 (N_653,In_184,In_775);
and U654 (N_654,In_916,In_814);
nor U655 (N_655,In_19,In_265);
or U656 (N_656,In_887,In_272);
or U657 (N_657,In_799,In_668);
nor U658 (N_658,In_501,In_577);
or U659 (N_659,In_990,In_65);
and U660 (N_660,In_148,In_710);
or U661 (N_661,In_120,In_614);
and U662 (N_662,In_273,In_976);
and U663 (N_663,In_881,In_600);
and U664 (N_664,In_49,In_705);
and U665 (N_665,In_214,In_871);
or U666 (N_666,In_239,In_939);
nor U667 (N_667,In_32,In_187);
nor U668 (N_668,In_273,In_950);
and U669 (N_669,In_346,In_690);
or U670 (N_670,In_948,In_752);
nor U671 (N_671,In_489,In_887);
nand U672 (N_672,In_411,In_501);
or U673 (N_673,In_461,In_120);
nand U674 (N_674,In_96,In_645);
or U675 (N_675,In_293,In_46);
nand U676 (N_676,In_360,In_268);
or U677 (N_677,In_372,In_977);
nand U678 (N_678,In_0,In_441);
nand U679 (N_679,In_696,In_19);
or U680 (N_680,In_547,In_490);
nand U681 (N_681,In_303,In_631);
nand U682 (N_682,In_769,In_218);
nor U683 (N_683,In_775,In_166);
and U684 (N_684,In_703,In_704);
and U685 (N_685,In_640,In_787);
nor U686 (N_686,In_369,In_491);
nand U687 (N_687,In_413,In_692);
or U688 (N_688,In_23,In_508);
nor U689 (N_689,In_121,In_676);
and U690 (N_690,In_529,In_488);
nor U691 (N_691,In_994,In_951);
nor U692 (N_692,In_814,In_843);
nand U693 (N_693,In_728,In_528);
nor U694 (N_694,In_519,In_177);
nor U695 (N_695,In_580,In_498);
nand U696 (N_696,In_554,In_149);
nand U697 (N_697,In_135,In_782);
and U698 (N_698,In_882,In_842);
nand U699 (N_699,In_570,In_115);
nand U700 (N_700,In_606,In_597);
and U701 (N_701,In_139,In_624);
nor U702 (N_702,In_655,In_771);
nand U703 (N_703,In_997,In_198);
nor U704 (N_704,In_968,In_318);
nand U705 (N_705,In_722,In_500);
nor U706 (N_706,In_611,In_946);
or U707 (N_707,In_2,In_645);
nor U708 (N_708,In_342,In_17);
nor U709 (N_709,In_855,In_455);
nor U710 (N_710,In_175,In_232);
nor U711 (N_711,In_229,In_927);
or U712 (N_712,In_35,In_795);
nor U713 (N_713,In_198,In_853);
and U714 (N_714,In_141,In_380);
and U715 (N_715,In_836,In_104);
nand U716 (N_716,In_328,In_610);
nor U717 (N_717,In_723,In_27);
and U718 (N_718,In_229,In_11);
and U719 (N_719,In_605,In_709);
and U720 (N_720,In_520,In_217);
nand U721 (N_721,In_946,In_421);
nand U722 (N_722,In_947,In_684);
nand U723 (N_723,In_246,In_689);
nor U724 (N_724,In_345,In_976);
and U725 (N_725,In_618,In_277);
and U726 (N_726,In_923,In_772);
nor U727 (N_727,In_772,In_614);
nand U728 (N_728,In_475,In_600);
nand U729 (N_729,In_869,In_813);
or U730 (N_730,In_801,In_167);
or U731 (N_731,In_643,In_764);
nor U732 (N_732,In_715,In_194);
nand U733 (N_733,In_886,In_635);
nand U734 (N_734,In_885,In_683);
or U735 (N_735,In_648,In_550);
nor U736 (N_736,In_853,In_274);
nor U737 (N_737,In_472,In_743);
nand U738 (N_738,In_863,In_788);
or U739 (N_739,In_23,In_425);
nor U740 (N_740,In_916,In_448);
nor U741 (N_741,In_470,In_784);
nor U742 (N_742,In_453,In_445);
nand U743 (N_743,In_528,In_988);
and U744 (N_744,In_34,In_162);
and U745 (N_745,In_930,In_360);
nor U746 (N_746,In_541,In_597);
and U747 (N_747,In_682,In_551);
nand U748 (N_748,In_777,In_794);
or U749 (N_749,In_213,In_362);
or U750 (N_750,In_961,In_648);
or U751 (N_751,In_480,In_114);
or U752 (N_752,In_846,In_549);
nand U753 (N_753,In_171,In_752);
or U754 (N_754,In_240,In_834);
or U755 (N_755,In_534,In_66);
and U756 (N_756,In_216,In_710);
and U757 (N_757,In_450,In_791);
nor U758 (N_758,In_672,In_566);
and U759 (N_759,In_373,In_202);
and U760 (N_760,In_772,In_466);
nand U761 (N_761,In_349,In_942);
or U762 (N_762,In_72,In_686);
or U763 (N_763,In_445,In_656);
and U764 (N_764,In_826,In_71);
and U765 (N_765,In_545,In_483);
nor U766 (N_766,In_725,In_894);
and U767 (N_767,In_458,In_621);
nor U768 (N_768,In_386,In_845);
or U769 (N_769,In_725,In_825);
nor U770 (N_770,In_515,In_489);
or U771 (N_771,In_189,In_183);
and U772 (N_772,In_866,In_535);
and U773 (N_773,In_712,In_378);
nand U774 (N_774,In_549,In_349);
and U775 (N_775,In_697,In_232);
or U776 (N_776,In_642,In_181);
nand U777 (N_777,In_175,In_23);
and U778 (N_778,In_322,In_296);
nand U779 (N_779,In_998,In_989);
or U780 (N_780,In_869,In_537);
or U781 (N_781,In_850,In_814);
nor U782 (N_782,In_979,In_168);
or U783 (N_783,In_438,In_110);
nand U784 (N_784,In_922,In_24);
or U785 (N_785,In_107,In_775);
and U786 (N_786,In_779,In_692);
nor U787 (N_787,In_67,In_646);
or U788 (N_788,In_957,In_775);
and U789 (N_789,In_38,In_205);
nor U790 (N_790,In_664,In_219);
nand U791 (N_791,In_545,In_726);
or U792 (N_792,In_592,In_904);
and U793 (N_793,In_364,In_978);
and U794 (N_794,In_4,In_671);
nand U795 (N_795,In_16,In_499);
or U796 (N_796,In_926,In_122);
or U797 (N_797,In_598,In_995);
or U798 (N_798,In_462,In_40);
or U799 (N_799,In_470,In_580);
nor U800 (N_800,In_722,In_78);
or U801 (N_801,In_588,In_378);
nor U802 (N_802,In_742,In_107);
or U803 (N_803,In_845,In_189);
and U804 (N_804,In_294,In_972);
xnor U805 (N_805,In_281,In_177);
nor U806 (N_806,In_791,In_602);
or U807 (N_807,In_68,In_772);
nor U808 (N_808,In_908,In_718);
nor U809 (N_809,In_621,In_352);
or U810 (N_810,In_719,In_702);
or U811 (N_811,In_521,In_625);
xnor U812 (N_812,In_936,In_231);
nand U813 (N_813,In_996,In_823);
and U814 (N_814,In_270,In_474);
and U815 (N_815,In_518,In_596);
and U816 (N_816,In_834,In_372);
nand U817 (N_817,In_463,In_45);
and U818 (N_818,In_721,In_133);
nor U819 (N_819,In_674,In_328);
and U820 (N_820,In_492,In_590);
nand U821 (N_821,In_867,In_646);
and U822 (N_822,In_605,In_622);
and U823 (N_823,In_162,In_249);
nor U824 (N_824,In_996,In_284);
or U825 (N_825,In_238,In_997);
nor U826 (N_826,In_907,In_58);
and U827 (N_827,In_186,In_592);
nor U828 (N_828,In_887,In_687);
nand U829 (N_829,In_852,In_762);
or U830 (N_830,In_793,In_70);
and U831 (N_831,In_41,In_215);
or U832 (N_832,In_592,In_650);
and U833 (N_833,In_313,In_711);
or U834 (N_834,In_883,In_63);
and U835 (N_835,In_174,In_528);
nor U836 (N_836,In_311,In_469);
or U837 (N_837,In_32,In_355);
and U838 (N_838,In_826,In_408);
nand U839 (N_839,In_467,In_219);
nor U840 (N_840,In_253,In_614);
nand U841 (N_841,In_436,In_279);
nand U842 (N_842,In_159,In_84);
nand U843 (N_843,In_617,In_741);
nand U844 (N_844,In_573,In_511);
and U845 (N_845,In_538,In_669);
nor U846 (N_846,In_772,In_525);
or U847 (N_847,In_463,In_381);
and U848 (N_848,In_813,In_330);
or U849 (N_849,In_311,In_946);
xor U850 (N_850,In_16,In_714);
nand U851 (N_851,In_756,In_916);
nor U852 (N_852,In_692,In_759);
or U853 (N_853,In_309,In_847);
or U854 (N_854,In_480,In_299);
nor U855 (N_855,In_837,In_35);
and U856 (N_856,In_289,In_57);
or U857 (N_857,In_909,In_265);
or U858 (N_858,In_626,In_159);
or U859 (N_859,In_374,In_15);
nand U860 (N_860,In_800,In_280);
nor U861 (N_861,In_413,In_859);
or U862 (N_862,In_990,In_436);
and U863 (N_863,In_397,In_277);
or U864 (N_864,In_27,In_909);
nand U865 (N_865,In_386,In_539);
or U866 (N_866,In_904,In_27);
or U867 (N_867,In_364,In_572);
or U868 (N_868,In_393,In_993);
nor U869 (N_869,In_253,In_567);
nor U870 (N_870,In_8,In_127);
and U871 (N_871,In_444,In_112);
and U872 (N_872,In_261,In_151);
or U873 (N_873,In_790,In_838);
or U874 (N_874,In_515,In_406);
and U875 (N_875,In_226,In_480);
nor U876 (N_876,In_262,In_303);
nor U877 (N_877,In_368,In_74);
nor U878 (N_878,In_491,In_979);
and U879 (N_879,In_313,In_695);
nor U880 (N_880,In_160,In_420);
nor U881 (N_881,In_72,In_764);
or U882 (N_882,In_493,In_47);
nand U883 (N_883,In_201,In_475);
nand U884 (N_884,In_696,In_776);
and U885 (N_885,In_687,In_499);
or U886 (N_886,In_540,In_46);
nand U887 (N_887,In_466,In_906);
nand U888 (N_888,In_423,In_779);
nor U889 (N_889,In_377,In_60);
nor U890 (N_890,In_889,In_466);
nand U891 (N_891,In_833,In_377);
and U892 (N_892,In_437,In_966);
and U893 (N_893,In_255,In_569);
nor U894 (N_894,In_98,In_166);
nand U895 (N_895,In_443,In_665);
nor U896 (N_896,In_743,In_999);
and U897 (N_897,In_627,In_512);
and U898 (N_898,In_403,In_336);
nand U899 (N_899,In_655,In_315);
nor U900 (N_900,In_193,In_235);
or U901 (N_901,In_731,In_775);
nor U902 (N_902,In_324,In_295);
or U903 (N_903,In_369,In_28);
or U904 (N_904,In_38,In_309);
nor U905 (N_905,In_370,In_295);
and U906 (N_906,In_503,In_910);
or U907 (N_907,In_244,In_162);
nor U908 (N_908,In_830,In_442);
and U909 (N_909,In_377,In_508);
and U910 (N_910,In_671,In_51);
nor U911 (N_911,In_57,In_623);
nand U912 (N_912,In_860,In_924);
xor U913 (N_913,In_501,In_855);
xor U914 (N_914,In_956,In_814);
and U915 (N_915,In_813,In_223);
and U916 (N_916,In_857,In_532);
or U917 (N_917,In_103,In_660);
nor U918 (N_918,In_158,In_623);
and U919 (N_919,In_987,In_575);
and U920 (N_920,In_199,In_256);
nor U921 (N_921,In_488,In_145);
or U922 (N_922,In_294,In_33);
nor U923 (N_923,In_944,In_241);
nand U924 (N_924,In_82,In_253);
nand U925 (N_925,In_543,In_137);
nor U926 (N_926,In_443,In_476);
nand U927 (N_927,In_829,In_333);
nor U928 (N_928,In_741,In_485);
nand U929 (N_929,In_699,In_11);
or U930 (N_930,In_75,In_920);
nor U931 (N_931,In_858,In_94);
nand U932 (N_932,In_372,In_493);
or U933 (N_933,In_770,In_906);
nor U934 (N_934,In_432,In_640);
nand U935 (N_935,In_39,In_736);
nand U936 (N_936,In_303,In_122);
and U937 (N_937,In_786,In_936);
nor U938 (N_938,In_139,In_693);
nand U939 (N_939,In_214,In_636);
and U940 (N_940,In_841,In_637);
and U941 (N_941,In_600,In_298);
and U942 (N_942,In_605,In_937);
nor U943 (N_943,In_973,In_350);
nor U944 (N_944,In_918,In_508);
or U945 (N_945,In_676,In_712);
and U946 (N_946,In_382,In_473);
nor U947 (N_947,In_530,In_469);
and U948 (N_948,In_921,In_909);
nand U949 (N_949,In_398,In_275);
or U950 (N_950,In_415,In_404);
nand U951 (N_951,In_270,In_879);
nor U952 (N_952,In_221,In_533);
xor U953 (N_953,In_190,In_601);
nor U954 (N_954,In_345,In_950);
nand U955 (N_955,In_262,In_156);
nor U956 (N_956,In_645,In_820);
or U957 (N_957,In_2,In_302);
nand U958 (N_958,In_473,In_608);
and U959 (N_959,In_4,In_246);
or U960 (N_960,In_54,In_827);
or U961 (N_961,In_603,In_423);
nand U962 (N_962,In_474,In_941);
nor U963 (N_963,In_990,In_622);
and U964 (N_964,In_834,In_709);
nand U965 (N_965,In_895,In_505);
xor U966 (N_966,In_698,In_799);
or U967 (N_967,In_405,In_294);
nand U968 (N_968,In_80,In_686);
or U969 (N_969,In_450,In_579);
nor U970 (N_970,In_944,In_607);
or U971 (N_971,In_473,In_218);
nor U972 (N_972,In_161,In_857);
and U973 (N_973,In_275,In_79);
or U974 (N_974,In_371,In_494);
nand U975 (N_975,In_938,In_415);
nor U976 (N_976,In_918,In_356);
or U977 (N_977,In_910,In_403);
and U978 (N_978,In_703,In_722);
nand U979 (N_979,In_98,In_991);
or U980 (N_980,In_168,In_7);
or U981 (N_981,In_182,In_258);
nor U982 (N_982,In_315,In_279);
and U983 (N_983,In_590,In_575);
and U984 (N_984,In_464,In_940);
xor U985 (N_985,In_253,In_43);
nand U986 (N_986,In_515,In_807);
nor U987 (N_987,In_343,In_474);
nor U988 (N_988,In_184,In_945);
nor U989 (N_989,In_364,In_648);
or U990 (N_990,In_452,In_784);
and U991 (N_991,In_13,In_311);
and U992 (N_992,In_826,In_333);
and U993 (N_993,In_260,In_852);
or U994 (N_994,In_437,In_691);
nor U995 (N_995,In_297,In_293);
nand U996 (N_996,In_818,In_835);
or U997 (N_997,In_167,In_400);
and U998 (N_998,In_153,In_890);
or U999 (N_999,In_201,In_828);
or U1000 (N_1000,In_297,In_822);
nor U1001 (N_1001,In_632,In_453);
or U1002 (N_1002,In_618,In_759);
nor U1003 (N_1003,In_12,In_568);
nor U1004 (N_1004,In_666,In_114);
xnor U1005 (N_1005,In_188,In_449);
and U1006 (N_1006,In_667,In_119);
nand U1007 (N_1007,In_96,In_612);
nor U1008 (N_1008,In_909,In_930);
nor U1009 (N_1009,In_794,In_847);
and U1010 (N_1010,In_77,In_696);
nor U1011 (N_1011,In_264,In_514);
or U1012 (N_1012,In_346,In_320);
and U1013 (N_1013,In_336,In_652);
nand U1014 (N_1014,In_693,In_627);
and U1015 (N_1015,In_44,In_991);
or U1016 (N_1016,In_900,In_911);
and U1017 (N_1017,In_490,In_567);
nand U1018 (N_1018,In_492,In_845);
and U1019 (N_1019,In_965,In_832);
nand U1020 (N_1020,In_949,In_827);
nor U1021 (N_1021,In_130,In_81);
nand U1022 (N_1022,In_669,In_274);
nor U1023 (N_1023,In_62,In_997);
nor U1024 (N_1024,In_968,In_464);
and U1025 (N_1025,In_847,In_805);
nor U1026 (N_1026,In_85,In_531);
nand U1027 (N_1027,In_803,In_990);
nand U1028 (N_1028,In_828,In_753);
nand U1029 (N_1029,In_932,In_810);
and U1030 (N_1030,In_175,In_340);
and U1031 (N_1031,In_682,In_648);
nor U1032 (N_1032,In_41,In_717);
and U1033 (N_1033,In_32,In_600);
nand U1034 (N_1034,In_924,In_442);
nor U1035 (N_1035,In_50,In_233);
and U1036 (N_1036,In_764,In_506);
nand U1037 (N_1037,In_634,In_418);
and U1038 (N_1038,In_140,In_384);
nand U1039 (N_1039,In_357,In_770);
or U1040 (N_1040,In_697,In_596);
and U1041 (N_1041,In_792,In_887);
nand U1042 (N_1042,In_328,In_318);
or U1043 (N_1043,In_996,In_820);
or U1044 (N_1044,In_938,In_654);
and U1045 (N_1045,In_505,In_892);
nor U1046 (N_1046,In_826,In_581);
nor U1047 (N_1047,In_656,In_588);
xnor U1048 (N_1048,In_311,In_146);
and U1049 (N_1049,In_459,In_80);
or U1050 (N_1050,In_868,In_658);
and U1051 (N_1051,In_377,In_192);
and U1052 (N_1052,In_288,In_865);
nand U1053 (N_1053,In_897,In_61);
and U1054 (N_1054,In_469,In_878);
nand U1055 (N_1055,In_787,In_594);
nand U1056 (N_1056,In_504,In_376);
and U1057 (N_1057,In_610,In_379);
and U1058 (N_1058,In_782,In_384);
nor U1059 (N_1059,In_556,In_5);
nand U1060 (N_1060,In_410,In_740);
or U1061 (N_1061,In_62,In_620);
and U1062 (N_1062,In_955,In_803);
nor U1063 (N_1063,In_536,In_101);
and U1064 (N_1064,In_174,In_532);
nand U1065 (N_1065,In_654,In_304);
nand U1066 (N_1066,In_555,In_252);
nor U1067 (N_1067,In_840,In_606);
nor U1068 (N_1068,In_284,In_652);
nor U1069 (N_1069,In_110,In_750);
or U1070 (N_1070,In_729,In_802);
nor U1071 (N_1071,In_397,In_351);
xor U1072 (N_1072,In_330,In_591);
nor U1073 (N_1073,In_880,In_413);
nand U1074 (N_1074,In_506,In_108);
and U1075 (N_1075,In_492,In_127);
and U1076 (N_1076,In_203,In_417);
nor U1077 (N_1077,In_289,In_297);
or U1078 (N_1078,In_54,In_37);
and U1079 (N_1079,In_889,In_872);
nor U1080 (N_1080,In_243,In_756);
nor U1081 (N_1081,In_94,In_359);
or U1082 (N_1082,In_420,In_305);
or U1083 (N_1083,In_862,In_38);
xor U1084 (N_1084,In_657,In_892);
or U1085 (N_1085,In_635,In_808);
or U1086 (N_1086,In_354,In_39);
or U1087 (N_1087,In_620,In_317);
or U1088 (N_1088,In_740,In_582);
or U1089 (N_1089,In_804,In_55);
nor U1090 (N_1090,In_1,In_586);
and U1091 (N_1091,In_8,In_555);
nor U1092 (N_1092,In_433,In_828);
nor U1093 (N_1093,In_897,In_13);
nor U1094 (N_1094,In_997,In_101);
nand U1095 (N_1095,In_599,In_12);
and U1096 (N_1096,In_228,In_489);
or U1097 (N_1097,In_981,In_787);
and U1098 (N_1098,In_812,In_130);
xor U1099 (N_1099,In_951,In_964);
nand U1100 (N_1100,In_685,In_901);
or U1101 (N_1101,In_964,In_587);
nor U1102 (N_1102,In_477,In_624);
and U1103 (N_1103,In_560,In_810);
nor U1104 (N_1104,In_960,In_82);
nand U1105 (N_1105,In_442,In_568);
and U1106 (N_1106,In_194,In_135);
nand U1107 (N_1107,In_378,In_366);
and U1108 (N_1108,In_85,In_788);
nand U1109 (N_1109,In_617,In_275);
and U1110 (N_1110,In_110,In_924);
nor U1111 (N_1111,In_65,In_890);
and U1112 (N_1112,In_466,In_238);
nor U1113 (N_1113,In_415,In_194);
nand U1114 (N_1114,In_529,In_94);
or U1115 (N_1115,In_365,In_808);
and U1116 (N_1116,In_315,In_744);
or U1117 (N_1117,In_245,In_745);
and U1118 (N_1118,In_37,In_662);
nand U1119 (N_1119,In_196,In_580);
nand U1120 (N_1120,In_872,In_432);
nand U1121 (N_1121,In_245,In_505);
nand U1122 (N_1122,In_495,In_527);
xor U1123 (N_1123,In_440,In_236);
and U1124 (N_1124,In_366,In_683);
or U1125 (N_1125,In_986,In_366);
nand U1126 (N_1126,In_132,In_564);
nand U1127 (N_1127,In_891,In_915);
or U1128 (N_1128,In_937,In_286);
nor U1129 (N_1129,In_198,In_810);
or U1130 (N_1130,In_155,In_10);
or U1131 (N_1131,In_730,In_923);
or U1132 (N_1132,In_359,In_835);
and U1133 (N_1133,In_559,In_288);
nand U1134 (N_1134,In_360,In_42);
and U1135 (N_1135,In_121,In_946);
nor U1136 (N_1136,In_941,In_272);
nor U1137 (N_1137,In_65,In_290);
nor U1138 (N_1138,In_116,In_444);
or U1139 (N_1139,In_999,In_580);
nand U1140 (N_1140,In_857,In_729);
nor U1141 (N_1141,In_647,In_825);
and U1142 (N_1142,In_804,In_526);
xor U1143 (N_1143,In_674,In_507);
nor U1144 (N_1144,In_20,In_427);
or U1145 (N_1145,In_103,In_468);
nand U1146 (N_1146,In_257,In_690);
and U1147 (N_1147,In_249,In_331);
and U1148 (N_1148,In_597,In_294);
or U1149 (N_1149,In_437,In_147);
nor U1150 (N_1150,In_339,In_824);
and U1151 (N_1151,In_743,In_111);
and U1152 (N_1152,In_654,In_340);
and U1153 (N_1153,In_246,In_400);
and U1154 (N_1154,In_717,In_165);
or U1155 (N_1155,In_532,In_421);
or U1156 (N_1156,In_955,In_290);
or U1157 (N_1157,In_936,In_175);
or U1158 (N_1158,In_709,In_47);
or U1159 (N_1159,In_139,In_511);
and U1160 (N_1160,In_966,In_164);
nor U1161 (N_1161,In_805,In_592);
nand U1162 (N_1162,In_79,In_383);
nand U1163 (N_1163,In_703,In_591);
or U1164 (N_1164,In_90,In_119);
and U1165 (N_1165,In_560,In_113);
nor U1166 (N_1166,In_371,In_655);
nor U1167 (N_1167,In_14,In_664);
or U1168 (N_1168,In_712,In_465);
and U1169 (N_1169,In_788,In_796);
nand U1170 (N_1170,In_253,In_520);
nand U1171 (N_1171,In_956,In_751);
or U1172 (N_1172,In_142,In_367);
nand U1173 (N_1173,In_129,In_854);
nor U1174 (N_1174,In_549,In_324);
and U1175 (N_1175,In_726,In_954);
nand U1176 (N_1176,In_81,In_662);
nor U1177 (N_1177,In_327,In_797);
nand U1178 (N_1178,In_546,In_401);
nand U1179 (N_1179,In_686,In_861);
nor U1180 (N_1180,In_820,In_590);
nand U1181 (N_1181,In_816,In_587);
or U1182 (N_1182,In_538,In_750);
or U1183 (N_1183,In_357,In_729);
nand U1184 (N_1184,In_545,In_826);
and U1185 (N_1185,In_795,In_219);
or U1186 (N_1186,In_401,In_12);
and U1187 (N_1187,In_424,In_950);
or U1188 (N_1188,In_429,In_64);
nand U1189 (N_1189,In_462,In_473);
nor U1190 (N_1190,In_515,In_113);
nand U1191 (N_1191,In_82,In_662);
and U1192 (N_1192,In_466,In_615);
or U1193 (N_1193,In_58,In_527);
nand U1194 (N_1194,In_811,In_287);
or U1195 (N_1195,In_754,In_541);
nor U1196 (N_1196,In_850,In_771);
or U1197 (N_1197,In_546,In_425);
or U1198 (N_1198,In_685,In_697);
nand U1199 (N_1199,In_525,In_863);
nor U1200 (N_1200,In_423,In_854);
nand U1201 (N_1201,In_352,In_543);
nor U1202 (N_1202,In_645,In_719);
or U1203 (N_1203,In_37,In_299);
nor U1204 (N_1204,In_770,In_718);
or U1205 (N_1205,In_723,In_262);
nor U1206 (N_1206,In_671,In_903);
or U1207 (N_1207,In_967,In_799);
xnor U1208 (N_1208,In_77,In_919);
and U1209 (N_1209,In_515,In_788);
or U1210 (N_1210,In_299,In_961);
nor U1211 (N_1211,In_905,In_551);
or U1212 (N_1212,In_840,In_985);
nor U1213 (N_1213,In_154,In_368);
xnor U1214 (N_1214,In_662,In_206);
or U1215 (N_1215,In_431,In_304);
nand U1216 (N_1216,In_234,In_229);
nor U1217 (N_1217,In_170,In_682);
and U1218 (N_1218,In_516,In_182);
nor U1219 (N_1219,In_752,In_677);
and U1220 (N_1220,In_968,In_138);
nand U1221 (N_1221,In_763,In_124);
or U1222 (N_1222,In_673,In_718);
or U1223 (N_1223,In_549,In_111);
and U1224 (N_1224,In_760,In_852);
nand U1225 (N_1225,In_577,In_144);
and U1226 (N_1226,In_529,In_954);
nand U1227 (N_1227,In_603,In_316);
or U1228 (N_1228,In_780,In_418);
and U1229 (N_1229,In_782,In_195);
or U1230 (N_1230,In_745,In_647);
and U1231 (N_1231,In_615,In_702);
nand U1232 (N_1232,In_89,In_661);
nor U1233 (N_1233,In_649,In_556);
nand U1234 (N_1234,In_81,In_537);
nor U1235 (N_1235,In_972,In_977);
or U1236 (N_1236,In_53,In_571);
or U1237 (N_1237,In_792,In_609);
nand U1238 (N_1238,In_565,In_785);
or U1239 (N_1239,In_213,In_454);
and U1240 (N_1240,In_92,In_80);
nor U1241 (N_1241,In_468,In_236);
nor U1242 (N_1242,In_952,In_120);
or U1243 (N_1243,In_155,In_987);
nand U1244 (N_1244,In_629,In_657);
and U1245 (N_1245,In_320,In_551);
nor U1246 (N_1246,In_832,In_900);
nand U1247 (N_1247,In_927,In_108);
and U1248 (N_1248,In_233,In_385);
nor U1249 (N_1249,In_479,In_27);
or U1250 (N_1250,In_197,In_336);
nor U1251 (N_1251,In_750,In_397);
nor U1252 (N_1252,In_956,In_205);
or U1253 (N_1253,In_323,In_55);
or U1254 (N_1254,In_312,In_818);
or U1255 (N_1255,In_839,In_212);
nor U1256 (N_1256,In_666,In_339);
nor U1257 (N_1257,In_34,In_494);
nand U1258 (N_1258,In_53,In_970);
and U1259 (N_1259,In_778,In_37);
nand U1260 (N_1260,In_865,In_738);
and U1261 (N_1261,In_165,In_132);
or U1262 (N_1262,In_475,In_737);
and U1263 (N_1263,In_743,In_280);
and U1264 (N_1264,In_802,In_627);
or U1265 (N_1265,In_449,In_196);
and U1266 (N_1266,In_499,In_56);
or U1267 (N_1267,In_52,In_563);
nor U1268 (N_1268,In_289,In_612);
nand U1269 (N_1269,In_192,In_875);
or U1270 (N_1270,In_551,In_346);
nand U1271 (N_1271,In_374,In_197);
or U1272 (N_1272,In_390,In_452);
or U1273 (N_1273,In_395,In_730);
or U1274 (N_1274,In_722,In_715);
or U1275 (N_1275,In_825,In_180);
or U1276 (N_1276,In_908,In_273);
nand U1277 (N_1277,In_730,In_293);
or U1278 (N_1278,In_350,In_985);
nand U1279 (N_1279,In_796,In_621);
and U1280 (N_1280,In_387,In_77);
nand U1281 (N_1281,In_272,In_380);
or U1282 (N_1282,In_31,In_409);
nor U1283 (N_1283,In_798,In_636);
or U1284 (N_1284,In_606,In_443);
nand U1285 (N_1285,In_829,In_554);
nand U1286 (N_1286,In_326,In_788);
or U1287 (N_1287,In_762,In_707);
nor U1288 (N_1288,In_968,In_181);
nand U1289 (N_1289,In_124,In_791);
and U1290 (N_1290,In_124,In_870);
and U1291 (N_1291,In_320,In_783);
nor U1292 (N_1292,In_217,In_302);
nand U1293 (N_1293,In_489,In_423);
nand U1294 (N_1294,In_39,In_761);
nand U1295 (N_1295,In_343,In_249);
and U1296 (N_1296,In_412,In_651);
or U1297 (N_1297,In_679,In_346);
nand U1298 (N_1298,In_691,In_89);
or U1299 (N_1299,In_556,In_790);
and U1300 (N_1300,In_962,In_65);
and U1301 (N_1301,In_367,In_623);
nand U1302 (N_1302,In_776,In_999);
or U1303 (N_1303,In_857,In_320);
nand U1304 (N_1304,In_859,In_389);
or U1305 (N_1305,In_972,In_494);
nand U1306 (N_1306,In_4,In_167);
and U1307 (N_1307,In_253,In_413);
or U1308 (N_1308,In_275,In_238);
nand U1309 (N_1309,In_34,In_944);
nand U1310 (N_1310,In_256,In_137);
nor U1311 (N_1311,In_90,In_923);
nor U1312 (N_1312,In_471,In_828);
nand U1313 (N_1313,In_361,In_517);
and U1314 (N_1314,In_894,In_11);
and U1315 (N_1315,In_43,In_155);
and U1316 (N_1316,In_870,In_275);
and U1317 (N_1317,In_586,In_504);
or U1318 (N_1318,In_191,In_545);
and U1319 (N_1319,In_306,In_608);
xor U1320 (N_1320,In_222,In_3);
nand U1321 (N_1321,In_757,In_791);
nand U1322 (N_1322,In_388,In_619);
and U1323 (N_1323,In_822,In_866);
or U1324 (N_1324,In_858,In_106);
nor U1325 (N_1325,In_612,In_575);
and U1326 (N_1326,In_621,In_308);
nand U1327 (N_1327,In_995,In_355);
nor U1328 (N_1328,In_725,In_388);
and U1329 (N_1329,In_27,In_594);
and U1330 (N_1330,In_775,In_64);
nor U1331 (N_1331,In_544,In_997);
nor U1332 (N_1332,In_208,In_484);
and U1333 (N_1333,In_376,In_180);
and U1334 (N_1334,In_657,In_175);
or U1335 (N_1335,In_705,In_636);
nand U1336 (N_1336,In_126,In_452);
nand U1337 (N_1337,In_308,In_821);
and U1338 (N_1338,In_852,In_932);
and U1339 (N_1339,In_741,In_777);
nor U1340 (N_1340,In_218,In_231);
nor U1341 (N_1341,In_475,In_667);
or U1342 (N_1342,In_980,In_254);
or U1343 (N_1343,In_252,In_697);
nor U1344 (N_1344,In_145,In_645);
or U1345 (N_1345,In_526,In_579);
or U1346 (N_1346,In_476,In_55);
nand U1347 (N_1347,In_940,In_849);
or U1348 (N_1348,In_850,In_876);
nand U1349 (N_1349,In_323,In_296);
and U1350 (N_1350,In_216,In_677);
or U1351 (N_1351,In_668,In_318);
and U1352 (N_1352,In_854,In_791);
and U1353 (N_1353,In_356,In_579);
and U1354 (N_1354,In_775,In_405);
and U1355 (N_1355,In_786,In_458);
nand U1356 (N_1356,In_59,In_197);
nand U1357 (N_1357,In_442,In_816);
nor U1358 (N_1358,In_8,In_951);
and U1359 (N_1359,In_981,In_835);
nor U1360 (N_1360,In_334,In_162);
and U1361 (N_1361,In_68,In_522);
or U1362 (N_1362,In_163,In_368);
nand U1363 (N_1363,In_533,In_437);
and U1364 (N_1364,In_589,In_770);
or U1365 (N_1365,In_993,In_32);
nand U1366 (N_1366,In_734,In_698);
and U1367 (N_1367,In_250,In_385);
nand U1368 (N_1368,In_738,In_395);
or U1369 (N_1369,In_602,In_772);
and U1370 (N_1370,In_131,In_656);
and U1371 (N_1371,In_484,In_957);
and U1372 (N_1372,In_903,In_78);
xor U1373 (N_1373,In_733,In_825);
or U1374 (N_1374,In_600,In_198);
and U1375 (N_1375,In_236,In_175);
and U1376 (N_1376,In_260,In_934);
nand U1377 (N_1377,In_201,In_86);
and U1378 (N_1378,In_353,In_735);
nor U1379 (N_1379,In_205,In_987);
nor U1380 (N_1380,In_27,In_356);
nand U1381 (N_1381,In_865,In_153);
nor U1382 (N_1382,In_847,In_926);
and U1383 (N_1383,In_679,In_37);
nor U1384 (N_1384,In_81,In_447);
and U1385 (N_1385,In_457,In_280);
or U1386 (N_1386,In_260,In_218);
or U1387 (N_1387,In_92,In_710);
nor U1388 (N_1388,In_956,In_74);
nor U1389 (N_1389,In_111,In_342);
nand U1390 (N_1390,In_614,In_807);
or U1391 (N_1391,In_260,In_485);
nand U1392 (N_1392,In_586,In_246);
and U1393 (N_1393,In_531,In_365);
or U1394 (N_1394,In_560,In_435);
nor U1395 (N_1395,In_542,In_295);
nand U1396 (N_1396,In_287,In_92);
nor U1397 (N_1397,In_380,In_511);
or U1398 (N_1398,In_544,In_306);
nor U1399 (N_1399,In_853,In_270);
and U1400 (N_1400,In_736,In_965);
nor U1401 (N_1401,In_398,In_39);
and U1402 (N_1402,In_637,In_575);
nand U1403 (N_1403,In_845,In_148);
and U1404 (N_1404,In_729,In_741);
and U1405 (N_1405,In_99,In_871);
and U1406 (N_1406,In_326,In_910);
and U1407 (N_1407,In_853,In_137);
nand U1408 (N_1408,In_261,In_477);
or U1409 (N_1409,In_169,In_12);
and U1410 (N_1410,In_438,In_733);
nor U1411 (N_1411,In_29,In_348);
nand U1412 (N_1412,In_428,In_567);
nand U1413 (N_1413,In_152,In_318);
and U1414 (N_1414,In_601,In_107);
nor U1415 (N_1415,In_734,In_551);
or U1416 (N_1416,In_311,In_642);
or U1417 (N_1417,In_709,In_650);
nand U1418 (N_1418,In_669,In_445);
nor U1419 (N_1419,In_951,In_699);
nand U1420 (N_1420,In_239,In_589);
nor U1421 (N_1421,In_501,In_212);
xor U1422 (N_1422,In_899,In_147);
nor U1423 (N_1423,In_334,In_105);
nand U1424 (N_1424,In_586,In_816);
xor U1425 (N_1425,In_116,In_604);
nand U1426 (N_1426,In_138,In_136);
nand U1427 (N_1427,In_924,In_168);
nand U1428 (N_1428,In_575,In_276);
and U1429 (N_1429,In_215,In_354);
nor U1430 (N_1430,In_742,In_887);
and U1431 (N_1431,In_738,In_895);
or U1432 (N_1432,In_637,In_895);
nand U1433 (N_1433,In_207,In_499);
and U1434 (N_1434,In_555,In_332);
nand U1435 (N_1435,In_605,In_302);
nor U1436 (N_1436,In_697,In_410);
nor U1437 (N_1437,In_297,In_947);
or U1438 (N_1438,In_807,In_780);
and U1439 (N_1439,In_264,In_810);
and U1440 (N_1440,In_370,In_427);
and U1441 (N_1441,In_120,In_295);
or U1442 (N_1442,In_820,In_9);
nor U1443 (N_1443,In_283,In_697);
nor U1444 (N_1444,In_860,In_578);
and U1445 (N_1445,In_707,In_723);
nand U1446 (N_1446,In_927,In_345);
nand U1447 (N_1447,In_677,In_335);
and U1448 (N_1448,In_608,In_754);
and U1449 (N_1449,In_528,In_627);
or U1450 (N_1450,In_143,In_486);
or U1451 (N_1451,In_352,In_718);
nand U1452 (N_1452,In_509,In_651);
and U1453 (N_1453,In_887,In_967);
nand U1454 (N_1454,In_808,In_905);
and U1455 (N_1455,In_691,In_216);
nor U1456 (N_1456,In_620,In_277);
and U1457 (N_1457,In_286,In_280);
nand U1458 (N_1458,In_858,In_610);
nand U1459 (N_1459,In_841,In_88);
nor U1460 (N_1460,In_748,In_955);
and U1461 (N_1461,In_104,In_535);
or U1462 (N_1462,In_425,In_579);
and U1463 (N_1463,In_480,In_516);
xor U1464 (N_1464,In_926,In_229);
nor U1465 (N_1465,In_346,In_121);
and U1466 (N_1466,In_114,In_73);
or U1467 (N_1467,In_428,In_988);
and U1468 (N_1468,In_660,In_717);
nor U1469 (N_1469,In_298,In_284);
nand U1470 (N_1470,In_898,In_440);
and U1471 (N_1471,In_321,In_64);
nor U1472 (N_1472,In_270,In_525);
and U1473 (N_1473,In_759,In_65);
or U1474 (N_1474,In_628,In_245);
xnor U1475 (N_1475,In_621,In_149);
and U1476 (N_1476,In_628,In_433);
and U1477 (N_1477,In_389,In_952);
nor U1478 (N_1478,In_600,In_134);
or U1479 (N_1479,In_604,In_445);
or U1480 (N_1480,In_415,In_642);
nor U1481 (N_1481,In_208,In_687);
nand U1482 (N_1482,In_368,In_545);
nor U1483 (N_1483,In_995,In_997);
and U1484 (N_1484,In_609,In_984);
nor U1485 (N_1485,In_488,In_738);
nand U1486 (N_1486,In_882,In_983);
nand U1487 (N_1487,In_834,In_401);
nand U1488 (N_1488,In_810,In_211);
nor U1489 (N_1489,In_209,In_261);
and U1490 (N_1490,In_595,In_597);
or U1491 (N_1491,In_330,In_225);
nand U1492 (N_1492,In_911,In_994);
nand U1493 (N_1493,In_706,In_325);
nand U1494 (N_1494,In_62,In_713);
xnor U1495 (N_1495,In_272,In_327);
or U1496 (N_1496,In_813,In_106);
nor U1497 (N_1497,In_93,In_825);
nor U1498 (N_1498,In_583,In_962);
or U1499 (N_1499,In_82,In_829);
nand U1500 (N_1500,In_112,In_554);
or U1501 (N_1501,In_375,In_80);
nand U1502 (N_1502,In_415,In_138);
nor U1503 (N_1503,In_393,In_97);
nand U1504 (N_1504,In_409,In_829);
nor U1505 (N_1505,In_877,In_692);
xor U1506 (N_1506,In_954,In_265);
xnor U1507 (N_1507,In_830,In_991);
or U1508 (N_1508,In_539,In_883);
and U1509 (N_1509,In_803,In_128);
and U1510 (N_1510,In_823,In_612);
or U1511 (N_1511,In_865,In_930);
or U1512 (N_1512,In_559,In_243);
or U1513 (N_1513,In_412,In_199);
nor U1514 (N_1514,In_186,In_816);
nor U1515 (N_1515,In_548,In_683);
nand U1516 (N_1516,In_982,In_546);
and U1517 (N_1517,In_112,In_717);
nor U1518 (N_1518,In_417,In_408);
nor U1519 (N_1519,In_516,In_30);
or U1520 (N_1520,In_18,In_823);
or U1521 (N_1521,In_298,In_669);
nand U1522 (N_1522,In_897,In_90);
and U1523 (N_1523,In_957,In_996);
and U1524 (N_1524,In_212,In_586);
nand U1525 (N_1525,In_405,In_994);
nand U1526 (N_1526,In_660,In_210);
nor U1527 (N_1527,In_499,In_137);
nand U1528 (N_1528,In_681,In_474);
nand U1529 (N_1529,In_359,In_615);
and U1530 (N_1530,In_588,In_401);
nor U1531 (N_1531,In_470,In_466);
and U1532 (N_1532,In_532,In_988);
nand U1533 (N_1533,In_651,In_644);
nand U1534 (N_1534,In_681,In_420);
and U1535 (N_1535,In_932,In_800);
or U1536 (N_1536,In_34,In_197);
or U1537 (N_1537,In_964,In_864);
nand U1538 (N_1538,In_593,In_263);
or U1539 (N_1539,In_806,In_32);
nand U1540 (N_1540,In_650,In_414);
nor U1541 (N_1541,In_114,In_81);
or U1542 (N_1542,In_790,In_38);
and U1543 (N_1543,In_28,In_885);
or U1544 (N_1544,In_75,In_358);
nand U1545 (N_1545,In_949,In_682);
and U1546 (N_1546,In_10,In_106);
nor U1547 (N_1547,In_718,In_487);
nand U1548 (N_1548,In_183,In_49);
and U1549 (N_1549,In_730,In_21);
or U1550 (N_1550,In_803,In_627);
nand U1551 (N_1551,In_465,In_161);
and U1552 (N_1552,In_855,In_767);
nor U1553 (N_1553,In_346,In_199);
nand U1554 (N_1554,In_993,In_253);
and U1555 (N_1555,In_421,In_727);
nand U1556 (N_1556,In_814,In_813);
nand U1557 (N_1557,In_766,In_850);
or U1558 (N_1558,In_876,In_459);
and U1559 (N_1559,In_953,In_352);
or U1560 (N_1560,In_755,In_152);
nor U1561 (N_1561,In_150,In_233);
nor U1562 (N_1562,In_253,In_545);
and U1563 (N_1563,In_348,In_650);
nand U1564 (N_1564,In_323,In_843);
or U1565 (N_1565,In_227,In_733);
nor U1566 (N_1566,In_214,In_912);
nor U1567 (N_1567,In_827,In_112);
nor U1568 (N_1568,In_909,In_736);
nand U1569 (N_1569,In_484,In_490);
and U1570 (N_1570,In_321,In_884);
and U1571 (N_1571,In_514,In_69);
and U1572 (N_1572,In_259,In_237);
nand U1573 (N_1573,In_574,In_919);
nand U1574 (N_1574,In_838,In_899);
nand U1575 (N_1575,In_150,In_895);
and U1576 (N_1576,In_100,In_299);
and U1577 (N_1577,In_820,In_634);
nand U1578 (N_1578,In_213,In_502);
nor U1579 (N_1579,In_951,In_130);
or U1580 (N_1580,In_603,In_698);
or U1581 (N_1581,In_724,In_836);
and U1582 (N_1582,In_305,In_418);
and U1583 (N_1583,In_526,In_465);
or U1584 (N_1584,In_334,In_217);
or U1585 (N_1585,In_814,In_899);
nor U1586 (N_1586,In_373,In_138);
nand U1587 (N_1587,In_762,In_321);
and U1588 (N_1588,In_173,In_90);
nor U1589 (N_1589,In_513,In_755);
or U1590 (N_1590,In_211,In_571);
nor U1591 (N_1591,In_119,In_311);
and U1592 (N_1592,In_63,In_862);
nor U1593 (N_1593,In_296,In_986);
or U1594 (N_1594,In_648,In_458);
nor U1595 (N_1595,In_798,In_228);
nand U1596 (N_1596,In_76,In_929);
or U1597 (N_1597,In_725,In_276);
and U1598 (N_1598,In_353,In_943);
nor U1599 (N_1599,In_406,In_480);
and U1600 (N_1600,In_537,In_306);
nand U1601 (N_1601,In_733,In_125);
and U1602 (N_1602,In_540,In_43);
nor U1603 (N_1603,In_17,In_294);
and U1604 (N_1604,In_89,In_347);
or U1605 (N_1605,In_655,In_334);
and U1606 (N_1606,In_994,In_504);
or U1607 (N_1607,In_958,In_143);
and U1608 (N_1608,In_46,In_403);
or U1609 (N_1609,In_384,In_36);
nor U1610 (N_1610,In_731,In_761);
and U1611 (N_1611,In_946,In_987);
nand U1612 (N_1612,In_303,In_132);
nand U1613 (N_1613,In_675,In_910);
or U1614 (N_1614,In_661,In_261);
nand U1615 (N_1615,In_639,In_305);
and U1616 (N_1616,In_126,In_554);
and U1617 (N_1617,In_867,In_216);
nor U1618 (N_1618,In_789,In_40);
or U1619 (N_1619,In_357,In_59);
and U1620 (N_1620,In_875,In_698);
nor U1621 (N_1621,In_682,In_494);
nor U1622 (N_1622,In_764,In_640);
nor U1623 (N_1623,In_701,In_767);
nor U1624 (N_1624,In_414,In_211);
and U1625 (N_1625,In_966,In_896);
or U1626 (N_1626,In_114,In_410);
and U1627 (N_1627,In_557,In_863);
and U1628 (N_1628,In_3,In_97);
nand U1629 (N_1629,In_628,In_299);
and U1630 (N_1630,In_448,In_233);
or U1631 (N_1631,In_732,In_578);
and U1632 (N_1632,In_550,In_9);
nand U1633 (N_1633,In_281,In_829);
nor U1634 (N_1634,In_251,In_570);
and U1635 (N_1635,In_614,In_16);
nor U1636 (N_1636,In_466,In_722);
nand U1637 (N_1637,In_240,In_636);
nor U1638 (N_1638,In_535,In_71);
or U1639 (N_1639,In_380,In_990);
and U1640 (N_1640,In_814,In_902);
or U1641 (N_1641,In_243,In_444);
nor U1642 (N_1642,In_86,In_429);
and U1643 (N_1643,In_450,In_853);
nand U1644 (N_1644,In_24,In_586);
or U1645 (N_1645,In_845,In_586);
and U1646 (N_1646,In_977,In_962);
or U1647 (N_1647,In_702,In_129);
nand U1648 (N_1648,In_558,In_403);
and U1649 (N_1649,In_520,In_220);
and U1650 (N_1650,In_852,In_353);
nor U1651 (N_1651,In_363,In_318);
or U1652 (N_1652,In_107,In_264);
and U1653 (N_1653,In_413,In_929);
or U1654 (N_1654,In_523,In_928);
or U1655 (N_1655,In_220,In_597);
or U1656 (N_1656,In_671,In_122);
nand U1657 (N_1657,In_13,In_906);
and U1658 (N_1658,In_636,In_177);
nor U1659 (N_1659,In_289,In_809);
xor U1660 (N_1660,In_939,In_382);
nor U1661 (N_1661,In_123,In_565);
or U1662 (N_1662,In_830,In_284);
and U1663 (N_1663,In_82,In_334);
or U1664 (N_1664,In_647,In_979);
and U1665 (N_1665,In_485,In_815);
nor U1666 (N_1666,In_39,In_759);
or U1667 (N_1667,In_386,In_844);
or U1668 (N_1668,In_400,In_283);
nand U1669 (N_1669,In_258,In_913);
or U1670 (N_1670,In_152,In_280);
and U1671 (N_1671,In_89,In_771);
nand U1672 (N_1672,In_254,In_619);
nand U1673 (N_1673,In_246,In_58);
nand U1674 (N_1674,In_762,In_57);
or U1675 (N_1675,In_33,In_803);
nor U1676 (N_1676,In_739,In_790);
nor U1677 (N_1677,In_869,In_983);
nand U1678 (N_1678,In_860,In_572);
and U1679 (N_1679,In_893,In_327);
and U1680 (N_1680,In_123,In_303);
nor U1681 (N_1681,In_146,In_995);
or U1682 (N_1682,In_255,In_166);
nand U1683 (N_1683,In_680,In_276);
or U1684 (N_1684,In_488,In_39);
and U1685 (N_1685,In_410,In_353);
or U1686 (N_1686,In_569,In_616);
or U1687 (N_1687,In_501,In_92);
or U1688 (N_1688,In_962,In_646);
and U1689 (N_1689,In_37,In_148);
nor U1690 (N_1690,In_162,In_77);
or U1691 (N_1691,In_356,In_273);
and U1692 (N_1692,In_457,In_448);
and U1693 (N_1693,In_154,In_327);
or U1694 (N_1694,In_521,In_689);
nor U1695 (N_1695,In_529,In_265);
and U1696 (N_1696,In_127,In_819);
nand U1697 (N_1697,In_92,In_537);
or U1698 (N_1698,In_22,In_199);
nor U1699 (N_1699,In_863,In_922);
nor U1700 (N_1700,In_792,In_996);
and U1701 (N_1701,In_209,In_826);
nand U1702 (N_1702,In_361,In_108);
nor U1703 (N_1703,In_211,In_872);
or U1704 (N_1704,In_301,In_116);
or U1705 (N_1705,In_138,In_903);
nand U1706 (N_1706,In_531,In_321);
or U1707 (N_1707,In_701,In_71);
nand U1708 (N_1708,In_382,In_464);
and U1709 (N_1709,In_743,In_62);
or U1710 (N_1710,In_756,In_631);
nand U1711 (N_1711,In_555,In_875);
and U1712 (N_1712,In_596,In_960);
or U1713 (N_1713,In_634,In_838);
nand U1714 (N_1714,In_842,In_617);
and U1715 (N_1715,In_639,In_134);
nor U1716 (N_1716,In_46,In_816);
nand U1717 (N_1717,In_529,In_689);
or U1718 (N_1718,In_402,In_359);
or U1719 (N_1719,In_717,In_440);
and U1720 (N_1720,In_749,In_391);
nand U1721 (N_1721,In_531,In_441);
nor U1722 (N_1722,In_472,In_27);
or U1723 (N_1723,In_740,In_400);
nand U1724 (N_1724,In_320,In_205);
nor U1725 (N_1725,In_829,In_356);
nand U1726 (N_1726,In_839,In_651);
nand U1727 (N_1727,In_884,In_164);
and U1728 (N_1728,In_238,In_667);
nand U1729 (N_1729,In_335,In_246);
nor U1730 (N_1730,In_546,In_909);
or U1731 (N_1731,In_853,In_793);
and U1732 (N_1732,In_40,In_59);
nor U1733 (N_1733,In_425,In_987);
or U1734 (N_1734,In_714,In_877);
nand U1735 (N_1735,In_324,In_18);
nor U1736 (N_1736,In_680,In_752);
nand U1737 (N_1737,In_580,In_921);
and U1738 (N_1738,In_376,In_1);
and U1739 (N_1739,In_511,In_291);
and U1740 (N_1740,In_679,In_296);
nor U1741 (N_1741,In_331,In_300);
nor U1742 (N_1742,In_378,In_817);
and U1743 (N_1743,In_457,In_173);
nor U1744 (N_1744,In_691,In_596);
and U1745 (N_1745,In_784,In_682);
nor U1746 (N_1746,In_798,In_661);
nor U1747 (N_1747,In_608,In_207);
nand U1748 (N_1748,In_342,In_544);
or U1749 (N_1749,In_503,In_863);
and U1750 (N_1750,In_463,In_79);
and U1751 (N_1751,In_375,In_716);
nand U1752 (N_1752,In_269,In_947);
or U1753 (N_1753,In_566,In_208);
or U1754 (N_1754,In_35,In_491);
nor U1755 (N_1755,In_385,In_23);
or U1756 (N_1756,In_454,In_997);
nand U1757 (N_1757,In_284,In_874);
and U1758 (N_1758,In_179,In_149);
nand U1759 (N_1759,In_314,In_656);
nor U1760 (N_1760,In_215,In_746);
and U1761 (N_1761,In_213,In_63);
nand U1762 (N_1762,In_643,In_605);
nor U1763 (N_1763,In_715,In_453);
and U1764 (N_1764,In_956,In_578);
nor U1765 (N_1765,In_685,In_319);
xor U1766 (N_1766,In_766,In_714);
nor U1767 (N_1767,In_159,In_547);
nor U1768 (N_1768,In_780,In_806);
and U1769 (N_1769,In_410,In_552);
and U1770 (N_1770,In_430,In_631);
and U1771 (N_1771,In_88,In_588);
xor U1772 (N_1772,In_843,In_829);
or U1773 (N_1773,In_701,In_352);
or U1774 (N_1774,In_200,In_501);
and U1775 (N_1775,In_713,In_482);
nand U1776 (N_1776,In_18,In_675);
nor U1777 (N_1777,In_755,In_723);
nand U1778 (N_1778,In_960,In_438);
nand U1779 (N_1779,In_940,In_491);
and U1780 (N_1780,In_254,In_916);
or U1781 (N_1781,In_130,In_917);
and U1782 (N_1782,In_894,In_856);
and U1783 (N_1783,In_610,In_676);
or U1784 (N_1784,In_640,In_493);
or U1785 (N_1785,In_239,In_814);
nand U1786 (N_1786,In_475,In_370);
nand U1787 (N_1787,In_56,In_238);
nand U1788 (N_1788,In_280,In_503);
nor U1789 (N_1789,In_158,In_484);
or U1790 (N_1790,In_578,In_871);
nand U1791 (N_1791,In_652,In_58);
and U1792 (N_1792,In_18,In_335);
and U1793 (N_1793,In_540,In_298);
nand U1794 (N_1794,In_118,In_605);
nand U1795 (N_1795,In_164,In_124);
and U1796 (N_1796,In_431,In_802);
or U1797 (N_1797,In_467,In_533);
nor U1798 (N_1798,In_394,In_645);
and U1799 (N_1799,In_293,In_206);
nand U1800 (N_1800,In_640,In_375);
and U1801 (N_1801,In_607,In_433);
nand U1802 (N_1802,In_785,In_774);
nor U1803 (N_1803,In_736,In_669);
nand U1804 (N_1804,In_509,In_44);
nand U1805 (N_1805,In_249,In_488);
nor U1806 (N_1806,In_442,In_584);
xnor U1807 (N_1807,In_91,In_986);
nor U1808 (N_1808,In_489,In_989);
or U1809 (N_1809,In_443,In_673);
or U1810 (N_1810,In_776,In_284);
nand U1811 (N_1811,In_615,In_66);
nand U1812 (N_1812,In_802,In_202);
or U1813 (N_1813,In_237,In_344);
and U1814 (N_1814,In_841,In_843);
or U1815 (N_1815,In_776,In_646);
or U1816 (N_1816,In_978,In_871);
or U1817 (N_1817,In_309,In_119);
nor U1818 (N_1818,In_801,In_692);
and U1819 (N_1819,In_376,In_520);
nor U1820 (N_1820,In_337,In_814);
or U1821 (N_1821,In_458,In_143);
nand U1822 (N_1822,In_194,In_69);
and U1823 (N_1823,In_711,In_789);
nor U1824 (N_1824,In_276,In_813);
nand U1825 (N_1825,In_515,In_2);
nor U1826 (N_1826,In_373,In_870);
nor U1827 (N_1827,In_142,In_392);
nand U1828 (N_1828,In_542,In_44);
and U1829 (N_1829,In_158,In_619);
nand U1830 (N_1830,In_121,In_106);
or U1831 (N_1831,In_807,In_250);
nor U1832 (N_1832,In_919,In_196);
or U1833 (N_1833,In_731,In_308);
or U1834 (N_1834,In_443,In_361);
xor U1835 (N_1835,In_276,In_45);
nand U1836 (N_1836,In_506,In_168);
nor U1837 (N_1837,In_726,In_448);
nor U1838 (N_1838,In_405,In_742);
nor U1839 (N_1839,In_10,In_790);
nor U1840 (N_1840,In_664,In_615);
nand U1841 (N_1841,In_856,In_263);
nand U1842 (N_1842,In_367,In_781);
and U1843 (N_1843,In_408,In_998);
nor U1844 (N_1844,In_61,In_308);
and U1845 (N_1845,In_693,In_44);
or U1846 (N_1846,In_80,In_946);
nand U1847 (N_1847,In_149,In_535);
nor U1848 (N_1848,In_646,In_431);
and U1849 (N_1849,In_178,In_215);
nand U1850 (N_1850,In_979,In_1);
nand U1851 (N_1851,In_131,In_67);
nand U1852 (N_1852,In_753,In_106);
or U1853 (N_1853,In_518,In_356);
nor U1854 (N_1854,In_901,In_752);
or U1855 (N_1855,In_415,In_477);
nand U1856 (N_1856,In_983,In_497);
or U1857 (N_1857,In_493,In_112);
and U1858 (N_1858,In_664,In_708);
nand U1859 (N_1859,In_967,In_837);
nand U1860 (N_1860,In_965,In_143);
nor U1861 (N_1861,In_584,In_985);
nand U1862 (N_1862,In_615,In_970);
nor U1863 (N_1863,In_645,In_707);
nor U1864 (N_1864,In_812,In_141);
nand U1865 (N_1865,In_148,In_374);
and U1866 (N_1866,In_401,In_962);
and U1867 (N_1867,In_176,In_371);
and U1868 (N_1868,In_399,In_890);
or U1869 (N_1869,In_881,In_48);
nor U1870 (N_1870,In_368,In_303);
nor U1871 (N_1871,In_771,In_160);
nor U1872 (N_1872,In_131,In_47);
or U1873 (N_1873,In_302,In_4);
nor U1874 (N_1874,In_671,In_152);
nand U1875 (N_1875,In_116,In_373);
or U1876 (N_1876,In_613,In_841);
nand U1877 (N_1877,In_146,In_894);
and U1878 (N_1878,In_895,In_20);
nand U1879 (N_1879,In_937,In_385);
nor U1880 (N_1880,In_486,In_464);
nor U1881 (N_1881,In_183,In_157);
nor U1882 (N_1882,In_26,In_939);
and U1883 (N_1883,In_42,In_406);
or U1884 (N_1884,In_906,In_521);
and U1885 (N_1885,In_124,In_242);
nor U1886 (N_1886,In_706,In_288);
and U1887 (N_1887,In_77,In_37);
nand U1888 (N_1888,In_599,In_817);
nor U1889 (N_1889,In_972,In_799);
nand U1890 (N_1890,In_61,In_92);
nand U1891 (N_1891,In_319,In_24);
nand U1892 (N_1892,In_255,In_175);
or U1893 (N_1893,In_821,In_780);
nor U1894 (N_1894,In_969,In_319);
nand U1895 (N_1895,In_641,In_87);
nand U1896 (N_1896,In_483,In_924);
and U1897 (N_1897,In_625,In_648);
nand U1898 (N_1898,In_788,In_183);
and U1899 (N_1899,In_519,In_954);
nand U1900 (N_1900,In_800,In_73);
nand U1901 (N_1901,In_409,In_104);
nor U1902 (N_1902,In_318,In_553);
or U1903 (N_1903,In_156,In_492);
or U1904 (N_1904,In_433,In_581);
or U1905 (N_1905,In_769,In_271);
and U1906 (N_1906,In_801,In_277);
or U1907 (N_1907,In_646,In_898);
nor U1908 (N_1908,In_111,In_197);
and U1909 (N_1909,In_301,In_975);
and U1910 (N_1910,In_118,In_576);
nand U1911 (N_1911,In_763,In_547);
or U1912 (N_1912,In_535,In_248);
or U1913 (N_1913,In_550,In_888);
and U1914 (N_1914,In_191,In_829);
and U1915 (N_1915,In_732,In_280);
or U1916 (N_1916,In_545,In_113);
nor U1917 (N_1917,In_794,In_234);
nand U1918 (N_1918,In_783,In_215);
and U1919 (N_1919,In_314,In_732);
and U1920 (N_1920,In_46,In_925);
and U1921 (N_1921,In_338,In_653);
nand U1922 (N_1922,In_143,In_282);
nor U1923 (N_1923,In_338,In_129);
and U1924 (N_1924,In_74,In_953);
nor U1925 (N_1925,In_342,In_21);
or U1926 (N_1926,In_788,In_958);
or U1927 (N_1927,In_583,In_774);
and U1928 (N_1928,In_924,In_187);
nand U1929 (N_1929,In_617,In_53);
and U1930 (N_1930,In_521,In_608);
and U1931 (N_1931,In_734,In_169);
or U1932 (N_1932,In_379,In_221);
nand U1933 (N_1933,In_296,In_402);
nand U1934 (N_1934,In_273,In_959);
nor U1935 (N_1935,In_237,In_486);
or U1936 (N_1936,In_122,In_566);
and U1937 (N_1937,In_440,In_341);
nand U1938 (N_1938,In_499,In_561);
nor U1939 (N_1939,In_114,In_967);
nor U1940 (N_1940,In_260,In_200);
nor U1941 (N_1941,In_559,In_828);
nor U1942 (N_1942,In_591,In_465);
nand U1943 (N_1943,In_187,In_43);
and U1944 (N_1944,In_966,In_811);
nor U1945 (N_1945,In_297,In_549);
nand U1946 (N_1946,In_527,In_484);
or U1947 (N_1947,In_433,In_622);
nand U1948 (N_1948,In_141,In_505);
and U1949 (N_1949,In_933,In_932);
and U1950 (N_1950,In_386,In_104);
nor U1951 (N_1951,In_117,In_928);
nand U1952 (N_1952,In_514,In_175);
and U1953 (N_1953,In_177,In_654);
nor U1954 (N_1954,In_732,In_318);
or U1955 (N_1955,In_569,In_814);
or U1956 (N_1956,In_598,In_194);
or U1957 (N_1957,In_876,In_636);
or U1958 (N_1958,In_969,In_560);
or U1959 (N_1959,In_806,In_458);
or U1960 (N_1960,In_498,In_636);
nand U1961 (N_1961,In_967,In_862);
nor U1962 (N_1962,In_709,In_653);
nor U1963 (N_1963,In_597,In_908);
and U1964 (N_1964,In_671,In_364);
or U1965 (N_1965,In_794,In_356);
nor U1966 (N_1966,In_472,In_738);
or U1967 (N_1967,In_527,In_733);
nand U1968 (N_1968,In_180,In_289);
nand U1969 (N_1969,In_208,In_888);
and U1970 (N_1970,In_41,In_170);
and U1971 (N_1971,In_325,In_463);
and U1972 (N_1972,In_626,In_148);
nand U1973 (N_1973,In_813,In_82);
nand U1974 (N_1974,In_734,In_732);
and U1975 (N_1975,In_968,In_945);
or U1976 (N_1976,In_224,In_13);
and U1977 (N_1977,In_485,In_398);
and U1978 (N_1978,In_848,In_958);
nand U1979 (N_1979,In_260,In_981);
or U1980 (N_1980,In_465,In_309);
or U1981 (N_1981,In_978,In_879);
nand U1982 (N_1982,In_899,In_792);
or U1983 (N_1983,In_358,In_408);
nor U1984 (N_1984,In_915,In_527);
or U1985 (N_1985,In_959,In_722);
nor U1986 (N_1986,In_14,In_47);
nand U1987 (N_1987,In_578,In_239);
and U1988 (N_1988,In_970,In_314);
or U1989 (N_1989,In_120,In_711);
or U1990 (N_1990,In_853,In_861);
and U1991 (N_1991,In_570,In_806);
nand U1992 (N_1992,In_759,In_350);
nand U1993 (N_1993,In_261,In_506);
nand U1994 (N_1994,In_480,In_461);
or U1995 (N_1995,In_394,In_261);
nor U1996 (N_1996,In_834,In_107);
and U1997 (N_1997,In_961,In_495);
and U1998 (N_1998,In_716,In_679);
nor U1999 (N_1999,In_931,In_393);
or U2000 (N_2000,In_710,In_658);
nor U2001 (N_2001,In_27,In_513);
nand U2002 (N_2002,In_65,In_71);
and U2003 (N_2003,In_254,In_273);
nor U2004 (N_2004,In_737,In_42);
nand U2005 (N_2005,In_38,In_754);
nor U2006 (N_2006,In_859,In_933);
and U2007 (N_2007,In_136,In_541);
nor U2008 (N_2008,In_495,In_532);
or U2009 (N_2009,In_210,In_335);
or U2010 (N_2010,In_243,In_751);
nand U2011 (N_2011,In_885,In_589);
or U2012 (N_2012,In_787,In_991);
nor U2013 (N_2013,In_247,In_272);
or U2014 (N_2014,In_100,In_420);
nor U2015 (N_2015,In_230,In_754);
nor U2016 (N_2016,In_133,In_688);
and U2017 (N_2017,In_94,In_263);
nand U2018 (N_2018,In_23,In_526);
and U2019 (N_2019,In_430,In_744);
nor U2020 (N_2020,In_655,In_4);
nor U2021 (N_2021,In_997,In_147);
and U2022 (N_2022,In_695,In_224);
nand U2023 (N_2023,In_15,In_368);
and U2024 (N_2024,In_42,In_382);
and U2025 (N_2025,In_75,In_295);
nor U2026 (N_2026,In_979,In_605);
nand U2027 (N_2027,In_639,In_362);
nand U2028 (N_2028,In_554,In_197);
nand U2029 (N_2029,In_741,In_742);
or U2030 (N_2030,In_303,In_965);
or U2031 (N_2031,In_860,In_717);
or U2032 (N_2032,In_932,In_652);
nand U2033 (N_2033,In_739,In_638);
and U2034 (N_2034,In_383,In_889);
and U2035 (N_2035,In_633,In_322);
nand U2036 (N_2036,In_373,In_650);
nand U2037 (N_2037,In_826,In_460);
nand U2038 (N_2038,In_834,In_62);
nor U2039 (N_2039,In_366,In_217);
and U2040 (N_2040,In_141,In_152);
or U2041 (N_2041,In_508,In_600);
nand U2042 (N_2042,In_918,In_787);
and U2043 (N_2043,In_422,In_517);
or U2044 (N_2044,In_292,In_590);
nand U2045 (N_2045,In_883,In_975);
or U2046 (N_2046,In_234,In_838);
and U2047 (N_2047,In_536,In_843);
nor U2048 (N_2048,In_49,In_438);
or U2049 (N_2049,In_252,In_904);
and U2050 (N_2050,In_173,In_663);
or U2051 (N_2051,In_439,In_277);
or U2052 (N_2052,In_889,In_70);
and U2053 (N_2053,In_409,In_759);
nor U2054 (N_2054,In_909,In_66);
and U2055 (N_2055,In_772,In_156);
nor U2056 (N_2056,In_992,In_588);
or U2057 (N_2057,In_413,In_614);
nor U2058 (N_2058,In_634,In_387);
and U2059 (N_2059,In_378,In_708);
or U2060 (N_2060,In_42,In_744);
and U2061 (N_2061,In_50,In_245);
nor U2062 (N_2062,In_650,In_758);
and U2063 (N_2063,In_356,In_411);
nor U2064 (N_2064,In_863,In_802);
or U2065 (N_2065,In_150,In_581);
and U2066 (N_2066,In_159,In_679);
and U2067 (N_2067,In_633,In_90);
and U2068 (N_2068,In_564,In_849);
and U2069 (N_2069,In_99,In_645);
or U2070 (N_2070,In_420,In_996);
or U2071 (N_2071,In_559,In_710);
nor U2072 (N_2072,In_520,In_117);
or U2073 (N_2073,In_818,In_612);
nor U2074 (N_2074,In_904,In_78);
and U2075 (N_2075,In_315,In_588);
nor U2076 (N_2076,In_506,In_295);
and U2077 (N_2077,In_442,In_276);
and U2078 (N_2078,In_132,In_440);
nand U2079 (N_2079,In_103,In_829);
and U2080 (N_2080,In_188,In_347);
nand U2081 (N_2081,In_286,In_340);
nand U2082 (N_2082,In_488,In_261);
nor U2083 (N_2083,In_359,In_182);
or U2084 (N_2084,In_671,In_767);
and U2085 (N_2085,In_556,In_375);
and U2086 (N_2086,In_612,In_803);
or U2087 (N_2087,In_249,In_847);
or U2088 (N_2088,In_927,In_79);
or U2089 (N_2089,In_822,In_490);
nand U2090 (N_2090,In_853,In_168);
nand U2091 (N_2091,In_690,In_524);
nand U2092 (N_2092,In_419,In_977);
nor U2093 (N_2093,In_49,In_531);
or U2094 (N_2094,In_573,In_703);
nor U2095 (N_2095,In_786,In_707);
nor U2096 (N_2096,In_904,In_678);
nand U2097 (N_2097,In_364,In_437);
nor U2098 (N_2098,In_991,In_336);
or U2099 (N_2099,In_285,In_60);
nand U2100 (N_2100,In_882,In_128);
or U2101 (N_2101,In_360,In_808);
nand U2102 (N_2102,In_49,In_608);
nand U2103 (N_2103,In_978,In_900);
nand U2104 (N_2104,In_908,In_484);
nand U2105 (N_2105,In_832,In_829);
or U2106 (N_2106,In_82,In_250);
nand U2107 (N_2107,In_101,In_655);
nor U2108 (N_2108,In_90,In_341);
and U2109 (N_2109,In_161,In_698);
nand U2110 (N_2110,In_600,In_319);
or U2111 (N_2111,In_534,In_923);
and U2112 (N_2112,In_63,In_942);
and U2113 (N_2113,In_591,In_92);
and U2114 (N_2114,In_426,In_887);
nand U2115 (N_2115,In_35,In_600);
nand U2116 (N_2116,In_775,In_794);
nand U2117 (N_2117,In_516,In_200);
nand U2118 (N_2118,In_958,In_714);
nand U2119 (N_2119,In_128,In_540);
and U2120 (N_2120,In_211,In_871);
and U2121 (N_2121,In_34,In_810);
nand U2122 (N_2122,In_89,In_805);
and U2123 (N_2123,In_558,In_820);
and U2124 (N_2124,In_321,In_259);
nand U2125 (N_2125,In_74,In_601);
nor U2126 (N_2126,In_306,In_600);
and U2127 (N_2127,In_240,In_521);
nor U2128 (N_2128,In_915,In_817);
nand U2129 (N_2129,In_124,In_931);
or U2130 (N_2130,In_990,In_473);
or U2131 (N_2131,In_485,In_645);
or U2132 (N_2132,In_945,In_972);
nand U2133 (N_2133,In_608,In_15);
and U2134 (N_2134,In_459,In_313);
nand U2135 (N_2135,In_617,In_163);
or U2136 (N_2136,In_398,In_747);
or U2137 (N_2137,In_201,In_879);
and U2138 (N_2138,In_262,In_540);
and U2139 (N_2139,In_326,In_294);
nand U2140 (N_2140,In_703,In_11);
nand U2141 (N_2141,In_6,In_433);
and U2142 (N_2142,In_678,In_997);
nand U2143 (N_2143,In_92,In_585);
and U2144 (N_2144,In_6,In_898);
nor U2145 (N_2145,In_396,In_726);
and U2146 (N_2146,In_380,In_558);
nor U2147 (N_2147,In_753,In_30);
nand U2148 (N_2148,In_31,In_308);
nor U2149 (N_2149,In_790,In_828);
nor U2150 (N_2150,In_228,In_481);
nor U2151 (N_2151,In_358,In_350);
nor U2152 (N_2152,In_464,In_837);
or U2153 (N_2153,In_445,In_778);
and U2154 (N_2154,In_515,In_42);
nor U2155 (N_2155,In_490,In_469);
nor U2156 (N_2156,In_7,In_125);
nand U2157 (N_2157,In_643,In_42);
nand U2158 (N_2158,In_117,In_968);
nor U2159 (N_2159,In_869,In_658);
xor U2160 (N_2160,In_301,In_504);
nor U2161 (N_2161,In_612,In_22);
or U2162 (N_2162,In_424,In_539);
and U2163 (N_2163,In_651,In_755);
and U2164 (N_2164,In_389,In_20);
or U2165 (N_2165,In_480,In_169);
or U2166 (N_2166,In_318,In_705);
nor U2167 (N_2167,In_296,In_644);
nand U2168 (N_2168,In_162,In_353);
nand U2169 (N_2169,In_761,In_678);
nor U2170 (N_2170,In_200,In_902);
or U2171 (N_2171,In_918,In_223);
and U2172 (N_2172,In_715,In_853);
and U2173 (N_2173,In_46,In_955);
or U2174 (N_2174,In_872,In_47);
and U2175 (N_2175,In_601,In_725);
nor U2176 (N_2176,In_293,In_340);
nor U2177 (N_2177,In_747,In_938);
or U2178 (N_2178,In_873,In_496);
and U2179 (N_2179,In_967,In_606);
or U2180 (N_2180,In_906,In_309);
nor U2181 (N_2181,In_606,In_158);
and U2182 (N_2182,In_539,In_676);
or U2183 (N_2183,In_298,In_556);
nor U2184 (N_2184,In_167,In_471);
or U2185 (N_2185,In_873,In_485);
nor U2186 (N_2186,In_925,In_610);
or U2187 (N_2187,In_907,In_542);
nor U2188 (N_2188,In_92,In_74);
nand U2189 (N_2189,In_537,In_343);
or U2190 (N_2190,In_152,In_389);
and U2191 (N_2191,In_909,In_181);
nand U2192 (N_2192,In_789,In_23);
nand U2193 (N_2193,In_615,In_83);
nand U2194 (N_2194,In_476,In_281);
nand U2195 (N_2195,In_679,In_894);
or U2196 (N_2196,In_376,In_499);
nor U2197 (N_2197,In_106,In_842);
nand U2198 (N_2198,In_987,In_738);
nand U2199 (N_2199,In_96,In_754);
nand U2200 (N_2200,In_350,In_551);
or U2201 (N_2201,In_650,In_782);
or U2202 (N_2202,In_187,In_160);
or U2203 (N_2203,In_551,In_520);
nor U2204 (N_2204,In_523,In_283);
nand U2205 (N_2205,In_659,In_747);
and U2206 (N_2206,In_962,In_174);
nand U2207 (N_2207,In_168,In_529);
or U2208 (N_2208,In_453,In_226);
and U2209 (N_2209,In_99,In_859);
nor U2210 (N_2210,In_368,In_123);
and U2211 (N_2211,In_709,In_238);
or U2212 (N_2212,In_240,In_649);
nand U2213 (N_2213,In_602,In_570);
or U2214 (N_2214,In_117,In_499);
and U2215 (N_2215,In_713,In_645);
or U2216 (N_2216,In_384,In_505);
and U2217 (N_2217,In_230,In_972);
nor U2218 (N_2218,In_179,In_652);
and U2219 (N_2219,In_621,In_147);
or U2220 (N_2220,In_299,In_369);
or U2221 (N_2221,In_689,In_114);
nor U2222 (N_2222,In_864,In_513);
and U2223 (N_2223,In_997,In_240);
nor U2224 (N_2224,In_221,In_394);
and U2225 (N_2225,In_871,In_798);
or U2226 (N_2226,In_616,In_552);
nor U2227 (N_2227,In_586,In_167);
nand U2228 (N_2228,In_716,In_509);
and U2229 (N_2229,In_839,In_899);
xnor U2230 (N_2230,In_945,In_231);
or U2231 (N_2231,In_954,In_477);
nand U2232 (N_2232,In_897,In_754);
nor U2233 (N_2233,In_612,In_434);
and U2234 (N_2234,In_503,In_253);
nor U2235 (N_2235,In_874,In_93);
and U2236 (N_2236,In_132,In_629);
and U2237 (N_2237,In_653,In_251);
or U2238 (N_2238,In_717,In_30);
or U2239 (N_2239,In_182,In_722);
or U2240 (N_2240,In_441,In_758);
and U2241 (N_2241,In_499,In_106);
and U2242 (N_2242,In_409,In_645);
xnor U2243 (N_2243,In_397,In_732);
nand U2244 (N_2244,In_444,In_234);
and U2245 (N_2245,In_591,In_297);
nor U2246 (N_2246,In_340,In_827);
or U2247 (N_2247,In_354,In_375);
and U2248 (N_2248,In_62,In_460);
nand U2249 (N_2249,In_191,In_810);
nand U2250 (N_2250,In_347,In_796);
and U2251 (N_2251,In_833,In_205);
or U2252 (N_2252,In_441,In_830);
nor U2253 (N_2253,In_187,In_457);
nand U2254 (N_2254,In_619,In_803);
or U2255 (N_2255,In_154,In_743);
and U2256 (N_2256,In_789,In_378);
and U2257 (N_2257,In_807,In_797);
or U2258 (N_2258,In_103,In_646);
and U2259 (N_2259,In_59,In_7);
or U2260 (N_2260,In_319,In_873);
or U2261 (N_2261,In_204,In_704);
nand U2262 (N_2262,In_539,In_959);
nand U2263 (N_2263,In_832,In_88);
or U2264 (N_2264,In_542,In_103);
and U2265 (N_2265,In_561,In_643);
and U2266 (N_2266,In_208,In_958);
nor U2267 (N_2267,In_781,In_868);
and U2268 (N_2268,In_867,In_101);
and U2269 (N_2269,In_643,In_40);
nand U2270 (N_2270,In_57,In_471);
or U2271 (N_2271,In_152,In_126);
nand U2272 (N_2272,In_60,In_595);
or U2273 (N_2273,In_724,In_363);
nor U2274 (N_2274,In_724,In_526);
nor U2275 (N_2275,In_619,In_651);
or U2276 (N_2276,In_5,In_596);
nand U2277 (N_2277,In_821,In_803);
or U2278 (N_2278,In_298,In_955);
and U2279 (N_2279,In_537,In_205);
nor U2280 (N_2280,In_934,In_305);
or U2281 (N_2281,In_703,In_336);
or U2282 (N_2282,In_617,In_995);
and U2283 (N_2283,In_296,In_12);
or U2284 (N_2284,In_320,In_914);
nand U2285 (N_2285,In_502,In_56);
or U2286 (N_2286,In_576,In_922);
nor U2287 (N_2287,In_415,In_770);
or U2288 (N_2288,In_140,In_457);
nor U2289 (N_2289,In_198,In_575);
and U2290 (N_2290,In_276,In_757);
and U2291 (N_2291,In_797,In_338);
and U2292 (N_2292,In_863,In_589);
nor U2293 (N_2293,In_511,In_847);
nand U2294 (N_2294,In_516,In_949);
and U2295 (N_2295,In_770,In_118);
or U2296 (N_2296,In_870,In_893);
nand U2297 (N_2297,In_16,In_446);
nor U2298 (N_2298,In_644,In_117);
and U2299 (N_2299,In_558,In_496);
and U2300 (N_2300,In_108,In_306);
and U2301 (N_2301,In_27,In_550);
nand U2302 (N_2302,In_687,In_140);
or U2303 (N_2303,In_153,In_487);
nand U2304 (N_2304,In_209,In_358);
and U2305 (N_2305,In_891,In_192);
nand U2306 (N_2306,In_643,In_233);
xnor U2307 (N_2307,In_257,In_267);
nand U2308 (N_2308,In_725,In_123);
or U2309 (N_2309,In_131,In_254);
and U2310 (N_2310,In_778,In_437);
or U2311 (N_2311,In_651,In_406);
and U2312 (N_2312,In_294,In_2);
or U2313 (N_2313,In_49,In_686);
nor U2314 (N_2314,In_33,In_827);
and U2315 (N_2315,In_552,In_795);
nand U2316 (N_2316,In_660,In_427);
or U2317 (N_2317,In_115,In_947);
and U2318 (N_2318,In_82,In_6);
and U2319 (N_2319,In_603,In_851);
or U2320 (N_2320,In_399,In_123);
and U2321 (N_2321,In_831,In_196);
and U2322 (N_2322,In_252,In_277);
and U2323 (N_2323,In_834,In_523);
and U2324 (N_2324,In_763,In_1);
nor U2325 (N_2325,In_606,In_125);
and U2326 (N_2326,In_233,In_878);
and U2327 (N_2327,In_299,In_488);
and U2328 (N_2328,In_485,In_119);
or U2329 (N_2329,In_135,In_118);
nor U2330 (N_2330,In_789,In_35);
and U2331 (N_2331,In_312,In_354);
nor U2332 (N_2332,In_544,In_110);
nor U2333 (N_2333,In_242,In_114);
nand U2334 (N_2334,In_62,In_747);
and U2335 (N_2335,In_708,In_889);
and U2336 (N_2336,In_524,In_490);
nand U2337 (N_2337,In_432,In_180);
and U2338 (N_2338,In_591,In_796);
nand U2339 (N_2339,In_36,In_288);
or U2340 (N_2340,In_318,In_378);
nor U2341 (N_2341,In_184,In_449);
and U2342 (N_2342,In_861,In_852);
nand U2343 (N_2343,In_564,In_964);
or U2344 (N_2344,In_350,In_50);
and U2345 (N_2345,In_936,In_959);
nand U2346 (N_2346,In_854,In_627);
nor U2347 (N_2347,In_813,In_658);
nand U2348 (N_2348,In_373,In_628);
nor U2349 (N_2349,In_156,In_716);
and U2350 (N_2350,In_488,In_177);
or U2351 (N_2351,In_381,In_540);
nand U2352 (N_2352,In_318,In_853);
nor U2353 (N_2353,In_568,In_493);
and U2354 (N_2354,In_186,In_66);
and U2355 (N_2355,In_202,In_912);
or U2356 (N_2356,In_680,In_25);
or U2357 (N_2357,In_79,In_788);
nand U2358 (N_2358,In_756,In_300);
and U2359 (N_2359,In_80,In_859);
and U2360 (N_2360,In_188,In_996);
and U2361 (N_2361,In_560,In_24);
and U2362 (N_2362,In_932,In_499);
nor U2363 (N_2363,In_425,In_703);
and U2364 (N_2364,In_899,In_576);
nand U2365 (N_2365,In_256,In_337);
nand U2366 (N_2366,In_149,In_317);
and U2367 (N_2367,In_690,In_179);
nand U2368 (N_2368,In_577,In_408);
or U2369 (N_2369,In_303,In_170);
or U2370 (N_2370,In_854,In_455);
nor U2371 (N_2371,In_300,In_587);
and U2372 (N_2372,In_720,In_979);
nand U2373 (N_2373,In_54,In_585);
nor U2374 (N_2374,In_344,In_934);
or U2375 (N_2375,In_200,In_523);
xor U2376 (N_2376,In_554,In_468);
or U2377 (N_2377,In_663,In_271);
or U2378 (N_2378,In_392,In_595);
nand U2379 (N_2379,In_789,In_211);
and U2380 (N_2380,In_55,In_493);
nand U2381 (N_2381,In_155,In_412);
or U2382 (N_2382,In_427,In_206);
nor U2383 (N_2383,In_970,In_227);
or U2384 (N_2384,In_267,In_185);
and U2385 (N_2385,In_729,In_7);
or U2386 (N_2386,In_443,In_541);
nor U2387 (N_2387,In_327,In_34);
nor U2388 (N_2388,In_560,In_879);
and U2389 (N_2389,In_909,In_578);
and U2390 (N_2390,In_399,In_415);
and U2391 (N_2391,In_229,In_958);
nor U2392 (N_2392,In_34,In_703);
nor U2393 (N_2393,In_350,In_614);
or U2394 (N_2394,In_328,In_675);
or U2395 (N_2395,In_97,In_187);
nand U2396 (N_2396,In_120,In_681);
or U2397 (N_2397,In_66,In_220);
or U2398 (N_2398,In_227,In_673);
nand U2399 (N_2399,In_15,In_808);
nor U2400 (N_2400,In_27,In_996);
or U2401 (N_2401,In_339,In_407);
nor U2402 (N_2402,In_466,In_883);
nand U2403 (N_2403,In_960,In_792);
or U2404 (N_2404,In_780,In_344);
or U2405 (N_2405,In_259,In_435);
xor U2406 (N_2406,In_149,In_28);
and U2407 (N_2407,In_307,In_955);
or U2408 (N_2408,In_963,In_529);
or U2409 (N_2409,In_578,In_105);
or U2410 (N_2410,In_688,In_923);
or U2411 (N_2411,In_114,In_99);
nor U2412 (N_2412,In_184,In_316);
nand U2413 (N_2413,In_837,In_174);
nor U2414 (N_2414,In_937,In_856);
or U2415 (N_2415,In_55,In_131);
nor U2416 (N_2416,In_974,In_222);
nand U2417 (N_2417,In_722,In_567);
or U2418 (N_2418,In_938,In_426);
or U2419 (N_2419,In_410,In_670);
nand U2420 (N_2420,In_260,In_940);
or U2421 (N_2421,In_121,In_215);
nand U2422 (N_2422,In_551,In_412);
and U2423 (N_2423,In_807,In_496);
and U2424 (N_2424,In_242,In_407);
and U2425 (N_2425,In_155,In_367);
nor U2426 (N_2426,In_798,In_499);
nand U2427 (N_2427,In_376,In_20);
or U2428 (N_2428,In_355,In_385);
nand U2429 (N_2429,In_975,In_929);
nand U2430 (N_2430,In_480,In_951);
nand U2431 (N_2431,In_374,In_513);
nand U2432 (N_2432,In_545,In_252);
nand U2433 (N_2433,In_122,In_477);
nand U2434 (N_2434,In_605,In_703);
and U2435 (N_2435,In_595,In_566);
or U2436 (N_2436,In_736,In_822);
or U2437 (N_2437,In_861,In_21);
or U2438 (N_2438,In_91,In_597);
or U2439 (N_2439,In_421,In_216);
or U2440 (N_2440,In_180,In_890);
xor U2441 (N_2441,In_535,In_209);
and U2442 (N_2442,In_504,In_621);
nand U2443 (N_2443,In_673,In_166);
or U2444 (N_2444,In_277,In_43);
or U2445 (N_2445,In_842,In_633);
nand U2446 (N_2446,In_795,In_213);
and U2447 (N_2447,In_224,In_756);
and U2448 (N_2448,In_858,In_757);
nor U2449 (N_2449,In_292,In_81);
or U2450 (N_2450,In_103,In_359);
nor U2451 (N_2451,In_961,In_732);
nor U2452 (N_2452,In_86,In_420);
nand U2453 (N_2453,In_833,In_996);
nand U2454 (N_2454,In_833,In_68);
and U2455 (N_2455,In_177,In_753);
nor U2456 (N_2456,In_512,In_450);
and U2457 (N_2457,In_502,In_893);
nor U2458 (N_2458,In_103,In_919);
nor U2459 (N_2459,In_516,In_278);
and U2460 (N_2460,In_564,In_118);
nor U2461 (N_2461,In_149,In_46);
and U2462 (N_2462,In_839,In_895);
or U2463 (N_2463,In_638,In_362);
nor U2464 (N_2464,In_58,In_604);
or U2465 (N_2465,In_796,In_367);
and U2466 (N_2466,In_520,In_49);
or U2467 (N_2467,In_43,In_185);
nand U2468 (N_2468,In_765,In_297);
or U2469 (N_2469,In_529,In_676);
and U2470 (N_2470,In_766,In_832);
nor U2471 (N_2471,In_45,In_894);
nand U2472 (N_2472,In_720,In_518);
nand U2473 (N_2473,In_252,In_623);
and U2474 (N_2474,In_319,In_952);
nand U2475 (N_2475,In_0,In_879);
and U2476 (N_2476,In_118,In_385);
nand U2477 (N_2477,In_48,In_779);
or U2478 (N_2478,In_714,In_143);
nand U2479 (N_2479,In_855,In_417);
nor U2480 (N_2480,In_95,In_110);
or U2481 (N_2481,In_713,In_110);
nor U2482 (N_2482,In_851,In_968);
nand U2483 (N_2483,In_12,In_572);
nand U2484 (N_2484,In_905,In_103);
nor U2485 (N_2485,In_140,In_601);
nand U2486 (N_2486,In_209,In_419);
and U2487 (N_2487,In_189,In_324);
nor U2488 (N_2488,In_766,In_224);
nor U2489 (N_2489,In_614,In_955);
nor U2490 (N_2490,In_117,In_932);
nor U2491 (N_2491,In_271,In_111);
or U2492 (N_2492,In_611,In_913);
nor U2493 (N_2493,In_199,In_699);
or U2494 (N_2494,In_177,In_797);
or U2495 (N_2495,In_661,In_449);
or U2496 (N_2496,In_90,In_237);
or U2497 (N_2497,In_688,In_201);
and U2498 (N_2498,In_625,In_280);
and U2499 (N_2499,In_397,In_577);
nand U2500 (N_2500,In_309,In_286);
and U2501 (N_2501,In_321,In_896);
and U2502 (N_2502,In_499,In_976);
and U2503 (N_2503,In_6,In_746);
nor U2504 (N_2504,In_272,In_10);
nor U2505 (N_2505,In_860,In_53);
or U2506 (N_2506,In_904,In_338);
and U2507 (N_2507,In_942,In_288);
and U2508 (N_2508,In_934,In_493);
and U2509 (N_2509,In_432,In_823);
or U2510 (N_2510,In_930,In_436);
and U2511 (N_2511,In_443,In_13);
or U2512 (N_2512,In_995,In_170);
nand U2513 (N_2513,In_2,In_721);
xor U2514 (N_2514,In_437,In_146);
nand U2515 (N_2515,In_861,In_195);
nor U2516 (N_2516,In_374,In_808);
nor U2517 (N_2517,In_623,In_581);
and U2518 (N_2518,In_834,In_348);
and U2519 (N_2519,In_762,In_574);
nor U2520 (N_2520,In_41,In_174);
or U2521 (N_2521,In_299,In_19);
nor U2522 (N_2522,In_766,In_520);
nor U2523 (N_2523,In_838,In_851);
and U2524 (N_2524,In_64,In_871);
nand U2525 (N_2525,In_891,In_295);
nor U2526 (N_2526,In_16,In_272);
or U2527 (N_2527,In_775,In_916);
or U2528 (N_2528,In_3,In_106);
or U2529 (N_2529,In_849,In_149);
nand U2530 (N_2530,In_969,In_248);
nor U2531 (N_2531,In_835,In_396);
or U2532 (N_2532,In_845,In_264);
nand U2533 (N_2533,In_747,In_112);
nand U2534 (N_2534,In_449,In_82);
nand U2535 (N_2535,In_821,In_652);
nor U2536 (N_2536,In_349,In_327);
nor U2537 (N_2537,In_660,In_796);
nor U2538 (N_2538,In_571,In_145);
and U2539 (N_2539,In_382,In_452);
or U2540 (N_2540,In_8,In_599);
xnor U2541 (N_2541,In_206,In_17);
nor U2542 (N_2542,In_989,In_551);
xnor U2543 (N_2543,In_982,In_405);
nand U2544 (N_2544,In_511,In_303);
nand U2545 (N_2545,In_62,In_320);
nor U2546 (N_2546,In_476,In_350);
nor U2547 (N_2547,In_235,In_145);
nand U2548 (N_2548,In_510,In_359);
nor U2549 (N_2549,In_506,In_898);
and U2550 (N_2550,In_557,In_238);
or U2551 (N_2551,In_1,In_686);
and U2552 (N_2552,In_507,In_571);
nor U2553 (N_2553,In_889,In_677);
nand U2554 (N_2554,In_166,In_425);
nor U2555 (N_2555,In_297,In_966);
nand U2556 (N_2556,In_234,In_608);
nor U2557 (N_2557,In_200,In_81);
or U2558 (N_2558,In_750,In_572);
nand U2559 (N_2559,In_288,In_387);
nor U2560 (N_2560,In_627,In_976);
or U2561 (N_2561,In_44,In_719);
nor U2562 (N_2562,In_38,In_382);
nor U2563 (N_2563,In_986,In_576);
nor U2564 (N_2564,In_628,In_619);
nand U2565 (N_2565,In_716,In_338);
and U2566 (N_2566,In_621,In_13);
or U2567 (N_2567,In_748,In_723);
or U2568 (N_2568,In_210,In_231);
nand U2569 (N_2569,In_789,In_102);
and U2570 (N_2570,In_800,In_964);
and U2571 (N_2571,In_246,In_700);
nor U2572 (N_2572,In_277,In_296);
nor U2573 (N_2573,In_321,In_21);
nor U2574 (N_2574,In_658,In_173);
or U2575 (N_2575,In_857,In_633);
nand U2576 (N_2576,In_138,In_840);
or U2577 (N_2577,In_443,In_498);
nor U2578 (N_2578,In_683,In_783);
nand U2579 (N_2579,In_404,In_38);
and U2580 (N_2580,In_909,In_398);
or U2581 (N_2581,In_899,In_758);
nor U2582 (N_2582,In_644,In_457);
and U2583 (N_2583,In_396,In_972);
nor U2584 (N_2584,In_776,In_232);
or U2585 (N_2585,In_645,In_637);
or U2586 (N_2586,In_608,In_317);
and U2587 (N_2587,In_15,In_444);
or U2588 (N_2588,In_909,In_165);
or U2589 (N_2589,In_260,In_569);
nor U2590 (N_2590,In_38,In_477);
and U2591 (N_2591,In_879,In_705);
nand U2592 (N_2592,In_520,In_976);
nand U2593 (N_2593,In_388,In_394);
or U2594 (N_2594,In_401,In_807);
nor U2595 (N_2595,In_797,In_9);
nand U2596 (N_2596,In_630,In_362);
or U2597 (N_2597,In_6,In_125);
or U2598 (N_2598,In_792,In_208);
and U2599 (N_2599,In_532,In_783);
nor U2600 (N_2600,In_878,In_767);
xor U2601 (N_2601,In_892,In_712);
and U2602 (N_2602,In_995,In_661);
and U2603 (N_2603,In_654,In_421);
nand U2604 (N_2604,In_910,In_229);
or U2605 (N_2605,In_62,In_97);
nand U2606 (N_2606,In_902,In_504);
and U2607 (N_2607,In_746,In_257);
nor U2608 (N_2608,In_326,In_318);
nand U2609 (N_2609,In_24,In_912);
or U2610 (N_2610,In_487,In_1);
or U2611 (N_2611,In_307,In_496);
nor U2612 (N_2612,In_727,In_98);
or U2613 (N_2613,In_678,In_475);
and U2614 (N_2614,In_853,In_523);
nand U2615 (N_2615,In_236,In_329);
or U2616 (N_2616,In_427,In_803);
nor U2617 (N_2617,In_307,In_938);
nand U2618 (N_2618,In_447,In_431);
and U2619 (N_2619,In_582,In_968);
and U2620 (N_2620,In_665,In_566);
nand U2621 (N_2621,In_579,In_657);
nand U2622 (N_2622,In_262,In_623);
or U2623 (N_2623,In_35,In_852);
nor U2624 (N_2624,In_77,In_646);
and U2625 (N_2625,In_916,In_390);
and U2626 (N_2626,In_585,In_405);
nand U2627 (N_2627,In_324,In_455);
nand U2628 (N_2628,In_202,In_301);
nand U2629 (N_2629,In_188,In_371);
nand U2630 (N_2630,In_911,In_785);
nor U2631 (N_2631,In_542,In_533);
nor U2632 (N_2632,In_724,In_246);
and U2633 (N_2633,In_299,In_83);
nand U2634 (N_2634,In_288,In_832);
and U2635 (N_2635,In_965,In_70);
nand U2636 (N_2636,In_827,In_249);
nor U2637 (N_2637,In_868,In_70);
nand U2638 (N_2638,In_581,In_555);
nor U2639 (N_2639,In_862,In_412);
or U2640 (N_2640,In_422,In_625);
or U2641 (N_2641,In_332,In_846);
or U2642 (N_2642,In_88,In_692);
and U2643 (N_2643,In_546,In_945);
and U2644 (N_2644,In_326,In_422);
nor U2645 (N_2645,In_27,In_3);
nand U2646 (N_2646,In_72,In_429);
nor U2647 (N_2647,In_990,In_928);
or U2648 (N_2648,In_878,In_674);
nor U2649 (N_2649,In_632,In_833);
and U2650 (N_2650,In_700,In_972);
nand U2651 (N_2651,In_983,In_739);
or U2652 (N_2652,In_315,In_428);
nand U2653 (N_2653,In_9,In_630);
and U2654 (N_2654,In_439,In_468);
or U2655 (N_2655,In_151,In_549);
xor U2656 (N_2656,In_565,In_797);
nor U2657 (N_2657,In_205,In_242);
or U2658 (N_2658,In_451,In_937);
or U2659 (N_2659,In_895,In_221);
nand U2660 (N_2660,In_20,In_331);
and U2661 (N_2661,In_560,In_471);
nor U2662 (N_2662,In_296,In_744);
and U2663 (N_2663,In_402,In_334);
or U2664 (N_2664,In_193,In_26);
or U2665 (N_2665,In_805,In_382);
or U2666 (N_2666,In_637,In_676);
nand U2667 (N_2667,In_711,In_484);
nand U2668 (N_2668,In_513,In_914);
nor U2669 (N_2669,In_142,In_956);
and U2670 (N_2670,In_744,In_947);
nand U2671 (N_2671,In_707,In_291);
and U2672 (N_2672,In_198,In_784);
nand U2673 (N_2673,In_603,In_492);
and U2674 (N_2674,In_529,In_763);
nand U2675 (N_2675,In_529,In_38);
and U2676 (N_2676,In_270,In_121);
nand U2677 (N_2677,In_800,In_514);
nor U2678 (N_2678,In_2,In_297);
or U2679 (N_2679,In_656,In_742);
and U2680 (N_2680,In_320,In_149);
and U2681 (N_2681,In_36,In_739);
nor U2682 (N_2682,In_843,In_310);
nand U2683 (N_2683,In_478,In_385);
or U2684 (N_2684,In_819,In_73);
or U2685 (N_2685,In_206,In_980);
nand U2686 (N_2686,In_869,In_937);
nand U2687 (N_2687,In_44,In_494);
nand U2688 (N_2688,In_412,In_795);
nand U2689 (N_2689,In_946,In_33);
nand U2690 (N_2690,In_912,In_331);
and U2691 (N_2691,In_592,In_113);
and U2692 (N_2692,In_717,In_58);
or U2693 (N_2693,In_878,In_827);
nand U2694 (N_2694,In_418,In_7);
nand U2695 (N_2695,In_104,In_454);
nor U2696 (N_2696,In_536,In_354);
or U2697 (N_2697,In_963,In_83);
nor U2698 (N_2698,In_626,In_424);
xor U2699 (N_2699,In_709,In_225);
nand U2700 (N_2700,In_933,In_636);
or U2701 (N_2701,In_96,In_882);
or U2702 (N_2702,In_963,In_713);
nand U2703 (N_2703,In_343,In_418);
or U2704 (N_2704,In_827,In_543);
nand U2705 (N_2705,In_445,In_261);
and U2706 (N_2706,In_14,In_186);
xor U2707 (N_2707,In_182,In_510);
or U2708 (N_2708,In_686,In_109);
and U2709 (N_2709,In_678,In_533);
and U2710 (N_2710,In_814,In_572);
and U2711 (N_2711,In_201,In_835);
and U2712 (N_2712,In_477,In_361);
nor U2713 (N_2713,In_179,In_425);
nand U2714 (N_2714,In_47,In_855);
nor U2715 (N_2715,In_208,In_101);
or U2716 (N_2716,In_882,In_543);
or U2717 (N_2717,In_94,In_468);
nand U2718 (N_2718,In_327,In_216);
and U2719 (N_2719,In_36,In_554);
nand U2720 (N_2720,In_886,In_769);
nor U2721 (N_2721,In_818,In_860);
and U2722 (N_2722,In_314,In_320);
and U2723 (N_2723,In_261,In_881);
nand U2724 (N_2724,In_265,In_794);
or U2725 (N_2725,In_506,In_182);
nor U2726 (N_2726,In_773,In_900);
nor U2727 (N_2727,In_67,In_791);
or U2728 (N_2728,In_809,In_818);
nor U2729 (N_2729,In_930,In_172);
or U2730 (N_2730,In_961,In_411);
nand U2731 (N_2731,In_621,In_477);
and U2732 (N_2732,In_911,In_959);
nor U2733 (N_2733,In_877,In_936);
and U2734 (N_2734,In_147,In_607);
or U2735 (N_2735,In_477,In_881);
and U2736 (N_2736,In_301,In_320);
or U2737 (N_2737,In_479,In_916);
and U2738 (N_2738,In_124,In_296);
nor U2739 (N_2739,In_400,In_163);
nand U2740 (N_2740,In_84,In_742);
or U2741 (N_2741,In_149,In_745);
or U2742 (N_2742,In_655,In_400);
nor U2743 (N_2743,In_212,In_989);
and U2744 (N_2744,In_835,In_444);
or U2745 (N_2745,In_390,In_856);
nand U2746 (N_2746,In_762,In_913);
or U2747 (N_2747,In_362,In_882);
nand U2748 (N_2748,In_323,In_615);
nor U2749 (N_2749,In_801,In_122);
or U2750 (N_2750,In_889,In_484);
nand U2751 (N_2751,In_200,In_28);
or U2752 (N_2752,In_811,In_946);
and U2753 (N_2753,In_498,In_117);
nand U2754 (N_2754,In_328,In_89);
nand U2755 (N_2755,In_196,In_884);
or U2756 (N_2756,In_666,In_545);
nor U2757 (N_2757,In_345,In_47);
nor U2758 (N_2758,In_635,In_617);
nand U2759 (N_2759,In_663,In_931);
nand U2760 (N_2760,In_329,In_437);
nand U2761 (N_2761,In_757,In_4);
and U2762 (N_2762,In_958,In_165);
nor U2763 (N_2763,In_722,In_529);
and U2764 (N_2764,In_446,In_619);
nand U2765 (N_2765,In_393,In_582);
nand U2766 (N_2766,In_823,In_817);
or U2767 (N_2767,In_923,In_137);
nor U2768 (N_2768,In_706,In_261);
nand U2769 (N_2769,In_824,In_373);
nand U2770 (N_2770,In_828,In_58);
and U2771 (N_2771,In_676,In_863);
or U2772 (N_2772,In_684,In_351);
and U2773 (N_2773,In_644,In_246);
xor U2774 (N_2774,In_860,In_8);
nand U2775 (N_2775,In_666,In_370);
nand U2776 (N_2776,In_334,In_255);
or U2777 (N_2777,In_815,In_145);
nand U2778 (N_2778,In_849,In_382);
nand U2779 (N_2779,In_220,In_576);
and U2780 (N_2780,In_325,In_363);
or U2781 (N_2781,In_124,In_919);
or U2782 (N_2782,In_629,In_24);
nor U2783 (N_2783,In_73,In_609);
and U2784 (N_2784,In_272,In_419);
or U2785 (N_2785,In_984,In_603);
nor U2786 (N_2786,In_104,In_958);
nand U2787 (N_2787,In_500,In_898);
and U2788 (N_2788,In_585,In_472);
or U2789 (N_2789,In_699,In_297);
nor U2790 (N_2790,In_337,In_622);
nand U2791 (N_2791,In_965,In_196);
or U2792 (N_2792,In_149,In_592);
nor U2793 (N_2793,In_814,In_906);
and U2794 (N_2794,In_523,In_516);
nor U2795 (N_2795,In_597,In_297);
nor U2796 (N_2796,In_745,In_215);
nor U2797 (N_2797,In_327,In_518);
nor U2798 (N_2798,In_618,In_468);
nor U2799 (N_2799,In_58,In_722);
nor U2800 (N_2800,In_210,In_118);
or U2801 (N_2801,In_386,In_167);
nor U2802 (N_2802,In_116,In_847);
and U2803 (N_2803,In_21,In_695);
nand U2804 (N_2804,In_857,In_273);
or U2805 (N_2805,In_122,In_365);
or U2806 (N_2806,In_911,In_760);
nand U2807 (N_2807,In_171,In_920);
or U2808 (N_2808,In_646,In_651);
nand U2809 (N_2809,In_441,In_978);
nand U2810 (N_2810,In_460,In_580);
nor U2811 (N_2811,In_197,In_587);
nor U2812 (N_2812,In_504,In_571);
and U2813 (N_2813,In_76,In_564);
nor U2814 (N_2814,In_860,In_332);
nand U2815 (N_2815,In_457,In_40);
or U2816 (N_2816,In_926,In_126);
nand U2817 (N_2817,In_114,In_760);
or U2818 (N_2818,In_692,In_39);
or U2819 (N_2819,In_816,In_690);
nand U2820 (N_2820,In_75,In_4);
or U2821 (N_2821,In_172,In_160);
nor U2822 (N_2822,In_129,In_153);
xnor U2823 (N_2823,In_33,In_597);
or U2824 (N_2824,In_927,In_675);
and U2825 (N_2825,In_311,In_837);
nor U2826 (N_2826,In_533,In_947);
or U2827 (N_2827,In_613,In_813);
and U2828 (N_2828,In_35,In_103);
or U2829 (N_2829,In_64,In_893);
or U2830 (N_2830,In_675,In_933);
nor U2831 (N_2831,In_593,In_552);
or U2832 (N_2832,In_386,In_501);
and U2833 (N_2833,In_146,In_480);
and U2834 (N_2834,In_429,In_345);
or U2835 (N_2835,In_408,In_610);
and U2836 (N_2836,In_975,In_957);
nor U2837 (N_2837,In_887,In_0);
or U2838 (N_2838,In_386,In_922);
and U2839 (N_2839,In_542,In_111);
nand U2840 (N_2840,In_224,In_287);
and U2841 (N_2841,In_561,In_888);
nor U2842 (N_2842,In_945,In_402);
and U2843 (N_2843,In_410,In_880);
and U2844 (N_2844,In_895,In_343);
nand U2845 (N_2845,In_725,In_303);
nor U2846 (N_2846,In_689,In_425);
nand U2847 (N_2847,In_991,In_666);
or U2848 (N_2848,In_538,In_100);
and U2849 (N_2849,In_335,In_569);
nand U2850 (N_2850,In_184,In_110);
nand U2851 (N_2851,In_64,In_563);
nor U2852 (N_2852,In_211,In_725);
nand U2853 (N_2853,In_553,In_594);
nor U2854 (N_2854,In_539,In_769);
nor U2855 (N_2855,In_800,In_273);
nor U2856 (N_2856,In_47,In_144);
nand U2857 (N_2857,In_370,In_777);
and U2858 (N_2858,In_667,In_297);
nand U2859 (N_2859,In_526,In_909);
nand U2860 (N_2860,In_996,In_399);
nand U2861 (N_2861,In_328,In_676);
or U2862 (N_2862,In_574,In_263);
nor U2863 (N_2863,In_639,In_735);
and U2864 (N_2864,In_29,In_253);
and U2865 (N_2865,In_817,In_384);
or U2866 (N_2866,In_517,In_754);
or U2867 (N_2867,In_135,In_842);
nand U2868 (N_2868,In_744,In_246);
or U2869 (N_2869,In_226,In_860);
nand U2870 (N_2870,In_366,In_43);
nor U2871 (N_2871,In_885,In_957);
or U2872 (N_2872,In_190,In_285);
and U2873 (N_2873,In_296,In_120);
nor U2874 (N_2874,In_678,In_843);
nand U2875 (N_2875,In_633,In_766);
nand U2876 (N_2876,In_215,In_35);
or U2877 (N_2877,In_938,In_949);
nand U2878 (N_2878,In_729,In_988);
nor U2879 (N_2879,In_247,In_309);
and U2880 (N_2880,In_867,In_249);
nand U2881 (N_2881,In_481,In_919);
and U2882 (N_2882,In_989,In_695);
nor U2883 (N_2883,In_307,In_536);
nand U2884 (N_2884,In_14,In_924);
nor U2885 (N_2885,In_701,In_349);
xor U2886 (N_2886,In_97,In_520);
and U2887 (N_2887,In_37,In_20);
nand U2888 (N_2888,In_563,In_596);
nand U2889 (N_2889,In_545,In_55);
nor U2890 (N_2890,In_246,In_542);
and U2891 (N_2891,In_445,In_837);
and U2892 (N_2892,In_792,In_470);
and U2893 (N_2893,In_515,In_861);
or U2894 (N_2894,In_377,In_47);
nand U2895 (N_2895,In_447,In_256);
and U2896 (N_2896,In_852,In_572);
nand U2897 (N_2897,In_264,In_935);
or U2898 (N_2898,In_64,In_413);
and U2899 (N_2899,In_507,In_771);
and U2900 (N_2900,In_269,In_57);
nand U2901 (N_2901,In_864,In_676);
nand U2902 (N_2902,In_542,In_233);
and U2903 (N_2903,In_555,In_565);
and U2904 (N_2904,In_901,In_79);
nor U2905 (N_2905,In_809,In_949);
and U2906 (N_2906,In_109,In_336);
nor U2907 (N_2907,In_494,In_841);
or U2908 (N_2908,In_486,In_910);
nor U2909 (N_2909,In_223,In_487);
nor U2910 (N_2910,In_731,In_295);
or U2911 (N_2911,In_326,In_407);
nand U2912 (N_2912,In_583,In_217);
or U2913 (N_2913,In_169,In_360);
or U2914 (N_2914,In_652,In_235);
nor U2915 (N_2915,In_358,In_397);
and U2916 (N_2916,In_819,In_280);
and U2917 (N_2917,In_961,In_550);
nor U2918 (N_2918,In_440,In_193);
or U2919 (N_2919,In_464,In_320);
nand U2920 (N_2920,In_677,In_587);
nor U2921 (N_2921,In_578,In_763);
nand U2922 (N_2922,In_406,In_397);
nand U2923 (N_2923,In_448,In_460);
nand U2924 (N_2924,In_129,In_23);
and U2925 (N_2925,In_23,In_848);
nor U2926 (N_2926,In_317,In_289);
or U2927 (N_2927,In_822,In_384);
nor U2928 (N_2928,In_930,In_680);
nor U2929 (N_2929,In_350,In_509);
and U2930 (N_2930,In_474,In_147);
and U2931 (N_2931,In_12,In_77);
nand U2932 (N_2932,In_154,In_503);
nand U2933 (N_2933,In_905,In_945);
nor U2934 (N_2934,In_158,In_895);
and U2935 (N_2935,In_938,In_907);
or U2936 (N_2936,In_493,In_696);
nand U2937 (N_2937,In_831,In_36);
or U2938 (N_2938,In_756,In_718);
or U2939 (N_2939,In_656,In_411);
nand U2940 (N_2940,In_314,In_85);
nor U2941 (N_2941,In_973,In_416);
and U2942 (N_2942,In_678,In_61);
or U2943 (N_2943,In_503,In_287);
and U2944 (N_2944,In_381,In_313);
nor U2945 (N_2945,In_916,In_796);
nand U2946 (N_2946,In_191,In_404);
or U2947 (N_2947,In_757,In_528);
nand U2948 (N_2948,In_263,In_102);
and U2949 (N_2949,In_238,In_81);
nor U2950 (N_2950,In_393,In_25);
nor U2951 (N_2951,In_945,In_915);
nor U2952 (N_2952,In_38,In_833);
nor U2953 (N_2953,In_130,In_97);
nand U2954 (N_2954,In_416,In_379);
or U2955 (N_2955,In_349,In_433);
nand U2956 (N_2956,In_463,In_438);
nand U2957 (N_2957,In_59,In_503);
nor U2958 (N_2958,In_986,In_605);
and U2959 (N_2959,In_565,In_27);
nand U2960 (N_2960,In_212,In_56);
nand U2961 (N_2961,In_532,In_784);
nor U2962 (N_2962,In_24,In_142);
or U2963 (N_2963,In_669,In_732);
and U2964 (N_2964,In_718,In_702);
nand U2965 (N_2965,In_955,In_41);
or U2966 (N_2966,In_959,In_396);
nand U2967 (N_2967,In_158,In_509);
and U2968 (N_2968,In_465,In_345);
or U2969 (N_2969,In_51,In_882);
or U2970 (N_2970,In_887,In_386);
nor U2971 (N_2971,In_262,In_761);
nor U2972 (N_2972,In_724,In_198);
nor U2973 (N_2973,In_358,In_859);
nor U2974 (N_2974,In_847,In_759);
nand U2975 (N_2975,In_442,In_487);
or U2976 (N_2976,In_242,In_14);
nand U2977 (N_2977,In_522,In_50);
nor U2978 (N_2978,In_476,In_0);
nand U2979 (N_2979,In_137,In_986);
or U2980 (N_2980,In_787,In_529);
nor U2981 (N_2981,In_413,In_806);
and U2982 (N_2982,In_7,In_644);
or U2983 (N_2983,In_927,In_328);
and U2984 (N_2984,In_883,In_834);
nand U2985 (N_2985,In_640,In_506);
nand U2986 (N_2986,In_572,In_591);
or U2987 (N_2987,In_192,In_348);
or U2988 (N_2988,In_463,In_303);
nor U2989 (N_2989,In_449,In_488);
and U2990 (N_2990,In_154,In_857);
nor U2991 (N_2991,In_812,In_137);
nand U2992 (N_2992,In_28,In_232);
nor U2993 (N_2993,In_657,In_126);
or U2994 (N_2994,In_521,In_587);
or U2995 (N_2995,In_67,In_810);
or U2996 (N_2996,In_834,In_14);
and U2997 (N_2997,In_382,In_557);
or U2998 (N_2998,In_108,In_854);
nand U2999 (N_2999,In_396,In_725);
or U3000 (N_3000,In_459,In_228);
or U3001 (N_3001,In_461,In_503);
nand U3002 (N_3002,In_919,In_525);
or U3003 (N_3003,In_696,In_606);
or U3004 (N_3004,In_909,In_966);
and U3005 (N_3005,In_108,In_66);
and U3006 (N_3006,In_133,In_815);
nand U3007 (N_3007,In_742,In_671);
nor U3008 (N_3008,In_979,In_515);
nor U3009 (N_3009,In_268,In_654);
and U3010 (N_3010,In_716,In_735);
nand U3011 (N_3011,In_615,In_661);
nand U3012 (N_3012,In_984,In_271);
or U3013 (N_3013,In_330,In_135);
or U3014 (N_3014,In_126,In_217);
nor U3015 (N_3015,In_424,In_874);
and U3016 (N_3016,In_711,In_435);
nand U3017 (N_3017,In_641,In_77);
nor U3018 (N_3018,In_361,In_84);
and U3019 (N_3019,In_493,In_183);
and U3020 (N_3020,In_699,In_960);
and U3021 (N_3021,In_616,In_852);
nand U3022 (N_3022,In_176,In_815);
or U3023 (N_3023,In_222,In_687);
and U3024 (N_3024,In_629,In_682);
nor U3025 (N_3025,In_821,In_323);
and U3026 (N_3026,In_158,In_362);
and U3027 (N_3027,In_498,In_260);
and U3028 (N_3028,In_579,In_8);
nand U3029 (N_3029,In_4,In_81);
and U3030 (N_3030,In_659,In_821);
and U3031 (N_3031,In_648,In_806);
nand U3032 (N_3032,In_319,In_446);
nand U3033 (N_3033,In_392,In_898);
nor U3034 (N_3034,In_944,In_682);
or U3035 (N_3035,In_545,In_864);
or U3036 (N_3036,In_87,In_737);
or U3037 (N_3037,In_304,In_455);
nor U3038 (N_3038,In_635,In_757);
and U3039 (N_3039,In_161,In_378);
or U3040 (N_3040,In_694,In_285);
or U3041 (N_3041,In_526,In_701);
and U3042 (N_3042,In_976,In_298);
and U3043 (N_3043,In_139,In_272);
and U3044 (N_3044,In_160,In_736);
or U3045 (N_3045,In_901,In_432);
and U3046 (N_3046,In_975,In_447);
nor U3047 (N_3047,In_136,In_144);
nor U3048 (N_3048,In_132,In_590);
or U3049 (N_3049,In_425,In_925);
or U3050 (N_3050,In_834,In_375);
or U3051 (N_3051,In_347,In_892);
nor U3052 (N_3052,In_808,In_620);
nand U3053 (N_3053,In_715,In_93);
nor U3054 (N_3054,In_376,In_162);
or U3055 (N_3055,In_217,In_133);
and U3056 (N_3056,In_154,In_52);
nor U3057 (N_3057,In_728,In_424);
nor U3058 (N_3058,In_144,In_763);
nor U3059 (N_3059,In_291,In_132);
nor U3060 (N_3060,In_928,In_683);
and U3061 (N_3061,In_259,In_799);
nand U3062 (N_3062,In_531,In_284);
and U3063 (N_3063,In_538,In_914);
or U3064 (N_3064,In_413,In_525);
and U3065 (N_3065,In_576,In_934);
and U3066 (N_3066,In_236,In_383);
or U3067 (N_3067,In_422,In_670);
nor U3068 (N_3068,In_779,In_83);
nand U3069 (N_3069,In_725,In_434);
nor U3070 (N_3070,In_970,In_574);
nand U3071 (N_3071,In_888,In_625);
or U3072 (N_3072,In_510,In_469);
nand U3073 (N_3073,In_691,In_523);
and U3074 (N_3074,In_519,In_296);
nor U3075 (N_3075,In_449,In_563);
and U3076 (N_3076,In_124,In_666);
and U3077 (N_3077,In_208,In_653);
nand U3078 (N_3078,In_564,In_963);
nand U3079 (N_3079,In_278,In_66);
and U3080 (N_3080,In_674,In_58);
and U3081 (N_3081,In_704,In_346);
nor U3082 (N_3082,In_278,In_32);
and U3083 (N_3083,In_477,In_596);
nor U3084 (N_3084,In_847,In_504);
nor U3085 (N_3085,In_75,In_119);
nand U3086 (N_3086,In_439,In_610);
nand U3087 (N_3087,In_212,In_600);
and U3088 (N_3088,In_406,In_658);
and U3089 (N_3089,In_206,In_853);
nand U3090 (N_3090,In_184,In_505);
nand U3091 (N_3091,In_405,In_283);
and U3092 (N_3092,In_75,In_645);
nor U3093 (N_3093,In_555,In_423);
and U3094 (N_3094,In_368,In_660);
xnor U3095 (N_3095,In_726,In_75);
nor U3096 (N_3096,In_272,In_363);
and U3097 (N_3097,In_836,In_11);
xor U3098 (N_3098,In_996,In_477);
and U3099 (N_3099,In_504,In_838);
or U3100 (N_3100,In_690,In_806);
nand U3101 (N_3101,In_582,In_822);
and U3102 (N_3102,In_201,In_356);
nor U3103 (N_3103,In_868,In_873);
nor U3104 (N_3104,In_286,In_470);
or U3105 (N_3105,In_901,In_593);
and U3106 (N_3106,In_48,In_170);
or U3107 (N_3107,In_877,In_431);
nand U3108 (N_3108,In_754,In_354);
or U3109 (N_3109,In_514,In_21);
nor U3110 (N_3110,In_294,In_732);
and U3111 (N_3111,In_345,In_973);
nor U3112 (N_3112,In_527,In_392);
nand U3113 (N_3113,In_528,In_145);
and U3114 (N_3114,In_546,In_802);
and U3115 (N_3115,In_124,In_82);
and U3116 (N_3116,In_532,In_37);
nor U3117 (N_3117,In_14,In_342);
nor U3118 (N_3118,In_508,In_161);
nor U3119 (N_3119,In_470,In_871);
nor U3120 (N_3120,In_568,In_899);
nand U3121 (N_3121,In_124,In_275);
and U3122 (N_3122,In_158,In_821);
nor U3123 (N_3123,In_999,In_384);
nor U3124 (N_3124,In_469,In_593);
or U3125 (N_3125,In_823,In_547);
nor U3126 (N_3126,In_705,In_697);
and U3127 (N_3127,In_914,In_756);
or U3128 (N_3128,In_268,In_533);
and U3129 (N_3129,In_269,In_85);
or U3130 (N_3130,In_403,In_441);
nand U3131 (N_3131,In_558,In_411);
nor U3132 (N_3132,In_636,In_835);
or U3133 (N_3133,In_179,In_883);
and U3134 (N_3134,In_3,In_571);
nor U3135 (N_3135,In_137,In_365);
nor U3136 (N_3136,In_483,In_236);
nand U3137 (N_3137,In_387,In_874);
nand U3138 (N_3138,In_973,In_409);
nand U3139 (N_3139,In_577,In_200);
or U3140 (N_3140,In_51,In_223);
or U3141 (N_3141,In_329,In_380);
xor U3142 (N_3142,In_105,In_952);
nand U3143 (N_3143,In_461,In_884);
nor U3144 (N_3144,In_144,In_831);
nand U3145 (N_3145,In_995,In_486);
and U3146 (N_3146,In_561,In_0);
nand U3147 (N_3147,In_762,In_331);
xnor U3148 (N_3148,In_687,In_666);
or U3149 (N_3149,In_383,In_853);
xnor U3150 (N_3150,In_958,In_594);
nor U3151 (N_3151,In_885,In_330);
and U3152 (N_3152,In_878,In_341);
or U3153 (N_3153,In_170,In_853);
or U3154 (N_3154,In_311,In_109);
and U3155 (N_3155,In_683,In_506);
or U3156 (N_3156,In_693,In_726);
and U3157 (N_3157,In_323,In_641);
and U3158 (N_3158,In_916,In_651);
nand U3159 (N_3159,In_705,In_749);
nor U3160 (N_3160,In_784,In_870);
nand U3161 (N_3161,In_943,In_392);
and U3162 (N_3162,In_150,In_405);
nand U3163 (N_3163,In_578,In_680);
and U3164 (N_3164,In_845,In_291);
or U3165 (N_3165,In_998,In_942);
and U3166 (N_3166,In_2,In_704);
or U3167 (N_3167,In_868,In_931);
and U3168 (N_3168,In_601,In_545);
nand U3169 (N_3169,In_525,In_173);
nor U3170 (N_3170,In_25,In_739);
and U3171 (N_3171,In_303,In_678);
or U3172 (N_3172,In_689,In_222);
or U3173 (N_3173,In_381,In_468);
nand U3174 (N_3174,In_62,In_731);
and U3175 (N_3175,In_939,In_800);
nand U3176 (N_3176,In_343,In_718);
nor U3177 (N_3177,In_106,In_565);
and U3178 (N_3178,In_913,In_886);
and U3179 (N_3179,In_355,In_112);
or U3180 (N_3180,In_864,In_803);
and U3181 (N_3181,In_225,In_730);
or U3182 (N_3182,In_675,In_474);
nand U3183 (N_3183,In_384,In_701);
or U3184 (N_3184,In_234,In_639);
or U3185 (N_3185,In_784,In_882);
or U3186 (N_3186,In_925,In_10);
and U3187 (N_3187,In_112,In_862);
or U3188 (N_3188,In_456,In_981);
nor U3189 (N_3189,In_793,In_353);
nor U3190 (N_3190,In_56,In_314);
and U3191 (N_3191,In_561,In_416);
or U3192 (N_3192,In_852,In_246);
and U3193 (N_3193,In_756,In_436);
or U3194 (N_3194,In_181,In_95);
or U3195 (N_3195,In_985,In_446);
and U3196 (N_3196,In_598,In_711);
nand U3197 (N_3197,In_173,In_51);
nand U3198 (N_3198,In_248,In_93);
nand U3199 (N_3199,In_150,In_900);
nor U3200 (N_3200,In_885,In_633);
and U3201 (N_3201,In_33,In_6);
or U3202 (N_3202,In_61,In_768);
or U3203 (N_3203,In_171,In_167);
nor U3204 (N_3204,In_364,In_934);
and U3205 (N_3205,In_29,In_37);
and U3206 (N_3206,In_74,In_752);
nand U3207 (N_3207,In_502,In_762);
nor U3208 (N_3208,In_278,In_458);
nand U3209 (N_3209,In_282,In_706);
nand U3210 (N_3210,In_877,In_602);
or U3211 (N_3211,In_783,In_218);
nor U3212 (N_3212,In_903,In_61);
nand U3213 (N_3213,In_18,In_30);
or U3214 (N_3214,In_107,In_999);
or U3215 (N_3215,In_877,In_623);
nand U3216 (N_3216,In_415,In_380);
nor U3217 (N_3217,In_793,In_596);
or U3218 (N_3218,In_938,In_232);
nand U3219 (N_3219,In_189,In_595);
nor U3220 (N_3220,In_20,In_282);
or U3221 (N_3221,In_125,In_819);
nand U3222 (N_3222,In_840,In_42);
or U3223 (N_3223,In_702,In_216);
and U3224 (N_3224,In_906,In_380);
and U3225 (N_3225,In_151,In_187);
nor U3226 (N_3226,In_940,In_334);
or U3227 (N_3227,In_708,In_722);
nand U3228 (N_3228,In_169,In_518);
and U3229 (N_3229,In_171,In_80);
nor U3230 (N_3230,In_424,In_535);
nor U3231 (N_3231,In_658,In_43);
or U3232 (N_3232,In_386,In_738);
or U3233 (N_3233,In_746,In_628);
xnor U3234 (N_3234,In_247,In_134);
and U3235 (N_3235,In_853,In_681);
nand U3236 (N_3236,In_792,In_935);
nand U3237 (N_3237,In_855,In_275);
and U3238 (N_3238,In_862,In_133);
or U3239 (N_3239,In_90,In_543);
or U3240 (N_3240,In_638,In_167);
nor U3241 (N_3241,In_522,In_615);
nand U3242 (N_3242,In_339,In_218);
nor U3243 (N_3243,In_987,In_626);
nor U3244 (N_3244,In_38,In_206);
nand U3245 (N_3245,In_850,In_913);
and U3246 (N_3246,In_498,In_566);
nor U3247 (N_3247,In_608,In_544);
nand U3248 (N_3248,In_10,In_75);
or U3249 (N_3249,In_372,In_901);
nor U3250 (N_3250,In_738,In_76);
nor U3251 (N_3251,In_364,In_806);
or U3252 (N_3252,In_308,In_849);
nor U3253 (N_3253,In_214,In_913);
nor U3254 (N_3254,In_207,In_908);
or U3255 (N_3255,In_783,In_422);
nor U3256 (N_3256,In_932,In_860);
nor U3257 (N_3257,In_151,In_304);
nor U3258 (N_3258,In_642,In_56);
and U3259 (N_3259,In_560,In_13);
nor U3260 (N_3260,In_502,In_329);
nand U3261 (N_3261,In_782,In_82);
nand U3262 (N_3262,In_754,In_353);
nand U3263 (N_3263,In_968,In_749);
nand U3264 (N_3264,In_495,In_985);
or U3265 (N_3265,In_158,In_465);
or U3266 (N_3266,In_959,In_385);
nor U3267 (N_3267,In_201,In_680);
nor U3268 (N_3268,In_53,In_963);
or U3269 (N_3269,In_182,In_117);
nor U3270 (N_3270,In_90,In_292);
or U3271 (N_3271,In_653,In_330);
nand U3272 (N_3272,In_410,In_763);
nor U3273 (N_3273,In_257,In_457);
nand U3274 (N_3274,In_794,In_275);
and U3275 (N_3275,In_739,In_361);
nor U3276 (N_3276,In_26,In_809);
nor U3277 (N_3277,In_720,In_650);
nor U3278 (N_3278,In_272,In_812);
nand U3279 (N_3279,In_24,In_450);
nand U3280 (N_3280,In_691,In_679);
nand U3281 (N_3281,In_788,In_876);
nor U3282 (N_3282,In_6,In_405);
and U3283 (N_3283,In_555,In_346);
nor U3284 (N_3284,In_725,In_414);
nand U3285 (N_3285,In_355,In_198);
nand U3286 (N_3286,In_65,In_52);
nor U3287 (N_3287,In_357,In_456);
nand U3288 (N_3288,In_525,In_456);
nor U3289 (N_3289,In_425,In_326);
nand U3290 (N_3290,In_811,In_972);
or U3291 (N_3291,In_689,In_676);
or U3292 (N_3292,In_258,In_759);
or U3293 (N_3293,In_698,In_501);
and U3294 (N_3294,In_615,In_803);
and U3295 (N_3295,In_426,In_677);
or U3296 (N_3296,In_855,In_647);
nor U3297 (N_3297,In_592,In_424);
nor U3298 (N_3298,In_698,In_611);
or U3299 (N_3299,In_740,In_17);
or U3300 (N_3300,In_118,In_858);
xnor U3301 (N_3301,In_729,In_547);
nor U3302 (N_3302,In_105,In_246);
nor U3303 (N_3303,In_442,In_562);
or U3304 (N_3304,In_398,In_854);
nand U3305 (N_3305,In_3,In_41);
nand U3306 (N_3306,In_353,In_610);
and U3307 (N_3307,In_401,In_723);
nand U3308 (N_3308,In_93,In_553);
nor U3309 (N_3309,In_245,In_43);
nor U3310 (N_3310,In_803,In_277);
nor U3311 (N_3311,In_333,In_222);
and U3312 (N_3312,In_873,In_920);
nor U3313 (N_3313,In_681,In_270);
nand U3314 (N_3314,In_444,In_308);
or U3315 (N_3315,In_374,In_320);
and U3316 (N_3316,In_803,In_709);
or U3317 (N_3317,In_238,In_587);
nor U3318 (N_3318,In_575,In_221);
or U3319 (N_3319,In_540,In_780);
and U3320 (N_3320,In_151,In_136);
nand U3321 (N_3321,In_257,In_825);
or U3322 (N_3322,In_657,In_396);
and U3323 (N_3323,In_50,In_610);
nand U3324 (N_3324,In_234,In_328);
nand U3325 (N_3325,In_376,In_803);
nand U3326 (N_3326,In_387,In_155);
nor U3327 (N_3327,In_901,In_672);
or U3328 (N_3328,In_277,In_600);
and U3329 (N_3329,In_834,In_965);
and U3330 (N_3330,In_143,In_482);
and U3331 (N_3331,In_850,In_555);
nor U3332 (N_3332,In_879,In_384);
or U3333 (N_3333,In_802,In_828);
or U3334 (N_3334,In_321,In_572);
and U3335 (N_3335,In_841,In_367);
and U3336 (N_3336,In_225,In_569);
nor U3337 (N_3337,In_593,In_845);
and U3338 (N_3338,In_129,In_315);
nor U3339 (N_3339,In_279,In_36);
nand U3340 (N_3340,In_659,In_805);
nand U3341 (N_3341,In_19,In_667);
and U3342 (N_3342,In_962,In_394);
nor U3343 (N_3343,In_543,In_900);
nor U3344 (N_3344,In_55,In_773);
or U3345 (N_3345,In_286,In_481);
and U3346 (N_3346,In_596,In_229);
nand U3347 (N_3347,In_53,In_40);
nand U3348 (N_3348,In_649,In_934);
nand U3349 (N_3349,In_419,In_462);
and U3350 (N_3350,In_646,In_609);
and U3351 (N_3351,In_650,In_600);
and U3352 (N_3352,In_840,In_156);
nor U3353 (N_3353,In_21,In_578);
nor U3354 (N_3354,In_629,In_840);
nand U3355 (N_3355,In_721,In_218);
nand U3356 (N_3356,In_226,In_564);
or U3357 (N_3357,In_412,In_4);
nand U3358 (N_3358,In_738,In_592);
and U3359 (N_3359,In_461,In_33);
nor U3360 (N_3360,In_111,In_101);
nor U3361 (N_3361,In_253,In_161);
nand U3362 (N_3362,In_650,In_82);
nand U3363 (N_3363,In_47,In_615);
nand U3364 (N_3364,In_879,In_510);
nand U3365 (N_3365,In_340,In_448);
nand U3366 (N_3366,In_806,In_312);
and U3367 (N_3367,In_860,In_125);
nor U3368 (N_3368,In_321,In_37);
nor U3369 (N_3369,In_856,In_80);
nor U3370 (N_3370,In_417,In_724);
and U3371 (N_3371,In_995,In_184);
and U3372 (N_3372,In_255,In_195);
or U3373 (N_3373,In_53,In_799);
nand U3374 (N_3374,In_455,In_901);
and U3375 (N_3375,In_827,In_492);
nor U3376 (N_3376,In_598,In_284);
nor U3377 (N_3377,In_587,In_398);
nor U3378 (N_3378,In_436,In_973);
or U3379 (N_3379,In_977,In_738);
nor U3380 (N_3380,In_325,In_364);
nand U3381 (N_3381,In_368,In_859);
or U3382 (N_3382,In_562,In_726);
or U3383 (N_3383,In_6,In_381);
and U3384 (N_3384,In_116,In_866);
nand U3385 (N_3385,In_288,In_667);
or U3386 (N_3386,In_645,In_871);
nand U3387 (N_3387,In_60,In_203);
nor U3388 (N_3388,In_765,In_634);
nor U3389 (N_3389,In_564,In_14);
or U3390 (N_3390,In_503,In_975);
and U3391 (N_3391,In_690,In_862);
and U3392 (N_3392,In_160,In_737);
nor U3393 (N_3393,In_393,In_944);
or U3394 (N_3394,In_485,In_618);
nand U3395 (N_3395,In_873,In_999);
xnor U3396 (N_3396,In_927,In_683);
nand U3397 (N_3397,In_756,In_183);
or U3398 (N_3398,In_508,In_651);
xor U3399 (N_3399,In_628,In_260);
and U3400 (N_3400,In_117,In_37);
and U3401 (N_3401,In_117,In_731);
nand U3402 (N_3402,In_377,In_539);
nor U3403 (N_3403,In_720,In_10);
nand U3404 (N_3404,In_674,In_335);
nor U3405 (N_3405,In_284,In_630);
or U3406 (N_3406,In_417,In_459);
or U3407 (N_3407,In_93,In_723);
nand U3408 (N_3408,In_834,In_702);
or U3409 (N_3409,In_214,In_249);
nor U3410 (N_3410,In_643,In_524);
nor U3411 (N_3411,In_595,In_427);
nor U3412 (N_3412,In_579,In_687);
nor U3413 (N_3413,In_969,In_481);
nor U3414 (N_3414,In_366,In_360);
nand U3415 (N_3415,In_738,In_61);
and U3416 (N_3416,In_216,In_475);
and U3417 (N_3417,In_810,In_143);
or U3418 (N_3418,In_530,In_173);
nor U3419 (N_3419,In_961,In_420);
nand U3420 (N_3420,In_355,In_796);
nand U3421 (N_3421,In_688,In_17);
nor U3422 (N_3422,In_870,In_747);
nor U3423 (N_3423,In_729,In_982);
and U3424 (N_3424,In_164,In_530);
nor U3425 (N_3425,In_17,In_336);
nor U3426 (N_3426,In_531,In_749);
nor U3427 (N_3427,In_527,In_803);
and U3428 (N_3428,In_234,In_984);
and U3429 (N_3429,In_16,In_901);
or U3430 (N_3430,In_419,In_330);
nor U3431 (N_3431,In_627,In_118);
and U3432 (N_3432,In_289,In_600);
or U3433 (N_3433,In_643,In_851);
nor U3434 (N_3434,In_711,In_252);
nand U3435 (N_3435,In_428,In_638);
and U3436 (N_3436,In_112,In_31);
nor U3437 (N_3437,In_118,In_6);
nor U3438 (N_3438,In_961,In_49);
nand U3439 (N_3439,In_929,In_667);
nor U3440 (N_3440,In_673,In_935);
and U3441 (N_3441,In_961,In_814);
nor U3442 (N_3442,In_810,In_431);
and U3443 (N_3443,In_986,In_71);
and U3444 (N_3444,In_896,In_537);
nand U3445 (N_3445,In_698,In_126);
nor U3446 (N_3446,In_591,In_654);
nand U3447 (N_3447,In_936,In_504);
or U3448 (N_3448,In_261,In_136);
nand U3449 (N_3449,In_525,In_135);
nand U3450 (N_3450,In_901,In_387);
and U3451 (N_3451,In_621,In_324);
or U3452 (N_3452,In_30,In_112);
and U3453 (N_3453,In_301,In_520);
nor U3454 (N_3454,In_373,In_581);
nor U3455 (N_3455,In_149,In_459);
nand U3456 (N_3456,In_909,In_583);
and U3457 (N_3457,In_937,In_601);
nand U3458 (N_3458,In_789,In_898);
and U3459 (N_3459,In_624,In_672);
and U3460 (N_3460,In_566,In_579);
or U3461 (N_3461,In_224,In_916);
or U3462 (N_3462,In_467,In_145);
nand U3463 (N_3463,In_303,In_234);
and U3464 (N_3464,In_108,In_935);
and U3465 (N_3465,In_253,In_19);
nor U3466 (N_3466,In_967,In_578);
and U3467 (N_3467,In_136,In_902);
and U3468 (N_3468,In_267,In_277);
nand U3469 (N_3469,In_355,In_905);
nand U3470 (N_3470,In_424,In_853);
nor U3471 (N_3471,In_592,In_838);
nor U3472 (N_3472,In_437,In_127);
nand U3473 (N_3473,In_88,In_244);
nand U3474 (N_3474,In_815,In_385);
and U3475 (N_3475,In_715,In_494);
nor U3476 (N_3476,In_140,In_169);
and U3477 (N_3477,In_452,In_856);
and U3478 (N_3478,In_34,In_371);
nor U3479 (N_3479,In_218,In_375);
nand U3480 (N_3480,In_513,In_875);
nor U3481 (N_3481,In_248,In_121);
and U3482 (N_3482,In_146,In_570);
or U3483 (N_3483,In_226,In_904);
and U3484 (N_3484,In_774,In_712);
or U3485 (N_3485,In_258,In_839);
and U3486 (N_3486,In_929,In_127);
and U3487 (N_3487,In_280,In_460);
nor U3488 (N_3488,In_901,In_991);
or U3489 (N_3489,In_338,In_905);
and U3490 (N_3490,In_106,In_891);
or U3491 (N_3491,In_662,In_173);
nor U3492 (N_3492,In_599,In_423);
nor U3493 (N_3493,In_877,In_347);
or U3494 (N_3494,In_438,In_964);
nand U3495 (N_3495,In_594,In_122);
and U3496 (N_3496,In_52,In_42);
or U3497 (N_3497,In_763,In_844);
nand U3498 (N_3498,In_920,In_78);
nor U3499 (N_3499,In_993,In_776);
and U3500 (N_3500,In_728,In_115);
nand U3501 (N_3501,In_942,In_671);
and U3502 (N_3502,In_364,In_469);
or U3503 (N_3503,In_625,In_142);
or U3504 (N_3504,In_101,In_31);
xor U3505 (N_3505,In_662,In_918);
nand U3506 (N_3506,In_44,In_723);
nand U3507 (N_3507,In_827,In_406);
nand U3508 (N_3508,In_279,In_319);
or U3509 (N_3509,In_380,In_591);
nor U3510 (N_3510,In_807,In_399);
nor U3511 (N_3511,In_8,In_984);
or U3512 (N_3512,In_815,In_465);
nand U3513 (N_3513,In_81,In_599);
or U3514 (N_3514,In_479,In_149);
nand U3515 (N_3515,In_396,In_651);
nand U3516 (N_3516,In_381,In_791);
nand U3517 (N_3517,In_964,In_798);
and U3518 (N_3518,In_713,In_299);
nor U3519 (N_3519,In_847,In_945);
and U3520 (N_3520,In_530,In_806);
xnor U3521 (N_3521,In_691,In_276);
nor U3522 (N_3522,In_432,In_841);
or U3523 (N_3523,In_943,In_436);
nand U3524 (N_3524,In_366,In_424);
or U3525 (N_3525,In_899,In_266);
or U3526 (N_3526,In_323,In_92);
nor U3527 (N_3527,In_549,In_771);
and U3528 (N_3528,In_972,In_313);
or U3529 (N_3529,In_443,In_684);
and U3530 (N_3530,In_441,In_291);
nor U3531 (N_3531,In_606,In_788);
and U3532 (N_3532,In_424,In_350);
nand U3533 (N_3533,In_936,In_703);
nand U3534 (N_3534,In_350,In_644);
or U3535 (N_3535,In_156,In_628);
nand U3536 (N_3536,In_816,In_941);
nand U3537 (N_3537,In_919,In_570);
nor U3538 (N_3538,In_401,In_84);
nor U3539 (N_3539,In_641,In_797);
nand U3540 (N_3540,In_115,In_278);
xnor U3541 (N_3541,In_945,In_892);
nor U3542 (N_3542,In_200,In_129);
or U3543 (N_3543,In_644,In_840);
nor U3544 (N_3544,In_727,In_608);
nand U3545 (N_3545,In_90,In_495);
and U3546 (N_3546,In_853,In_977);
or U3547 (N_3547,In_381,In_4);
or U3548 (N_3548,In_356,In_403);
nor U3549 (N_3549,In_622,In_455);
nand U3550 (N_3550,In_706,In_757);
or U3551 (N_3551,In_760,In_339);
nand U3552 (N_3552,In_32,In_292);
nor U3553 (N_3553,In_656,In_78);
and U3554 (N_3554,In_212,In_430);
nor U3555 (N_3555,In_749,In_17);
and U3556 (N_3556,In_359,In_994);
xnor U3557 (N_3557,In_943,In_280);
nor U3558 (N_3558,In_598,In_331);
and U3559 (N_3559,In_579,In_806);
nor U3560 (N_3560,In_791,In_459);
or U3561 (N_3561,In_626,In_122);
nor U3562 (N_3562,In_755,In_449);
xor U3563 (N_3563,In_3,In_218);
or U3564 (N_3564,In_229,In_547);
or U3565 (N_3565,In_176,In_913);
nand U3566 (N_3566,In_255,In_320);
nor U3567 (N_3567,In_90,In_741);
or U3568 (N_3568,In_364,In_681);
or U3569 (N_3569,In_565,In_260);
nor U3570 (N_3570,In_290,In_916);
nand U3571 (N_3571,In_683,In_968);
nand U3572 (N_3572,In_2,In_891);
and U3573 (N_3573,In_894,In_25);
nand U3574 (N_3574,In_405,In_425);
nand U3575 (N_3575,In_168,In_995);
nor U3576 (N_3576,In_338,In_388);
or U3577 (N_3577,In_262,In_845);
or U3578 (N_3578,In_265,In_636);
nor U3579 (N_3579,In_371,In_715);
nand U3580 (N_3580,In_529,In_999);
nor U3581 (N_3581,In_759,In_265);
and U3582 (N_3582,In_59,In_713);
or U3583 (N_3583,In_755,In_38);
nor U3584 (N_3584,In_296,In_923);
nor U3585 (N_3585,In_565,In_507);
nor U3586 (N_3586,In_935,In_866);
nor U3587 (N_3587,In_530,In_250);
and U3588 (N_3588,In_741,In_393);
or U3589 (N_3589,In_801,In_941);
and U3590 (N_3590,In_893,In_707);
nand U3591 (N_3591,In_932,In_95);
nand U3592 (N_3592,In_928,In_459);
nand U3593 (N_3593,In_555,In_878);
and U3594 (N_3594,In_487,In_850);
and U3595 (N_3595,In_161,In_362);
and U3596 (N_3596,In_237,In_275);
nor U3597 (N_3597,In_910,In_21);
or U3598 (N_3598,In_453,In_146);
and U3599 (N_3599,In_22,In_740);
and U3600 (N_3600,In_913,In_442);
and U3601 (N_3601,In_324,In_425);
and U3602 (N_3602,In_546,In_575);
or U3603 (N_3603,In_767,In_433);
nor U3604 (N_3604,In_648,In_491);
xnor U3605 (N_3605,In_665,In_879);
nor U3606 (N_3606,In_503,In_459);
or U3607 (N_3607,In_699,In_430);
or U3608 (N_3608,In_648,In_990);
and U3609 (N_3609,In_76,In_242);
nand U3610 (N_3610,In_394,In_201);
and U3611 (N_3611,In_950,In_493);
or U3612 (N_3612,In_105,In_634);
or U3613 (N_3613,In_32,In_631);
or U3614 (N_3614,In_798,In_698);
and U3615 (N_3615,In_322,In_74);
nor U3616 (N_3616,In_908,In_195);
and U3617 (N_3617,In_749,In_335);
nor U3618 (N_3618,In_793,In_316);
nand U3619 (N_3619,In_558,In_614);
nor U3620 (N_3620,In_834,In_48);
nor U3621 (N_3621,In_288,In_364);
nand U3622 (N_3622,In_595,In_218);
and U3623 (N_3623,In_262,In_653);
nand U3624 (N_3624,In_580,In_488);
and U3625 (N_3625,In_49,In_757);
nor U3626 (N_3626,In_452,In_77);
nor U3627 (N_3627,In_4,In_745);
or U3628 (N_3628,In_543,In_366);
or U3629 (N_3629,In_150,In_157);
nor U3630 (N_3630,In_76,In_406);
nor U3631 (N_3631,In_291,In_619);
nor U3632 (N_3632,In_97,In_103);
or U3633 (N_3633,In_492,In_278);
xnor U3634 (N_3634,In_179,In_776);
nand U3635 (N_3635,In_175,In_598);
nor U3636 (N_3636,In_72,In_165);
nand U3637 (N_3637,In_944,In_584);
and U3638 (N_3638,In_760,In_508);
nand U3639 (N_3639,In_265,In_885);
nand U3640 (N_3640,In_833,In_286);
nand U3641 (N_3641,In_846,In_941);
nor U3642 (N_3642,In_37,In_163);
or U3643 (N_3643,In_829,In_803);
nor U3644 (N_3644,In_164,In_919);
nor U3645 (N_3645,In_45,In_842);
and U3646 (N_3646,In_805,In_333);
or U3647 (N_3647,In_180,In_732);
and U3648 (N_3648,In_852,In_39);
or U3649 (N_3649,In_192,In_798);
nor U3650 (N_3650,In_591,In_933);
or U3651 (N_3651,In_258,In_465);
nor U3652 (N_3652,In_636,In_486);
and U3653 (N_3653,In_919,In_39);
nor U3654 (N_3654,In_575,In_90);
or U3655 (N_3655,In_175,In_0);
and U3656 (N_3656,In_891,In_835);
and U3657 (N_3657,In_222,In_911);
nand U3658 (N_3658,In_290,In_663);
nand U3659 (N_3659,In_509,In_446);
nor U3660 (N_3660,In_649,In_61);
and U3661 (N_3661,In_64,In_863);
or U3662 (N_3662,In_22,In_7);
nor U3663 (N_3663,In_129,In_994);
nor U3664 (N_3664,In_622,In_378);
and U3665 (N_3665,In_680,In_615);
and U3666 (N_3666,In_331,In_53);
or U3667 (N_3667,In_994,In_303);
nor U3668 (N_3668,In_190,In_957);
and U3669 (N_3669,In_856,In_999);
nand U3670 (N_3670,In_433,In_740);
and U3671 (N_3671,In_787,In_347);
or U3672 (N_3672,In_498,In_265);
nand U3673 (N_3673,In_467,In_966);
nor U3674 (N_3674,In_175,In_421);
nand U3675 (N_3675,In_492,In_300);
nor U3676 (N_3676,In_676,In_964);
or U3677 (N_3677,In_92,In_455);
or U3678 (N_3678,In_335,In_686);
and U3679 (N_3679,In_741,In_547);
nand U3680 (N_3680,In_621,In_510);
nor U3681 (N_3681,In_561,In_853);
and U3682 (N_3682,In_366,In_598);
and U3683 (N_3683,In_907,In_97);
or U3684 (N_3684,In_483,In_865);
and U3685 (N_3685,In_516,In_208);
and U3686 (N_3686,In_998,In_221);
nand U3687 (N_3687,In_455,In_723);
or U3688 (N_3688,In_13,In_565);
and U3689 (N_3689,In_149,In_932);
nor U3690 (N_3690,In_838,In_412);
and U3691 (N_3691,In_903,In_766);
or U3692 (N_3692,In_800,In_604);
nor U3693 (N_3693,In_210,In_446);
and U3694 (N_3694,In_464,In_989);
nand U3695 (N_3695,In_669,In_694);
nor U3696 (N_3696,In_650,In_985);
or U3697 (N_3697,In_158,In_615);
nor U3698 (N_3698,In_508,In_319);
and U3699 (N_3699,In_832,In_197);
and U3700 (N_3700,In_489,In_282);
and U3701 (N_3701,In_889,In_629);
or U3702 (N_3702,In_360,In_190);
and U3703 (N_3703,In_245,In_870);
nor U3704 (N_3704,In_72,In_23);
nor U3705 (N_3705,In_569,In_607);
or U3706 (N_3706,In_1,In_342);
nand U3707 (N_3707,In_137,In_402);
or U3708 (N_3708,In_364,In_877);
nor U3709 (N_3709,In_360,In_104);
or U3710 (N_3710,In_21,In_491);
nand U3711 (N_3711,In_955,In_526);
or U3712 (N_3712,In_208,In_236);
and U3713 (N_3713,In_762,In_903);
and U3714 (N_3714,In_469,In_848);
nor U3715 (N_3715,In_750,In_833);
nand U3716 (N_3716,In_395,In_14);
nor U3717 (N_3717,In_257,In_513);
and U3718 (N_3718,In_179,In_737);
nand U3719 (N_3719,In_725,In_644);
and U3720 (N_3720,In_334,In_21);
and U3721 (N_3721,In_659,In_35);
nor U3722 (N_3722,In_892,In_863);
nor U3723 (N_3723,In_805,In_871);
and U3724 (N_3724,In_144,In_837);
nor U3725 (N_3725,In_279,In_502);
or U3726 (N_3726,In_872,In_66);
and U3727 (N_3727,In_38,In_369);
xnor U3728 (N_3728,In_228,In_331);
nor U3729 (N_3729,In_386,In_940);
nand U3730 (N_3730,In_311,In_338);
nand U3731 (N_3731,In_963,In_175);
nand U3732 (N_3732,In_176,In_699);
nand U3733 (N_3733,In_160,In_358);
nor U3734 (N_3734,In_369,In_760);
or U3735 (N_3735,In_736,In_192);
and U3736 (N_3736,In_868,In_80);
nor U3737 (N_3737,In_809,In_745);
and U3738 (N_3738,In_129,In_869);
nor U3739 (N_3739,In_413,In_970);
or U3740 (N_3740,In_234,In_988);
nand U3741 (N_3741,In_120,In_738);
or U3742 (N_3742,In_986,In_737);
and U3743 (N_3743,In_201,In_213);
and U3744 (N_3744,In_871,In_957);
and U3745 (N_3745,In_602,In_48);
nor U3746 (N_3746,In_557,In_970);
nor U3747 (N_3747,In_681,In_20);
nand U3748 (N_3748,In_178,In_906);
nor U3749 (N_3749,In_321,In_486);
nor U3750 (N_3750,In_727,In_358);
nand U3751 (N_3751,In_56,In_622);
or U3752 (N_3752,In_972,In_30);
nand U3753 (N_3753,In_546,In_114);
and U3754 (N_3754,In_626,In_949);
nor U3755 (N_3755,In_252,In_396);
nand U3756 (N_3756,In_635,In_533);
or U3757 (N_3757,In_745,In_187);
nand U3758 (N_3758,In_169,In_258);
or U3759 (N_3759,In_297,In_982);
nor U3760 (N_3760,In_145,In_61);
and U3761 (N_3761,In_900,In_155);
or U3762 (N_3762,In_33,In_560);
nor U3763 (N_3763,In_27,In_655);
and U3764 (N_3764,In_856,In_34);
and U3765 (N_3765,In_652,In_21);
nor U3766 (N_3766,In_814,In_644);
nor U3767 (N_3767,In_937,In_51);
xor U3768 (N_3768,In_102,In_753);
and U3769 (N_3769,In_138,In_585);
nand U3770 (N_3770,In_656,In_496);
or U3771 (N_3771,In_773,In_959);
and U3772 (N_3772,In_12,In_293);
or U3773 (N_3773,In_121,In_774);
and U3774 (N_3774,In_43,In_701);
nand U3775 (N_3775,In_836,In_613);
nor U3776 (N_3776,In_551,In_793);
nor U3777 (N_3777,In_747,In_486);
nand U3778 (N_3778,In_157,In_538);
or U3779 (N_3779,In_196,In_768);
or U3780 (N_3780,In_811,In_102);
or U3781 (N_3781,In_607,In_390);
nor U3782 (N_3782,In_340,In_669);
nand U3783 (N_3783,In_994,In_275);
nand U3784 (N_3784,In_8,In_372);
nor U3785 (N_3785,In_711,In_621);
nor U3786 (N_3786,In_979,In_258);
and U3787 (N_3787,In_810,In_140);
and U3788 (N_3788,In_515,In_564);
nor U3789 (N_3789,In_872,In_352);
nor U3790 (N_3790,In_164,In_163);
and U3791 (N_3791,In_699,In_860);
nor U3792 (N_3792,In_155,In_274);
nor U3793 (N_3793,In_773,In_825);
nand U3794 (N_3794,In_824,In_962);
or U3795 (N_3795,In_802,In_211);
and U3796 (N_3796,In_623,In_110);
and U3797 (N_3797,In_678,In_135);
nand U3798 (N_3798,In_57,In_2);
and U3799 (N_3799,In_38,In_831);
nand U3800 (N_3800,In_477,In_635);
or U3801 (N_3801,In_22,In_4);
or U3802 (N_3802,In_979,In_441);
nor U3803 (N_3803,In_542,In_416);
or U3804 (N_3804,In_908,In_448);
and U3805 (N_3805,In_786,In_510);
and U3806 (N_3806,In_888,In_985);
nand U3807 (N_3807,In_477,In_671);
and U3808 (N_3808,In_914,In_989);
and U3809 (N_3809,In_859,In_103);
and U3810 (N_3810,In_286,In_855);
nand U3811 (N_3811,In_823,In_370);
and U3812 (N_3812,In_485,In_911);
and U3813 (N_3813,In_946,In_37);
and U3814 (N_3814,In_921,In_890);
nand U3815 (N_3815,In_708,In_360);
nor U3816 (N_3816,In_929,In_783);
nor U3817 (N_3817,In_298,In_457);
nor U3818 (N_3818,In_363,In_119);
nand U3819 (N_3819,In_551,In_209);
nand U3820 (N_3820,In_613,In_173);
and U3821 (N_3821,In_268,In_761);
nand U3822 (N_3822,In_132,In_643);
nor U3823 (N_3823,In_389,In_757);
nand U3824 (N_3824,In_187,In_108);
and U3825 (N_3825,In_976,In_872);
nor U3826 (N_3826,In_178,In_668);
or U3827 (N_3827,In_918,In_457);
nor U3828 (N_3828,In_110,In_200);
and U3829 (N_3829,In_275,In_299);
and U3830 (N_3830,In_97,In_622);
nor U3831 (N_3831,In_113,In_697);
or U3832 (N_3832,In_452,In_273);
or U3833 (N_3833,In_364,In_957);
and U3834 (N_3834,In_113,In_810);
nor U3835 (N_3835,In_673,In_620);
nand U3836 (N_3836,In_176,In_351);
nand U3837 (N_3837,In_708,In_491);
or U3838 (N_3838,In_87,In_284);
nor U3839 (N_3839,In_394,In_750);
nand U3840 (N_3840,In_423,In_338);
nand U3841 (N_3841,In_6,In_501);
and U3842 (N_3842,In_918,In_591);
and U3843 (N_3843,In_694,In_179);
nand U3844 (N_3844,In_572,In_417);
and U3845 (N_3845,In_138,In_201);
and U3846 (N_3846,In_906,In_556);
and U3847 (N_3847,In_719,In_482);
or U3848 (N_3848,In_277,In_684);
nor U3849 (N_3849,In_797,In_493);
or U3850 (N_3850,In_239,In_208);
or U3851 (N_3851,In_603,In_714);
and U3852 (N_3852,In_815,In_74);
or U3853 (N_3853,In_708,In_182);
nor U3854 (N_3854,In_976,In_506);
and U3855 (N_3855,In_203,In_153);
or U3856 (N_3856,In_931,In_416);
and U3857 (N_3857,In_931,In_642);
or U3858 (N_3858,In_532,In_700);
nor U3859 (N_3859,In_229,In_14);
or U3860 (N_3860,In_497,In_937);
nor U3861 (N_3861,In_139,In_518);
or U3862 (N_3862,In_216,In_61);
nor U3863 (N_3863,In_317,In_954);
and U3864 (N_3864,In_999,In_287);
and U3865 (N_3865,In_612,In_366);
nand U3866 (N_3866,In_179,In_856);
nor U3867 (N_3867,In_45,In_194);
and U3868 (N_3868,In_356,In_910);
and U3869 (N_3869,In_968,In_373);
and U3870 (N_3870,In_403,In_38);
or U3871 (N_3871,In_160,In_272);
nand U3872 (N_3872,In_76,In_507);
or U3873 (N_3873,In_877,In_97);
nand U3874 (N_3874,In_282,In_378);
nand U3875 (N_3875,In_348,In_556);
and U3876 (N_3876,In_460,In_813);
nand U3877 (N_3877,In_246,In_766);
nand U3878 (N_3878,In_545,In_462);
nand U3879 (N_3879,In_619,In_215);
or U3880 (N_3880,In_199,In_235);
nand U3881 (N_3881,In_186,In_853);
or U3882 (N_3882,In_17,In_656);
nand U3883 (N_3883,In_377,In_932);
nand U3884 (N_3884,In_22,In_574);
nor U3885 (N_3885,In_383,In_992);
nand U3886 (N_3886,In_889,In_711);
or U3887 (N_3887,In_276,In_550);
nor U3888 (N_3888,In_832,In_708);
nand U3889 (N_3889,In_669,In_186);
nand U3890 (N_3890,In_846,In_937);
nand U3891 (N_3891,In_568,In_743);
or U3892 (N_3892,In_182,In_419);
and U3893 (N_3893,In_296,In_868);
xnor U3894 (N_3894,In_204,In_582);
nor U3895 (N_3895,In_398,In_224);
nand U3896 (N_3896,In_781,In_417);
nand U3897 (N_3897,In_237,In_427);
or U3898 (N_3898,In_397,In_931);
nand U3899 (N_3899,In_773,In_152);
nand U3900 (N_3900,In_203,In_746);
or U3901 (N_3901,In_733,In_492);
or U3902 (N_3902,In_213,In_705);
nor U3903 (N_3903,In_655,In_647);
nand U3904 (N_3904,In_462,In_307);
nand U3905 (N_3905,In_133,In_810);
nand U3906 (N_3906,In_640,In_927);
nor U3907 (N_3907,In_564,In_843);
and U3908 (N_3908,In_617,In_827);
nor U3909 (N_3909,In_782,In_803);
and U3910 (N_3910,In_540,In_351);
and U3911 (N_3911,In_715,In_551);
or U3912 (N_3912,In_822,In_933);
nor U3913 (N_3913,In_96,In_121);
nor U3914 (N_3914,In_161,In_977);
nand U3915 (N_3915,In_536,In_915);
and U3916 (N_3916,In_369,In_753);
or U3917 (N_3917,In_264,In_694);
or U3918 (N_3918,In_575,In_150);
nor U3919 (N_3919,In_343,In_622);
nor U3920 (N_3920,In_248,In_236);
or U3921 (N_3921,In_363,In_108);
or U3922 (N_3922,In_698,In_785);
nor U3923 (N_3923,In_996,In_209);
or U3924 (N_3924,In_725,In_574);
or U3925 (N_3925,In_426,In_818);
and U3926 (N_3926,In_8,In_383);
and U3927 (N_3927,In_309,In_471);
or U3928 (N_3928,In_399,In_263);
xnor U3929 (N_3929,In_686,In_694);
nor U3930 (N_3930,In_10,In_902);
nand U3931 (N_3931,In_192,In_655);
nand U3932 (N_3932,In_618,In_574);
nor U3933 (N_3933,In_517,In_968);
or U3934 (N_3934,In_881,In_296);
nand U3935 (N_3935,In_154,In_616);
or U3936 (N_3936,In_473,In_639);
or U3937 (N_3937,In_195,In_854);
nor U3938 (N_3938,In_884,In_231);
and U3939 (N_3939,In_29,In_934);
or U3940 (N_3940,In_441,In_706);
or U3941 (N_3941,In_195,In_625);
nand U3942 (N_3942,In_814,In_187);
or U3943 (N_3943,In_764,In_921);
nor U3944 (N_3944,In_252,In_167);
and U3945 (N_3945,In_40,In_287);
nand U3946 (N_3946,In_642,In_874);
or U3947 (N_3947,In_738,In_260);
nand U3948 (N_3948,In_304,In_213);
nor U3949 (N_3949,In_687,In_338);
and U3950 (N_3950,In_578,In_296);
nor U3951 (N_3951,In_911,In_461);
and U3952 (N_3952,In_637,In_130);
nor U3953 (N_3953,In_943,In_584);
nor U3954 (N_3954,In_15,In_990);
nand U3955 (N_3955,In_697,In_926);
and U3956 (N_3956,In_136,In_842);
or U3957 (N_3957,In_211,In_963);
and U3958 (N_3958,In_406,In_112);
and U3959 (N_3959,In_556,In_432);
nor U3960 (N_3960,In_211,In_29);
and U3961 (N_3961,In_318,In_599);
nor U3962 (N_3962,In_779,In_987);
nand U3963 (N_3963,In_308,In_97);
nor U3964 (N_3964,In_626,In_436);
nand U3965 (N_3965,In_997,In_94);
and U3966 (N_3966,In_306,In_272);
nor U3967 (N_3967,In_108,In_90);
or U3968 (N_3968,In_217,In_115);
nor U3969 (N_3969,In_502,In_629);
nor U3970 (N_3970,In_707,In_724);
and U3971 (N_3971,In_852,In_201);
nor U3972 (N_3972,In_588,In_86);
nor U3973 (N_3973,In_899,In_563);
and U3974 (N_3974,In_496,In_268);
nand U3975 (N_3975,In_219,In_223);
nand U3976 (N_3976,In_747,In_364);
and U3977 (N_3977,In_970,In_720);
nor U3978 (N_3978,In_186,In_484);
nand U3979 (N_3979,In_875,In_186);
or U3980 (N_3980,In_857,In_612);
nand U3981 (N_3981,In_151,In_949);
or U3982 (N_3982,In_184,In_524);
or U3983 (N_3983,In_165,In_713);
or U3984 (N_3984,In_140,In_282);
or U3985 (N_3985,In_785,In_967);
and U3986 (N_3986,In_78,In_723);
nand U3987 (N_3987,In_688,In_604);
or U3988 (N_3988,In_674,In_620);
nor U3989 (N_3989,In_266,In_201);
nand U3990 (N_3990,In_343,In_775);
nand U3991 (N_3991,In_186,In_852);
and U3992 (N_3992,In_82,In_780);
xor U3993 (N_3993,In_903,In_41);
nor U3994 (N_3994,In_412,In_416);
nand U3995 (N_3995,In_132,In_753);
nor U3996 (N_3996,In_178,In_893);
xor U3997 (N_3997,In_569,In_963);
and U3998 (N_3998,In_845,In_995);
nand U3999 (N_3999,In_855,In_482);
nor U4000 (N_4000,In_220,In_370);
nand U4001 (N_4001,In_647,In_313);
nand U4002 (N_4002,In_963,In_416);
or U4003 (N_4003,In_311,In_51);
nand U4004 (N_4004,In_558,In_611);
or U4005 (N_4005,In_94,In_28);
or U4006 (N_4006,In_965,In_198);
or U4007 (N_4007,In_428,In_664);
nand U4008 (N_4008,In_370,In_274);
or U4009 (N_4009,In_178,In_299);
nand U4010 (N_4010,In_94,In_781);
nor U4011 (N_4011,In_304,In_876);
and U4012 (N_4012,In_878,In_371);
and U4013 (N_4013,In_365,In_369);
and U4014 (N_4014,In_446,In_173);
and U4015 (N_4015,In_252,In_990);
and U4016 (N_4016,In_238,In_815);
nor U4017 (N_4017,In_807,In_184);
and U4018 (N_4018,In_387,In_406);
and U4019 (N_4019,In_194,In_124);
nand U4020 (N_4020,In_952,In_138);
or U4021 (N_4021,In_598,In_373);
nor U4022 (N_4022,In_930,In_527);
and U4023 (N_4023,In_797,In_112);
and U4024 (N_4024,In_447,In_697);
nor U4025 (N_4025,In_704,In_885);
or U4026 (N_4026,In_42,In_679);
and U4027 (N_4027,In_972,In_692);
and U4028 (N_4028,In_777,In_193);
nand U4029 (N_4029,In_120,In_329);
nor U4030 (N_4030,In_825,In_660);
or U4031 (N_4031,In_322,In_794);
nor U4032 (N_4032,In_441,In_976);
and U4033 (N_4033,In_519,In_281);
and U4034 (N_4034,In_665,In_946);
nor U4035 (N_4035,In_630,In_703);
and U4036 (N_4036,In_280,In_694);
nor U4037 (N_4037,In_323,In_280);
and U4038 (N_4038,In_697,In_550);
or U4039 (N_4039,In_935,In_434);
or U4040 (N_4040,In_376,In_667);
and U4041 (N_4041,In_930,In_433);
or U4042 (N_4042,In_38,In_288);
and U4043 (N_4043,In_373,In_403);
nand U4044 (N_4044,In_140,In_953);
nor U4045 (N_4045,In_537,In_523);
nand U4046 (N_4046,In_842,In_455);
or U4047 (N_4047,In_576,In_150);
nor U4048 (N_4048,In_199,In_234);
nor U4049 (N_4049,In_533,In_604);
nor U4050 (N_4050,In_159,In_501);
nor U4051 (N_4051,In_86,In_143);
nand U4052 (N_4052,In_79,In_39);
nand U4053 (N_4053,In_624,In_238);
nor U4054 (N_4054,In_249,In_23);
nand U4055 (N_4055,In_658,In_98);
nand U4056 (N_4056,In_934,In_303);
or U4057 (N_4057,In_600,In_140);
or U4058 (N_4058,In_272,In_238);
or U4059 (N_4059,In_76,In_49);
and U4060 (N_4060,In_153,In_736);
nand U4061 (N_4061,In_538,In_398);
and U4062 (N_4062,In_662,In_264);
nand U4063 (N_4063,In_894,In_691);
nand U4064 (N_4064,In_458,In_443);
or U4065 (N_4065,In_977,In_95);
nand U4066 (N_4066,In_207,In_348);
and U4067 (N_4067,In_49,In_732);
nor U4068 (N_4068,In_6,In_229);
and U4069 (N_4069,In_675,In_37);
nand U4070 (N_4070,In_551,In_857);
nor U4071 (N_4071,In_297,In_160);
and U4072 (N_4072,In_782,In_175);
and U4073 (N_4073,In_43,In_910);
and U4074 (N_4074,In_93,In_856);
and U4075 (N_4075,In_439,In_92);
and U4076 (N_4076,In_804,In_831);
or U4077 (N_4077,In_778,In_981);
or U4078 (N_4078,In_201,In_6);
or U4079 (N_4079,In_488,In_446);
nor U4080 (N_4080,In_246,In_111);
or U4081 (N_4081,In_840,In_691);
nor U4082 (N_4082,In_267,In_546);
or U4083 (N_4083,In_48,In_490);
nor U4084 (N_4084,In_266,In_246);
nor U4085 (N_4085,In_320,In_876);
nor U4086 (N_4086,In_77,In_819);
nor U4087 (N_4087,In_327,In_693);
nand U4088 (N_4088,In_785,In_193);
nand U4089 (N_4089,In_828,In_104);
nor U4090 (N_4090,In_47,In_33);
nand U4091 (N_4091,In_197,In_580);
and U4092 (N_4092,In_778,In_782);
nor U4093 (N_4093,In_164,In_690);
nand U4094 (N_4094,In_837,In_257);
nor U4095 (N_4095,In_77,In_25);
or U4096 (N_4096,In_438,In_854);
or U4097 (N_4097,In_456,In_614);
nand U4098 (N_4098,In_816,In_187);
and U4099 (N_4099,In_97,In_577);
and U4100 (N_4100,In_288,In_934);
or U4101 (N_4101,In_310,In_312);
or U4102 (N_4102,In_606,In_620);
or U4103 (N_4103,In_525,In_532);
and U4104 (N_4104,In_526,In_527);
nand U4105 (N_4105,In_423,In_98);
nor U4106 (N_4106,In_774,In_83);
or U4107 (N_4107,In_546,In_876);
or U4108 (N_4108,In_316,In_818);
or U4109 (N_4109,In_649,In_159);
and U4110 (N_4110,In_772,In_839);
and U4111 (N_4111,In_403,In_379);
nor U4112 (N_4112,In_348,In_138);
nor U4113 (N_4113,In_549,In_317);
nand U4114 (N_4114,In_565,In_609);
and U4115 (N_4115,In_110,In_60);
nor U4116 (N_4116,In_25,In_222);
or U4117 (N_4117,In_975,In_801);
and U4118 (N_4118,In_267,In_98);
and U4119 (N_4119,In_280,In_731);
and U4120 (N_4120,In_15,In_57);
and U4121 (N_4121,In_237,In_253);
and U4122 (N_4122,In_56,In_336);
nand U4123 (N_4123,In_230,In_239);
nand U4124 (N_4124,In_63,In_775);
and U4125 (N_4125,In_652,In_756);
nor U4126 (N_4126,In_532,In_128);
nor U4127 (N_4127,In_829,In_633);
nor U4128 (N_4128,In_609,In_655);
and U4129 (N_4129,In_679,In_660);
or U4130 (N_4130,In_751,In_219);
nand U4131 (N_4131,In_914,In_31);
and U4132 (N_4132,In_548,In_775);
nand U4133 (N_4133,In_117,In_632);
or U4134 (N_4134,In_607,In_596);
or U4135 (N_4135,In_748,In_978);
nand U4136 (N_4136,In_717,In_138);
or U4137 (N_4137,In_827,In_44);
nand U4138 (N_4138,In_523,In_985);
nor U4139 (N_4139,In_913,In_605);
and U4140 (N_4140,In_569,In_343);
nand U4141 (N_4141,In_84,In_434);
nand U4142 (N_4142,In_84,In_594);
nand U4143 (N_4143,In_742,In_853);
and U4144 (N_4144,In_599,In_521);
nor U4145 (N_4145,In_747,In_696);
and U4146 (N_4146,In_795,In_123);
and U4147 (N_4147,In_110,In_422);
or U4148 (N_4148,In_217,In_199);
and U4149 (N_4149,In_179,In_537);
and U4150 (N_4150,In_509,In_676);
nor U4151 (N_4151,In_918,In_518);
or U4152 (N_4152,In_971,In_831);
nor U4153 (N_4153,In_336,In_830);
nor U4154 (N_4154,In_244,In_973);
and U4155 (N_4155,In_980,In_720);
and U4156 (N_4156,In_27,In_97);
and U4157 (N_4157,In_970,In_461);
nand U4158 (N_4158,In_515,In_582);
nand U4159 (N_4159,In_967,In_591);
or U4160 (N_4160,In_652,In_620);
and U4161 (N_4161,In_439,In_67);
or U4162 (N_4162,In_445,In_495);
nand U4163 (N_4163,In_994,In_877);
or U4164 (N_4164,In_628,In_764);
nand U4165 (N_4165,In_699,In_686);
and U4166 (N_4166,In_926,In_97);
or U4167 (N_4167,In_313,In_437);
nor U4168 (N_4168,In_488,In_929);
nor U4169 (N_4169,In_351,In_64);
or U4170 (N_4170,In_189,In_456);
and U4171 (N_4171,In_319,In_785);
nor U4172 (N_4172,In_927,In_129);
and U4173 (N_4173,In_926,In_169);
nand U4174 (N_4174,In_599,In_253);
nor U4175 (N_4175,In_779,In_542);
nand U4176 (N_4176,In_915,In_192);
and U4177 (N_4177,In_769,In_254);
or U4178 (N_4178,In_229,In_974);
nand U4179 (N_4179,In_143,In_715);
nor U4180 (N_4180,In_573,In_185);
nand U4181 (N_4181,In_317,In_819);
and U4182 (N_4182,In_236,In_980);
and U4183 (N_4183,In_894,In_538);
or U4184 (N_4184,In_36,In_861);
nand U4185 (N_4185,In_373,In_449);
nor U4186 (N_4186,In_329,In_94);
nor U4187 (N_4187,In_570,In_543);
and U4188 (N_4188,In_594,In_270);
nor U4189 (N_4189,In_990,In_681);
or U4190 (N_4190,In_5,In_373);
or U4191 (N_4191,In_725,In_582);
nand U4192 (N_4192,In_545,In_155);
or U4193 (N_4193,In_304,In_941);
nand U4194 (N_4194,In_216,In_647);
and U4195 (N_4195,In_200,In_264);
nand U4196 (N_4196,In_325,In_928);
and U4197 (N_4197,In_160,In_980);
and U4198 (N_4198,In_922,In_349);
nand U4199 (N_4199,In_266,In_953);
xnor U4200 (N_4200,In_313,In_682);
or U4201 (N_4201,In_231,In_204);
and U4202 (N_4202,In_708,In_228);
or U4203 (N_4203,In_875,In_170);
nand U4204 (N_4204,In_606,In_485);
or U4205 (N_4205,In_758,In_504);
nand U4206 (N_4206,In_791,In_128);
and U4207 (N_4207,In_588,In_479);
nor U4208 (N_4208,In_867,In_574);
nand U4209 (N_4209,In_251,In_258);
nor U4210 (N_4210,In_0,In_934);
or U4211 (N_4211,In_179,In_107);
nand U4212 (N_4212,In_67,In_508);
and U4213 (N_4213,In_677,In_64);
and U4214 (N_4214,In_965,In_363);
or U4215 (N_4215,In_172,In_294);
and U4216 (N_4216,In_372,In_542);
nand U4217 (N_4217,In_700,In_819);
and U4218 (N_4218,In_623,In_80);
and U4219 (N_4219,In_55,In_464);
nor U4220 (N_4220,In_305,In_557);
nand U4221 (N_4221,In_458,In_242);
nor U4222 (N_4222,In_298,In_902);
and U4223 (N_4223,In_476,In_127);
or U4224 (N_4224,In_75,In_567);
nand U4225 (N_4225,In_349,In_845);
and U4226 (N_4226,In_965,In_387);
or U4227 (N_4227,In_346,In_397);
nand U4228 (N_4228,In_717,In_687);
nand U4229 (N_4229,In_838,In_368);
and U4230 (N_4230,In_390,In_589);
or U4231 (N_4231,In_248,In_697);
and U4232 (N_4232,In_511,In_57);
nand U4233 (N_4233,In_461,In_601);
and U4234 (N_4234,In_551,In_947);
and U4235 (N_4235,In_27,In_791);
or U4236 (N_4236,In_769,In_262);
or U4237 (N_4237,In_412,In_226);
and U4238 (N_4238,In_868,In_28);
nor U4239 (N_4239,In_38,In_294);
nor U4240 (N_4240,In_853,In_379);
nor U4241 (N_4241,In_789,In_231);
nor U4242 (N_4242,In_284,In_853);
and U4243 (N_4243,In_283,In_344);
and U4244 (N_4244,In_3,In_193);
nand U4245 (N_4245,In_235,In_195);
nand U4246 (N_4246,In_502,In_993);
and U4247 (N_4247,In_676,In_827);
and U4248 (N_4248,In_271,In_252);
nor U4249 (N_4249,In_376,In_836);
or U4250 (N_4250,In_734,In_102);
nor U4251 (N_4251,In_33,In_795);
or U4252 (N_4252,In_388,In_675);
nor U4253 (N_4253,In_412,In_431);
nor U4254 (N_4254,In_303,In_495);
nor U4255 (N_4255,In_525,In_95);
nand U4256 (N_4256,In_777,In_543);
or U4257 (N_4257,In_486,In_100);
nor U4258 (N_4258,In_247,In_239);
nand U4259 (N_4259,In_288,In_581);
nand U4260 (N_4260,In_631,In_933);
and U4261 (N_4261,In_771,In_47);
nand U4262 (N_4262,In_822,In_873);
nor U4263 (N_4263,In_431,In_666);
nor U4264 (N_4264,In_279,In_540);
nand U4265 (N_4265,In_404,In_286);
nand U4266 (N_4266,In_345,In_592);
and U4267 (N_4267,In_952,In_323);
or U4268 (N_4268,In_759,In_825);
or U4269 (N_4269,In_507,In_254);
nor U4270 (N_4270,In_367,In_490);
or U4271 (N_4271,In_215,In_89);
or U4272 (N_4272,In_337,In_411);
and U4273 (N_4273,In_506,In_704);
nand U4274 (N_4274,In_892,In_202);
or U4275 (N_4275,In_827,In_757);
nor U4276 (N_4276,In_144,In_461);
nor U4277 (N_4277,In_859,In_640);
xor U4278 (N_4278,In_180,In_996);
or U4279 (N_4279,In_566,In_18);
and U4280 (N_4280,In_914,In_860);
and U4281 (N_4281,In_462,In_328);
nor U4282 (N_4282,In_539,In_19);
and U4283 (N_4283,In_260,In_124);
nand U4284 (N_4284,In_104,In_691);
nor U4285 (N_4285,In_380,In_959);
or U4286 (N_4286,In_479,In_234);
nor U4287 (N_4287,In_611,In_26);
nand U4288 (N_4288,In_117,In_661);
and U4289 (N_4289,In_292,In_852);
nor U4290 (N_4290,In_769,In_971);
xnor U4291 (N_4291,In_242,In_727);
nor U4292 (N_4292,In_963,In_894);
nor U4293 (N_4293,In_106,In_750);
nor U4294 (N_4294,In_244,In_986);
nand U4295 (N_4295,In_323,In_336);
nor U4296 (N_4296,In_98,In_470);
or U4297 (N_4297,In_497,In_470);
nand U4298 (N_4298,In_50,In_439);
nor U4299 (N_4299,In_663,In_71);
nor U4300 (N_4300,In_687,In_729);
and U4301 (N_4301,In_450,In_433);
or U4302 (N_4302,In_364,In_909);
nor U4303 (N_4303,In_937,In_32);
and U4304 (N_4304,In_959,In_531);
or U4305 (N_4305,In_242,In_59);
or U4306 (N_4306,In_974,In_322);
nand U4307 (N_4307,In_444,In_590);
or U4308 (N_4308,In_547,In_651);
nand U4309 (N_4309,In_288,In_520);
and U4310 (N_4310,In_935,In_961);
nand U4311 (N_4311,In_983,In_730);
nor U4312 (N_4312,In_446,In_737);
nor U4313 (N_4313,In_496,In_114);
and U4314 (N_4314,In_463,In_206);
or U4315 (N_4315,In_193,In_478);
or U4316 (N_4316,In_308,In_393);
nor U4317 (N_4317,In_449,In_738);
and U4318 (N_4318,In_67,In_797);
nor U4319 (N_4319,In_581,In_847);
and U4320 (N_4320,In_321,In_16);
xnor U4321 (N_4321,In_590,In_656);
nor U4322 (N_4322,In_451,In_229);
nor U4323 (N_4323,In_834,In_404);
nand U4324 (N_4324,In_31,In_145);
nand U4325 (N_4325,In_408,In_643);
and U4326 (N_4326,In_792,In_243);
or U4327 (N_4327,In_376,In_998);
nand U4328 (N_4328,In_861,In_544);
nor U4329 (N_4329,In_120,In_795);
or U4330 (N_4330,In_205,In_509);
or U4331 (N_4331,In_677,In_118);
and U4332 (N_4332,In_901,In_134);
nand U4333 (N_4333,In_369,In_941);
nor U4334 (N_4334,In_315,In_983);
or U4335 (N_4335,In_783,In_550);
nand U4336 (N_4336,In_159,In_426);
and U4337 (N_4337,In_303,In_263);
nor U4338 (N_4338,In_406,In_511);
or U4339 (N_4339,In_616,In_166);
and U4340 (N_4340,In_319,In_774);
or U4341 (N_4341,In_394,In_380);
and U4342 (N_4342,In_997,In_758);
nor U4343 (N_4343,In_270,In_350);
nand U4344 (N_4344,In_976,In_816);
nor U4345 (N_4345,In_127,In_919);
or U4346 (N_4346,In_59,In_630);
nand U4347 (N_4347,In_738,In_771);
or U4348 (N_4348,In_692,In_512);
and U4349 (N_4349,In_585,In_834);
and U4350 (N_4350,In_616,In_829);
nand U4351 (N_4351,In_104,In_861);
nand U4352 (N_4352,In_261,In_414);
and U4353 (N_4353,In_271,In_469);
and U4354 (N_4354,In_93,In_103);
nor U4355 (N_4355,In_7,In_902);
nor U4356 (N_4356,In_782,In_473);
or U4357 (N_4357,In_431,In_388);
and U4358 (N_4358,In_208,In_285);
and U4359 (N_4359,In_964,In_926);
or U4360 (N_4360,In_305,In_511);
nand U4361 (N_4361,In_628,In_672);
and U4362 (N_4362,In_999,In_101);
nand U4363 (N_4363,In_346,In_560);
xnor U4364 (N_4364,In_130,In_164);
and U4365 (N_4365,In_442,In_718);
or U4366 (N_4366,In_993,In_702);
nor U4367 (N_4367,In_503,In_142);
or U4368 (N_4368,In_515,In_506);
and U4369 (N_4369,In_433,In_518);
or U4370 (N_4370,In_93,In_33);
and U4371 (N_4371,In_452,In_123);
nand U4372 (N_4372,In_745,In_168);
or U4373 (N_4373,In_148,In_440);
and U4374 (N_4374,In_472,In_837);
nor U4375 (N_4375,In_741,In_51);
nand U4376 (N_4376,In_316,In_9);
nand U4377 (N_4377,In_374,In_85);
nor U4378 (N_4378,In_662,In_576);
nand U4379 (N_4379,In_806,In_543);
and U4380 (N_4380,In_113,In_833);
and U4381 (N_4381,In_509,In_648);
and U4382 (N_4382,In_916,In_154);
and U4383 (N_4383,In_531,In_53);
nand U4384 (N_4384,In_900,In_926);
nand U4385 (N_4385,In_213,In_643);
and U4386 (N_4386,In_594,In_839);
nand U4387 (N_4387,In_947,In_147);
or U4388 (N_4388,In_147,In_888);
or U4389 (N_4389,In_23,In_936);
nor U4390 (N_4390,In_433,In_985);
xor U4391 (N_4391,In_252,In_665);
or U4392 (N_4392,In_284,In_929);
nor U4393 (N_4393,In_102,In_497);
nor U4394 (N_4394,In_552,In_193);
nand U4395 (N_4395,In_419,In_51);
or U4396 (N_4396,In_85,In_397);
and U4397 (N_4397,In_410,In_801);
or U4398 (N_4398,In_350,In_44);
nor U4399 (N_4399,In_992,In_108);
nor U4400 (N_4400,In_397,In_126);
nand U4401 (N_4401,In_229,In_386);
nor U4402 (N_4402,In_784,In_490);
nor U4403 (N_4403,In_752,In_186);
or U4404 (N_4404,In_46,In_748);
or U4405 (N_4405,In_19,In_533);
nand U4406 (N_4406,In_748,In_371);
and U4407 (N_4407,In_387,In_657);
or U4408 (N_4408,In_789,In_100);
or U4409 (N_4409,In_429,In_876);
nand U4410 (N_4410,In_731,In_663);
nand U4411 (N_4411,In_135,In_23);
or U4412 (N_4412,In_410,In_497);
nand U4413 (N_4413,In_453,In_651);
nand U4414 (N_4414,In_328,In_840);
nor U4415 (N_4415,In_318,In_642);
nand U4416 (N_4416,In_529,In_782);
nor U4417 (N_4417,In_230,In_980);
and U4418 (N_4418,In_968,In_978);
and U4419 (N_4419,In_577,In_171);
or U4420 (N_4420,In_753,In_44);
nand U4421 (N_4421,In_406,In_146);
and U4422 (N_4422,In_502,In_999);
or U4423 (N_4423,In_706,In_68);
nor U4424 (N_4424,In_336,In_138);
nor U4425 (N_4425,In_1,In_410);
nor U4426 (N_4426,In_923,In_194);
and U4427 (N_4427,In_959,In_812);
and U4428 (N_4428,In_410,In_546);
and U4429 (N_4429,In_385,In_629);
nor U4430 (N_4430,In_97,In_193);
nand U4431 (N_4431,In_938,In_766);
or U4432 (N_4432,In_844,In_802);
nand U4433 (N_4433,In_710,In_513);
nand U4434 (N_4434,In_109,In_278);
and U4435 (N_4435,In_241,In_128);
or U4436 (N_4436,In_333,In_501);
or U4437 (N_4437,In_207,In_787);
or U4438 (N_4438,In_720,In_201);
or U4439 (N_4439,In_720,In_89);
nand U4440 (N_4440,In_243,In_286);
nand U4441 (N_4441,In_965,In_296);
nand U4442 (N_4442,In_50,In_75);
and U4443 (N_4443,In_697,In_331);
and U4444 (N_4444,In_198,In_29);
nand U4445 (N_4445,In_658,In_971);
and U4446 (N_4446,In_912,In_221);
nor U4447 (N_4447,In_945,In_45);
or U4448 (N_4448,In_880,In_968);
nor U4449 (N_4449,In_853,In_513);
or U4450 (N_4450,In_807,In_574);
nor U4451 (N_4451,In_8,In_683);
and U4452 (N_4452,In_362,In_828);
or U4453 (N_4453,In_857,In_318);
and U4454 (N_4454,In_294,In_878);
or U4455 (N_4455,In_424,In_97);
nor U4456 (N_4456,In_472,In_643);
nand U4457 (N_4457,In_892,In_51);
and U4458 (N_4458,In_241,In_161);
nand U4459 (N_4459,In_246,In_847);
or U4460 (N_4460,In_692,In_615);
or U4461 (N_4461,In_638,In_193);
or U4462 (N_4462,In_676,In_62);
nand U4463 (N_4463,In_817,In_896);
or U4464 (N_4464,In_529,In_208);
or U4465 (N_4465,In_928,In_755);
and U4466 (N_4466,In_237,In_752);
nand U4467 (N_4467,In_600,In_401);
or U4468 (N_4468,In_696,In_357);
or U4469 (N_4469,In_738,In_881);
and U4470 (N_4470,In_476,In_190);
or U4471 (N_4471,In_925,In_599);
nand U4472 (N_4472,In_949,In_941);
nand U4473 (N_4473,In_555,In_678);
nand U4474 (N_4474,In_277,In_233);
nor U4475 (N_4475,In_253,In_765);
nor U4476 (N_4476,In_140,In_811);
nor U4477 (N_4477,In_394,In_195);
and U4478 (N_4478,In_105,In_927);
and U4479 (N_4479,In_174,In_46);
or U4480 (N_4480,In_432,In_584);
or U4481 (N_4481,In_161,In_722);
and U4482 (N_4482,In_633,In_452);
or U4483 (N_4483,In_610,In_546);
nand U4484 (N_4484,In_742,In_268);
or U4485 (N_4485,In_544,In_31);
nor U4486 (N_4486,In_488,In_189);
nand U4487 (N_4487,In_908,In_657);
nor U4488 (N_4488,In_411,In_698);
nor U4489 (N_4489,In_674,In_467);
and U4490 (N_4490,In_311,In_440);
and U4491 (N_4491,In_926,In_339);
or U4492 (N_4492,In_542,In_402);
and U4493 (N_4493,In_670,In_548);
nand U4494 (N_4494,In_328,In_978);
nand U4495 (N_4495,In_993,In_255);
or U4496 (N_4496,In_897,In_930);
or U4497 (N_4497,In_551,In_769);
and U4498 (N_4498,In_277,In_667);
and U4499 (N_4499,In_889,In_816);
or U4500 (N_4500,In_401,In_924);
nand U4501 (N_4501,In_699,In_650);
nand U4502 (N_4502,In_500,In_557);
and U4503 (N_4503,In_916,In_66);
nand U4504 (N_4504,In_378,In_747);
xnor U4505 (N_4505,In_75,In_779);
and U4506 (N_4506,In_575,In_674);
or U4507 (N_4507,In_711,In_233);
xor U4508 (N_4508,In_944,In_620);
or U4509 (N_4509,In_429,In_343);
or U4510 (N_4510,In_962,In_686);
and U4511 (N_4511,In_277,In_858);
and U4512 (N_4512,In_45,In_541);
and U4513 (N_4513,In_222,In_130);
and U4514 (N_4514,In_233,In_849);
nor U4515 (N_4515,In_106,In_686);
nand U4516 (N_4516,In_682,In_171);
nor U4517 (N_4517,In_244,In_617);
nand U4518 (N_4518,In_448,In_98);
nand U4519 (N_4519,In_20,In_761);
nand U4520 (N_4520,In_569,In_575);
nand U4521 (N_4521,In_953,In_504);
xnor U4522 (N_4522,In_894,In_194);
or U4523 (N_4523,In_706,In_399);
or U4524 (N_4524,In_480,In_53);
nor U4525 (N_4525,In_336,In_72);
or U4526 (N_4526,In_592,In_436);
and U4527 (N_4527,In_434,In_860);
nand U4528 (N_4528,In_136,In_312);
and U4529 (N_4529,In_523,In_607);
and U4530 (N_4530,In_315,In_881);
and U4531 (N_4531,In_601,In_931);
nor U4532 (N_4532,In_9,In_690);
and U4533 (N_4533,In_817,In_814);
nand U4534 (N_4534,In_703,In_207);
nor U4535 (N_4535,In_948,In_105);
and U4536 (N_4536,In_794,In_192);
or U4537 (N_4537,In_679,In_276);
and U4538 (N_4538,In_247,In_586);
or U4539 (N_4539,In_974,In_969);
nor U4540 (N_4540,In_258,In_475);
nand U4541 (N_4541,In_747,In_954);
or U4542 (N_4542,In_359,In_86);
nor U4543 (N_4543,In_961,In_808);
and U4544 (N_4544,In_813,In_325);
nand U4545 (N_4545,In_761,In_560);
nor U4546 (N_4546,In_516,In_924);
and U4547 (N_4547,In_229,In_419);
nor U4548 (N_4548,In_926,In_811);
or U4549 (N_4549,In_643,In_947);
or U4550 (N_4550,In_603,In_114);
and U4551 (N_4551,In_327,In_1);
xor U4552 (N_4552,In_450,In_663);
nand U4553 (N_4553,In_714,In_564);
nand U4554 (N_4554,In_253,In_761);
nor U4555 (N_4555,In_740,In_101);
nand U4556 (N_4556,In_525,In_813);
or U4557 (N_4557,In_166,In_784);
and U4558 (N_4558,In_47,In_39);
nand U4559 (N_4559,In_897,In_733);
or U4560 (N_4560,In_636,In_438);
nor U4561 (N_4561,In_245,In_979);
nand U4562 (N_4562,In_519,In_126);
nand U4563 (N_4563,In_403,In_752);
nor U4564 (N_4564,In_197,In_123);
and U4565 (N_4565,In_411,In_802);
and U4566 (N_4566,In_991,In_812);
and U4567 (N_4567,In_898,In_176);
or U4568 (N_4568,In_922,In_619);
nor U4569 (N_4569,In_508,In_143);
or U4570 (N_4570,In_521,In_781);
nand U4571 (N_4571,In_893,In_863);
nor U4572 (N_4572,In_348,In_349);
or U4573 (N_4573,In_596,In_956);
or U4574 (N_4574,In_593,In_165);
or U4575 (N_4575,In_809,In_393);
nand U4576 (N_4576,In_59,In_316);
or U4577 (N_4577,In_41,In_986);
nor U4578 (N_4578,In_118,In_354);
and U4579 (N_4579,In_225,In_927);
nor U4580 (N_4580,In_651,In_67);
nand U4581 (N_4581,In_355,In_449);
or U4582 (N_4582,In_173,In_512);
and U4583 (N_4583,In_582,In_227);
and U4584 (N_4584,In_296,In_140);
or U4585 (N_4585,In_520,In_959);
nand U4586 (N_4586,In_741,In_457);
or U4587 (N_4587,In_354,In_279);
nand U4588 (N_4588,In_406,In_110);
and U4589 (N_4589,In_669,In_418);
and U4590 (N_4590,In_181,In_188);
or U4591 (N_4591,In_618,In_490);
nand U4592 (N_4592,In_197,In_906);
and U4593 (N_4593,In_754,In_746);
or U4594 (N_4594,In_316,In_478);
and U4595 (N_4595,In_254,In_773);
or U4596 (N_4596,In_584,In_490);
nand U4597 (N_4597,In_456,In_962);
nand U4598 (N_4598,In_494,In_529);
or U4599 (N_4599,In_664,In_289);
or U4600 (N_4600,In_944,In_303);
nand U4601 (N_4601,In_540,In_167);
nor U4602 (N_4602,In_625,In_267);
nand U4603 (N_4603,In_801,In_614);
nor U4604 (N_4604,In_693,In_743);
and U4605 (N_4605,In_117,In_596);
nand U4606 (N_4606,In_563,In_370);
or U4607 (N_4607,In_573,In_24);
and U4608 (N_4608,In_461,In_319);
or U4609 (N_4609,In_895,In_983);
and U4610 (N_4610,In_364,In_527);
nand U4611 (N_4611,In_522,In_304);
or U4612 (N_4612,In_719,In_41);
and U4613 (N_4613,In_476,In_892);
nor U4614 (N_4614,In_142,In_460);
and U4615 (N_4615,In_689,In_34);
and U4616 (N_4616,In_956,In_837);
and U4617 (N_4617,In_823,In_589);
nor U4618 (N_4618,In_907,In_89);
or U4619 (N_4619,In_172,In_93);
nor U4620 (N_4620,In_744,In_405);
nor U4621 (N_4621,In_319,In_318);
nand U4622 (N_4622,In_81,In_640);
or U4623 (N_4623,In_878,In_810);
nand U4624 (N_4624,In_137,In_956);
nand U4625 (N_4625,In_912,In_4);
nand U4626 (N_4626,In_611,In_555);
nand U4627 (N_4627,In_830,In_124);
and U4628 (N_4628,In_787,In_419);
nor U4629 (N_4629,In_929,In_347);
and U4630 (N_4630,In_614,In_14);
or U4631 (N_4631,In_181,In_376);
nand U4632 (N_4632,In_719,In_568);
nand U4633 (N_4633,In_289,In_149);
nor U4634 (N_4634,In_980,In_373);
or U4635 (N_4635,In_91,In_564);
or U4636 (N_4636,In_709,In_609);
nand U4637 (N_4637,In_343,In_475);
nor U4638 (N_4638,In_938,In_267);
or U4639 (N_4639,In_282,In_998);
nor U4640 (N_4640,In_584,In_675);
nor U4641 (N_4641,In_534,In_717);
or U4642 (N_4642,In_956,In_781);
nor U4643 (N_4643,In_502,In_309);
or U4644 (N_4644,In_966,In_641);
or U4645 (N_4645,In_478,In_498);
nor U4646 (N_4646,In_90,In_796);
or U4647 (N_4647,In_429,In_632);
and U4648 (N_4648,In_53,In_22);
nor U4649 (N_4649,In_756,In_575);
or U4650 (N_4650,In_730,In_846);
or U4651 (N_4651,In_179,In_452);
nand U4652 (N_4652,In_273,In_499);
nor U4653 (N_4653,In_361,In_962);
nor U4654 (N_4654,In_108,In_222);
and U4655 (N_4655,In_982,In_237);
or U4656 (N_4656,In_484,In_347);
nand U4657 (N_4657,In_907,In_476);
nor U4658 (N_4658,In_864,In_423);
nor U4659 (N_4659,In_807,In_101);
or U4660 (N_4660,In_996,In_34);
nor U4661 (N_4661,In_205,In_594);
nor U4662 (N_4662,In_437,In_365);
and U4663 (N_4663,In_752,In_380);
xnor U4664 (N_4664,In_227,In_99);
nor U4665 (N_4665,In_195,In_942);
nand U4666 (N_4666,In_236,In_191);
nor U4667 (N_4667,In_930,In_448);
or U4668 (N_4668,In_752,In_414);
and U4669 (N_4669,In_25,In_78);
nand U4670 (N_4670,In_191,In_119);
and U4671 (N_4671,In_317,In_942);
nor U4672 (N_4672,In_214,In_773);
nand U4673 (N_4673,In_669,In_590);
nor U4674 (N_4674,In_542,In_513);
nor U4675 (N_4675,In_486,In_562);
or U4676 (N_4676,In_766,In_327);
nand U4677 (N_4677,In_257,In_71);
or U4678 (N_4678,In_149,In_673);
and U4679 (N_4679,In_220,In_54);
and U4680 (N_4680,In_978,In_803);
nor U4681 (N_4681,In_993,In_504);
and U4682 (N_4682,In_249,In_525);
nor U4683 (N_4683,In_317,In_779);
nand U4684 (N_4684,In_63,In_575);
and U4685 (N_4685,In_611,In_750);
or U4686 (N_4686,In_560,In_558);
nor U4687 (N_4687,In_103,In_235);
nor U4688 (N_4688,In_144,In_768);
nand U4689 (N_4689,In_352,In_415);
nand U4690 (N_4690,In_847,In_599);
or U4691 (N_4691,In_46,In_805);
and U4692 (N_4692,In_385,In_419);
nor U4693 (N_4693,In_500,In_402);
nand U4694 (N_4694,In_944,In_804);
or U4695 (N_4695,In_612,In_4);
nand U4696 (N_4696,In_412,In_126);
nor U4697 (N_4697,In_210,In_776);
nor U4698 (N_4698,In_899,In_62);
or U4699 (N_4699,In_624,In_440);
and U4700 (N_4700,In_316,In_40);
nand U4701 (N_4701,In_103,In_680);
and U4702 (N_4702,In_913,In_699);
nand U4703 (N_4703,In_244,In_422);
nand U4704 (N_4704,In_725,In_655);
nand U4705 (N_4705,In_888,In_922);
and U4706 (N_4706,In_701,In_232);
nand U4707 (N_4707,In_591,In_34);
nor U4708 (N_4708,In_339,In_43);
nand U4709 (N_4709,In_486,In_770);
nor U4710 (N_4710,In_236,In_610);
nor U4711 (N_4711,In_519,In_189);
nand U4712 (N_4712,In_127,In_240);
nor U4713 (N_4713,In_700,In_832);
nor U4714 (N_4714,In_293,In_55);
or U4715 (N_4715,In_734,In_228);
and U4716 (N_4716,In_89,In_704);
nor U4717 (N_4717,In_513,In_169);
and U4718 (N_4718,In_231,In_977);
nor U4719 (N_4719,In_278,In_142);
and U4720 (N_4720,In_612,In_457);
nand U4721 (N_4721,In_583,In_267);
and U4722 (N_4722,In_258,In_274);
and U4723 (N_4723,In_701,In_556);
nand U4724 (N_4724,In_172,In_632);
nand U4725 (N_4725,In_818,In_95);
nand U4726 (N_4726,In_694,In_975);
nor U4727 (N_4727,In_771,In_565);
and U4728 (N_4728,In_873,In_741);
nor U4729 (N_4729,In_49,In_473);
nand U4730 (N_4730,In_518,In_64);
or U4731 (N_4731,In_705,In_239);
nor U4732 (N_4732,In_242,In_513);
nand U4733 (N_4733,In_113,In_197);
nor U4734 (N_4734,In_687,In_620);
or U4735 (N_4735,In_125,In_127);
or U4736 (N_4736,In_946,In_729);
nand U4737 (N_4737,In_134,In_711);
or U4738 (N_4738,In_824,In_251);
nor U4739 (N_4739,In_585,In_151);
nor U4740 (N_4740,In_351,In_660);
and U4741 (N_4741,In_573,In_687);
nand U4742 (N_4742,In_213,In_379);
nor U4743 (N_4743,In_751,In_798);
or U4744 (N_4744,In_98,In_191);
nor U4745 (N_4745,In_968,In_860);
nor U4746 (N_4746,In_264,In_69);
nor U4747 (N_4747,In_600,In_7);
nand U4748 (N_4748,In_997,In_287);
xnor U4749 (N_4749,In_997,In_804);
nor U4750 (N_4750,In_264,In_210);
and U4751 (N_4751,In_82,In_438);
nor U4752 (N_4752,In_134,In_179);
and U4753 (N_4753,In_105,In_368);
nand U4754 (N_4754,In_440,In_438);
nor U4755 (N_4755,In_30,In_302);
nand U4756 (N_4756,In_497,In_81);
nand U4757 (N_4757,In_895,In_157);
nor U4758 (N_4758,In_370,In_797);
nand U4759 (N_4759,In_147,In_125);
nor U4760 (N_4760,In_975,In_726);
nor U4761 (N_4761,In_350,In_965);
nand U4762 (N_4762,In_477,In_431);
or U4763 (N_4763,In_250,In_450);
nand U4764 (N_4764,In_74,In_471);
and U4765 (N_4765,In_253,In_342);
or U4766 (N_4766,In_323,In_318);
nor U4767 (N_4767,In_22,In_806);
nor U4768 (N_4768,In_835,In_199);
and U4769 (N_4769,In_410,In_676);
and U4770 (N_4770,In_374,In_910);
and U4771 (N_4771,In_647,In_658);
or U4772 (N_4772,In_939,In_846);
or U4773 (N_4773,In_107,In_352);
or U4774 (N_4774,In_647,In_634);
or U4775 (N_4775,In_853,In_413);
or U4776 (N_4776,In_293,In_100);
nand U4777 (N_4777,In_596,In_968);
or U4778 (N_4778,In_605,In_519);
nor U4779 (N_4779,In_445,In_191);
nor U4780 (N_4780,In_352,In_351);
or U4781 (N_4781,In_537,In_436);
nand U4782 (N_4782,In_15,In_428);
nor U4783 (N_4783,In_210,In_718);
or U4784 (N_4784,In_753,In_387);
nor U4785 (N_4785,In_671,In_32);
or U4786 (N_4786,In_259,In_603);
nand U4787 (N_4787,In_848,In_934);
nor U4788 (N_4788,In_4,In_120);
nor U4789 (N_4789,In_490,In_899);
nand U4790 (N_4790,In_429,In_0);
nor U4791 (N_4791,In_941,In_62);
nor U4792 (N_4792,In_904,In_581);
nor U4793 (N_4793,In_377,In_458);
or U4794 (N_4794,In_408,In_451);
nand U4795 (N_4795,In_687,In_713);
or U4796 (N_4796,In_278,In_238);
or U4797 (N_4797,In_117,In_342);
nand U4798 (N_4798,In_152,In_648);
or U4799 (N_4799,In_870,In_488);
xor U4800 (N_4800,In_329,In_43);
and U4801 (N_4801,In_678,In_643);
and U4802 (N_4802,In_975,In_192);
nor U4803 (N_4803,In_623,In_807);
nor U4804 (N_4804,In_847,In_386);
or U4805 (N_4805,In_746,In_125);
nand U4806 (N_4806,In_659,In_541);
and U4807 (N_4807,In_503,In_508);
or U4808 (N_4808,In_577,In_9);
or U4809 (N_4809,In_794,In_40);
and U4810 (N_4810,In_735,In_756);
or U4811 (N_4811,In_32,In_269);
and U4812 (N_4812,In_510,In_569);
or U4813 (N_4813,In_253,In_412);
nor U4814 (N_4814,In_354,In_21);
and U4815 (N_4815,In_450,In_872);
nand U4816 (N_4816,In_546,In_151);
nor U4817 (N_4817,In_611,In_751);
and U4818 (N_4818,In_320,In_350);
or U4819 (N_4819,In_498,In_884);
and U4820 (N_4820,In_692,In_966);
and U4821 (N_4821,In_801,In_997);
or U4822 (N_4822,In_983,In_698);
nand U4823 (N_4823,In_605,In_35);
or U4824 (N_4824,In_896,In_291);
nor U4825 (N_4825,In_491,In_738);
and U4826 (N_4826,In_94,In_269);
and U4827 (N_4827,In_911,In_320);
nor U4828 (N_4828,In_961,In_890);
nor U4829 (N_4829,In_145,In_726);
nand U4830 (N_4830,In_680,In_204);
and U4831 (N_4831,In_330,In_317);
nand U4832 (N_4832,In_960,In_538);
or U4833 (N_4833,In_317,In_676);
nand U4834 (N_4834,In_65,In_771);
or U4835 (N_4835,In_807,In_134);
nor U4836 (N_4836,In_258,In_592);
nand U4837 (N_4837,In_62,In_708);
nor U4838 (N_4838,In_238,In_730);
or U4839 (N_4839,In_853,In_589);
and U4840 (N_4840,In_836,In_23);
nand U4841 (N_4841,In_378,In_692);
or U4842 (N_4842,In_311,In_738);
nand U4843 (N_4843,In_484,In_659);
and U4844 (N_4844,In_66,In_292);
and U4845 (N_4845,In_815,In_40);
or U4846 (N_4846,In_838,In_298);
or U4847 (N_4847,In_469,In_340);
nor U4848 (N_4848,In_948,In_20);
or U4849 (N_4849,In_348,In_51);
and U4850 (N_4850,In_68,In_629);
or U4851 (N_4851,In_760,In_481);
xnor U4852 (N_4852,In_210,In_392);
nand U4853 (N_4853,In_481,In_85);
nand U4854 (N_4854,In_687,In_379);
nand U4855 (N_4855,In_114,In_502);
xor U4856 (N_4856,In_335,In_400);
and U4857 (N_4857,In_237,In_497);
nor U4858 (N_4858,In_891,In_162);
or U4859 (N_4859,In_695,In_771);
and U4860 (N_4860,In_60,In_493);
nand U4861 (N_4861,In_268,In_637);
nand U4862 (N_4862,In_453,In_928);
and U4863 (N_4863,In_536,In_894);
or U4864 (N_4864,In_972,In_567);
xnor U4865 (N_4865,In_237,In_814);
or U4866 (N_4866,In_600,In_939);
nor U4867 (N_4867,In_379,In_592);
nor U4868 (N_4868,In_947,In_650);
nor U4869 (N_4869,In_594,In_924);
nor U4870 (N_4870,In_173,In_983);
or U4871 (N_4871,In_85,In_183);
and U4872 (N_4872,In_226,In_704);
or U4873 (N_4873,In_433,In_690);
nand U4874 (N_4874,In_215,In_627);
and U4875 (N_4875,In_595,In_904);
nand U4876 (N_4876,In_488,In_657);
or U4877 (N_4877,In_800,In_211);
nand U4878 (N_4878,In_325,In_770);
nor U4879 (N_4879,In_372,In_844);
and U4880 (N_4880,In_587,In_825);
or U4881 (N_4881,In_141,In_616);
nor U4882 (N_4882,In_790,In_83);
nand U4883 (N_4883,In_797,In_14);
or U4884 (N_4884,In_658,In_957);
and U4885 (N_4885,In_159,In_134);
or U4886 (N_4886,In_283,In_787);
nand U4887 (N_4887,In_948,In_915);
nor U4888 (N_4888,In_54,In_451);
and U4889 (N_4889,In_455,In_558);
and U4890 (N_4890,In_904,In_900);
or U4891 (N_4891,In_27,In_951);
or U4892 (N_4892,In_344,In_253);
nand U4893 (N_4893,In_673,In_400);
and U4894 (N_4894,In_784,In_261);
nor U4895 (N_4895,In_145,In_88);
nand U4896 (N_4896,In_333,In_507);
nand U4897 (N_4897,In_641,In_67);
or U4898 (N_4898,In_604,In_901);
and U4899 (N_4899,In_576,In_877);
or U4900 (N_4900,In_641,In_771);
nor U4901 (N_4901,In_59,In_673);
and U4902 (N_4902,In_831,In_800);
nand U4903 (N_4903,In_334,In_12);
and U4904 (N_4904,In_753,In_886);
and U4905 (N_4905,In_583,In_108);
nand U4906 (N_4906,In_736,In_352);
and U4907 (N_4907,In_391,In_977);
and U4908 (N_4908,In_807,In_227);
nand U4909 (N_4909,In_202,In_80);
or U4910 (N_4910,In_339,In_134);
and U4911 (N_4911,In_779,In_62);
nor U4912 (N_4912,In_993,In_100);
nand U4913 (N_4913,In_158,In_674);
nor U4914 (N_4914,In_547,In_902);
nor U4915 (N_4915,In_64,In_305);
or U4916 (N_4916,In_494,In_957);
nor U4917 (N_4917,In_481,In_458);
nand U4918 (N_4918,In_93,In_964);
or U4919 (N_4919,In_949,In_536);
nor U4920 (N_4920,In_970,In_664);
or U4921 (N_4921,In_911,In_702);
nor U4922 (N_4922,In_560,In_452);
or U4923 (N_4923,In_98,In_963);
nor U4924 (N_4924,In_358,In_992);
nand U4925 (N_4925,In_584,In_451);
or U4926 (N_4926,In_80,In_855);
xor U4927 (N_4927,In_471,In_810);
or U4928 (N_4928,In_935,In_56);
nand U4929 (N_4929,In_430,In_315);
and U4930 (N_4930,In_575,In_210);
nand U4931 (N_4931,In_378,In_830);
or U4932 (N_4932,In_104,In_683);
nor U4933 (N_4933,In_513,In_159);
nand U4934 (N_4934,In_300,In_523);
or U4935 (N_4935,In_653,In_876);
nor U4936 (N_4936,In_251,In_550);
or U4937 (N_4937,In_632,In_167);
or U4938 (N_4938,In_8,In_66);
or U4939 (N_4939,In_983,In_46);
nor U4940 (N_4940,In_38,In_35);
or U4941 (N_4941,In_579,In_203);
or U4942 (N_4942,In_271,In_671);
nor U4943 (N_4943,In_140,In_324);
nor U4944 (N_4944,In_506,In_452);
nand U4945 (N_4945,In_513,In_691);
or U4946 (N_4946,In_932,In_706);
nor U4947 (N_4947,In_955,In_566);
and U4948 (N_4948,In_768,In_235);
or U4949 (N_4949,In_49,In_833);
xnor U4950 (N_4950,In_318,In_340);
or U4951 (N_4951,In_355,In_543);
nand U4952 (N_4952,In_322,In_125);
nor U4953 (N_4953,In_437,In_530);
nand U4954 (N_4954,In_430,In_863);
and U4955 (N_4955,In_8,In_249);
nor U4956 (N_4956,In_48,In_146);
nand U4957 (N_4957,In_416,In_996);
or U4958 (N_4958,In_655,In_562);
or U4959 (N_4959,In_844,In_1);
nand U4960 (N_4960,In_532,In_327);
nand U4961 (N_4961,In_443,In_656);
nand U4962 (N_4962,In_842,In_277);
nand U4963 (N_4963,In_827,In_525);
nor U4964 (N_4964,In_15,In_314);
nand U4965 (N_4965,In_616,In_692);
or U4966 (N_4966,In_819,In_992);
or U4967 (N_4967,In_96,In_108);
nand U4968 (N_4968,In_835,In_10);
nor U4969 (N_4969,In_760,In_656);
nor U4970 (N_4970,In_909,In_80);
nand U4971 (N_4971,In_885,In_3);
nor U4972 (N_4972,In_933,In_222);
nor U4973 (N_4973,In_613,In_253);
and U4974 (N_4974,In_685,In_931);
nand U4975 (N_4975,In_407,In_175);
and U4976 (N_4976,In_230,In_75);
nand U4977 (N_4977,In_178,In_519);
nand U4978 (N_4978,In_1,In_507);
and U4979 (N_4979,In_22,In_804);
and U4980 (N_4980,In_63,In_12);
or U4981 (N_4981,In_549,In_830);
nor U4982 (N_4982,In_296,In_673);
or U4983 (N_4983,In_438,In_545);
or U4984 (N_4984,In_353,In_891);
xnor U4985 (N_4985,In_170,In_581);
and U4986 (N_4986,In_643,In_185);
and U4987 (N_4987,In_663,In_66);
or U4988 (N_4988,In_528,In_95);
nor U4989 (N_4989,In_666,In_586);
nand U4990 (N_4990,In_12,In_594);
and U4991 (N_4991,In_610,In_840);
or U4992 (N_4992,In_850,In_168);
nand U4993 (N_4993,In_887,In_509);
and U4994 (N_4994,In_879,In_928);
or U4995 (N_4995,In_109,In_884);
nand U4996 (N_4996,In_796,In_643);
and U4997 (N_4997,In_807,In_216);
nor U4998 (N_4998,In_235,In_370);
or U4999 (N_4999,In_592,In_881);
nor U5000 (N_5000,N_1020,N_2120);
or U5001 (N_5001,N_4374,N_2345);
nor U5002 (N_5002,N_151,N_2103);
and U5003 (N_5003,N_3689,N_1065);
nand U5004 (N_5004,N_263,N_2157);
and U5005 (N_5005,N_3350,N_3398);
and U5006 (N_5006,N_45,N_599);
and U5007 (N_5007,N_4688,N_1660);
nand U5008 (N_5008,N_4272,N_4657);
xor U5009 (N_5009,N_3354,N_2156);
nand U5010 (N_5010,N_870,N_2375);
or U5011 (N_5011,N_4140,N_3209);
nand U5012 (N_5012,N_3942,N_1176);
or U5013 (N_5013,N_4427,N_4426);
or U5014 (N_5014,N_2264,N_4292);
nor U5015 (N_5015,N_4932,N_1721);
nand U5016 (N_5016,N_1758,N_3248);
nand U5017 (N_5017,N_4060,N_1729);
nand U5018 (N_5018,N_4455,N_714);
nor U5019 (N_5019,N_1671,N_969);
or U5020 (N_5020,N_2234,N_3871);
and U5021 (N_5021,N_594,N_1338);
nand U5022 (N_5022,N_1172,N_4569);
nor U5023 (N_5023,N_29,N_3904);
nor U5024 (N_5024,N_3466,N_4852);
nand U5025 (N_5025,N_4953,N_2782);
or U5026 (N_5026,N_15,N_4127);
nand U5027 (N_5027,N_32,N_1099);
nor U5028 (N_5028,N_3539,N_2384);
and U5029 (N_5029,N_603,N_4122);
nand U5030 (N_5030,N_2024,N_785);
nand U5031 (N_5031,N_1770,N_3719);
xnor U5032 (N_5032,N_2818,N_563);
nand U5033 (N_5033,N_2618,N_4760);
nand U5034 (N_5034,N_4447,N_3771);
or U5035 (N_5035,N_2277,N_3302);
nor U5036 (N_5036,N_3017,N_1279);
or U5037 (N_5037,N_2140,N_4612);
nor U5038 (N_5038,N_1627,N_3512);
or U5039 (N_5039,N_25,N_4303);
nand U5040 (N_5040,N_1732,N_135);
or U5041 (N_5041,N_848,N_1173);
or U5042 (N_5042,N_1522,N_1268);
nor U5043 (N_5043,N_4049,N_4897);
or U5044 (N_5044,N_4345,N_381);
nor U5045 (N_5045,N_2305,N_4836);
nand U5046 (N_5046,N_4962,N_4989);
nor U5047 (N_5047,N_139,N_422);
and U5048 (N_5048,N_2418,N_1854);
and U5049 (N_5049,N_2703,N_1407);
nand U5050 (N_5050,N_1037,N_3450);
nand U5051 (N_5051,N_1736,N_1511);
nand U5052 (N_5052,N_2280,N_3985);
or U5053 (N_5053,N_4386,N_4848);
nand U5054 (N_5054,N_4914,N_1587);
and U5055 (N_5055,N_2047,N_1067);
nand U5056 (N_5056,N_2398,N_1723);
or U5057 (N_5057,N_4238,N_1015);
and U5058 (N_5058,N_1963,N_4246);
nand U5059 (N_5059,N_1615,N_3821);
nand U5060 (N_5060,N_4767,N_4279);
nand U5061 (N_5061,N_4458,N_1210);
and U5062 (N_5062,N_1321,N_4838);
and U5063 (N_5063,N_4369,N_956);
xnor U5064 (N_5064,N_4092,N_1490);
or U5065 (N_5065,N_3419,N_162);
nand U5066 (N_5066,N_4438,N_4300);
and U5067 (N_5067,N_470,N_1967);
and U5068 (N_5068,N_2530,N_4142);
and U5069 (N_5069,N_1394,N_4687);
nor U5070 (N_5070,N_3929,N_4739);
and U5071 (N_5071,N_3016,N_4547);
and U5072 (N_5072,N_2975,N_4436);
and U5073 (N_5073,N_1492,N_52);
and U5074 (N_5074,N_1678,N_817);
nand U5075 (N_5075,N_1055,N_2983);
nand U5076 (N_5076,N_4772,N_886);
nand U5077 (N_5077,N_1433,N_878);
nor U5078 (N_5078,N_2516,N_3632);
nor U5079 (N_5079,N_3170,N_31);
and U5080 (N_5080,N_3988,N_4437);
and U5081 (N_5081,N_2141,N_3358);
and U5082 (N_5082,N_2665,N_2393);
or U5083 (N_5083,N_3702,N_2396);
and U5084 (N_5084,N_1102,N_4580);
nand U5085 (N_5085,N_4890,N_690);
nor U5086 (N_5086,N_3515,N_4723);
or U5087 (N_5087,N_106,N_4245);
nand U5088 (N_5088,N_857,N_2945);
nand U5089 (N_5089,N_3649,N_637);
nand U5090 (N_5090,N_1423,N_3437);
or U5091 (N_5091,N_3744,N_3353);
nor U5092 (N_5092,N_342,N_97);
or U5093 (N_5093,N_18,N_4108);
nor U5094 (N_5094,N_1884,N_1366);
and U5095 (N_5095,N_4529,N_3662);
and U5096 (N_5096,N_2736,N_3543);
nor U5097 (N_5097,N_503,N_4994);
nand U5098 (N_5098,N_4229,N_4656);
and U5099 (N_5099,N_4750,N_1186);
or U5100 (N_5100,N_1160,N_331);
and U5101 (N_5101,N_1273,N_323);
nor U5102 (N_5102,N_3734,N_3714);
and U5103 (N_5103,N_4576,N_695);
nor U5104 (N_5104,N_3725,N_99);
and U5105 (N_5105,N_1529,N_4783);
and U5106 (N_5106,N_3535,N_2315);
or U5107 (N_5107,N_2642,N_625);
or U5108 (N_5108,N_1710,N_4343);
or U5109 (N_5109,N_2682,N_2121);
nor U5110 (N_5110,N_3410,N_4434);
nand U5111 (N_5111,N_767,N_3080);
nor U5112 (N_5112,N_3157,N_209);
nor U5113 (N_5113,N_3884,N_2136);
or U5114 (N_5114,N_88,N_4482);
and U5115 (N_5115,N_2771,N_2143);
and U5116 (N_5116,N_2399,N_204);
nor U5117 (N_5117,N_3105,N_2940);
or U5118 (N_5118,N_4075,N_2804);
nor U5119 (N_5119,N_4907,N_92);
nand U5120 (N_5120,N_4693,N_2297);
or U5121 (N_5121,N_825,N_474);
nor U5122 (N_5122,N_4441,N_3832);
and U5123 (N_5123,N_838,N_726);
nor U5124 (N_5124,N_961,N_4360);
nand U5125 (N_5125,N_3798,N_2791);
nor U5126 (N_5126,N_4544,N_1969);
or U5127 (N_5127,N_1914,N_1759);
nand U5128 (N_5128,N_1701,N_4083);
nand U5129 (N_5129,N_3004,N_3723);
nand U5130 (N_5130,N_1794,N_3745);
nand U5131 (N_5131,N_4814,N_4942);
nor U5132 (N_5132,N_2144,N_2509);
nor U5133 (N_5133,N_4534,N_1140);
or U5134 (N_5134,N_3562,N_1124);
nor U5135 (N_5135,N_2973,N_1110);
nor U5136 (N_5136,N_163,N_1591);
or U5137 (N_5137,N_1760,N_3160);
nor U5138 (N_5138,N_3200,N_2481);
nor U5139 (N_5139,N_4596,N_4645);
and U5140 (N_5140,N_3309,N_1088);
or U5141 (N_5141,N_1436,N_3506);
or U5142 (N_5142,N_1948,N_4530);
or U5143 (N_5143,N_3197,N_1127);
nor U5144 (N_5144,N_286,N_2584);
nor U5145 (N_5145,N_2592,N_3769);
nand U5146 (N_5146,N_4100,N_2355);
nor U5147 (N_5147,N_3447,N_2927);
or U5148 (N_5148,N_868,N_1157);
xnor U5149 (N_5149,N_3322,N_3328);
or U5150 (N_5150,N_3005,N_4834);
and U5151 (N_5151,N_4433,N_2366);
or U5152 (N_5152,N_1636,N_5);
nor U5153 (N_5153,N_1456,N_2574);
nor U5154 (N_5154,N_639,N_4863);
or U5155 (N_5155,N_4764,N_2414);
and U5156 (N_5156,N_2358,N_3807);
nand U5157 (N_5157,N_3012,N_2891);
nand U5158 (N_5158,N_3083,N_4940);
or U5159 (N_5159,N_3387,N_2201);
nand U5160 (N_5160,N_4188,N_680);
and U5161 (N_5161,N_2337,N_1445);
and U5162 (N_5162,N_4562,N_2200);
nand U5163 (N_5163,N_1457,N_2555);
nor U5164 (N_5164,N_2554,N_4903);
nand U5165 (N_5165,N_4102,N_2360);
and U5166 (N_5166,N_1304,N_986);
nor U5167 (N_5167,N_2562,N_3079);
nand U5168 (N_5168,N_653,N_627);
and U5169 (N_5169,N_1296,N_4929);
nand U5170 (N_5170,N_2594,N_433);
or U5171 (N_5171,N_4881,N_3971);
and U5172 (N_5172,N_1161,N_4790);
nand U5173 (N_5173,N_1850,N_662);
nand U5174 (N_5174,N_1198,N_1968);
and U5175 (N_5175,N_1586,N_4079);
and U5176 (N_5176,N_4261,N_1889);
or U5177 (N_5177,N_909,N_3351);
and U5178 (N_5178,N_861,N_1043);
nand U5179 (N_5179,N_1653,N_1670);
and U5180 (N_5180,N_757,N_4996);
and U5181 (N_5181,N_673,N_3169);
or U5182 (N_5182,N_2836,N_176);
or U5183 (N_5183,N_755,N_2857);
or U5184 (N_5184,N_4061,N_435);
nor U5185 (N_5185,N_1887,N_1530);
nand U5186 (N_5186,N_4672,N_4780);
nand U5187 (N_5187,N_1558,N_1285);
and U5188 (N_5188,N_2893,N_4243);
nor U5189 (N_5189,N_3476,N_3068);
and U5190 (N_5190,N_4009,N_391);
or U5191 (N_5191,N_4330,N_207);
nor U5192 (N_5192,N_3448,N_2388);
and U5193 (N_5193,N_4701,N_3009);
or U5194 (N_5194,N_421,N_1917);
and U5195 (N_5195,N_3499,N_4682);
and U5196 (N_5196,N_3425,N_265);
and U5197 (N_5197,N_4763,N_3203);
nor U5198 (N_5198,N_569,N_2332);
or U5199 (N_5199,N_1897,N_1345);
nand U5200 (N_5200,N_3810,N_562);
nor U5201 (N_5201,N_2069,N_4904);
or U5202 (N_5202,N_2578,N_508);
nand U5203 (N_5203,N_3164,N_4133);
or U5204 (N_5204,N_480,N_4307);
nor U5205 (N_5205,N_2934,N_4706);
or U5206 (N_5206,N_1957,N_3824);
or U5207 (N_5207,N_763,N_137);
and U5208 (N_5208,N_4889,N_1773);
nor U5209 (N_5209,N_4404,N_2988);
and U5210 (N_5210,N_2013,N_4543);
and U5211 (N_5211,N_3802,N_1420);
or U5212 (N_5212,N_4844,N_1931);
or U5213 (N_5213,N_4632,N_2435);
and U5214 (N_5214,N_3845,N_3869);
nor U5215 (N_5215,N_3758,N_3071);
nand U5216 (N_5216,N_3603,N_1021);
nand U5217 (N_5217,N_1940,N_3031);
nor U5218 (N_5218,N_4414,N_1898);
or U5219 (N_5219,N_1488,N_3308);
nor U5220 (N_5220,N_2513,N_2247);
or U5221 (N_5221,N_2646,N_1720);
nor U5222 (N_5222,N_1668,N_892);
nand U5223 (N_5223,N_1594,N_363);
or U5224 (N_5224,N_3396,N_2668);
nand U5225 (N_5225,N_2276,N_1471);
nor U5226 (N_5226,N_1482,N_3850);
nor U5227 (N_5227,N_1971,N_4479);
nand U5228 (N_5228,N_947,N_4028);
nor U5229 (N_5229,N_78,N_4538);
nand U5230 (N_5230,N_3040,N_285);
and U5231 (N_5231,N_3381,N_2050);
nor U5232 (N_5232,N_4765,N_1498);
nand U5233 (N_5233,N_1106,N_2735);
nor U5234 (N_5234,N_1076,N_4905);
nand U5235 (N_5235,N_3705,N_1430);
nor U5236 (N_5236,N_4830,N_195);
nand U5237 (N_5237,N_4804,N_1754);
nand U5238 (N_5238,N_2401,N_1374);
nor U5239 (N_5239,N_169,N_2801);
or U5240 (N_5240,N_4705,N_4798);
nor U5241 (N_5241,N_2471,N_4990);
or U5242 (N_5242,N_2607,N_1191);
nand U5243 (N_5243,N_1978,N_461);
nand U5244 (N_5244,N_4112,N_4743);
nor U5245 (N_5245,N_2174,N_416);
or U5246 (N_5246,N_874,N_3388);
or U5247 (N_5247,N_4356,N_2601);
and U5248 (N_5248,N_3885,N_2128);
nor U5249 (N_5249,N_4240,N_107);
nor U5250 (N_5250,N_397,N_3670);
nand U5251 (N_5251,N_4016,N_2627);
nor U5252 (N_5252,N_3347,N_548);
nor U5253 (N_5253,N_398,N_1614);
or U5254 (N_5254,N_2636,N_555);
or U5255 (N_5255,N_394,N_2429);
nor U5256 (N_5256,N_4314,N_3436);
and U5257 (N_5257,N_999,N_1427);
and U5258 (N_5258,N_2158,N_3464);
nand U5259 (N_5259,N_1112,N_3795);
and U5260 (N_5260,N_2210,N_4638);
or U5261 (N_5261,N_4203,N_4741);
nand U5262 (N_5262,N_2752,N_3013);
or U5263 (N_5263,N_2477,N_1777);
nor U5264 (N_5264,N_2076,N_3742);
or U5265 (N_5265,N_3604,N_87);
nand U5266 (N_5266,N_2135,N_3973);
and U5267 (N_5267,N_1060,N_241);
or U5268 (N_5268,N_1454,N_4690);
nand U5269 (N_5269,N_621,N_3362);
and U5270 (N_5270,N_4726,N_2869);
and U5271 (N_5271,N_1918,N_2840);
or U5272 (N_5272,N_4503,N_3107);
or U5273 (N_5273,N_3806,N_898);
or U5274 (N_5274,N_2595,N_3356);
xnor U5275 (N_5275,N_3747,N_2541);
nor U5276 (N_5276,N_4017,N_3010);
and U5277 (N_5277,N_4317,N_993);
nor U5278 (N_5278,N_4526,N_759);
xor U5279 (N_5279,N_1937,N_1063);
and U5280 (N_5280,N_2048,N_738);
nor U5281 (N_5281,N_2591,N_3591);
nand U5282 (N_5282,N_3680,N_980);
and U5283 (N_5283,N_1453,N_1905);
and U5284 (N_5284,N_4802,N_2908);
nand U5285 (N_5285,N_4887,N_1237);
and U5286 (N_5286,N_1410,N_3323);
or U5287 (N_5287,N_64,N_3324);
and U5288 (N_5288,N_4024,N_379);
nand U5289 (N_5289,N_2218,N_4459);
nand U5290 (N_5290,N_4190,N_2998);
nand U5291 (N_5291,N_4435,N_4954);
nand U5292 (N_5292,N_2783,N_498);
nor U5293 (N_5293,N_1271,N_1838);
and U5294 (N_5294,N_2968,N_3111);
or U5295 (N_5295,N_3483,N_834);
or U5296 (N_5296,N_2299,N_3945);
or U5297 (N_5297,N_1380,N_120);
nand U5298 (N_5298,N_2670,N_3870);
nor U5299 (N_5299,N_452,N_1925);
and U5300 (N_5300,N_3380,N_3274);
nor U5301 (N_5301,N_1399,N_4560);
and U5302 (N_5302,N_4147,N_3421);
nor U5303 (N_5303,N_2316,N_349);
or U5304 (N_5304,N_650,N_1483);
nor U5305 (N_5305,N_1799,N_4922);
or U5306 (N_5306,N_2550,N_1510);
or U5307 (N_5307,N_2630,N_4185);
or U5308 (N_5308,N_370,N_310);
and U5309 (N_5309,N_1942,N_3600);
nand U5310 (N_5310,N_2311,N_4875);
and U5311 (N_5311,N_2767,N_1531);
and U5312 (N_5312,N_4058,N_4336);
and U5313 (N_5313,N_3774,N_688);
nor U5314 (N_5314,N_2291,N_3902);
and U5315 (N_5315,N_1182,N_4368);
nor U5316 (N_5316,N_2197,N_114);
or U5317 (N_5317,N_4952,N_890);
xnor U5318 (N_5318,N_3379,N_4231);
nand U5319 (N_5319,N_4902,N_3936);
nor U5320 (N_5320,N_2362,N_2613);
nor U5321 (N_5321,N_4388,N_3831);
nor U5322 (N_5322,N_227,N_3921);
nand U5323 (N_5323,N_3136,N_1601);
nand U5324 (N_5324,N_2520,N_4398);
and U5325 (N_5325,N_4618,N_4719);
nor U5326 (N_5326,N_3053,N_4335);
nor U5327 (N_5327,N_184,N_155);
or U5328 (N_5328,N_2118,N_4679);
nor U5329 (N_5329,N_710,N_749);
or U5330 (N_5330,N_4807,N_2495);
nor U5331 (N_5331,N_3580,N_876);
and U5332 (N_5332,N_560,N_495);
or U5333 (N_5333,N_1752,N_847);
or U5334 (N_5334,N_589,N_2223);
nand U5335 (N_5335,N_4327,N_4465);
or U5336 (N_5336,N_3553,N_2486);
and U5337 (N_5337,N_2647,N_2923);
and U5338 (N_5338,N_2307,N_3428);
nor U5339 (N_5339,N_4648,N_3960);
nor U5340 (N_5340,N_1334,N_1416);
or U5341 (N_5341,N_2078,N_3837);
and U5342 (N_5342,N_3234,N_3249);
nand U5343 (N_5343,N_3946,N_1373);
nor U5344 (N_5344,N_459,N_4756);
nand U5345 (N_5345,N_1090,N_4019);
nor U5346 (N_5346,N_3541,N_1691);
nor U5347 (N_5347,N_2074,N_68);
nor U5348 (N_5348,N_4787,N_238);
nor U5349 (N_5349,N_995,N_2907);
nor U5350 (N_5350,N_794,N_2597);
nand U5351 (N_5351,N_3932,N_190);
and U5352 (N_5352,N_3687,N_3363);
nor U5353 (N_5353,N_2057,N_375);
nand U5354 (N_5354,N_368,N_1502);
or U5355 (N_5355,N_3494,N_4866);
and U5356 (N_5356,N_2845,N_3517);
nor U5357 (N_5357,N_2610,N_3633);
nand U5358 (N_5358,N_2081,N_2717);
nand U5359 (N_5359,N_2428,N_1346);
or U5360 (N_5360,N_558,N_4253);
and U5361 (N_5361,N_3441,N_697);
or U5362 (N_5362,N_4715,N_1461);
xnor U5363 (N_5363,N_214,N_4077);
and U5364 (N_5364,N_2914,N_4766);
or U5365 (N_5365,N_1936,N_3269);
or U5366 (N_5366,N_2890,N_1542);
nand U5367 (N_5367,N_4110,N_2371);
nor U5368 (N_5368,N_4288,N_3311);
or U5369 (N_5369,N_3015,N_3895);
and U5370 (N_5370,N_3839,N_808);
and U5371 (N_5371,N_4971,N_4540);
nand U5372 (N_5372,N_3305,N_1728);
and U5373 (N_5373,N_2871,N_1733);
nand U5374 (N_5374,N_2391,N_3424);
or U5375 (N_5375,N_329,N_671);
nand U5376 (N_5376,N_2547,N_3968);
nor U5377 (N_5377,N_3475,N_2750);
nand U5378 (N_5378,N_4789,N_1158);
nand U5379 (N_5379,N_2424,N_4702);
nand U5380 (N_5380,N_4341,N_1867);
or U5381 (N_5381,N_2522,N_1938);
or U5382 (N_5382,N_4453,N_473);
nand U5383 (N_5383,N_3147,N_515);
or U5384 (N_5384,N_193,N_1223);
or U5385 (N_5385,N_4030,N_339);
and U5386 (N_5386,N_2267,N_2850);
and U5387 (N_5387,N_577,N_4520);
nor U5388 (N_5388,N_3051,N_1113);
nand U5389 (N_5389,N_1707,N_1569);
and U5390 (N_5390,N_2901,N_2667);
nor U5391 (N_5391,N_1362,N_822);
or U5392 (N_5392,N_2108,N_1387);
nor U5393 (N_5393,N_1893,N_1537);
and U5394 (N_5394,N_1094,N_113);
nand U5395 (N_5395,N_1797,N_1050);
and U5396 (N_5396,N_4043,N_1214);
and U5397 (N_5397,N_1452,N_4877);
and U5398 (N_5398,N_3630,N_1330);
xnor U5399 (N_5399,N_651,N_1421);
or U5400 (N_5400,N_1254,N_4865);
nand U5401 (N_5401,N_4389,N_2814);
and U5402 (N_5402,N_4457,N_1805);
nand U5403 (N_5403,N_1676,N_4759);
nor U5404 (N_5404,N_4072,N_4210);
nand U5405 (N_5405,N_2748,N_4412);
nor U5406 (N_5406,N_4949,N_1910);
or U5407 (N_5407,N_2385,N_4869);
and U5408 (N_5408,N_2022,N_741);
nand U5409 (N_5409,N_922,N_63);
and U5410 (N_5410,N_3913,N_3155);
nor U5411 (N_5411,N_1538,N_2702);
or U5412 (N_5412,N_968,N_1351);
and U5413 (N_5413,N_1982,N_3935);
xnor U5414 (N_5414,N_3052,N_4938);
nand U5415 (N_5415,N_3551,N_3438);
or U5416 (N_5416,N_4349,N_4306);
nand U5417 (N_5417,N_1293,N_4358);
nor U5418 (N_5418,N_4299,N_35);
or U5419 (N_5419,N_3726,N_3596);
and U5420 (N_5420,N_682,N_1316);
or U5421 (N_5421,N_1166,N_91);
and U5422 (N_5422,N_833,N_4716);
or U5423 (N_5423,N_1183,N_4284);
nand U5424 (N_5424,N_1751,N_2811);
and U5425 (N_5425,N_4208,N_4069);
nor U5426 (N_5426,N_4555,N_1882);
or U5427 (N_5427,N_1269,N_4753);
and U5428 (N_5428,N_771,N_1169);
nand U5429 (N_5429,N_1204,N_1170);
and U5430 (N_5430,N_2700,N_3455);
nor U5431 (N_5431,N_333,N_4101);
or U5432 (N_5432,N_2018,N_2444);
and U5433 (N_5433,N_2408,N_2443);
nand U5434 (N_5434,N_2454,N_3178);
and U5435 (N_5435,N_483,N_3877);
nor U5436 (N_5436,N_543,N_2160);
nand U5437 (N_5437,N_3916,N_842);
and U5438 (N_5438,N_2965,N_4496);
nor U5439 (N_5439,N_4597,N_2580);
and U5440 (N_5440,N_1540,N_2483);
or U5441 (N_5441,N_1054,N_2905);
or U5442 (N_5442,N_1403,N_3020);
nand U5443 (N_5443,N_1702,N_3360);
and U5444 (N_5444,N_1181,N_2870);
nand U5445 (N_5445,N_2942,N_889);
nand U5446 (N_5446,N_1425,N_437);
nand U5447 (N_5447,N_1038,N_1988);
nand U5448 (N_5448,N_1029,N_3153);
or U5449 (N_5449,N_2777,N_552);
or U5450 (N_5450,N_2394,N_2230);
or U5451 (N_5451,N_2616,N_2012);
or U5452 (N_5452,N_4181,N_4067);
nor U5453 (N_5453,N_4329,N_3648);
nand U5454 (N_5454,N_239,N_739);
xnor U5455 (N_5455,N_2786,N_1946);
nor U5456 (N_5456,N_4423,N_213);
or U5457 (N_5457,N_1294,N_668);
and U5458 (N_5458,N_3752,N_4390);
or U5459 (N_5459,N_4563,N_494);
nand U5460 (N_5460,N_1605,N_3498);
or U5461 (N_5461,N_4777,N_378);
nand U5462 (N_5462,N_3149,N_602);
nor U5463 (N_5463,N_3874,N_4167);
nand U5464 (N_5464,N_429,N_3526);
or U5465 (N_5465,N_358,N_937);
nor U5466 (N_5466,N_4213,N_1699);
xor U5467 (N_5467,N_1953,N_3749);
or U5468 (N_5468,N_4403,N_643);
nand U5469 (N_5469,N_1286,N_2809);
and U5470 (N_5470,N_4833,N_4146);
and U5471 (N_5471,N_1132,N_351);
nor U5472 (N_5472,N_2663,N_3781);
or U5473 (N_5473,N_4888,N_2656);
nor U5474 (N_5474,N_3531,N_1414);
or U5475 (N_5475,N_2812,N_962);
or U5476 (N_5476,N_262,N_1137);
or U5477 (N_5477,N_325,N_615);
nor U5478 (N_5478,N_2301,N_2154);
nor U5479 (N_5479,N_1667,N_3629);
or U5480 (N_5480,N_4500,N_887);
nor U5481 (N_5481,N_2575,N_2284);
nor U5482 (N_5482,N_4411,N_3467);
nand U5483 (N_5483,N_1566,N_3355);
or U5484 (N_5484,N_1785,N_1836);
nand U5485 (N_5485,N_4405,N_3899);
nand U5486 (N_5486,N_3631,N_4258);
nor U5487 (N_5487,N_1541,N_2115);
and U5488 (N_5488,N_4254,N_72);
and U5489 (N_5489,N_2802,N_2586);
nor U5490 (N_5490,N_3325,N_4915);
and U5491 (N_5491,N_1300,N_2623);
nor U5492 (N_5492,N_1926,N_3727);
or U5493 (N_5493,N_2505,N_2961);
and U5494 (N_5494,N_4218,N_1692);
xor U5495 (N_5495,N_1952,N_3784);
and U5496 (N_5496,N_3740,N_4373);
nor U5497 (N_5497,N_2126,N_4786);
or U5498 (N_5498,N_1283,N_2402);
nor U5499 (N_5499,N_3431,N_3433);
nor U5500 (N_5500,N_4007,N_4960);
nand U5501 (N_5501,N_1044,N_530);
nand U5502 (N_5502,N_2031,N_4986);
and U5503 (N_5503,N_413,N_872);
nand U5504 (N_5504,N_115,N_604);
nand U5505 (N_5505,N_3857,N_1449);
and U5506 (N_5506,N_1257,N_4152);
nand U5507 (N_5507,N_3418,N_3693);
or U5508 (N_5508,N_950,N_989);
and U5509 (N_5509,N_4132,N_4571);
nand U5510 (N_5510,N_2219,N_3417);
nand U5511 (N_5511,N_2084,N_3847);
nand U5512 (N_5512,N_4085,N_894);
nand U5513 (N_5513,N_3247,N_3375);
nor U5514 (N_5514,N_1326,N_4471);
and U5515 (N_5515,N_3284,N_2635);
or U5516 (N_5516,N_4955,N_3691);
or U5517 (N_5517,N_1508,N_705);
nor U5518 (N_5518,N_2040,N_1155);
and U5519 (N_5519,N_4602,N_24);
or U5520 (N_5520,N_1229,N_531);
or U5521 (N_5521,N_4531,N_3442);
nand U5522 (N_5522,N_4084,N_4326);
nor U5523 (N_5523,N_1100,N_1983);
and U5524 (N_5524,N_1767,N_2014);
nor U5525 (N_5525,N_3926,N_1539);
nand U5526 (N_5526,N_4975,N_891);
or U5527 (N_5527,N_2744,N_939);
or U5528 (N_5528,N_1830,N_2149);
nand U5529 (N_5529,N_985,N_3289);
nand U5530 (N_5530,N_4733,N_2238);
nor U5531 (N_5531,N_2270,N_1557);
or U5532 (N_5532,N_0,N_4059);
and U5533 (N_5533,N_1645,N_2847);
nand U5534 (N_5534,N_4985,N_2242);
nand U5535 (N_5535,N_2123,N_1860);
and U5536 (N_5536,N_1298,N_3150);
nor U5537 (N_5537,N_1772,N_4197);
and U5538 (N_5538,N_2930,N_983);
nand U5539 (N_5539,N_1381,N_2758);
or U5540 (N_5540,N_1793,N_2631);
and U5541 (N_5541,N_4809,N_2041);
nor U5542 (N_5542,N_3801,N_1116);
or U5543 (N_5543,N_837,N_318);
nand U5544 (N_5544,N_4451,N_852);
and U5545 (N_5545,N_1136,N_4583);
nor U5546 (N_5546,N_1547,N_2922);
nor U5547 (N_5547,N_1255,N_2387);
nand U5548 (N_5548,N_3788,N_1574);
nor U5549 (N_5549,N_4277,N_337);
nand U5550 (N_5550,N_3905,N_716);
nand U5551 (N_5551,N_4365,N_2348);
and U5552 (N_5552,N_1307,N_1363);
and U5553 (N_5553,N_3341,N_524);
or U5554 (N_5554,N_3563,N_1842);
and U5555 (N_5555,N_3779,N_4799);
and U5556 (N_5556,N_1190,N_4921);
or U5557 (N_5557,N_3659,N_3711);
nand U5558 (N_5558,N_4988,N_2763);
nand U5559 (N_5559,N_2926,N_2484);
nor U5560 (N_5560,N_405,N_1074);
nand U5561 (N_5561,N_4627,N_875);
nand U5562 (N_5562,N_4510,N_3909);
and U5563 (N_5563,N_3304,N_645);
and U5564 (N_5564,N_4755,N_1618);
nor U5565 (N_5565,N_3695,N_3637);
nor U5566 (N_5566,N_4681,N_1187);
and U5567 (N_5567,N_3549,N_997);
nor U5568 (N_5568,N_3759,N_2021);
nor U5569 (N_5569,N_824,N_287);
nand U5570 (N_5570,N_3148,N_79);
nor U5571 (N_5571,N_526,N_4784);
or U5572 (N_5572,N_2917,N_4778);
nor U5573 (N_5573,N_4609,N_3622);
or U5574 (N_5574,N_1159,N_3663);
nor U5575 (N_5575,N_4042,N_250);
and U5576 (N_5576,N_2312,N_4125);
nand U5577 (N_5577,N_4397,N_1369);
nand U5578 (N_5578,N_3962,N_4517);
and U5579 (N_5579,N_4150,N_2848);
nand U5580 (N_5580,N_2641,N_841);
nor U5581 (N_5581,N_2220,N_3470);
and U5582 (N_5582,N_2864,N_4965);
nor U5583 (N_5583,N_44,N_167);
and U5584 (N_5584,N_344,N_3523);
or U5585 (N_5585,N_41,N_1985);
or U5586 (N_5586,N_4832,N_3678);
and U5587 (N_5587,N_918,N_1189);
or U5588 (N_5588,N_1841,N_1520);
and U5589 (N_5589,N_1372,N_929);
nor U5590 (N_5590,N_3041,N_3595);
or U5591 (N_5591,N_1990,N_2339);
xnor U5592 (N_5592,N_4325,N_3420);
and U5593 (N_5593,N_353,N_4585);
nor U5594 (N_5594,N_3684,N_4823);
nand U5595 (N_5595,N_1310,N_3236);
and U5596 (N_5596,N_466,N_967);
or U5597 (N_5597,N_4293,N_3540);
or U5598 (N_5598,N_3422,N_1075);
nor U5599 (N_5599,N_4925,N_4029);
nand U5600 (N_5600,N_3995,N_2209);
nand U5601 (N_5601,N_4383,N_393);
nor U5602 (N_5602,N_367,N_3703);
and U5603 (N_5603,N_4376,N_2617);
nand U5604 (N_5604,N_4663,N_1516);
or U5605 (N_5605,N_2473,N_4183);
nand U5606 (N_5606,N_3273,N_259);
nand U5607 (N_5607,N_172,N_856);
nor U5608 (N_5608,N_410,N_2094);
nand U5609 (N_5609,N_2405,N_3760);
nand U5610 (N_5610,N_2564,N_4039);
nand U5611 (N_5611,N_2976,N_1322);
nand U5612 (N_5612,N_2379,N_3919);
nand U5613 (N_5613,N_4725,N_3235);
and U5614 (N_5614,N_2560,N_3565);
or U5615 (N_5615,N_815,N_254);
nand U5616 (N_5616,N_1727,N_2981);
nor U5617 (N_5617,N_3014,N_991);
nor U5618 (N_5618,N_2889,N_2807);
and U5619 (N_5619,N_1146,N_3461);
and U5620 (N_5620,N_2993,N_4281);
nor U5621 (N_5621,N_895,N_1129);
xor U5622 (N_5622,N_1804,N_2446);
or U5623 (N_5623,N_1779,N_3212);
nor U5624 (N_5624,N_4499,N_341);
nand U5625 (N_5625,N_4984,N_1536);
nor U5626 (N_5626,N_2828,N_521);
nand U5627 (N_5627,N_4420,N_39);
nand U5628 (N_5628,N_4677,N_4614);
or U5629 (N_5629,N_3141,N_4346);
nand U5630 (N_5630,N_4164,N_1979);
nand U5631 (N_5631,N_3792,N_3577);
nand U5632 (N_5632,N_4773,N_3616);
nor U5633 (N_5633,N_90,N_1703);
and U5634 (N_5634,N_4347,N_4919);
or U5635 (N_5635,N_3953,N_1650);
and U5636 (N_5636,N_2637,N_826);
or U5637 (N_5637,N_1486,N_3975);
xor U5638 (N_5638,N_3757,N_146);
and U5639 (N_5639,N_4126,N_2704);
and U5640 (N_5640,N_3271,N_4651);
nor U5641 (N_5641,N_3260,N_3521);
xor U5642 (N_5642,N_4315,N_361);
and U5643 (N_5643,N_1481,N_1504);
nand U5644 (N_5644,N_3836,N_126);
nand U5645 (N_5645,N_2304,N_1426);
nor U5646 (N_5646,N_2390,N_3701);
and U5647 (N_5647,N_3963,N_1588);
nor U5648 (N_5648,N_355,N_3830);
and U5649 (N_5649,N_2886,N_2112);
or U5650 (N_5650,N_3074,N_4533);
nor U5651 (N_5651,N_2415,N_3028);
nand U5652 (N_5652,N_4828,N_2372);
or U5653 (N_5653,N_1045,N_4797);
nor U5654 (N_5654,N_522,N_4394);
or U5655 (N_5655,N_1117,N_3189);
nand U5656 (N_5656,N_4806,N_201);
and U5657 (N_5657,N_2127,N_990);
nor U5658 (N_5658,N_3280,N_2579);
and U5659 (N_5659,N_4273,N_1774);
or U5660 (N_5660,N_1422,N_1658);
nor U5661 (N_5661,N_3947,N_2898);
nand U5662 (N_5662,N_1750,N_1911);
or U5663 (N_5663,N_2456,N_4035);
and U5664 (N_5664,N_4913,N_3961);
and U5665 (N_5665,N_2778,N_1222);
nand U5666 (N_5666,N_4066,N_3025);
nand U5667 (N_5667,N_1994,N_654);
nor U5668 (N_5668,N_1951,N_931);
nor U5669 (N_5669,N_2448,N_3849);
nor U5670 (N_5670,N_1619,N_2824);
nand U5671 (N_5671,N_4579,N_2107);
and U5672 (N_5672,N_4769,N_1518);
or U5673 (N_5673,N_2897,N_1999);
and U5674 (N_5674,N_1485,N_655);
nand U5675 (N_5675,N_3664,N_684);
and U5676 (N_5676,N_1207,N_2491);
nor U5677 (N_5677,N_2919,N_4744);
or U5678 (N_5678,N_4257,N_202);
nor U5679 (N_5679,N_4324,N_1388);
and U5680 (N_5680,N_2195,N_4056);
or U5681 (N_5681,N_2971,N_1009);
and U5682 (N_5682,N_3775,N_1525);
or U5683 (N_5683,N_4232,N_3712);
or U5684 (N_5684,N_3881,N_4709);
or U5685 (N_5685,N_3854,N_893);
nor U5686 (N_5686,N_127,N_4055);
nand U5687 (N_5687,N_3454,N_3065);
nand U5688 (N_5688,N_4582,N_636);
or U5689 (N_5689,N_622,N_831);
and U5690 (N_5690,N_4136,N_4355);
nor U5691 (N_5691,N_3805,N_462);
nor U5692 (N_5692,N_4372,N_2410);
or U5693 (N_5693,N_2990,N_3718);
or U5694 (N_5694,N_3762,N_2878);
nor U5695 (N_5695,N_3883,N_2492);
or U5696 (N_5696,N_619,N_4977);
nor U5697 (N_5697,N_1496,N_2088);
and U5698 (N_5698,N_1135,N_3797);
or U5699 (N_5699,N_4660,N_2208);
nor U5700 (N_5700,N_3930,N_4361);
nand U5701 (N_5701,N_4721,N_4931);
and U5702 (N_5702,N_2461,N_2055);
or U5703 (N_5703,N_324,N_3627);
nor U5704 (N_5704,N_3699,N_1103);
or U5705 (N_5705,N_3282,N_2873);
and U5706 (N_5706,N_4217,N_1034);
nor U5707 (N_5707,N_192,N_715);
or U5708 (N_5708,N_4170,N_2518);
nor U5709 (N_5709,N_3529,N_4973);
nor U5710 (N_5710,N_4595,N_2543);
nor U5711 (N_5711,N_920,N_408);
xnor U5712 (N_5712,N_4377,N_3538);
and U5713 (N_5713,N_2761,N_4608);
or U5714 (N_5714,N_326,N_3113);
or U5715 (N_5715,N_3660,N_4393);
nand U5716 (N_5716,N_1499,N_1107);
and U5717 (N_5717,N_4930,N_516);
or U5718 (N_5718,N_3034,N_3463);
nor U5719 (N_5719,N_2723,N_4666);
and U5720 (N_5720,N_2581,N_2900);
nor U5721 (N_5721,N_67,N_1956);
nor U5722 (N_5722,N_490,N_3011);
nor U5723 (N_5723,N_3495,N_4957);
nor U5724 (N_5724,N_2322,N_3796);
or U5725 (N_5725,N_27,N_449);
and U5726 (N_5726,N_4312,N_2254);
nand U5727 (N_5727,N_2148,N_587);
or U5728 (N_5728,N_3043,N_1347);
xnor U5729 (N_5729,N_496,N_211);
and U5730 (N_5730,N_1628,N_3102);
and U5731 (N_5731,N_1756,N_2915);
nor U5732 (N_5732,N_701,N_3263);
nor U5733 (N_5733,N_4737,N_2510);
and U5734 (N_5734,N_2314,N_4086);
nor U5735 (N_5735,N_2892,N_1258);
and U5736 (N_5736,N_2985,N_2259);
or U5737 (N_5737,N_2517,N_751);
and U5738 (N_5738,N_3096,N_4626);
and U5739 (N_5739,N_553,N_4617);
nor U5740 (N_5740,N_4570,N_1562);
or U5741 (N_5741,N_4839,N_3270);
nor U5742 (N_5742,N_4621,N_3791);
and U5743 (N_5743,N_2773,N_2369);
nand U5744 (N_5744,N_2251,N_147);
nand U5745 (N_5745,N_383,N_4850);
nand U5746 (N_5746,N_3704,N_4811);
and U5747 (N_5747,N_423,N_4255);
and U5748 (N_5748,N_2680,N_1309);
or U5749 (N_5749,N_2110,N_3602);
nand U5750 (N_5750,N_3307,N_2295);
nand U5751 (N_5751,N_4600,N_607);
and U5752 (N_5752,N_4856,N_536);
and U5753 (N_5753,N_3608,N_3359);
or U5754 (N_5754,N_3569,N_1833);
nand U5755 (N_5755,N_4249,N_3250);
and U5756 (N_5756,N_2754,N_1813);
nor U5757 (N_5757,N_578,N_1960);
nand U5758 (N_5758,N_58,N_4144);
nor U5759 (N_5759,N_2794,N_196);
xnor U5760 (N_5760,N_3116,N_1661);
and U5761 (N_5761,N_1317,N_1644);
and U5762 (N_5762,N_468,N_4022);
nor U5763 (N_5763,N_1150,N_1795);
or U5764 (N_5764,N_3578,N_4542);
and U5765 (N_5765,N_4053,N_3124);
and U5766 (N_5766,N_647,N_532);
nor U5767 (N_5767,N_2052,N_1944);
or U5768 (N_5768,N_240,N_1339);
nand U5769 (N_5769,N_3044,N_3315);
and U5770 (N_5770,N_4948,N_4918);
nor U5771 (N_5771,N_3572,N_3951);
nor U5772 (N_5772,N_2300,N_3611);
nand U5773 (N_5773,N_295,N_457);
nand U5774 (N_5774,N_1580,N_2470);
and U5775 (N_5775,N_4171,N_1709);
nor U5776 (N_5776,N_1320,N_4174);
and U5777 (N_5777,N_4124,N_693);
and U5778 (N_5778,N_4539,N_4976);
nand U5779 (N_5779,N_3860,N_2317);
nand U5780 (N_5780,N_185,N_4031);
nand U5781 (N_5781,N_2895,N_3685);
nor U5782 (N_5782,N_3756,N_1262);
and U5783 (N_5783,N_1122,N_1684);
or U5784 (N_5784,N_440,N_1178);
nor U5785 (N_5785,N_95,N_2831);
or U5786 (N_5786,N_2095,N_4639);
or U5787 (N_5787,N_4810,N_3330);
and U5788 (N_5788,N_2779,N_2512);
and U5789 (N_5789,N_1472,N_2309);
nand U5790 (N_5790,N_3844,N_289);
nand U5791 (N_5791,N_3165,N_3692);
or U5792 (N_5792,N_4207,N_1371);
nor U5793 (N_5793,N_4549,N_3440);
and U5794 (N_5794,N_158,N_3337);
or U5795 (N_5795,N_4586,N_3897);
or U5796 (N_5796,N_3038,N_404);
nor U5797 (N_5797,N_4179,N_2035);
nand U5798 (N_5798,N_2732,N_4815);
nand U5799 (N_5799,N_1115,N_4551);
nand U5800 (N_5800,N_3898,N_601);
or U5801 (N_5801,N_3676,N_631);
and U5802 (N_5802,N_232,N_3334);
or U5803 (N_5803,N_3265,N_3502);
and U5804 (N_5804,N_2913,N_4934);
and U5805 (N_5805,N_2916,N_3059);
or U5806 (N_5806,N_305,N_3661);
nor U5807 (N_5807,N_3114,N_3528);
nor U5808 (N_5808,N_2933,N_1809);
or U5809 (N_5809,N_3872,N_915);
or U5810 (N_5810,N_1869,N_4532);
nor U5811 (N_5811,N_879,N_4912);
xor U5812 (N_5812,N_2827,N_4634);
and U5813 (N_5813,N_761,N_4096);
nor U5814 (N_5814,N_3667,N_2738);
and U5815 (N_5815,N_1843,N_835);
nor U5816 (N_5816,N_4259,N_1290);
and U5817 (N_5817,N_1806,N_853);
nand U5818 (N_5818,N_276,N_3518);
nor U5819 (N_5819,N_858,N_4490);
and U5820 (N_5820,N_2911,N_2876);
nor U5821 (N_5821,N_3119,N_2793);
or U5822 (N_5822,N_1031,N_948);
nand U5823 (N_5823,N_4649,N_609);
and U5824 (N_5824,N_1359,N_3076);
or U5825 (N_5825,N_3343,N_1154);
xor U5826 (N_5826,N_4993,N_1177);
and U5827 (N_5827,N_3135,N_3790);
nand U5828 (N_5828,N_2774,N_1206);
and U5829 (N_5829,N_624,N_2507);
nand U5830 (N_5830,N_829,N_4872);
or U5831 (N_5831,N_1782,N_3384);
and U5832 (N_5832,N_3199,N_2175);
nor U5833 (N_5833,N_3026,N_4409);
nand U5834 (N_5834,N_606,N_3266);
nand U5835 (N_5835,N_3889,N_1348);
or U5836 (N_5836,N_1688,N_2053);
nor U5837 (N_5837,N_4812,N_261);
nor U5838 (N_5838,N_528,N_1224);
nor U5839 (N_5839,N_3713,N_86);
and U5840 (N_5840,N_1941,N_2169);
nor U5841 (N_5841,N_3613,N_3144);
nor U5842 (N_5842,N_2268,N_66);
or U5843 (N_5843,N_3003,N_3842);
or U5844 (N_5844,N_3378,N_3996);
and U5845 (N_5845,N_1977,N_1396);
nor U5846 (N_5846,N_839,N_685);
or U5847 (N_5847,N_1677,N_3903);
or U5848 (N_5848,N_2370,N_3510);
or U5849 (N_5849,N_1,N_2569);
or U5850 (N_5850,N_4071,N_2183);
nand U5851 (N_5851,N_2743,N_1716);
nor U5852 (N_5852,N_2097,N_4244);
nand U5853 (N_5853,N_813,N_401);
or U5854 (N_5854,N_2970,N_380);
nor U5855 (N_5855,N_3918,N_1442);
nor U5856 (N_5856,N_2003,N_1517);
or U5857 (N_5857,N_4094,N_1631);
and U5858 (N_5858,N_1778,N_1563);
nand U5859 (N_5859,N_4521,N_3777);
nand U5860 (N_5860,N_377,N_1718);
or U5861 (N_5861,N_1883,N_236);
or U5862 (N_5862,N_2902,N_2086);
and U5863 (N_5863,N_1635,N_3207);
and U5864 (N_5864,N_523,N_3992);
or U5865 (N_5865,N_467,N_694);
nor U5866 (N_5866,N_2296,N_4751);
or U5867 (N_5867,N_4221,N_133);
nor U5868 (N_5868,N_1662,N_2687);
nor U5869 (N_5869,N_4105,N_247);
nor U5870 (N_5870,N_2180,N_1881);
nor U5871 (N_5871,N_3880,N_3027);
nor U5872 (N_5872,N_3556,N_2669);
and U5873 (N_5873,N_3827,N_2237);
nor U5874 (N_5874,N_4481,N_2679);
or U5875 (N_5875,N_420,N_492);
nor U5876 (N_5876,N_1199,N_4633);
nor U5877 (N_5877,N_2005,N_796);
nand U5878 (N_5878,N_3598,N_683);
and U5879 (N_5879,N_764,N_2521);
nor U5880 (N_5880,N_2328,N_1891);
nor U5881 (N_5881,N_4200,N_865);
and U5882 (N_5882,N_2324,N_3614);
and U5883 (N_5883,N_3125,N_884);
or U5884 (N_5884,N_3977,N_3901);
and U5885 (N_5885,N_3293,N_4186);
and U5886 (N_5886,N_1284,N_458);
nor U5887 (N_5887,N_3524,N_2426);
nor U5888 (N_5888,N_2712,N_215);
or U5889 (N_5889,N_4223,N_3671);
nand U5890 (N_5890,N_789,N_4091);
or U5891 (N_5891,N_460,N_1260);
and U5892 (N_5892,N_4054,N_4270);
nand U5893 (N_5893,N_4002,N_3650);
and U5894 (N_5894,N_3644,N_108);
nand U5895 (N_5895,N_664,N_2787);
nor U5896 (N_5896,N_3570,N_1437);
nor U5897 (N_5897,N_1451,N_1282);
and U5898 (N_5898,N_1392,N_4241);
nand U5899 (N_5899,N_4320,N_731);
nor U5900 (N_5900,N_1266,N_4023);
nor U5901 (N_5901,N_3145,N_657);
nand U5902 (N_5902,N_4518,N_3679);
and U5903 (N_5903,N_2912,N_1082);
or U5904 (N_5904,N_4015,N_4738);
and U5905 (N_5905,N_1391,N_1477);
or U5906 (N_5906,N_4868,N_4310);
or U5907 (N_5907,N_2034,N_199);
and U5908 (N_5908,N_4524,N_721);
and U5909 (N_5909,N_400,N_1203);
or U5910 (N_5910,N_2666,N_53);
and U5911 (N_5911,N_4637,N_3835);
nand U5912 (N_5912,N_4008,N_3999);
and U5913 (N_5913,N_3340,N_1570);
nor U5914 (N_5914,N_2285,N_220);
and U5915 (N_5915,N_119,N_3227);
or U5916 (N_5916,N_3046,N_575);
nor U5917 (N_5917,N_489,N_2186);
nor U5918 (N_5918,N_1665,N_4422);
nor U5919 (N_5919,N_125,N_3423);
nand U5920 (N_5920,N_4757,N_1855);
nand U5921 (N_5921,N_1332,N_50);
or U5922 (N_5922,N_3937,N_3765);
or U5923 (N_5923,N_596,N_2956);
and U5924 (N_5924,N_1197,N_546);
and U5925 (N_5925,N_610,N_1487);
nand U5926 (N_5926,N_3944,N_4339);
nor U5927 (N_5927,N_1019,N_1324);
nand U5928 (N_5928,N_248,N_4044);
nor U5929 (N_5929,N_4474,N_559);
or U5930 (N_5930,N_3914,N_226);
or U5931 (N_5931,N_4062,N_55);
nand U5932 (N_5932,N_745,N_2765);
nor U5933 (N_5933,N_1996,N_2308);
or U5934 (N_5934,N_1340,N_4646);
nor U5935 (N_5935,N_1787,N_4722);
nand U5936 (N_5936,N_2286,N_899);
nor U5937 (N_5937,N_581,N_2017);
nor U5938 (N_5938,N_4088,N_1353);
or U5939 (N_5939,N_1997,N_4078);
or U5940 (N_5940,N_1895,N_669);
or U5941 (N_5941,N_2760,N_3675);
nand U5942 (N_5942,N_4808,N_2929);
nand U5943 (N_5943,N_2533,N_2137);
and U5944 (N_5944,N_4076,N_83);
nand U5945 (N_5945,N_4662,N_445);
and U5946 (N_5946,N_1418,N_3743);
or U5947 (N_5947,N_3093,N_1724);
or U5948 (N_5948,N_1965,N_2515);
and U5949 (N_5949,N_965,N_3060);
nand U5950 (N_5950,N_2966,N_479);
nand U5951 (N_5951,N_1377,N_4419);
nor U5952 (N_5952,N_2114,N_497);
nor U5953 (N_5953,N_2457,N_3585);
nor U5954 (N_5954,N_1680,N_2867);
and U5955 (N_5955,N_2480,N_2000);
or U5956 (N_5956,N_3439,N_3369);
nor U5957 (N_5957,N_4138,N_1617);
nor U5958 (N_5958,N_2272,N_3943);
nand U5959 (N_5959,N_1311,N_2239);
and U5960 (N_5960,N_3032,N_4309);
nor U5961 (N_5961,N_3176,N_4717);
and U5962 (N_5962,N_4762,N_2351);
nor U5963 (N_5963,N_3268,N_512);
or U5964 (N_5964,N_2619,N_3391);
nor U5965 (N_5965,N_4642,N_4981);
or U5966 (N_5966,N_1598,N_1448);
or U5967 (N_5967,N_3576,N_2462);
nor U5968 (N_5968,N_1848,N_660);
nand U5969 (N_5969,N_1270,N_3112);
nor U5970 (N_5970,N_1098,N_3115);
nor U5971 (N_5971,N_2422,N_4224);
nand U5972 (N_5972,N_3816,N_3245);
and U5973 (N_5973,N_1892,N_4923);
nand U5974 (N_5974,N_3414,N_3925);
or U5975 (N_5975,N_1171,N_1383);
nor U5976 (N_5976,N_205,N_81);
nor U5977 (N_5977,N_4048,N_798);
and U5978 (N_5978,N_3101,N_2859);
nand U5979 (N_5979,N_1633,N_4697);
or U5980 (N_5980,N_988,N_2083);
nand U5981 (N_5981,N_455,N_1125);
and U5982 (N_5982,N_3401,N_3216);
nand U5983 (N_5983,N_1220,N_3156);
or U5984 (N_5984,N_3139,N_1781);
nand U5985 (N_5985,N_4822,N_869);
and U5986 (N_5986,N_3232,N_2488);
and U5987 (N_5987,N_1250,N_3416);
nand U5988 (N_5988,N_2746,N_2742);
nor U5989 (N_5989,N_2184,N_200);
nand U5990 (N_5990,N_4817,N_3333);
and U5991 (N_5991,N_1468,N_4280);
and U5992 (N_5992,N_40,N_4871);
nor U5993 (N_5993,N_1046,N_1080);
xor U5994 (N_5994,N_597,N_2032);
or U5995 (N_5995,N_3297,N_1613);
nand U5996 (N_5996,N_1640,N_4943);
or U5997 (N_5997,N_3786,N_2525);
nor U5998 (N_5998,N_1863,N_4406);
or U5999 (N_5999,N_4916,N_385);
or U6000 (N_6000,N_633,N_529);
and U6001 (N_6001,N_387,N_1981);
nand U6002 (N_6002,N_3707,N_2256);
or U6003 (N_6003,N_1059,N_3778);
nor U6004 (N_6004,N_2060,N_2250);
nand U6005 (N_6005,N_2553,N_281);
and U6006 (N_6006,N_1634,N_271);
nand U6007 (N_6007,N_382,N_4120);
and U6008 (N_6008,N_4109,N_60);
and U6009 (N_6009,N_2951,N_3301);
nand U6010 (N_6010,N_4689,N_1864);
nor U6011 (N_6011,N_3829,N_2701);
and U6012 (N_6012,N_1556,N_1244);
and U6013 (N_6013,N_1467,N_3761);
nor U6014 (N_6014,N_47,N_1213);
nand U6015 (N_6015,N_691,N_1976);
and U6016 (N_6016,N_4640,N_4963);
or U6017 (N_6017,N_2936,N_4215);
and U6018 (N_6018,N_1603,N_3504);
nand U6019 (N_6019,N_3403,N_1337);
and U6020 (N_6020,N_568,N_1144);
and U6021 (N_6021,N_2288,N_3406);
nand U6022 (N_6022,N_2978,N_65);
xor U6023 (N_6023,N_3090,N_2066);
nor U6024 (N_6024,N_1526,N_912);
nor U6025 (N_6025,N_4430,N_540);
nand U6026 (N_6026,N_3407,N_4643);
and U6027 (N_6027,N_4969,N_327);
or U6028 (N_6028,N_1240,N_1577);
nand U6029 (N_6029,N_2856,N_1505);
nor U6030 (N_6030,N_4992,N_2188);
or U6031 (N_6031,N_2576,N_1011);
or U6032 (N_6032,N_2652,N_3690);
or U6033 (N_6033,N_1474,N_1010);
nor U6034 (N_6034,N_98,N_156);
nand U6035 (N_6035,N_2099,N_2839);
nand U6036 (N_6036,N_1934,N_2731);
and U6037 (N_6037,N_4130,N_3137);
or U6038 (N_6038,N_1185,N_4564);
or U6039 (N_6039,N_4610,N_1675);
xnor U6040 (N_6040,N_1991,N_2546);
nand U6041 (N_6041,N_2960,N_3110);
nor U6042 (N_6042,N_2633,N_1784);
or U6043 (N_6043,N_981,N_2645);
or U6044 (N_6044,N_3720,N_4578);
or U6045 (N_6045,N_3182,N_4380);
nor U6046 (N_6046,N_2894,N_2755);
and U6047 (N_6047,N_3952,N_3738);
nand U6048 (N_6048,N_316,N_4311);
nand U6049 (N_6049,N_3415,N_2502);
nor U6050 (N_6050,N_187,N_811);
nor U6051 (N_6051,N_1023,N_565);
nand U6052 (N_6052,N_3706,N_2883);
and U6053 (N_6053,N_3099,N_3606);
nor U6054 (N_6054,N_1989,N_1834);
or U6055 (N_6055,N_712,N_116);
nand U6056 (N_6056,N_1101,N_2567);
nand U6057 (N_6057,N_1145,N_4712);
and U6058 (N_6058,N_4899,N_4286);
and U6059 (N_6059,N_2189,N_2948);
nand U6060 (N_6060,N_1245,N_949);
nand U6061 (N_6061,N_1783,N_4502);
nand U6062 (N_6062,N_3130,N_2117);
nor U6063 (N_6063,N_778,N_941);
nor U6064 (N_6064,N_1673,N_4858);
or U6065 (N_6065,N_2987,N_396);
or U6066 (N_6066,N_130,N_3365);
nor U6067 (N_6067,N_33,N_1022);
or U6068 (N_6068,N_3258,N_978);
nor U6069 (N_6069,N_2329,N_2672);
or U6070 (N_6070,N_2784,N_1832);
nor U6071 (N_6071,N_4851,N_2815);
and U6072 (N_6072,N_3318,N_827);
nand U6073 (N_6073,N_4352,N_1165);
and U6074 (N_6074,N_3492,N_1695);
and U6075 (N_6075,N_260,N_1295);
nor U6076 (N_6076,N_56,N_3728);
nor U6077 (N_6077,N_4298,N_676);
nand U6078 (N_6078,N_554,N_3451);
nor U6079 (N_6079,N_1578,N_1450);
nor U6080 (N_6080,N_544,N_2173);
nor U6081 (N_6081,N_3819,N_1666);
nor U6082 (N_6082,N_1444,N_2622);
or U6083 (N_6083,N_3037,N_4468);
nor U6084 (N_6084,N_3033,N_3185);
or U6085 (N_6085,N_4089,N_788);
or U6086 (N_6086,N_1327,N_4978);
or U6087 (N_6087,N_4445,N_206);
or U6088 (N_6088,N_352,N_348);
nor U6089 (N_6089,N_2352,N_1429);
or U6090 (N_6090,N_3838,N_1315);
and U6091 (N_6091,N_2155,N_3218);
nand U6092 (N_6092,N_2092,N_4967);
nand U6093 (N_6093,N_3296,N_1501);
nand U6094 (N_6094,N_2837,N_3049);
nand U6095 (N_6095,N_4493,N_4334);
nor U6096 (N_6096,N_933,N_104);
nor U6097 (N_6097,N_74,N_4081);
and U6098 (N_6098,N_4615,N_1851);
and U6099 (N_6099,N_1233,N_1281);
nor U6100 (N_6100,N_1620,N_2153);
nor U6101 (N_6101,N_101,N_4883);
nand U6102 (N_6102,N_1071,N_3412);
and U6103 (N_6103,N_777,N_2102);
nand U6104 (N_6104,N_987,N_472);
or U6105 (N_6105,N_2689,N_830);
and U6106 (N_6106,N_3581,N_2969);
or U6107 (N_6107,N_4425,N_3453);
or U6108 (N_6108,N_1364,N_3395);
xnor U6109 (N_6109,N_1600,N_4581);
and U6110 (N_6110,N_4641,N_1534);
nor U6111 (N_6111,N_4671,N_1972);
or U6112 (N_6112,N_3709,N_572);
or U6113 (N_6113,N_1013,N_818);
nor U6114 (N_6114,N_786,N_3174);
or U6115 (N_6115,N_237,N_3997);
nand U6116 (N_6116,N_4699,N_2938);
nor U6117 (N_6117,N_3782,N_3729);
or U6118 (N_6118,N_436,N_2695);
and U6119 (N_6119,N_820,N_2659);
or U6120 (N_6120,N_1943,N_1331);
nor U6121 (N_6121,N_1859,N_4093);
nand U6122 (N_6122,N_453,N_124);
xnor U6123 (N_6123,N_4745,N_219);
and U6124 (N_6124,N_1217,N_2101);
and U6125 (N_6125,N_3098,N_2458);
and U6126 (N_6126,N_4882,N_849);
nand U6127 (N_6127,N_2269,N_520);
nor U6128 (N_6128,N_3809,N_123);
nor U6129 (N_6129,N_2226,N_4898);
or U6130 (N_6130,N_4489,N_3490);
nor U6131 (N_6131,N_3204,N_854);
or U6132 (N_6132,N_4148,N_598);
nand U6133 (N_6133,N_4328,N_2338);
nand U6134 (N_6134,N_4461,N_274);
and U6135 (N_6135,N_364,N_4118);
or U6136 (N_6136,N_2994,N_4658);
nand U6137 (N_6137,N_1431,N_2487);
and U6138 (N_6138,N_4038,N_328);
or U6139 (N_6139,N_1479,N_234);
nand U6140 (N_6140,N_3906,N_3056);
or U6141 (N_6141,N_4065,N_666);
nor U6142 (N_6142,N_1769,N_3910);
nand U6143 (N_6143,N_1776,N_280);
or U6144 (N_6144,N_1231,N_3507);
or U6145 (N_6145,N_3405,N_293);
nor U6146 (N_6146,N_3817,N_4840);
nor U6147 (N_6147,N_3338,N_451);
and U6148 (N_6148,N_689,N_1458);
and U6149 (N_6149,N_4927,N_4819);
and U6150 (N_6150,N_4870,N_1611);
and U6151 (N_6151,N_4250,N_850);
or U6152 (N_6152,N_4587,N_487);
and U6153 (N_6153,N_2271,N_1032);
or U6154 (N_6154,N_3158,N_571);
and U6155 (N_6155,N_4824,N_1228);
nor U6156 (N_6156,N_4020,N_432);
nand U6157 (N_6157,N_4454,N_3408);
nor U6158 (N_6158,N_4282,N_2838);
nand U6159 (N_6159,N_4113,N_4525);
or U6160 (N_6160,N_952,N_3717);
nor U6161 (N_6161,N_1419,N_4342);
and U6162 (N_6162,N_3281,N_3366);
nand U6163 (N_6163,N_4333,N_4956);
nor U6164 (N_6164,N_402,N_233);
or U6165 (N_6165,N_2741,N_911);
nor U6166 (N_6166,N_4515,N_505);
or U6167 (N_6167,N_2235,N_3228);
nand U6168 (N_6168,N_1441,N_1409);
nor U6169 (N_6169,N_1036,N_1026);
nand U6170 (N_6170,N_2884,N_4686);
nor U6171 (N_6171,N_3481,N_2386);
nor U6172 (N_6172,N_1845,N_4308);
and U6173 (N_6173,N_3626,N_1630);
nand U6174 (N_6174,N_2205,N_3716);
nor U6175 (N_6175,N_38,N_3399);
and U6176 (N_6176,N_2589,N_17);
or U6177 (N_6177,N_3537,N_2718);
nand U6178 (N_6178,N_4391,N_4842);
nor U6179 (N_6179,N_3339,N_307);
nor U6180 (N_6180,N_1945,N_2528);
nand U6181 (N_6181,N_2232,N_454);
nand U6182 (N_6182,N_1253,N_925);
nor U6183 (N_6183,N_1001,N_73);
nor U6184 (N_6184,N_3489,N_4854);
and U6185 (N_6185,N_1328,N_1292);
or U6186 (N_6186,N_4477,N_2715);
nand U6187 (N_6187,N_4668,N_4768);
and U6188 (N_6188,N_4225,N_3924);
nand U6189 (N_6189,N_4385,N_2170);
and U6190 (N_6190,N_2124,N_582);
nor U6191 (N_6191,N_3240,N_2350);
nand U6192 (N_6192,N_4206,N_832);
xnor U6193 (N_6193,N_2162,N_1484);
nor U6194 (N_6194,N_1877,N_976);
or U6195 (N_6195,N_4901,N_2946);
and U6196 (N_6196,N_4700,N_3298);
and U6197 (N_6197,N_4193,N_2739);
or U6198 (N_6198,N_1693,N_3372);
or U6199 (N_6199,N_13,N_1196);
nand U6200 (N_6200,N_2751,N_2207);
nor U6201 (N_6201,N_1119,N_4129);
or U6202 (N_6202,N_1555,N_4367);
nor U6203 (N_6203,N_1480,N_2536);
nor U6204 (N_6204,N_3192,N_510);
nor U6205 (N_6205,N_132,N_282);
and U6206 (N_6206,N_3131,N_4939);
nand U6207 (N_6207,N_1935,N_4878);
nand U6208 (N_6208,N_2273,N_940);
nand U6209 (N_6209,N_4775,N_2335);
or U6210 (N_6210,N_216,N_3469);
or U6211 (N_6211,N_1962,N_1975);
or U6212 (N_6212,N_2770,N_253);
and U6213 (N_6213,N_2374,N_269);
nand U6214 (N_6214,N_1344,N_3908);
nand U6215 (N_6215,N_3064,N_1970);
and U6216 (N_6216,N_1616,N_1274);
or U6217 (N_6217,N_3091,N_2298);
nand U6218 (N_6218,N_4900,N_4006);
and U6219 (N_6219,N_2868,N_2113);
nor U6220 (N_6220,N_3993,N_4236);
or U6221 (N_6221,N_2989,N_567);
or U6222 (N_6222,N_1138,N_1734);
or U6223 (N_6223,N_4271,N_971);
and U6224 (N_6224,N_3983,N_513);
and U6225 (N_6225,N_2474,N_170);
or U6226 (N_6226,N_2628,N_2514);
or U6227 (N_6227,N_2561,N_2805);
nor U6228 (N_6228,N_4505,N_1259);
and U6229 (N_6229,N_386,N_374);
nand U6230 (N_6230,N_1514,N_1543);
and U6231 (N_6231,N_3915,N_2588);
or U6232 (N_6232,N_4268,N_257);
and U6233 (N_6233,N_3542,N_203);
nand U6234 (N_6234,N_415,N_3097);
or U6235 (N_6235,N_3175,N_3081);
nand U6236 (N_6236,N_371,N_3390);
and U6237 (N_6237,N_143,N_2125);
or U6238 (N_6238,N_2644,N_292);
and U6239 (N_6239,N_600,N_863);
or U6240 (N_6240,N_579,N_309);
or U6241 (N_6241,N_702,N_2033);
nor U6242 (N_6242,N_700,N_753);
and U6243 (N_6243,N_3948,N_2651);
or U6244 (N_6244,N_3773,N_1674);
nor U6245 (N_6245,N_3893,N_4318);
and U6246 (N_6246,N_3177,N_3023);
and U6247 (N_6247,N_4876,N_3374);
nor U6248 (N_6248,N_43,N_4348);
nor U6249 (N_6249,N_2823,N_3652);
nand U6250 (N_6250,N_343,N_3638);
or U6251 (N_6251,N_4111,N_4285);
or U6252 (N_6252,N_1932,N_2389);
nor U6253 (N_6253,N_2719,N_4653);
and U6254 (N_6254,N_1583,N_535);
nor U6255 (N_6255,N_1507,N_2442);
and U6256 (N_6256,N_4891,N_1743);
xnor U6257 (N_6257,N_2079,N_2841);
and U6258 (N_6258,N_118,N_2049);
and U6259 (N_6259,N_4886,N_3552);
or U6260 (N_6260,N_2364,N_4995);
or U6261 (N_6261,N_3826,N_3673);
or U6262 (N_6262,N_179,N_4344);
or U6263 (N_6263,N_3077,N_138);
and U6264 (N_6264,N_3462,N_2138);
nand U6265 (N_6265,N_3770,N_2548);
nor U6266 (N_6266,N_923,N_1656);
nand U6267 (N_6267,N_1402,N_801);
and U6268 (N_6268,N_843,N_4873);
nand U6269 (N_6269,N_1415,N_3303);
nor U6270 (N_6270,N_48,N_4590);
or U6271 (N_6271,N_4399,N_1698);
or U6272 (N_6272,N_59,N_1913);
nor U6273 (N_6273,N_1700,N_1406);
nand U6274 (N_6274,N_4983,N_2445);
or U6275 (N_6275,N_2164,N_963);
nor U6276 (N_6276,N_3750,N_1024);
or U6277 (N_6277,N_20,N_2059);
nor U6278 (N_6278,N_3558,N_3892);
and U6279 (N_6279,N_3519,N_2626);
nand U6280 (N_6280,N_173,N_2343);
or U6281 (N_6281,N_732,N_3488);
or U6282 (N_6282,N_3287,N_4248);
and U6283 (N_6283,N_2678,N_51);
and U6284 (N_6284,N_3950,N_3286);
nand U6285 (N_6285,N_2624,N_2132);
nand U6286 (N_6286,N_4754,N_4297);
nor U6287 (N_6287,N_4252,N_2590);
nand U6288 (N_6288,N_2279,N_4669);
nand U6289 (N_6289,N_3313,N_464);
nand U6290 (N_6290,N_1853,N_2091);
nor U6291 (N_6291,N_3058,N_3787);
nor U6292 (N_6292,N_4227,N_4163);
or U6293 (N_6293,N_1175,N_539);
nand U6294 (N_6294,N_425,N_3851);
nor U6295 (N_6295,N_414,N_75);
and U6296 (N_6296,N_904,N_1040);
nand U6297 (N_6297,N_3900,N_3152);
nand U6298 (N_6298,N_3668,N_450);
nand U6299 (N_6299,N_2638,N_1714);
nand U6300 (N_6300,N_3352,N_1395);
and U6301 (N_6301,N_2325,N_3907);
and U6302 (N_6302,N_4607,N_3666);
nand U6303 (N_6303,N_1221,N_3195);
or U6304 (N_6304,N_4636,N_1297);
and U6305 (N_6305,N_37,N_1440);
or U6306 (N_6306,N_1056,N_3086);
nand U6307 (N_6307,N_1738,N_2163);
and U6308 (N_6308,N_3047,N_3800);
nor U6309 (N_6309,N_1906,N_4483);
nor U6310 (N_6310,N_4117,N_2433);
nand U6311 (N_6311,N_1261,N_4613);
nor U6312 (N_6312,N_2313,N_3220);
or U6313 (N_6313,N_2072,N_1986);
and U6314 (N_6314,N_4407,N_942);
and U6315 (N_6315,N_1079,N_1792);
or U6316 (N_6316,N_1167,N_1064);
and U6317 (N_6317,N_1195,N_2077);
and U6318 (N_6318,N_1272,N_2959);
nand U6319 (N_6319,N_2294,N_1109);
nor U6320 (N_6320,N_2542,N_481);
nand U6321 (N_6321,N_1599,N_3715);
nor U6322 (N_6322,N_249,N_2246);
nand U6323 (N_6323,N_3867,N_3890);
nor U6324 (N_6324,N_1057,N_2939);
nand U6325 (N_6325,N_4266,N_2585);
nor U6326 (N_6326,N_3045,N_4974);
nand U6327 (N_6327,N_3316,N_804);
and U6328 (N_6328,N_2785,N_1739);
nor U6329 (N_6329,N_4026,N_3327);
nor U6330 (N_6330,N_3568,N_4979);
nand U6331 (N_6331,N_141,N_3084);
or U6332 (N_6332,N_4123,N_4748);
or U6333 (N_6333,N_2844,N_2463);
nand U6334 (N_6334,N_4704,N_1890);
nor U6335 (N_6335,N_4235,N_4884);
nor U6336 (N_6336,N_1376,N_463);
nor U6337 (N_6337,N_4917,N_1051);
and U6338 (N_6338,N_2216,N_2196);
and U6339 (N_6339,N_2204,N_744);
and U6340 (N_6340,N_3525,N_4514);
nand U6341 (N_6341,N_2504,N_1839);
and U6342 (N_6342,N_2557,N_2330);
nor U6343 (N_6343,N_3933,N_1184);
nor U6344 (N_6344,N_2037,N_586);
or U6345 (N_6345,N_2439,N_2658);
and U6346 (N_6346,N_388,N_1909);
and U6347 (N_6347,N_2503,N_4431);
or U6348 (N_6348,N_4103,N_4413);
or U6349 (N_6349,N_272,N_1478);
and U6350 (N_6350,N_1866,N_2111);
nor U6351 (N_6351,N_2775,N_1072);
nand U6352 (N_6352,N_304,N_3066);
and U6353 (N_6353,N_62,N_3793);
nand U6354 (N_6354,N_880,N_2583);
or U6355 (N_6355,N_659,N_4196);
and U6356 (N_6356,N_2464,N_1354);
nor U6357 (N_6357,N_4402,N_4684);
nor U6358 (N_6358,N_2863,N_1120);
or U6359 (N_6359,N_2063,N_4535);
and U6360 (N_6360,N_3868,N_641);
and U6361 (N_6361,N_1606,N_1147);
or U6362 (N_6362,N_3561,N_1393);
or U6363 (N_6363,N_189,N_2303);
nor U6364 (N_6364,N_717,N_3310);
nor U6365 (N_6365,N_4443,N_4073);
or U6366 (N_6366,N_4137,N_566);
nand U6367 (N_6367,N_727,N_4452);
and U6368 (N_6368,N_1302,N_4831);
and U6369 (N_6369,N_2478,N_1005);
nor U6370 (N_6370,N_1188,N_1239);
nand U6371 (N_6371,N_951,N_1595);
and U6372 (N_6372,N_4486,N_3246);
or U6373 (N_6373,N_3958,N_3641);
nand U6374 (N_6374,N_1033,N_3048);
and U6375 (N_6375,N_806,N_2935);
or U6376 (N_6376,N_57,N_4381);
nand U6377 (N_6377,N_1489,N_805);
and U6378 (N_6378,N_3371,N_2058);
and U6379 (N_6379,N_4337,N_3166);
nand U6380 (N_6380,N_2649,N_780);
nor U6381 (N_6381,N_3967,N_165);
nand U6382 (N_6382,N_1737,N_4387);
or U6383 (N_6383,N_4448,N_2851);
nand U6384 (N_6384,N_4463,N_1319);
and U6385 (N_6385,N_2796,N_2217);
nand U6386 (N_6386,N_4351,N_4924);
or U6387 (N_6387,N_630,N_4509);
nor U6388 (N_6388,N_3544,N_3969);
nand U6389 (N_6389,N_704,N_3656);
or U6390 (N_6390,N_2051,N_585);
nor U6391 (N_6391,N_2357,N_2733);
and U6392 (N_6392,N_617,N_648);
or U6393 (N_6393,N_984,N_21);
nand U6394 (N_6394,N_2249,N_1134);
nand U6395 (N_6395,N_1565,N_71);
nand U6396 (N_6396,N_3615,N_3640);
and U6397 (N_6397,N_663,N_4894);
or U6398 (N_6398,N_1949,N_4498);
nand U6399 (N_6399,N_2726,N_2093);
nand U6400 (N_6400,N_4131,N_2281);
or U6401 (N_6401,N_3783,N_3959);
or U6402 (N_6402,N_1202,N_2941);
nand U6403 (N_6403,N_4857,N_1904);
and U6404 (N_6404,N_754,N_737);
nor U6405 (N_6405,N_4623,N_4504);
and U6406 (N_6406,N_2982,N_2243);
nand U6407 (N_6407,N_2860,N_4119);
nor U6408 (N_6408,N_4316,N_3474);
nor U6409 (N_6409,N_970,N_4506);
nand U6410 (N_6410,N_4233,N_932);
nand U6411 (N_6411,N_3672,N_1470);
or U6412 (N_6412,N_3306,N_84);
and U6413 (N_6413,N_4982,N_725);
nand U6414 (N_6414,N_4321,N_2552);
nor U6415 (N_6415,N_2745,N_4604);
nor U6416 (N_6416,N_149,N_2612);
and U6417 (N_6417,N_1741,N_4278);
and U6418 (N_6418,N_1546,N_1149);
or U6419 (N_6419,N_4161,N_2846);
nand U6420 (N_6420,N_4680,N_4363);
nor U6421 (N_6421,N_1108,N_1554);
nand U6422 (N_6422,N_3855,N_1123);
nand U6423 (N_6423,N_3724,N_1697);
nor U6424 (N_6424,N_4302,N_150);
nor U6425 (N_6425,N_3128,N_2650);
nand U6426 (N_6426,N_3987,N_4516);
nor U6427 (N_6427,N_2073,N_1087);
and U6428 (N_6428,N_36,N_1657);
and U6429 (N_6429,N_1435,N_4998);
nor U6430 (N_6430,N_2532,N_3601);
xor U6431 (N_6431,N_3920,N_4305);
or U6432 (N_6432,N_4816,N_4635);
and U6433 (N_6433,N_3949,N_1007);
or U6434 (N_6434,N_4488,N_3123);
nand U6435 (N_6435,N_3142,N_2833);
or U6436 (N_6436,N_1629,N_4675);
or U6437 (N_6437,N_136,N_1568);
or U6438 (N_6438,N_3434,N_770);
or U6439 (N_6439,N_1846,N_1497);
nand U6440 (N_6440,N_1126,N_756);
and U6441 (N_6441,N_430,N_729);
or U6442 (N_6442,N_217,N_2185);
nand U6443 (N_6443,N_1571,N_799);
nand U6444 (N_6444,N_4707,N_2085);
and U6445 (N_6445,N_4265,N_779);
nand U6446 (N_6446,N_1014,N_3954);
and U6447 (N_6447,N_2082,N_765);
and U6448 (N_6448,N_2866,N_3002);
nor U6449 (N_6449,N_3560,N_4987);
nor U6450 (N_6450,N_1070,N_3482);
and U6451 (N_6451,N_972,N_3094);
and U6452 (N_6452,N_1192,N_1690);
and U6453 (N_6453,N_2686,N_4792);
or U6454 (N_6454,N_1235,N_3731);
and U6455 (N_6455,N_3514,N_491);
or U6456 (N_6456,N_2950,N_2953);
and U6457 (N_6457,N_4710,N_3822);
or U6458 (N_6458,N_1131,N_3698);
and U6459 (N_6459,N_2413,N_2764);
and U6460 (N_6460,N_692,N_2320);
or U6461 (N_6461,N_3,N_2872);
and U6462 (N_6462,N_1114,N_2821);
xnor U6463 (N_6463,N_1111,N_3575);
nor U6464 (N_6464,N_3008,N_4864);
or U6465 (N_6465,N_2660,N_797);
nand U6466 (N_6466,N_4944,N_110);
or U6467 (N_6467,N_178,N_1405);
and U6468 (N_6468,N_2563,N_3427);
and U6469 (N_6469,N_954,N_3180);
or U6470 (N_6470,N_1459,N_4415);
nand U6471 (N_6471,N_2506,N_345);
nand U6472 (N_6472,N_4226,N_2676);
or U6473 (N_6473,N_4400,N_1287);
nand U6474 (N_6474,N_3088,N_4867);
nor U6475 (N_6475,N_2566,N_3922);
nand U6476 (N_6476,N_4251,N_2147);
nor U6477 (N_6477,N_1740,N_1358);
nor U6478 (N_6478,N_2490,N_3367);
nor U6479 (N_6479,N_3193,N_4892);
or U6480 (N_6480,N_3062,N_538);
and U6481 (N_6481,N_2949,N_3940);
nor U6482 (N_6482,N_2608,N_4242);
nand U6483 (N_6483,N_2434,N_1434);
or U6484 (N_6484,N_1639,N_556);
or U6485 (N_6485,N_730,N_1567);
nor U6486 (N_6486,N_2046,N_411);
and U6487 (N_6487,N_1713,N_3694);
or U6488 (N_6488,N_4074,N_2211);
nand U6489 (N_6489,N_1163,N_2903);
or U6490 (N_6490,N_2331,N_4323);
nor U6491 (N_6491,N_406,N_3373);
nand U6492 (N_6492,N_4064,N_2265);
nor U6493 (N_6493,N_308,N_1637);
and U6494 (N_6494,N_485,N_3217);
and U6495 (N_6495,N_1894,N_2222);
or U6496 (N_6496,N_2865,N_1927);
nand U6497 (N_6497,N_836,N_319);
nand U6498 (N_6498,N_802,N_2696);
nand U6499 (N_6499,N_3834,N_3319);
and U6500 (N_6500,N_389,N_4168);
nor U6501 (N_6501,N_2452,N_3653);
or U6502 (N_6502,N_517,N_4805);
or U6503 (N_6503,N_297,N_1907);
or U6504 (N_6504,N_1880,N_2327);
nor U6505 (N_6505,N_3589,N_258);
and U6506 (N_6506,N_166,N_3054);
or U6507 (N_6507,N_2466,N_2240);
nand U6508 (N_6508,N_4718,N_4156);
nor U6509 (N_6509,N_4301,N_795);
and U6510 (N_6510,N_1550,N_4625);
nor U6511 (N_6511,N_1876,N_4095);
and U6512 (N_6512,N_1624,N_1095);
nor U6513 (N_6513,N_2803,N_3095);
nor U6514 (N_6514,N_360,N_3329);
and U6515 (N_6515,N_2202,N_1579);
nor U6516 (N_6516,N_3368,N_1821);
nor U6517 (N_6517,N_845,N_946);
nand U6518 (N_6518,N_557,N_2697);
and U6519 (N_6519,N_3386,N_1006);
and U6520 (N_6520,N_444,N_3823);
and U6521 (N_6521,N_2054,N_2241);
nor U6522 (N_6522,N_1901,N_12);
and U6523 (N_6523,N_3383,N_964);
nand U6524 (N_6524,N_1973,N_2756);
and U6525 (N_6525,N_3658,N_128);
and U6526 (N_6526,N_2931,N_2292);
or U6527 (N_6527,N_4980,N_2056);
or U6528 (N_6528,N_2925,N_4466);
and U6529 (N_6529,N_881,N_1156);
nor U6530 (N_6530,N_3516,N_332);
nor U6531 (N_6531,N_4591,N_1226);
and U6532 (N_6532,N_2109,N_1885);
nand U6533 (N_6533,N_3222,N_3276);
or U6534 (N_6534,N_2455,N_1305);
nand U6535 (N_6535,N_221,N_2129);
nor U6536 (N_6536,N_4331,N_4247);
or U6537 (N_6537,N_16,N_4290);
nand U6538 (N_6538,N_3618,N_2962);
and U6539 (N_6539,N_22,N_164);
and U6540 (N_6540,N_1827,N_3106);
nor U6541 (N_6541,N_4713,N_1748);
and U6542 (N_6542,N_1959,N_3605);
nor U6543 (N_6543,N_1641,N_2019);
or U6544 (N_6544,N_790,N_3477);
nor U6545 (N_6545,N_2421,N_302);
nand U6546 (N_6546,N_2228,N_533);
nand U6547 (N_6547,N_2245,N_4665);
or U6548 (N_6548,N_3642,N_3223);
and U6549 (N_6549,N_4051,N_1717);
or U6550 (N_6550,N_1582,N_3896);
nor U6551 (N_6551,N_2955,N_2015);
nand U6552 (N_6552,N_2694,N_2816);
and U6553 (N_6553,N_1742,N_1465);
nand U6554 (N_6554,N_2888,N_3487);
nand U6555 (N_6555,N_4556,N_3876);
nand U6556 (N_6556,N_105,N_3151);
and U6557 (N_6557,N_930,N_4198);
nand U6558 (N_6558,N_2453,N_3980);
and U6559 (N_6559,N_708,N_1041);
nand U6560 (N_6560,N_350,N_4827);
nor U6561 (N_6561,N_2498,N_1730);
nor U6562 (N_6562,N_4450,N_448);
nand U6563 (N_6563,N_4046,N_2614);
or U6564 (N_6564,N_542,N_728);
nand U6565 (N_6565,N_2984,N_1092);
or U6566 (N_6566,N_471,N_4114);
nor U6567 (N_6567,N_1749,N_2749);
nand U6568 (N_6568,N_2862,N_4294);
or U6569 (N_6569,N_2302,N_3624);
and U6570 (N_6570,N_4205,N_687);
nor U6571 (N_6571,N_3534,N_4631);
and U6572 (N_6572,N_4194,N_2412);
nor U6573 (N_6573,N_4661,N_1745);
nand U6574 (N_6574,N_2544,N_1649);
nand U6575 (N_6575,N_3848,N_3007);
or U6576 (N_6576,N_3579,N_3143);
nor U6577 (N_6577,N_537,N_4926);
and U6578 (N_6578,N_2423,N_365);
or U6579 (N_6579,N_3669,N_2075);
nor U6580 (N_6580,N_733,N_611);
and U6581 (N_6581,N_3813,N_4735);
or U6582 (N_6582,N_2130,N_3108);
nor U6583 (N_6583,N_4264,N_1278);
nand U6584 (N_6584,N_157,N_574);
nor U6585 (N_6585,N_1652,N_3965);
nand U6586 (N_6586,N_3545,N_903);
nor U6587 (N_6587,N_3894,N_2451);
and U6588 (N_6588,N_4683,N_4464);
or U6589 (N_6589,N_1256,N_678);
nor U6590 (N_6590,N_573,N_3089);
and U6591 (N_6591,N_584,N_3292);
and U6592 (N_6592,N_4691,N_1704);
nor U6593 (N_6593,N_3768,N_724);
nand U6594 (N_6594,N_871,N_4087);
nor U6595 (N_6595,N_1622,N_2008);
nor U6596 (N_6596,N_3776,N_3278);
nand U6597 (N_6597,N_2431,N_4432);
or U6598 (N_6598,N_4027,N_2671);
nor U6599 (N_6599,N_2190,N_3206);
and U6600 (N_6600,N_412,N_4442);
nand U6601 (N_6601,N_3179,N_2832);
nor U6602 (N_6602,N_938,N_576);
xor U6603 (N_6603,N_4040,N_1626);
or U6604 (N_6604,N_1002,N_1385);
nand U6605 (N_6605,N_4157,N_3607);
and U6606 (N_6606,N_4862,N_4262);
and U6607 (N_6607,N_2707,N_1476);
and U6608 (N_6608,N_2967,N_916);
or U6609 (N_6609,N_2568,N_4685);
nand U6610 (N_6610,N_303,N_2045);
nand U6611 (N_6611,N_4154,N_4269);
and U6612 (N_6612,N_1974,N_336);
and U6613 (N_6613,N_2734,N_1227);
nand U6614 (N_6614,N_3612,N_3154);
nor U6615 (N_6615,N_1246,N_4845);
nand U6616 (N_6616,N_109,N_752);
and U6617 (N_6617,N_4752,N_2632);
or U6618 (N_6618,N_1607,N_3617);
nand U6619 (N_6619,N_1561,N_3231);
nor U6620 (N_6620,N_4508,N_1575);
and U6621 (N_6621,N_736,N_2167);
and U6622 (N_6622,N_3479,N_1276);
and U6623 (N_6623,N_1873,N_1267);
or U6624 (N_6624,N_3840,N_266);
or U6625 (N_6625,N_4557,N_2531);
and U6626 (N_6626,N_1831,N_3259);
and U6627 (N_6627,N_679,N_590);
or U6628 (N_6628,N_973,N_1725);
or U6629 (N_6629,N_2150,N_3072);
or U6630 (N_6630,N_4475,N_760);
xor U6631 (N_6631,N_735,N_1104);
nand U6632 (N_6632,N_2629,N_4572);
and U6633 (N_6633,N_3456,N_4961);
nor U6634 (N_6634,N_198,N_4801);
nor U6635 (N_6635,N_734,N_3196);
and U6636 (N_6636,N_1896,N_2957);
nand U6637 (N_6637,N_1096,N_1201);
nand U6638 (N_6638,N_4714,N_709);
and U6639 (N_6639,N_3021,N_3103);
nand U6640 (N_6640,N_23,N_372);
nor U6641 (N_6641,N_3686,N_2634);
nand U6642 (N_6642,N_1685,N_4239);
nand U6643 (N_6643,N_807,N_2852);
and U6644 (N_6644,N_3314,N_4021);
or U6645 (N_6645,N_1091,N_2002);
or U6646 (N_6646,N_2,N_3320);
and U6647 (N_6647,N_642,N_908);
nor U6648 (N_6648,N_4304,N_2964);
nor U6649 (N_6649,N_1849,N_42);
and U6650 (N_6650,N_4849,N_1473);
nand U6651 (N_6651,N_2772,N_3219);
nand U6652 (N_6652,N_2501,N_270);
nand U6653 (N_6653,N_443,N_3254);
and U6654 (N_6654,N_527,N_3376);
or U6655 (N_6655,N_212,N_2598);
or U6656 (N_6656,N_957,N_4501);
nand U6657 (N_6657,N_1638,N_2714);
and U6658 (N_6658,N_148,N_2725);
or U6659 (N_6659,N_1200,N_4276);
or U6660 (N_6660,N_914,N_94);
nor U6661 (N_6661,N_877,N_955);
nand U6662 (N_6662,N_644,N_3121);
nor U6663 (N_6663,N_2459,N_3818);
nand U6664 (N_6664,N_2896,N_913);
nor U6665 (N_6665,N_2508,N_4322);
and U6666 (N_6666,N_1335,N_4012);
nand U6667 (N_6667,N_1408,N_3584);
nand U6668 (N_6668,N_3241,N_3409);
and U6669 (N_6669,N_1168,N_4559);
nand U6670 (N_6670,N_111,N_3018);
nand U6671 (N_6671,N_1814,N_3735);
and U6672 (N_6672,N_1966,N_3126);
or U6673 (N_6673,N_2795,N_1868);
or U6674 (N_6674,N_2354,N_4291);
nor U6675 (N_6675,N_2664,N_2599);
or U6676 (N_6676,N_246,N_3859);
or U6677 (N_6677,N_1062,N_509);
nor U6678 (N_6678,N_1775,N_4401);
and U6679 (N_6679,N_3511,N_2416);
or U6680 (N_6680,N_1766,N_2365);
nor U6681 (N_6681,N_2427,N_1523);
or U6682 (N_6682,N_4063,N_1035);
or U6683 (N_6683,N_4162,N_2363);
xnor U6684 (N_6684,N_2511,N_376);
nand U6685 (N_6685,N_1164,N_882);
or U6686 (N_6686,N_1572,N_4606);
or U6687 (N_6687,N_3751,N_171);
nor U6688 (N_6688,N_2282,N_1355);
nand U6689 (N_6689,N_2029,N_2479);
nand U6690 (N_6690,N_2425,N_1438);
nor U6691 (N_6691,N_2972,N_3082);
nor U6692 (N_6692,N_4567,N_1922);
and U6693 (N_6693,N_1610,N_776);
or U6694 (N_6694,N_672,N_428);
nand U6695 (N_6695,N_3262,N_3557);
nor U6696 (N_6696,N_4821,N_2028);
and U6697 (N_6697,N_469,N_828);
nand U6698 (N_6698,N_2806,N_3846);
or U6699 (N_6699,N_793,N_1819);
and U6700 (N_6700,N_2036,N_1612);
and U6701 (N_6701,N_294,N_3587);
and U6702 (N_6702,N_1549,N_3345);
and U6703 (N_6703,N_2392,N_3233);
nand U6704 (N_6704,N_3753,N_1242);
and U6705 (N_6705,N_181,N_4776);
nor U6706 (N_6706,N_3966,N_3722);
nor U6707 (N_6707,N_1643,N_3912);
nor U6708 (N_6708,N_4855,N_477);
nor U6709 (N_6709,N_4652,N_3766);
or U6710 (N_6710,N_229,N_3394);
and U6711 (N_6711,N_4664,N_1648);
or U6712 (N_6712,N_19,N_2643);
nand U6713 (N_6713,N_1413,N_927);
nand U6714 (N_6714,N_1012,N_2621);
or U6715 (N_6715,N_4728,N_4678);
and U6716 (N_6716,N_2882,N_1844);
nor U6717 (N_6717,N_1241,N_3326);
nor U6718 (N_6718,N_1545,N_3377);
or U6719 (N_6719,N_748,N_623);
nor U6720 (N_6720,N_3852,N_224);
nand U6721 (N_6721,N_1818,N_1964);
and U6722 (N_6722,N_2467,N_698);
nand U6723 (N_6723,N_2489,N_3134);
and U6724 (N_6724,N_2673,N_707);
nor U6725 (N_6725,N_1495,N_2657);
nand U6726 (N_6726,N_3100,N_373);
and U6727 (N_6727,N_2909,N_2395);
or U6728 (N_6728,N_3501,N_1857);
or U6729 (N_6729,N_4782,N_4650);
nand U6730 (N_6730,N_2724,N_3508);
or U6731 (N_6731,N_2485,N_3866);
or U6732 (N_6732,N_791,N_2577);
or U6733 (N_6733,N_4584,N_1912);
and U6734 (N_6734,N_1142,N_4536);
and U6735 (N_6735,N_357,N_4800);
nor U6736 (N_6736,N_2080,N_3460);
and U6737 (N_6737,N_3986,N_1655);
nor U6738 (N_6738,N_677,N_4176);
nand U6739 (N_6739,N_4234,N_251);
and U6740 (N_6740,N_1576,N_3808);
nor U6741 (N_6741,N_1608,N_3183);
nor U6742 (N_6742,N_4175,N_4936);
and U6743 (N_6743,N_4820,N_4577);
or U6744 (N_6744,N_4000,N_2854);
or U6745 (N_6745,N_2181,N_3820);
and U6746 (N_6746,N_1564,N_3159);
or U6747 (N_6747,N_442,N_2096);
or U6748 (N_6748,N_2829,N_3272);
or U6749 (N_6749,N_2708,N_2849);
or U6750 (N_6750,N_499,N_2026);
and U6751 (N_6751,N_3864,N_4014);
or U6752 (N_6752,N_1632,N_4237);
nand U6753 (N_6753,N_1003,N_4275);
nor U6754 (N_6754,N_2460,N_3764);
nand U6755 (N_6755,N_1365,N_1824);
nor U6756 (N_6756,N_4880,N_4201);
nor U6757 (N_6757,N_2342,N_4097);
nand U6758 (N_6758,N_3457,N_4439);
nor U6759 (N_6759,N_3473,N_279);
or U6760 (N_6760,N_1544,N_134);
or U6761 (N_6761,N_1672,N_699);
nor U6762 (N_6762,N_2106,N_3238);
and U6763 (N_6763,N_1386,N_4470);
nand U6764 (N_6764,N_1592,N_2105);
nand U6765 (N_6765,N_1325,N_787);
nor U6766 (N_6766,N_3588,N_3348);
and U6767 (N_6767,N_3493,N_4695);
and U6768 (N_6768,N_3882,N_230);
or U6769 (N_6769,N_3688,N_2450);
and U6770 (N_6770,N_4734,N_2710);
nand U6771 (N_6771,N_4392,N_1058);
and U6772 (N_6772,N_2874,N_706);
nand U6773 (N_6773,N_4230,N_4749);
nand U6774 (N_6774,N_851,N_2825);
and U6775 (N_6775,N_781,N_2709);
and U6776 (N_6776,N_1251,N_2974);
nand U6777 (N_6777,N_3075,N_117);
and U6778 (N_6778,N_3843,N_2261);
nand U6779 (N_6779,N_3755,N_4145);
nand U6780 (N_6780,N_3634,N_3582);
or U6781 (N_6781,N_1903,N_4003);
nand U6782 (N_6782,N_3370,N_2176);
nor U6783 (N_6783,N_1642,N_1789);
nor U6784 (N_6784,N_2604,N_175);
nand U6785 (N_6785,N_1475,N_2253);
nand U6786 (N_6786,N_4444,N_2899);
nor U6787 (N_6787,N_652,N_4966);
nor U6788 (N_6788,N_1921,N_3392);
nor U6789 (N_6789,N_1796,N_2404);
and U6790 (N_6790,N_1747,N_2535);
and U6791 (N_6791,N_4366,N_4837);
and U6792 (N_6792,N_3599,N_4553);
and U6793 (N_6793,N_917,N_3665);
and U6794 (N_6794,N_2753,N_4573);
nor U6795 (N_6795,N_2065,N_183);
and U6796 (N_6796,N_2928,N_2766);
nand U6797 (N_6797,N_1771,N_419);
or U6798 (N_6798,N_34,N_3229);
nor U6799 (N_6799,N_2361,N_1299);
nand U6800 (N_6800,N_1400,N_2920);
nand U6801 (N_6801,N_3998,N_3191);
nor U6802 (N_6802,N_1929,N_3497);
and U6803 (N_6803,N_4598,N_340);
nor U6804 (N_6804,N_3244,N_3285);
and U6805 (N_6805,N_96,N_3989);
or U6806 (N_6806,N_4698,N_3181);
or U6807 (N_6807,N_4644,N_2790);
nor U6808 (N_6808,N_1061,N_2145);
nand U6809 (N_6809,N_275,N_3865);
or U6810 (N_6810,N_545,N_4620);
nand U6811 (N_6811,N_2545,N_4353);
or U6812 (N_6812,N_322,N_61);
or U6813 (N_6813,N_1042,N_2131);
nand U6814 (N_6814,N_486,N_1382);
or U6815 (N_6815,N_4462,N_618);
nand U6816 (N_6816,N_4274,N_231);
or U6817 (N_6817,N_2146,N_4523);
or U6818 (N_6818,N_2798,N_2438);
nor U6819 (N_6819,N_1512,N_4519);
nor U6820 (N_6820,N_1238,N_1902);
nand U6821 (N_6821,N_3484,N_1950);
nand U6822 (N_6822,N_4947,N_2721);
and U6823 (N_6823,N_252,N_2159);
nand U6824 (N_6824,N_2023,N_1230);
or U6825 (N_6825,N_4724,N_2061);
and U6826 (N_6826,N_3261,N_1312);
nand U6827 (N_6827,N_4182,N_4192);
nand U6828 (N_6828,N_612,N_3486);
nand U6829 (N_6829,N_1357,N_665);
nor U6830 (N_6830,N_2722,N_907);
or U6831 (N_6831,N_4853,N_4829);
nand U6832 (N_6832,N_4153,N_3811);
nor U6833 (N_6833,N_896,N_4364);
nand U6834 (N_6834,N_3957,N_3171);
nand U6835 (N_6835,N_800,N_541);
and U6836 (N_6836,N_2496,N_1623);
nor U6837 (N_6837,N_1265,N_417);
and U6838 (N_6838,N_855,N_4513);
and U6839 (N_6839,N_2820,N_1105);
nand U6840 (N_6840,N_3976,N_2380);
or U6841 (N_6841,N_547,N_2194);
nor U6842 (N_6842,N_1000,N_273);
xnor U6843 (N_6843,N_992,N_3754);
or U6844 (N_6844,N_1390,N_1086);
nor U6845 (N_6845,N_1664,N_4180);
and U6846 (N_6846,N_4134,N_1078);
nor U6847 (N_6847,N_3858,N_1755);
nand U6848 (N_6848,N_2319,N_160);
or U6849 (N_6849,N_2004,N_4416);
or U6850 (N_6850,N_11,N_3187);
nand U6851 (N_6851,N_862,N_3574);
nand U6852 (N_6852,N_1367,N_1705);
nor U6853 (N_6853,N_4370,N_2944);
nand U6854 (N_6854,N_1368,N_626);
or U6855 (N_6855,N_2383,N_2781);
nor U6856 (N_6856,N_888,N_1681);
nand U6857 (N_6857,N_2359,N_103);
nand U6858 (N_6858,N_4670,N_3841);
nand U6859 (N_6859,N_89,N_1958);
or U6860 (N_6860,N_4742,N_1560);
nor U6861 (N_6861,N_2681,N_3548);
nor U6862 (N_6862,N_3057,N_3140);
nand U6863 (N_6863,N_635,N_122);
and U6864 (N_6864,N_3132,N_2861);
or U6865 (N_6865,N_1194,N_1208);
nand U6866 (N_6866,N_1389,N_14);
and U6867 (N_6867,N_1768,N_4143);
or U6868 (N_6868,N_608,N_3522);
nand U6869 (N_6869,N_3710,N_2539);
nor U6870 (N_6870,N_3210,N_4861);
or U6871 (N_6871,N_1143,N_4189);
and U6872 (N_6872,N_2819,N_1148);
nand U6873 (N_6873,N_1780,N_3472);
nand U6874 (N_6874,N_928,N_1524);
and U6875 (N_6875,N_2356,N_1820);
nand U6876 (N_6876,N_3224,N_3739);
nand U6877 (N_6877,N_1275,N_2768);
nor U6878 (N_6878,N_112,N_3001);
nand U6879 (N_6879,N_4478,N_996);
nand U6880 (N_6880,N_3789,N_1837);
nand U6881 (N_6881,N_1715,N_3346);
nor U6882 (N_6882,N_3024,N_1646);
and U6883 (N_6883,N_4005,N_145);
or U6884 (N_6884,N_4165,N_3104);
and U6885 (N_6885,N_2116,N_1800);
nand U6886 (N_6886,N_4204,N_4362);
nor U6887 (N_6887,N_4731,N_4545);
nor U6888 (N_6888,N_670,N_3917);
nand U6889 (N_6889,N_1939,N_4313);
or U6890 (N_6890,N_3878,N_1039);
or U6891 (N_6891,N_2068,N_1694);
and U6892 (N_6892,N_696,N_1249);
nor U6893 (N_6893,N_1121,N_2104);
nor U6894 (N_6894,N_3815,N_2737);
and U6895 (N_6895,N_2600,N_1336);
nand U6896 (N_6896,N_1248,N_3643);
nand U6897 (N_6897,N_4920,N_3931);
and U6898 (N_6898,N_3092,N_3446);
nand U6899 (N_6899,N_2730,N_2958);
or U6900 (N_6900,N_1858,N_70);
and U6901 (N_6901,N_1533,N_4972);
or U6902 (N_6902,N_4771,N_902);
nor U6903 (N_6903,N_320,N_403);
or U6904 (N_6904,N_2367,N_3061);
nor U6905 (N_6905,N_2368,N_2639);
and U6906 (N_6906,N_4283,N_2493);
nor U6907 (N_6907,N_3674,N_2030);
or U6908 (N_6908,N_873,N_2690);
or U6909 (N_6909,N_1342,N_4793);
and U6910 (N_6910,N_4910,N_2432);
nor U6911 (N_6911,N_3213,N_4202);
or U6912 (N_6912,N_2417,N_2353);
or U6913 (N_6913,N_317,N_1493);
nor U6914 (N_6914,N_3331,N_2199);
nand U6915 (N_6915,N_2826,N_4941);
nor U6916 (N_6916,N_3636,N_4169);
and U6917 (N_6917,N_4495,N_2729);
nor U6918 (N_6918,N_2293,N_2178);
nand U6919 (N_6919,N_4909,N_2349);
nand U6920 (N_6920,N_2654,N_2089);
and U6921 (N_6921,N_4624,N_2215);
nand U6922 (N_6922,N_982,N_2100);
or U6923 (N_6923,N_1746,N_291);
and U6924 (N_6924,N_1919,N_1211);
nand U6925 (N_6925,N_3070,N_719);
nor U6926 (N_6926,N_4033,N_3198);
and U6927 (N_6927,N_1513,N_4408);
nand U6928 (N_6928,N_2519,N_8);
nor U6929 (N_6929,N_3530,N_2193);
and U6930 (N_6930,N_953,N_2378);
nor U6931 (N_6931,N_4099,N_593);
or U6932 (N_6932,N_4761,N_4155);
and U6933 (N_6933,N_2759,N_1993);
nor U6934 (N_6934,N_2952,N_2877);
nand U6935 (N_6935,N_4770,N_3471);
nor U6936 (N_6936,N_823,N_369);
or U6937 (N_6937,N_3990,N_4497);
nand U6938 (N_6938,N_2716,N_3875);
nor U6939 (N_6939,N_1874,N_3573);
nand U6940 (N_6940,N_3623,N_2274);
or U6941 (N_6941,N_4611,N_4440);
and U6942 (N_6942,N_819,N_2027);
and U6943 (N_6943,N_2221,N_507);
or U6944 (N_6944,N_3435,N_2191);
nor U6945 (N_6945,N_4375,N_4379);
nand U6946 (N_6946,N_2992,N_1234);
and U6947 (N_6947,N_3681,N_4968);
and U6948 (N_6948,N_1753,N_975);
nor U6949 (N_6949,N_1923,N_1152);
or U6950 (N_6950,N_885,N_1954);
nor U6951 (N_6951,N_3291,N_4507);
and U6952 (N_6952,N_3697,N_1604);
and U6953 (N_6953,N_616,N_2769);
nor U6954 (N_6954,N_501,N_4727);
and U6955 (N_6955,N_3288,N_2640);
nor U6956 (N_6956,N_656,N_1397);
or U6957 (N_6957,N_2236,N_3208);
nor U6958 (N_6958,N_1093,N_2996);
nand U6959 (N_6959,N_3411,N_2991);
nor U6960 (N_6960,N_3078,N_945);
and U6961 (N_6961,N_1763,N_93);
and U6962 (N_6962,N_1073,N_711);
or U6963 (N_6963,N_3733,N_399);
or U6964 (N_6964,N_1384,N_3067);
or U6965 (N_6965,N_3138,N_720);
nor U6966 (N_6966,N_1469,N_356);
nor U6967 (N_6967,N_614,N_514);
nand U6968 (N_6968,N_4950,N_4654);
nand U6969 (N_6969,N_395,N_1899);
and U6970 (N_6970,N_4561,N_3862);
nor U6971 (N_6971,N_4813,N_4485);
or U6972 (N_6972,N_4359,N_4378);
and U6973 (N_6973,N_4622,N_1049);
nor U6974 (N_6974,N_243,N_26);
nor U6975 (N_6975,N_1826,N_3055);
nand U6976 (N_6976,N_1264,N_46);
nor U6977 (N_6977,N_3491,N_2326);
nand U6978 (N_6978,N_1455,N_1141);
or U6979 (N_6979,N_4945,N_1180);
and U6980 (N_6980,N_3122,N_3146);
or U6981 (N_6981,N_1712,N_859);
nor U6982 (N_6982,N_2403,N_3799);
nand U6983 (N_6983,N_2441,N_4958);
or U6984 (N_6984,N_943,N_919);
and U6985 (N_6985,N_3465,N_2706);
nor U6986 (N_6986,N_3393,N_844);
nor U6987 (N_6987,N_4421,N_3625);
or U6988 (N_6988,N_2407,N_2549);
or U6989 (N_6989,N_2677,N_3533);
and U6990 (N_6990,N_482,N_944);
nand U6991 (N_6991,N_550,N_2252);
or U6992 (N_6992,N_244,N_2954);
or U6993 (N_6993,N_2648,N_3449);
nand U6994 (N_6994,N_3342,N_1535);
nand U6995 (N_6995,N_2430,N_142);
nor U6996 (N_6996,N_3972,N_2168);
nand U6997 (N_6997,N_1682,N_3635);
nand U6998 (N_6998,N_4588,N_3628);
or U6999 (N_6999,N_4172,N_2203);
or U7000 (N_7000,N_4788,N_1439);
nor U7001 (N_7001,N_2044,N_4541);
and U7002 (N_7002,N_4214,N_1066);
and U7003 (N_7003,N_3385,N_3382);
or U7004 (N_7004,N_3888,N_629);
and U7005 (N_7005,N_4011,N_222);
nand U7006 (N_7006,N_809,N_814);
and U7007 (N_7007,N_772,N_2310);
and U7008 (N_7008,N_4047,N_2336);
nand U7009 (N_7009,N_1089,N_3336);
and U7010 (N_7010,N_49,N_3194);
nand U7011 (N_7011,N_1955,N_3645);
nor U7012 (N_7012,N_288,N_2688);
nand U7013 (N_7013,N_1924,N_3527);
and U7014 (N_7014,N_4135,N_3035);
and U7015 (N_7015,N_2334,N_1870);
nand U7016 (N_7016,N_2606,N_2152);
nand U7017 (N_7017,N_3243,N_2683);
nand U7018 (N_7018,N_3654,N_3532);
and U7019 (N_7019,N_2675,N_3349);
or U7020 (N_7020,N_1961,N_1428);
xor U7021 (N_7021,N_4594,N_4835);
and U7022 (N_7022,N_4149,N_4340);
nand U7023 (N_7023,N_3853,N_3730);
nand U7024 (N_7024,N_3050,N_3443);
or U7025 (N_7025,N_69,N_1596);
or U7026 (N_7026,N_3256,N_2693);
or U7027 (N_7027,N_3042,N_3879);
nor U7028 (N_7028,N_4896,N_4527);
and U7029 (N_7029,N_4603,N_2321);
and U7030 (N_7030,N_1621,N_4494);
or U7031 (N_7031,N_2691,N_4558);
or U7032 (N_7032,N_4032,N_1589);
nand U7033 (N_7033,N_3564,N_2227);
nand U7034 (N_7034,N_4959,N_3979);
or U7035 (N_7035,N_4057,N_4173);
nand U7036 (N_7036,N_620,N_3721);
nor U7037 (N_7037,N_1765,N_3239);
nand U7038 (N_7038,N_3592,N_866);
or U7039 (N_7039,N_561,N_4082);
and U7040 (N_7040,N_661,N_634);
nand U7041 (N_7041,N_2440,N_4484);
nor U7042 (N_7042,N_1333,N_4574);
nor U7043 (N_7043,N_4216,N_3927);
nor U7044 (N_7044,N_2788,N_743);
and U7045 (N_7045,N_3873,N_605);
or U7046 (N_7046,N_4220,N_1218);
and U7047 (N_7047,N_1761,N_4703);
and U7048 (N_7048,N_3404,N_2810);
nand U7049 (N_7049,N_3619,N_1928);
nor U7050 (N_7050,N_2615,N_2142);
nand U7051 (N_7051,N_1803,N_703);
nor U7052 (N_7052,N_177,N_1708);
and U7053 (N_7053,N_2853,N_1047);
nor U7054 (N_7054,N_1829,N_1764);
and U7055 (N_7055,N_3938,N_2119);
nor U7056 (N_7056,N_2979,N_3201);
nor U7057 (N_7057,N_2475,N_82);
nand U7058 (N_7058,N_628,N_4843);
nor U7059 (N_7059,N_588,N_1052);
or U7060 (N_7060,N_4616,N_3172);
nor U7061 (N_7061,N_4694,N_3586);
or U7062 (N_7062,N_4874,N_1417);
or U7063 (N_7063,N_2602,N_3283);
nor U7064 (N_7064,N_2212,N_335);
nand U7065 (N_7065,N_1528,N_4791);
nor U7066 (N_7066,N_3594,N_3856);
nor U7067 (N_7067,N_2476,N_475);
or U7068 (N_7068,N_2655,N_4396);
or U7069 (N_7069,N_2381,N_792);
nor U7070 (N_7070,N_2306,N_2420);
or U7071 (N_7071,N_2275,N_4628);
or U7072 (N_7072,N_2206,N_4667);
nand U7073 (N_7073,N_210,N_3063);
nor U7074 (N_7074,N_197,N_4456);
and U7075 (N_7075,N_2025,N_2376);
and U7076 (N_7076,N_2921,N_4018);
nor U7077 (N_7077,N_2887,N_1215);
nand U7078 (N_7078,N_4050,N_1995);
nand U7079 (N_7079,N_2177,N_2346);
and U7080 (N_7080,N_2684,N_3994);
nand U7081 (N_7081,N_1828,N_3163);
and U7082 (N_7082,N_4711,N_434);
or U7083 (N_7083,N_2192,N_1791);
and U7084 (N_7084,N_2879,N_1349);
and U7085 (N_7085,N_418,N_1205);
and U7086 (N_7086,N_4476,N_4492);
or U7087 (N_7087,N_1816,N_3984);
and U7088 (N_7088,N_3825,N_511);
and U7089 (N_7089,N_910,N_1236);
nor U7090 (N_7090,N_255,N_1069);
nor U7091 (N_7091,N_1084,N_4158);
or U7092 (N_7092,N_1509,N_3344);
nand U7093 (N_7093,N_4166,N_4528);
xor U7094 (N_7094,N_1553,N_640);
nand U7095 (N_7095,N_2986,N_1998);
and U7096 (N_7096,N_4141,N_583);
and U7097 (N_7097,N_564,N_223);
and U7098 (N_7098,N_4199,N_1081);
nand U7099 (N_7099,N_3389,N_4696);
and U7100 (N_7100,N_301,N_346);
nand U7101 (N_7101,N_277,N_3785);
nand U7102 (N_7102,N_1280,N_2780);
and U7103 (N_7103,N_1659,N_2571);
nor U7104 (N_7104,N_1822,N_4575);
nor U7105 (N_7105,N_1915,N_4647);
or U7106 (N_7106,N_1992,N_1350);
and U7107 (N_7107,N_4263,N_174);
nor U7108 (N_7108,N_409,N_284);
or U7109 (N_7109,N_2419,N_3509);
or U7110 (N_7110,N_1277,N_4211);
nor U7111 (N_7111,N_1840,N_3109);
and U7112 (N_7112,N_3459,N_77);
nor U7113 (N_7113,N_3267,N_1303);
or U7114 (N_7114,N_2843,N_3978);
or U7115 (N_7115,N_2039,N_3361);
and U7116 (N_7116,N_1323,N_3230);
nand U7117 (N_7117,N_4184,N_3226);
nor U7118 (N_7118,N_2133,N_300);
or U7119 (N_7119,N_2382,N_2347);
or U7120 (N_7120,N_3639,N_3312);
nand U7121 (N_7121,N_4999,N_311);
and U7122 (N_7122,N_1689,N_3485);
nor U7123 (N_7123,N_2698,N_3974);
and U7124 (N_7124,N_2213,N_2262);
nor U7125 (N_7125,N_977,N_1515);
nand U7126 (N_7126,N_1318,N_3794);
xnor U7127 (N_7127,N_4446,N_3069);
nor U7128 (N_7128,N_2198,N_4178);
nand U7129 (N_7129,N_4070,N_228);
nand U7130 (N_7130,N_1762,N_225);
nand U7131 (N_7131,N_1590,N_488);
or U7132 (N_7132,N_2792,N_3571);
nor U7133 (N_7133,N_2244,N_1133);
nand U7134 (N_7134,N_2436,N_2166);
or U7135 (N_7135,N_1027,N_638);
or U7136 (N_7136,N_1139,N_504);
nor U7137 (N_7137,N_3242,N_675);
nor U7138 (N_7138,N_4605,N_28);
and U7139 (N_7139,N_2134,N_900);
and U7140 (N_7140,N_4708,N_1212);
nand U7141 (N_7141,N_4847,N_2570);
and U7142 (N_7142,N_2906,N_2963);
nand U7143 (N_7143,N_525,N_1519);
nand U7144 (N_7144,N_3700,N_3651);
and U7145 (N_7145,N_4601,N_2171);
nand U7146 (N_7146,N_2258,N_3335);
and U7147 (N_7147,N_2740,N_2995);
nor U7148 (N_7148,N_1987,N_3444);
or U7149 (N_7149,N_3732,N_1817);
and U7150 (N_7150,N_4859,N_821);
nor U7151 (N_7151,N_1947,N_3006);
nand U7152 (N_7152,N_2558,N_4730);
and U7153 (N_7153,N_427,N_3567);
and U7154 (N_7154,N_3891,N_4267);
and U7155 (N_7155,N_3429,N_1735);
nor U7156 (N_7156,N_2225,N_2062);
nand U7157 (N_7157,N_1378,N_390);
and U7158 (N_7158,N_208,N_1288);
or U7159 (N_7159,N_4219,N_4593);
nand U7160 (N_7160,N_2437,N_3221);
nor U7161 (N_7161,N_76,N_4758);
or U7162 (N_7162,N_846,N_1861);
nor U7163 (N_7163,N_306,N_3357);
nand U7164 (N_7164,N_313,N_3480);
or U7165 (N_7165,N_1663,N_4041);
and U7166 (N_7166,N_4747,N_2997);
nand U7167 (N_7167,N_4,N_1247);
or U7168 (N_7168,N_1878,N_3167);
or U7169 (N_7169,N_1559,N_2472);
and U7170 (N_7170,N_3275,N_1356);
or U7171 (N_7171,N_2161,N_3430);
nor U7172 (N_7172,N_4732,N_2904);
nand U7173 (N_7173,N_299,N_4004);
or U7174 (N_7174,N_1077,N_1153);
and U7175 (N_7175,N_4893,N_438);
or U7176 (N_7176,N_188,N_2179);
nor U7177 (N_7177,N_2713,N_3863);
and U7178 (N_7178,N_3610,N_456);
or U7179 (N_7179,N_338,N_1647);
xor U7180 (N_7180,N_1291,N_3162);
and U7181 (N_7181,N_2800,N_784);
and U7182 (N_7182,N_632,N_3886);
and U7183 (N_7183,N_3087,N_4629);
nand U7184 (N_7184,N_3657,N_186);
nand U7185 (N_7185,N_2318,N_773);
nor U7186 (N_7186,N_1306,N_1862);
nand U7187 (N_7187,N_1815,N_1930);
nor U7188 (N_7188,N_658,N_3780);
nand U7189 (N_7189,N_3400,N_3452);
and U7190 (N_7190,N_4350,N_1597);
nand U7191 (N_7191,N_1651,N_2609);
nand U7192 (N_7192,N_1900,N_3696);
nand U7193 (N_7193,N_4885,N_2593);
nor U7194 (N_7194,N_4473,N_2400);
nor U7195 (N_7195,N_3300,N_921);
or U7196 (N_7196,N_2098,N_235);
nand U7197 (N_7197,N_746,N_1068);
and U7198 (N_7198,N_4491,N_4522);
or U7199 (N_7199,N_580,N_1609);
nor U7200 (N_7200,N_3173,N_3934);
and U7201 (N_7201,N_1151,N_762);
nor U7202 (N_7202,N_2020,N_3513);
and U7203 (N_7203,N_3767,N_1447);
nand U7204 (N_7204,N_3290,N_1085);
or U7205 (N_7205,N_3255,N_4296);
nand U7206 (N_7206,N_1798,N_518);
and U7207 (N_7207,N_242,N_1314);
nand U7208 (N_7208,N_1871,N_447);
and U7209 (N_7209,N_3332,N_519);
nor U7210 (N_7210,N_2257,N_3364);
nand U7211 (N_7211,N_4460,N_3621);
or U7212 (N_7212,N_424,N_2229);
nand U7213 (N_7213,N_392,N_2090);
and U7214 (N_7214,N_2943,N_4826);
nor U7215 (N_7215,N_1209,N_2070);
and U7216 (N_7216,N_4946,N_2260);
or U7217 (N_7217,N_2537,N_1757);
nor U7218 (N_7218,N_2556,N_2499);
or U7219 (N_7219,N_4013,N_3683);
nor U7220 (N_7220,N_366,N_4036);
nor U7221 (N_7221,N_3708,N_4354);
and U7222 (N_7222,N_4469,N_2187);
xor U7223 (N_7223,N_2497,N_312);
nor U7224 (N_7224,N_3432,N_446);
or U7225 (N_7225,N_812,N_1872);
and U7226 (N_7226,N_2858,N_218);
nand U7227 (N_7227,N_1808,N_613);
or U7228 (N_7228,N_3190,N_194);
or U7229 (N_7229,N_4037,N_4552);
nor U7230 (N_7230,N_1726,N_267);
nor U7231 (N_7231,N_3294,N_85);
nand U7232 (N_7232,N_362,N_1225);
nand U7233 (N_7233,N_426,N_1521);
and U7234 (N_7234,N_766,N_1744);
nand U7235 (N_7235,N_1446,N_1788);
or U7236 (N_7236,N_3478,N_966);
nor U7237 (N_7237,N_1375,N_1722);
nand U7238 (N_7238,N_4589,N_740);
and U7239 (N_7239,N_2214,N_484);
and U7240 (N_7240,N_1687,N_3264);
and U7241 (N_7241,N_3928,N_3085);
nor U7242 (N_7242,N_1008,N_4151);
or U7243 (N_7243,N_2776,N_3225);
or U7244 (N_7244,N_4160,N_1219);
nand U7245 (N_7245,N_3468,N_646);
or U7246 (N_7246,N_936,N_1852);
nor U7247 (N_7247,N_1301,N_3202);
or U7248 (N_7248,N_3736,N_3505);
and U7249 (N_7249,N_3609,N_960);
nor U7250 (N_7250,N_3682,N_1016);
nand U7251 (N_7251,N_4785,N_1823);
nor U7252 (N_7252,N_3939,N_1825);
nor U7253 (N_7253,N_649,N_3118);
nand U7254 (N_7254,N_4991,N_4630);
nor U7255 (N_7255,N_935,N_3036);
nor U7256 (N_7256,N_3496,N_4673);
and U7257 (N_7257,N_3550,N_1370);
and U7258 (N_7258,N_3413,N_2834);
nand U7259 (N_7259,N_10,N_4295);
nand U7260 (N_7260,N_3911,N_159);
and U7261 (N_7261,N_2042,N_2789);
or U7262 (N_7262,N_2875,N_2526);
nor U7263 (N_7263,N_1179,N_2529);
nor U7264 (N_7264,N_4803,N_3127);
nand U7265 (N_7265,N_3186,N_3073);
and U7266 (N_7266,N_2344,N_3763);
and U7267 (N_7267,N_4090,N_3237);
and U7268 (N_7268,N_4796,N_2255);
and U7269 (N_7269,N_1811,N_2248);
nor U7270 (N_7270,N_4879,N_4928);
nor U7271 (N_7271,N_4159,N_1243);
or U7272 (N_7272,N_2447,N_4104);
and U7273 (N_7273,N_2323,N_3555);
nor U7274 (N_7274,N_1352,N_4068);
and U7275 (N_7275,N_2603,N_6);
or U7276 (N_7276,N_4599,N_2817);
nand U7277 (N_7277,N_758,N_2534);
and U7278 (N_7278,N_2151,N_4001);
and U7279 (N_7279,N_4860,N_2071);
nor U7280 (N_7280,N_2727,N_2932);
nand U7281 (N_7281,N_2559,N_674);
and U7282 (N_7282,N_4537,N_264);
and U7283 (N_7283,N_3956,N_441);
and U7284 (N_7284,N_860,N_1920);
nand U7285 (N_7285,N_4781,N_102);
and U7286 (N_7286,N_506,N_7);
nor U7287 (N_7287,N_2283,N_1916);
nor U7288 (N_7288,N_723,N_4566);
nor U7289 (N_7289,N_1551,N_1018);
and U7290 (N_7290,N_4746,N_2937);
nand U7291 (N_7291,N_2377,N_2449);
or U7292 (N_7292,N_314,N_4964);
or U7293 (N_7293,N_4906,N_4256);
or U7294 (N_7294,N_570,N_1865);
nor U7295 (N_7295,N_2289,N_4139);
or U7296 (N_7296,N_3772,N_2469);
or U7297 (N_7297,N_2340,N_4655);
nand U7298 (N_7298,N_2572,N_1030);
or U7299 (N_7299,N_3677,N_2087);
or U7300 (N_7300,N_2880,N_1361);
and U7301 (N_7301,N_4568,N_4177);
and U7302 (N_7302,N_2661,N_500);
and U7303 (N_7303,N_3741,N_774);
xor U7304 (N_7304,N_1584,N_1696);
xor U7305 (N_7305,N_2266,N_3655);
or U7306 (N_7306,N_2278,N_4846);
nor U7307 (N_7307,N_3257,N_1443);
or U7308 (N_7308,N_4449,N_2182);
nor U7309 (N_7309,N_80,N_3445);
and U7310 (N_7310,N_4676,N_1313);
and U7311 (N_7311,N_283,N_1412);
nor U7312 (N_7312,N_840,N_1193);
or U7313 (N_7313,N_1856,N_3955);
and U7314 (N_7314,N_4428,N_2067);
or U7315 (N_7315,N_3188,N_1686);
nor U7316 (N_7316,N_1411,N_551);
or U7317 (N_7317,N_1083,N_4825);
and U7318 (N_7318,N_783,N_1602);
nand U7319 (N_7319,N_152,N_2010);
and U7320 (N_7320,N_3833,N_934);
nand U7321 (N_7321,N_2007,N_3941);
or U7322 (N_7322,N_1329,N_3215);
nor U7323 (N_7323,N_1216,N_3547);
nor U7324 (N_7324,N_4338,N_2822);
xnor U7325 (N_7325,N_1232,N_897);
and U7326 (N_7326,N_2842,N_2263);
and U7327 (N_7327,N_3129,N_4935);
nand U7328 (N_7328,N_4480,N_2397);
nor U7329 (N_7329,N_4970,N_4384);
nor U7330 (N_7330,N_3503,N_2224);
nand U7331 (N_7331,N_4098,N_998);
and U7332 (N_7332,N_2333,N_4228);
or U7333 (N_7333,N_182,N_3964);
xnor U7334 (N_7334,N_2523,N_1731);
and U7335 (N_7335,N_2373,N_1984);
nand U7336 (N_7336,N_2524,N_4554);
nor U7337 (N_7337,N_4511,N_901);
nand U7338 (N_7338,N_1401,N_4417);
or U7339 (N_7339,N_4841,N_3426);
and U7340 (N_7340,N_439,N_4212);
or U7341 (N_7341,N_1503,N_1263);
and U7342 (N_7342,N_4128,N_144);
nor U7343 (N_7343,N_3277,N_180);
nand U7344 (N_7344,N_2038,N_4720);
nand U7345 (N_7345,N_2411,N_2910);
nand U7346 (N_7346,N_2674,N_2813);
or U7347 (N_7347,N_2165,N_3748);
and U7348 (N_7348,N_3812,N_1424);
nor U7349 (N_7349,N_1790,N_2172);
and U7350 (N_7350,N_2685,N_4222);
and U7351 (N_7351,N_905,N_2540);
nand U7352 (N_7352,N_3536,N_1847);
nand U7353 (N_7353,N_3970,N_4395);
and U7354 (N_7354,N_315,N_3030);
or U7355 (N_7355,N_298,N_3981);
or U7356 (N_7356,N_1683,N_591);
nand U7357 (N_7357,N_4487,N_3299);
nand U7358 (N_7358,N_359,N_3646);
xor U7359 (N_7359,N_2538,N_1593);
nand U7360 (N_7360,N_4550,N_3991);
and U7361 (N_7361,N_747,N_4429);
and U7362 (N_7362,N_1017,N_2924);
and U7363 (N_7363,N_2016,N_4729);
and U7364 (N_7364,N_2596,N_3000);
or U7365 (N_7365,N_1548,N_4937);
and U7366 (N_7366,N_4116,N_2705);
nand U7367 (N_7367,N_3803,N_334);
and U7368 (N_7368,N_3397,N_2855);
or U7369 (N_7369,N_465,N_2064);
or U7370 (N_7370,N_3029,N_1048);
or U7371 (N_7371,N_3295,N_4736);
or U7372 (N_7372,N_4191,N_4779);
and U7373 (N_7373,N_816,N_2625);
nor U7374 (N_7374,N_2139,N_121);
or U7375 (N_7375,N_131,N_384);
or U7376 (N_7376,N_883,N_2620);
nand U7377 (N_7377,N_1464,N_2011);
nand U7378 (N_7378,N_1573,N_2587);
and U7379 (N_7379,N_2808,N_3253);
nor U7380 (N_7380,N_3317,N_1933);
nand U7381 (N_7381,N_4467,N_3804);
nand U7382 (N_7382,N_1802,N_191);
and U7383 (N_7383,N_2043,N_1252);
or U7384 (N_7384,N_1980,N_2980);
or U7385 (N_7385,N_2287,N_4010);
and U7386 (N_7386,N_3161,N_979);
nor U7387 (N_7387,N_1654,N_2500);
nand U7388 (N_7388,N_742,N_4034);
and U7389 (N_7389,N_1812,N_3279);
and U7390 (N_7390,N_3590,N_4774);
or U7391 (N_7391,N_153,N_9);
nand U7392 (N_7392,N_1886,N_1879);
or U7393 (N_7393,N_2653,N_1810);
nor U7394 (N_7394,N_1908,N_924);
nor U7395 (N_7395,N_4908,N_2009);
nand U7396 (N_7396,N_2999,N_3746);
or U7397 (N_7397,N_1308,N_296);
or U7398 (N_7398,N_3039,N_2799);
and U7399 (N_7399,N_3120,N_1491);
and U7400 (N_7400,N_1130,N_3458);
and U7401 (N_7401,N_2762,N_478);
or U7402 (N_7402,N_4592,N_2728);
or U7403 (N_7403,N_1097,N_4052);
nor U7404 (N_7404,N_1581,N_4187);
or U7405 (N_7405,N_4674,N_431);
nand U7406 (N_7406,N_3251,N_2341);
or U7407 (N_7407,N_718,N_1875);
nand U7408 (N_7408,N_1801,N_2231);
nand U7409 (N_7409,N_4911,N_595);
nand U7410 (N_7410,N_722,N_347);
nor U7411 (N_7411,N_2797,N_1506);
or U7412 (N_7412,N_3168,N_4418);
and U7413 (N_7413,N_290,N_1343);
or U7414 (N_7414,N_1719,N_2122);
and U7415 (N_7415,N_54,N_4106);
nor U7416 (N_7416,N_256,N_1028);
or U7417 (N_7417,N_1025,N_2551);
and U7418 (N_7418,N_3923,N_4107);
nor U7419 (N_7419,N_1532,N_1807);
nor U7420 (N_7420,N_3022,N_4287);
nor U7421 (N_7421,N_4289,N_2835);
and U7422 (N_7422,N_4121,N_4997);
nand U7423 (N_7423,N_3814,N_3252);
nor U7424 (N_7424,N_2699,N_4357);
or U7425 (N_7425,N_4371,N_1835);
nand U7426 (N_7426,N_3554,N_2233);
nand U7427 (N_7427,N_768,N_493);
or U7428 (N_7428,N_354,N_2482);
nand U7429 (N_7429,N_2757,N_2947);
and U7430 (N_7430,N_4115,N_867);
nand U7431 (N_7431,N_959,N_4565);
and U7432 (N_7432,N_864,N_168);
nor U7433 (N_7433,N_2662,N_3133);
nand U7434 (N_7434,N_1711,N_268);
nor U7435 (N_7435,N_2006,N_4472);
and U7436 (N_7436,N_4659,N_4692);
nor U7437 (N_7437,N_4512,N_2290);
and U7438 (N_7438,N_534,N_2881);
or U7439 (N_7439,N_3828,N_1432);
nand U7440 (N_7440,N_2573,N_2692);
nor U7441 (N_7441,N_2001,N_958);
nor U7442 (N_7442,N_100,N_3620);
nand U7443 (N_7443,N_4195,N_1527);
nand U7444 (N_7444,N_1679,N_926);
nand U7445 (N_7445,N_2711,N_2468);
or U7446 (N_7446,N_330,N_994);
nand U7447 (N_7447,N_1460,N_3500);
or U7448 (N_7448,N_502,N_1360);
nand U7449 (N_7449,N_1162,N_4740);
nor U7450 (N_7450,N_4795,N_3184);
or U7451 (N_7451,N_4025,N_4319);
nor U7452 (N_7452,N_4546,N_3887);
nand U7453 (N_7453,N_1128,N_1552);
nor U7454 (N_7454,N_4818,N_1706);
nand U7455 (N_7455,N_803,N_3559);
nor U7456 (N_7456,N_974,N_1118);
and U7457 (N_7457,N_3737,N_3861);
and U7458 (N_7458,N_2494,N_1462);
and U7459 (N_7459,N_1888,N_4410);
nand U7460 (N_7460,N_4951,N_1463);
or U7461 (N_7461,N_3211,N_3566);
xnor U7462 (N_7462,N_2406,N_3402);
nor U7463 (N_7463,N_3583,N_1786);
and U7464 (N_7464,N_2611,N_2885);
nand U7465 (N_7465,N_1053,N_1585);
and U7466 (N_7466,N_713,N_810);
nor U7467 (N_7467,N_3597,N_4045);
nor U7468 (N_7468,N_278,N_1289);
or U7469 (N_7469,N_2720,N_2527);
or U7470 (N_7470,N_750,N_407);
nand U7471 (N_7471,N_4895,N_3117);
and U7472 (N_7472,N_667,N_2977);
nor U7473 (N_7473,N_549,N_769);
and U7474 (N_7474,N_30,N_1669);
and U7475 (N_7475,N_245,N_782);
nor U7476 (N_7476,N_686,N_4619);
nor U7477 (N_7477,N_321,N_3593);
nand U7478 (N_7478,N_1466,N_3321);
nand U7479 (N_7479,N_2409,N_3647);
nand U7480 (N_7480,N_4382,N_681);
nand U7481 (N_7481,N_4209,N_2830);
and U7482 (N_7482,N_4080,N_775);
or U7483 (N_7483,N_4933,N_4260);
or U7484 (N_7484,N_1398,N_4794);
nor U7485 (N_7485,N_1004,N_3205);
or U7486 (N_7486,N_1494,N_161);
nor U7487 (N_7487,N_906,N_3982);
nand U7488 (N_7488,N_2565,N_154);
or U7489 (N_7489,N_140,N_592);
nand U7490 (N_7490,N_4548,N_2465);
nand U7491 (N_7491,N_129,N_1500);
nor U7492 (N_7492,N_3546,N_2582);
nor U7493 (N_7493,N_1341,N_3520);
or U7494 (N_7494,N_1379,N_1174);
nand U7495 (N_7495,N_3019,N_4332);
nor U7496 (N_7496,N_2918,N_2747);
and U7497 (N_7497,N_3214,N_476);
nand U7498 (N_7498,N_4424,N_2605);
and U7499 (N_7499,N_1625,N_1404);
and U7500 (N_7500,N_2462,N_4970);
nand U7501 (N_7501,N_3629,N_3944);
nand U7502 (N_7502,N_3798,N_4036);
nand U7503 (N_7503,N_3736,N_4236);
and U7504 (N_7504,N_1208,N_4911);
nor U7505 (N_7505,N_410,N_3125);
and U7506 (N_7506,N_4251,N_544);
nor U7507 (N_7507,N_1946,N_1650);
and U7508 (N_7508,N_385,N_4768);
nor U7509 (N_7509,N_3135,N_3650);
nor U7510 (N_7510,N_1047,N_1902);
nor U7511 (N_7511,N_3910,N_4078);
nand U7512 (N_7512,N_308,N_4318);
or U7513 (N_7513,N_1378,N_3430);
nand U7514 (N_7514,N_4110,N_349);
or U7515 (N_7515,N_1452,N_1773);
or U7516 (N_7516,N_3442,N_2280);
and U7517 (N_7517,N_3057,N_4584);
or U7518 (N_7518,N_1450,N_1463);
and U7519 (N_7519,N_205,N_4157);
or U7520 (N_7520,N_2175,N_1658);
and U7521 (N_7521,N_4030,N_119);
nor U7522 (N_7522,N_4411,N_3508);
or U7523 (N_7523,N_2007,N_3285);
and U7524 (N_7524,N_4426,N_4687);
and U7525 (N_7525,N_316,N_4635);
nand U7526 (N_7526,N_2702,N_1752);
xnor U7527 (N_7527,N_4098,N_611);
or U7528 (N_7528,N_795,N_3589);
nor U7529 (N_7529,N_1829,N_625);
nand U7530 (N_7530,N_4149,N_3293);
nor U7531 (N_7531,N_4854,N_4741);
nand U7532 (N_7532,N_4866,N_3096);
nand U7533 (N_7533,N_1904,N_2442);
nand U7534 (N_7534,N_2569,N_4956);
and U7535 (N_7535,N_2509,N_1938);
nor U7536 (N_7536,N_1687,N_301);
or U7537 (N_7537,N_1930,N_4225);
nor U7538 (N_7538,N_609,N_1170);
or U7539 (N_7539,N_797,N_3900);
or U7540 (N_7540,N_3165,N_3536);
nor U7541 (N_7541,N_3366,N_35);
nand U7542 (N_7542,N_4073,N_4993);
and U7543 (N_7543,N_2390,N_1355);
nand U7544 (N_7544,N_1681,N_780);
nor U7545 (N_7545,N_16,N_1902);
nand U7546 (N_7546,N_4287,N_665);
and U7547 (N_7547,N_4943,N_1138);
or U7548 (N_7548,N_3145,N_598);
or U7549 (N_7549,N_4605,N_939);
and U7550 (N_7550,N_4109,N_3371);
nor U7551 (N_7551,N_1574,N_1163);
nor U7552 (N_7552,N_4603,N_4940);
or U7553 (N_7553,N_3714,N_180);
nand U7554 (N_7554,N_109,N_4580);
xor U7555 (N_7555,N_2773,N_2604);
and U7556 (N_7556,N_4988,N_1980);
and U7557 (N_7557,N_1297,N_4508);
and U7558 (N_7558,N_1226,N_3505);
nor U7559 (N_7559,N_3108,N_2155);
nor U7560 (N_7560,N_664,N_4932);
nor U7561 (N_7561,N_4878,N_917);
nor U7562 (N_7562,N_2098,N_4444);
and U7563 (N_7563,N_4832,N_1769);
nor U7564 (N_7564,N_1629,N_2567);
nor U7565 (N_7565,N_1884,N_3392);
nand U7566 (N_7566,N_2277,N_1143);
nand U7567 (N_7567,N_2568,N_4364);
nand U7568 (N_7568,N_3081,N_4078);
nor U7569 (N_7569,N_955,N_2384);
and U7570 (N_7570,N_2394,N_2928);
nand U7571 (N_7571,N_4175,N_955);
nand U7572 (N_7572,N_4027,N_3548);
and U7573 (N_7573,N_4397,N_2557);
and U7574 (N_7574,N_4607,N_4242);
and U7575 (N_7575,N_937,N_4192);
nand U7576 (N_7576,N_3892,N_3274);
nand U7577 (N_7577,N_118,N_3068);
and U7578 (N_7578,N_1032,N_3078);
and U7579 (N_7579,N_657,N_1712);
nor U7580 (N_7580,N_1487,N_1121);
and U7581 (N_7581,N_1334,N_2574);
nor U7582 (N_7582,N_4784,N_2199);
nand U7583 (N_7583,N_2300,N_4049);
nor U7584 (N_7584,N_2659,N_3777);
or U7585 (N_7585,N_3915,N_2723);
nand U7586 (N_7586,N_1597,N_3027);
nor U7587 (N_7587,N_2568,N_3978);
or U7588 (N_7588,N_3017,N_2579);
nor U7589 (N_7589,N_1306,N_4407);
and U7590 (N_7590,N_3888,N_968);
and U7591 (N_7591,N_174,N_111);
nand U7592 (N_7592,N_3313,N_780);
nor U7593 (N_7593,N_3669,N_3019);
nor U7594 (N_7594,N_191,N_273);
nor U7595 (N_7595,N_741,N_2273);
or U7596 (N_7596,N_4389,N_3915);
or U7597 (N_7597,N_1720,N_4416);
and U7598 (N_7598,N_4602,N_372);
nand U7599 (N_7599,N_338,N_1195);
nor U7600 (N_7600,N_4836,N_623);
nand U7601 (N_7601,N_3594,N_4761);
and U7602 (N_7602,N_2087,N_708);
and U7603 (N_7603,N_3089,N_4556);
or U7604 (N_7604,N_2830,N_2082);
xor U7605 (N_7605,N_848,N_2577);
or U7606 (N_7606,N_3297,N_1531);
nor U7607 (N_7607,N_2759,N_3608);
nand U7608 (N_7608,N_2328,N_3710);
nand U7609 (N_7609,N_2340,N_2181);
and U7610 (N_7610,N_873,N_4354);
nor U7611 (N_7611,N_1881,N_784);
nand U7612 (N_7612,N_1097,N_3159);
nor U7613 (N_7613,N_1361,N_2087);
nor U7614 (N_7614,N_3527,N_4561);
and U7615 (N_7615,N_2894,N_1977);
and U7616 (N_7616,N_3617,N_1300);
nand U7617 (N_7617,N_4664,N_4114);
or U7618 (N_7618,N_2097,N_4341);
nand U7619 (N_7619,N_324,N_2255);
nand U7620 (N_7620,N_2153,N_198);
nor U7621 (N_7621,N_2841,N_2732);
nor U7622 (N_7622,N_1909,N_2939);
nand U7623 (N_7623,N_2535,N_2476);
nand U7624 (N_7624,N_2049,N_2586);
or U7625 (N_7625,N_4944,N_3471);
and U7626 (N_7626,N_1596,N_1663);
nand U7627 (N_7627,N_1849,N_3870);
nor U7628 (N_7628,N_1147,N_2418);
nor U7629 (N_7629,N_4496,N_688);
and U7630 (N_7630,N_3353,N_4252);
nand U7631 (N_7631,N_600,N_2887);
and U7632 (N_7632,N_346,N_2545);
or U7633 (N_7633,N_1394,N_1971);
nand U7634 (N_7634,N_4507,N_2339);
xnor U7635 (N_7635,N_3058,N_1266);
or U7636 (N_7636,N_663,N_325);
nand U7637 (N_7637,N_4397,N_4378);
nor U7638 (N_7638,N_49,N_2631);
nor U7639 (N_7639,N_4810,N_4633);
and U7640 (N_7640,N_2376,N_2628);
nand U7641 (N_7641,N_2969,N_2100);
and U7642 (N_7642,N_3987,N_3080);
or U7643 (N_7643,N_589,N_1647);
nand U7644 (N_7644,N_873,N_1113);
nand U7645 (N_7645,N_2060,N_2710);
or U7646 (N_7646,N_1601,N_1998);
nor U7647 (N_7647,N_2896,N_447);
nand U7648 (N_7648,N_4358,N_1719);
and U7649 (N_7649,N_1258,N_4975);
nor U7650 (N_7650,N_672,N_4773);
nand U7651 (N_7651,N_3856,N_2920);
or U7652 (N_7652,N_1543,N_3463);
and U7653 (N_7653,N_3776,N_3250);
or U7654 (N_7654,N_1009,N_3399);
and U7655 (N_7655,N_3049,N_2024);
or U7656 (N_7656,N_352,N_2641);
or U7657 (N_7657,N_2980,N_2790);
nand U7658 (N_7658,N_1682,N_202);
nor U7659 (N_7659,N_4774,N_1366);
nand U7660 (N_7660,N_2679,N_3120);
and U7661 (N_7661,N_2200,N_4724);
nor U7662 (N_7662,N_74,N_2229);
nor U7663 (N_7663,N_2364,N_1229);
nand U7664 (N_7664,N_2398,N_2665);
and U7665 (N_7665,N_1700,N_2554);
and U7666 (N_7666,N_495,N_2557);
nor U7667 (N_7667,N_1020,N_1760);
nand U7668 (N_7668,N_741,N_2684);
nand U7669 (N_7669,N_3392,N_1095);
or U7670 (N_7670,N_4154,N_1771);
nor U7671 (N_7671,N_459,N_4423);
and U7672 (N_7672,N_4489,N_2781);
nand U7673 (N_7673,N_2443,N_3114);
nor U7674 (N_7674,N_2447,N_944);
nor U7675 (N_7675,N_1318,N_1522);
nor U7676 (N_7676,N_2123,N_686);
nand U7677 (N_7677,N_2081,N_577);
or U7678 (N_7678,N_3382,N_122);
nor U7679 (N_7679,N_4229,N_2799);
nand U7680 (N_7680,N_4759,N_4928);
or U7681 (N_7681,N_4551,N_2198);
nor U7682 (N_7682,N_568,N_2121);
and U7683 (N_7683,N_2326,N_4489);
and U7684 (N_7684,N_82,N_3159);
nand U7685 (N_7685,N_1877,N_3250);
nand U7686 (N_7686,N_617,N_3226);
nand U7687 (N_7687,N_2593,N_4785);
and U7688 (N_7688,N_3660,N_421);
nor U7689 (N_7689,N_4328,N_827);
and U7690 (N_7690,N_2419,N_1584);
and U7691 (N_7691,N_1727,N_3482);
nand U7692 (N_7692,N_2543,N_834);
nand U7693 (N_7693,N_336,N_3408);
and U7694 (N_7694,N_3957,N_114);
or U7695 (N_7695,N_971,N_1773);
nor U7696 (N_7696,N_4309,N_2185);
nand U7697 (N_7697,N_2090,N_4035);
or U7698 (N_7698,N_4108,N_4300);
nor U7699 (N_7699,N_656,N_2348);
nor U7700 (N_7700,N_4952,N_3160);
and U7701 (N_7701,N_4086,N_3222);
nor U7702 (N_7702,N_1957,N_2810);
and U7703 (N_7703,N_2242,N_1311);
and U7704 (N_7704,N_552,N_1810);
or U7705 (N_7705,N_280,N_306);
nor U7706 (N_7706,N_2186,N_3099);
and U7707 (N_7707,N_92,N_25);
nor U7708 (N_7708,N_1643,N_2966);
or U7709 (N_7709,N_3271,N_2520);
nand U7710 (N_7710,N_1913,N_4688);
or U7711 (N_7711,N_1000,N_3749);
or U7712 (N_7712,N_2419,N_4153);
or U7713 (N_7713,N_53,N_3451);
and U7714 (N_7714,N_3074,N_2110);
and U7715 (N_7715,N_2143,N_126);
or U7716 (N_7716,N_1696,N_2566);
xnor U7717 (N_7717,N_1503,N_664);
or U7718 (N_7718,N_4597,N_2176);
and U7719 (N_7719,N_3576,N_3945);
and U7720 (N_7720,N_4349,N_3581);
and U7721 (N_7721,N_2157,N_3284);
nor U7722 (N_7722,N_2829,N_1527);
and U7723 (N_7723,N_103,N_822);
nor U7724 (N_7724,N_1790,N_3023);
and U7725 (N_7725,N_3974,N_1483);
nand U7726 (N_7726,N_3072,N_4367);
nand U7727 (N_7727,N_3610,N_1474);
nand U7728 (N_7728,N_3636,N_4459);
and U7729 (N_7729,N_648,N_4610);
and U7730 (N_7730,N_4304,N_2774);
or U7731 (N_7731,N_1118,N_2674);
nand U7732 (N_7732,N_1953,N_4270);
or U7733 (N_7733,N_334,N_4139);
nor U7734 (N_7734,N_741,N_2255);
and U7735 (N_7735,N_3621,N_4883);
and U7736 (N_7736,N_609,N_4794);
and U7737 (N_7737,N_4581,N_2385);
nor U7738 (N_7738,N_590,N_2670);
nand U7739 (N_7739,N_2800,N_2556);
nand U7740 (N_7740,N_3602,N_1804);
or U7741 (N_7741,N_2120,N_2149);
nand U7742 (N_7742,N_2067,N_2903);
nand U7743 (N_7743,N_4693,N_36);
nand U7744 (N_7744,N_207,N_2563);
and U7745 (N_7745,N_1857,N_4935);
nand U7746 (N_7746,N_4626,N_2601);
nor U7747 (N_7747,N_2158,N_151);
nor U7748 (N_7748,N_1113,N_2628);
nand U7749 (N_7749,N_1374,N_2672);
and U7750 (N_7750,N_1320,N_3927);
nand U7751 (N_7751,N_2999,N_3608);
nor U7752 (N_7752,N_4571,N_1385);
or U7753 (N_7753,N_3976,N_1807);
nor U7754 (N_7754,N_537,N_1462);
and U7755 (N_7755,N_4871,N_397);
nand U7756 (N_7756,N_4893,N_3359);
nand U7757 (N_7757,N_1688,N_2208);
and U7758 (N_7758,N_3503,N_4977);
and U7759 (N_7759,N_379,N_2949);
nand U7760 (N_7760,N_3405,N_20);
nor U7761 (N_7761,N_3140,N_3917);
and U7762 (N_7762,N_2690,N_3259);
nor U7763 (N_7763,N_4367,N_371);
nor U7764 (N_7764,N_2077,N_4315);
or U7765 (N_7765,N_3341,N_567);
nor U7766 (N_7766,N_269,N_1955);
or U7767 (N_7767,N_4794,N_4474);
nand U7768 (N_7768,N_4682,N_1435);
nand U7769 (N_7769,N_4332,N_2392);
nand U7770 (N_7770,N_286,N_3853);
nor U7771 (N_7771,N_802,N_3183);
and U7772 (N_7772,N_4117,N_1617);
nand U7773 (N_7773,N_2120,N_2497);
or U7774 (N_7774,N_2037,N_1867);
and U7775 (N_7775,N_2486,N_1109);
or U7776 (N_7776,N_1264,N_3078);
and U7777 (N_7777,N_4921,N_3297);
or U7778 (N_7778,N_3933,N_1551);
nor U7779 (N_7779,N_2595,N_195);
nor U7780 (N_7780,N_4942,N_2326);
nor U7781 (N_7781,N_1866,N_506);
or U7782 (N_7782,N_4596,N_882);
nand U7783 (N_7783,N_3409,N_991);
nand U7784 (N_7784,N_854,N_4922);
nor U7785 (N_7785,N_1202,N_110);
and U7786 (N_7786,N_1957,N_2531);
or U7787 (N_7787,N_4767,N_742);
or U7788 (N_7788,N_2270,N_1521);
nand U7789 (N_7789,N_937,N_2194);
nor U7790 (N_7790,N_2658,N_154);
nor U7791 (N_7791,N_1687,N_1536);
nor U7792 (N_7792,N_676,N_2063);
and U7793 (N_7793,N_551,N_682);
and U7794 (N_7794,N_3450,N_2992);
and U7795 (N_7795,N_3242,N_1279);
nand U7796 (N_7796,N_1771,N_126);
nand U7797 (N_7797,N_495,N_3656);
or U7798 (N_7798,N_1157,N_4439);
and U7799 (N_7799,N_2029,N_3399);
or U7800 (N_7800,N_1204,N_3338);
nand U7801 (N_7801,N_3726,N_4287);
nor U7802 (N_7802,N_2504,N_2497);
and U7803 (N_7803,N_1730,N_3960);
nor U7804 (N_7804,N_3057,N_583);
nor U7805 (N_7805,N_258,N_381);
or U7806 (N_7806,N_1038,N_4396);
or U7807 (N_7807,N_3643,N_2521);
or U7808 (N_7808,N_2049,N_567);
nand U7809 (N_7809,N_2266,N_2370);
and U7810 (N_7810,N_855,N_1741);
or U7811 (N_7811,N_4371,N_4987);
and U7812 (N_7812,N_4975,N_2522);
or U7813 (N_7813,N_1629,N_708);
and U7814 (N_7814,N_4768,N_762);
or U7815 (N_7815,N_634,N_1203);
nand U7816 (N_7816,N_1232,N_692);
nor U7817 (N_7817,N_1,N_439);
nor U7818 (N_7818,N_2811,N_1251);
nor U7819 (N_7819,N_108,N_2086);
or U7820 (N_7820,N_3957,N_1914);
and U7821 (N_7821,N_3830,N_2173);
nor U7822 (N_7822,N_4811,N_1421);
nand U7823 (N_7823,N_1746,N_239);
nand U7824 (N_7824,N_4703,N_1805);
nor U7825 (N_7825,N_1668,N_1580);
and U7826 (N_7826,N_2331,N_637);
nor U7827 (N_7827,N_200,N_1154);
and U7828 (N_7828,N_4613,N_1129);
nand U7829 (N_7829,N_1159,N_3520);
nand U7830 (N_7830,N_2009,N_2644);
nor U7831 (N_7831,N_2035,N_519);
and U7832 (N_7832,N_591,N_4295);
or U7833 (N_7833,N_3989,N_4487);
or U7834 (N_7834,N_1545,N_4641);
nor U7835 (N_7835,N_2605,N_345);
nand U7836 (N_7836,N_540,N_3080);
and U7837 (N_7837,N_3724,N_2358);
and U7838 (N_7838,N_1935,N_2637);
and U7839 (N_7839,N_3135,N_857);
nor U7840 (N_7840,N_859,N_4141);
and U7841 (N_7841,N_4002,N_584);
nor U7842 (N_7842,N_1733,N_514);
or U7843 (N_7843,N_2379,N_2694);
or U7844 (N_7844,N_2151,N_4568);
and U7845 (N_7845,N_529,N_734);
nor U7846 (N_7846,N_704,N_4500);
or U7847 (N_7847,N_2232,N_4284);
nor U7848 (N_7848,N_3812,N_1598);
nor U7849 (N_7849,N_1106,N_1926);
and U7850 (N_7850,N_4982,N_2274);
or U7851 (N_7851,N_3675,N_2061);
and U7852 (N_7852,N_2424,N_914);
or U7853 (N_7853,N_34,N_1110);
and U7854 (N_7854,N_3395,N_3689);
and U7855 (N_7855,N_1727,N_4527);
nor U7856 (N_7856,N_1101,N_932);
or U7857 (N_7857,N_673,N_1213);
nor U7858 (N_7858,N_4489,N_835);
nor U7859 (N_7859,N_3320,N_308);
or U7860 (N_7860,N_2039,N_3991);
and U7861 (N_7861,N_3962,N_2600);
and U7862 (N_7862,N_3014,N_2688);
nand U7863 (N_7863,N_3303,N_228);
nand U7864 (N_7864,N_3604,N_3704);
or U7865 (N_7865,N_424,N_3816);
xor U7866 (N_7866,N_1991,N_3009);
nor U7867 (N_7867,N_3200,N_563);
nor U7868 (N_7868,N_1365,N_1149);
or U7869 (N_7869,N_1292,N_1629);
nand U7870 (N_7870,N_1146,N_3956);
nand U7871 (N_7871,N_1328,N_2567);
nand U7872 (N_7872,N_3224,N_4593);
or U7873 (N_7873,N_4215,N_579);
and U7874 (N_7874,N_650,N_195);
nor U7875 (N_7875,N_1045,N_4419);
nor U7876 (N_7876,N_2111,N_3378);
or U7877 (N_7877,N_4060,N_2528);
and U7878 (N_7878,N_2703,N_3770);
nor U7879 (N_7879,N_591,N_2931);
nand U7880 (N_7880,N_3710,N_1854);
and U7881 (N_7881,N_1607,N_2769);
nor U7882 (N_7882,N_360,N_3819);
or U7883 (N_7883,N_874,N_2999);
nand U7884 (N_7884,N_1728,N_3458);
or U7885 (N_7885,N_3173,N_483);
or U7886 (N_7886,N_4302,N_3030);
nand U7887 (N_7887,N_2927,N_1106);
and U7888 (N_7888,N_602,N_1464);
and U7889 (N_7889,N_1439,N_2085);
nand U7890 (N_7890,N_3984,N_3495);
nor U7891 (N_7891,N_2959,N_2685);
and U7892 (N_7892,N_2853,N_3231);
and U7893 (N_7893,N_2705,N_1949);
and U7894 (N_7894,N_3760,N_4075);
or U7895 (N_7895,N_2107,N_4604);
and U7896 (N_7896,N_3037,N_3555);
and U7897 (N_7897,N_1910,N_2355);
or U7898 (N_7898,N_3008,N_4296);
and U7899 (N_7899,N_3181,N_4505);
nor U7900 (N_7900,N_3724,N_3136);
nand U7901 (N_7901,N_981,N_2992);
nor U7902 (N_7902,N_1331,N_3690);
nor U7903 (N_7903,N_3819,N_1090);
nor U7904 (N_7904,N_3898,N_2493);
or U7905 (N_7905,N_739,N_1515);
or U7906 (N_7906,N_4270,N_2379);
and U7907 (N_7907,N_152,N_2313);
nor U7908 (N_7908,N_2002,N_2561);
nand U7909 (N_7909,N_4712,N_4497);
nor U7910 (N_7910,N_4703,N_947);
nand U7911 (N_7911,N_4531,N_4409);
nor U7912 (N_7912,N_3908,N_428);
nor U7913 (N_7913,N_2291,N_833);
nand U7914 (N_7914,N_4488,N_596);
nor U7915 (N_7915,N_3252,N_4044);
nand U7916 (N_7916,N_2372,N_2456);
nand U7917 (N_7917,N_2889,N_4793);
or U7918 (N_7918,N_1050,N_3347);
or U7919 (N_7919,N_458,N_4703);
nand U7920 (N_7920,N_3610,N_2637);
nor U7921 (N_7921,N_2815,N_4639);
nor U7922 (N_7922,N_2337,N_4107);
nor U7923 (N_7923,N_4069,N_2034);
nand U7924 (N_7924,N_2177,N_1744);
or U7925 (N_7925,N_4811,N_171);
or U7926 (N_7926,N_1900,N_3075);
or U7927 (N_7927,N_1312,N_2831);
or U7928 (N_7928,N_2076,N_816);
and U7929 (N_7929,N_4089,N_456);
nor U7930 (N_7930,N_4860,N_4586);
nor U7931 (N_7931,N_1653,N_1175);
nor U7932 (N_7932,N_4754,N_4710);
nand U7933 (N_7933,N_4114,N_3242);
and U7934 (N_7934,N_1330,N_3076);
and U7935 (N_7935,N_360,N_3930);
and U7936 (N_7936,N_2680,N_1780);
nor U7937 (N_7937,N_1040,N_3481);
or U7938 (N_7938,N_3047,N_1444);
and U7939 (N_7939,N_1370,N_1718);
nand U7940 (N_7940,N_3595,N_1505);
nor U7941 (N_7941,N_3950,N_4590);
nand U7942 (N_7942,N_2839,N_709);
or U7943 (N_7943,N_3461,N_3329);
or U7944 (N_7944,N_4313,N_3046);
and U7945 (N_7945,N_4614,N_1559);
nor U7946 (N_7946,N_912,N_1452);
nand U7947 (N_7947,N_4403,N_4108);
nand U7948 (N_7948,N_2398,N_3975);
or U7949 (N_7949,N_144,N_4122);
or U7950 (N_7950,N_1223,N_4042);
nand U7951 (N_7951,N_884,N_1430);
and U7952 (N_7952,N_1365,N_3797);
or U7953 (N_7953,N_132,N_2537);
nor U7954 (N_7954,N_4121,N_4674);
and U7955 (N_7955,N_3773,N_2231);
or U7956 (N_7956,N_2310,N_3389);
or U7957 (N_7957,N_4802,N_2238);
nor U7958 (N_7958,N_4827,N_3159);
nor U7959 (N_7959,N_2458,N_90);
nor U7960 (N_7960,N_1154,N_459);
and U7961 (N_7961,N_192,N_4672);
or U7962 (N_7962,N_2799,N_1325);
nor U7963 (N_7963,N_2874,N_4712);
nand U7964 (N_7964,N_4911,N_3054);
or U7965 (N_7965,N_4424,N_3629);
or U7966 (N_7966,N_1004,N_2492);
nand U7967 (N_7967,N_1196,N_1738);
or U7968 (N_7968,N_3900,N_2522);
nor U7969 (N_7969,N_4707,N_542);
and U7970 (N_7970,N_4274,N_1556);
or U7971 (N_7971,N_1723,N_2437);
and U7972 (N_7972,N_3365,N_2689);
and U7973 (N_7973,N_3662,N_804);
and U7974 (N_7974,N_4238,N_3661);
nand U7975 (N_7975,N_4399,N_1405);
nor U7976 (N_7976,N_3166,N_1047);
and U7977 (N_7977,N_1559,N_367);
or U7978 (N_7978,N_2258,N_3799);
nand U7979 (N_7979,N_2468,N_3029);
or U7980 (N_7980,N_4455,N_4759);
nor U7981 (N_7981,N_3340,N_2237);
nor U7982 (N_7982,N_1328,N_922);
nand U7983 (N_7983,N_1403,N_4004);
or U7984 (N_7984,N_4147,N_3163);
or U7985 (N_7985,N_4100,N_3801);
and U7986 (N_7986,N_4535,N_1838);
or U7987 (N_7987,N_1603,N_3816);
nand U7988 (N_7988,N_3570,N_2264);
and U7989 (N_7989,N_1496,N_1203);
and U7990 (N_7990,N_1148,N_1068);
nor U7991 (N_7991,N_404,N_1663);
nor U7992 (N_7992,N_3724,N_3198);
nor U7993 (N_7993,N_958,N_58);
nor U7994 (N_7994,N_3900,N_3907);
nand U7995 (N_7995,N_405,N_941);
nor U7996 (N_7996,N_4049,N_3896);
and U7997 (N_7997,N_1636,N_3650);
nor U7998 (N_7998,N_686,N_3140);
nor U7999 (N_7999,N_1114,N_3466);
nand U8000 (N_8000,N_2385,N_2296);
and U8001 (N_8001,N_1290,N_2596);
and U8002 (N_8002,N_4618,N_4781);
nor U8003 (N_8003,N_1259,N_4762);
and U8004 (N_8004,N_2029,N_815);
nor U8005 (N_8005,N_814,N_4403);
and U8006 (N_8006,N_4569,N_3149);
or U8007 (N_8007,N_309,N_4839);
nor U8008 (N_8008,N_939,N_3814);
nand U8009 (N_8009,N_1904,N_496);
nand U8010 (N_8010,N_2393,N_1829);
and U8011 (N_8011,N_290,N_1294);
nand U8012 (N_8012,N_2030,N_3696);
nor U8013 (N_8013,N_624,N_5);
nor U8014 (N_8014,N_1886,N_800);
nor U8015 (N_8015,N_4059,N_2924);
nor U8016 (N_8016,N_3359,N_2480);
nand U8017 (N_8017,N_4001,N_4945);
or U8018 (N_8018,N_4206,N_383);
nor U8019 (N_8019,N_3326,N_1662);
and U8020 (N_8020,N_1684,N_748);
and U8021 (N_8021,N_123,N_2668);
or U8022 (N_8022,N_3175,N_4675);
and U8023 (N_8023,N_155,N_1340);
and U8024 (N_8024,N_2227,N_3689);
and U8025 (N_8025,N_3241,N_2647);
or U8026 (N_8026,N_2091,N_3279);
or U8027 (N_8027,N_43,N_2777);
nor U8028 (N_8028,N_1593,N_3238);
or U8029 (N_8029,N_4186,N_2361);
or U8030 (N_8030,N_3900,N_826);
and U8031 (N_8031,N_489,N_1498);
and U8032 (N_8032,N_1837,N_1946);
nand U8033 (N_8033,N_2604,N_3875);
nand U8034 (N_8034,N_190,N_3493);
nand U8035 (N_8035,N_4027,N_2889);
nor U8036 (N_8036,N_389,N_3231);
nand U8037 (N_8037,N_4283,N_3363);
nand U8038 (N_8038,N_288,N_1832);
and U8039 (N_8039,N_2274,N_4139);
nor U8040 (N_8040,N_4203,N_4444);
and U8041 (N_8041,N_2947,N_1413);
nand U8042 (N_8042,N_4330,N_366);
and U8043 (N_8043,N_2863,N_2395);
nand U8044 (N_8044,N_913,N_3076);
and U8045 (N_8045,N_3775,N_2505);
or U8046 (N_8046,N_1775,N_4014);
and U8047 (N_8047,N_2257,N_580);
nor U8048 (N_8048,N_3004,N_217);
or U8049 (N_8049,N_2899,N_89);
nand U8050 (N_8050,N_2009,N_2404);
and U8051 (N_8051,N_2045,N_2721);
nor U8052 (N_8052,N_615,N_2831);
or U8053 (N_8053,N_1427,N_1348);
nor U8054 (N_8054,N_4237,N_4955);
and U8055 (N_8055,N_4942,N_95);
or U8056 (N_8056,N_915,N_2160);
nand U8057 (N_8057,N_3200,N_4179);
or U8058 (N_8058,N_757,N_3346);
and U8059 (N_8059,N_2224,N_3369);
or U8060 (N_8060,N_2839,N_2402);
nor U8061 (N_8061,N_3210,N_1276);
and U8062 (N_8062,N_4420,N_2345);
or U8063 (N_8063,N_490,N_3812);
and U8064 (N_8064,N_1818,N_235);
nand U8065 (N_8065,N_2179,N_3082);
nand U8066 (N_8066,N_4761,N_2725);
or U8067 (N_8067,N_342,N_951);
nor U8068 (N_8068,N_285,N_4934);
nand U8069 (N_8069,N_914,N_695);
and U8070 (N_8070,N_4635,N_1973);
nand U8071 (N_8071,N_1906,N_448);
and U8072 (N_8072,N_2341,N_3318);
nor U8073 (N_8073,N_2019,N_3927);
nand U8074 (N_8074,N_367,N_1782);
or U8075 (N_8075,N_554,N_3493);
nor U8076 (N_8076,N_1058,N_2735);
or U8077 (N_8077,N_1830,N_4835);
and U8078 (N_8078,N_841,N_2323);
nand U8079 (N_8079,N_2855,N_2745);
or U8080 (N_8080,N_1871,N_2439);
nor U8081 (N_8081,N_1773,N_3960);
nor U8082 (N_8082,N_4097,N_2267);
nor U8083 (N_8083,N_1418,N_3402);
xnor U8084 (N_8084,N_4128,N_2270);
nor U8085 (N_8085,N_1757,N_3619);
or U8086 (N_8086,N_3870,N_4600);
nand U8087 (N_8087,N_3377,N_2554);
nand U8088 (N_8088,N_4289,N_2743);
or U8089 (N_8089,N_4272,N_147);
nand U8090 (N_8090,N_3968,N_870);
or U8091 (N_8091,N_161,N_4712);
or U8092 (N_8092,N_1388,N_2527);
nor U8093 (N_8093,N_3499,N_2661);
nor U8094 (N_8094,N_3546,N_3144);
or U8095 (N_8095,N_796,N_3943);
or U8096 (N_8096,N_2618,N_4260);
and U8097 (N_8097,N_3565,N_2285);
or U8098 (N_8098,N_1076,N_4277);
nand U8099 (N_8099,N_262,N_581);
or U8100 (N_8100,N_3633,N_0);
nand U8101 (N_8101,N_731,N_940);
nand U8102 (N_8102,N_2646,N_2675);
nand U8103 (N_8103,N_4876,N_1418);
or U8104 (N_8104,N_2409,N_3328);
nand U8105 (N_8105,N_4221,N_3240);
nand U8106 (N_8106,N_290,N_4655);
nor U8107 (N_8107,N_4937,N_3919);
or U8108 (N_8108,N_2388,N_1631);
nor U8109 (N_8109,N_1791,N_4726);
nand U8110 (N_8110,N_2701,N_744);
and U8111 (N_8111,N_573,N_2183);
and U8112 (N_8112,N_375,N_3893);
nand U8113 (N_8113,N_3513,N_4617);
nand U8114 (N_8114,N_2840,N_317);
nor U8115 (N_8115,N_1238,N_777);
and U8116 (N_8116,N_2165,N_4232);
nand U8117 (N_8117,N_2458,N_1064);
nand U8118 (N_8118,N_2680,N_3091);
or U8119 (N_8119,N_891,N_1219);
and U8120 (N_8120,N_3809,N_3008);
and U8121 (N_8121,N_4752,N_980);
nor U8122 (N_8122,N_2954,N_4357);
and U8123 (N_8123,N_938,N_3490);
xnor U8124 (N_8124,N_1579,N_1634);
and U8125 (N_8125,N_4040,N_3557);
nand U8126 (N_8126,N_2290,N_4666);
nand U8127 (N_8127,N_641,N_4232);
nand U8128 (N_8128,N_1298,N_2554);
or U8129 (N_8129,N_1117,N_1960);
nand U8130 (N_8130,N_700,N_762);
nand U8131 (N_8131,N_773,N_506);
nor U8132 (N_8132,N_4167,N_228);
nor U8133 (N_8133,N_320,N_769);
and U8134 (N_8134,N_2508,N_2378);
and U8135 (N_8135,N_3051,N_4953);
and U8136 (N_8136,N_3704,N_1077);
nand U8137 (N_8137,N_2779,N_2107);
nor U8138 (N_8138,N_342,N_3439);
nand U8139 (N_8139,N_3101,N_1337);
and U8140 (N_8140,N_2240,N_3081);
nor U8141 (N_8141,N_4696,N_943);
and U8142 (N_8142,N_2697,N_3019);
nor U8143 (N_8143,N_522,N_4795);
nand U8144 (N_8144,N_470,N_4620);
or U8145 (N_8145,N_1194,N_1219);
nor U8146 (N_8146,N_627,N_3689);
and U8147 (N_8147,N_2573,N_4537);
nor U8148 (N_8148,N_440,N_933);
nor U8149 (N_8149,N_553,N_1476);
and U8150 (N_8150,N_2814,N_307);
or U8151 (N_8151,N_4592,N_3167);
nor U8152 (N_8152,N_932,N_2147);
or U8153 (N_8153,N_4340,N_1376);
nand U8154 (N_8154,N_1968,N_4636);
nand U8155 (N_8155,N_1345,N_3286);
nand U8156 (N_8156,N_2009,N_4818);
nor U8157 (N_8157,N_1778,N_3194);
or U8158 (N_8158,N_2528,N_1083);
nor U8159 (N_8159,N_1237,N_4353);
nor U8160 (N_8160,N_2948,N_3814);
and U8161 (N_8161,N_3637,N_2201);
nand U8162 (N_8162,N_182,N_364);
nand U8163 (N_8163,N_953,N_623);
or U8164 (N_8164,N_4395,N_1707);
nor U8165 (N_8165,N_1283,N_292);
nor U8166 (N_8166,N_490,N_369);
or U8167 (N_8167,N_1181,N_1248);
and U8168 (N_8168,N_4445,N_1601);
nand U8169 (N_8169,N_4819,N_4250);
or U8170 (N_8170,N_645,N_4848);
nand U8171 (N_8171,N_2533,N_4863);
nor U8172 (N_8172,N_2460,N_3162);
nand U8173 (N_8173,N_4406,N_300);
nor U8174 (N_8174,N_3650,N_2894);
nor U8175 (N_8175,N_2090,N_4840);
nor U8176 (N_8176,N_1703,N_4754);
nor U8177 (N_8177,N_1638,N_4467);
and U8178 (N_8178,N_1627,N_1431);
and U8179 (N_8179,N_4237,N_1219);
and U8180 (N_8180,N_1183,N_578);
nand U8181 (N_8181,N_923,N_866);
or U8182 (N_8182,N_1287,N_2044);
nor U8183 (N_8183,N_3942,N_1002);
and U8184 (N_8184,N_3793,N_891);
nor U8185 (N_8185,N_4952,N_4640);
nand U8186 (N_8186,N_562,N_3105);
nor U8187 (N_8187,N_2861,N_2606);
nor U8188 (N_8188,N_3561,N_1832);
nor U8189 (N_8189,N_3832,N_3292);
nor U8190 (N_8190,N_1807,N_1505);
and U8191 (N_8191,N_2866,N_1438);
and U8192 (N_8192,N_2531,N_4117);
and U8193 (N_8193,N_912,N_2265);
and U8194 (N_8194,N_2929,N_4446);
xnor U8195 (N_8195,N_2048,N_1227);
nand U8196 (N_8196,N_4505,N_3546);
nand U8197 (N_8197,N_3191,N_3380);
nand U8198 (N_8198,N_222,N_3913);
nor U8199 (N_8199,N_2555,N_4810);
and U8200 (N_8200,N_3694,N_4283);
or U8201 (N_8201,N_2311,N_3255);
and U8202 (N_8202,N_894,N_1369);
or U8203 (N_8203,N_778,N_1361);
nand U8204 (N_8204,N_760,N_3387);
nor U8205 (N_8205,N_4544,N_3754);
or U8206 (N_8206,N_962,N_1841);
or U8207 (N_8207,N_3433,N_4670);
nand U8208 (N_8208,N_2414,N_3232);
and U8209 (N_8209,N_1239,N_401);
and U8210 (N_8210,N_222,N_1341);
or U8211 (N_8211,N_4234,N_3948);
xor U8212 (N_8212,N_595,N_1859);
or U8213 (N_8213,N_500,N_435);
and U8214 (N_8214,N_1378,N_1898);
and U8215 (N_8215,N_3239,N_1805);
and U8216 (N_8216,N_3582,N_2499);
and U8217 (N_8217,N_1765,N_4214);
nor U8218 (N_8218,N_1650,N_283);
nand U8219 (N_8219,N_4504,N_409);
or U8220 (N_8220,N_153,N_671);
nor U8221 (N_8221,N_3523,N_1727);
or U8222 (N_8222,N_3985,N_3913);
nand U8223 (N_8223,N_3060,N_4297);
or U8224 (N_8224,N_227,N_2311);
or U8225 (N_8225,N_1999,N_4567);
nor U8226 (N_8226,N_2968,N_1622);
nand U8227 (N_8227,N_1698,N_2730);
or U8228 (N_8228,N_3996,N_2474);
and U8229 (N_8229,N_99,N_2491);
and U8230 (N_8230,N_3156,N_2865);
nand U8231 (N_8231,N_1390,N_4928);
nor U8232 (N_8232,N_2073,N_3664);
nand U8233 (N_8233,N_4417,N_2011);
nor U8234 (N_8234,N_3788,N_2402);
nand U8235 (N_8235,N_1423,N_2656);
nor U8236 (N_8236,N_333,N_1099);
nand U8237 (N_8237,N_4499,N_649);
nor U8238 (N_8238,N_2009,N_4327);
or U8239 (N_8239,N_1675,N_42);
nand U8240 (N_8240,N_1241,N_412);
nor U8241 (N_8241,N_2601,N_3744);
or U8242 (N_8242,N_1495,N_1623);
nor U8243 (N_8243,N_215,N_1471);
nand U8244 (N_8244,N_174,N_365);
nor U8245 (N_8245,N_4468,N_1309);
nand U8246 (N_8246,N_625,N_1095);
or U8247 (N_8247,N_4647,N_4163);
and U8248 (N_8248,N_1642,N_4790);
nor U8249 (N_8249,N_1061,N_2503);
or U8250 (N_8250,N_4590,N_1311);
nand U8251 (N_8251,N_781,N_845);
nand U8252 (N_8252,N_4806,N_4084);
and U8253 (N_8253,N_1722,N_2309);
nor U8254 (N_8254,N_3335,N_2661);
nor U8255 (N_8255,N_1701,N_2288);
nor U8256 (N_8256,N_4645,N_793);
nor U8257 (N_8257,N_1347,N_3335);
or U8258 (N_8258,N_2084,N_1306);
nand U8259 (N_8259,N_2932,N_1486);
nand U8260 (N_8260,N_3546,N_243);
nand U8261 (N_8261,N_1286,N_4181);
nand U8262 (N_8262,N_3585,N_2464);
or U8263 (N_8263,N_2850,N_3401);
nand U8264 (N_8264,N_739,N_1403);
or U8265 (N_8265,N_4862,N_3434);
nor U8266 (N_8266,N_2094,N_2757);
nand U8267 (N_8267,N_152,N_821);
or U8268 (N_8268,N_3869,N_2289);
or U8269 (N_8269,N_152,N_2896);
and U8270 (N_8270,N_4002,N_683);
and U8271 (N_8271,N_3409,N_3530);
nor U8272 (N_8272,N_2293,N_4965);
or U8273 (N_8273,N_1062,N_426);
and U8274 (N_8274,N_3114,N_4737);
and U8275 (N_8275,N_713,N_4418);
nand U8276 (N_8276,N_4107,N_4145);
or U8277 (N_8277,N_4543,N_2956);
or U8278 (N_8278,N_3530,N_759);
or U8279 (N_8279,N_4458,N_2601);
and U8280 (N_8280,N_1680,N_4844);
nor U8281 (N_8281,N_155,N_2533);
nor U8282 (N_8282,N_1474,N_345);
or U8283 (N_8283,N_1811,N_3233);
and U8284 (N_8284,N_2421,N_1791);
nor U8285 (N_8285,N_994,N_2329);
and U8286 (N_8286,N_465,N_2937);
and U8287 (N_8287,N_1012,N_3981);
or U8288 (N_8288,N_3058,N_3381);
nand U8289 (N_8289,N_1582,N_1269);
or U8290 (N_8290,N_3831,N_103);
or U8291 (N_8291,N_3333,N_213);
and U8292 (N_8292,N_3806,N_680);
nor U8293 (N_8293,N_1588,N_4044);
or U8294 (N_8294,N_3010,N_4760);
nand U8295 (N_8295,N_3009,N_2296);
nand U8296 (N_8296,N_101,N_1587);
nor U8297 (N_8297,N_3972,N_2149);
or U8298 (N_8298,N_3674,N_4081);
nand U8299 (N_8299,N_3976,N_1754);
or U8300 (N_8300,N_1595,N_1405);
nand U8301 (N_8301,N_3098,N_3811);
nand U8302 (N_8302,N_4963,N_281);
and U8303 (N_8303,N_3094,N_647);
nand U8304 (N_8304,N_191,N_3255);
nor U8305 (N_8305,N_4381,N_363);
or U8306 (N_8306,N_1555,N_4441);
and U8307 (N_8307,N_259,N_203);
nor U8308 (N_8308,N_2588,N_1802);
or U8309 (N_8309,N_4522,N_3539);
and U8310 (N_8310,N_3436,N_2623);
nand U8311 (N_8311,N_1223,N_130);
or U8312 (N_8312,N_2504,N_1341);
nor U8313 (N_8313,N_947,N_4628);
nor U8314 (N_8314,N_1460,N_3919);
and U8315 (N_8315,N_760,N_2729);
nand U8316 (N_8316,N_1140,N_2935);
nand U8317 (N_8317,N_3279,N_1828);
nor U8318 (N_8318,N_180,N_3143);
and U8319 (N_8319,N_4182,N_3573);
and U8320 (N_8320,N_4258,N_153);
nand U8321 (N_8321,N_2754,N_3572);
nand U8322 (N_8322,N_3046,N_2226);
and U8323 (N_8323,N_2216,N_2623);
or U8324 (N_8324,N_1910,N_3294);
nor U8325 (N_8325,N_4279,N_1231);
nor U8326 (N_8326,N_3096,N_482);
nand U8327 (N_8327,N_2550,N_2618);
or U8328 (N_8328,N_1666,N_1056);
and U8329 (N_8329,N_4906,N_530);
nand U8330 (N_8330,N_4967,N_778);
or U8331 (N_8331,N_2910,N_3461);
nor U8332 (N_8332,N_819,N_3384);
or U8333 (N_8333,N_1896,N_3432);
and U8334 (N_8334,N_2302,N_1139);
and U8335 (N_8335,N_56,N_4000);
or U8336 (N_8336,N_3235,N_987);
nor U8337 (N_8337,N_2589,N_662);
and U8338 (N_8338,N_738,N_371);
nor U8339 (N_8339,N_4687,N_1334);
nor U8340 (N_8340,N_2980,N_276);
nor U8341 (N_8341,N_2332,N_727);
xnor U8342 (N_8342,N_1241,N_1078);
and U8343 (N_8343,N_3266,N_2509);
and U8344 (N_8344,N_1357,N_3903);
nor U8345 (N_8345,N_1727,N_3211);
nand U8346 (N_8346,N_3772,N_3332);
nand U8347 (N_8347,N_2194,N_4726);
nand U8348 (N_8348,N_2800,N_1719);
or U8349 (N_8349,N_952,N_1464);
nand U8350 (N_8350,N_2306,N_2021);
nand U8351 (N_8351,N_4475,N_1307);
and U8352 (N_8352,N_3289,N_1345);
nand U8353 (N_8353,N_120,N_3874);
nor U8354 (N_8354,N_2023,N_4881);
nand U8355 (N_8355,N_4373,N_3417);
and U8356 (N_8356,N_1646,N_2078);
or U8357 (N_8357,N_2039,N_175);
or U8358 (N_8358,N_613,N_2759);
and U8359 (N_8359,N_2225,N_299);
nor U8360 (N_8360,N_495,N_3477);
and U8361 (N_8361,N_2754,N_1360);
nor U8362 (N_8362,N_2461,N_3390);
or U8363 (N_8363,N_2836,N_830);
nor U8364 (N_8364,N_420,N_845);
or U8365 (N_8365,N_1073,N_835);
nor U8366 (N_8366,N_2785,N_2830);
nand U8367 (N_8367,N_429,N_2188);
nor U8368 (N_8368,N_1238,N_3399);
nor U8369 (N_8369,N_2783,N_2163);
nand U8370 (N_8370,N_1445,N_2112);
or U8371 (N_8371,N_1156,N_1188);
nor U8372 (N_8372,N_1431,N_99);
and U8373 (N_8373,N_1326,N_3630);
nand U8374 (N_8374,N_2131,N_119);
nor U8375 (N_8375,N_3060,N_4832);
and U8376 (N_8376,N_3030,N_505);
or U8377 (N_8377,N_2226,N_3419);
and U8378 (N_8378,N_4105,N_3452);
nand U8379 (N_8379,N_547,N_2689);
or U8380 (N_8380,N_2980,N_2413);
nor U8381 (N_8381,N_229,N_3480);
nand U8382 (N_8382,N_4070,N_3564);
nor U8383 (N_8383,N_761,N_3379);
or U8384 (N_8384,N_890,N_1366);
and U8385 (N_8385,N_2274,N_3935);
or U8386 (N_8386,N_4315,N_1768);
nand U8387 (N_8387,N_1399,N_2519);
nand U8388 (N_8388,N_3696,N_2113);
nand U8389 (N_8389,N_4962,N_537);
and U8390 (N_8390,N_1472,N_2046);
or U8391 (N_8391,N_1137,N_2233);
and U8392 (N_8392,N_806,N_3681);
and U8393 (N_8393,N_2293,N_4355);
nand U8394 (N_8394,N_4692,N_92);
or U8395 (N_8395,N_2359,N_3873);
nand U8396 (N_8396,N_1589,N_3688);
nand U8397 (N_8397,N_64,N_2920);
and U8398 (N_8398,N_2466,N_3583);
nor U8399 (N_8399,N_3748,N_2468);
and U8400 (N_8400,N_3845,N_781);
nor U8401 (N_8401,N_822,N_4853);
nand U8402 (N_8402,N_1295,N_2027);
or U8403 (N_8403,N_3280,N_1003);
and U8404 (N_8404,N_1471,N_2212);
and U8405 (N_8405,N_2564,N_254);
nand U8406 (N_8406,N_4631,N_2583);
nor U8407 (N_8407,N_3903,N_1708);
nor U8408 (N_8408,N_4002,N_2346);
nand U8409 (N_8409,N_2329,N_71);
and U8410 (N_8410,N_4390,N_2095);
nand U8411 (N_8411,N_824,N_1306);
or U8412 (N_8412,N_1804,N_3461);
nand U8413 (N_8413,N_3180,N_1203);
and U8414 (N_8414,N_1706,N_3904);
nand U8415 (N_8415,N_2695,N_4271);
nor U8416 (N_8416,N_4235,N_4930);
nand U8417 (N_8417,N_593,N_1552);
nor U8418 (N_8418,N_3452,N_4342);
and U8419 (N_8419,N_1863,N_679);
nand U8420 (N_8420,N_415,N_3667);
nand U8421 (N_8421,N_1916,N_3574);
or U8422 (N_8422,N_3755,N_3185);
nand U8423 (N_8423,N_3102,N_2578);
nand U8424 (N_8424,N_463,N_4371);
nand U8425 (N_8425,N_1067,N_392);
nand U8426 (N_8426,N_1850,N_1472);
nand U8427 (N_8427,N_1828,N_3746);
nor U8428 (N_8428,N_222,N_733);
and U8429 (N_8429,N_2671,N_471);
and U8430 (N_8430,N_3853,N_626);
nor U8431 (N_8431,N_2573,N_3472);
nand U8432 (N_8432,N_3701,N_3432);
nand U8433 (N_8433,N_3530,N_2754);
nor U8434 (N_8434,N_377,N_4885);
and U8435 (N_8435,N_3091,N_3124);
nand U8436 (N_8436,N_1391,N_67);
or U8437 (N_8437,N_4414,N_3179);
and U8438 (N_8438,N_4906,N_2705);
nand U8439 (N_8439,N_173,N_3801);
nand U8440 (N_8440,N_2767,N_4062);
nand U8441 (N_8441,N_980,N_1862);
and U8442 (N_8442,N_4111,N_4742);
nand U8443 (N_8443,N_4386,N_3537);
nand U8444 (N_8444,N_2468,N_3351);
nand U8445 (N_8445,N_2419,N_4989);
nand U8446 (N_8446,N_1934,N_3515);
or U8447 (N_8447,N_2083,N_2560);
nand U8448 (N_8448,N_2240,N_828);
and U8449 (N_8449,N_446,N_4664);
and U8450 (N_8450,N_2632,N_3435);
and U8451 (N_8451,N_3698,N_3785);
or U8452 (N_8452,N_1965,N_3553);
and U8453 (N_8453,N_4773,N_1229);
and U8454 (N_8454,N_712,N_3634);
and U8455 (N_8455,N_4862,N_3775);
nand U8456 (N_8456,N_2979,N_3031);
nor U8457 (N_8457,N_3087,N_4115);
or U8458 (N_8458,N_3146,N_3929);
or U8459 (N_8459,N_3274,N_3228);
and U8460 (N_8460,N_1276,N_3829);
nand U8461 (N_8461,N_4629,N_115);
and U8462 (N_8462,N_2243,N_2148);
and U8463 (N_8463,N_3074,N_1527);
nand U8464 (N_8464,N_157,N_4899);
and U8465 (N_8465,N_548,N_2269);
and U8466 (N_8466,N_1711,N_4375);
or U8467 (N_8467,N_552,N_3754);
and U8468 (N_8468,N_847,N_611);
nor U8469 (N_8469,N_2376,N_3169);
or U8470 (N_8470,N_24,N_1022);
and U8471 (N_8471,N_3640,N_842);
and U8472 (N_8472,N_3972,N_4162);
or U8473 (N_8473,N_159,N_3636);
nor U8474 (N_8474,N_4722,N_282);
nor U8475 (N_8475,N_1725,N_4931);
or U8476 (N_8476,N_2308,N_2856);
nor U8477 (N_8477,N_4792,N_1397);
xor U8478 (N_8478,N_2577,N_3811);
nand U8479 (N_8479,N_1604,N_1891);
or U8480 (N_8480,N_1738,N_1154);
nor U8481 (N_8481,N_2178,N_3670);
or U8482 (N_8482,N_2112,N_1242);
nand U8483 (N_8483,N_4654,N_368);
or U8484 (N_8484,N_359,N_2650);
nor U8485 (N_8485,N_3247,N_2925);
nor U8486 (N_8486,N_685,N_3154);
nor U8487 (N_8487,N_128,N_4636);
and U8488 (N_8488,N_428,N_50);
or U8489 (N_8489,N_4295,N_2727);
or U8490 (N_8490,N_1251,N_515);
nor U8491 (N_8491,N_551,N_2830);
nor U8492 (N_8492,N_2508,N_607);
nand U8493 (N_8493,N_33,N_2979);
and U8494 (N_8494,N_2962,N_3182);
nor U8495 (N_8495,N_4242,N_4089);
or U8496 (N_8496,N_3002,N_1048);
or U8497 (N_8497,N_4686,N_294);
or U8498 (N_8498,N_1671,N_938);
nand U8499 (N_8499,N_1740,N_4353);
nor U8500 (N_8500,N_2930,N_1997);
nor U8501 (N_8501,N_3913,N_3728);
nor U8502 (N_8502,N_1062,N_772);
nand U8503 (N_8503,N_781,N_689);
nor U8504 (N_8504,N_722,N_2165);
nand U8505 (N_8505,N_4514,N_3108);
and U8506 (N_8506,N_1733,N_2215);
xor U8507 (N_8507,N_2385,N_3626);
and U8508 (N_8508,N_4703,N_2945);
nor U8509 (N_8509,N_1053,N_1294);
nand U8510 (N_8510,N_577,N_2103);
nand U8511 (N_8511,N_14,N_3782);
or U8512 (N_8512,N_2756,N_1482);
or U8513 (N_8513,N_1183,N_1386);
nor U8514 (N_8514,N_551,N_53);
nor U8515 (N_8515,N_1544,N_3775);
or U8516 (N_8516,N_4934,N_3899);
nand U8517 (N_8517,N_526,N_6);
and U8518 (N_8518,N_3117,N_1066);
and U8519 (N_8519,N_4943,N_4584);
nor U8520 (N_8520,N_3316,N_3553);
nor U8521 (N_8521,N_3265,N_3232);
or U8522 (N_8522,N_1416,N_95);
nand U8523 (N_8523,N_4065,N_3704);
or U8524 (N_8524,N_2358,N_2398);
or U8525 (N_8525,N_3808,N_2866);
and U8526 (N_8526,N_3763,N_3099);
and U8527 (N_8527,N_1562,N_1840);
nand U8528 (N_8528,N_4210,N_2276);
or U8529 (N_8529,N_1706,N_1015);
xnor U8530 (N_8530,N_2703,N_925);
nor U8531 (N_8531,N_2645,N_843);
or U8532 (N_8532,N_3258,N_1955);
nand U8533 (N_8533,N_4089,N_2147);
nand U8534 (N_8534,N_4566,N_4427);
or U8535 (N_8535,N_1018,N_1537);
or U8536 (N_8536,N_3097,N_2170);
and U8537 (N_8537,N_4210,N_3630);
nor U8538 (N_8538,N_3752,N_24);
and U8539 (N_8539,N_327,N_3117);
nand U8540 (N_8540,N_3543,N_2791);
and U8541 (N_8541,N_4430,N_1927);
or U8542 (N_8542,N_4906,N_3636);
nor U8543 (N_8543,N_4325,N_2716);
and U8544 (N_8544,N_4238,N_1807);
and U8545 (N_8545,N_2054,N_1044);
nand U8546 (N_8546,N_2372,N_4874);
nand U8547 (N_8547,N_2178,N_148);
and U8548 (N_8548,N_4918,N_2557);
and U8549 (N_8549,N_711,N_3116);
nand U8550 (N_8550,N_141,N_3326);
nand U8551 (N_8551,N_4332,N_3861);
nand U8552 (N_8552,N_2754,N_2066);
nand U8553 (N_8553,N_1587,N_4471);
nand U8554 (N_8554,N_2827,N_3593);
nand U8555 (N_8555,N_1834,N_3995);
or U8556 (N_8556,N_1826,N_1328);
or U8557 (N_8557,N_941,N_1193);
or U8558 (N_8558,N_3284,N_2762);
and U8559 (N_8559,N_630,N_1287);
nand U8560 (N_8560,N_3506,N_4798);
and U8561 (N_8561,N_395,N_1849);
nand U8562 (N_8562,N_772,N_3639);
nor U8563 (N_8563,N_4489,N_3123);
nand U8564 (N_8564,N_2422,N_2515);
nor U8565 (N_8565,N_4199,N_4410);
nor U8566 (N_8566,N_4759,N_4537);
nand U8567 (N_8567,N_3881,N_4931);
nand U8568 (N_8568,N_1073,N_2681);
or U8569 (N_8569,N_4996,N_1037);
and U8570 (N_8570,N_2074,N_2713);
nand U8571 (N_8571,N_2567,N_1231);
nand U8572 (N_8572,N_3322,N_1330);
nor U8573 (N_8573,N_3043,N_2612);
nand U8574 (N_8574,N_797,N_4396);
or U8575 (N_8575,N_181,N_2172);
nor U8576 (N_8576,N_3679,N_4618);
nor U8577 (N_8577,N_2141,N_3762);
nand U8578 (N_8578,N_4652,N_2553);
and U8579 (N_8579,N_2615,N_4590);
or U8580 (N_8580,N_3906,N_2173);
xnor U8581 (N_8581,N_3227,N_1021);
nor U8582 (N_8582,N_937,N_1212);
or U8583 (N_8583,N_1724,N_2412);
and U8584 (N_8584,N_1611,N_417);
and U8585 (N_8585,N_2235,N_318);
nor U8586 (N_8586,N_1084,N_832);
nor U8587 (N_8587,N_959,N_2627);
and U8588 (N_8588,N_4209,N_1645);
or U8589 (N_8589,N_4808,N_220);
nor U8590 (N_8590,N_1237,N_4320);
or U8591 (N_8591,N_1552,N_2638);
nand U8592 (N_8592,N_331,N_2303);
nor U8593 (N_8593,N_3475,N_2962);
nor U8594 (N_8594,N_2179,N_135);
or U8595 (N_8595,N_631,N_1025);
and U8596 (N_8596,N_541,N_4029);
nor U8597 (N_8597,N_4675,N_843);
nand U8598 (N_8598,N_2664,N_4759);
nor U8599 (N_8599,N_4454,N_3734);
and U8600 (N_8600,N_4731,N_1443);
or U8601 (N_8601,N_3946,N_3778);
nor U8602 (N_8602,N_3072,N_2906);
and U8603 (N_8603,N_971,N_4608);
and U8604 (N_8604,N_4901,N_3051);
or U8605 (N_8605,N_4707,N_2453);
or U8606 (N_8606,N_57,N_3175);
and U8607 (N_8607,N_1459,N_974);
nor U8608 (N_8608,N_3467,N_1835);
nand U8609 (N_8609,N_222,N_3774);
and U8610 (N_8610,N_1646,N_1466);
nand U8611 (N_8611,N_4807,N_1334);
nor U8612 (N_8612,N_3276,N_3759);
or U8613 (N_8613,N_1932,N_975);
nand U8614 (N_8614,N_2130,N_4552);
nand U8615 (N_8615,N_2065,N_531);
nand U8616 (N_8616,N_4622,N_2079);
nand U8617 (N_8617,N_3927,N_4398);
or U8618 (N_8618,N_4948,N_3930);
and U8619 (N_8619,N_2950,N_712);
nor U8620 (N_8620,N_1530,N_3637);
or U8621 (N_8621,N_580,N_2946);
xor U8622 (N_8622,N_3748,N_4220);
or U8623 (N_8623,N_3203,N_2515);
or U8624 (N_8624,N_3710,N_669);
nand U8625 (N_8625,N_3968,N_55);
and U8626 (N_8626,N_4125,N_4563);
or U8627 (N_8627,N_2889,N_2539);
and U8628 (N_8628,N_2718,N_4956);
nor U8629 (N_8629,N_898,N_2969);
nand U8630 (N_8630,N_269,N_568);
and U8631 (N_8631,N_1781,N_3828);
or U8632 (N_8632,N_3481,N_3940);
and U8633 (N_8633,N_1794,N_1042);
and U8634 (N_8634,N_4887,N_1609);
or U8635 (N_8635,N_4294,N_529);
nand U8636 (N_8636,N_140,N_307);
nor U8637 (N_8637,N_2061,N_2371);
nor U8638 (N_8638,N_4918,N_475);
nand U8639 (N_8639,N_4883,N_4229);
nand U8640 (N_8640,N_1226,N_14);
or U8641 (N_8641,N_4980,N_1818);
nand U8642 (N_8642,N_3397,N_2960);
and U8643 (N_8643,N_2352,N_3591);
nand U8644 (N_8644,N_1320,N_88);
or U8645 (N_8645,N_1888,N_1298);
or U8646 (N_8646,N_705,N_2494);
or U8647 (N_8647,N_3230,N_454);
and U8648 (N_8648,N_3226,N_3366);
nor U8649 (N_8649,N_1172,N_397);
and U8650 (N_8650,N_1418,N_3300);
or U8651 (N_8651,N_532,N_1124);
or U8652 (N_8652,N_3260,N_4950);
nor U8653 (N_8653,N_3710,N_1765);
nor U8654 (N_8654,N_1053,N_4473);
or U8655 (N_8655,N_3740,N_3787);
and U8656 (N_8656,N_1332,N_2672);
or U8657 (N_8657,N_4233,N_2249);
nor U8658 (N_8658,N_4549,N_1293);
and U8659 (N_8659,N_3727,N_483);
nor U8660 (N_8660,N_2131,N_3164);
nor U8661 (N_8661,N_726,N_3106);
and U8662 (N_8662,N_222,N_3474);
or U8663 (N_8663,N_2233,N_1435);
or U8664 (N_8664,N_1161,N_1326);
or U8665 (N_8665,N_2488,N_1700);
nand U8666 (N_8666,N_3470,N_2925);
or U8667 (N_8667,N_4112,N_3409);
nor U8668 (N_8668,N_3053,N_881);
nand U8669 (N_8669,N_2642,N_114);
and U8670 (N_8670,N_4906,N_1301);
or U8671 (N_8671,N_3641,N_3599);
or U8672 (N_8672,N_2468,N_3429);
or U8673 (N_8673,N_679,N_63);
or U8674 (N_8674,N_305,N_228);
or U8675 (N_8675,N_3753,N_4625);
nor U8676 (N_8676,N_3613,N_864);
and U8677 (N_8677,N_4776,N_1297);
nor U8678 (N_8678,N_2209,N_2551);
nor U8679 (N_8679,N_1490,N_2364);
and U8680 (N_8680,N_4812,N_3331);
nor U8681 (N_8681,N_567,N_1602);
nor U8682 (N_8682,N_4869,N_1537);
or U8683 (N_8683,N_1779,N_4881);
or U8684 (N_8684,N_2409,N_4443);
nand U8685 (N_8685,N_1821,N_1983);
and U8686 (N_8686,N_2190,N_1020);
and U8687 (N_8687,N_1055,N_3398);
nand U8688 (N_8688,N_1401,N_3128);
nand U8689 (N_8689,N_4338,N_3903);
and U8690 (N_8690,N_3718,N_2569);
and U8691 (N_8691,N_1394,N_3692);
or U8692 (N_8692,N_4089,N_713);
nor U8693 (N_8693,N_211,N_4631);
or U8694 (N_8694,N_1036,N_2713);
or U8695 (N_8695,N_1517,N_1024);
or U8696 (N_8696,N_2532,N_4672);
nor U8697 (N_8697,N_23,N_996);
nand U8698 (N_8698,N_1368,N_4246);
nand U8699 (N_8699,N_4784,N_2329);
or U8700 (N_8700,N_656,N_2780);
and U8701 (N_8701,N_272,N_1389);
and U8702 (N_8702,N_4300,N_3470);
nor U8703 (N_8703,N_2625,N_4878);
and U8704 (N_8704,N_2914,N_658);
nand U8705 (N_8705,N_1649,N_890);
and U8706 (N_8706,N_979,N_2959);
and U8707 (N_8707,N_4275,N_4572);
and U8708 (N_8708,N_1826,N_3529);
nand U8709 (N_8709,N_3582,N_283);
nor U8710 (N_8710,N_3407,N_2790);
nand U8711 (N_8711,N_2814,N_2671);
nand U8712 (N_8712,N_221,N_618);
and U8713 (N_8713,N_4412,N_2762);
nand U8714 (N_8714,N_3006,N_3801);
xor U8715 (N_8715,N_4739,N_495);
nand U8716 (N_8716,N_1215,N_1814);
or U8717 (N_8717,N_587,N_2122);
nor U8718 (N_8718,N_4662,N_2952);
nand U8719 (N_8719,N_2118,N_2929);
or U8720 (N_8720,N_2692,N_1096);
nor U8721 (N_8721,N_2057,N_1396);
nand U8722 (N_8722,N_3357,N_313);
nand U8723 (N_8723,N_1361,N_3762);
nor U8724 (N_8724,N_2254,N_4934);
nor U8725 (N_8725,N_550,N_1141);
nand U8726 (N_8726,N_203,N_3027);
and U8727 (N_8727,N_3505,N_1480);
and U8728 (N_8728,N_4594,N_1550);
or U8729 (N_8729,N_18,N_3939);
or U8730 (N_8730,N_216,N_2030);
or U8731 (N_8731,N_807,N_2804);
nor U8732 (N_8732,N_4755,N_4836);
and U8733 (N_8733,N_2199,N_4807);
and U8734 (N_8734,N_2877,N_1547);
and U8735 (N_8735,N_334,N_4650);
and U8736 (N_8736,N_238,N_3047);
and U8737 (N_8737,N_4512,N_3781);
nand U8738 (N_8738,N_2660,N_1679);
or U8739 (N_8739,N_3395,N_246);
nand U8740 (N_8740,N_3460,N_3017);
and U8741 (N_8741,N_2625,N_2353);
or U8742 (N_8742,N_4582,N_2629);
nand U8743 (N_8743,N_950,N_3090);
and U8744 (N_8744,N_847,N_1037);
nor U8745 (N_8745,N_2281,N_2370);
and U8746 (N_8746,N_1913,N_3097);
and U8747 (N_8747,N_3268,N_3911);
or U8748 (N_8748,N_4524,N_3770);
nand U8749 (N_8749,N_2518,N_4920);
nand U8750 (N_8750,N_2347,N_1809);
and U8751 (N_8751,N_3321,N_2278);
or U8752 (N_8752,N_708,N_1286);
and U8753 (N_8753,N_1705,N_1889);
and U8754 (N_8754,N_3048,N_1208);
and U8755 (N_8755,N_3066,N_1410);
nand U8756 (N_8756,N_3505,N_3480);
and U8757 (N_8757,N_85,N_4202);
nand U8758 (N_8758,N_3490,N_831);
nand U8759 (N_8759,N_2561,N_4904);
nor U8760 (N_8760,N_770,N_2212);
or U8761 (N_8761,N_3925,N_3973);
nand U8762 (N_8762,N_409,N_3041);
and U8763 (N_8763,N_3133,N_4165);
or U8764 (N_8764,N_3970,N_2278);
or U8765 (N_8765,N_3522,N_3123);
or U8766 (N_8766,N_3740,N_2690);
nor U8767 (N_8767,N_3188,N_3014);
nor U8768 (N_8768,N_905,N_2923);
nand U8769 (N_8769,N_2534,N_199);
and U8770 (N_8770,N_4702,N_2897);
or U8771 (N_8771,N_123,N_4331);
and U8772 (N_8772,N_4865,N_2408);
nor U8773 (N_8773,N_3233,N_55);
nand U8774 (N_8774,N_3898,N_993);
nor U8775 (N_8775,N_3472,N_2371);
nand U8776 (N_8776,N_2875,N_2865);
nor U8777 (N_8777,N_3885,N_2507);
and U8778 (N_8778,N_3308,N_3296);
nand U8779 (N_8779,N_674,N_4377);
and U8780 (N_8780,N_322,N_3544);
nand U8781 (N_8781,N_1616,N_120);
and U8782 (N_8782,N_2255,N_1470);
or U8783 (N_8783,N_1606,N_440);
nand U8784 (N_8784,N_230,N_1669);
and U8785 (N_8785,N_3747,N_1035);
or U8786 (N_8786,N_142,N_806);
or U8787 (N_8787,N_4967,N_147);
nor U8788 (N_8788,N_4355,N_3036);
and U8789 (N_8789,N_1733,N_751);
and U8790 (N_8790,N_4371,N_1079);
nor U8791 (N_8791,N_2549,N_1562);
and U8792 (N_8792,N_310,N_961);
nor U8793 (N_8793,N_626,N_4220);
and U8794 (N_8794,N_1769,N_2966);
nor U8795 (N_8795,N_2531,N_648);
or U8796 (N_8796,N_3070,N_180);
nand U8797 (N_8797,N_2153,N_2154);
or U8798 (N_8798,N_3954,N_2447);
or U8799 (N_8799,N_422,N_3262);
nor U8800 (N_8800,N_1774,N_1492);
nand U8801 (N_8801,N_3979,N_3456);
nand U8802 (N_8802,N_2130,N_3520);
nand U8803 (N_8803,N_832,N_4869);
nor U8804 (N_8804,N_1526,N_3654);
nand U8805 (N_8805,N_3631,N_4945);
nor U8806 (N_8806,N_2039,N_4999);
nand U8807 (N_8807,N_276,N_4325);
or U8808 (N_8808,N_3540,N_1421);
or U8809 (N_8809,N_1424,N_3636);
nand U8810 (N_8810,N_4479,N_424);
or U8811 (N_8811,N_3105,N_2526);
nand U8812 (N_8812,N_2484,N_904);
or U8813 (N_8813,N_958,N_3664);
and U8814 (N_8814,N_1511,N_4004);
nor U8815 (N_8815,N_4910,N_3475);
nor U8816 (N_8816,N_4483,N_3280);
nor U8817 (N_8817,N_2560,N_973);
nor U8818 (N_8818,N_172,N_883);
nor U8819 (N_8819,N_4853,N_188);
or U8820 (N_8820,N_1412,N_1636);
nor U8821 (N_8821,N_748,N_1622);
nor U8822 (N_8822,N_1203,N_509);
or U8823 (N_8823,N_3165,N_2896);
nor U8824 (N_8824,N_2717,N_1582);
nor U8825 (N_8825,N_1708,N_532);
and U8826 (N_8826,N_1109,N_590);
or U8827 (N_8827,N_2973,N_2139);
nand U8828 (N_8828,N_4584,N_3402);
nor U8829 (N_8829,N_3818,N_575);
nor U8830 (N_8830,N_4724,N_4427);
and U8831 (N_8831,N_3387,N_1748);
and U8832 (N_8832,N_947,N_3425);
and U8833 (N_8833,N_856,N_1045);
nand U8834 (N_8834,N_946,N_97);
nor U8835 (N_8835,N_4643,N_4863);
or U8836 (N_8836,N_3541,N_678);
and U8837 (N_8837,N_3997,N_1453);
or U8838 (N_8838,N_2623,N_1338);
and U8839 (N_8839,N_1902,N_4418);
and U8840 (N_8840,N_4923,N_2166);
nor U8841 (N_8841,N_1762,N_336);
nor U8842 (N_8842,N_4774,N_1557);
and U8843 (N_8843,N_375,N_2223);
nor U8844 (N_8844,N_1528,N_192);
or U8845 (N_8845,N_4213,N_1818);
nor U8846 (N_8846,N_1571,N_1152);
nor U8847 (N_8847,N_4162,N_1467);
nand U8848 (N_8848,N_4064,N_1984);
or U8849 (N_8849,N_1624,N_841);
nand U8850 (N_8850,N_4280,N_4497);
nand U8851 (N_8851,N_1720,N_3371);
nand U8852 (N_8852,N_1893,N_2159);
nand U8853 (N_8853,N_4257,N_2596);
nand U8854 (N_8854,N_616,N_3349);
nand U8855 (N_8855,N_293,N_788);
nor U8856 (N_8856,N_1662,N_1347);
nand U8857 (N_8857,N_4604,N_4538);
nor U8858 (N_8858,N_3833,N_4782);
xnor U8859 (N_8859,N_3021,N_1097);
and U8860 (N_8860,N_3404,N_4288);
and U8861 (N_8861,N_1475,N_1577);
nand U8862 (N_8862,N_4769,N_4944);
nor U8863 (N_8863,N_2326,N_1652);
nor U8864 (N_8864,N_195,N_499);
nor U8865 (N_8865,N_3432,N_1052);
and U8866 (N_8866,N_2914,N_2091);
nand U8867 (N_8867,N_1807,N_2651);
nand U8868 (N_8868,N_2895,N_994);
nor U8869 (N_8869,N_4073,N_2388);
and U8870 (N_8870,N_4347,N_2007);
nand U8871 (N_8871,N_519,N_1657);
and U8872 (N_8872,N_675,N_2045);
nand U8873 (N_8873,N_1424,N_655);
nor U8874 (N_8874,N_1414,N_4333);
and U8875 (N_8875,N_4688,N_3336);
xnor U8876 (N_8876,N_4565,N_4023);
or U8877 (N_8877,N_1274,N_671);
xor U8878 (N_8878,N_3156,N_1428);
nand U8879 (N_8879,N_4443,N_2205);
or U8880 (N_8880,N_928,N_479);
nor U8881 (N_8881,N_4636,N_4573);
or U8882 (N_8882,N_1688,N_164);
nand U8883 (N_8883,N_852,N_1509);
nor U8884 (N_8884,N_1623,N_4423);
nand U8885 (N_8885,N_3236,N_1066);
and U8886 (N_8886,N_106,N_119);
nand U8887 (N_8887,N_3092,N_211);
nand U8888 (N_8888,N_19,N_1826);
nand U8889 (N_8889,N_4033,N_922);
or U8890 (N_8890,N_4127,N_4464);
nand U8891 (N_8891,N_3879,N_3281);
nor U8892 (N_8892,N_4232,N_847);
or U8893 (N_8893,N_803,N_4676);
or U8894 (N_8894,N_929,N_2715);
nand U8895 (N_8895,N_2860,N_689);
nand U8896 (N_8896,N_3500,N_2175);
nor U8897 (N_8897,N_3174,N_2934);
or U8898 (N_8898,N_630,N_4984);
xnor U8899 (N_8899,N_4748,N_3775);
nand U8900 (N_8900,N_1678,N_714);
or U8901 (N_8901,N_1730,N_3884);
and U8902 (N_8902,N_2975,N_2304);
nand U8903 (N_8903,N_2386,N_248);
nor U8904 (N_8904,N_291,N_798);
nor U8905 (N_8905,N_3395,N_1016);
and U8906 (N_8906,N_881,N_1835);
and U8907 (N_8907,N_4183,N_248);
nor U8908 (N_8908,N_4126,N_4395);
and U8909 (N_8909,N_2057,N_1636);
and U8910 (N_8910,N_341,N_3503);
nor U8911 (N_8911,N_1762,N_4150);
nand U8912 (N_8912,N_2011,N_3048);
and U8913 (N_8913,N_3658,N_2962);
or U8914 (N_8914,N_2341,N_13);
nor U8915 (N_8915,N_1122,N_641);
and U8916 (N_8916,N_94,N_495);
and U8917 (N_8917,N_4608,N_152);
or U8918 (N_8918,N_1804,N_3392);
nand U8919 (N_8919,N_2698,N_3162);
nor U8920 (N_8920,N_3823,N_916);
nand U8921 (N_8921,N_2369,N_2108);
nand U8922 (N_8922,N_2203,N_3550);
or U8923 (N_8923,N_1895,N_2197);
or U8924 (N_8924,N_3088,N_3895);
and U8925 (N_8925,N_3089,N_3189);
nand U8926 (N_8926,N_2121,N_1020);
nand U8927 (N_8927,N_1370,N_1089);
xor U8928 (N_8928,N_3271,N_1310);
nand U8929 (N_8929,N_1983,N_3696);
nor U8930 (N_8930,N_3256,N_2557);
xnor U8931 (N_8931,N_1832,N_3502);
nand U8932 (N_8932,N_3884,N_3008);
nor U8933 (N_8933,N_4713,N_4349);
nor U8934 (N_8934,N_3848,N_3916);
nand U8935 (N_8935,N_1833,N_2836);
nor U8936 (N_8936,N_2742,N_1652);
or U8937 (N_8937,N_4325,N_2186);
or U8938 (N_8938,N_915,N_126);
or U8939 (N_8939,N_4824,N_2584);
and U8940 (N_8940,N_3588,N_3399);
or U8941 (N_8941,N_1491,N_2198);
nand U8942 (N_8942,N_4621,N_4838);
nor U8943 (N_8943,N_3669,N_3776);
and U8944 (N_8944,N_4645,N_69);
or U8945 (N_8945,N_1444,N_231);
nand U8946 (N_8946,N_1738,N_3533);
nor U8947 (N_8947,N_1980,N_303);
and U8948 (N_8948,N_1454,N_3785);
nor U8949 (N_8949,N_3266,N_3285);
and U8950 (N_8950,N_4283,N_3701);
nor U8951 (N_8951,N_181,N_3233);
or U8952 (N_8952,N_4214,N_4936);
and U8953 (N_8953,N_2664,N_3303);
nor U8954 (N_8954,N_1503,N_1892);
nand U8955 (N_8955,N_3130,N_2129);
or U8956 (N_8956,N_4392,N_251);
nand U8957 (N_8957,N_2454,N_1006);
or U8958 (N_8958,N_4161,N_554);
or U8959 (N_8959,N_4490,N_2868);
or U8960 (N_8960,N_2651,N_1884);
and U8961 (N_8961,N_2897,N_2575);
nor U8962 (N_8962,N_2866,N_917);
or U8963 (N_8963,N_3525,N_4804);
or U8964 (N_8964,N_3563,N_4452);
or U8965 (N_8965,N_4838,N_69);
and U8966 (N_8966,N_1866,N_1097);
and U8967 (N_8967,N_3773,N_3811);
nor U8968 (N_8968,N_500,N_1014);
and U8969 (N_8969,N_1092,N_204);
or U8970 (N_8970,N_2742,N_2179);
and U8971 (N_8971,N_3742,N_4526);
nor U8972 (N_8972,N_1800,N_398);
or U8973 (N_8973,N_3299,N_3462);
or U8974 (N_8974,N_2601,N_1204);
nor U8975 (N_8975,N_3531,N_1511);
nand U8976 (N_8976,N_1743,N_1962);
nand U8977 (N_8977,N_437,N_1921);
and U8978 (N_8978,N_3745,N_4353);
and U8979 (N_8979,N_1354,N_4513);
and U8980 (N_8980,N_4168,N_2034);
nor U8981 (N_8981,N_2799,N_3964);
and U8982 (N_8982,N_3920,N_3034);
or U8983 (N_8983,N_1138,N_2957);
nor U8984 (N_8984,N_2320,N_641);
and U8985 (N_8985,N_2120,N_2225);
and U8986 (N_8986,N_4361,N_285);
nor U8987 (N_8987,N_3271,N_300);
nor U8988 (N_8988,N_72,N_4879);
nand U8989 (N_8989,N_1357,N_1211);
and U8990 (N_8990,N_1792,N_2904);
nor U8991 (N_8991,N_1270,N_3930);
and U8992 (N_8992,N_3572,N_3354);
or U8993 (N_8993,N_49,N_3031);
nand U8994 (N_8994,N_3504,N_3338);
or U8995 (N_8995,N_2015,N_3487);
nor U8996 (N_8996,N_2213,N_3273);
and U8997 (N_8997,N_1915,N_3288);
nand U8998 (N_8998,N_1764,N_538);
nand U8999 (N_8999,N_4817,N_1193);
nand U9000 (N_9000,N_4026,N_563);
or U9001 (N_9001,N_107,N_4755);
nor U9002 (N_9002,N_155,N_4017);
and U9003 (N_9003,N_1724,N_893);
nor U9004 (N_9004,N_4058,N_1615);
and U9005 (N_9005,N_2382,N_1642);
nor U9006 (N_9006,N_644,N_2622);
or U9007 (N_9007,N_177,N_937);
and U9008 (N_9008,N_2593,N_195);
and U9009 (N_9009,N_1650,N_3534);
nor U9010 (N_9010,N_3144,N_4494);
nand U9011 (N_9011,N_505,N_3918);
or U9012 (N_9012,N_92,N_1124);
nand U9013 (N_9013,N_4249,N_4865);
or U9014 (N_9014,N_1766,N_2197);
nor U9015 (N_9015,N_4649,N_573);
and U9016 (N_9016,N_3944,N_1254);
nand U9017 (N_9017,N_1947,N_2970);
nand U9018 (N_9018,N_626,N_2002);
and U9019 (N_9019,N_4609,N_976);
nand U9020 (N_9020,N_658,N_3767);
and U9021 (N_9021,N_2386,N_4399);
nor U9022 (N_9022,N_4290,N_4281);
nor U9023 (N_9023,N_255,N_2610);
nor U9024 (N_9024,N_2158,N_4976);
and U9025 (N_9025,N_3628,N_3250);
or U9026 (N_9026,N_4714,N_1644);
and U9027 (N_9027,N_4394,N_4969);
and U9028 (N_9028,N_668,N_2856);
or U9029 (N_9029,N_1781,N_3712);
or U9030 (N_9030,N_479,N_867);
and U9031 (N_9031,N_4619,N_1371);
nor U9032 (N_9032,N_4525,N_2835);
and U9033 (N_9033,N_294,N_1738);
or U9034 (N_9034,N_1683,N_2740);
or U9035 (N_9035,N_147,N_2015);
nor U9036 (N_9036,N_3628,N_4172);
nand U9037 (N_9037,N_4327,N_617);
nand U9038 (N_9038,N_773,N_2802);
nor U9039 (N_9039,N_126,N_1683);
or U9040 (N_9040,N_2607,N_1844);
nand U9041 (N_9041,N_3509,N_4332);
or U9042 (N_9042,N_231,N_2521);
or U9043 (N_9043,N_1363,N_805);
and U9044 (N_9044,N_2254,N_1511);
and U9045 (N_9045,N_3198,N_4530);
nand U9046 (N_9046,N_2793,N_45);
or U9047 (N_9047,N_4552,N_1080);
and U9048 (N_9048,N_343,N_1423);
and U9049 (N_9049,N_1133,N_3413);
nor U9050 (N_9050,N_2596,N_4730);
or U9051 (N_9051,N_3552,N_1919);
and U9052 (N_9052,N_1297,N_2832);
nor U9053 (N_9053,N_2430,N_4214);
nand U9054 (N_9054,N_4678,N_3457);
nand U9055 (N_9055,N_3442,N_2943);
and U9056 (N_9056,N_730,N_148);
nor U9057 (N_9057,N_3518,N_3180);
or U9058 (N_9058,N_2834,N_1966);
and U9059 (N_9059,N_519,N_280);
nor U9060 (N_9060,N_187,N_3934);
and U9061 (N_9061,N_2760,N_4922);
or U9062 (N_9062,N_925,N_3279);
and U9063 (N_9063,N_794,N_1173);
nand U9064 (N_9064,N_2604,N_4440);
or U9065 (N_9065,N_4002,N_2184);
nor U9066 (N_9066,N_3102,N_2917);
nand U9067 (N_9067,N_4193,N_4790);
nor U9068 (N_9068,N_3010,N_4970);
nor U9069 (N_9069,N_68,N_2749);
nand U9070 (N_9070,N_3667,N_2133);
nand U9071 (N_9071,N_4231,N_1565);
and U9072 (N_9072,N_1058,N_2783);
and U9073 (N_9073,N_4296,N_4672);
nand U9074 (N_9074,N_1663,N_3925);
nand U9075 (N_9075,N_3236,N_3831);
nand U9076 (N_9076,N_2688,N_2265);
xor U9077 (N_9077,N_4717,N_125);
and U9078 (N_9078,N_3919,N_3267);
or U9079 (N_9079,N_3452,N_3480);
or U9080 (N_9080,N_3763,N_2978);
nor U9081 (N_9081,N_4110,N_2531);
nand U9082 (N_9082,N_4580,N_2884);
nand U9083 (N_9083,N_2978,N_4416);
and U9084 (N_9084,N_245,N_3938);
or U9085 (N_9085,N_799,N_4183);
nor U9086 (N_9086,N_1757,N_3148);
and U9087 (N_9087,N_3286,N_3604);
nand U9088 (N_9088,N_370,N_2825);
nand U9089 (N_9089,N_2584,N_1437);
nor U9090 (N_9090,N_3111,N_3478);
and U9091 (N_9091,N_4872,N_1359);
nor U9092 (N_9092,N_538,N_3413);
nand U9093 (N_9093,N_4515,N_4942);
and U9094 (N_9094,N_3259,N_4524);
nor U9095 (N_9095,N_4293,N_943);
nor U9096 (N_9096,N_4695,N_2786);
or U9097 (N_9097,N_327,N_3822);
nand U9098 (N_9098,N_1513,N_3982);
xnor U9099 (N_9099,N_1118,N_3210);
and U9100 (N_9100,N_3732,N_4283);
and U9101 (N_9101,N_2340,N_2791);
or U9102 (N_9102,N_372,N_2760);
nor U9103 (N_9103,N_3508,N_3013);
or U9104 (N_9104,N_2961,N_752);
nor U9105 (N_9105,N_994,N_2347);
and U9106 (N_9106,N_1434,N_1308);
nand U9107 (N_9107,N_3847,N_2923);
or U9108 (N_9108,N_545,N_803);
and U9109 (N_9109,N_1577,N_2434);
or U9110 (N_9110,N_2463,N_496);
nor U9111 (N_9111,N_1882,N_2351);
and U9112 (N_9112,N_3747,N_1980);
nand U9113 (N_9113,N_2306,N_3772);
and U9114 (N_9114,N_4993,N_2589);
nand U9115 (N_9115,N_4454,N_845);
or U9116 (N_9116,N_2740,N_4325);
nor U9117 (N_9117,N_241,N_1098);
or U9118 (N_9118,N_4090,N_253);
and U9119 (N_9119,N_3348,N_1241);
and U9120 (N_9120,N_1003,N_4776);
and U9121 (N_9121,N_2159,N_776);
nor U9122 (N_9122,N_3492,N_3412);
nor U9123 (N_9123,N_4890,N_2081);
nor U9124 (N_9124,N_3171,N_3998);
or U9125 (N_9125,N_179,N_2380);
nor U9126 (N_9126,N_814,N_4599);
or U9127 (N_9127,N_788,N_1312);
or U9128 (N_9128,N_3950,N_1434);
or U9129 (N_9129,N_229,N_765);
nor U9130 (N_9130,N_4434,N_1153);
and U9131 (N_9131,N_4180,N_26);
and U9132 (N_9132,N_4552,N_3196);
xor U9133 (N_9133,N_1876,N_2019);
nand U9134 (N_9134,N_577,N_4228);
nor U9135 (N_9135,N_4241,N_2576);
and U9136 (N_9136,N_4182,N_4759);
nand U9137 (N_9137,N_534,N_2652);
nor U9138 (N_9138,N_4336,N_3616);
or U9139 (N_9139,N_1682,N_1951);
and U9140 (N_9140,N_253,N_4572);
and U9141 (N_9141,N_1394,N_3862);
nor U9142 (N_9142,N_416,N_107);
and U9143 (N_9143,N_1197,N_1652);
nand U9144 (N_9144,N_1633,N_1079);
or U9145 (N_9145,N_391,N_1874);
nor U9146 (N_9146,N_933,N_59);
or U9147 (N_9147,N_356,N_297);
nand U9148 (N_9148,N_3178,N_4914);
nand U9149 (N_9149,N_4134,N_2776);
and U9150 (N_9150,N_2153,N_4675);
and U9151 (N_9151,N_2674,N_4654);
or U9152 (N_9152,N_3064,N_1275);
or U9153 (N_9153,N_3098,N_2864);
and U9154 (N_9154,N_352,N_3693);
and U9155 (N_9155,N_1622,N_2508);
and U9156 (N_9156,N_1652,N_2827);
nand U9157 (N_9157,N_3624,N_4567);
nor U9158 (N_9158,N_1862,N_1368);
and U9159 (N_9159,N_3561,N_3788);
nand U9160 (N_9160,N_3058,N_2224);
or U9161 (N_9161,N_3239,N_4525);
or U9162 (N_9162,N_2514,N_820);
and U9163 (N_9163,N_1651,N_4584);
and U9164 (N_9164,N_1547,N_2014);
nor U9165 (N_9165,N_730,N_1197);
or U9166 (N_9166,N_289,N_3336);
or U9167 (N_9167,N_2122,N_2046);
and U9168 (N_9168,N_2842,N_2643);
or U9169 (N_9169,N_4387,N_3344);
and U9170 (N_9170,N_817,N_257);
and U9171 (N_9171,N_4013,N_859);
or U9172 (N_9172,N_2839,N_2445);
nand U9173 (N_9173,N_4672,N_667);
or U9174 (N_9174,N_1055,N_421);
and U9175 (N_9175,N_3195,N_2575);
and U9176 (N_9176,N_1962,N_1449);
and U9177 (N_9177,N_3745,N_4760);
or U9178 (N_9178,N_2118,N_3921);
or U9179 (N_9179,N_595,N_4230);
and U9180 (N_9180,N_1810,N_3394);
or U9181 (N_9181,N_4014,N_941);
nand U9182 (N_9182,N_2732,N_2902);
and U9183 (N_9183,N_569,N_1004);
nand U9184 (N_9184,N_4387,N_2669);
nand U9185 (N_9185,N_4956,N_993);
xnor U9186 (N_9186,N_2004,N_4743);
nand U9187 (N_9187,N_4918,N_1872);
nand U9188 (N_9188,N_2878,N_1034);
nor U9189 (N_9189,N_4083,N_604);
nand U9190 (N_9190,N_4896,N_4725);
nand U9191 (N_9191,N_2509,N_4311);
and U9192 (N_9192,N_4829,N_3480);
nand U9193 (N_9193,N_580,N_2274);
and U9194 (N_9194,N_796,N_362);
or U9195 (N_9195,N_254,N_1923);
nand U9196 (N_9196,N_2574,N_173);
and U9197 (N_9197,N_220,N_4516);
nor U9198 (N_9198,N_2388,N_1883);
nor U9199 (N_9199,N_3383,N_3540);
nand U9200 (N_9200,N_1386,N_60);
and U9201 (N_9201,N_2787,N_1546);
or U9202 (N_9202,N_4258,N_2448);
nor U9203 (N_9203,N_2109,N_3105);
or U9204 (N_9204,N_783,N_404);
and U9205 (N_9205,N_2096,N_2170);
nand U9206 (N_9206,N_4675,N_1605);
or U9207 (N_9207,N_1591,N_4030);
nor U9208 (N_9208,N_993,N_753);
or U9209 (N_9209,N_364,N_1275);
nor U9210 (N_9210,N_1409,N_3706);
or U9211 (N_9211,N_1395,N_2762);
nor U9212 (N_9212,N_3873,N_4312);
or U9213 (N_9213,N_4643,N_1264);
and U9214 (N_9214,N_1173,N_1212);
or U9215 (N_9215,N_4755,N_4980);
and U9216 (N_9216,N_4624,N_2045);
nand U9217 (N_9217,N_2307,N_1821);
and U9218 (N_9218,N_3746,N_3780);
nand U9219 (N_9219,N_1047,N_401);
nor U9220 (N_9220,N_997,N_2741);
nor U9221 (N_9221,N_3304,N_2845);
or U9222 (N_9222,N_698,N_1285);
nand U9223 (N_9223,N_3167,N_11);
or U9224 (N_9224,N_1277,N_475);
and U9225 (N_9225,N_2898,N_2464);
and U9226 (N_9226,N_4761,N_4547);
nand U9227 (N_9227,N_525,N_606);
nor U9228 (N_9228,N_1809,N_4477);
and U9229 (N_9229,N_584,N_4867);
or U9230 (N_9230,N_1727,N_815);
or U9231 (N_9231,N_3787,N_788);
and U9232 (N_9232,N_2801,N_732);
nand U9233 (N_9233,N_4006,N_1148);
and U9234 (N_9234,N_2575,N_1832);
or U9235 (N_9235,N_2610,N_3021);
or U9236 (N_9236,N_647,N_1536);
and U9237 (N_9237,N_4241,N_2142);
or U9238 (N_9238,N_3896,N_2825);
or U9239 (N_9239,N_4306,N_3426);
and U9240 (N_9240,N_2589,N_2679);
nand U9241 (N_9241,N_344,N_1500);
and U9242 (N_9242,N_1710,N_1053);
nor U9243 (N_9243,N_263,N_3971);
nor U9244 (N_9244,N_1808,N_2073);
and U9245 (N_9245,N_2378,N_3453);
nand U9246 (N_9246,N_3597,N_3547);
nor U9247 (N_9247,N_3469,N_1234);
nor U9248 (N_9248,N_148,N_796);
nor U9249 (N_9249,N_1642,N_954);
nor U9250 (N_9250,N_524,N_3940);
nand U9251 (N_9251,N_725,N_2160);
or U9252 (N_9252,N_22,N_299);
nor U9253 (N_9253,N_4635,N_1526);
nor U9254 (N_9254,N_4204,N_3532);
nand U9255 (N_9255,N_4095,N_4936);
xnor U9256 (N_9256,N_4489,N_1713);
nor U9257 (N_9257,N_2524,N_4984);
nor U9258 (N_9258,N_4517,N_1804);
nor U9259 (N_9259,N_4131,N_1978);
nand U9260 (N_9260,N_2424,N_4655);
and U9261 (N_9261,N_450,N_489);
or U9262 (N_9262,N_2296,N_2869);
nor U9263 (N_9263,N_95,N_2487);
nand U9264 (N_9264,N_402,N_1397);
or U9265 (N_9265,N_3677,N_709);
or U9266 (N_9266,N_4817,N_4790);
or U9267 (N_9267,N_94,N_4643);
or U9268 (N_9268,N_894,N_3634);
nor U9269 (N_9269,N_2335,N_2914);
or U9270 (N_9270,N_1770,N_458);
nand U9271 (N_9271,N_3767,N_3538);
nor U9272 (N_9272,N_2251,N_4522);
or U9273 (N_9273,N_2485,N_4667);
nand U9274 (N_9274,N_161,N_2490);
or U9275 (N_9275,N_3927,N_1345);
and U9276 (N_9276,N_1866,N_418);
or U9277 (N_9277,N_2499,N_1936);
or U9278 (N_9278,N_1116,N_1641);
nand U9279 (N_9279,N_1197,N_2348);
or U9280 (N_9280,N_4937,N_1048);
nor U9281 (N_9281,N_4651,N_2072);
or U9282 (N_9282,N_1047,N_3539);
nand U9283 (N_9283,N_3103,N_2157);
or U9284 (N_9284,N_3897,N_2980);
nand U9285 (N_9285,N_2438,N_3010);
or U9286 (N_9286,N_2061,N_4873);
or U9287 (N_9287,N_198,N_293);
nor U9288 (N_9288,N_4086,N_2153);
and U9289 (N_9289,N_1660,N_2663);
or U9290 (N_9290,N_3586,N_3687);
or U9291 (N_9291,N_2193,N_4092);
nor U9292 (N_9292,N_4225,N_338);
nor U9293 (N_9293,N_1058,N_855);
nand U9294 (N_9294,N_2301,N_4642);
nand U9295 (N_9295,N_2811,N_2088);
and U9296 (N_9296,N_1839,N_4033);
nand U9297 (N_9297,N_4368,N_1849);
and U9298 (N_9298,N_1529,N_1301);
and U9299 (N_9299,N_2028,N_2598);
nand U9300 (N_9300,N_3412,N_990);
or U9301 (N_9301,N_3770,N_4092);
or U9302 (N_9302,N_533,N_1512);
or U9303 (N_9303,N_2856,N_2766);
nor U9304 (N_9304,N_667,N_707);
or U9305 (N_9305,N_3169,N_1598);
and U9306 (N_9306,N_4131,N_2708);
nand U9307 (N_9307,N_4999,N_2435);
or U9308 (N_9308,N_2312,N_1896);
or U9309 (N_9309,N_129,N_676);
or U9310 (N_9310,N_1363,N_2692);
or U9311 (N_9311,N_3794,N_658);
and U9312 (N_9312,N_4474,N_3288);
nor U9313 (N_9313,N_1276,N_1872);
nor U9314 (N_9314,N_438,N_1025);
and U9315 (N_9315,N_2057,N_4706);
nand U9316 (N_9316,N_3152,N_3293);
or U9317 (N_9317,N_4519,N_1533);
nand U9318 (N_9318,N_1690,N_4924);
and U9319 (N_9319,N_4552,N_1509);
nand U9320 (N_9320,N_4917,N_2077);
nor U9321 (N_9321,N_2265,N_509);
or U9322 (N_9322,N_2795,N_3659);
nand U9323 (N_9323,N_978,N_3628);
nand U9324 (N_9324,N_2518,N_1354);
or U9325 (N_9325,N_2597,N_1951);
nor U9326 (N_9326,N_1054,N_1753);
nand U9327 (N_9327,N_2435,N_1181);
nand U9328 (N_9328,N_4925,N_158);
nand U9329 (N_9329,N_2653,N_3171);
and U9330 (N_9330,N_3591,N_3025);
nand U9331 (N_9331,N_1722,N_3905);
and U9332 (N_9332,N_2007,N_1458);
and U9333 (N_9333,N_988,N_2515);
or U9334 (N_9334,N_311,N_4716);
or U9335 (N_9335,N_4120,N_1775);
nor U9336 (N_9336,N_1455,N_1871);
nand U9337 (N_9337,N_2086,N_1746);
or U9338 (N_9338,N_1790,N_1396);
and U9339 (N_9339,N_4692,N_2178);
nor U9340 (N_9340,N_3758,N_2196);
nand U9341 (N_9341,N_1164,N_2754);
nand U9342 (N_9342,N_495,N_1645);
nor U9343 (N_9343,N_4439,N_1953);
nand U9344 (N_9344,N_117,N_3452);
nor U9345 (N_9345,N_4987,N_3834);
nand U9346 (N_9346,N_759,N_2867);
or U9347 (N_9347,N_49,N_2441);
nand U9348 (N_9348,N_2689,N_2045);
nand U9349 (N_9349,N_3088,N_2373);
nor U9350 (N_9350,N_2031,N_3905);
nor U9351 (N_9351,N_1376,N_4139);
or U9352 (N_9352,N_263,N_2415);
nand U9353 (N_9353,N_155,N_3626);
nor U9354 (N_9354,N_2096,N_4399);
nor U9355 (N_9355,N_2762,N_3917);
and U9356 (N_9356,N_2088,N_2115);
nor U9357 (N_9357,N_596,N_1137);
and U9358 (N_9358,N_3544,N_1782);
and U9359 (N_9359,N_483,N_3598);
or U9360 (N_9360,N_3008,N_4921);
or U9361 (N_9361,N_213,N_4783);
nor U9362 (N_9362,N_488,N_4955);
nand U9363 (N_9363,N_1621,N_1109);
or U9364 (N_9364,N_1479,N_2580);
nand U9365 (N_9365,N_2576,N_2485);
nand U9366 (N_9366,N_4081,N_4587);
nand U9367 (N_9367,N_796,N_2467);
or U9368 (N_9368,N_400,N_3505);
or U9369 (N_9369,N_1949,N_4517);
or U9370 (N_9370,N_288,N_1482);
or U9371 (N_9371,N_2460,N_45);
nand U9372 (N_9372,N_460,N_3240);
nand U9373 (N_9373,N_1356,N_2315);
or U9374 (N_9374,N_2050,N_3031);
or U9375 (N_9375,N_2322,N_4577);
or U9376 (N_9376,N_1519,N_1506);
and U9377 (N_9377,N_1560,N_4184);
nand U9378 (N_9378,N_4896,N_4471);
and U9379 (N_9379,N_541,N_4337);
nor U9380 (N_9380,N_26,N_3173);
nand U9381 (N_9381,N_1884,N_3013);
and U9382 (N_9382,N_4048,N_3519);
nand U9383 (N_9383,N_1556,N_1389);
or U9384 (N_9384,N_2884,N_1561);
or U9385 (N_9385,N_1246,N_2295);
nor U9386 (N_9386,N_527,N_3947);
and U9387 (N_9387,N_3472,N_862);
nor U9388 (N_9388,N_2572,N_2193);
or U9389 (N_9389,N_4325,N_2902);
and U9390 (N_9390,N_3360,N_3850);
or U9391 (N_9391,N_3544,N_1858);
nand U9392 (N_9392,N_207,N_811);
nand U9393 (N_9393,N_2001,N_3266);
nor U9394 (N_9394,N_4549,N_4583);
nand U9395 (N_9395,N_2378,N_4793);
nand U9396 (N_9396,N_717,N_807);
and U9397 (N_9397,N_2753,N_782);
or U9398 (N_9398,N_415,N_4100);
and U9399 (N_9399,N_1902,N_2720);
nor U9400 (N_9400,N_141,N_3973);
nor U9401 (N_9401,N_2759,N_274);
nand U9402 (N_9402,N_2055,N_3706);
nor U9403 (N_9403,N_586,N_3090);
or U9404 (N_9404,N_1054,N_2631);
or U9405 (N_9405,N_1505,N_579);
nand U9406 (N_9406,N_4978,N_4216);
and U9407 (N_9407,N_1296,N_1382);
and U9408 (N_9408,N_2017,N_2449);
or U9409 (N_9409,N_4296,N_2682);
and U9410 (N_9410,N_4114,N_4274);
or U9411 (N_9411,N_1616,N_1495);
and U9412 (N_9412,N_4776,N_78);
or U9413 (N_9413,N_3961,N_3324);
and U9414 (N_9414,N_1896,N_2684);
or U9415 (N_9415,N_2994,N_3547);
and U9416 (N_9416,N_2190,N_136);
or U9417 (N_9417,N_2302,N_66);
nor U9418 (N_9418,N_1918,N_4547);
nor U9419 (N_9419,N_3883,N_4487);
or U9420 (N_9420,N_3087,N_2385);
xor U9421 (N_9421,N_1589,N_4907);
or U9422 (N_9422,N_2579,N_2250);
and U9423 (N_9423,N_2949,N_3130);
nor U9424 (N_9424,N_234,N_2708);
xnor U9425 (N_9425,N_682,N_516);
and U9426 (N_9426,N_1299,N_3185);
or U9427 (N_9427,N_2605,N_4920);
or U9428 (N_9428,N_4686,N_4812);
nand U9429 (N_9429,N_4773,N_1074);
nor U9430 (N_9430,N_1270,N_328);
nand U9431 (N_9431,N_3895,N_2552);
and U9432 (N_9432,N_3476,N_92);
and U9433 (N_9433,N_4943,N_4498);
or U9434 (N_9434,N_2778,N_344);
nor U9435 (N_9435,N_3522,N_244);
nor U9436 (N_9436,N_4665,N_951);
nor U9437 (N_9437,N_4444,N_1394);
and U9438 (N_9438,N_1437,N_4194);
and U9439 (N_9439,N_2711,N_3090);
or U9440 (N_9440,N_2364,N_632);
or U9441 (N_9441,N_2781,N_867);
nor U9442 (N_9442,N_2543,N_2978);
and U9443 (N_9443,N_4389,N_4625);
nor U9444 (N_9444,N_487,N_225);
and U9445 (N_9445,N_1413,N_1627);
nand U9446 (N_9446,N_2509,N_3756);
and U9447 (N_9447,N_2671,N_4114);
or U9448 (N_9448,N_3081,N_4479);
nand U9449 (N_9449,N_108,N_1145);
and U9450 (N_9450,N_2700,N_4739);
nand U9451 (N_9451,N_1432,N_2445);
nand U9452 (N_9452,N_3033,N_186);
nor U9453 (N_9453,N_4508,N_4697);
or U9454 (N_9454,N_380,N_1053);
and U9455 (N_9455,N_1417,N_88);
or U9456 (N_9456,N_215,N_1694);
and U9457 (N_9457,N_1469,N_2185);
or U9458 (N_9458,N_652,N_2697);
and U9459 (N_9459,N_4028,N_3510);
and U9460 (N_9460,N_2522,N_4001);
nand U9461 (N_9461,N_405,N_3323);
and U9462 (N_9462,N_3364,N_3983);
nand U9463 (N_9463,N_1060,N_4566);
nor U9464 (N_9464,N_4774,N_1024);
and U9465 (N_9465,N_4926,N_1001);
or U9466 (N_9466,N_1525,N_791);
nand U9467 (N_9467,N_2961,N_2484);
or U9468 (N_9468,N_1440,N_2084);
nand U9469 (N_9469,N_501,N_2359);
and U9470 (N_9470,N_2902,N_3962);
and U9471 (N_9471,N_4938,N_1637);
nor U9472 (N_9472,N_1738,N_1153);
or U9473 (N_9473,N_3742,N_1859);
or U9474 (N_9474,N_4261,N_3780);
or U9475 (N_9475,N_964,N_4674);
and U9476 (N_9476,N_4201,N_872);
nand U9477 (N_9477,N_406,N_178);
nor U9478 (N_9478,N_17,N_212);
nor U9479 (N_9479,N_1796,N_379);
nor U9480 (N_9480,N_591,N_4759);
nand U9481 (N_9481,N_4378,N_2172);
nor U9482 (N_9482,N_3163,N_128);
nand U9483 (N_9483,N_408,N_2424);
and U9484 (N_9484,N_1626,N_2744);
nand U9485 (N_9485,N_173,N_4555);
and U9486 (N_9486,N_3227,N_3648);
and U9487 (N_9487,N_2665,N_1708);
xor U9488 (N_9488,N_2103,N_4314);
nor U9489 (N_9489,N_2360,N_2258);
xnor U9490 (N_9490,N_4293,N_4096);
or U9491 (N_9491,N_3834,N_2878);
and U9492 (N_9492,N_2791,N_498);
nor U9493 (N_9493,N_4523,N_4416);
or U9494 (N_9494,N_4752,N_4880);
nor U9495 (N_9495,N_2806,N_22);
and U9496 (N_9496,N_2919,N_2558);
nor U9497 (N_9497,N_4060,N_2484);
nand U9498 (N_9498,N_3866,N_1861);
and U9499 (N_9499,N_2994,N_372);
and U9500 (N_9500,N_641,N_1095);
and U9501 (N_9501,N_4444,N_4272);
and U9502 (N_9502,N_204,N_1901);
and U9503 (N_9503,N_1568,N_3531);
or U9504 (N_9504,N_2074,N_2897);
or U9505 (N_9505,N_2160,N_1499);
nor U9506 (N_9506,N_963,N_3239);
nand U9507 (N_9507,N_4990,N_4928);
nand U9508 (N_9508,N_390,N_532);
and U9509 (N_9509,N_1241,N_3016);
or U9510 (N_9510,N_2738,N_1258);
nand U9511 (N_9511,N_3175,N_1209);
and U9512 (N_9512,N_3204,N_2813);
or U9513 (N_9513,N_4188,N_2260);
nor U9514 (N_9514,N_3169,N_628);
or U9515 (N_9515,N_876,N_4673);
or U9516 (N_9516,N_4038,N_308);
nand U9517 (N_9517,N_2488,N_712);
or U9518 (N_9518,N_1978,N_1266);
nand U9519 (N_9519,N_1291,N_2581);
and U9520 (N_9520,N_3973,N_1558);
nand U9521 (N_9521,N_514,N_4746);
and U9522 (N_9522,N_1517,N_754);
or U9523 (N_9523,N_2624,N_984);
and U9524 (N_9524,N_3874,N_2467);
or U9525 (N_9525,N_265,N_2141);
nand U9526 (N_9526,N_1807,N_4821);
nand U9527 (N_9527,N_2464,N_4923);
nand U9528 (N_9528,N_2889,N_599);
and U9529 (N_9529,N_6,N_407);
nand U9530 (N_9530,N_2826,N_2335);
nor U9531 (N_9531,N_3230,N_3939);
nor U9532 (N_9532,N_3685,N_605);
or U9533 (N_9533,N_3991,N_4683);
or U9534 (N_9534,N_3029,N_2605);
or U9535 (N_9535,N_3418,N_2101);
or U9536 (N_9536,N_468,N_498);
nand U9537 (N_9537,N_4069,N_2339);
and U9538 (N_9538,N_4540,N_4377);
nand U9539 (N_9539,N_3929,N_4190);
or U9540 (N_9540,N_2658,N_450);
nand U9541 (N_9541,N_950,N_624);
or U9542 (N_9542,N_1908,N_1140);
and U9543 (N_9543,N_4510,N_146);
and U9544 (N_9544,N_1072,N_3422);
or U9545 (N_9545,N_525,N_2163);
and U9546 (N_9546,N_3781,N_442);
nor U9547 (N_9547,N_1301,N_4081);
nand U9548 (N_9548,N_3218,N_845);
nor U9549 (N_9549,N_1905,N_2687);
nand U9550 (N_9550,N_4971,N_2741);
and U9551 (N_9551,N_1650,N_3724);
nand U9552 (N_9552,N_4884,N_1550);
and U9553 (N_9553,N_4330,N_278);
nand U9554 (N_9554,N_397,N_3812);
or U9555 (N_9555,N_4789,N_1035);
nand U9556 (N_9556,N_1311,N_2897);
nand U9557 (N_9557,N_4666,N_1203);
nor U9558 (N_9558,N_3962,N_2602);
or U9559 (N_9559,N_4152,N_3973);
and U9560 (N_9560,N_2997,N_3352);
nor U9561 (N_9561,N_458,N_4472);
nand U9562 (N_9562,N_1386,N_1291);
or U9563 (N_9563,N_708,N_1959);
and U9564 (N_9564,N_1527,N_3111);
nor U9565 (N_9565,N_4282,N_4979);
and U9566 (N_9566,N_671,N_554);
or U9567 (N_9567,N_1010,N_32);
nand U9568 (N_9568,N_1521,N_65);
and U9569 (N_9569,N_3072,N_3046);
nor U9570 (N_9570,N_4594,N_1735);
nor U9571 (N_9571,N_1497,N_1659);
nor U9572 (N_9572,N_4799,N_1065);
or U9573 (N_9573,N_3987,N_295);
and U9574 (N_9574,N_1645,N_2447);
or U9575 (N_9575,N_1464,N_4912);
and U9576 (N_9576,N_845,N_2803);
and U9577 (N_9577,N_3833,N_2658);
and U9578 (N_9578,N_1578,N_11);
and U9579 (N_9579,N_4730,N_1986);
nor U9580 (N_9580,N_999,N_1657);
xor U9581 (N_9581,N_4916,N_2569);
and U9582 (N_9582,N_4460,N_3797);
nor U9583 (N_9583,N_3124,N_218);
nor U9584 (N_9584,N_3593,N_4637);
nand U9585 (N_9585,N_2074,N_123);
or U9586 (N_9586,N_161,N_3350);
nor U9587 (N_9587,N_678,N_3271);
nand U9588 (N_9588,N_837,N_2444);
and U9589 (N_9589,N_780,N_4539);
or U9590 (N_9590,N_3551,N_146);
and U9591 (N_9591,N_3843,N_3267);
or U9592 (N_9592,N_3102,N_1854);
or U9593 (N_9593,N_1852,N_2197);
nand U9594 (N_9594,N_1969,N_1310);
nand U9595 (N_9595,N_23,N_1344);
or U9596 (N_9596,N_355,N_85);
nor U9597 (N_9597,N_1496,N_1571);
and U9598 (N_9598,N_1958,N_868);
nor U9599 (N_9599,N_3682,N_2550);
nand U9600 (N_9600,N_4103,N_1728);
nor U9601 (N_9601,N_2138,N_4263);
nor U9602 (N_9602,N_1127,N_1566);
and U9603 (N_9603,N_1459,N_2561);
nor U9604 (N_9604,N_1868,N_4729);
nor U9605 (N_9605,N_4044,N_3667);
nand U9606 (N_9606,N_827,N_4137);
and U9607 (N_9607,N_1502,N_965);
or U9608 (N_9608,N_4556,N_1399);
nor U9609 (N_9609,N_81,N_4614);
nor U9610 (N_9610,N_2512,N_1141);
and U9611 (N_9611,N_2557,N_3474);
or U9612 (N_9612,N_443,N_2324);
nor U9613 (N_9613,N_2712,N_4897);
nand U9614 (N_9614,N_969,N_4327);
nor U9615 (N_9615,N_1862,N_2046);
nand U9616 (N_9616,N_4290,N_4378);
nand U9617 (N_9617,N_3507,N_2009);
nand U9618 (N_9618,N_89,N_4464);
nor U9619 (N_9619,N_2280,N_3715);
and U9620 (N_9620,N_201,N_2692);
nand U9621 (N_9621,N_1763,N_167);
nand U9622 (N_9622,N_1024,N_2243);
xnor U9623 (N_9623,N_3420,N_4897);
or U9624 (N_9624,N_4911,N_130);
or U9625 (N_9625,N_4758,N_4066);
or U9626 (N_9626,N_4388,N_390);
nand U9627 (N_9627,N_4874,N_936);
nand U9628 (N_9628,N_4479,N_4048);
and U9629 (N_9629,N_2569,N_4437);
or U9630 (N_9630,N_1283,N_3433);
xnor U9631 (N_9631,N_3919,N_2402);
and U9632 (N_9632,N_4438,N_1735);
nor U9633 (N_9633,N_4350,N_3136);
and U9634 (N_9634,N_3378,N_3423);
or U9635 (N_9635,N_3876,N_2494);
and U9636 (N_9636,N_2765,N_182);
and U9637 (N_9637,N_1170,N_2958);
nand U9638 (N_9638,N_1658,N_566);
or U9639 (N_9639,N_2494,N_3080);
nand U9640 (N_9640,N_3432,N_2493);
or U9641 (N_9641,N_537,N_3423);
or U9642 (N_9642,N_1036,N_2963);
or U9643 (N_9643,N_1477,N_3725);
or U9644 (N_9644,N_3609,N_4875);
nor U9645 (N_9645,N_2467,N_747);
or U9646 (N_9646,N_4513,N_3130);
nor U9647 (N_9647,N_453,N_4074);
nand U9648 (N_9648,N_1983,N_1653);
or U9649 (N_9649,N_4311,N_4090);
or U9650 (N_9650,N_2713,N_249);
xnor U9651 (N_9651,N_3857,N_1904);
nand U9652 (N_9652,N_543,N_3268);
nand U9653 (N_9653,N_1469,N_4565);
nor U9654 (N_9654,N_4935,N_3941);
and U9655 (N_9655,N_2688,N_3593);
nor U9656 (N_9656,N_334,N_1835);
and U9657 (N_9657,N_4756,N_1633);
or U9658 (N_9658,N_917,N_2386);
nand U9659 (N_9659,N_3528,N_1315);
or U9660 (N_9660,N_128,N_54);
or U9661 (N_9661,N_142,N_3352);
and U9662 (N_9662,N_148,N_4227);
nor U9663 (N_9663,N_2632,N_1972);
or U9664 (N_9664,N_1930,N_4574);
or U9665 (N_9665,N_3745,N_3665);
nand U9666 (N_9666,N_2258,N_3072);
nor U9667 (N_9667,N_825,N_4754);
and U9668 (N_9668,N_1287,N_2451);
nor U9669 (N_9669,N_4453,N_3163);
and U9670 (N_9670,N_2981,N_3979);
or U9671 (N_9671,N_3248,N_439);
nor U9672 (N_9672,N_4044,N_2463);
or U9673 (N_9673,N_2755,N_4444);
nand U9674 (N_9674,N_128,N_2010);
and U9675 (N_9675,N_2982,N_249);
nor U9676 (N_9676,N_3164,N_4795);
nand U9677 (N_9677,N_270,N_2130);
and U9678 (N_9678,N_4080,N_3106);
nand U9679 (N_9679,N_804,N_3423);
and U9680 (N_9680,N_4886,N_2348);
and U9681 (N_9681,N_3083,N_3776);
nor U9682 (N_9682,N_290,N_2566);
nor U9683 (N_9683,N_3314,N_1699);
and U9684 (N_9684,N_3033,N_1663);
nand U9685 (N_9685,N_2723,N_3137);
nand U9686 (N_9686,N_3616,N_2876);
nor U9687 (N_9687,N_1590,N_3191);
or U9688 (N_9688,N_3339,N_3097);
nand U9689 (N_9689,N_1182,N_2975);
nor U9690 (N_9690,N_97,N_2106);
nor U9691 (N_9691,N_1098,N_3097);
nor U9692 (N_9692,N_4526,N_2298);
nor U9693 (N_9693,N_4968,N_1385);
or U9694 (N_9694,N_3783,N_2637);
and U9695 (N_9695,N_3279,N_3392);
or U9696 (N_9696,N_2383,N_731);
nand U9697 (N_9697,N_162,N_4728);
or U9698 (N_9698,N_3953,N_3911);
nor U9699 (N_9699,N_309,N_508);
nand U9700 (N_9700,N_2038,N_2866);
or U9701 (N_9701,N_2787,N_3763);
and U9702 (N_9702,N_2310,N_1864);
and U9703 (N_9703,N_624,N_3122);
and U9704 (N_9704,N_2226,N_2165);
nand U9705 (N_9705,N_3152,N_2533);
or U9706 (N_9706,N_2804,N_544);
and U9707 (N_9707,N_3455,N_1895);
or U9708 (N_9708,N_3218,N_4993);
nor U9709 (N_9709,N_3370,N_4920);
nor U9710 (N_9710,N_1916,N_609);
nand U9711 (N_9711,N_2107,N_4809);
and U9712 (N_9712,N_1110,N_4163);
nor U9713 (N_9713,N_3962,N_2494);
nor U9714 (N_9714,N_2371,N_1216);
or U9715 (N_9715,N_4322,N_4772);
or U9716 (N_9716,N_2495,N_3872);
nand U9717 (N_9717,N_4299,N_912);
or U9718 (N_9718,N_388,N_4443);
nand U9719 (N_9719,N_2177,N_3321);
and U9720 (N_9720,N_1333,N_1786);
nor U9721 (N_9721,N_232,N_3034);
and U9722 (N_9722,N_3276,N_4911);
nand U9723 (N_9723,N_3834,N_2321);
and U9724 (N_9724,N_3533,N_2600);
nand U9725 (N_9725,N_3327,N_3126);
nand U9726 (N_9726,N_228,N_3265);
and U9727 (N_9727,N_2753,N_2836);
and U9728 (N_9728,N_3308,N_1861);
and U9729 (N_9729,N_3929,N_4623);
or U9730 (N_9730,N_3494,N_3830);
nor U9731 (N_9731,N_2036,N_2291);
nor U9732 (N_9732,N_1122,N_3658);
or U9733 (N_9733,N_4708,N_4008);
and U9734 (N_9734,N_604,N_3498);
or U9735 (N_9735,N_125,N_2189);
nor U9736 (N_9736,N_4866,N_3637);
nor U9737 (N_9737,N_790,N_851);
nor U9738 (N_9738,N_4285,N_1173);
nor U9739 (N_9739,N_1760,N_2627);
nor U9740 (N_9740,N_648,N_3096);
nor U9741 (N_9741,N_1248,N_2996);
or U9742 (N_9742,N_4675,N_3083);
nand U9743 (N_9743,N_4224,N_757);
nand U9744 (N_9744,N_3002,N_4011);
and U9745 (N_9745,N_3603,N_3695);
nor U9746 (N_9746,N_502,N_3428);
nor U9747 (N_9747,N_2786,N_1352);
nor U9748 (N_9748,N_2804,N_883);
nand U9749 (N_9749,N_1554,N_2891);
nor U9750 (N_9750,N_3568,N_560);
or U9751 (N_9751,N_4544,N_1061);
or U9752 (N_9752,N_1394,N_2517);
or U9753 (N_9753,N_4472,N_3913);
or U9754 (N_9754,N_564,N_1021);
nand U9755 (N_9755,N_4350,N_2151);
nand U9756 (N_9756,N_2364,N_1821);
and U9757 (N_9757,N_3383,N_1430);
nand U9758 (N_9758,N_4437,N_2042);
nor U9759 (N_9759,N_1530,N_4814);
nand U9760 (N_9760,N_4617,N_2565);
nand U9761 (N_9761,N_2447,N_3327);
or U9762 (N_9762,N_404,N_366);
nor U9763 (N_9763,N_3225,N_1264);
or U9764 (N_9764,N_475,N_4852);
xor U9765 (N_9765,N_859,N_4444);
and U9766 (N_9766,N_1798,N_3220);
nor U9767 (N_9767,N_2593,N_764);
nand U9768 (N_9768,N_869,N_736);
and U9769 (N_9769,N_659,N_1174);
or U9770 (N_9770,N_4490,N_1643);
and U9771 (N_9771,N_381,N_2161);
or U9772 (N_9772,N_3943,N_1163);
or U9773 (N_9773,N_402,N_4567);
or U9774 (N_9774,N_492,N_335);
xnor U9775 (N_9775,N_2746,N_3721);
and U9776 (N_9776,N_2119,N_268);
nand U9777 (N_9777,N_1471,N_3761);
nand U9778 (N_9778,N_4132,N_3020);
or U9779 (N_9779,N_41,N_1979);
or U9780 (N_9780,N_3188,N_324);
and U9781 (N_9781,N_2661,N_1550);
nor U9782 (N_9782,N_2486,N_2497);
nand U9783 (N_9783,N_87,N_3313);
nand U9784 (N_9784,N_2313,N_4423);
nand U9785 (N_9785,N_3221,N_4118);
nand U9786 (N_9786,N_518,N_3796);
and U9787 (N_9787,N_2180,N_4836);
nor U9788 (N_9788,N_1562,N_3855);
and U9789 (N_9789,N_3783,N_2066);
nor U9790 (N_9790,N_2957,N_669);
nand U9791 (N_9791,N_2891,N_1402);
nand U9792 (N_9792,N_337,N_225);
and U9793 (N_9793,N_1239,N_1339);
or U9794 (N_9794,N_1840,N_4113);
nand U9795 (N_9795,N_605,N_860);
and U9796 (N_9796,N_1520,N_4579);
nand U9797 (N_9797,N_2441,N_560);
or U9798 (N_9798,N_4787,N_568);
and U9799 (N_9799,N_4139,N_4392);
nor U9800 (N_9800,N_3297,N_4523);
nor U9801 (N_9801,N_2883,N_1825);
or U9802 (N_9802,N_654,N_336);
nand U9803 (N_9803,N_842,N_2687);
and U9804 (N_9804,N_253,N_3655);
or U9805 (N_9805,N_293,N_3487);
nand U9806 (N_9806,N_4706,N_4632);
nand U9807 (N_9807,N_2402,N_4372);
and U9808 (N_9808,N_597,N_2303);
nand U9809 (N_9809,N_1020,N_2599);
nor U9810 (N_9810,N_4124,N_786);
nor U9811 (N_9811,N_2929,N_2878);
nor U9812 (N_9812,N_4179,N_4442);
nor U9813 (N_9813,N_2621,N_3597);
nand U9814 (N_9814,N_2221,N_4006);
nor U9815 (N_9815,N_1443,N_967);
nand U9816 (N_9816,N_3952,N_4875);
nand U9817 (N_9817,N_137,N_3186);
nand U9818 (N_9818,N_4190,N_2643);
nand U9819 (N_9819,N_2334,N_2275);
nor U9820 (N_9820,N_2648,N_2078);
nor U9821 (N_9821,N_3698,N_3975);
xnor U9822 (N_9822,N_273,N_4568);
nor U9823 (N_9823,N_1821,N_1933);
and U9824 (N_9824,N_4832,N_3883);
nor U9825 (N_9825,N_4966,N_68);
nor U9826 (N_9826,N_2843,N_2454);
nor U9827 (N_9827,N_3788,N_1991);
or U9828 (N_9828,N_1494,N_836);
nand U9829 (N_9829,N_2537,N_4913);
and U9830 (N_9830,N_1134,N_1842);
nor U9831 (N_9831,N_662,N_1040);
nor U9832 (N_9832,N_2374,N_2463);
or U9833 (N_9833,N_4835,N_1776);
and U9834 (N_9834,N_629,N_794);
and U9835 (N_9835,N_1214,N_2994);
and U9836 (N_9836,N_4201,N_1650);
nand U9837 (N_9837,N_4975,N_3147);
or U9838 (N_9838,N_2917,N_4113);
and U9839 (N_9839,N_4362,N_4682);
nor U9840 (N_9840,N_134,N_4416);
and U9841 (N_9841,N_2122,N_4592);
or U9842 (N_9842,N_1525,N_4121);
or U9843 (N_9843,N_15,N_968);
or U9844 (N_9844,N_3888,N_3421);
and U9845 (N_9845,N_1665,N_3845);
nor U9846 (N_9846,N_4063,N_3216);
and U9847 (N_9847,N_2940,N_1100);
and U9848 (N_9848,N_1022,N_3469);
nand U9849 (N_9849,N_2230,N_4719);
or U9850 (N_9850,N_2856,N_2436);
and U9851 (N_9851,N_4294,N_2290);
nand U9852 (N_9852,N_3402,N_1393);
nand U9853 (N_9853,N_4640,N_2152);
nor U9854 (N_9854,N_3240,N_4241);
nand U9855 (N_9855,N_3800,N_1025);
nor U9856 (N_9856,N_1098,N_2330);
and U9857 (N_9857,N_1334,N_1985);
or U9858 (N_9858,N_546,N_1039);
nand U9859 (N_9859,N_4874,N_1334);
and U9860 (N_9860,N_678,N_3099);
nor U9861 (N_9861,N_2795,N_2265);
nor U9862 (N_9862,N_3210,N_512);
or U9863 (N_9863,N_1000,N_4146);
nor U9864 (N_9864,N_300,N_1918);
or U9865 (N_9865,N_2211,N_4268);
nor U9866 (N_9866,N_3860,N_922);
nand U9867 (N_9867,N_3688,N_4753);
nor U9868 (N_9868,N_708,N_4691);
nand U9869 (N_9869,N_3873,N_1008);
nor U9870 (N_9870,N_21,N_3361);
and U9871 (N_9871,N_3795,N_1419);
or U9872 (N_9872,N_1419,N_924);
nor U9873 (N_9873,N_3465,N_3805);
nand U9874 (N_9874,N_2497,N_3082);
or U9875 (N_9875,N_925,N_4650);
nor U9876 (N_9876,N_319,N_2320);
or U9877 (N_9877,N_4183,N_4047);
nor U9878 (N_9878,N_2256,N_4057);
and U9879 (N_9879,N_3847,N_1396);
or U9880 (N_9880,N_3469,N_3515);
or U9881 (N_9881,N_3290,N_3254);
xnor U9882 (N_9882,N_2156,N_4259);
nor U9883 (N_9883,N_1372,N_1625);
nand U9884 (N_9884,N_3609,N_4972);
nor U9885 (N_9885,N_383,N_4265);
or U9886 (N_9886,N_3136,N_4394);
nor U9887 (N_9887,N_3362,N_4050);
and U9888 (N_9888,N_4007,N_4345);
or U9889 (N_9889,N_3038,N_2306);
and U9890 (N_9890,N_1266,N_869);
nor U9891 (N_9891,N_4877,N_2608);
nor U9892 (N_9892,N_4002,N_3994);
and U9893 (N_9893,N_623,N_41);
or U9894 (N_9894,N_4968,N_3396);
nor U9895 (N_9895,N_1424,N_952);
or U9896 (N_9896,N_2937,N_2603);
nor U9897 (N_9897,N_4246,N_2148);
nand U9898 (N_9898,N_529,N_1258);
nand U9899 (N_9899,N_1549,N_1602);
nor U9900 (N_9900,N_1505,N_3920);
nand U9901 (N_9901,N_2191,N_1211);
nor U9902 (N_9902,N_3361,N_3754);
nor U9903 (N_9903,N_4915,N_3775);
and U9904 (N_9904,N_870,N_4104);
and U9905 (N_9905,N_692,N_3149);
or U9906 (N_9906,N_2762,N_740);
or U9907 (N_9907,N_3963,N_438);
nand U9908 (N_9908,N_697,N_524);
nand U9909 (N_9909,N_3941,N_2785);
nor U9910 (N_9910,N_2808,N_325);
and U9911 (N_9911,N_3491,N_1521);
nor U9912 (N_9912,N_4087,N_4650);
nor U9913 (N_9913,N_3290,N_3554);
nand U9914 (N_9914,N_4953,N_2464);
nor U9915 (N_9915,N_2586,N_2980);
nand U9916 (N_9916,N_929,N_106);
nand U9917 (N_9917,N_3025,N_2772);
or U9918 (N_9918,N_2711,N_4752);
or U9919 (N_9919,N_192,N_3375);
nand U9920 (N_9920,N_2810,N_4055);
and U9921 (N_9921,N_3322,N_4143);
or U9922 (N_9922,N_3490,N_198);
or U9923 (N_9923,N_1575,N_2180);
nor U9924 (N_9924,N_1595,N_91);
or U9925 (N_9925,N_1101,N_564);
nor U9926 (N_9926,N_174,N_2656);
nand U9927 (N_9927,N_3301,N_2052);
nand U9928 (N_9928,N_4743,N_1399);
nor U9929 (N_9929,N_3650,N_1272);
nor U9930 (N_9930,N_3715,N_4387);
nand U9931 (N_9931,N_1125,N_3749);
nand U9932 (N_9932,N_4346,N_4412);
nor U9933 (N_9933,N_2007,N_1149);
and U9934 (N_9934,N_576,N_648);
nor U9935 (N_9935,N_4379,N_1729);
and U9936 (N_9936,N_3408,N_1083);
or U9937 (N_9937,N_1486,N_3520);
and U9938 (N_9938,N_3362,N_1282);
nor U9939 (N_9939,N_669,N_3438);
or U9940 (N_9940,N_1891,N_2785);
xor U9941 (N_9941,N_4969,N_229);
or U9942 (N_9942,N_2621,N_4514);
or U9943 (N_9943,N_2109,N_2609);
and U9944 (N_9944,N_3442,N_4266);
or U9945 (N_9945,N_2581,N_2409);
nor U9946 (N_9946,N_1781,N_1266);
and U9947 (N_9947,N_832,N_3580);
or U9948 (N_9948,N_3202,N_148);
nand U9949 (N_9949,N_4936,N_1612);
nor U9950 (N_9950,N_1962,N_4750);
nand U9951 (N_9951,N_2598,N_1158);
and U9952 (N_9952,N_2417,N_1130);
nor U9953 (N_9953,N_1601,N_822);
nor U9954 (N_9954,N_2873,N_4079);
nor U9955 (N_9955,N_401,N_551);
or U9956 (N_9956,N_1494,N_448);
and U9957 (N_9957,N_812,N_1413);
or U9958 (N_9958,N_2214,N_101);
and U9959 (N_9959,N_4969,N_3398);
or U9960 (N_9960,N_2580,N_3522);
and U9961 (N_9961,N_984,N_663);
and U9962 (N_9962,N_967,N_2357);
nand U9963 (N_9963,N_766,N_4947);
nor U9964 (N_9964,N_3471,N_347);
nor U9965 (N_9965,N_649,N_1450);
and U9966 (N_9966,N_77,N_1865);
or U9967 (N_9967,N_1434,N_374);
or U9968 (N_9968,N_228,N_2679);
nand U9969 (N_9969,N_1053,N_678);
nand U9970 (N_9970,N_3967,N_1006);
or U9971 (N_9971,N_1428,N_3235);
or U9972 (N_9972,N_693,N_4746);
nand U9973 (N_9973,N_3237,N_2246);
nor U9974 (N_9974,N_1966,N_4813);
nor U9975 (N_9975,N_1648,N_215);
or U9976 (N_9976,N_3543,N_824);
nor U9977 (N_9977,N_2076,N_912);
or U9978 (N_9978,N_2328,N_2325);
and U9979 (N_9979,N_4713,N_482);
nand U9980 (N_9980,N_1218,N_4258);
nand U9981 (N_9981,N_1594,N_915);
or U9982 (N_9982,N_3086,N_3466);
and U9983 (N_9983,N_3569,N_3924);
and U9984 (N_9984,N_185,N_2230);
and U9985 (N_9985,N_2994,N_2400);
and U9986 (N_9986,N_3943,N_2154);
nor U9987 (N_9987,N_1292,N_1827);
and U9988 (N_9988,N_1558,N_2223);
or U9989 (N_9989,N_4564,N_3920);
nor U9990 (N_9990,N_690,N_4084);
or U9991 (N_9991,N_3216,N_2973);
or U9992 (N_9992,N_4636,N_779);
or U9993 (N_9993,N_142,N_1148);
nor U9994 (N_9994,N_1420,N_2143);
and U9995 (N_9995,N_3934,N_613);
and U9996 (N_9996,N_1413,N_4831);
and U9997 (N_9997,N_2489,N_2341);
or U9998 (N_9998,N_945,N_2961);
nor U9999 (N_9999,N_2591,N_3932);
nand UO_0 (O_0,N_9617,N_9918);
or UO_1 (O_1,N_8541,N_8101);
nand UO_2 (O_2,N_8463,N_5168);
nor UO_3 (O_3,N_7859,N_5446);
nand UO_4 (O_4,N_5321,N_6324);
or UO_5 (O_5,N_6274,N_8486);
and UO_6 (O_6,N_8628,N_8364);
nand UO_7 (O_7,N_7190,N_8376);
xnor UO_8 (O_8,N_7758,N_5827);
or UO_9 (O_9,N_6626,N_5891);
or UO_10 (O_10,N_5796,N_8894);
and UO_11 (O_11,N_5125,N_7608);
nor UO_12 (O_12,N_9357,N_6802);
and UO_13 (O_13,N_6267,N_8270);
or UO_14 (O_14,N_8654,N_7324);
nor UO_15 (O_15,N_6557,N_9407);
or UO_16 (O_16,N_9295,N_8638);
and UO_17 (O_17,N_8965,N_7193);
or UO_18 (O_18,N_9195,N_7399);
nor UO_19 (O_19,N_9866,N_5846);
nand UO_20 (O_20,N_7499,N_9704);
or UO_21 (O_21,N_9742,N_5972);
and UO_22 (O_22,N_8273,N_8271);
or UO_23 (O_23,N_5402,N_5589);
or UO_24 (O_24,N_5400,N_8586);
nand UO_25 (O_25,N_7341,N_9077);
nor UO_26 (O_26,N_5170,N_7586);
nand UO_27 (O_27,N_8526,N_9961);
and UO_28 (O_28,N_9960,N_9771);
nor UO_29 (O_29,N_9598,N_5723);
or UO_30 (O_30,N_9666,N_5099);
nand UO_31 (O_31,N_5555,N_6874);
or UO_32 (O_32,N_7055,N_7483);
and UO_33 (O_33,N_6656,N_6576);
and UO_34 (O_34,N_7185,N_7947);
and UO_35 (O_35,N_7099,N_5098);
and UO_36 (O_36,N_9735,N_7290);
nand UO_37 (O_37,N_6131,N_7302);
and UO_38 (O_38,N_8839,N_9684);
or UO_39 (O_39,N_5887,N_5287);
and UO_40 (O_40,N_8266,N_7613);
or UO_41 (O_41,N_9507,N_9629);
or UO_42 (O_42,N_6484,N_7315);
nand UO_43 (O_43,N_8931,N_5829);
or UO_44 (O_44,N_7899,N_8967);
or UO_45 (O_45,N_7760,N_9221);
or UO_46 (O_46,N_6581,N_9733);
nor UO_47 (O_47,N_7125,N_5705);
or UO_48 (O_48,N_5883,N_7982);
nor UO_49 (O_49,N_8168,N_8972);
xnor UO_50 (O_50,N_6548,N_9972);
nor UO_51 (O_51,N_9651,N_7590);
and UO_52 (O_52,N_8567,N_5305);
and UO_53 (O_53,N_6586,N_5495);
or UO_54 (O_54,N_6280,N_9418);
nor UO_55 (O_55,N_5938,N_9243);
and UO_56 (O_56,N_9159,N_9180);
and UO_57 (O_57,N_7391,N_5593);
or UO_58 (O_58,N_9571,N_9103);
nand UO_59 (O_59,N_8989,N_8629);
nand UO_60 (O_60,N_5571,N_9572);
and UO_61 (O_61,N_7879,N_8464);
or UO_62 (O_62,N_6781,N_7766);
nand UO_63 (O_63,N_6887,N_5376);
nand UO_64 (O_64,N_9309,N_7034);
nand UO_65 (O_65,N_8620,N_8410);
and UO_66 (O_66,N_5563,N_5022);
nand UO_67 (O_67,N_5508,N_5897);
nand UO_68 (O_68,N_7756,N_8532);
nor UO_69 (O_69,N_9577,N_9130);
and UO_70 (O_70,N_5033,N_5173);
nand UO_71 (O_71,N_7460,N_6596);
nor UO_72 (O_72,N_6703,N_8911);
nor UO_73 (O_73,N_6620,N_7116);
nand UO_74 (O_74,N_7439,N_9658);
nand UO_75 (O_75,N_5194,N_7227);
nand UO_76 (O_76,N_5175,N_6789);
nand UO_77 (O_77,N_8724,N_9226);
nand UO_78 (O_78,N_5227,N_7726);
and UO_79 (O_79,N_6224,N_8071);
nor UO_80 (O_80,N_6774,N_9475);
and UO_81 (O_81,N_8878,N_6796);
and UO_82 (O_82,N_8535,N_8513);
nand UO_83 (O_83,N_7910,N_8889);
and UO_84 (O_84,N_9211,N_7925);
or UO_85 (O_85,N_7102,N_7408);
or UO_86 (O_86,N_8781,N_9324);
nor UO_87 (O_87,N_6508,N_8505);
nand UO_88 (O_88,N_6634,N_7486);
nand UO_89 (O_89,N_7043,N_5832);
and UO_90 (O_90,N_6697,N_8664);
nor UO_91 (O_91,N_5306,N_6725);
nand UO_92 (O_92,N_6378,N_8073);
nand UO_93 (O_93,N_7968,N_5439);
nor UO_94 (O_94,N_6441,N_6692);
nor UO_95 (O_95,N_8793,N_6005);
nand UO_96 (O_96,N_6260,N_9959);
or UO_97 (O_97,N_9163,N_8250);
or UO_98 (O_98,N_7208,N_6010);
and UO_99 (O_99,N_6716,N_6648);
or UO_100 (O_100,N_8375,N_5190);
or UO_101 (O_101,N_7348,N_7442);
and UO_102 (O_102,N_5754,N_8487);
and UO_103 (O_103,N_8278,N_6522);
nor UO_104 (O_104,N_6875,N_5310);
nor UO_105 (O_105,N_9857,N_5279);
nand UO_106 (O_106,N_9583,N_5152);
nor UO_107 (O_107,N_7216,N_5521);
nand UO_108 (O_108,N_6353,N_7707);
nand UO_109 (O_109,N_6934,N_7334);
or UO_110 (O_110,N_5119,N_6138);
or UO_111 (O_111,N_9852,N_7914);
nor UO_112 (O_112,N_9930,N_6202);
or UO_113 (O_113,N_7830,N_9779);
nor UO_114 (O_114,N_8838,N_8117);
nor UO_115 (O_115,N_7904,N_5730);
nand UO_116 (O_116,N_8444,N_6011);
nor UO_117 (O_117,N_7274,N_6915);
nand UO_118 (O_118,N_9308,N_9848);
and UO_119 (O_119,N_8470,N_9619);
nor UO_120 (O_120,N_8699,N_7962);
nand UO_121 (O_121,N_7413,N_8539);
and UO_122 (O_122,N_8493,N_8466);
and UO_123 (O_123,N_7307,N_8885);
nor UO_124 (O_124,N_8515,N_8194);
nand UO_125 (O_125,N_6564,N_6180);
nand UO_126 (O_126,N_9956,N_5676);
nor UO_127 (O_127,N_5468,N_7073);
and UO_128 (O_128,N_5387,N_8384);
and UO_129 (O_129,N_5879,N_5256);
or UO_130 (O_130,N_5381,N_7054);
or UO_131 (O_131,N_8106,N_5795);
or UO_132 (O_132,N_8239,N_7838);
nor UO_133 (O_133,N_7459,N_8852);
nor UO_134 (O_134,N_7430,N_5612);
or UO_135 (O_135,N_5659,N_6719);
and UO_136 (O_136,N_6676,N_7386);
or UO_137 (O_137,N_6165,N_7207);
nor UO_138 (O_138,N_8434,N_6357);
and UO_139 (O_139,N_8000,N_9647);
and UO_140 (O_140,N_6503,N_8481);
nand UO_141 (O_141,N_8743,N_8403);
nand UO_142 (O_142,N_5020,N_5813);
nor UO_143 (O_143,N_8844,N_5300);
nand UO_144 (O_144,N_7471,N_7365);
nand UO_145 (O_145,N_9714,N_9068);
nand UO_146 (O_146,N_9729,N_8834);
nand UO_147 (O_147,N_6426,N_9654);
nor UO_148 (O_148,N_5939,N_8879);
and UO_149 (O_149,N_9002,N_5538);
nor UO_150 (O_150,N_7031,N_9313);
and UO_151 (O_151,N_7071,N_6848);
xor UO_152 (O_152,N_9081,N_8676);
or UO_153 (O_153,N_5875,N_9410);
nand UO_154 (O_154,N_6297,N_8409);
nor UO_155 (O_155,N_8886,N_8075);
nor UO_156 (O_156,N_5774,N_5814);
or UO_157 (O_157,N_7177,N_7346);
nor UO_158 (O_158,N_7600,N_7523);
and UO_159 (O_159,N_7870,N_5716);
and UO_160 (O_160,N_9037,N_8225);
nand UO_161 (O_161,N_9281,N_5100);
or UO_162 (O_162,N_5789,N_9982);
or UO_163 (O_163,N_6625,N_7111);
nor UO_164 (O_164,N_5569,N_7584);
or UO_165 (O_165,N_8749,N_8891);
nor UO_166 (O_166,N_7735,N_6452);
nor UO_167 (O_167,N_6575,N_5710);
or UO_168 (O_168,N_5664,N_9765);
or UO_169 (O_169,N_8241,N_6955);
or UO_170 (O_170,N_9371,N_9758);
or UO_171 (O_171,N_6938,N_6006);
or UO_172 (O_172,N_9707,N_9656);
nand UO_173 (O_173,N_5613,N_9799);
and UO_174 (O_174,N_6619,N_6531);
nor UO_175 (O_175,N_5463,N_5103);
or UO_176 (O_176,N_5665,N_9540);
nand UO_177 (O_177,N_6336,N_7350);
nor UO_178 (O_178,N_7538,N_9715);
nand UO_179 (O_179,N_6122,N_8167);
nand UO_180 (O_180,N_6231,N_5097);
or UO_181 (O_181,N_7980,N_6245);
and UO_182 (O_182,N_8305,N_7298);
nor UO_183 (O_183,N_9178,N_5385);
or UO_184 (O_184,N_8746,N_7814);
nand UO_185 (O_185,N_8517,N_6356);
and UO_186 (O_186,N_7537,N_6407);
and UO_187 (O_187,N_6904,N_8415);
nand UO_188 (O_188,N_8276,N_8129);
and UO_189 (O_189,N_8530,N_8518);
or UO_190 (O_190,N_5161,N_8359);
nor UO_191 (O_191,N_6886,N_9905);
nor UO_192 (O_192,N_6445,N_7355);
and UO_193 (O_193,N_7509,N_5630);
nor UO_194 (O_194,N_7567,N_6504);
or UO_195 (O_195,N_8870,N_5285);
nand UO_196 (O_196,N_9929,N_8576);
nor UO_197 (O_197,N_9471,N_6382);
nand UO_198 (O_198,N_8590,N_9067);
nor UO_199 (O_199,N_5977,N_8902);
nand UO_200 (O_200,N_8607,N_5819);
nand UO_201 (O_201,N_8748,N_6398);
and UO_202 (O_202,N_7998,N_5627);
or UO_203 (O_203,N_9196,N_8303);
and UO_204 (O_204,N_6119,N_8286);
or UO_205 (O_205,N_8367,N_7051);
nor UO_206 (O_206,N_8501,N_7654);
or UO_207 (O_207,N_7546,N_5023);
or UO_208 (O_208,N_9635,N_5148);
nor UO_209 (O_209,N_7070,N_9479);
and UO_210 (O_210,N_7137,N_8301);
xnor UO_211 (O_211,N_5900,N_9209);
and UO_212 (O_212,N_7715,N_9529);
and UO_213 (O_213,N_9708,N_6271);
nand UO_214 (O_214,N_9155,N_7616);
and UO_215 (O_215,N_9939,N_8933);
nand UO_216 (O_216,N_9794,N_8385);
nand UO_217 (O_217,N_8491,N_7564);
nor UO_218 (O_218,N_8121,N_6281);
and UO_219 (O_219,N_9753,N_9859);
nand UO_220 (O_220,N_8943,N_6709);
nand UO_221 (O_221,N_6594,N_6704);
or UO_222 (O_222,N_5492,N_8059);
nor UO_223 (O_223,N_5480,N_6374);
nor UO_224 (O_224,N_5982,N_8740);
and UO_225 (O_225,N_6239,N_7625);
and UO_226 (O_226,N_8881,N_7003);
nor UO_227 (O_227,N_6219,N_5541);
nor UO_228 (O_228,N_7222,N_9431);
nand UO_229 (O_229,N_7176,N_6695);
nand UO_230 (O_230,N_5505,N_7196);
and UO_231 (O_231,N_6027,N_7474);
nor UO_232 (O_232,N_7607,N_6609);
nor UO_233 (O_233,N_8206,N_9193);
nand UO_234 (O_234,N_5224,N_9136);
nand UO_235 (O_235,N_7440,N_8826);
and UO_236 (O_236,N_6817,N_8701);
or UO_237 (O_237,N_9833,N_9473);
or UO_238 (O_238,N_7557,N_7542);
or UO_239 (O_239,N_6921,N_8296);
and UO_240 (O_240,N_5136,N_5257);
nor UO_241 (O_241,N_6605,N_7017);
nor UO_242 (O_242,N_6543,N_7993);
and UO_243 (O_243,N_7595,N_9916);
nor UO_244 (O_244,N_5978,N_7646);
nor UO_245 (O_245,N_7873,N_5767);
and UO_246 (O_246,N_6135,N_6276);
and UO_247 (O_247,N_6468,N_8437);
and UO_248 (O_248,N_7952,N_5297);
and UO_249 (O_249,N_9146,N_8723);
nor UO_250 (O_250,N_7249,N_7284);
and UO_251 (O_251,N_7175,N_8521);
or UO_252 (O_252,N_5961,N_7181);
nor UO_253 (O_253,N_9141,N_9219);
or UO_254 (O_254,N_7576,N_8649);
or UO_255 (O_255,N_6460,N_7012);
and UO_256 (O_256,N_8761,N_7833);
or UO_257 (O_257,N_9908,N_7242);
nor UO_258 (O_258,N_5466,N_8002);
nand UO_259 (O_259,N_9400,N_9108);
and UO_260 (O_260,N_9311,N_5561);
and UO_261 (O_261,N_8419,N_7064);
and UO_262 (O_262,N_6065,N_7895);
nor UO_263 (O_263,N_9695,N_5373);
or UO_264 (O_264,N_8231,N_6649);
and UO_265 (O_265,N_9125,N_5549);
or UO_266 (O_266,N_7695,N_8549);
and UO_267 (O_267,N_9781,N_7352);
and UO_268 (O_268,N_7347,N_6777);
or UO_269 (O_269,N_7067,N_6246);
and UO_270 (O_270,N_7513,N_6477);
nand UO_271 (O_271,N_6261,N_9274);
or UO_272 (O_272,N_9924,N_9596);
or UO_273 (O_273,N_5512,N_7087);
nand UO_274 (O_274,N_8494,N_8163);
and UO_275 (O_275,N_8402,N_9297);
or UO_276 (O_276,N_7907,N_9456);
nand UO_277 (O_277,N_9417,N_6410);
or UO_278 (O_278,N_8265,N_9256);
and UO_279 (O_279,N_6370,N_5479);
or UO_280 (O_280,N_6125,N_5501);
or UO_281 (O_281,N_7632,N_9296);
and UO_282 (O_282,N_5974,N_5631);
or UO_283 (O_283,N_6818,N_9249);
and UO_284 (O_284,N_5391,N_7572);
nor UO_285 (O_285,N_9926,N_6804);
and UO_286 (O_286,N_8057,N_9592);
and UO_287 (O_287,N_6783,N_5014);
or UO_288 (O_288,N_9277,N_8908);
and UO_289 (O_289,N_7198,N_9528);
nor UO_290 (O_290,N_7319,N_5700);
nor UO_291 (O_291,N_5526,N_5874);
nor UO_292 (O_292,N_9156,N_8139);
nand UO_293 (O_293,N_9705,N_7209);
nor UO_294 (O_294,N_9639,N_5335);
or UO_295 (O_295,N_9828,N_9406);
nand UO_296 (O_296,N_5812,N_8828);
nand UO_297 (O_297,N_5447,N_6545);
nand UO_298 (O_298,N_7581,N_8441);
nor UO_299 (O_299,N_7157,N_8019);
and UO_300 (O_300,N_6330,N_5678);
nand UO_301 (O_301,N_9028,N_9754);
nand UO_302 (O_302,N_5139,N_8288);
nor UO_303 (O_303,N_7610,N_9603);
nand UO_304 (O_304,N_7018,N_8929);
or UO_305 (O_305,N_6113,N_9320);
nand UO_306 (O_306,N_6092,N_5497);
or UO_307 (O_307,N_7566,N_7687);
or UO_308 (O_308,N_9590,N_8246);
or UO_309 (O_309,N_6063,N_6186);
or UO_310 (O_310,N_8986,N_6474);
nor UO_311 (O_311,N_9760,N_9743);
nand UO_312 (O_312,N_8680,N_8910);
nor UO_313 (O_313,N_8528,N_9750);
or UO_314 (O_314,N_7390,N_8609);
or UO_315 (O_315,N_6559,N_9537);
and UO_316 (O_316,N_8783,N_8604);
or UO_317 (O_317,N_5338,N_6034);
or UO_318 (O_318,N_7144,N_5433);
or UO_319 (O_319,N_9120,N_7432);
or UO_320 (O_320,N_6435,N_9553);
nor UO_321 (O_321,N_9096,N_7972);
and UO_322 (O_322,N_7162,N_7349);
nand UO_323 (O_323,N_9716,N_5046);
or UO_324 (O_324,N_5482,N_7053);
nor UO_325 (O_325,N_9845,N_6813);
nor UO_326 (O_326,N_8416,N_6222);
and UO_327 (O_327,N_5250,N_5339);
nor UO_328 (O_328,N_5089,N_7955);
nand UO_329 (O_329,N_9662,N_7010);
or UO_330 (O_330,N_7373,N_8674);
and UO_331 (O_331,N_9800,N_7517);
or UO_332 (O_332,N_6950,N_8906);
or UO_333 (O_333,N_5616,N_5210);
and UO_334 (O_334,N_8217,N_8390);
and UO_335 (O_335,N_5126,N_7097);
and UO_336 (O_336,N_5513,N_5365);
nor UO_337 (O_337,N_6419,N_7936);
nand UO_338 (O_338,N_8824,N_9841);
nand UO_339 (O_339,N_8076,N_5719);
nand UO_340 (O_340,N_8312,N_9310);
and UO_341 (O_341,N_5601,N_6442);
nor UO_342 (O_342,N_5945,N_5000);
nor UO_343 (O_343,N_5451,N_6612);
or UO_344 (O_344,N_6486,N_7123);
and UO_345 (O_345,N_9575,N_7147);
or UO_346 (O_346,N_5069,N_9838);
and UO_347 (O_347,N_7820,N_5470);
and UO_348 (O_348,N_8603,N_6106);
and UO_349 (O_349,N_9027,N_9558);
nand UO_350 (O_350,N_5314,N_5452);
and UO_351 (O_351,N_5048,N_5861);
nor UO_352 (O_352,N_5346,N_9892);
nand UO_353 (O_353,N_5718,N_6029);
nand UO_354 (O_354,N_6475,N_7536);
and UO_355 (O_355,N_7637,N_8594);
nor UO_356 (O_356,N_8924,N_9913);
nor UO_357 (O_357,N_6583,N_7287);
nand UO_358 (O_358,N_6025,N_7964);
and UO_359 (O_359,N_8600,N_6761);
or UO_360 (O_360,N_8540,N_6590);
nor UO_361 (O_361,N_6850,N_5378);
nand UO_362 (O_362,N_8457,N_8363);
nor UO_363 (O_363,N_5764,N_6220);
nand UO_364 (O_364,N_7827,N_8936);
and UO_365 (O_365,N_8326,N_7488);
or UO_366 (O_366,N_9582,N_5539);
and UO_367 (O_367,N_9440,N_6792);
nand UO_368 (O_368,N_5588,N_7154);
xor UO_369 (O_369,N_7730,N_7612);
xnor UO_370 (O_370,N_5362,N_6665);
nand UO_371 (O_371,N_9951,N_7890);
and UO_372 (O_372,N_8962,N_5193);
nand UO_373 (O_373,N_7640,N_9021);
nand UO_374 (O_374,N_5773,N_7478);
nor UO_375 (O_375,N_9175,N_6595);
and UO_376 (O_376,N_7400,N_5850);
or UO_377 (O_377,N_5454,N_7623);
nor UO_378 (O_378,N_8332,N_6121);
or UO_379 (O_379,N_6973,N_7950);
nand UO_380 (O_380,N_9361,N_5049);
nor UO_381 (O_381,N_9183,N_9761);
nor UO_382 (O_382,N_6942,N_9349);
nand UO_383 (O_383,N_5399,N_6898);
nor UO_384 (O_384,N_6133,N_5301);
nand UO_385 (O_385,N_9258,N_7344);
nand UO_386 (O_386,N_5295,N_9791);
or UO_387 (O_387,N_6288,N_8072);
nor UO_388 (O_388,N_8978,N_9774);
nor UO_389 (O_389,N_5707,N_9009);
or UO_390 (O_390,N_6439,N_7452);
nand UO_391 (O_391,N_8811,N_9341);
and UO_392 (O_392,N_5576,N_9726);
or UO_393 (O_393,N_5890,N_8439);
and UO_394 (O_394,N_6462,N_8477);
or UO_395 (O_395,N_6570,N_6616);
nand UO_396 (O_396,N_9114,N_8968);
nor UO_397 (O_397,N_6929,N_7529);
nand UO_398 (O_398,N_9401,N_5870);
nor UO_399 (O_399,N_5318,N_5394);
nand UO_400 (O_400,N_7024,N_5776);
or UO_401 (O_401,N_5502,N_5230);
or UO_402 (O_402,N_8938,N_7038);
and UO_403 (O_403,N_8435,N_7634);
or UO_404 (O_404,N_5107,N_7056);
nand UO_405 (O_405,N_9446,N_9054);
nor UO_406 (O_406,N_7363,N_6427);
or UO_407 (O_407,N_9749,N_5980);
and UO_408 (O_408,N_9262,N_7280);
nor UO_409 (O_409,N_9556,N_9441);
xnor UO_410 (O_410,N_5232,N_9105);
or UO_411 (O_411,N_9300,N_9057);
nand UO_412 (O_412,N_7113,N_7001);
or UO_413 (O_413,N_7960,N_9517);
or UO_414 (O_414,N_9673,N_5903);
and UO_415 (O_415,N_8392,N_5461);
nand UO_416 (O_416,N_8144,N_7694);
or UO_417 (O_417,N_5281,N_9991);
nand UO_418 (O_418,N_8670,N_5895);
or UO_419 (O_419,N_9513,N_7301);
nor UO_420 (O_420,N_5729,N_5464);
and UO_421 (O_421,N_6322,N_8450);
and UO_422 (O_422,N_7167,N_5650);
and UO_423 (O_423,N_9024,N_5457);
and UO_424 (O_424,N_5715,N_5003);
nand UO_425 (O_425,N_5264,N_8346);
or UO_426 (O_426,N_7809,N_8658);
nand UO_427 (O_427,N_8056,N_9861);
and UO_428 (O_428,N_6146,N_5834);
nor UO_429 (O_429,N_9805,N_8316);
nand UO_430 (O_430,N_9071,N_9784);
or UO_431 (O_431,N_9897,N_5652);
nand UO_432 (O_432,N_5633,N_7443);
and UO_433 (O_433,N_8903,N_5954);
nand UO_434 (O_434,N_8928,N_8030);
or UO_435 (O_435,N_8560,N_8127);
or UO_436 (O_436,N_5516,N_5288);
nor UO_437 (O_437,N_9177,N_9316);
and UO_438 (O_438,N_9957,N_9188);
or UO_439 (O_439,N_9672,N_6300);
and UO_440 (O_440,N_5149,N_6728);
nand UO_441 (O_441,N_5607,N_5236);
nand UO_442 (O_442,N_5941,N_9215);
and UO_443 (O_443,N_8920,N_9107);
nand UO_444 (O_444,N_6688,N_6362);
nor UO_445 (O_445,N_7680,N_5626);
and UO_446 (O_446,N_8111,N_8134);
xnor UO_447 (O_447,N_7849,N_7655);
or UO_448 (O_448,N_5772,N_6217);
nor UO_449 (O_449,N_7729,N_6748);
nand UO_450 (O_450,N_5422,N_6572);
or UO_451 (O_451,N_8880,N_6775);
or UO_452 (O_452,N_8883,N_7676);
or UO_453 (O_453,N_6153,N_7638);
nor UO_454 (O_454,N_9523,N_9533);
and UO_455 (O_455,N_7651,N_7913);
and UO_456 (O_456,N_8492,N_6831);
nor UO_457 (O_457,N_5159,N_9377);
or UO_458 (O_458,N_7482,N_5746);
or UO_459 (O_459,N_8417,N_7690);
nor UO_460 (O_460,N_6808,N_8692);
nand UO_461 (O_461,N_6284,N_5927);
nor UO_462 (O_462,N_8706,N_9364);
nor UO_463 (O_463,N_6126,N_5490);
nor UO_464 (O_464,N_8079,N_5517);
nor UO_465 (O_465,N_6499,N_7807);
or UO_466 (O_466,N_5253,N_7911);
and UO_467 (O_467,N_6747,N_5481);
and UO_468 (O_468,N_5839,N_5775);
or UO_469 (O_469,N_6601,N_7932);
nor UO_470 (O_470,N_7258,N_9661);
or UO_471 (O_471,N_6345,N_5459);
or UO_472 (O_472,N_9778,N_8480);
xnor UO_473 (O_473,N_9664,N_8370);
nor UO_474 (O_474,N_5684,N_9542);
nand UO_475 (O_475,N_7130,N_8065);
or UO_476 (O_476,N_9643,N_6629);
nor UO_477 (O_477,N_7543,N_8133);
nand UO_478 (O_478,N_5228,N_5742);
and UO_479 (O_479,N_6105,N_6036);
nor UO_480 (O_480,N_5367,N_8110);
nand UO_481 (O_481,N_5114,N_5043);
or UO_482 (O_482,N_6204,N_7896);
or UO_483 (O_483,N_7383,N_9538);
or UO_484 (O_484,N_8284,N_9531);
nor UO_485 (O_485,N_8559,N_5327);
nand UO_486 (O_486,N_8090,N_8511);
nand UO_487 (O_487,N_8702,N_5044);
or UO_488 (O_488,N_7540,N_8190);
nor UO_489 (O_489,N_7839,N_5535);
or UO_490 (O_490,N_5120,N_9690);
nand UO_491 (O_491,N_7412,N_9266);
nand UO_492 (O_492,N_9140,N_8814);
and UO_493 (O_493,N_9786,N_9802);
nand UO_494 (O_494,N_7021,N_7455);
or UO_495 (O_495,N_6917,N_5453);
and UO_496 (O_496,N_8961,N_5265);
nand UO_497 (O_497,N_7406,N_6582);
nor UO_498 (O_498,N_7205,N_7518);
or UO_499 (O_499,N_5074,N_5604);
or UO_500 (O_500,N_5291,N_5837);
and UO_501 (O_501,N_5025,N_8488);
or UO_502 (O_502,N_7372,N_9070);
nand UO_503 (O_503,N_9932,N_5144);
nand UO_504 (O_504,N_9813,N_8525);
nand UO_505 (O_505,N_5406,N_7132);
and UO_506 (O_506,N_7182,N_5423);
nor UO_507 (O_507,N_8484,N_8596);
or UO_508 (O_508,N_9046,N_7796);
and UO_509 (O_509,N_7402,N_7325);
or UO_510 (O_510,N_7493,N_8672);
and UO_511 (O_511,N_5866,N_7906);
nand UO_512 (O_512,N_5268,N_5559);
nand UO_513 (O_513,N_5375,N_5197);
nor UO_514 (O_514,N_7016,N_8784);
or UO_515 (O_515,N_6263,N_9245);
and UO_516 (O_516,N_9969,N_6226);
nand UO_517 (O_517,N_5262,N_8461);
and UO_518 (O_518,N_9712,N_6323);
or UO_519 (O_519,N_7520,N_6303);
xnor UO_520 (O_520,N_7541,N_6355);
and UO_521 (O_521,N_6638,N_5552);
and UO_522 (O_522,N_8454,N_6966);
and UO_523 (O_523,N_5644,N_6578);
nor UO_524 (O_524,N_7554,N_6529);
nor UO_525 (O_525,N_7791,N_9711);
or UO_526 (O_526,N_8971,N_8342);
nand UO_527 (O_527,N_7203,N_6054);
nor UO_528 (O_528,N_6311,N_6843);
nor UO_529 (O_529,N_6320,N_7742);
nand UO_530 (O_530,N_9593,N_9906);
nor UO_531 (O_531,N_5309,N_7370);
nand UO_532 (O_532,N_9472,N_5759);
nand UO_533 (O_533,N_8950,N_9880);
nor UO_534 (O_534,N_6163,N_7059);
or UO_535 (O_535,N_6306,N_9220);
nor UO_536 (O_536,N_5611,N_6599);
and UO_537 (O_537,N_6053,N_6307);
or UO_538 (O_538,N_7553,N_6782);
nor UO_539 (O_539,N_8423,N_7987);
nand UO_540 (O_540,N_6314,N_5987);
and UO_541 (O_541,N_7605,N_5821);
nor UO_542 (O_542,N_8613,N_5350);
and UO_543 (O_543,N_5902,N_7418);
nand UO_544 (O_544,N_8038,N_5838);
nor UO_545 (O_545,N_7573,N_9263);
nand UO_546 (O_546,N_6720,N_7263);
and UO_547 (O_547,N_9580,N_6839);
nand UO_548 (O_548,N_6633,N_6571);
and UO_549 (O_549,N_5360,N_5935);
or UO_550 (O_550,N_7971,N_5205);
and UO_551 (O_551,N_9270,N_6936);
nand UO_552 (O_552,N_7155,N_8745);
nor UO_553 (O_553,N_6050,N_7958);
nor UO_554 (O_554,N_6088,N_9010);
nor UO_555 (O_555,N_6655,N_5782);
nor UO_556 (O_556,N_7531,N_6534);
and UO_557 (O_557,N_7069,N_5275);
and UO_558 (O_558,N_7746,N_6235);
and UO_559 (O_559,N_8799,N_5693);
nor UO_560 (O_560,N_9445,N_7744);
nor UO_561 (O_561,N_8837,N_8094);
and UO_562 (O_562,N_8907,N_9139);
and UO_563 (O_563,N_7140,N_8563);
nor UO_564 (O_564,N_6338,N_5888);
or UO_565 (O_565,N_7211,N_8136);
or UO_566 (O_566,N_7515,N_7674);
or UO_567 (O_567,N_6147,N_8285);
nand UO_568 (O_568,N_9030,N_8218);
or UO_569 (O_569,N_5817,N_7570);
nand UO_570 (O_570,N_6549,N_5818);
nor UO_571 (O_571,N_5184,N_6089);
nor UO_572 (O_572,N_5862,N_7392);
and UO_573 (O_573,N_8703,N_9963);
nand UO_574 (O_574,N_6193,N_9005);
nand UO_575 (O_575,N_9484,N_9135);
nor UO_576 (O_576,N_8275,N_7832);
and UO_577 (O_577,N_7108,N_6325);
nor UO_578 (O_578,N_8349,N_5856);
and UO_579 (O_579,N_7453,N_7858);
and UO_580 (O_580,N_5249,N_9398);
nand UO_581 (O_581,N_5229,N_8498);
or UO_582 (O_582,N_8710,N_5021);
nand UO_583 (O_583,N_9231,N_8923);
and UO_584 (O_584,N_8188,N_5868);
or UO_585 (O_585,N_9217,N_5050);
and UO_586 (O_586,N_6383,N_8716);
or UO_587 (O_587,N_9881,N_5226);
nand UO_588 (O_588,N_6997,N_8489);
nand UO_589 (O_589,N_7969,N_6537);
and UO_590 (O_590,N_7359,N_7732);
nand UO_591 (O_591,N_8728,N_5147);
or UO_592 (O_592,N_6563,N_9518);
nor UO_593 (O_593,N_6472,N_7984);
and UO_594 (O_594,N_8172,N_5810);
and UO_595 (O_595,N_5597,N_5735);
nor UO_596 (O_596,N_6256,N_6677);
and UO_597 (O_597,N_8998,N_6883);
and UO_598 (O_598,N_5386,N_9477);
or UO_599 (O_599,N_8502,N_6807);
and UO_600 (O_600,N_7533,N_6520);
nor UO_601 (O_601,N_6067,N_9115);
or UO_602 (O_602,N_8531,N_8195);
nor UO_603 (O_603,N_6448,N_9796);
nand UO_604 (O_604,N_7909,N_6873);
nor UO_605 (O_605,N_8325,N_8918);
and UO_606 (O_606,N_9380,N_7286);
and UO_607 (O_607,N_9914,N_5084);
and UO_608 (O_608,N_7023,N_7086);
nand UO_609 (O_609,N_7942,N_6400);
nor UO_610 (O_610,N_7552,N_5802);
or UO_611 (O_611,N_9623,N_6456);
nand UO_612 (O_612,N_7239,N_5484);
nor UO_613 (O_613,N_7077,N_8546);
nand UO_614 (O_614,N_5396,N_7121);
or UO_615 (O_615,N_8915,N_8029);
or UO_616 (O_616,N_7066,N_8142);
or UO_617 (O_617,N_6983,N_9449);
or UO_618 (O_618,N_7218,N_8042);
or UO_619 (O_619,N_5738,N_5176);
nand UO_620 (O_620,N_9143,N_6169);
and UO_621 (O_621,N_9996,N_7384);
nand UO_622 (O_622,N_7824,N_5403);
and UO_623 (O_623,N_6865,N_6440);
and UO_624 (O_624,N_7975,N_9303);
nand UO_625 (O_625,N_7261,N_5047);
nand UO_626 (O_626,N_9934,N_8391);
nand UO_627 (O_627,N_6858,N_7764);
nor UO_628 (O_628,N_7733,N_5784);
or UO_629 (O_629,N_9172,N_6861);
nand UO_630 (O_630,N_5263,N_6556);
and UO_631 (O_631,N_7454,N_5973);
nand UO_632 (O_632,N_6488,N_6937);
or UO_633 (O_633,N_8180,N_5682);
and UO_634 (O_634,N_9228,N_9809);
or UO_635 (O_635,N_9491,N_7611);
nor UO_636 (O_636,N_8130,N_6056);
nand UO_637 (O_637,N_8196,N_7750);
or UO_638 (O_638,N_5600,N_9649);
nand UO_639 (O_639,N_5598,N_8896);
nor UO_640 (O_640,N_5859,N_6658);
and UO_641 (O_641,N_9375,N_9970);
nand UO_642 (O_642,N_9663,N_7669);
nand UO_643 (O_643,N_5911,N_8046);
and UO_644 (O_644,N_9942,N_8817);
and UO_645 (O_645,N_5636,N_5212);
or UO_646 (O_646,N_7338,N_7403);
nand UO_647 (O_647,N_7081,N_7374);
nor UO_648 (O_648,N_6923,N_7648);
or UO_649 (O_649,N_6070,N_7855);
or UO_650 (O_650,N_7367,N_8446);
and UO_651 (O_651,N_9610,N_6758);
or UO_652 (O_652,N_8659,N_8882);
nor UO_653 (O_653,N_6068,N_7787);
or UO_654 (O_654,N_6301,N_7270);
and UO_655 (O_655,N_7456,N_8138);
xnor UO_656 (O_656,N_5909,N_5556);
and UO_657 (O_657,N_6237,N_6071);
and UO_658 (O_658,N_5965,N_7201);
or UO_659 (O_659,N_6199,N_8145);
nand UO_660 (O_660,N_7358,N_5203);
and UO_661 (O_661,N_7277,N_8203);
and UO_662 (O_662,N_8892,N_7743);
or UO_663 (O_663,N_6528,N_5998);
nand UO_664 (O_664,N_9818,N_7396);
nand UO_665 (O_665,N_7436,N_5077);
or UO_666 (O_666,N_5284,N_8854);
nand UO_667 (O_667,N_8321,N_5445);
and UO_668 (O_668,N_6592,N_6509);
and UO_669 (O_669,N_8107,N_6476);
or UO_670 (O_670,N_5697,N_8916);
nor UO_671 (O_671,N_6809,N_8548);
and UO_672 (O_672,N_8039,N_6853);
nor UO_673 (O_673,N_5345,N_6877);
or UO_674 (O_674,N_6910,N_5522);
nor UO_675 (O_675,N_9314,N_5267);
nand UO_676 (O_676,N_5727,N_8396);
nand UO_677 (O_677,N_5679,N_7166);
nand UO_678 (O_678,N_7663,N_8258);
nor UO_679 (O_679,N_5996,N_8732);
or UO_680 (O_680,N_7401,N_8865);
or UO_681 (O_681,N_7507,N_8197);
nor UO_682 (O_682,N_9198,N_8412);
and UO_683 (O_683,N_5657,N_6552);
or UO_684 (O_684,N_6905,N_5504);
nor UO_685 (O_685,N_5615,N_5083);
and UO_686 (O_686,N_8780,N_6478);
and UO_687 (O_687,N_8418,N_6350);
and UO_688 (O_688,N_7898,N_9073);
and UO_689 (O_689,N_9589,N_8631);
nor UO_690 (O_690,N_8520,N_5312);
nand UO_691 (O_691,N_9207,N_7438);
and UO_692 (O_692,N_5661,N_5520);
nor UO_693 (O_693,N_5163,N_7622);
or UO_694 (O_694,N_8084,N_5398);
nand UO_695 (O_695,N_9736,N_5336);
or UO_696 (O_696,N_8705,N_6339);
nand UO_697 (O_697,N_9359,N_7060);
or UO_698 (O_698,N_6009,N_7985);
or UO_699 (O_699,N_7803,N_8954);
nor UO_700 (O_700,N_6513,N_5546);
or UO_701 (O_701,N_9713,N_9127);
nor UO_702 (O_702,N_6851,N_7505);
or UO_703 (O_703,N_5706,N_5116);
nor UO_704 (O_704,N_5940,N_6832);
and UO_705 (O_705,N_9560,N_9903);
or UO_706 (O_706,N_5441,N_7093);
or UO_707 (O_707,N_5530,N_7706);
or UO_708 (O_708,N_7096,N_8832);
and UO_709 (O_709,N_9133,N_8436);
nor UO_710 (O_710,N_7068,N_6659);
nor UO_711 (O_711,N_5213,N_8874);
or UO_712 (O_712,N_9605,N_7271);
and UO_713 (O_713,N_8380,N_5036);
and UO_714 (O_714,N_6055,N_6588);
or UO_715 (O_715,N_5282,N_8185);
and UO_716 (O_716,N_7084,N_7825);
and UO_717 (O_717,N_7229,N_6144);
and UO_718 (O_718,N_9490,N_5558);
or UO_719 (O_719,N_5572,N_8768);
nand UO_720 (O_720,N_5401,N_5624);
or UO_721 (O_721,N_8372,N_9142);
or UO_722 (O_722,N_8820,N_9795);
and UO_723 (O_723,N_9082,N_9185);
nand UO_724 (O_724,N_6299,N_5877);
or UO_725 (O_725,N_9092,N_5390);
nor UO_726 (O_726,N_8473,N_9741);
or UO_727 (O_727,N_8554,N_8776);
nor UO_728 (O_728,N_7686,N_7058);
and UO_729 (O_729,N_6227,N_7977);
xnor UO_730 (O_730,N_5496,N_5785);
and UO_731 (O_731,N_9299,N_7826);
nand UO_732 (O_732,N_9482,N_7966);
nor UO_733 (O_733,N_5560,N_9990);
and UO_734 (O_734,N_7015,N_5341);
nor UO_735 (O_735,N_7892,N_9954);
and UO_736 (O_736,N_6168,N_7847);
and UO_737 (O_737,N_7601,N_8300);
or UO_738 (O_738,N_7697,N_5356);
and UO_739 (O_739,N_8766,N_8584);
nand UO_740 (O_740,N_6480,N_8371);
nor UO_741 (O_741,N_7219,N_5112);
nor UO_742 (O_742,N_8756,N_6396);
nand UO_743 (O_743,N_5620,N_9044);
or UO_744 (O_744,N_9283,N_7473);
xor UO_745 (O_745,N_8078,N_8458);
and UO_746 (O_746,N_6083,N_5436);
or UO_747 (O_747,N_8352,N_5456);
nand UO_748 (O_748,N_9405,N_6819);
nand UO_749 (O_749,N_7639,N_6229);
nor UO_750 (O_750,N_7311,N_9746);
nand UO_751 (O_751,N_7492,N_8566);
or UO_752 (O_752,N_5113,N_6262);
and UO_753 (O_753,N_9645,N_5815);
and UO_754 (O_754,N_7210,N_8264);
and UO_755 (O_755,N_7924,N_9272);
nand UO_756 (O_756,N_7558,N_7313);
nor UO_757 (O_757,N_8044,N_5095);
nand UO_758 (O_758,N_6705,N_5731);
or UO_759 (O_759,N_8578,N_7628);
and UO_760 (O_760,N_9074,N_8337);
nor UO_761 (O_761,N_9100,N_5207);
nor UO_762 (O_762,N_9830,N_5547);
nand UO_763 (O_763,N_6021,N_9016);
nor UO_764 (O_764,N_9506,N_7889);
nor UO_765 (O_765,N_6190,N_7801);
and UO_766 (O_766,N_9584,N_6593);
or UO_767 (O_767,N_6157,N_9353);
nor UO_768 (O_768,N_9896,N_5248);
nand UO_769 (O_769,N_5509,N_9350);
or UO_770 (O_770,N_7696,N_5483);
nor UO_771 (O_771,N_7703,N_8858);
and UO_772 (O_772,N_9757,N_7918);
and UO_773 (O_773,N_9524,N_9015);
and UO_774 (O_774,N_7698,N_9689);
nand UO_775 (O_775,N_6107,N_9247);
nor UO_776 (O_776,N_7404,N_6892);
and UO_777 (O_777,N_5799,N_7186);
or UO_778 (O_778,N_5619,N_7431);
nand UO_779 (O_779,N_8753,N_7779);
nand UO_780 (O_780,N_8867,N_6814);
or UO_781 (O_781,N_9174,N_5592);
nor UO_782 (O_782,N_7802,N_6555);
and UO_783 (O_783,N_7485,N_6672);
nand UO_784 (O_784,N_7117,N_6822);
nor UO_785 (O_785,N_6176,N_9782);
nand UO_786 (O_786,N_6252,N_9053);
nor UO_787 (O_787,N_8500,N_8442);
and UO_788 (O_788,N_9395,N_7656);
nand UO_789 (O_789,N_7421,N_6541);
nor UO_790 (O_790,N_7619,N_9898);
nor UO_791 (O_791,N_6060,N_8819);
nand UO_792 (O_792,N_6072,N_8016);
nor UO_793 (O_793,N_7761,N_9087);
nand UO_794 (O_794,N_6137,N_7444);
nor UO_795 (O_795,N_8181,N_9527);
nand UO_796 (O_796,N_5002,N_7931);
nand UO_797 (O_797,N_9420,N_9650);
or UO_798 (O_798,N_5304,N_7617);
nor UO_799 (O_799,N_9362,N_9697);
nand UO_800 (O_800,N_7609,N_9739);
nand UO_801 (O_801,N_8244,N_6479);
nand UO_802 (O_802,N_6430,N_6432);
and UO_803 (O_803,N_5914,N_6738);
or UO_804 (O_804,N_8957,N_8610);
xnor UO_805 (O_805,N_5146,N_8827);
or UO_806 (O_806,N_8711,N_7948);
and UO_807 (O_807,N_7700,N_5407);
nor UO_808 (O_808,N_5960,N_9566);
nor UO_809 (O_809,N_9230,N_9197);
and UO_810 (O_810,N_5059,N_7883);
or UO_811 (O_811,N_7326,N_6591);
or UO_812 (O_812,N_5930,N_5219);
nor UO_813 (O_813,N_7441,N_8420);
or UO_814 (O_814,N_8148,N_6505);
nor UO_815 (O_815,N_5728,N_5292);
or UO_816 (O_816,N_6820,N_7502);
nand UO_817 (O_817,N_6264,N_9494);
nand UO_818 (O_818,N_8252,N_9578);
or UO_819 (O_819,N_9681,N_6295);
xor UO_820 (O_820,N_5725,N_9873);
nand UO_821 (O_821,N_8334,N_7151);
or UO_822 (O_822,N_7713,N_5359);
nand UO_823 (O_823,N_8561,N_9233);
or UO_824 (O_824,N_5849,N_9492);
nand UO_825 (O_825,N_8612,N_9936);
or UO_826 (O_826,N_7854,N_6870);
and UO_827 (O_827,N_9250,N_6603);
nand UO_828 (O_828,N_5313,N_9090);
and UO_829 (O_829,N_9770,N_9331);
and UO_830 (O_830,N_9273,N_8178);
nor UO_831 (O_831,N_7266,N_8105);
nand UO_832 (O_832,N_9001,N_5354);
or UO_833 (O_833,N_8818,N_5214);
or UO_834 (O_834,N_5734,N_8456);
nand UO_835 (O_835,N_9275,N_5486);
and UO_836 (O_836,N_6097,N_9203);
and UO_837 (O_837,N_7770,N_5952);
or UO_838 (O_838,N_6368,N_5653);
or UO_839 (O_839,N_7772,N_9824);
nor UO_840 (O_840,N_7449,N_6657);
nand UO_841 (O_841,N_5805,N_6712);
and UO_842 (O_842,N_5340,N_7100);
nor UO_843 (O_843,N_8856,N_6734);
nand UO_844 (O_844,N_8608,N_7153);
nor UO_845 (O_845,N_9562,N_8718);
and UO_846 (O_846,N_6753,N_5337);
and UO_847 (O_847,N_5514,N_6444);
nor UO_848 (O_848,N_6714,N_8080);
and UO_849 (O_849,N_6913,N_6108);
nor UO_850 (O_850,N_7225,N_9858);
and UO_851 (O_851,N_9549,N_8999);
nand UO_852 (O_852,N_7009,N_8757);
or UO_853 (O_853,N_8021,N_9065);
or UO_854 (O_854,N_7875,N_5510);
and UO_855 (O_855,N_8381,N_9412);
nor UO_856 (O_856,N_8033,N_5854);
or UO_857 (O_857,N_9979,N_6238);
or UO_858 (O_858,N_9007,N_9512);
and UO_859 (O_859,N_6399,N_8991);
nor UO_860 (O_860,N_6114,N_8905);
nand UO_861 (O_861,N_6879,N_8086);
xnor UO_862 (O_862,N_6726,N_7664);
nor UO_863 (O_863,N_6933,N_7083);
nor UO_864 (O_864,N_8447,N_7410);
nor UO_865 (O_865,N_8893,N_8063);
and UO_866 (O_866,N_6924,N_6367);
and UO_867 (O_867,N_8070,N_8785);
nand UO_868 (O_868,N_8636,N_9872);
or UO_869 (O_869,N_6888,N_9455);
or UO_870 (O_870,N_5878,N_7305);
nor UO_871 (O_871,N_8913,N_9166);
or UO_872 (O_872,N_9801,N_9952);
or UO_873 (O_873,N_7717,N_8149);
or UO_874 (O_874,N_7545,N_7468);
and UO_875 (O_875,N_7152,N_5416);
or UO_876 (O_876,N_8762,N_6660);
and UO_877 (O_877,N_9430,N_6255);
nand UO_878 (O_878,N_9399,N_7682);
and UO_879 (O_879,N_9093,N_9026);
nor UO_880 (O_880,N_5017,N_7379);
and UO_881 (O_881,N_9338,N_9788);
nand UO_882 (O_882,N_6766,N_9312);
or UO_883 (O_883,N_6481,N_5135);
and UO_884 (O_884,N_8299,N_6630);
nor UO_885 (O_885,N_6663,N_7291);
nand UO_886 (O_886,N_6124,N_8682);
and UO_887 (O_887,N_6364,N_5415);
and UO_888 (O_888,N_9980,N_7528);
or UO_889 (O_889,N_5901,N_9535);
and UO_890 (O_890,N_8678,N_9448);
or UO_891 (O_891,N_6461,N_6236);
and UO_892 (O_892,N_5428,N_8506);
nor UO_893 (O_893,N_7888,N_5708);
nand UO_894 (O_894,N_9702,N_6961);
and UO_895 (O_895,N_7477,N_6882);
or UO_896 (O_896,N_8279,N_6679);
nor UO_897 (O_897,N_5384,N_7044);
or UO_898 (O_898,N_7965,N_9466);
and UO_899 (O_899,N_9720,N_9307);
and UO_900 (O_900,N_6512,N_5581);
nor UO_901 (O_901,N_6698,N_5680);
nor UO_902 (O_902,N_9928,N_8601);
or UO_903 (O_903,N_5752,N_5872);
nor UO_904 (O_904,N_8490,N_9718);
nor UO_905 (O_905,N_8027,N_7296);
nand UO_906 (O_906,N_7727,N_6836);
or UO_907 (O_907,N_8193,N_7991);
and UO_908 (O_908,N_6895,N_7264);
and UO_909 (O_909,N_9480,N_6962);
nor UO_910 (O_910,N_9822,N_7643);
nor UO_911 (O_911,N_9116,N_6884);
nand UO_912 (O_912,N_8407,N_5066);
nand UO_913 (O_913,N_6161,N_8621);
and UO_914 (O_914,N_8170,N_6177);
or UO_915 (O_915,N_8980,N_6823);
and UO_916 (O_916,N_9938,N_6402);
nor UO_917 (O_917,N_9031,N_9600);
nand UO_918 (O_918,N_7668,N_8657);
and UO_919 (O_919,N_7868,N_7228);
nor UO_920 (O_920,N_6207,N_9426);
and UO_921 (O_921,N_8324,N_9551);
and UO_922 (O_922,N_7591,N_6840);
nor UO_923 (O_923,N_8634,N_8298);
nor UO_924 (O_924,N_6179,N_8164);
nor UO_925 (O_925,N_5944,N_9059);
nand UO_926 (O_926,N_7195,N_5524);
and UO_927 (O_927,N_6864,N_6151);
nand UO_928 (O_928,N_9269,N_6487);
nand UO_929 (O_929,N_9384,N_9393);
nor UO_930 (O_930,N_9863,N_6554);
nor UO_931 (O_931,N_9793,N_9192);
or UO_932 (O_932,N_7052,N_6428);
nor UO_933 (O_933,N_8483,N_6538);
nand UO_934 (O_934,N_7731,N_7548);
or UO_935 (O_935,N_8096,N_9315);
or UO_936 (O_936,N_8553,N_5876);
nand UO_937 (O_937,N_5529,N_6579);
nand UO_938 (O_938,N_8474,N_7476);
or UO_939 (O_939,N_8775,N_6903);
nand UO_940 (O_940,N_6527,N_8790);
and UO_941 (O_941,N_8460,N_7992);
nor UO_942 (O_942,N_9363,N_9365);
nor UO_943 (O_943,N_5140,N_6379);
nand UO_944 (O_944,N_5762,N_8222);
and UO_945 (O_945,N_7724,N_9501);
nor UO_946 (O_946,N_6272,N_8660);
nand UO_947 (O_947,N_9798,N_9725);
and UO_948 (O_948,N_5153,N_7136);
nand UO_949 (O_949,N_9637,N_9981);
or UO_950 (O_950,N_7496,N_6536);
or UO_951 (O_951,N_7489,N_9000);
nand UO_952 (O_952,N_6490,N_9387);
nand UO_953 (O_953,N_5990,N_7293);
or UO_954 (O_954,N_7484,N_8795);
and UO_955 (O_955,N_7150,N_5685);
and UO_956 (O_956,N_8770,N_7110);
or UO_957 (O_957,N_7448,N_9543);
nor UO_958 (O_958,N_7636,N_8162);
nor UO_959 (O_959,N_9604,N_7323);
or UO_960 (O_960,N_7289,N_6184);
nand UO_961 (O_961,N_5955,N_8529);
or UO_962 (O_962,N_6344,N_7788);
nor UO_963 (O_963,N_8786,N_7624);
or UO_964 (O_964,N_5918,N_8268);
and UO_965 (O_965,N_8791,N_9205);
nand UO_966 (O_966,N_8058,N_5052);
or UO_967 (O_967,N_8871,N_8340);
and UO_968 (O_968,N_7967,N_9413);
nor UO_969 (O_969,N_8238,N_9642);
and UO_970 (O_970,N_9890,N_9397);
nor UO_971 (O_971,N_7281,N_9727);
or UO_972 (O_972,N_5234,N_7159);
nor UO_973 (O_973,N_8012,N_7935);
nand UO_974 (O_974,N_6772,N_5349);
nor UO_975 (O_975,N_5127,N_5179);
and UO_976 (O_976,N_7168,N_6446);
and UO_977 (O_977,N_6008,N_5358);
or UO_978 (O_978,N_6044,N_6511);
nand UO_979 (O_979,N_8947,N_7380);
or UO_980 (O_980,N_6469,N_6717);
nor UO_981 (O_981,N_5430,N_9888);
nand UO_982 (O_982,N_8626,N_5791);
and UO_983 (O_983,N_5166,N_8803);
and UO_984 (O_984,N_7079,N_7214);
nor UO_985 (O_985,N_5929,N_6473);
and UO_986 (O_986,N_5933,N_7382);
nand UO_987 (O_987,N_8341,N_6906);
nor UO_988 (O_988,N_5222,N_9900);
nor UO_989 (O_989,N_7405,N_8214);
and UO_990 (O_990,N_7681,N_6403);
nor UO_991 (O_991,N_9669,N_7491);
or UO_992 (O_992,N_8901,N_6674);
and UO_993 (O_993,N_8642,N_8405);
or UO_994 (O_994,N_8377,N_9176);
and UO_995 (O_995,N_8453,N_9235);
nor UO_996 (O_996,N_8606,N_9875);
nand UO_997 (O_997,N_8686,N_5372);
and UO_998 (O_998,N_8126,N_8433);
nand UO_999 (O_999,N_9985,N_8026);
and UO_1000 (O_1000,N_5557,N_7549);
or UO_1001 (O_1001,N_7085,N_6833);
nand UO_1002 (O_1002,N_6562,N_9179);
nor UO_1003 (O_1003,N_5991,N_9920);
and UO_1004 (O_1004,N_9462,N_5884);
or UO_1005 (O_1005,N_6406,N_6287);
or UO_1006 (O_1006,N_8137,N_9921);
nand UO_1007 (O_1007,N_5231,N_7495);
nand UO_1008 (O_1008,N_6686,N_5864);
or UO_1009 (O_1009,N_9304,N_8179);
nor UO_1010 (O_1010,N_9827,N_9334);
or UO_1011 (O_1011,N_5925,N_7811);
and UO_1012 (O_1012,N_8994,N_8125);
or UO_1013 (O_1013,N_9958,N_8034);
nand UO_1014 (O_1014,N_8051,N_5369);
and UO_1015 (O_1015,N_8245,N_9853);
xor UO_1016 (O_1016,N_9842,N_5289);
or UO_1017 (O_1017,N_8835,N_5326);
or UO_1018 (O_1018,N_6265,N_5984);
and UO_1019 (O_1019,N_8496,N_9469);
and UO_1020 (O_1020,N_7303,N_5185);
nand UO_1021 (O_1021,N_6449,N_9868);
or UO_1022 (O_1022,N_7223,N_7927);
nor UO_1023 (O_1023,N_7784,N_6666);
nand UO_1024 (O_1024,N_8043,N_6532);
nor UO_1025 (O_1025,N_6333,N_9941);
or UO_1026 (O_1026,N_7532,N_6434);
nor UO_1027 (O_1027,N_7197,N_7465);
nor UO_1028 (O_1028,N_5076,N_5698);
and UO_1029 (O_1029,N_9182,N_6800);
and UO_1030 (O_1030,N_9812,N_5830);
nor UO_1031 (O_1031,N_8176,N_9927);
and UO_1032 (O_1032,N_8643,N_7728);
and UO_1033 (O_1033,N_6437,N_7752);
nand UO_1034 (O_1034,N_9369,N_9238);
nor UO_1035 (O_1035,N_9783,N_8485);
nor UO_1036 (O_1036,N_8556,N_6149);
nand UO_1037 (O_1037,N_9162,N_6742);
nand UO_1038 (O_1038,N_9550,N_9748);
nand UO_1039 (O_1039,N_6982,N_6967);
nand UO_1040 (O_1040,N_7213,N_5670);
or UO_1041 (O_1041,N_5915,N_5666);
nor UO_1042 (O_1042,N_9493,N_6062);
nand UO_1043 (O_1043,N_9901,N_6533);
nor UO_1044 (O_1044,N_6852,N_7869);
nor UO_1045 (O_1045,N_7719,N_8752);
or UO_1046 (O_1046,N_6335,N_7789);
or UO_1047 (O_1047,N_7504,N_9814);
and UO_1048 (O_1048,N_7670,N_5237);
nor UO_1049 (O_1049,N_6812,N_8379);
nand UO_1050 (O_1050,N_7329,N_5610);
nor UO_1051 (O_1051,N_6073,N_6348);
and UO_1052 (O_1052,N_8205,N_9019);
or UO_1053 (O_1053,N_9276,N_6415);
or UO_1054 (O_1054,N_9056,N_5921);
or UO_1055 (O_1055,N_8429,N_9302);
nor UO_1056 (O_1056,N_5129,N_6150);
or UO_1057 (O_1057,N_8995,N_8622);
nand UO_1058 (O_1058,N_6751,N_6454);
or UO_1059 (O_1059,N_8704,N_9126);
nand UO_1060 (O_1060,N_9504,N_9388);
and UO_1061 (O_1061,N_8736,N_7351);
or UO_1062 (O_1062,N_7659,N_9950);
or UO_1063 (O_1063,N_5080,N_5780);
nand UO_1064 (O_1064,N_7224,N_6492);
or UO_1065 (O_1065,N_9436,N_7865);
nor UO_1066 (O_1066,N_6727,N_5018);
nor UO_1067 (O_1067,N_5649,N_9564);
nand UO_1068 (O_1068,N_8849,N_6385);
and UO_1069 (O_1069,N_5582,N_7256);
nor UO_1070 (O_1070,N_8884,N_6645);
and UO_1071 (O_1071,N_5270,N_6431);
nor UO_1072 (O_1072,N_6930,N_5577);
or UO_1073 (O_1073,N_5352,N_9216);
nor UO_1074 (O_1074,N_8120,N_5739);
or UO_1075 (O_1075,N_8524,N_8917);
nand UO_1076 (O_1076,N_7806,N_6259);
or UO_1077 (O_1077,N_5733,N_6205);
or UO_1078 (O_1078,N_6943,N_8154);
and UO_1079 (O_1079,N_8542,N_6835);
nand UO_1080 (O_1080,N_5498,N_5442);
or UO_1081 (O_1081,N_9119,N_6130);
and UO_1082 (O_1082,N_5660,N_8006);
and UO_1083 (O_1083,N_6881,N_5244);
or UO_1084 (O_1084,N_5761,N_7929);
or UO_1085 (O_1085,N_6376,N_5964);
nand UO_1086 (O_1086,N_5051,N_5898);
nor UO_1087 (O_1087,N_9820,N_9665);
or UO_1088 (O_1088,N_8669,N_6110);
and UO_1089 (O_1089,N_6363,N_9062);
and UO_1090 (O_1090,N_9644,N_6496);
nand UO_1091 (O_1091,N_8788,N_5635);
or UO_1092 (O_1092,N_9676,N_7560);
or UO_1093 (O_1093,N_9688,N_9485);
nor UO_1094 (O_1094,N_5995,N_6049);
and UO_1095 (O_1095,N_5273,N_5432);
and UO_1096 (O_1096,N_5621,N_9255);
and UO_1097 (O_1097,N_6788,N_8675);
nor UO_1098 (O_1098,N_6318,N_5117);
nand UO_1099 (O_1099,N_9955,N_8544);
and UO_1100 (O_1100,N_5078,N_6059);
nor UO_1101 (O_1101,N_7976,N_9429);
nand UO_1102 (O_1102,N_5086,N_7361);
or UO_1103 (O_1103,N_7739,N_5726);
or UO_1104 (O_1104,N_9045,N_7781);
nor UO_1105 (O_1105,N_9613,N_9667);
nor UO_1106 (O_1106,N_5424,N_8890);
nand UO_1107 (O_1107,N_9157,N_6544);
nand UO_1108 (O_1108,N_6332,N_8357);
nor UO_1109 (O_1109,N_8260,N_7963);
nand UO_1110 (O_1110,N_8851,N_6710);
nor UO_1111 (O_1111,N_7867,N_9862);
or UO_1112 (O_1112,N_5703,N_5523);
nor UO_1113 (O_1113,N_7173,N_8591);
or UO_1114 (O_1114,N_6954,N_6497);
nor UO_1115 (O_1115,N_8293,N_9169);
nor UO_1116 (O_1116,N_6855,N_6115);
nor UO_1117 (O_1117,N_5629,N_6453);
and UO_1118 (O_1118,N_6136,N_5923);
nand UO_1119 (O_1119,N_5763,N_9851);
nand UO_1120 (O_1120,N_5691,N_8302);
and UO_1121 (O_1121,N_9882,N_8237);
nand UO_1122 (O_1122,N_9394,N_7065);
nor UO_1123 (O_1123,N_8290,N_6051);
xor UO_1124 (O_1124,N_9486,N_6450);
or UO_1125 (O_1125,N_6003,N_5953);
and UO_1126 (O_1126,N_5943,N_9088);
nand UO_1127 (O_1127,N_6694,N_8011);
or UO_1128 (O_1128,N_9104,N_6856);
or UO_1129 (O_1129,N_8697,N_9123);
or UO_1130 (O_1130,N_8236,N_9879);
and UO_1131 (O_1131,N_8635,N_5924);
and UO_1132 (O_1132,N_7688,N_6740);
nor UO_1133 (O_1133,N_6174,N_5073);
nor UO_1134 (O_1134,N_9831,N_5181);
nor UO_1135 (O_1135,N_6201,N_7720);
xor UO_1136 (O_1136,N_9986,N_8904);
or UO_1137 (O_1137,N_6897,N_9641);
and UO_1138 (O_1138,N_8374,N_5531);
and UO_1139 (O_1139,N_8365,N_5389);
and UO_1140 (O_1140,N_7903,N_7260);
nor UO_1141 (O_1141,N_8846,N_9378);
or UO_1142 (O_1142,N_9025,N_8443);
nor UO_1143 (O_1143,N_9993,N_8388);
and UO_1144 (O_1144,N_7041,N_9510);
or UO_1145 (O_1145,N_7823,N_6243);
nor UO_1146 (O_1146,N_7300,N_8209);
nand UO_1147 (O_1147,N_5931,N_7641);
and UO_1148 (O_1148,N_6340,N_7259);
or UO_1149 (O_1149,N_6643,N_7094);
and UO_1150 (O_1150,N_8755,N_9997);
nand UO_1151 (O_1151,N_6366,N_9336);
nand UO_1152 (O_1152,N_6941,N_7675);
nor UO_1153 (O_1153,N_6618,N_6621);
or UO_1154 (O_1154,N_7199,N_5590);
nor UO_1155 (O_1155,N_8061,N_9481);
nor UO_1156 (O_1156,N_6076,N_8592);
nor UO_1157 (O_1157,N_7782,N_7457);
or UO_1158 (O_1158,N_5096,N_8821);
nor UO_1159 (O_1159,N_7268,N_9291);
nand UO_1160 (O_1160,N_7705,N_6994);
nor UO_1161 (O_1161,N_5507,N_7751);
and UO_1162 (O_1162,N_9498,N_5225);
nor UO_1163 (O_1163,N_9554,N_5525);
nand UO_1164 (O_1164,N_9762,N_6080);
nand UO_1165 (O_1165,N_5928,N_5093);
and UO_1166 (O_1166,N_5434,N_5957);
or UO_1167 (O_1167,N_8650,N_7593);
and UO_1168 (O_1168,N_9694,N_6871);
nor UO_1169 (O_1169,N_8714,N_8644);
or UO_1170 (O_1170,N_6568,N_6273);
or UO_1171 (O_1171,N_8625,N_9525);
nand UO_1172 (O_1172,N_9035,N_6769);
nand UO_1173 (O_1173,N_6421,N_8552);
or UO_1174 (O_1174,N_6687,N_5269);
or UO_1175 (O_1175,N_8256,N_8213);
or UO_1176 (O_1176,N_6408,N_9587);
and UO_1177 (O_1177,N_6500,N_9424);
or UO_1178 (O_1178,N_5469,N_8320);
or UO_1179 (O_1179,N_5797,N_5792);
and UO_1180 (O_1180,N_9124,N_5894);
or UO_1181 (O_1181,N_6642,N_7606);
nor UO_1182 (O_1182,N_7704,N_8523);
or UO_1183 (O_1183,N_7008,N_7881);
nand UO_1184 (O_1184,N_6091,N_6191);
and UO_1185 (O_1185,N_8455,N_7377);
nand UO_1186 (O_1186,N_8304,N_5331);
nor UO_1187 (O_1187,N_6047,N_9003);
and UO_1188 (O_1188,N_7004,N_9502);
nand UO_1189 (O_1189,N_7304,N_8719);
nand UO_1190 (O_1190,N_8645,N_8616);
nor UO_1191 (O_1191,N_7603,N_5567);
nand UO_1192 (O_1192,N_5721,N_9840);
nor UO_1193 (O_1193,N_9254,N_8132);
or UO_1194 (O_1194,N_5503,N_6756);
nor UO_1195 (O_1195,N_8872,N_8280);
nand UO_1196 (O_1196,N_7645,N_7184);
and UO_1197 (O_1197,N_5970,N_6652);
nor UO_1198 (O_1198,N_5757,N_6540);
or UO_1199 (O_1199,N_6880,N_5494);
nor UO_1200 (O_1200,N_6946,N_7172);
and UO_1201 (O_1201,N_7928,N_9464);
nand UO_1202 (O_1202,N_6977,N_6885);
or UO_1203 (O_1203,N_9131,N_5157);
or UO_1204 (O_1204,N_8665,N_5388);
or UO_1205 (O_1205,N_8507,N_8565);
and UO_1206 (O_1206,N_5873,N_7028);
or UO_1207 (O_1207,N_7555,N_6866);
nor UO_1208 (O_1208,N_7206,N_5056);
nor UO_1209 (O_1209,N_8328,N_8927);
or UO_1210 (O_1210,N_9161,N_9442);
and UO_1211 (O_1211,N_5765,N_8912);
or UO_1212 (O_1212,N_9759,N_6253);
nor UO_1213 (O_1213,N_9675,N_8247);
nor UO_1214 (O_1214,N_6004,N_9036);
and UO_1215 (O_1215,N_5798,N_8919);
nor UO_1216 (O_1216,N_5133,N_6602);
or UO_1217 (O_1217,N_9776,N_5809);
nand UO_1218 (O_1218,N_9222,N_7371);
nand UO_1219 (O_1219,N_9415,N_5001);
nand UO_1220 (O_1220,N_7279,N_6371);
nand UO_1221 (O_1221,N_5701,N_7422);
nor UO_1222 (O_1222,N_5717,N_8049);
nor UO_1223 (O_1223,N_8930,N_7997);
nor UO_1224 (O_1224,N_6566,N_6120);
and UO_1225 (O_1225,N_9766,N_7799);
nor UO_1226 (O_1226,N_8853,N_6706);
nand UO_1227 (O_1227,N_6971,N_9971);
or UO_1228 (O_1228,N_6123,N_9919);
or UO_1229 (O_1229,N_6018,N_7247);
nor UO_1230 (O_1230,N_5444,N_7785);
nand UO_1231 (O_1231,N_7915,N_8572);
and UO_1232 (O_1232,N_6001,N_9843);
nor UO_1233 (O_1233,N_5150,N_5848);
nand UO_1234 (O_1234,N_8475,N_6773);
nor UO_1235 (O_1235,N_7397,N_6631);
and UO_1236 (O_1236,N_7828,N_5491);
or UO_1237 (O_1237,N_5142,N_5663);
nand UO_1238 (O_1238,N_8373,N_6329);
and UO_1239 (O_1239,N_6098,N_6413);
or UO_1240 (O_1240,N_7314,N_9624);
and UO_1241 (O_1241,N_5242,N_9909);
nor UO_1242 (O_1242,N_5732,N_9634);
and UO_1243 (O_1243,N_7767,N_8157);
and UO_1244 (O_1244,N_6278,N_9075);
and UO_1245 (O_1245,N_7583,N_9912);
nor UO_1246 (O_1246,N_9755,N_8408);
or UO_1247 (O_1247,N_6890,N_7131);
nand UO_1248 (O_1248,N_8759,N_5431);
nand UO_1249 (O_1249,N_5843,N_8467);
or UO_1250 (O_1250,N_5478,N_6291);
and UO_1251 (O_1251,N_7032,N_5667);
nor UO_1252 (O_1252,N_8249,N_6337);
and UO_1253 (O_1253,N_9439,N_5460);
nand UO_1254 (O_1254,N_8615,N_8873);
nor UO_1255 (O_1255,N_5199,N_5348);
nor UO_1256 (O_1256,N_9700,N_5737);
nand UO_1257 (O_1257,N_8773,N_8679);
nor UO_1258 (O_1258,N_6308,N_5788);
nand UO_1259 (O_1259,N_5647,N_7148);
or UO_1260 (O_1260,N_8017,N_5216);
or UO_1261 (O_1261,N_6867,N_7853);
nor UO_1262 (O_1262,N_9547,N_6111);
nor UO_1263 (O_1263,N_9229,N_5608);
nor UO_1264 (O_1264,N_5704,N_7217);
and UO_1265 (O_1265,N_9252,N_5315);
nor UO_1266 (O_1266,N_5110,N_8868);
nor UO_1267 (O_1267,N_9390,N_5934);
and UO_1268 (O_1268,N_8097,N_6200);
and UO_1269 (O_1269,N_9358,N_8401);
and UO_1270 (O_1270,N_5155,N_7817);
or UO_1271 (O_1271,N_7105,N_5841);
nor UO_1272 (O_1272,N_5124,N_5605);
nand UO_1273 (O_1273,N_6127,N_9768);
and UO_1274 (O_1274,N_9327,N_7943);
nor UO_1275 (O_1275,N_6976,N_6745);
or UO_1276 (O_1276,N_6670,N_6516);
and UO_1277 (O_1277,N_7385,N_6285);
and UO_1278 (O_1278,N_5857,N_9925);
nand UO_1279 (O_1279,N_9998,N_9433);
nand UO_1280 (O_1280,N_6902,N_5042);
nor UO_1281 (O_1281,N_6637,N_7769);
nand UO_1282 (O_1282,N_6845,N_8472);
or UO_1283 (O_1283,N_6391,N_5922);
nand UO_1284 (O_1284,N_7317,N_5409);
and UO_1285 (O_1285,N_5926,N_5342);
nor UO_1286 (O_1286,N_8509,N_6172);
or UO_1287 (O_1287,N_9568,N_6617);
nor UO_1288 (O_1288,N_5364,N_9404);
nand UO_1289 (O_1289,N_8174,N_9244);
nor UO_1290 (O_1290,N_5551,N_9777);
and UO_1291 (O_1291,N_8653,N_7926);
or UO_1292 (O_1292,N_6206,N_9330);
and UO_1293 (O_1293,N_6494,N_8847);
nand UO_1294 (O_1294,N_5298,N_9039);
nand UO_1295 (O_1295,N_7226,N_7525);
and UO_1296 (O_1296,N_8772,N_5963);
or UO_1297 (O_1297,N_5450,N_8582);
nor UO_1298 (O_1298,N_6771,N_7027);
nand UO_1299 (O_1299,N_8720,N_8850);
or UO_1300 (O_1300,N_9922,N_8156);
nand UO_1301 (O_1301,N_8898,N_6017);
or UO_1302 (O_1302,N_8727,N_9346);
and UO_1303 (O_1303,N_9144,N_6485);
and UO_1304 (O_1304,N_9438,N_7846);
nor UO_1305 (O_1305,N_6996,N_5371);
or UO_1306 (O_1306,N_8754,N_5867);
nand UO_1307 (O_1307,N_7797,N_9751);
nand UO_1308 (O_1308,N_6785,N_8666);
or UO_1309 (O_1309,N_5221,N_7075);
or UO_1310 (O_1310,N_5515,N_7763);
nor UO_1311 (O_1311,N_9165,N_8282);
or UO_1312 (O_1312,N_7561,N_7158);
nand UO_1313 (O_1313,N_5031,N_9321);
or UO_1314 (O_1314,N_7143,N_6372);
nand UO_1315 (O_1315,N_8926,N_7212);
nand UO_1316 (O_1316,N_9627,N_5749);
and UO_1317 (O_1317,N_8274,N_8640);
or UO_1318 (O_1318,N_9094,N_8580);
nor UO_1319 (O_1319,N_7642,N_5540);
xor UO_1320 (O_1320,N_5215,N_9808);
or UO_1321 (O_1321,N_6289,N_8859);
nand UO_1322 (O_1322,N_6390,N_8397);
or UO_1323 (O_1323,N_7588,N_8721);
and UO_1324 (O_1324,N_9051,N_7088);
or UO_1325 (O_1325,N_7844,N_7416);
nand UO_1326 (O_1326,N_7805,N_9992);
or UO_1327 (O_1327,N_8333,N_8688);
or UO_1328 (O_1328,N_6844,N_6662);
or UO_1329 (O_1329,N_5180,N_6358);
and UO_1330 (O_1330,N_9660,N_9008);
nand UO_1331 (O_1331,N_7461,N_5465);
and UO_1332 (O_1332,N_6502,N_8318);
nor UO_1333 (O_1333,N_5564,N_9474);
nand UO_1334 (O_1334,N_6316,N_8816);
or UO_1335 (O_1335,N_7039,N_9772);
and UO_1336 (O_1336,N_9461,N_8782);
nand UO_1337 (O_1337,N_5736,N_5544);
and UO_1338 (O_1338,N_9773,N_7563);
and UO_1339 (O_1339,N_8681,N_8876);
nor UO_1340 (O_1340,N_7426,N_9447);
nor UO_1341 (O_1341,N_6798,N_9709);
nand UO_1342 (O_1342,N_7996,N_7295);
and UO_1343 (O_1343,N_5011,N_8102);
nand UO_1344 (O_1344,N_6632,N_5361);
nor UO_1345 (O_1345,N_7983,N_9111);
and UO_1346 (O_1346,N_6711,N_5642);
and UO_1347 (O_1347,N_8344,N_6953);
nor UO_1348 (O_1348,N_9014,N_5638);
nor UO_1349 (O_1349,N_5641,N_7718);
and UO_1350 (O_1350,N_6574,N_8074);
or UO_1351 (O_1351,N_5101,N_7506);
and UO_1352 (O_1352,N_8813,N_5986);
and UO_1353 (O_1353,N_5906,N_5681);
and UO_1354 (O_1354,N_9373,N_5882);
nor UO_1355 (O_1355,N_9110,N_9076);
nor UO_1356 (O_1356,N_6292,N_6989);
and UO_1357 (O_1357,N_5472,N_6565);
and UO_1358 (O_1358,N_6302,N_7427);
or UO_1359 (O_1359,N_7912,N_7878);
nor UO_1360 (O_1360,N_5324,N_6254);
or UO_1361 (O_1361,N_5578,N_9301);
nor UO_1362 (O_1362,N_8224,N_5183);
and UO_1363 (O_1363,N_5565,N_6197);
or UO_1364 (O_1364,N_6577,N_6899);
and UO_1365 (O_1365,N_7237,N_5082);
nor UO_1366 (O_1366,N_6900,N_6393);
nand UO_1367 (O_1367,N_9356,N_5363);
nand UO_1368 (O_1368,N_9744,N_5206);
and UO_1369 (O_1369,N_9792,N_8315);
or UO_1370 (O_1370,N_6928,N_9984);
and UO_1371 (O_1371,N_9190,N_6969);
nand UO_1372 (O_1372,N_6669,N_9876);
and UO_1373 (O_1373,N_5323,N_9573);
xnor UO_1374 (O_1374,N_5090,N_7146);
nand UO_1375 (O_1375,N_7979,N_8362);
nor UO_1376 (O_1376,N_6389,N_5255);
nand UO_1377 (O_1377,N_6279,N_7666);
or UO_1378 (O_1378,N_5672,N_7458);
nand UO_1379 (O_1379,N_7472,N_9889);
and UO_1380 (O_1380,N_7961,N_8574);
nor UO_1381 (O_1381,N_8587,N_9940);
nand UO_1382 (O_1382,N_8624,N_9574);
and UO_1383 (O_1383,N_8864,N_9671);
and UO_1384 (O_1384,N_5845,N_6780);
nor UO_1385 (O_1385,N_7091,N_7318);
or UO_1386 (O_1386,N_7535,N_7970);
nor UO_1387 (O_1387,N_7650,N_9680);
and UO_1388 (O_1388,N_5353,N_8970);
nor UO_1389 (O_1389,N_9298,N_8652);
and UO_1390 (O_1390,N_7501,N_8731);
or UO_1391 (O_1391,N_6654,N_6521);
and UO_1392 (O_1392,N_5188,N_6334);
nor UO_1393 (O_1393,N_7090,N_6404);
and UO_1394 (O_1394,N_5912,N_6995);
or UO_1395 (O_1395,N_6691,N_6515);
and UO_1396 (O_1396,N_8522,N_8147);
nor UO_1397 (O_1397,N_5240,N_6922);
nand UO_1398 (O_1398,N_8527,N_8583);
or UO_1399 (O_1399,N_6623,N_7463);
or UO_1400 (O_1400,N_5853,N_8122);
nor UO_1401 (O_1401,N_5808,N_8764);
nor UO_1402 (O_1402,N_9355,N_8935);
and UO_1403 (O_1403,N_5744,N_7202);
nand UO_1404 (O_1404,N_8614,N_5067);
nor UO_1405 (O_1405,N_6296,N_6041);
and UO_1406 (O_1406,N_8655,N_8330);
or UO_1407 (O_1407,N_5058,N_8993);
nor UO_1408 (O_1408,N_5137,N_9983);
and UO_1409 (O_1409,N_5280,N_7036);
nor UO_1410 (O_1410,N_9565,N_8228);
nand UO_1411 (O_1411,N_5393,N_9332);
or UO_1412 (O_1412,N_9780,N_7292);
or UO_1413 (O_1413,N_6225,N_7283);
or UO_1414 (O_1414,N_9964,N_8263);
and UO_1415 (O_1415,N_7180,N_8009);
nor UO_1416 (O_1416,N_7773,N_9516);
and UO_1417 (O_1417,N_9224,N_8018);
nor UO_1418 (O_1418,N_7134,N_9895);
or UO_1419 (O_1419,N_7524,N_6170);
and UO_1420 (O_1420,N_8696,N_5061);
and UO_1421 (O_1421,N_6932,N_5686);
nor UO_1422 (O_1422,N_6980,N_6920);
or UO_1423 (O_1423,N_8877,N_6022);
nand UO_1424 (O_1424,N_9150,N_9038);
and UO_1425 (O_1425,N_6290,N_8953);
nor UO_1426 (O_1426,N_5254,N_9154);
or UO_1427 (O_1427,N_7033,N_9839);
and UO_1428 (O_1428,N_7120,N_9478);
and UO_1429 (O_1429,N_8478,N_9043);
nor UO_1430 (O_1430,N_7040,N_8577);
and UO_1431 (O_1431,N_5005,N_6525);
nor UO_1432 (O_1432,N_8569,N_6891);
and UO_1433 (O_1433,N_7701,N_5724);
or UO_1434 (O_1434,N_8741,N_7521);
nand UO_1435 (O_1435,N_6837,N_5412);
nand UO_1436 (O_1436,N_6729,N_7022);
or UO_1437 (O_1437,N_8792,N_5458);
nand UO_1438 (O_1438,N_8003,N_7316);
nand UO_1439 (O_1439,N_6013,N_6026);
nor UO_1440 (O_1440,N_6493,N_8430);
nor UO_1441 (O_1441,N_7275,N_7109);
nor UO_1442 (O_1442,N_6102,N_9618);
nor UO_1443 (O_1443,N_6104,N_9427);
nand UO_1444 (O_1444,N_7451,N_7145);
and UO_1445 (O_1445,N_7062,N_5893);
nor UO_1446 (O_1446,N_5296,N_7845);
or UO_1447 (O_1447,N_7530,N_6158);
or UO_1448 (O_1448,N_8794,N_8060);
nand UO_1449 (O_1449,N_8589,N_6094);
or UO_1450 (O_1450,N_8946,N_7800);
or UO_1451 (O_1451,N_5007,N_5603);
nor UO_1452 (O_1452,N_6678,N_7978);
or UO_1453 (O_1453,N_9239,N_9248);
or UO_1454 (O_1454,N_5671,N_9616);
and UO_1455 (O_1455,N_9946,N_9630);
or UO_1456 (O_1456,N_9561,N_7343);
and UO_1457 (O_1457,N_5039,N_9292);
nand UO_1458 (O_1458,N_5351,N_8054);
nand UO_1459 (O_1459,N_7512,N_5413);
nand UO_1460 (O_1460,N_6038,N_8114);
nand UO_1461 (O_1461,N_6315,N_5689);
nor UO_1462 (O_1462,N_8235,N_5278);
nor UO_1463 (O_1463,N_5769,N_7526);
nor UO_1464 (O_1464,N_6234,N_9326);
or UO_1465 (O_1465,N_6211,N_5054);
or UO_1466 (O_1466,N_5198,N_5102);
or UO_1467 (O_1467,N_9191,N_7014);
and UO_1468 (O_1468,N_8571,N_6965);
and UO_1469 (O_1469,N_6696,N_7020);
and UO_1470 (O_1470,N_6181,N_8958);
and UO_1471 (O_1471,N_5740,N_8914);
nand UO_1472 (O_1472,N_8677,N_8128);
nor UO_1473 (O_1473,N_9422,N_7246);
nor UO_1474 (O_1474,N_8155,N_9837);
or UO_1475 (O_1475,N_7741,N_9022);
or UO_1476 (O_1476,N_7299,N_8974);
and UO_1477 (O_1477,N_8806,N_8715);
and UO_1478 (O_1478,N_8382,N_5041);
nor UO_1479 (O_1479,N_6935,N_7336);
or UO_1480 (O_1480,N_7620,N_7527);
or UO_1481 (O_1481,N_5260,N_6635);
nor UO_1482 (O_1482,N_5634,N_5344);
and UO_1483 (O_1483,N_8568,N_9883);
nand UO_1484 (O_1484,N_7076,N_9402);
or UO_1485 (O_1485,N_5420,N_6826);
nor UO_1486 (O_1486,N_5863,N_5370);
or UO_1487 (O_1487,N_5655,N_5217);
nor UO_1488 (O_1488,N_7679,N_5889);
nor UO_1489 (O_1489,N_5196,N_5012);
or UO_1490 (O_1490,N_8242,N_6801);
and UO_1491 (O_1491,N_9854,N_6615);
nand UO_1492 (O_1492,N_5108,N_5550);
nand UO_1493 (O_1493,N_9581,N_9611);
nand UO_1494 (O_1494,N_6321,N_9134);
nor UO_1495 (O_1495,N_9937,N_9345);
nand UO_1496 (O_1496,N_9452,N_5302);
nand UO_1497 (O_1497,N_6721,N_9408);
xnor UO_1498 (O_1498,N_9083,N_7757);
or UO_1499 (O_1499,N_7597,N_8860);
endmodule