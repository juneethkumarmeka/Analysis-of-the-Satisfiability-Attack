module basic_1500_15000_2000_60_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_139,In_16);
and U1 (N_1,In_731,In_187);
xor U2 (N_2,In_1179,In_640);
and U3 (N_3,In_760,In_1092);
nor U4 (N_4,In_615,In_251);
or U5 (N_5,In_1242,In_856);
nor U6 (N_6,In_517,In_709);
or U7 (N_7,In_582,In_652);
or U8 (N_8,In_446,In_372);
or U9 (N_9,In_911,In_1352);
nand U10 (N_10,In_577,In_510);
and U11 (N_11,In_110,In_889);
or U12 (N_12,In_899,In_1151);
or U13 (N_13,In_272,In_280);
nor U14 (N_14,In_89,In_1026);
or U15 (N_15,In_204,In_1012);
xnor U16 (N_16,In_815,In_1375);
nand U17 (N_17,In_1146,In_1195);
xor U18 (N_18,In_299,In_1013);
nand U19 (N_19,In_1088,In_1311);
nor U20 (N_20,In_1389,In_365);
xor U21 (N_21,In_1203,In_823);
nor U22 (N_22,In_1212,In_1287);
or U23 (N_23,In_779,In_613);
or U24 (N_24,In_407,In_1142);
nor U25 (N_25,In_560,In_1492);
or U26 (N_26,In_1010,In_216);
nand U27 (N_27,In_151,In_1218);
nand U28 (N_28,In_1217,In_245);
and U29 (N_29,In_527,In_818);
nor U30 (N_30,In_881,In_33);
xnor U31 (N_31,In_1374,In_1402);
xor U32 (N_32,In_434,In_1450);
and U33 (N_33,In_898,In_226);
or U34 (N_34,In_489,In_1284);
or U35 (N_35,In_524,In_79);
and U36 (N_36,In_437,In_798);
xnor U37 (N_37,In_822,In_684);
or U38 (N_38,In_782,In_598);
xor U39 (N_39,In_706,In_1249);
nor U40 (N_40,In_237,In_669);
nor U41 (N_41,In_1124,In_1063);
nor U42 (N_42,In_1486,In_1274);
and U43 (N_43,In_637,In_1465);
or U44 (N_44,In_411,In_330);
nor U45 (N_45,In_1476,In_970);
or U46 (N_46,In_21,In_1087);
and U47 (N_47,In_1388,In_890);
xor U48 (N_48,In_631,In_750);
or U49 (N_49,In_174,In_937);
nor U50 (N_50,In_1317,In_693);
or U51 (N_51,In_364,In_182);
and U52 (N_52,In_633,In_1250);
nor U53 (N_53,In_695,In_550);
and U54 (N_54,In_1137,In_676);
or U55 (N_55,In_113,In_1008);
and U56 (N_56,In_250,In_513);
nor U57 (N_57,In_1040,In_925);
xor U58 (N_58,In_374,In_1048);
xor U59 (N_59,In_328,In_1477);
xor U60 (N_60,In_66,In_1094);
or U61 (N_61,In_109,In_773);
nor U62 (N_62,In_1366,In_474);
nor U63 (N_63,In_367,In_260);
nand U64 (N_64,In_192,In_303);
xor U65 (N_65,In_1115,In_843);
or U66 (N_66,In_155,In_1347);
xnor U67 (N_67,In_100,In_1213);
nor U68 (N_68,In_741,In_1164);
nor U69 (N_69,In_453,In_841);
and U70 (N_70,In_1310,In_1441);
and U71 (N_71,In_1020,In_740);
nor U72 (N_72,In_1334,In_757);
nor U73 (N_73,In_968,In_1403);
or U74 (N_74,In_1415,In_229);
nand U75 (N_75,In_569,In_1257);
xnor U76 (N_76,In_479,In_356);
nor U77 (N_77,In_339,In_632);
and U78 (N_78,In_327,In_785);
and U79 (N_79,In_72,In_78);
nor U80 (N_80,In_404,In_654);
xor U81 (N_81,In_289,In_467);
nor U82 (N_82,In_1315,In_964);
or U83 (N_83,In_344,In_468);
and U84 (N_84,In_1245,In_1396);
or U85 (N_85,In_564,In_1207);
nand U86 (N_86,In_459,In_101);
or U87 (N_87,In_991,In_77);
and U88 (N_88,In_730,In_247);
nand U89 (N_89,In_1130,In_973);
xnor U90 (N_90,In_412,In_959);
xor U91 (N_91,In_179,In_470);
nand U92 (N_92,In_724,In_213);
or U93 (N_93,In_267,In_1439);
nand U94 (N_94,In_1078,In_1320);
xor U95 (N_95,In_1271,In_961);
nand U96 (N_96,In_111,In_1225);
or U97 (N_97,In_1099,In_1417);
nand U98 (N_98,In_138,In_1073);
xnor U99 (N_99,In_645,In_162);
or U100 (N_100,In_166,In_274);
or U101 (N_101,In_482,In_848);
and U102 (N_102,In_1062,In_142);
or U103 (N_103,In_0,In_715);
xnor U104 (N_104,In_571,In_771);
and U105 (N_105,In_13,In_48);
xnor U106 (N_106,In_386,In_698);
xnor U107 (N_107,In_1043,In_621);
nor U108 (N_108,In_430,In_1230);
nor U109 (N_109,In_1172,In_92);
nor U110 (N_110,In_1184,In_3);
nand U111 (N_111,In_1167,In_293);
nand U112 (N_112,In_1468,In_1244);
or U113 (N_113,In_912,In_1237);
nand U114 (N_114,In_41,In_1022);
and U115 (N_115,In_1114,In_783);
nor U116 (N_116,In_219,In_1251);
and U117 (N_117,In_923,In_537);
or U118 (N_118,In_416,In_708);
or U119 (N_119,In_1160,In_1);
or U120 (N_120,In_1425,In_1173);
and U121 (N_121,In_30,In_619);
nor U122 (N_122,In_825,In_362);
nor U123 (N_123,In_1252,In_85);
or U124 (N_124,In_197,In_61);
xnor U125 (N_125,In_477,In_520);
and U126 (N_126,In_545,In_1261);
or U127 (N_127,In_1085,In_665);
or U128 (N_128,In_1256,In_478);
and U129 (N_129,In_1359,In_1368);
or U130 (N_130,In_507,In_784);
nand U131 (N_131,In_974,In_1409);
nor U132 (N_132,In_1060,In_369);
nor U133 (N_133,In_218,In_150);
and U134 (N_134,In_1358,In_840);
nand U135 (N_135,In_1144,In_1279);
or U136 (N_136,In_1057,In_508);
nand U137 (N_137,In_878,In_1333);
and U138 (N_138,In_1384,In_685);
xnor U139 (N_139,In_1436,In_1491);
and U140 (N_140,In_410,In_506);
or U141 (N_141,In_742,In_185);
or U142 (N_142,In_389,In_1498);
and U143 (N_143,In_1482,In_644);
xnor U144 (N_144,In_707,In_648);
xor U145 (N_145,In_148,In_1329);
or U146 (N_146,In_348,In_523);
or U147 (N_147,In_1174,In_1463);
nand U148 (N_148,In_826,In_1170);
xor U149 (N_149,In_397,In_81);
or U150 (N_150,In_804,In_942);
nand U151 (N_151,In_261,In_1181);
nand U152 (N_152,In_1229,In_868);
xnor U153 (N_153,In_200,In_592);
nor U154 (N_154,In_512,In_960);
nand U155 (N_155,In_1042,In_625);
and U156 (N_156,In_980,In_370);
and U157 (N_157,In_1024,In_565);
or U158 (N_158,In_301,In_1206);
nand U159 (N_159,In_1293,In_1109);
xor U160 (N_160,In_678,In_516);
xnor U161 (N_161,In_1177,In_157);
and U162 (N_162,In_1095,In_605);
or U163 (N_163,In_896,In_1233);
nand U164 (N_164,In_1291,In_1289);
and U165 (N_165,In_1460,In_472);
or U166 (N_166,In_780,In_855);
and U167 (N_167,In_1161,In_1005);
xnor U168 (N_168,In_1175,In_994);
and U169 (N_169,In_765,In_546);
or U170 (N_170,In_1176,In_1079);
xnor U171 (N_171,In_927,In_319);
and U172 (N_172,In_1003,In_1157);
nand U173 (N_173,In_1053,In_672);
xor U174 (N_174,In_190,In_761);
and U175 (N_175,In_1393,In_1202);
xor U176 (N_176,In_775,In_342);
nand U177 (N_177,In_322,In_1267);
nor U178 (N_178,In_548,In_1275);
nand U179 (N_179,In_1059,In_488);
nand U180 (N_180,In_1285,In_1470);
and U181 (N_181,In_1258,In_1325);
or U182 (N_182,In_745,In_340);
and U183 (N_183,In_1466,In_976);
and U184 (N_184,In_1447,In_955);
and U185 (N_185,In_793,In_1350);
and U186 (N_186,In_1050,In_831);
or U187 (N_187,In_833,In_1434);
or U188 (N_188,In_908,In_1152);
or U189 (N_189,In_722,In_304);
nor U190 (N_190,In_505,In_236);
nand U191 (N_191,In_1322,In_649);
xor U192 (N_192,In_1452,In_1210);
xor U193 (N_193,In_275,In_651);
nor U194 (N_194,In_816,In_531);
or U195 (N_195,In_169,In_222);
xnor U196 (N_196,In_596,In_1145);
nor U197 (N_197,In_1037,In_989);
and U198 (N_198,In_1038,In_9);
nor U199 (N_199,In_653,In_1238);
xor U200 (N_200,In_324,In_660);
nand U201 (N_201,In_492,In_701);
or U202 (N_202,In_786,In_201);
nor U203 (N_203,In_306,In_1045);
xor U204 (N_204,In_1228,In_949);
xor U205 (N_205,In_290,In_861);
or U206 (N_206,In_418,In_1019);
nand U207 (N_207,In_664,In_954);
nor U208 (N_208,In_1002,In_1223);
xor U209 (N_209,In_1101,In_906);
xnor U210 (N_210,In_1182,In_1097);
xor U211 (N_211,In_969,In_688);
nor U212 (N_212,In_316,In_829);
nand U213 (N_213,In_1398,In_1108);
xnor U214 (N_214,In_1487,In_929);
or U215 (N_215,In_80,In_1306);
or U216 (N_216,In_136,In_1316);
or U217 (N_217,In_1016,In_907);
or U218 (N_218,In_788,In_145);
xnor U219 (N_219,In_55,In_429);
xor U220 (N_220,In_338,In_1422);
nor U221 (N_221,In_643,In_876);
nor U222 (N_222,In_1474,In_65);
and U223 (N_223,In_975,In_1070);
nor U224 (N_224,In_1496,In_754);
nor U225 (N_225,In_1483,In_500);
nor U226 (N_226,In_1169,In_207);
xnor U227 (N_227,In_869,In_585);
xnor U228 (N_228,In_1361,In_534);
or U229 (N_229,In_186,In_17);
and U230 (N_230,In_1096,In_373);
or U231 (N_231,In_535,In_1072);
or U232 (N_232,In_2,In_1369);
xnor U233 (N_233,In_1296,In_1335);
nor U234 (N_234,In_1292,In_230);
nand U235 (N_235,In_1103,In_1379);
and U236 (N_236,In_309,In_1451);
xor U237 (N_237,In_628,In_259);
xor U238 (N_238,In_1282,In_1156);
xnor U239 (N_239,In_58,In_1423);
nor U240 (N_240,In_752,In_1104);
nand U241 (N_241,In_278,In_295);
nor U242 (N_242,In_770,In_727);
or U243 (N_243,In_842,In_705);
nor U244 (N_244,In_315,In_175);
nor U245 (N_245,In_343,In_153);
nor U246 (N_246,In_176,In_666);
or U247 (N_247,In_872,In_420);
nor U248 (N_248,In_893,In_552);
xnor U249 (N_249,In_992,In_1165);
nor U250 (N_250,In_160,N_21);
nand U251 (N_251,In_1001,In_1318);
nand U252 (N_252,In_68,In_436);
and U253 (N_253,In_903,In_849);
xnor U254 (N_254,In_1138,In_114);
or U255 (N_255,In_71,In_1259);
xor U256 (N_256,In_528,N_191);
nor U257 (N_257,In_1435,In_986);
nand U258 (N_258,In_1052,In_1105);
or U259 (N_259,In_119,In_396);
or U260 (N_260,In_1338,In_496);
xor U261 (N_261,In_495,In_1139);
nand U262 (N_262,In_1083,N_79);
nand U263 (N_263,In_1426,In_1254);
or U264 (N_264,In_753,In_380);
xnor U265 (N_265,In_1294,In_739);
or U266 (N_266,In_650,In_681);
xnor U267 (N_267,In_774,In_242);
nand U268 (N_268,In_450,In_361);
and U269 (N_269,In_811,In_183);
xor U270 (N_270,In_957,In_35);
and U271 (N_271,In_1471,In_1337);
and U272 (N_272,In_972,In_1234);
xnor U273 (N_273,In_887,In_945);
nand U274 (N_274,In_1007,In_509);
and U275 (N_275,In_946,In_874);
and U276 (N_276,In_417,N_71);
and U277 (N_277,In_593,In_600);
and U278 (N_278,In_828,In_736);
or U279 (N_279,In_471,In_624);
nor U280 (N_280,In_1260,In_1061);
xor U281 (N_281,N_73,In_42);
or U282 (N_282,In_1220,In_1021);
or U283 (N_283,In_941,In_1241);
nand U284 (N_284,In_891,In_171);
and U285 (N_285,In_1268,In_161);
xor U286 (N_286,In_800,N_110);
and U287 (N_287,N_2,In_363);
and U288 (N_288,N_152,In_1123);
or U289 (N_289,In_987,In_608);
nor U290 (N_290,In_144,In_1090);
xor U291 (N_291,In_832,In_642);
or U292 (N_292,N_111,In_74);
xor U293 (N_293,In_400,N_58);
nor U294 (N_294,In_1385,In_694);
xor U295 (N_295,In_892,In_1178);
nor U296 (N_296,In_687,In_262);
nand U297 (N_297,In_696,In_595);
nor U298 (N_298,In_56,In_751);
nand U299 (N_299,In_526,N_122);
xor U300 (N_300,N_160,N_130);
or U301 (N_301,In_735,In_916);
xor U302 (N_302,In_808,In_1004);
xor U303 (N_303,In_156,In_1356);
nor U304 (N_304,In_623,In_963);
nand U305 (N_305,In_1199,In_423);
xor U306 (N_306,In_46,In_817);
xor U307 (N_307,In_1091,In_1277);
or U308 (N_308,N_93,N_141);
and U309 (N_309,In_323,In_895);
or U310 (N_310,In_965,In_1006);
xnor U311 (N_311,In_900,In_82);
and U312 (N_312,In_231,In_378);
or U313 (N_313,In_801,In_298);
nand U314 (N_314,In_1416,In_778);
nor U315 (N_315,In_590,In_26);
nand U316 (N_316,N_146,In_1150);
nand U317 (N_317,N_159,In_932);
nand U318 (N_318,In_321,In_830);
nand U319 (N_319,In_297,In_64);
nor U320 (N_320,N_116,In_544);
or U321 (N_321,In_425,N_121);
nor U322 (N_322,In_844,In_1495);
and U323 (N_323,In_1343,N_28);
nand U324 (N_324,N_106,In_1035);
or U325 (N_325,N_224,N_208);
or U326 (N_326,In_533,In_1437);
nand U327 (N_327,In_457,In_276);
nor U328 (N_328,In_382,In_313);
nor U329 (N_329,N_45,In_1272);
nand U330 (N_330,In_217,In_1118);
xnor U331 (N_331,In_1263,In_1159);
and U332 (N_332,In_462,N_226);
and U333 (N_333,In_821,N_15);
nor U334 (N_334,In_966,N_44);
xnor U335 (N_335,In_108,In_1340);
xor U336 (N_336,N_68,In_790);
or U337 (N_337,N_137,In_766);
or U338 (N_338,In_748,In_1065);
or U339 (N_339,In_982,N_173);
nor U340 (N_340,In_803,In_549);
or U341 (N_341,N_119,In_1081);
xor U342 (N_342,N_78,N_244);
xor U343 (N_343,In_198,In_689);
or U344 (N_344,In_210,In_104);
or U345 (N_345,In_951,In_971);
nand U346 (N_346,N_176,In_1448);
nand U347 (N_347,In_839,In_257);
xor U348 (N_348,In_381,In_985);
nor U349 (N_349,In_515,In_1168);
nor U350 (N_350,In_583,N_16);
or U351 (N_351,In_376,In_195);
nand U352 (N_352,N_216,N_230);
or U353 (N_353,In_679,N_87);
or U354 (N_354,In_738,In_962);
and U355 (N_355,In_1281,In_938);
xnor U356 (N_356,N_113,In_854);
and U357 (N_357,In_725,In_1362);
or U358 (N_358,In_377,In_859);
and U359 (N_359,In_279,In_173);
xnor U360 (N_360,N_193,In_20);
nand U361 (N_361,In_7,In_168);
xor U362 (N_362,In_1269,N_194);
xor U363 (N_363,In_1209,In_292);
nand U364 (N_364,In_885,In_432);
or U365 (N_365,In_1373,In_240);
nor U366 (N_366,In_163,In_703);
and U367 (N_367,In_776,N_185);
nor U368 (N_368,In_431,In_112);
xor U369 (N_369,N_213,In_852);
and U370 (N_370,In_1493,In_1226);
nand U371 (N_371,In_921,In_851);
or U372 (N_372,N_105,In_820);
nand U373 (N_373,In_346,In_1453);
xor U374 (N_374,In_209,In_630);
nand U375 (N_375,In_265,In_627);
nand U376 (N_376,In_636,N_150);
xnor U377 (N_377,In_44,In_194);
and U378 (N_378,N_144,In_543);
xor U379 (N_379,N_82,In_387);
or U380 (N_380,In_998,N_183);
nor U381 (N_381,In_447,In_1353);
nand U382 (N_382,N_240,In_719);
nand U383 (N_383,In_939,In_997);
nor U384 (N_384,In_1255,In_682);
xnor U385 (N_385,In_445,In_1128);
nand U386 (N_386,N_30,In_1106);
and U387 (N_387,In_116,In_690);
xor U388 (N_388,N_210,In_622);
nor U389 (N_389,In_728,N_232);
xnor U390 (N_390,In_806,In_1056);
xnor U391 (N_391,In_45,In_354);
nand U392 (N_392,In_170,In_1286);
nor U393 (N_393,N_242,In_87);
nand U394 (N_394,In_680,In_62);
and U395 (N_395,In_246,In_1330);
nor U396 (N_396,In_444,In_146);
nand U397 (N_397,In_1321,In_248);
or U398 (N_398,In_710,N_236);
nor U399 (N_399,In_180,N_163);
and U400 (N_400,In_225,In_43);
xnor U401 (N_401,In_36,In_167);
nand U402 (N_402,In_540,In_76);
xor U403 (N_403,In_11,In_1488);
nand U404 (N_404,In_184,In_455);
nand U405 (N_405,In_439,In_853);
xnor U406 (N_406,In_603,In_586);
xor U407 (N_407,In_578,In_281);
or U408 (N_408,In_602,In_1049);
xnor U409 (N_409,In_129,In_1148);
or U410 (N_410,In_199,In_384);
nand U411 (N_411,In_29,In_368);
xnor U412 (N_412,In_814,In_1288);
nand U413 (N_413,In_918,In_1454);
and U414 (N_414,In_124,In_196);
nor U415 (N_415,In_294,In_332);
xnor U416 (N_416,N_174,In_31);
nand U417 (N_417,In_674,In_208);
nand U418 (N_418,In_658,N_132);
nand U419 (N_419,In_1240,In_440);
or U420 (N_420,In_1084,In_6);
or U421 (N_421,In_310,In_936);
and U422 (N_422,In_575,In_1300);
nand U423 (N_423,In_1399,N_126);
nor U424 (N_424,In_314,In_677);
or U425 (N_425,In_1438,In_1116);
nor U426 (N_426,In_1407,N_157);
nand U427 (N_427,In_922,In_884);
or U428 (N_428,In_563,N_48);
nand U429 (N_429,In_399,In_647);
and U430 (N_430,In_950,In_334);
and U431 (N_431,In_1071,In_32);
or U432 (N_432,In_883,In_1421);
or U433 (N_433,In_1068,In_882);
nand U434 (N_434,In_1339,In_347);
and U435 (N_435,In_408,N_20);
or U436 (N_436,In_12,In_1490);
or U437 (N_437,N_241,In_662);
nor U438 (N_438,N_39,In_1283);
and U439 (N_439,In_629,In_931);
nand U440 (N_440,In_463,In_351);
xor U441 (N_441,In_530,N_142);
nor U442 (N_442,In_888,In_718);
nor U443 (N_443,N_203,In_8);
nand U444 (N_444,In_494,In_609);
or U445 (N_445,In_253,In_105);
nor U446 (N_446,In_1370,N_211);
or U447 (N_447,In_1367,In_809);
nand U448 (N_448,In_1180,In_860);
xor U449 (N_449,In_977,N_175);
and U450 (N_450,In_1376,In_1033);
and U451 (N_451,In_456,N_53);
and U452 (N_452,N_70,N_35);
xnor U453 (N_453,In_799,In_433);
nor U454 (N_454,In_1395,In_287);
and U455 (N_455,N_89,In_1080);
xor U456 (N_456,In_1265,In_93);
or U457 (N_457,N_206,In_1187);
nand U458 (N_458,In_746,In_919);
or U459 (N_459,N_128,N_22);
and U460 (N_460,In_867,N_98);
and U461 (N_461,In_1413,In_850);
and U462 (N_462,In_1047,In_1135);
or U463 (N_463,In_390,N_56);
xor U464 (N_464,In_570,In_756);
or U465 (N_465,N_136,In_606);
nor U466 (N_466,N_103,In_729);
nand U467 (N_467,N_23,In_483);
and U468 (N_468,In_743,In_1382);
xnor U469 (N_469,In_614,N_246);
xor U470 (N_470,In_125,In_704);
and U471 (N_471,In_791,In_318);
xnor U472 (N_472,In_73,In_943);
and U473 (N_473,In_928,In_1221);
or U474 (N_474,In_713,In_1069);
or U475 (N_475,In_574,In_1132);
nor U476 (N_476,In_1025,In_1023);
nand U477 (N_477,In_291,N_200);
xnor U478 (N_478,In_1401,In_1355);
xor U479 (N_479,N_75,In_317);
nor U480 (N_480,In_1149,In_1485);
nand U481 (N_481,In_409,In_383);
nand U482 (N_482,N_26,In_519);
nand U483 (N_483,In_475,In_875);
xnor U484 (N_484,In_588,In_1064);
xor U485 (N_485,In_1280,In_1499);
nor U486 (N_486,In_835,In_402);
and U487 (N_487,In_834,In_300);
and U488 (N_488,In_1377,N_69);
or U489 (N_489,N_102,In_979);
and U490 (N_490,In_769,In_326);
and U491 (N_491,In_795,In_661);
or U492 (N_492,In_1459,In_59);
xor U493 (N_493,In_732,In_126);
nor U494 (N_494,In_249,In_47);
xor U495 (N_495,In_1074,In_1028);
and U496 (N_496,In_522,N_235);
or U497 (N_497,In_568,In_529);
nand U498 (N_498,In_1186,In_1314);
xor U499 (N_499,In_358,In_83);
nand U500 (N_500,N_228,In_940);
nand U501 (N_501,In_518,In_967);
nor U502 (N_502,In_902,In_1107);
and U503 (N_503,In_52,In_1469);
nand U504 (N_504,In_131,N_86);
nand U505 (N_505,N_454,N_360);
xnor U506 (N_506,N_263,N_96);
and U507 (N_507,In_1270,N_43);
xor U508 (N_508,N_380,In_355);
or U509 (N_509,In_716,In_102);
nand U510 (N_510,In_1364,In_759);
or U511 (N_511,N_428,In_758);
or U512 (N_512,N_85,In_371);
xor U513 (N_513,In_838,In_1029);
nand U514 (N_514,N_95,N_301);
and U515 (N_515,N_46,In_75);
and U516 (N_516,In_1231,N_425);
nand U517 (N_517,N_294,In_120);
or U518 (N_518,N_385,N_371);
nor U519 (N_519,In_422,N_375);
nand U520 (N_520,In_772,In_1430);
and U521 (N_521,In_525,In_1331);
nor U522 (N_522,In_1262,In_1298);
or U523 (N_523,In_140,N_483);
and U524 (N_524,N_316,In_1232);
or U525 (N_525,N_91,N_397);
nand U526 (N_526,In_23,In_215);
or U527 (N_527,In_1011,In_1134);
or U528 (N_528,In_285,In_107);
or U529 (N_529,In_1126,In_541);
and U530 (N_530,N_265,In_490);
nor U531 (N_531,N_239,In_1066);
and U532 (N_532,In_587,N_457);
nand U533 (N_533,In_1075,In_149);
nand U534 (N_534,In_449,N_223);
xor U535 (N_535,N_287,N_237);
xor U536 (N_536,N_391,In_686);
xor U537 (N_537,N_318,N_38);
or U538 (N_538,In_819,In_283);
xor U539 (N_539,N_298,N_456);
and U540 (N_540,N_84,In_767);
or U541 (N_541,In_345,In_1461);
and U542 (N_542,In_638,N_461);
or U543 (N_543,In_88,In_1391);
nor U544 (N_544,In_426,N_229);
or U545 (N_545,N_178,In_311);
and U546 (N_546,In_211,N_195);
nand U547 (N_547,In_762,In_1204);
xnor U548 (N_548,In_375,In_905);
xnor U549 (N_549,In_873,N_248);
or U550 (N_550,N_233,In_657);
nand U551 (N_551,N_1,N_169);
xor U552 (N_552,In_1308,N_444);
nand U553 (N_553,In_18,In_558);
or U554 (N_554,N_282,In_1445);
or U555 (N_555,N_349,N_347);
nand U556 (N_556,N_495,N_204);
or U557 (N_557,In_1349,N_114);
nor U558 (N_558,In_1328,N_383);
xnor U559 (N_559,In_1478,N_463);
nor U560 (N_560,N_134,In_721);
nand U561 (N_561,In_266,In_398);
nor U562 (N_562,In_1185,In_1051);
and U563 (N_563,In_67,In_14);
nor U564 (N_564,In_511,N_260);
and U565 (N_565,In_787,In_10);
nand U566 (N_566,In_749,N_418);
or U567 (N_567,In_286,In_1222);
or U568 (N_568,N_470,In_1346);
and U569 (N_569,In_427,In_1127);
and U570 (N_570,In_1383,N_443);
and U571 (N_571,In_214,N_382);
xor U572 (N_572,N_24,In_601);
or U573 (N_573,N_27,In_865);
nand U574 (N_574,N_65,In_1098);
nand U575 (N_575,N_481,N_479);
xnor U576 (N_576,In_1030,In_115);
nor U577 (N_577,In_837,In_205);
xnor U578 (N_578,In_618,In_352);
or U579 (N_579,In_1100,In_37);
nand U580 (N_580,N_11,N_429);
nor U581 (N_581,In_428,In_421);
nand U582 (N_582,N_414,N_390);
nand U583 (N_583,In_158,N_459);
xnor U584 (N_584,In_539,In_845);
nand U585 (N_585,In_353,In_734);
nand U586 (N_586,In_1131,In_847);
nand U587 (N_587,In_49,N_372);
nand U588 (N_588,In_70,In_1336);
xor U589 (N_589,N_450,N_36);
and U590 (N_590,In_909,In_188);
and U591 (N_591,In_40,In_141);
and U592 (N_592,In_1121,In_604);
or U593 (N_593,In_395,In_827);
and U594 (N_594,N_368,In_391);
or U595 (N_595,N_147,In_118);
and U596 (N_596,N_217,In_802);
or U597 (N_597,In_700,In_763);
or U598 (N_598,N_135,In_1044);
nand U599 (N_599,N_162,In_1190);
nand U600 (N_600,In_96,In_128);
and U601 (N_601,N_381,In_1424);
or U602 (N_602,N_170,N_275);
and U603 (N_603,In_234,In_594);
xnor U604 (N_604,N_285,In_536);
nor U605 (N_605,In_559,N_149);
and U606 (N_606,In_1458,N_437);
nor U607 (N_607,N_120,In_1307);
nand U608 (N_608,N_231,In_1332);
or U609 (N_609,In_956,In_359);
or U610 (N_610,N_12,N_139);
nor U611 (N_611,In_1215,In_424);
and U612 (N_612,In_164,N_467);
nor U613 (N_613,In_1197,N_482);
nor U614 (N_614,N_346,N_222);
nor U615 (N_615,N_5,In_1036);
or U616 (N_616,N_445,In_697);
nor U617 (N_617,N_336,In_877);
xor U618 (N_618,In_532,N_186);
xnor U619 (N_619,N_430,N_407);
xor U620 (N_620,In_1054,In_824);
or U621 (N_621,In_1431,In_1208);
nand U622 (N_622,In_39,In_1432);
xnor U623 (N_623,In_1481,N_31);
nand U624 (N_624,In_454,N_225);
xor U625 (N_625,In_178,In_933);
nand U626 (N_626,In_1201,In_1196);
or U627 (N_627,In_1341,In_1193);
xor U628 (N_628,N_6,N_440);
nand U629 (N_629,N_192,In_988);
nor U630 (N_630,N_370,In_1420);
xnor U631 (N_631,In_503,In_1189);
nand U632 (N_632,In_308,N_496);
nor U633 (N_633,N_484,N_51);
nor U634 (N_634,In_484,In_1086);
and U635 (N_635,In_1351,In_451);
and U636 (N_636,In_1143,In_1194);
xor U637 (N_637,In_233,N_376);
and U638 (N_638,N_328,In_1304);
and U639 (N_639,N_267,N_497);
xnor U640 (N_640,N_42,N_269);
or U641 (N_641,In_235,In_1248);
nor U642 (N_642,In_1433,N_409);
nor U643 (N_643,In_610,In_244);
and U644 (N_644,In_252,N_251);
or U645 (N_645,In_1371,N_488);
and U646 (N_646,N_266,N_337);
xnor U647 (N_647,In_1155,N_464);
or U648 (N_648,N_280,N_357);
nand U649 (N_649,In_481,N_412);
nand U650 (N_650,N_389,N_158);
nor U651 (N_651,In_862,In_1119);
xor U652 (N_652,In_224,N_476);
nand U653 (N_653,In_572,N_62);
nand U654 (N_654,N_289,In_777);
and U655 (N_655,In_1494,N_491);
nand U656 (N_656,In_1387,N_306);
nor U657 (N_657,N_311,In_1017);
xnor U658 (N_658,In_448,N_129);
nor U659 (N_659,N_164,N_261);
xor U660 (N_660,In_223,N_345);
xor U661 (N_661,In_999,In_897);
or U662 (N_662,N_40,In_617);
nor U663 (N_663,In_1113,N_92);
or U664 (N_664,N_100,In_913);
nor U665 (N_665,N_319,N_177);
nor U666 (N_666,N_247,In_435);
nor U667 (N_667,In_915,In_1301);
and U668 (N_668,In_438,In_591);
nor U669 (N_669,N_325,In_538);
nand U670 (N_670,N_471,N_0);
and U671 (N_671,In_1457,N_295);
and U672 (N_672,N_292,In_768);
and U673 (N_673,In_781,N_55);
nand U674 (N_674,In_794,In_1032);
xnor U675 (N_675,N_52,In_562);
nand U676 (N_676,In_63,N_256);
or U677 (N_677,In_385,N_436);
or U678 (N_678,N_281,In_1110);
or U679 (N_679,In_487,In_228);
or U680 (N_680,N_10,In_106);
or U681 (N_681,N_379,N_215);
xnor U682 (N_682,In_202,N_438);
or U683 (N_683,N_377,N_97);
nor U684 (N_684,N_300,In_1455);
or U685 (N_685,N_303,N_350);
and U686 (N_686,N_140,In_1273);
and U687 (N_687,In_117,In_1429);
or U688 (N_688,In_159,N_378);
nor U689 (N_689,N_83,In_812);
and U690 (N_690,In_1214,In_810);
and U691 (N_691,In_1276,In_983);
or U692 (N_692,In_1410,In_1397);
nand U693 (N_693,In_264,N_171);
xor U694 (N_694,In_675,In_1227);
and U695 (N_695,N_131,N_180);
and U696 (N_696,N_413,In_1018);
nand U697 (N_697,In_97,N_331);
nor U698 (N_698,In_94,In_1166);
or U699 (N_699,In_4,N_4);
nor U700 (N_700,In_1067,N_104);
nor U701 (N_701,N_81,In_547);
or U702 (N_702,N_270,N_394);
and U703 (N_703,In_993,N_451);
xor U704 (N_704,N_353,In_567);
and U705 (N_705,N_458,In_646);
nor U706 (N_706,N_88,In_401);
nand U707 (N_707,N_478,N_313);
xor U708 (N_708,N_17,N_181);
xor U709 (N_709,In_726,N_57);
nor U710 (N_710,In_1404,N_227);
nor U711 (N_711,In_1400,In_917);
and U712 (N_712,In_86,In_673);
and U713 (N_713,In_626,In_84);
xor U714 (N_714,N_477,In_1014);
xor U715 (N_715,In_1125,N_364);
xnor U716 (N_716,N_486,In_464);
xor U717 (N_717,In_19,In_239);
nand U718 (N_718,In_341,In_926);
nor U719 (N_719,In_329,In_702);
or U720 (N_720,In_241,In_553);
nor U721 (N_721,N_32,In_1163);
nand U722 (N_722,In_469,In_551);
nor U723 (N_723,N_421,N_367);
nand U724 (N_724,In_904,In_947);
and U725 (N_725,N_138,N_369);
xnor U726 (N_726,N_420,In_493);
xor U727 (N_727,In_415,N_309);
or U728 (N_728,In_255,N_393);
nand U729 (N_729,N_123,N_76);
and U730 (N_730,In_659,N_387);
and U731 (N_731,In_270,In_805);
nor U732 (N_732,N_417,In_733);
xnor U733 (N_733,In_656,N_67);
or U734 (N_734,N_446,N_474);
nand U735 (N_735,In_406,In_393);
xor U736 (N_736,N_422,In_557);
xnor U737 (N_737,In_394,In_302);
xor U738 (N_738,In_1323,In_894);
or U739 (N_739,In_53,In_147);
or U740 (N_740,In_1158,N_148);
or U741 (N_741,In_1191,N_351);
nand U742 (N_742,In_442,N_314);
nor U743 (N_743,N_431,In_607);
and U744 (N_744,N_419,In_1041);
and U745 (N_745,In_296,N_34);
nand U746 (N_746,In_1326,In_1122);
nor U747 (N_747,N_334,In_502);
and U748 (N_748,In_1077,In_1365);
and U749 (N_749,In_1133,N_453);
xor U750 (N_750,N_468,N_365);
and U751 (N_751,N_675,N_728);
or U752 (N_752,In_263,N_684);
and U753 (N_753,N_502,In_1243);
or U754 (N_754,N_361,In_1313);
nor U755 (N_755,N_50,In_1473);
nand U756 (N_756,In_392,In_744);
or U757 (N_757,In_879,N_613);
nand U758 (N_758,N_212,In_50);
nor U759 (N_759,In_611,N_60);
nand U760 (N_760,N_625,In_403);
nand U761 (N_761,In_1440,N_492);
nor U762 (N_762,N_670,In_668);
xor U763 (N_763,N_523,In_573);
and U764 (N_764,N_439,N_646);
and U765 (N_765,N_290,N_631);
xnor U766 (N_766,N_665,N_663);
xor U767 (N_767,N_424,N_435);
nor U768 (N_768,N_615,In_1345);
nor U769 (N_769,In_1480,N_538);
nor U770 (N_770,N_628,In_1082);
nand U771 (N_771,In_103,In_1419);
nand U772 (N_772,N_688,N_745);
or U773 (N_773,In_271,N_220);
and U774 (N_774,N_644,In_1046);
and U775 (N_775,N_243,N_589);
xnor U776 (N_776,N_354,N_343);
xor U777 (N_777,N_513,N_530);
nand U778 (N_778,N_214,N_168);
or U779 (N_779,N_259,N_277);
or U780 (N_780,In_414,N_645);
nand U781 (N_781,In_691,In_441);
and U782 (N_782,N_592,N_472);
nand U783 (N_783,In_1211,N_549);
xnor U784 (N_784,In_1246,N_410);
and U785 (N_785,In_57,N_587);
or U786 (N_786,N_59,N_218);
nor U787 (N_787,N_499,In_1380);
nand U788 (N_788,N_706,In_699);
nand U789 (N_789,N_386,N_503);
nor U790 (N_790,In_1235,N_677);
and U791 (N_791,In_1089,N_524);
nand U792 (N_792,In_203,In_1394);
xor U793 (N_793,N_61,N_332);
xor U794 (N_794,In_499,N_661);
and U795 (N_795,N_18,In_1386);
nor U796 (N_796,N_542,In_1405);
and U797 (N_797,In_1449,In_1129);
nor U798 (N_798,In_996,In_277);
xor U799 (N_799,N_520,In_1392);
xnor U800 (N_800,N_599,N_356);
xor U801 (N_801,In_132,In_130);
and U802 (N_802,In_1015,In_38);
nor U803 (N_803,N_432,N_465);
nand U804 (N_804,In_683,In_1489);
and U805 (N_805,N_304,In_581);
nor U806 (N_806,N_655,N_209);
xnor U807 (N_807,In_282,N_278);
or U808 (N_808,In_1147,In_934);
xnor U809 (N_809,In_1312,In_655);
nor U810 (N_810,N_54,N_299);
nor U811 (N_811,In_172,N_643);
xnor U812 (N_812,N_531,In_320);
and U813 (N_813,In_634,N_545);
nand U814 (N_814,In_337,N_339);
or U815 (N_815,In_465,N_7);
or U816 (N_816,N_585,In_307);
nor U817 (N_817,N_603,N_609);
nand U818 (N_818,In_486,In_1247);
or U819 (N_819,In_846,N_532);
or U820 (N_820,In_717,In_221);
xor U821 (N_821,N_358,In_1354);
nand U822 (N_822,In_1076,N_279);
and U823 (N_823,N_252,N_307);
nor U824 (N_824,N_565,In_948);
nor U825 (N_825,In_181,N_683);
and U826 (N_826,N_741,N_154);
or U827 (N_827,N_709,In_1112);
nor U828 (N_828,N_711,N_533);
xor U829 (N_829,N_500,In_461);
nand U830 (N_830,N_553,In_366);
and U831 (N_831,N_600,N_253);
nor U832 (N_832,N_355,N_634);
xor U833 (N_833,In_177,N_546);
or U834 (N_834,In_1412,N_448);
and U835 (N_835,In_639,N_340);
nor U836 (N_836,N_401,N_554);
xor U837 (N_837,N_704,N_501);
xor U838 (N_838,N_384,N_199);
or U839 (N_839,N_548,N_535);
nand U840 (N_840,N_49,In_981);
and U841 (N_841,N_161,N_656);
nor U842 (N_842,N_466,In_1140);
and U843 (N_843,N_221,In_22);
nor U844 (N_844,N_489,In_24);
or U845 (N_845,N_514,N_708);
or U846 (N_846,In_443,N_629);
or U847 (N_847,N_713,In_137);
nand U848 (N_848,N_258,In_667);
nor U849 (N_849,In_952,N_274);
nor U850 (N_850,N_189,N_664);
nand U851 (N_851,In_797,N_598);
or U852 (N_852,N_597,N_408);
or U853 (N_853,In_1162,In_1219);
or U854 (N_854,In_90,N_201);
or U855 (N_855,In_671,In_995);
xnor U856 (N_856,N_544,In_243);
or U857 (N_857,In_1239,N_701);
xor U858 (N_858,In_747,N_680);
nor U859 (N_859,In_1236,In_880);
nand U860 (N_860,N_526,N_66);
or U861 (N_861,In_485,N_678);
xnor U862 (N_862,N_725,In_349);
or U863 (N_863,N_262,In_1278);
xnor U864 (N_864,N_99,In_15);
or U865 (N_865,N_272,In_254);
nand U866 (N_866,N_584,In_91);
or U867 (N_867,N_543,In_1327);
xnor U868 (N_868,In_1475,In_723);
and U869 (N_869,In_1411,N_145);
or U870 (N_870,N_403,N_507);
nor U871 (N_871,N_550,N_616);
or U872 (N_872,In_953,N_652);
and U873 (N_873,N_540,N_373);
or U874 (N_874,In_1154,N_617);
nor U875 (N_875,In_333,In_312);
nand U876 (N_876,In_597,N_341);
and U877 (N_877,In_789,N_167);
and U878 (N_878,N_187,In_901);
xnor U879 (N_879,N_731,In_978);
xor U880 (N_880,In_755,N_33);
nor U881 (N_881,N_747,N_567);
xor U882 (N_882,N_581,N_344);
nand U883 (N_883,N_516,N_698);
and U884 (N_884,In_1198,N_101);
nand U885 (N_885,N_722,N_254);
nor U886 (N_886,N_433,N_515);
nor U887 (N_887,N_310,In_1120);
nand U888 (N_888,N_672,N_321);
xnor U889 (N_889,N_143,N_297);
xnor U890 (N_890,N_547,In_27);
or U891 (N_891,N_635,In_1303);
and U892 (N_892,In_863,N_156);
or U893 (N_893,N_653,N_712);
or U894 (N_894,N_674,N_723);
or U895 (N_895,In_886,N_566);
and U896 (N_896,N_707,N_579);
or U897 (N_897,In_924,In_288);
xor U898 (N_898,N_124,N_742);
nor U899 (N_899,In_268,N_527);
and U900 (N_900,In_357,N_19);
xor U901 (N_901,N_574,N_583);
nand U902 (N_902,N_117,In_1357);
or U903 (N_903,N_506,In_620);
xnor U904 (N_904,In_54,N_250);
xnor U905 (N_905,In_1309,In_458);
nand U906 (N_906,N_423,In_1446);
or U907 (N_907,N_234,In_28);
and U908 (N_908,N_462,In_1102);
xnor U909 (N_909,In_1344,N_729);
or U910 (N_910,In_521,In_405);
and U911 (N_911,N_667,N_649);
and U912 (N_912,N_697,N_607);
xor U913 (N_913,N_658,N_359);
nor U914 (N_914,N_727,N_518);
nand U915 (N_915,N_608,N_650);
and U916 (N_916,N_362,N_434);
and U917 (N_917,N_315,In_599);
or U918 (N_918,In_497,In_1058);
nor U919 (N_919,N_718,In_1467);
nand U920 (N_920,N_586,N_366);
nand U921 (N_921,In_134,N_730);
nand U922 (N_922,N_402,N_322);
nand U923 (N_923,In_712,In_1000);
or U924 (N_924,In_1479,N_312);
nor U925 (N_925,N_541,In_95);
nand U926 (N_926,N_396,N_659);
nand U927 (N_927,N_330,In_1378);
or U928 (N_928,N_172,N_692);
xor U929 (N_929,N_198,N_657);
or U930 (N_930,N_560,N_196);
or U931 (N_931,N_571,N_539);
or U932 (N_932,In_1360,In_127);
and U933 (N_933,N_639,N_739);
xnor U934 (N_934,N_165,N_473);
xnor U935 (N_935,In_714,N_691);
nand U936 (N_936,N_41,N_626);
xor U937 (N_937,N_696,In_51);
xor U938 (N_938,In_1031,N_679);
nor U939 (N_939,In_227,N_529);
xnor U940 (N_940,N_504,In_335);
or U941 (N_941,N_575,In_1111);
xnor U942 (N_942,N_460,N_638);
and U943 (N_943,N_525,N_320);
and U944 (N_944,N_669,N_284);
nand U945 (N_945,N_681,N_77);
or U946 (N_946,N_323,In_1136);
or U947 (N_947,In_576,N_155);
or U948 (N_948,N_740,In_232);
xnor U949 (N_949,N_534,N_569);
xor U950 (N_950,N_293,In_1464);
nor U951 (N_951,N_184,N_426);
xor U952 (N_952,N_449,N_642);
and U953 (N_953,In_857,N_363);
and U954 (N_954,N_109,N_288);
xnor U955 (N_955,N_268,N_699);
xor U956 (N_956,In_336,In_555);
and U957 (N_957,In_1264,N_333);
and U958 (N_958,N_416,N_654);
or U959 (N_959,In_836,N_559);
xnor U960 (N_960,N_400,In_191);
nor U961 (N_961,In_1319,N_564);
and U962 (N_962,N_286,In_1039);
and U963 (N_963,In_1253,N_612);
xor U964 (N_964,In_1141,N_694);
nor U965 (N_965,N_562,N_264);
xor U966 (N_966,N_14,N_633);
or U967 (N_967,In_1009,In_1414);
nor U968 (N_968,In_1472,N_291);
nand U969 (N_969,In_1266,In_920);
and U970 (N_970,N_3,N_207);
nand U971 (N_971,In_711,In_466);
xor U972 (N_972,In_1200,N_510);
nand U973 (N_973,In_491,In_670);
nor U974 (N_974,In_419,N_735);
or U975 (N_975,In_1372,In_498);
or U976 (N_976,In_542,In_480);
and U977 (N_977,In_566,In_388);
xnor U978 (N_978,N_594,In_123);
nand U979 (N_979,In_1216,In_273);
nand U980 (N_980,In_616,N_327);
or U981 (N_981,N_338,N_245);
nand U982 (N_982,N_606,In_871);
xnor U983 (N_983,N_743,N_632);
nand U984 (N_984,N_509,N_687);
and U985 (N_985,In_165,In_121);
nor U986 (N_986,N_411,N_29);
xor U987 (N_987,N_74,N_257);
nand U988 (N_988,N_399,In_589);
xnor U989 (N_989,In_870,N_614);
or U990 (N_990,N_442,N_455);
and U991 (N_991,N_153,N_427);
nor U992 (N_992,N_563,N_703);
nor U993 (N_993,In_1484,N_705);
nor U994 (N_994,N_179,N_577);
nor U995 (N_995,In_764,N_552);
xor U996 (N_996,In_580,N_591);
xor U997 (N_997,N_202,N_630);
or U998 (N_998,In_206,In_554);
and U999 (N_999,In_796,N_485);
or U1000 (N_1000,N_13,In_360);
nor U1001 (N_1001,N_949,N_984);
nand U1002 (N_1002,In_813,N_788);
nor U1003 (N_1003,N_981,N_825);
xnor U1004 (N_1004,N_480,N_794);
nor U1005 (N_1005,In_584,In_1302);
xnor U1006 (N_1006,N_878,N_919);
xnor U1007 (N_1007,N_786,N_811);
nand U1008 (N_1008,N_950,N_537);
and U1009 (N_1009,N_975,In_99);
or U1010 (N_1010,N_960,N_800);
xor U1011 (N_1011,N_829,N_576);
or U1012 (N_1012,N_816,N_415);
or U1013 (N_1013,N_795,N_782);
or U1014 (N_1014,In_413,N_582);
nor U1015 (N_1015,N_997,N_989);
or U1016 (N_1016,N_737,N_108);
and U1017 (N_1017,N_792,In_269);
or U1018 (N_1018,N_865,N_570);
or U1019 (N_1019,N_980,N_920);
and U1020 (N_1020,N_882,N_901);
xnor U1021 (N_1021,N_849,N_889);
nor U1022 (N_1022,N_700,N_686);
or U1023 (N_1023,N_760,N_807);
or U1024 (N_1024,N_778,N_374);
and U1025 (N_1025,N_884,N_335);
and U1026 (N_1026,N_621,N_819);
and U1027 (N_1027,N_803,N_846);
xor U1028 (N_1028,In_5,N_871);
or U1029 (N_1029,N_441,In_331);
or U1030 (N_1030,In_133,N_648);
nor U1031 (N_1031,N_219,N_127);
and U1032 (N_1032,N_831,In_1055);
nor U1033 (N_1033,N_886,In_1406);
or U1034 (N_1034,N_944,N_863);
and U1035 (N_1035,N_388,N_757);
nor U1036 (N_1036,N_519,N_899);
or U1037 (N_1037,N_750,N_915);
nand U1038 (N_1038,N_815,N_996);
or U1039 (N_1039,N_37,N_494);
nor U1040 (N_1040,N_982,N_879);
nand U1041 (N_1041,N_283,In_258);
xor U1042 (N_1042,N_904,N_992);
xor U1043 (N_1043,N_787,N_832);
nor U1044 (N_1044,In_914,N_765);
nand U1045 (N_1045,N_964,N_693);
nand U1046 (N_1046,N_604,N_593);
nand U1047 (N_1047,In_612,N_115);
xor U1048 (N_1048,In_1443,N_767);
xnor U1049 (N_1049,N_798,In_220);
xor U1050 (N_1050,N_805,In_910);
nor U1051 (N_1051,N_715,N_862);
or U1052 (N_1052,N_945,N_557);
or U1053 (N_1053,N_490,N_977);
nand U1054 (N_1054,N_536,N_676);
nand U1055 (N_1055,N_726,N_893);
xnor U1056 (N_1056,In_256,N_806);
or U1057 (N_1057,In_501,N_768);
xor U1058 (N_1058,N_808,N_936);
xnor U1059 (N_1059,N_682,In_720);
and U1060 (N_1060,N_973,N_776);
and U1061 (N_1061,N_752,N_857);
nand U1062 (N_1062,N_967,N_721);
or U1063 (N_1063,N_72,N_627);
xor U1064 (N_1064,In_866,N_888);
nand U1065 (N_1065,N_796,N_761);
nor U1066 (N_1066,N_818,N_935);
nand U1067 (N_1067,N_923,In_143);
nor U1068 (N_1068,N_308,N_870);
nand U1069 (N_1069,N_942,In_1408);
nand U1070 (N_1070,N_820,In_663);
or U1071 (N_1071,N_452,In_958);
xnor U1072 (N_1072,N_637,In_1034);
nand U1073 (N_1073,N_107,N_758);
and U1074 (N_1074,N_753,N_809);
xor U1075 (N_1075,N_125,N_8);
and U1076 (N_1076,N_955,N_671);
or U1077 (N_1077,N_873,In_1192);
nor U1078 (N_1078,N_907,N_80);
xnor U1079 (N_1079,N_916,N_342);
or U1080 (N_1080,N_965,N_25);
xnor U1081 (N_1081,N_573,N_970);
xor U1082 (N_1082,N_948,N_605);
nand U1083 (N_1083,N_998,In_556);
or U1084 (N_1084,N_939,N_521);
nand U1085 (N_1085,N_914,N_859);
nor U1086 (N_1086,N_517,N_881);
nand U1087 (N_1087,N_744,N_732);
nor U1088 (N_1088,N_848,N_395);
or U1089 (N_1089,In_579,N_190);
and U1090 (N_1090,N_601,N_733);
or U1091 (N_1091,N_572,N_854);
nor U1092 (N_1092,N_611,N_668);
and U1093 (N_1093,N_951,N_766);
nor U1094 (N_1094,N_962,In_1171);
and U1095 (N_1095,N_769,N_837);
nand U1096 (N_1096,N_954,In_193);
xor U1097 (N_1097,N_911,In_990);
or U1098 (N_1098,N_205,N_910);
xnor U1099 (N_1099,N_824,N_814);
or U1100 (N_1100,N_717,N_918);
and U1101 (N_1101,In_60,N_690);
nand U1102 (N_1102,N_590,In_1205);
or U1103 (N_1103,N_821,N_685);
xnor U1104 (N_1104,N_166,N_928);
nand U1105 (N_1105,N_930,N_983);
or U1106 (N_1106,N_913,In_305);
or U1107 (N_1107,N_941,N_588);
nor U1108 (N_1108,N_511,In_514);
nor U1109 (N_1109,In_1348,In_238);
or U1110 (N_1110,N_861,N_892);
xor U1111 (N_1111,N_522,In_1427);
nand U1112 (N_1112,In_641,N_968);
nand U1113 (N_1113,In_212,In_135);
nand U1114 (N_1114,N_791,In_1224);
and U1115 (N_1115,N_898,N_620);
nand U1116 (N_1116,N_763,N_112);
nor U1117 (N_1117,In_1324,N_469);
or U1118 (N_1118,N_780,N_802);
and U1119 (N_1119,In_69,N_775);
nand U1120 (N_1120,N_773,N_556);
nor U1121 (N_1121,N_961,N_487);
nor U1122 (N_1122,N_835,N_770);
nor U1123 (N_1123,N_781,N_969);
and U1124 (N_1124,N_963,N_673);
xor U1125 (N_1125,N_797,N_905);
and U1126 (N_1126,N_512,N_249);
nor U1127 (N_1127,N_937,N_799);
or U1128 (N_1128,In_152,N_874);
or U1129 (N_1129,N_895,N_958);
or U1130 (N_1130,In_737,N_595);
xnor U1131 (N_1131,N_720,N_636);
or U1132 (N_1132,In_473,N_891);
or U1133 (N_1133,N_398,N_271);
xnor U1134 (N_1134,N_842,N_926);
nor U1135 (N_1135,N_352,N_755);
nor U1136 (N_1136,N_880,N_561);
and U1137 (N_1137,N_839,In_1093);
and U1138 (N_1138,N_804,N_858);
xor U1139 (N_1139,N_406,N_689);
xnor U1140 (N_1140,N_508,N_853);
xnor U1141 (N_1141,N_903,N_894);
and U1142 (N_1142,N_714,In_325);
nand U1143 (N_1143,N_302,N_852);
xnor U1144 (N_1144,In_692,N_749);
or U1145 (N_1145,In_864,N_908);
nor U1146 (N_1146,N_756,N_822);
nand U1147 (N_1147,N_623,N_917);
or U1148 (N_1148,N_956,In_1290);
xnor U1149 (N_1149,N_568,N_188);
nor U1150 (N_1150,N_953,N_666);
nand U1151 (N_1151,N_771,N_867);
or U1152 (N_1152,N_777,N_710);
or U1153 (N_1153,In_1305,N_877);
xnor U1154 (N_1154,N_790,In_1027);
or U1155 (N_1155,N_971,N_660);
nand U1156 (N_1156,N_759,N_931);
and U1157 (N_1157,N_329,N_855);
or U1158 (N_1158,N_887,N_827);
and U1159 (N_1159,N_976,In_98);
nor U1160 (N_1160,N_841,N_823);
nand U1161 (N_1161,N_348,N_986);
xnor U1162 (N_1162,N_813,N_838);
and U1163 (N_1163,N_927,N_909);
or U1164 (N_1164,In_1442,N_974);
xor U1165 (N_1165,N_943,N_779);
or U1166 (N_1166,N_810,N_558);
and U1167 (N_1167,N_622,N_578);
nor U1168 (N_1168,In_858,N_860);
or U1169 (N_1169,N_843,N_833);
nor U1170 (N_1170,In_1297,In_1342);
xor U1171 (N_1171,In_1381,N_922);
nor U1172 (N_1172,N_933,N_990);
and U1173 (N_1173,N_528,N_991);
or U1174 (N_1174,In_1418,In_1117);
or U1175 (N_1175,N_197,In_930);
xnor U1176 (N_1176,In_122,N_902);
nor U1177 (N_1177,N_555,N_868);
nor U1178 (N_1178,N_182,N_988);
xnor U1179 (N_1179,In_1295,N_876);
nor U1180 (N_1180,N_890,N_695);
xor U1181 (N_1181,N_851,N_883);
or U1182 (N_1182,N_772,In_635);
and U1183 (N_1183,N_826,N_947);
nor U1184 (N_1184,N_610,N_885);
or U1185 (N_1185,In_1363,N_793);
nor U1186 (N_1186,In_452,In_792);
nand U1187 (N_1187,In_460,N_995);
or U1188 (N_1188,N_906,N_872);
xnor U1189 (N_1189,In_1456,N_118);
nor U1190 (N_1190,N_498,N_850);
or U1191 (N_1191,N_801,N_912);
or U1192 (N_1192,N_651,N_764);
or U1193 (N_1193,N_47,N_774);
nand U1194 (N_1194,In_34,N_746);
xor U1195 (N_1195,N_641,N_938);
nand U1196 (N_1196,N_812,N_64);
and U1197 (N_1197,In_944,N_840);
and U1198 (N_1198,N_978,N_702);
nand U1199 (N_1199,N_276,N_94);
nor U1200 (N_1200,N_834,In_561);
or U1201 (N_1201,In_1497,N_719);
or U1202 (N_1202,N_828,N_640);
nor U1203 (N_1203,N_925,In_379);
or U1204 (N_1204,In_807,N_957);
and U1205 (N_1205,N_866,N_999);
or U1206 (N_1206,N_856,N_924);
or U1207 (N_1207,N_505,N_836);
nand U1208 (N_1208,N_932,In_504);
nor U1209 (N_1209,N_830,In_476);
nor U1210 (N_1210,N_255,N_987);
xor U1211 (N_1211,N_921,N_900);
xor U1212 (N_1212,N_875,N_596);
or U1213 (N_1213,N_845,N_993);
and U1214 (N_1214,N_946,N_736);
xor U1215 (N_1215,N_896,N_296);
nor U1216 (N_1216,In_1462,In_1428);
or U1217 (N_1217,N_324,N_789);
nor U1218 (N_1218,N_624,N_748);
and U1219 (N_1219,N_551,N_133);
xnor U1220 (N_1220,N_864,N_618);
xor U1221 (N_1221,N_392,N_326);
nand U1222 (N_1222,N_151,N_90);
xnor U1223 (N_1223,N_619,N_897);
xor U1224 (N_1224,N_972,N_662);
and U1225 (N_1225,In_1183,N_929);
nand U1226 (N_1226,N_934,N_580);
nor U1227 (N_1227,N_869,N_994);
or U1228 (N_1228,In_154,N_940);
and U1229 (N_1229,N_9,N_273);
nand U1230 (N_1230,In_1299,N_785);
and U1231 (N_1231,In_935,In_189);
nor U1232 (N_1232,N_751,N_716);
or U1233 (N_1233,N_762,N_238);
or U1234 (N_1234,N_979,N_985);
and U1235 (N_1235,N_475,In_1444);
nand U1236 (N_1236,N_844,In_984);
nand U1237 (N_1237,N_647,In_1153);
xnor U1238 (N_1238,In_350,N_305);
or U1239 (N_1239,N_317,N_405);
xor U1240 (N_1240,N_817,In_25);
and U1241 (N_1241,N_784,N_959);
or U1242 (N_1242,N_447,N_952);
and U1243 (N_1243,N_738,N_63);
or U1244 (N_1244,N_602,In_1188);
xor U1245 (N_1245,N_724,In_1390);
nor U1246 (N_1246,N_847,N_404);
nor U1247 (N_1247,N_493,In_284);
and U1248 (N_1248,N_966,N_754);
xor U1249 (N_1249,N_734,N_783);
nor U1250 (N_1250,N_1184,N_1066);
nor U1251 (N_1251,N_1107,N_1018);
nand U1252 (N_1252,N_1053,N_1002);
and U1253 (N_1253,N_1167,N_1198);
or U1254 (N_1254,N_1084,N_1113);
nand U1255 (N_1255,N_1197,N_1099);
or U1256 (N_1256,N_1248,N_1009);
and U1257 (N_1257,N_1145,N_1075);
and U1258 (N_1258,N_1153,N_1191);
nor U1259 (N_1259,N_1051,N_1090);
nand U1260 (N_1260,N_1148,N_1019);
or U1261 (N_1261,N_1209,N_1242);
or U1262 (N_1262,N_1166,N_1015);
and U1263 (N_1263,N_1029,N_1213);
xnor U1264 (N_1264,N_1062,N_1149);
nand U1265 (N_1265,N_1120,N_1079);
nand U1266 (N_1266,N_1243,N_1183);
xnor U1267 (N_1267,N_1189,N_1231);
xnor U1268 (N_1268,N_1142,N_1026);
or U1269 (N_1269,N_1226,N_1080);
and U1270 (N_1270,N_1116,N_1160);
nor U1271 (N_1271,N_1196,N_1118);
xor U1272 (N_1272,N_1060,N_1049);
xor U1273 (N_1273,N_1194,N_1082);
xnor U1274 (N_1274,N_1152,N_1203);
and U1275 (N_1275,N_1176,N_1050);
or U1276 (N_1276,N_1156,N_1110);
and U1277 (N_1277,N_1058,N_1147);
xor U1278 (N_1278,N_1008,N_1232);
xor U1279 (N_1279,N_1087,N_1219);
or U1280 (N_1280,N_1144,N_1130);
xor U1281 (N_1281,N_1013,N_1020);
and U1282 (N_1282,N_1022,N_1047);
nor U1283 (N_1283,N_1127,N_1239);
xor U1284 (N_1284,N_1229,N_1109);
nand U1285 (N_1285,N_1102,N_1212);
nand U1286 (N_1286,N_1180,N_1112);
xor U1287 (N_1287,N_1223,N_1138);
xnor U1288 (N_1288,N_1055,N_1052);
and U1289 (N_1289,N_1240,N_1048);
nand U1290 (N_1290,N_1092,N_1115);
and U1291 (N_1291,N_1068,N_1201);
nand U1292 (N_1292,N_1085,N_1143);
or U1293 (N_1293,N_1067,N_1244);
nor U1294 (N_1294,N_1225,N_1161);
or U1295 (N_1295,N_1042,N_1037);
nor U1296 (N_1296,N_1216,N_1218);
nand U1297 (N_1297,N_1230,N_1033);
nor U1298 (N_1298,N_1070,N_1207);
nand U1299 (N_1299,N_1086,N_1101);
xnor U1300 (N_1300,N_1076,N_1247);
nand U1301 (N_1301,N_1124,N_1246);
or U1302 (N_1302,N_1030,N_1165);
nand U1303 (N_1303,N_1121,N_1214);
or U1304 (N_1304,N_1200,N_1117);
nand U1305 (N_1305,N_1221,N_1179);
nand U1306 (N_1306,N_1135,N_1111);
and U1307 (N_1307,N_1077,N_1036);
nand U1308 (N_1308,N_1027,N_1164);
or U1309 (N_1309,N_1175,N_1202);
nor U1310 (N_1310,N_1227,N_1151);
nand U1311 (N_1311,N_1100,N_1210);
or U1312 (N_1312,N_1224,N_1063);
nand U1313 (N_1313,N_1155,N_1106);
and U1314 (N_1314,N_1010,N_1035);
or U1315 (N_1315,N_1072,N_1083);
and U1316 (N_1316,N_1162,N_1159);
and U1317 (N_1317,N_1040,N_1056);
xor U1318 (N_1318,N_1134,N_1217);
xnor U1319 (N_1319,N_1074,N_1146);
nand U1320 (N_1320,N_1158,N_1136);
nor U1321 (N_1321,N_1094,N_1185);
xor U1322 (N_1322,N_1215,N_1054);
or U1323 (N_1323,N_1173,N_1091);
xnor U1324 (N_1324,N_1057,N_1028);
and U1325 (N_1325,N_1025,N_1133);
or U1326 (N_1326,N_1140,N_1154);
xnor U1327 (N_1327,N_1237,N_1187);
nor U1328 (N_1328,N_1193,N_1114);
or U1329 (N_1329,N_1182,N_1093);
nand U1330 (N_1330,N_1238,N_1129);
nor U1331 (N_1331,N_1192,N_1016);
nand U1332 (N_1332,N_1041,N_1178);
xnor U1333 (N_1333,N_1097,N_1123);
nand U1334 (N_1334,N_1064,N_1012);
nor U1335 (N_1335,N_1199,N_1188);
xor U1336 (N_1336,N_1032,N_1071);
nand U1337 (N_1337,N_1132,N_1017);
xnor U1338 (N_1338,N_1186,N_1069);
and U1339 (N_1339,N_1011,N_1061);
nor U1340 (N_1340,N_1001,N_1103);
and U1341 (N_1341,N_1220,N_1004);
and U1342 (N_1342,N_1021,N_1031);
nand U1343 (N_1343,N_1128,N_1007);
xor U1344 (N_1344,N_1234,N_1131);
nand U1345 (N_1345,N_1171,N_1122);
nor U1346 (N_1346,N_1190,N_1043);
xor U1347 (N_1347,N_1005,N_1038);
and U1348 (N_1348,N_1089,N_1108);
or U1349 (N_1349,N_1003,N_1044);
nor U1350 (N_1350,N_1088,N_1228);
and U1351 (N_1351,N_1039,N_1098);
nor U1352 (N_1352,N_1177,N_1233);
or U1353 (N_1353,N_1006,N_1014);
nand U1354 (N_1354,N_1024,N_1241);
xnor U1355 (N_1355,N_1150,N_1169);
nand U1356 (N_1356,N_1126,N_1170);
xnor U1357 (N_1357,N_1181,N_1125);
nor U1358 (N_1358,N_1034,N_1078);
nand U1359 (N_1359,N_1206,N_1096);
nand U1360 (N_1360,N_1023,N_1168);
xnor U1361 (N_1361,N_1174,N_1195);
xnor U1362 (N_1362,N_1205,N_1222);
and U1363 (N_1363,N_1045,N_1172);
nor U1364 (N_1364,N_1236,N_1157);
nor U1365 (N_1365,N_1065,N_1119);
and U1366 (N_1366,N_1235,N_1104);
nor U1367 (N_1367,N_1137,N_1249);
nor U1368 (N_1368,N_1139,N_1059);
nand U1369 (N_1369,N_1163,N_1000);
nand U1370 (N_1370,N_1208,N_1095);
nand U1371 (N_1371,N_1081,N_1211);
or U1372 (N_1372,N_1204,N_1046);
nand U1373 (N_1373,N_1073,N_1245);
and U1374 (N_1374,N_1141,N_1105);
nand U1375 (N_1375,N_1177,N_1234);
nor U1376 (N_1376,N_1027,N_1003);
and U1377 (N_1377,N_1142,N_1106);
and U1378 (N_1378,N_1175,N_1090);
xor U1379 (N_1379,N_1227,N_1078);
nor U1380 (N_1380,N_1247,N_1140);
or U1381 (N_1381,N_1187,N_1113);
xnor U1382 (N_1382,N_1057,N_1003);
nor U1383 (N_1383,N_1231,N_1183);
or U1384 (N_1384,N_1007,N_1226);
or U1385 (N_1385,N_1097,N_1230);
xnor U1386 (N_1386,N_1215,N_1181);
or U1387 (N_1387,N_1128,N_1214);
xnor U1388 (N_1388,N_1075,N_1058);
nand U1389 (N_1389,N_1067,N_1078);
and U1390 (N_1390,N_1011,N_1206);
nand U1391 (N_1391,N_1091,N_1015);
xor U1392 (N_1392,N_1096,N_1063);
nand U1393 (N_1393,N_1107,N_1032);
nor U1394 (N_1394,N_1241,N_1053);
nand U1395 (N_1395,N_1133,N_1231);
nand U1396 (N_1396,N_1075,N_1061);
xor U1397 (N_1397,N_1065,N_1052);
xor U1398 (N_1398,N_1068,N_1155);
and U1399 (N_1399,N_1048,N_1111);
or U1400 (N_1400,N_1108,N_1016);
xor U1401 (N_1401,N_1196,N_1163);
and U1402 (N_1402,N_1156,N_1174);
nor U1403 (N_1403,N_1176,N_1111);
nor U1404 (N_1404,N_1020,N_1068);
nand U1405 (N_1405,N_1140,N_1099);
nor U1406 (N_1406,N_1223,N_1035);
nand U1407 (N_1407,N_1051,N_1143);
xor U1408 (N_1408,N_1053,N_1071);
nand U1409 (N_1409,N_1180,N_1178);
or U1410 (N_1410,N_1105,N_1058);
nand U1411 (N_1411,N_1235,N_1046);
nand U1412 (N_1412,N_1189,N_1061);
or U1413 (N_1413,N_1242,N_1053);
or U1414 (N_1414,N_1086,N_1169);
xnor U1415 (N_1415,N_1000,N_1182);
or U1416 (N_1416,N_1061,N_1115);
nor U1417 (N_1417,N_1015,N_1142);
nand U1418 (N_1418,N_1136,N_1108);
nor U1419 (N_1419,N_1176,N_1161);
nand U1420 (N_1420,N_1230,N_1067);
nor U1421 (N_1421,N_1192,N_1190);
xnor U1422 (N_1422,N_1243,N_1086);
nor U1423 (N_1423,N_1202,N_1020);
nand U1424 (N_1424,N_1151,N_1154);
nand U1425 (N_1425,N_1068,N_1139);
xnor U1426 (N_1426,N_1052,N_1123);
xnor U1427 (N_1427,N_1087,N_1018);
xnor U1428 (N_1428,N_1122,N_1081);
and U1429 (N_1429,N_1055,N_1193);
nand U1430 (N_1430,N_1160,N_1143);
nand U1431 (N_1431,N_1178,N_1172);
nor U1432 (N_1432,N_1016,N_1180);
nand U1433 (N_1433,N_1183,N_1152);
and U1434 (N_1434,N_1145,N_1008);
xor U1435 (N_1435,N_1094,N_1106);
nand U1436 (N_1436,N_1022,N_1170);
nand U1437 (N_1437,N_1247,N_1209);
nand U1438 (N_1438,N_1150,N_1172);
xor U1439 (N_1439,N_1198,N_1207);
xnor U1440 (N_1440,N_1187,N_1148);
nand U1441 (N_1441,N_1056,N_1080);
and U1442 (N_1442,N_1208,N_1020);
nor U1443 (N_1443,N_1222,N_1195);
and U1444 (N_1444,N_1186,N_1014);
nor U1445 (N_1445,N_1195,N_1169);
xnor U1446 (N_1446,N_1139,N_1030);
and U1447 (N_1447,N_1091,N_1138);
or U1448 (N_1448,N_1019,N_1175);
nand U1449 (N_1449,N_1159,N_1196);
nor U1450 (N_1450,N_1233,N_1078);
nor U1451 (N_1451,N_1236,N_1048);
and U1452 (N_1452,N_1186,N_1115);
and U1453 (N_1453,N_1052,N_1163);
nand U1454 (N_1454,N_1130,N_1166);
xnor U1455 (N_1455,N_1138,N_1079);
nor U1456 (N_1456,N_1223,N_1068);
nand U1457 (N_1457,N_1105,N_1235);
nand U1458 (N_1458,N_1202,N_1227);
nand U1459 (N_1459,N_1061,N_1065);
nor U1460 (N_1460,N_1198,N_1074);
or U1461 (N_1461,N_1000,N_1052);
or U1462 (N_1462,N_1157,N_1107);
nor U1463 (N_1463,N_1097,N_1023);
and U1464 (N_1464,N_1193,N_1165);
nand U1465 (N_1465,N_1188,N_1034);
nand U1466 (N_1466,N_1210,N_1226);
xor U1467 (N_1467,N_1191,N_1217);
nor U1468 (N_1468,N_1030,N_1236);
and U1469 (N_1469,N_1088,N_1167);
or U1470 (N_1470,N_1160,N_1046);
and U1471 (N_1471,N_1230,N_1188);
or U1472 (N_1472,N_1145,N_1012);
nor U1473 (N_1473,N_1138,N_1028);
nand U1474 (N_1474,N_1157,N_1144);
or U1475 (N_1475,N_1204,N_1187);
xnor U1476 (N_1476,N_1241,N_1017);
xor U1477 (N_1477,N_1077,N_1091);
or U1478 (N_1478,N_1054,N_1178);
nand U1479 (N_1479,N_1146,N_1091);
or U1480 (N_1480,N_1243,N_1112);
nor U1481 (N_1481,N_1059,N_1034);
or U1482 (N_1482,N_1042,N_1228);
or U1483 (N_1483,N_1073,N_1052);
or U1484 (N_1484,N_1134,N_1202);
xor U1485 (N_1485,N_1179,N_1082);
nand U1486 (N_1486,N_1056,N_1175);
xor U1487 (N_1487,N_1130,N_1161);
or U1488 (N_1488,N_1197,N_1062);
nand U1489 (N_1489,N_1110,N_1233);
and U1490 (N_1490,N_1124,N_1146);
or U1491 (N_1491,N_1109,N_1057);
and U1492 (N_1492,N_1134,N_1098);
nor U1493 (N_1493,N_1030,N_1170);
nor U1494 (N_1494,N_1051,N_1101);
or U1495 (N_1495,N_1139,N_1119);
xnor U1496 (N_1496,N_1238,N_1038);
xor U1497 (N_1497,N_1128,N_1113);
xor U1498 (N_1498,N_1111,N_1233);
nand U1499 (N_1499,N_1215,N_1000);
nand U1500 (N_1500,N_1454,N_1336);
or U1501 (N_1501,N_1364,N_1285);
or U1502 (N_1502,N_1483,N_1282);
nand U1503 (N_1503,N_1304,N_1474);
and U1504 (N_1504,N_1398,N_1449);
and U1505 (N_1505,N_1404,N_1498);
xor U1506 (N_1506,N_1305,N_1411);
nor U1507 (N_1507,N_1452,N_1359);
xnor U1508 (N_1508,N_1340,N_1400);
or U1509 (N_1509,N_1347,N_1435);
or U1510 (N_1510,N_1280,N_1492);
xor U1511 (N_1511,N_1324,N_1490);
or U1512 (N_1512,N_1433,N_1473);
xor U1513 (N_1513,N_1393,N_1372);
or U1514 (N_1514,N_1312,N_1329);
and U1515 (N_1515,N_1466,N_1374);
xnor U1516 (N_1516,N_1300,N_1290);
nor U1517 (N_1517,N_1496,N_1289);
xor U1518 (N_1518,N_1427,N_1277);
and U1519 (N_1519,N_1258,N_1426);
xor U1520 (N_1520,N_1256,N_1379);
xnor U1521 (N_1521,N_1338,N_1399);
or U1522 (N_1522,N_1255,N_1261);
nor U1523 (N_1523,N_1457,N_1371);
nand U1524 (N_1524,N_1269,N_1472);
or U1525 (N_1525,N_1414,N_1497);
nor U1526 (N_1526,N_1327,N_1319);
or U1527 (N_1527,N_1373,N_1273);
and U1528 (N_1528,N_1302,N_1428);
and U1529 (N_1529,N_1403,N_1477);
or U1530 (N_1530,N_1395,N_1313);
xor U1531 (N_1531,N_1270,N_1360);
nand U1532 (N_1532,N_1357,N_1378);
or U1533 (N_1533,N_1476,N_1432);
and U1534 (N_1534,N_1406,N_1361);
nand U1535 (N_1535,N_1401,N_1262);
and U1536 (N_1536,N_1299,N_1341);
nand U1537 (N_1537,N_1482,N_1448);
or U1538 (N_1538,N_1303,N_1475);
nand U1539 (N_1539,N_1461,N_1423);
xnor U1540 (N_1540,N_1354,N_1293);
and U1541 (N_1541,N_1298,N_1356);
xnor U1542 (N_1542,N_1478,N_1388);
or U1543 (N_1543,N_1268,N_1418);
nand U1544 (N_1544,N_1460,N_1479);
nand U1545 (N_1545,N_1380,N_1250);
nor U1546 (N_1546,N_1253,N_1459);
nor U1547 (N_1547,N_1484,N_1387);
xor U1548 (N_1548,N_1405,N_1499);
nor U1549 (N_1549,N_1464,N_1480);
and U1550 (N_1550,N_1320,N_1470);
nand U1551 (N_1551,N_1310,N_1366);
nor U1552 (N_1552,N_1430,N_1494);
or U1553 (N_1553,N_1352,N_1389);
or U1554 (N_1554,N_1311,N_1297);
xor U1555 (N_1555,N_1381,N_1349);
nand U1556 (N_1556,N_1444,N_1487);
or U1557 (N_1557,N_1442,N_1334);
and U1558 (N_1558,N_1259,N_1316);
xor U1559 (N_1559,N_1471,N_1437);
and U1560 (N_1560,N_1429,N_1402);
nand U1561 (N_1561,N_1295,N_1391);
or U1562 (N_1562,N_1410,N_1462);
xor U1563 (N_1563,N_1485,N_1351);
nand U1564 (N_1564,N_1325,N_1332);
or U1565 (N_1565,N_1301,N_1276);
or U1566 (N_1566,N_1275,N_1467);
nor U1567 (N_1567,N_1330,N_1314);
and U1568 (N_1568,N_1443,N_1451);
and U1569 (N_1569,N_1252,N_1415);
and U1570 (N_1570,N_1416,N_1333);
xor U1571 (N_1571,N_1383,N_1363);
or U1572 (N_1572,N_1343,N_1409);
and U1573 (N_1573,N_1279,N_1390);
nor U1574 (N_1574,N_1394,N_1337);
or U1575 (N_1575,N_1315,N_1413);
nand U1576 (N_1576,N_1417,N_1450);
or U1577 (N_1577,N_1436,N_1440);
xor U1578 (N_1578,N_1488,N_1382);
or U1579 (N_1579,N_1441,N_1377);
nand U1580 (N_1580,N_1445,N_1263);
nand U1581 (N_1581,N_1264,N_1278);
and U1582 (N_1582,N_1368,N_1425);
nand U1583 (N_1583,N_1424,N_1292);
nor U1584 (N_1584,N_1254,N_1369);
or U1585 (N_1585,N_1346,N_1495);
nand U1586 (N_1586,N_1272,N_1481);
or U1587 (N_1587,N_1335,N_1358);
and U1588 (N_1588,N_1434,N_1446);
and U1589 (N_1589,N_1322,N_1260);
and U1590 (N_1590,N_1266,N_1318);
nand U1591 (N_1591,N_1339,N_1321);
or U1592 (N_1592,N_1345,N_1455);
nor U1593 (N_1593,N_1348,N_1342);
nor U1594 (N_1594,N_1365,N_1251);
nor U1595 (N_1595,N_1469,N_1422);
nand U1596 (N_1596,N_1412,N_1420);
or U1597 (N_1597,N_1308,N_1317);
nor U1598 (N_1598,N_1486,N_1326);
xnor U1599 (N_1599,N_1274,N_1362);
or U1600 (N_1600,N_1421,N_1493);
and U1601 (N_1601,N_1331,N_1294);
nand U1602 (N_1602,N_1353,N_1323);
xnor U1603 (N_1603,N_1291,N_1350);
nand U1604 (N_1604,N_1306,N_1447);
xnor U1605 (N_1605,N_1288,N_1491);
nor U1606 (N_1606,N_1463,N_1375);
and U1607 (N_1607,N_1328,N_1456);
xnor U1608 (N_1608,N_1489,N_1307);
xor U1609 (N_1609,N_1468,N_1370);
and U1610 (N_1610,N_1465,N_1344);
or U1611 (N_1611,N_1453,N_1408);
and U1612 (N_1612,N_1287,N_1257);
nor U1613 (N_1613,N_1265,N_1458);
xor U1614 (N_1614,N_1296,N_1392);
nor U1615 (N_1615,N_1286,N_1367);
and U1616 (N_1616,N_1267,N_1439);
or U1617 (N_1617,N_1407,N_1271);
and U1618 (N_1618,N_1281,N_1284);
xnor U1619 (N_1619,N_1355,N_1283);
and U1620 (N_1620,N_1376,N_1431);
nand U1621 (N_1621,N_1309,N_1385);
nor U1622 (N_1622,N_1419,N_1396);
nor U1623 (N_1623,N_1438,N_1397);
nor U1624 (N_1624,N_1386,N_1384);
or U1625 (N_1625,N_1367,N_1391);
or U1626 (N_1626,N_1383,N_1391);
nor U1627 (N_1627,N_1462,N_1323);
nand U1628 (N_1628,N_1389,N_1438);
nand U1629 (N_1629,N_1309,N_1269);
nor U1630 (N_1630,N_1413,N_1394);
nand U1631 (N_1631,N_1290,N_1402);
nor U1632 (N_1632,N_1317,N_1357);
xor U1633 (N_1633,N_1434,N_1453);
nor U1634 (N_1634,N_1302,N_1405);
xor U1635 (N_1635,N_1409,N_1411);
and U1636 (N_1636,N_1419,N_1494);
or U1637 (N_1637,N_1377,N_1316);
nor U1638 (N_1638,N_1272,N_1367);
or U1639 (N_1639,N_1348,N_1458);
nor U1640 (N_1640,N_1442,N_1341);
and U1641 (N_1641,N_1484,N_1256);
nor U1642 (N_1642,N_1254,N_1402);
xor U1643 (N_1643,N_1315,N_1340);
nand U1644 (N_1644,N_1420,N_1363);
or U1645 (N_1645,N_1454,N_1459);
nor U1646 (N_1646,N_1371,N_1330);
nand U1647 (N_1647,N_1326,N_1400);
xor U1648 (N_1648,N_1320,N_1362);
nand U1649 (N_1649,N_1252,N_1257);
and U1650 (N_1650,N_1392,N_1280);
and U1651 (N_1651,N_1398,N_1416);
and U1652 (N_1652,N_1319,N_1361);
and U1653 (N_1653,N_1373,N_1266);
nor U1654 (N_1654,N_1432,N_1356);
nand U1655 (N_1655,N_1424,N_1253);
nor U1656 (N_1656,N_1303,N_1456);
or U1657 (N_1657,N_1462,N_1492);
and U1658 (N_1658,N_1399,N_1257);
xnor U1659 (N_1659,N_1391,N_1342);
xnor U1660 (N_1660,N_1462,N_1494);
and U1661 (N_1661,N_1427,N_1256);
and U1662 (N_1662,N_1364,N_1289);
and U1663 (N_1663,N_1428,N_1474);
nor U1664 (N_1664,N_1313,N_1325);
nand U1665 (N_1665,N_1306,N_1427);
xor U1666 (N_1666,N_1422,N_1347);
or U1667 (N_1667,N_1484,N_1349);
xor U1668 (N_1668,N_1361,N_1322);
xor U1669 (N_1669,N_1461,N_1367);
or U1670 (N_1670,N_1371,N_1346);
or U1671 (N_1671,N_1480,N_1445);
xnor U1672 (N_1672,N_1267,N_1358);
nor U1673 (N_1673,N_1282,N_1462);
nand U1674 (N_1674,N_1313,N_1480);
xnor U1675 (N_1675,N_1494,N_1424);
and U1676 (N_1676,N_1310,N_1412);
xor U1677 (N_1677,N_1309,N_1460);
nor U1678 (N_1678,N_1451,N_1404);
and U1679 (N_1679,N_1341,N_1392);
nor U1680 (N_1680,N_1414,N_1345);
nand U1681 (N_1681,N_1324,N_1381);
and U1682 (N_1682,N_1325,N_1475);
nand U1683 (N_1683,N_1436,N_1474);
nand U1684 (N_1684,N_1270,N_1323);
nor U1685 (N_1685,N_1494,N_1348);
nor U1686 (N_1686,N_1480,N_1470);
and U1687 (N_1687,N_1251,N_1340);
xor U1688 (N_1688,N_1447,N_1465);
and U1689 (N_1689,N_1492,N_1366);
or U1690 (N_1690,N_1374,N_1339);
nand U1691 (N_1691,N_1303,N_1263);
nor U1692 (N_1692,N_1417,N_1303);
nand U1693 (N_1693,N_1473,N_1314);
or U1694 (N_1694,N_1271,N_1263);
nor U1695 (N_1695,N_1397,N_1313);
or U1696 (N_1696,N_1495,N_1460);
nor U1697 (N_1697,N_1403,N_1447);
or U1698 (N_1698,N_1396,N_1331);
xnor U1699 (N_1699,N_1292,N_1465);
nand U1700 (N_1700,N_1380,N_1362);
or U1701 (N_1701,N_1381,N_1435);
and U1702 (N_1702,N_1443,N_1309);
nor U1703 (N_1703,N_1355,N_1335);
xnor U1704 (N_1704,N_1329,N_1379);
xor U1705 (N_1705,N_1417,N_1340);
nand U1706 (N_1706,N_1335,N_1445);
nor U1707 (N_1707,N_1482,N_1260);
nand U1708 (N_1708,N_1406,N_1262);
nand U1709 (N_1709,N_1266,N_1299);
xnor U1710 (N_1710,N_1383,N_1392);
nand U1711 (N_1711,N_1466,N_1416);
nand U1712 (N_1712,N_1477,N_1414);
or U1713 (N_1713,N_1270,N_1462);
xnor U1714 (N_1714,N_1475,N_1406);
xor U1715 (N_1715,N_1284,N_1489);
nand U1716 (N_1716,N_1252,N_1301);
or U1717 (N_1717,N_1383,N_1439);
xnor U1718 (N_1718,N_1472,N_1323);
nor U1719 (N_1719,N_1419,N_1409);
or U1720 (N_1720,N_1252,N_1336);
nor U1721 (N_1721,N_1498,N_1315);
nor U1722 (N_1722,N_1256,N_1294);
and U1723 (N_1723,N_1334,N_1489);
xnor U1724 (N_1724,N_1290,N_1413);
and U1725 (N_1725,N_1397,N_1333);
nand U1726 (N_1726,N_1489,N_1291);
and U1727 (N_1727,N_1495,N_1330);
xnor U1728 (N_1728,N_1455,N_1271);
nor U1729 (N_1729,N_1370,N_1338);
nand U1730 (N_1730,N_1341,N_1262);
or U1731 (N_1731,N_1387,N_1491);
nor U1732 (N_1732,N_1366,N_1499);
nand U1733 (N_1733,N_1289,N_1480);
nand U1734 (N_1734,N_1293,N_1358);
and U1735 (N_1735,N_1457,N_1309);
nor U1736 (N_1736,N_1274,N_1264);
nand U1737 (N_1737,N_1315,N_1454);
nand U1738 (N_1738,N_1324,N_1481);
and U1739 (N_1739,N_1383,N_1346);
and U1740 (N_1740,N_1392,N_1344);
or U1741 (N_1741,N_1397,N_1469);
xnor U1742 (N_1742,N_1262,N_1431);
and U1743 (N_1743,N_1492,N_1472);
nand U1744 (N_1744,N_1417,N_1462);
nor U1745 (N_1745,N_1458,N_1374);
and U1746 (N_1746,N_1434,N_1360);
xor U1747 (N_1747,N_1294,N_1363);
nor U1748 (N_1748,N_1466,N_1446);
and U1749 (N_1749,N_1395,N_1296);
nor U1750 (N_1750,N_1572,N_1505);
and U1751 (N_1751,N_1624,N_1668);
nand U1752 (N_1752,N_1545,N_1503);
nand U1753 (N_1753,N_1663,N_1507);
nand U1754 (N_1754,N_1592,N_1719);
xnor U1755 (N_1755,N_1565,N_1675);
xor U1756 (N_1756,N_1538,N_1659);
nor U1757 (N_1757,N_1611,N_1744);
and U1758 (N_1758,N_1510,N_1656);
nand U1759 (N_1759,N_1740,N_1693);
xor U1760 (N_1760,N_1513,N_1734);
or U1761 (N_1761,N_1534,N_1588);
or U1762 (N_1762,N_1688,N_1543);
nor U1763 (N_1763,N_1702,N_1612);
and U1764 (N_1764,N_1748,N_1524);
and U1765 (N_1765,N_1680,N_1587);
nand U1766 (N_1766,N_1536,N_1615);
nor U1767 (N_1767,N_1699,N_1729);
nand U1768 (N_1768,N_1716,N_1626);
nor U1769 (N_1769,N_1730,N_1523);
nand U1770 (N_1770,N_1749,N_1664);
nand U1771 (N_1771,N_1589,N_1614);
nor U1772 (N_1772,N_1689,N_1720);
nor U1773 (N_1773,N_1636,N_1590);
nor U1774 (N_1774,N_1700,N_1617);
or U1775 (N_1775,N_1576,N_1629);
xor U1776 (N_1776,N_1738,N_1618);
nor U1777 (N_1777,N_1666,N_1672);
and U1778 (N_1778,N_1613,N_1676);
nand U1779 (N_1779,N_1745,N_1637);
and U1780 (N_1780,N_1569,N_1527);
or U1781 (N_1781,N_1564,N_1597);
xnor U1782 (N_1782,N_1646,N_1623);
nor U1783 (N_1783,N_1573,N_1562);
or U1784 (N_1784,N_1639,N_1712);
xor U1785 (N_1785,N_1655,N_1667);
xnor U1786 (N_1786,N_1652,N_1514);
and U1787 (N_1787,N_1728,N_1657);
or U1788 (N_1788,N_1661,N_1743);
nor U1789 (N_1789,N_1705,N_1724);
nor U1790 (N_1790,N_1580,N_1746);
and U1791 (N_1791,N_1677,N_1581);
and U1792 (N_1792,N_1521,N_1665);
xnor U1793 (N_1793,N_1701,N_1698);
xor U1794 (N_1794,N_1598,N_1602);
or U1795 (N_1795,N_1708,N_1604);
nand U1796 (N_1796,N_1658,N_1501);
nor U1797 (N_1797,N_1500,N_1731);
nor U1798 (N_1798,N_1540,N_1625);
and U1799 (N_1799,N_1508,N_1509);
and U1800 (N_1800,N_1567,N_1556);
or U1801 (N_1801,N_1577,N_1605);
or U1802 (N_1802,N_1711,N_1547);
xnor U1803 (N_1803,N_1696,N_1603);
nor U1804 (N_1804,N_1586,N_1558);
or U1805 (N_1805,N_1541,N_1707);
nor U1806 (N_1806,N_1528,N_1529);
nor U1807 (N_1807,N_1742,N_1694);
nand U1808 (N_1808,N_1643,N_1504);
xnor U1809 (N_1809,N_1518,N_1713);
nor U1810 (N_1810,N_1531,N_1560);
nor U1811 (N_1811,N_1517,N_1553);
and U1812 (N_1812,N_1566,N_1662);
or U1813 (N_1813,N_1593,N_1721);
and U1814 (N_1814,N_1578,N_1522);
xor U1815 (N_1815,N_1715,N_1649);
and U1816 (N_1816,N_1609,N_1579);
or U1817 (N_1817,N_1570,N_1640);
and U1818 (N_1818,N_1679,N_1549);
nor U1819 (N_1819,N_1559,N_1684);
xnor U1820 (N_1820,N_1733,N_1519);
or U1821 (N_1821,N_1634,N_1747);
or U1822 (N_1822,N_1678,N_1606);
or U1823 (N_1823,N_1648,N_1551);
nor U1824 (N_1824,N_1526,N_1601);
nor U1825 (N_1825,N_1622,N_1520);
nand U1826 (N_1826,N_1555,N_1627);
nand U1827 (N_1827,N_1539,N_1717);
and U1828 (N_1828,N_1544,N_1722);
nand U1829 (N_1829,N_1718,N_1608);
xor U1830 (N_1830,N_1511,N_1714);
nand U1831 (N_1831,N_1591,N_1709);
nand U1832 (N_1832,N_1619,N_1727);
or U1833 (N_1833,N_1735,N_1635);
nor U1834 (N_1834,N_1532,N_1568);
nor U1835 (N_1835,N_1561,N_1736);
and U1836 (N_1836,N_1732,N_1692);
xor U1837 (N_1837,N_1681,N_1506);
or U1838 (N_1838,N_1633,N_1645);
nor U1839 (N_1839,N_1620,N_1660);
xnor U1840 (N_1840,N_1641,N_1584);
nand U1841 (N_1841,N_1653,N_1552);
and U1842 (N_1842,N_1631,N_1574);
nand U1843 (N_1843,N_1695,N_1704);
and U1844 (N_1844,N_1616,N_1703);
nor U1845 (N_1845,N_1670,N_1548);
or U1846 (N_1846,N_1739,N_1630);
and U1847 (N_1847,N_1638,N_1687);
and U1848 (N_1848,N_1542,N_1582);
and U1849 (N_1849,N_1595,N_1690);
nor U1850 (N_1850,N_1632,N_1697);
nand U1851 (N_1851,N_1583,N_1644);
nand U1852 (N_1852,N_1533,N_1686);
nand U1853 (N_1853,N_1671,N_1651);
and U1854 (N_1854,N_1557,N_1585);
nand U1855 (N_1855,N_1600,N_1530);
nor U1856 (N_1856,N_1682,N_1726);
nand U1857 (N_1857,N_1537,N_1647);
nand U1858 (N_1858,N_1710,N_1725);
and U1859 (N_1859,N_1628,N_1512);
xor U1860 (N_1860,N_1594,N_1571);
and U1861 (N_1861,N_1691,N_1596);
or U1862 (N_1862,N_1741,N_1706);
xor U1863 (N_1863,N_1535,N_1610);
or U1864 (N_1864,N_1607,N_1516);
nand U1865 (N_1865,N_1515,N_1673);
or U1866 (N_1866,N_1674,N_1546);
xnor U1867 (N_1867,N_1550,N_1525);
nand U1868 (N_1868,N_1502,N_1683);
xnor U1869 (N_1869,N_1654,N_1669);
and U1870 (N_1870,N_1563,N_1554);
xor U1871 (N_1871,N_1723,N_1621);
xnor U1872 (N_1872,N_1737,N_1642);
xnor U1873 (N_1873,N_1685,N_1599);
or U1874 (N_1874,N_1650,N_1575);
and U1875 (N_1875,N_1530,N_1701);
xnor U1876 (N_1876,N_1693,N_1670);
or U1877 (N_1877,N_1575,N_1519);
or U1878 (N_1878,N_1603,N_1699);
xor U1879 (N_1879,N_1681,N_1523);
nand U1880 (N_1880,N_1505,N_1622);
nand U1881 (N_1881,N_1630,N_1565);
nand U1882 (N_1882,N_1637,N_1668);
xnor U1883 (N_1883,N_1578,N_1625);
nor U1884 (N_1884,N_1714,N_1575);
nand U1885 (N_1885,N_1609,N_1605);
and U1886 (N_1886,N_1744,N_1621);
or U1887 (N_1887,N_1612,N_1508);
or U1888 (N_1888,N_1535,N_1722);
or U1889 (N_1889,N_1536,N_1594);
nor U1890 (N_1890,N_1528,N_1678);
nand U1891 (N_1891,N_1677,N_1565);
nand U1892 (N_1892,N_1641,N_1676);
nor U1893 (N_1893,N_1741,N_1586);
nand U1894 (N_1894,N_1663,N_1670);
and U1895 (N_1895,N_1574,N_1616);
and U1896 (N_1896,N_1509,N_1528);
and U1897 (N_1897,N_1608,N_1686);
and U1898 (N_1898,N_1726,N_1549);
xnor U1899 (N_1899,N_1559,N_1585);
or U1900 (N_1900,N_1622,N_1531);
and U1901 (N_1901,N_1521,N_1540);
xnor U1902 (N_1902,N_1509,N_1668);
and U1903 (N_1903,N_1682,N_1713);
nor U1904 (N_1904,N_1596,N_1699);
xor U1905 (N_1905,N_1543,N_1728);
or U1906 (N_1906,N_1507,N_1530);
xor U1907 (N_1907,N_1545,N_1700);
nand U1908 (N_1908,N_1661,N_1703);
nor U1909 (N_1909,N_1539,N_1532);
or U1910 (N_1910,N_1685,N_1592);
nand U1911 (N_1911,N_1502,N_1664);
or U1912 (N_1912,N_1500,N_1642);
nand U1913 (N_1913,N_1519,N_1508);
nand U1914 (N_1914,N_1550,N_1744);
nor U1915 (N_1915,N_1529,N_1735);
and U1916 (N_1916,N_1508,N_1672);
and U1917 (N_1917,N_1668,N_1576);
xor U1918 (N_1918,N_1703,N_1554);
or U1919 (N_1919,N_1686,N_1621);
or U1920 (N_1920,N_1711,N_1632);
nand U1921 (N_1921,N_1662,N_1522);
nor U1922 (N_1922,N_1614,N_1644);
and U1923 (N_1923,N_1541,N_1571);
and U1924 (N_1924,N_1665,N_1684);
nand U1925 (N_1925,N_1530,N_1516);
and U1926 (N_1926,N_1507,N_1635);
nand U1927 (N_1927,N_1629,N_1526);
nor U1928 (N_1928,N_1580,N_1670);
or U1929 (N_1929,N_1686,N_1703);
nand U1930 (N_1930,N_1712,N_1674);
nor U1931 (N_1931,N_1684,N_1568);
and U1932 (N_1932,N_1559,N_1647);
or U1933 (N_1933,N_1516,N_1604);
nand U1934 (N_1934,N_1738,N_1598);
xnor U1935 (N_1935,N_1513,N_1622);
nor U1936 (N_1936,N_1564,N_1701);
nand U1937 (N_1937,N_1627,N_1518);
nand U1938 (N_1938,N_1685,N_1533);
or U1939 (N_1939,N_1538,N_1545);
and U1940 (N_1940,N_1541,N_1629);
nor U1941 (N_1941,N_1621,N_1623);
and U1942 (N_1942,N_1713,N_1616);
xor U1943 (N_1943,N_1656,N_1559);
nand U1944 (N_1944,N_1584,N_1636);
and U1945 (N_1945,N_1735,N_1673);
xor U1946 (N_1946,N_1735,N_1570);
nor U1947 (N_1947,N_1727,N_1657);
or U1948 (N_1948,N_1706,N_1584);
nor U1949 (N_1949,N_1713,N_1681);
nor U1950 (N_1950,N_1656,N_1518);
nor U1951 (N_1951,N_1649,N_1588);
or U1952 (N_1952,N_1613,N_1580);
xnor U1953 (N_1953,N_1682,N_1502);
nor U1954 (N_1954,N_1541,N_1640);
nor U1955 (N_1955,N_1732,N_1574);
or U1956 (N_1956,N_1581,N_1683);
nand U1957 (N_1957,N_1535,N_1502);
or U1958 (N_1958,N_1527,N_1502);
and U1959 (N_1959,N_1701,N_1651);
or U1960 (N_1960,N_1637,N_1537);
and U1961 (N_1961,N_1582,N_1659);
nand U1962 (N_1962,N_1590,N_1645);
xnor U1963 (N_1963,N_1680,N_1720);
or U1964 (N_1964,N_1523,N_1684);
or U1965 (N_1965,N_1530,N_1606);
nand U1966 (N_1966,N_1716,N_1583);
xor U1967 (N_1967,N_1702,N_1513);
and U1968 (N_1968,N_1694,N_1631);
and U1969 (N_1969,N_1718,N_1586);
nor U1970 (N_1970,N_1689,N_1611);
or U1971 (N_1971,N_1643,N_1721);
nor U1972 (N_1972,N_1697,N_1661);
or U1973 (N_1973,N_1647,N_1673);
nor U1974 (N_1974,N_1687,N_1572);
or U1975 (N_1975,N_1504,N_1554);
xor U1976 (N_1976,N_1525,N_1543);
nor U1977 (N_1977,N_1555,N_1610);
and U1978 (N_1978,N_1729,N_1563);
nor U1979 (N_1979,N_1667,N_1729);
xnor U1980 (N_1980,N_1606,N_1566);
or U1981 (N_1981,N_1616,N_1626);
or U1982 (N_1982,N_1685,N_1613);
and U1983 (N_1983,N_1526,N_1588);
xnor U1984 (N_1984,N_1723,N_1517);
xor U1985 (N_1985,N_1652,N_1698);
nor U1986 (N_1986,N_1578,N_1574);
xnor U1987 (N_1987,N_1717,N_1575);
or U1988 (N_1988,N_1737,N_1618);
or U1989 (N_1989,N_1632,N_1644);
nor U1990 (N_1990,N_1504,N_1609);
or U1991 (N_1991,N_1599,N_1579);
xnor U1992 (N_1992,N_1537,N_1564);
nor U1993 (N_1993,N_1712,N_1534);
nor U1994 (N_1994,N_1587,N_1562);
and U1995 (N_1995,N_1715,N_1741);
nor U1996 (N_1996,N_1695,N_1667);
nand U1997 (N_1997,N_1557,N_1668);
and U1998 (N_1998,N_1670,N_1531);
xor U1999 (N_1999,N_1736,N_1678);
or U2000 (N_2000,N_1950,N_1817);
xnor U2001 (N_2001,N_1947,N_1932);
xor U2002 (N_2002,N_1989,N_1752);
or U2003 (N_2003,N_1956,N_1972);
nor U2004 (N_2004,N_1814,N_1974);
or U2005 (N_2005,N_1751,N_1949);
xnor U2006 (N_2006,N_1962,N_1866);
nor U2007 (N_2007,N_1875,N_1939);
or U2008 (N_2008,N_1801,N_1973);
nand U2009 (N_2009,N_1919,N_1755);
nand U2010 (N_2010,N_1969,N_1887);
nand U2011 (N_2011,N_1933,N_1807);
or U2012 (N_2012,N_1916,N_1978);
xnor U2013 (N_2013,N_1941,N_1851);
nor U2014 (N_2014,N_1929,N_1859);
nand U2015 (N_2015,N_1821,N_1874);
or U2016 (N_2016,N_1832,N_1824);
or U2017 (N_2017,N_1831,N_1786);
xnor U2018 (N_2018,N_1912,N_1990);
or U2019 (N_2019,N_1775,N_1849);
and U2020 (N_2020,N_1971,N_1861);
or U2021 (N_2021,N_1762,N_1881);
nor U2022 (N_2022,N_1797,N_1837);
nand U2023 (N_2023,N_1901,N_1776);
nand U2024 (N_2024,N_1938,N_1810);
nor U2025 (N_2025,N_1795,N_1966);
or U2026 (N_2026,N_1799,N_1967);
and U2027 (N_2027,N_1769,N_1753);
and U2028 (N_2028,N_1785,N_1910);
or U2029 (N_2029,N_1825,N_1899);
or U2030 (N_2030,N_1854,N_1925);
xnor U2031 (N_2031,N_1986,N_1920);
xnor U2032 (N_2032,N_1922,N_1889);
and U2033 (N_2033,N_1853,N_1763);
or U2034 (N_2034,N_1987,N_1835);
nor U2035 (N_2035,N_1894,N_1789);
nor U2036 (N_2036,N_1777,N_1819);
nor U2037 (N_2037,N_1771,N_1946);
nor U2038 (N_2038,N_1888,N_1766);
and U2039 (N_2039,N_1984,N_1996);
xor U2040 (N_2040,N_1848,N_1794);
nand U2041 (N_2041,N_1995,N_1897);
xor U2042 (N_2042,N_1815,N_1906);
or U2043 (N_2043,N_1796,N_1780);
xor U2044 (N_2044,N_1924,N_1997);
nand U2045 (N_2045,N_1768,N_1940);
nand U2046 (N_2046,N_1855,N_1908);
nand U2047 (N_2047,N_1860,N_1781);
and U2048 (N_2048,N_1890,N_1830);
or U2049 (N_2049,N_1847,N_1968);
xnor U2050 (N_2050,N_1970,N_1823);
xor U2051 (N_2051,N_1943,N_1878);
or U2052 (N_2052,N_1958,N_1806);
nand U2053 (N_2053,N_1877,N_1857);
xnor U2054 (N_2054,N_1809,N_1951);
nand U2055 (N_2055,N_1783,N_1761);
nor U2056 (N_2056,N_1800,N_1862);
xnor U2057 (N_2057,N_1994,N_1820);
xor U2058 (N_2058,N_1979,N_1900);
nand U2059 (N_2059,N_1905,N_1952);
or U2060 (N_2060,N_1765,N_1954);
nor U2061 (N_2061,N_1921,N_1965);
xor U2062 (N_2062,N_1915,N_1788);
xnor U2063 (N_2063,N_1991,N_1834);
nor U2064 (N_2064,N_1867,N_1988);
xnor U2065 (N_2065,N_1829,N_1879);
and U2066 (N_2066,N_1914,N_1770);
nor U2067 (N_2067,N_1864,N_1784);
xnor U2068 (N_2068,N_1975,N_1931);
nor U2069 (N_2069,N_1833,N_1778);
and U2070 (N_2070,N_1870,N_1816);
nor U2071 (N_2071,N_1883,N_1805);
xor U2072 (N_2072,N_1793,N_1827);
or U2073 (N_2073,N_1982,N_1934);
nand U2074 (N_2074,N_1959,N_1773);
xor U2075 (N_2075,N_1981,N_1955);
or U2076 (N_2076,N_1907,N_1893);
xor U2077 (N_2077,N_1911,N_1798);
xor U2078 (N_2078,N_1872,N_1953);
xor U2079 (N_2079,N_1977,N_1868);
and U2080 (N_2080,N_1803,N_1896);
nand U2081 (N_2081,N_1826,N_1985);
or U2082 (N_2082,N_1756,N_1964);
nor U2083 (N_2083,N_1948,N_1892);
or U2084 (N_2084,N_1873,N_1863);
nand U2085 (N_2085,N_1790,N_1757);
xnor U2086 (N_2086,N_1992,N_1936);
nor U2087 (N_2087,N_1802,N_1865);
or U2088 (N_2088,N_1998,N_1818);
xor U2089 (N_2089,N_1840,N_1836);
nor U2090 (N_2090,N_1882,N_1942);
xnor U2091 (N_2091,N_1850,N_1945);
xnor U2092 (N_2092,N_1845,N_1852);
and U2093 (N_2093,N_1963,N_1880);
or U2094 (N_2094,N_1792,N_1759);
xor U2095 (N_2095,N_1844,N_1774);
nor U2096 (N_2096,N_1944,N_1779);
or U2097 (N_2097,N_1884,N_1976);
and U2098 (N_2098,N_1927,N_1937);
xnor U2099 (N_2099,N_1895,N_1917);
nand U2100 (N_2100,N_1904,N_1760);
and U2101 (N_2101,N_1935,N_1750);
nand U2102 (N_2102,N_1842,N_1903);
and U2103 (N_2103,N_1960,N_1886);
or U2104 (N_2104,N_1838,N_1983);
xnor U2105 (N_2105,N_1869,N_1913);
nand U2106 (N_2106,N_1928,N_1841);
nor U2107 (N_2107,N_1891,N_1764);
and U2108 (N_2108,N_1957,N_1858);
or U2109 (N_2109,N_1754,N_1839);
xor U2110 (N_2110,N_1999,N_1787);
nor U2111 (N_2111,N_1930,N_1811);
xnor U2112 (N_2112,N_1876,N_1923);
nor U2113 (N_2113,N_1980,N_1804);
and U2114 (N_2114,N_1813,N_1909);
and U2115 (N_2115,N_1782,N_1767);
xor U2116 (N_2116,N_1843,N_1926);
xor U2117 (N_2117,N_1993,N_1885);
nor U2118 (N_2118,N_1871,N_1846);
nor U2119 (N_2119,N_1808,N_1961);
and U2120 (N_2120,N_1772,N_1791);
nor U2121 (N_2121,N_1856,N_1918);
nand U2122 (N_2122,N_1898,N_1828);
and U2123 (N_2123,N_1758,N_1902);
nor U2124 (N_2124,N_1812,N_1822);
xnor U2125 (N_2125,N_1774,N_1958);
nor U2126 (N_2126,N_1879,N_1954);
nor U2127 (N_2127,N_1825,N_1911);
nand U2128 (N_2128,N_1815,N_1845);
nor U2129 (N_2129,N_1786,N_1979);
nor U2130 (N_2130,N_1899,N_1955);
nand U2131 (N_2131,N_1882,N_1858);
and U2132 (N_2132,N_1888,N_1976);
xor U2133 (N_2133,N_1992,N_1966);
or U2134 (N_2134,N_1813,N_1892);
nor U2135 (N_2135,N_1933,N_1766);
or U2136 (N_2136,N_1969,N_1783);
nand U2137 (N_2137,N_1969,N_1758);
nand U2138 (N_2138,N_1861,N_1926);
nand U2139 (N_2139,N_1755,N_1834);
xnor U2140 (N_2140,N_1791,N_1944);
nor U2141 (N_2141,N_1972,N_1887);
xor U2142 (N_2142,N_1888,N_1918);
or U2143 (N_2143,N_1753,N_1952);
nand U2144 (N_2144,N_1942,N_1814);
and U2145 (N_2145,N_1884,N_1870);
or U2146 (N_2146,N_1825,N_1999);
nor U2147 (N_2147,N_1940,N_1888);
and U2148 (N_2148,N_1902,N_1933);
and U2149 (N_2149,N_1993,N_1962);
xnor U2150 (N_2150,N_1937,N_1824);
xnor U2151 (N_2151,N_1784,N_1818);
and U2152 (N_2152,N_1993,N_1783);
and U2153 (N_2153,N_1759,N_1814);
or U2154 (N_2154,N_1793,N_1771);
nand U2155 (N_2155,N_1786,N_1811);
nand U2156 (N_2156,N_1967,N_1792);
and U2157 (N_2157,N_1914,N_1850);
and U2158 (N_2158,N_1936,N_1851);
or U2159 (N_2159,N_1790,N_1964);
nand U2160 (N_2160,N_1810,N_1785);
and U2161 (N_2161,N_1845,N_1977);
and U2162 (N_2162,N_1976,N_1974);
or U2163 (N_2163,N_1951,N_1926);
nand U2164 (N_2164,N_1788,N_1822);
nor U2165 (N_2165,N_1931,N_1824);
nor U2166 (N_2166,N_1834,N_1899);
nand U2167 (N_2167,N_1849,N_1931);
nor U2168 (N_2168,N_1932,N_1921);
or U2169 (N_2169,N_1764,N_1890);
xor U2170 (N_2170,N_1927,N_1841);
and U2171 (N_2171,N_1992,N_1881);
or U2172 (N_2172,N_1789,N_1949);
nor U2173 (N_2173,N_1830,N_1939);
and U2174 (N_2174,N_1833,N_1765);
or U2175 (N_2175,N_1983,N_1754);
or U2176 (N_2176,N_1918,N_1928);
xnor U2177 (N_2177,N_1799,N_1876);
and U2178 (N_2178,N_1780,N_1828);
nand U2179 (N_2179,N_1952,N_1767);
nor U2180 (N_2180,N_1850,N_1889);
xnor U2181 (N_2181,N_1985,N_1863);
nor U2182 (N_2182,N_1839,N_1877);
nand U2183 (N_2183,N_1965,N_1814);
or U2184 (N_2184,N_1777,N_1973);
nor U2185 (N_2185,N_1960,N_1829);
or U2186 (N_2186,N_1861,N_1773);
and U2187 (N_2187,N_1989,N_1905);
nand U2188 (N_2188,N_1836,N_1818);
nor U2189 (N_2189,N_1774,N_1868);
or U2190 (N_2190,N_1871,N_1855);
or U2191 (N_2191,N_1892,N_1861);
nor U2192 (N_2192,N_1966,N_1791);
or U2193 (N_2193,N_1809,N_1912);
nand U2194 (N_2194,N_1983,N_1993);
or U2195 (N_2195,N_1860,N_1919);
nand U2196 (N_2196,N_1843,N_1941);
nand U2197 (N_2197,N_1890,N_1973);
and U2198 (N_2198,N_1751,N_1764);
and U2199 (N_2199,N_1792,N_1770);
nand U2200 (N_2200,N_1926,N_1974);
nand U2201 (N_2201,N_1871,N_1864);
or U2202 (N_2202,N_1883,N_1872);
nor U2203 (N_2203,N_1986,N_1784);
and U2204 (N_2204,N_1931,N_1983);
xnor U2205 (N_2205,N_1963,N_1969);
and U2206 (N_2206,N_1996,N_1910);
nand U2207 (N_2207,N_1873,N_1868);
and U2208 (N_2208,N_1899,N_1812);
nor U2209 (N_2209,N_1956,N_1755);
nor U2210 (N_2210,N_1844,N_1880);
nand U2211 (N_2211,N_1816,N_1974);
or U2212 (N_2212,N_1922,N_1880);
xor U2213 (N_2213,N_1777,N_1976);
nor U2214 (N_2214,N_1894,N_1916);
xor U2215 (N_2215,N_1974,N_1850);
or U2216 (N_2216,N_1895,N_1956);
xnor U2217 (N_2217,N_1994,N_1892);
and U2218 (N_2218,N_1975,N_1980);
nand U2219 (N_2219,N_1998,N_1864);
xnor U2220 (N_2220,N_1912,N_1996);
xor U2221 (N_2221,N_1922,N_1850);
xnor U2222 (N_2222,N_1842,N_1777);
nor U2223 (N_2223,N_1941,N_1899);
nand U2224 (N_2224,N_1858,N_1972);
or U2225 (N_2225,N_1785,N_1819);
or U2226 (N_2226,N_1833,N_1771);
or U2227 (N_2227,N_1995,N_1955);
or U2228 (N_2228,N_1892,N_1755);
and U2229 (N_2229,N_1995,N_1799);
nand U2230 (N_2230,N_1757,N_1880);
or U2231 (N_2231,N_1878,N_1975);
nand U2232 (N_2232,N_1758,N_1943);
nor U2233 (N_2233,N_1835,N_1758);
xor U2234 (N_2234,N_1854,N_1915);
and U2235 (N_2235,N_1817,N_1837);
xor U2236 (N_2236,N_1787,N_1832);
nor U2237 (N_2237,N_1799,N_1774);
xnor U2238 (N_2238,N_1784,N_1774);
nand U2239 (N_2239,N_1755,N_1912);
or U2240 (N_2240,N_1922,N_1943);
and U2241 (N_2241,N_1976,N_1950);
or U2242 (N_2242,N_1774,N_1750);
nand U2243 (N_2243,N_1850,N_1983);
nand U2244 (N_2244,N_1787,N_1810);
nand U2245 (N_2245,N_1779,N_1884);
or U2246 (N_2246,N_1787,N_1797);
and U2247 (N_2247,N_1820,N_1751);
and U2248 (N_2248,N_1766,N_1850);
xor U2249 (N_2249,N_1906,N_1820);
xor U2250 (N_2250,N_2018,N_2016);
and U2251 (N_2251,N_2216,N_2012);
or U2252 (N_2252,N_2112,N_2059);
and U2253 (N_2253,N_2143,N_2239);
nor U2254 (N_2254,N_2064,N_2214);
xnor U2255 (N_2255,N_2120,N_2185);
nor U2256 (N_2256,N_2087,N_2027);
xor U2257 (N_2257,N_2128,N_2060);
or U2258 (N_2258,N_2031,N_2209);
and U2259 (N_2259,N_2138,N_2080);
nand U2260 (N_2260,N_2084,N_2189);
or U2261 (N_2261,N_2061,N_2040);
or U2262 (N_2262,N_2184,N_2142);
or U2263 (N_2263,N_2045,N_2034);
xnor U2264 (N_2264,N_2062,N_2009);
or U2265 (N_2265,N_2025,N_2033);
or U2266 (N_2266,N_2134,N_2162);
or U2267 (N_2267,N_2075,N_2237);
nor U2268 (N_2268,N_2160,N_2053);
or U2269 (N_2269,N_2085,N_2020);
nor U2270 (N_2270,N_2213,N_2171);
nor U2271 (N_2271,N_2065,N_2072);
or U2272 (N_2272,N_2179,N_2182);
and U2273 (N_2273,N_2131,N_2124);
and U2274 (N_2274,N_2243,N_2021);
nor U2275 (N_2275,N_2206,N_2028);
xor U2276 (N_2276,N_2105,N_2132);
or U2277 (N_2277,N_2156,N_2043);
nor U2278 (N_2278,N_2229,N_2133);
and U2279 (N_2279,N_2161,N_2153);
or U2280 (N_2280,N_2205,N_2234);
and U2281 (N_2281,N_2078,N_2198);
and U2282 (N_2282,N_2057,N_2249);
xnor U2283 (N_2283,N_2026,N_2041);
and U2284 (N_2284,N_2163,N_2202);
xnor U2285 (N_2285,N_2173,N_2200);
nand U2286 (N_2286,N_2103,N_2042);
or U2287 (N_2287,N_2109,N_2199);
nor U2288 (N_2288,N_2052,N_2236);
or U2289 (N_2289,N_2119,N_2145);
xnor U2290 (N_2290,N_2187,N_2240);
and U2291 (N_2291,N_2165,N_2180);
xnor U2292 (N_2292,N_2242,N_2168);
and U2293 (N_2293,N_2019,N_2190);
or U2294 (N_2294,N_2097,N_2118);
xor U2295 (N_2295,N_2104,N_2129);
nand U2296 (N_2296,N_2096,N_2241);
and U2297 (N_2297,N_2159,N_2246);
and U2298 (N_2298,N_2125,N_2247);
nor U2299 (N_2299,N_2024,N_2152);
and U2300 (N_2300,N_2147,N_2164);
xnor U2301 (N_2301,N_2203,N_2055);
nand U2302 (N_2302,N_2110,N_2066);
nor U2303 (N_2303,N_2196,N_2224);
xnor U2304 (N_2304,N_2005,N_2010);
and U2305 (N_2305,N_2093,N_2039);
and U2306 (N_2306,N_2003,N_2225);
nor U2307 (N_2307,N_2174,N_2178);
nor U2308 (N_2308,N_2232,N_2068);
nor U2309 (N_2309,N_2051,N_2011);
xor U2310 (N_2310,N_2014,N_2230);
and U2311 (N_2311,N_2023,N_2150);
or U2312 (N_2312,N_2036,N_2035);
nor U2313 (N_2313,N_2222,N_2077);
nand U2314 (N_2314,N_2007,N_2015);
nor U2315 (N_2315,N_2191,N_2155);
xnor U2316 (N_2316,N_2056,N_2101);
and U2317 (N_2317,N_2223,N_2049);
or U2318 (N_2318,N_2217,N_2211);
or U2319 (N_2319,N_2221,N_2047);
and U2320 (N_2320,N_2095,N_2227);
and U2321 (N_2321,N_2017,N_2192);
or U2322 (N_2322,N_2092,N_2212);
nor U2323 (N_2323,N_2151,N_2022);
nor U2324 (N_2324,N_2086,N_2090);
or U2325 (N_2325,N_2201,N_2215);
and U2326 (N_2326,N_2148,N_2063);
nor U2327 (N_2327,N_2122,N_2244);
and U2328 (N_2328,N_2186,N_2245);
and U2329 (N_2329,N_2181,N_2231);
xnor U2330 (N_2330,N_2137,N_2074);
nand U2331 (N_2331,N_2032,N_2115);
or U2332 (N_2332,N_2140,N_2111);
nand U2333 (N_2333,N_2113,N_2013);
nand U2334 (N_2334,N_2070,N_2116);
nor U2335 (N_2335,N_2094,N_2228);
nor U2336 (N_2336,N_2001,N_2006);
nor U2337 (N_2337,N_2204,N_2008);
nor U2338 (N_2338,N_2220,N_2208);
and U2339 (N_2339,N_2107,N_2102);
xor U2340 (N_2340,N_2038,N_2037);
or U2341 (N_2341,N_2108,N_2050);
xor U2342 (N_2342,N_2235,N_2135);
or U2343 (N_2343,N_2166,N_2069);
and U2344 (N_2344,N_2226,N_2054);
and U2345 (N_2345,N_2177,N_2188);
and U2346 (N_2346,N_2126,N_2139);
and U2347 (N_2347,N_2158,N_2130);
nor U2348 (N_2348,N_2046,N_2071);
and U2349 (N_2349,N_2004,N_2210);
nand U2350 (N_2350,N_2141,N_2176);
or U2351 (N_2351,N_2167,N_2121);
nand U2352 (N_2352,N_2076,N_2195);
nor U2353 (N_2353,N_2194,N_2154);
and U2354 (N_2354,N_2248,N_2157);
or U2355 (N_2355,N_2172,N_2207);
nand U2356 (N_2356,N_2099,N_2193);
xnor U2357 (N_2357,N_2100,N_2123);
and U2358 (N_2358,N_2219,N_2058);
or U2359 (N_2359,N_2238,N_2170);
or U2360 (N_2360,N_2106,N_2089);
and U2361 (N_2361,N_2197,N_2073);
xor U2362 (N_2362,N_2067,N_2029);
nand U2363 (N_2363,N_2044,N_2091);
nor U2364 (N_2364,N_2117,N_2048);
nand U2365 (N_2365,N_2030,N_2082);
or U2366 (N_2366,N_2146,N_2218);
nand U2367 (N_2367,N_2088,N_2081);
nand U2368 (N_2368,N_2079,N_2175);
nor U2369 (N_2369,N_2002,N_2136);
and U2370 (N_2370,N_2098,N_2127);
nand U2371 (N_2371,N_2144,N_2149);
nand U2372 (N_2372,N_2083,N_2114);
and U2373 (N_2373,N_2000,N_2233);
nor U2374 (N_2374,N_2183,N_2169);
nand U2375 (N_2375,N_2106,N_2012);
and U2376 (N_2376,N_2086,N_2168);
or U2377 (N_2377,N_2197,N_2055);
and U2378 (N_2378,N_2087,N_2226);
nand U2379 (N_2379,N_2073,N_2051);
or U2380 (N_2380,N_2127,N_2061);
or U2381 (N_2381,N_2187,N_2144);
nand U2382 (N_2382,N_2043,N_2054);
nor U2383 (N_2383,N_2054,N_2053);
xnor U2384 (N_2384,N_2071,N_2211);
xnor U2385 (N_2385,N_2143,N_2214);
nand U2386 (N_2386,N_2129,N_2044);
nand U2387 (N_2387,N_2219,N_2103);
or U2388 (N_2388,N_2087,N_2235);
nand U2389 (N_2389,N_2009,N_2238);
and U2390 (N_2390,N_2097,N_2237);
nand U2391 (N_2391,N_2061,N_2146);
or U2392 (N_2392,N_2022,N_2177);
and U2393 (N_2393,N_2207,N_2181);
nand U2394 (N_2394,N_2043,N_2060);
and U2395 (N_2395,N_2090,N_2149);
nor U2396 (N_2396,N_2221,N_2080);
or U2397 (N_2397,N_2086,N_2189);
nand U2398 (N_2398,N_2100,N_2128);
nand U2399 (N_2399,N_2106,N_2150);
nand U2400 (N_2400,N_2126,N_2007);
nor U2401 (N_2401,N_2130,N_2092);
or U2402 (N_2402,N_2049,N_2064);
nand U2403 (N_2403,N_2005,N_2104);
or U2404 (N_2404,N_2190,N_2061);
or U2405 (N_2405,N_2023,N_2248);
and U2406 (N_2406,N_2044,N_2054);
nand U2407 (N_2407,N_2169,N_2072);
and U2408 (N_2408,N_2191,N_2232);
nor U2409 (N_2409,N_2220,N_2015);
or U2410 (N_2410,N_2143,N_2066);
nand U2411 (N_2411,N_2134,N_2085);
xnor U2412 (N_2412,N_2145,N_2224);
or U2413 (N_2413,N_2227,N_2033);
or U2414 (N_2414,N_2101,N_2118);
xnor U2415 (N_2415,N_2170,N_2133);
xor U2416 (N_2416,N_2167,N_2093);
nand U2417 (N_2417,N_2220,N_2033);
and U2418 (N_2418,N_2086,N_2170);
nand U2419 (N_2419,N_2008,N_2246);
xnor U2420 (N_2420,N_2107,N_2026);
nand U2421 (N_2421,N_2098,N_2194);
nand U2422 (N_2422,N_2009,N_2116);
and U2423 (N_2423,N_2231,N_2075);
and U2424 (N_2424,N_2126,N_2190);
and U2425 (N_2425,N_2003,N_2237);
or U2426 (N_2426,N_2165,N_2011);
xor U2427 (N_2427,N_2021,N_2128);
xnor U2428 (N_2428,N_2005,N_2192);
and U2429 (N_2429,N_2241,N_2074);
xor U2430 (N_2430,N_2091,N_2020);
and U2431 (N_2431,N_2053,N_2149);
or U2432 (N_2432,N_2009,N_2121);
or U2433 (N_2433,N_2029,N_2100);
xor U2434 (N_2434,N_2085,N_2185);
and U2435 (N_2435,N_2080,N_2228);
nand U2436 (N_2436,N_2248,N_2008);
or U2437 (N_2437,N_2213,N_2041);
and U2438 (N_2438,N_2036,N_2220);
nor U2439 (N_2439,N_2108,N_2216);
nand U2440 (N_2440,N_2039,N_2026);
nor U2441 (N_2441,N_2231,N_2246);
xnor U2442 (N_2442,N_2083,N_2067);
nor U2443 (N_2443,N_2094,N_2011);
xor U2444 (N_2444,N_2091,N_2114);
nor U2445 (N_2445,N_2244,N_2191);
nand U2446 (N_2446,N_2245,N_2048);
and U2447 (N_2447,N_2038,N_2055);
or U2448 (N_2448,N_2243,N_2090);
or U2449 (N_2449,N_2073,N_2187);
and U2450 (N_2450,N_2231,N_2174);
xor U2451 (N_2451,N_2041,N_2111);
or U2452 (N_2452,N_2084,N_2063);
and U2453 (N_2453,N_2118,N_2243);
or U2454 (N_2454,N_2171,N_2108);
xnor U2455 (N_2455,N_2158,N_2193);
and U2456 (N_2456,N_2072,N_2023);
nand U2457 (N_2457,N_2017,N_2168);
nand U2458 (N_2458,N_2209,N_2081);
and U2459 (N_2459,N_2087,N_2230);
nand U2460 (N_2460,N_2207,N_2196);
xnor U2461 (N_2461,N_2024,N_2215);
nor U2462 (N_2462,N_2014,N_2118);
nor U2463 (N_2463,N_2040,N_2112);
nor U2464 (N_2464,N_2066,N_2027);
xnor U2465 (N_2465,N_2246,N_2081);
nor U2466 (N_2466,N_2007,N_2102);
nand U2467 (N_2467,N_2108,N_2105);
and U2468 (N_2468,N_2150,N_2186);
nand U2469 (N_2469,N_2226,N_2106);
nand U2470 (N_2470,N_2249,N_2199);
nand U2471 (N_2471,N_2032,N_2215);
xor U2472 (N_2472,N_2190,N_2194);
or U2473 (N_2473,N_2060,N_2139);
nor U2474 (N_2474,N_2164,N_2134);
nor U2475 (N_2475,N_2171,N_2100);
nor U2476 (N_2476,N_2141,N_2104);
and U2477 (N_2477,N_2008,N_2016);
and U2478 (N_2478,N_2074,N_2197);
nor U2479 (N_2479,N_2081,N_2185);
or U2480 (N_2480,N_2060,N_2210);
or U2481 (N_2481,N_2229,N_2042);
and U2482 (N_2482,N_2153,N_2029);
nand U2483 (N_2483,N_2209,N_2099);
and U2484 (N_2484,N_2160,N_2225);
and U2485 (N_2485,N_2038,N_2084);
xnor U2486 (N_2486,N_2042,N_2047);
nor U2487 (N_2487,N_2150,N_2237);
or U2488 (N_2488,N_2009,N_2197);
nor U2489 (N_2489,N_2081,N_2086);
and U2490 (N_2490,N_2138,N_2187);
and U2491 (N_2491,N_2161,N_2132);
nor U2492 (N_2492,N_2100,N_2219);
nand U2493 (N_2493,N_2056,N_2063);
nor U2494 (N_2494,N_2101,N_2216);
xor U2495 (N_2495,N_2110,N_2219);
xnor U2496 (N_2496,N_2092,N_2211);
nand U2497 (N_2497,N_2056,N_2175);
nand U2498 (N_2498,N_2204,N_2164);
or U2499 (N_2499,N_2039,N_2087);
nor U2500 (N_2500,N_2358,N_2386);
nor U2501 (N_2501,N_2261,N_2339);
nor U2502 (N_2502,N_2364,N_2421);
nor U2503 (N_2503,N_2300,N_2461);
nor U2504 (N_2504,N_2411,N_2474);
nor U2505 (N_2505,N_2438,N_2455);
xor U2506 (N_2506,N_2468,N_2304);
or U2507 (N_2507,N_2344,N_2490);
xor U2508 (N_2508,N_2382,N_2340);
nor U2509 (N_2509,N_2273,N_2478);
and U2510 (N_2510,N_2472,N_2329);
nor U2511 (N_2511,N_2426,N_2464);
nand U2512 (N_2512,N_2345,N_2416);
or U2513 (N_2513,N_2264,N_2487);
nand U2514 (N_2514,N_2310,N_2308);
nor U2515 (N_2515,N_2362,N_2370);
nor U2516 (N_2516,N_2491,N_2425);
nand U2517 (N_2517,N_2473,N_2497);
xor U2518 (N_2518,N_2326,N_2267);
nor U2519 (N_2519,N_2439,N_2289);
nand U2520 (N_2520,N_2436,N_2318);
xor U2521 (N_2521,N_2453,N_2260);
nor U2522 (N_2522,N_2315,N_2409);
xnor U2523 (N_2523,N_2299,N_2337);
and U2524 (N_2524,N_2263,N_2395);
nand U2525 (N_2525,N_2332,N_2417);
or U2526 (N_2526,N_2458,N_2429);
nor U2527 (N_2527,N_2305,N_2306);
xor U2528 (N_2528,N_2302,N_2493);
and U2529 (N_2529,N_2369,N_2482);
xor U2530 (N_2530,N_2283,N_2367);
nand U2531 (N_2531,N_2287,N_2422);
xor U2532 (N_2532,N_2400,N_2291);
xnor U2533 (N_2533,N_2488,N_2418);
nand U2534 (N_2534,N_2286,N_2266);
nor U2535 (N_2535,N_2277,N_2408);
or U2536 (N_2536,N_2385,N_2486);
xnor U2537 (N_2537,N_2448,N_2419);
or U2538 (N_2538,N_2377,N_2250);
xnor U2539 (N_2539,N_2324,N_2272);
and U2540 (N_2540,N_2372,N_2351);
nor U2541 (N_2541,N_2251,N_2450);
or U2542 (N_2542,N_2341,N_2252);
and U2543 (N_2543,N_2398,N_2432);
and U2544 (N_2544,N_2405,N_2471);
and U2545 (N_2545,N_2465,N_2470);
and U2546 (N_2546,N_2262,N_2288);
nor U2547 (N_2547,N_2394,N_2281);
or U2548 (N_2548,N_2285,N_2402);
nand U2549 (N_2549,N_2446,N_2295);
nor U2550 (N_2550,N_2357,N_2414);
and U2551 (N_2551,N_2375,N_2442);
or U2552 (N_2552,N_2483,N_2457);
and U2553 (N_2553,N_2327,N_2335);
nor U2554 (N_2554,N_2356,N_2420);
xnor U2555 (N_2555,N_2397,N_2368);
or U2556 (N_2556,N_2371,N_2480);
xnor U2557 (N_2557,N_2447,N_2390);
and U2558 (N_2558,N_2391,N_2309);
and U2559 (N_2559,N_2477,N_2469);
nor U2560 (N_2560,N_2325,N_2270);
nand U2561 (N_2561,N_2431,N_2338);
nand U2562 (N_2562,N_2254,N_2349);
and U2563 (N_2563,N_2437,N_2415);
and U2564 (N_2564,N_2492,N_2380);
nand U2565 (N_2565,N_2336,N_2365);
nor U2566 (N_2566,N_2342,N_2494);
or U2567 (N_2567,N_2354,N_2451);
or U2568 (N_2568,N_2423,N_2284);
or U2569 (N_2569,N_2430,N_2279);
and U2570 (N_2570,N_2406,N_2258);
or U2571 (N_2571,N_2361,N_2403);
nand U2572 (N_2572,N_2489,N_2294);
and U2573 (N_2573,N_2347,N_2481);
nand U2574 (N_2574,N_2399,N_2388);
xnor U2575 (N_2575,N_2434,N_2296);
and U2576 (N_2576,N_2352,N_2293);
or U2577 (N_2577,N_2343,N_2498);
nor U2578 (N_2578,N_2333,N_2407);
and U2579 (N_2579,N_2313,N_2381);
nor U2580 (N_2580,N_2499,N_2387);
and U2581 (N_2581,N_2307,N_2275);
or U2582 (N_2582,N_2435,N_2330);
nand U2583 (N_2583,N_2355,N_2459);
and U2584 (N_2584,N_2314,N_2441);
or U2585 (N_2585,N_2462,N_2320);
xor U2586 (N_2586,N_2374,N_2378);
and U2587 (N_2587,N_2280,N_2401);
xor U2588 (N_2588,N_2346,N_2350);
nor U2589 (N_2589,N_2476,N_2392);
or U2590 (N_2590,N_2445,N_2466);
or U2591 (N_2591,N_2383,N_2323);
nor U2592 (N_2592,N_2256,N_2449);
or U2593 (N_2593,N_2297,N_2312);
xor U2594 (N_2594,N_2298,N_2290);
xnor U2595 (N_2595,N_2485,N_2276);
or U2596 (N_2596,N_2257,N_2452);
nand U2597 (N_2597,N_2278,N_2301);
nand U2598 (N_2598,N_2467,N_2376);
or U2599 (N_2599,N_2389,N_2255);
or U2600 (N_2600,N_2440,N_2443);
xnor U2601 (N_2601,N_2410,N_2424);
nor U2602 (N_2602,N_2316,N_2463);
nand U2603 (N_2603,N_2363,N_2303);
nand U2604 (N_2604,N_2433,N_2396);
nor U2605 (N_2605,N_2331,N_2484);
nand U2606 (N_2606,N_2366,N_2384);
xnor U2607 (N_2607,N_2456,N_2322);
and U2608 (N_2608,N_2427,N_2269);
and U2609 (N_2609,N_2454,N_2274);
nor U2610 (N_2610,N_2348,N_2311);
xnor U2611 (N_2611,N_2259,N_2496);
nor U2612 (N_2612,N_2271,N_2268);
nand U2613 (N_2613,N_2479,N_2444);
and U2614 (N_2614,N_2328,N_2373);
nor U2615 (N_2615,N_2319,N_2413);
nand U2616 (N_2616,N_2282,N_2253);
nand U2617 (N_2617,N_2292,N_2428);
and U2618 (N_2618,N_2334,N_2379);
nand U2619 (N_2619,N_2495,N_2359);
xor U2620 (N_2620,N_2412,N_2317);
and U2621 (N_2621,N_2475,N_2393);
and U2622 (N_2622,N_2265,N_2404);
xnor U2623 (N_2623,N_2460,N_2353);
and U2624 (N_2624,N_2321,N_2360);
xnor U2625 (N_2625,N_2326,N_2379);
xor U2626 (N_2626,N_2455,N_2307);
xor U2627 (N_2627,N_2251,N_2302);
nor U2628 (N_2628,N_2402,N_2406);
xnor U2629 (N_2629,N_2358,N_2256);
nor U2630 (N_2630,N_2321,N_2446);
nor U2631 (N_2631,N_2480,N_2466);
or U2632 (N_2632,N_2396,N_2469);
nor U2633 (N_2633,N_2425,N_2372);
or U2634 (N_2634,N_2410,N_2423);
nor U2635 (N_2635,N_2303,N_2428);
or U2636 (N_2636,N_2344,N_2444);
nand U2637 (N_2637,N_2287,N_2258);
xnor U2638 (N_2638,N_2428,N_2431);
nor U2639 (N_2639,N_2283,N_2262);
nand U2640 (N_2640,N_2481,N_2475);
nor U2641 (N_2641,N_2307,N_2274);
nand U2642 (N_2642,N_2279,N_2374);
xnor U2643 (N_2643,N_2363,N_2480);
xnor U2644 (N_2644,N_2379,N_2408);
nor U2645 (N_2645,N_2418,N_2378);
and U2646 (N_2646,N_2385,N_2270);
nand U2647 (N_2647,N_2261,N_2445);
or U2648 (N_2648,N_2283,N_2452);
nand U2649 (N_2649,N_2433,N_2299);
nand U2650 (N_2650,N_2327,N_2453);
xor U2651 (N_2651,N_2274,N_2300);
xor U2652 (N_2652,N_2320,N_2437);
xor U2653 (N_2653,N_2346,N_2362);
xnor U2654 (N_2654,N_2411,N_2320);
and U2655 (N_2655,N_2438,N_2380);
nor U2656 (N_2656,N_2301,N_2474);
xnor U2657 (N_2657,N_2313,N_2278);
nand U2658 (N_2658,N_2428,N_2398);
nand U2659 (N_2659,N_2385,N_2268);
nor U2660 (N_2660,N_2443,N_2326);
nor U2661 (N_2661,N_2264,N_2308);
nand U2662 (N_2662,N_2436,N_2344);
or U2663 (N_2663,N_2327,N_2467);
nor U2664 (N_2664,N_2341,N_2285);
xnor U2665 (N_2665,N_2453,N_2325);
xnor U2666 (N_2666,N_2412,N_2321);
xor U2667 (N_2667,N_2490,N_2451);
nand U2668 (N_2668,N_2406,N_2279);
nand U2669 (N_2669,N_2450,N_2407);
nor U2670 (N_2670,N_2440,N_2282);
nand U2671 (N_2671,N_2299,N_2341);
nor U2672 (N_2672,N_2356,N_2345);
and U2673 (N_2673,N_2273,N_2363);
xnor U2674 (N_2674,N_2316,N_2482);
or U2675 (N_2675,N_2299,N_2357);
nor U2676 (N_2676,N_2261,N_2315);
nor U2677 (N_2677,N_2448,N_2383);
nor U2678 (N_2678,N_2495,N_2479);
nand U2679 (N_2679,N_2411,N_2368);
or U2680 (N_2680,N_2382,N_2272);
or U2681 (N_2681,N_2464,N_2497);
or U2682 (N_2682,N_2281,N_2491);
and U2683 (N_2683,N_2315,N_2424);
or U2684 (N_2684,N_2324,N_2282);
xor U2685 (N_2685,N_2340,N_2424);
nand U2686 (N_2686,N_2475,N_2432);
or U2687 (N_2687,N_2263,N_2274);
and U2688 (N_2688,N_2250,N_2442);
and U2689 (N_2689,N_2336,N_2361);
nand U2690 (N_2690,N_2343,N_2320);
nor U2691 (N_2691,N_2331,N_2321);
or U2692 (N_2692,N_2265,N_2389);
nand U2693 (N_2693,N_2287,N_2359);
xnor U2694 (N_2694,N_2467,N_2492);
nor U2695 (N_2695,N_2290,N_2475);
nand U2696 (N_2696,N_2417,N_2287);
nor U2697 (N_2697,N_2490,N_2325);
nand U2698 (N_2698,N_2457,N_2429);
xnor U2699 (N_2699,N_2343,N_2371);
or U2700 (N_2700,N_2385,N_2323);
nand U2701 (N_2701,N_2316,N_2479);
or U2702 (N_2702,N_2446,N_2491);
and U2703 (N_2703,N_2385,N_2279);
or U2704 (N_2704,N_2337,N_2343);
and U2705 (N_2705,N_2489,N_2443);
xor U2706 (N_2706,N_2279,N_2276);
nor U2707 (N_2707,N_2452,N_2451);
and U2708 (N_2708,N_2259,N_2352);
nand U2709 (N_2709,N_2466,N_2410);
nor U2710 (N_2710,N_2323,N_2262);
nand U2711 (N_2711,N_2464,N_2488);
nand U2712 (N_2712,N_2279,N_2405);
or U2713 (N_2713,N_2479,N_2307);
or U2714 (N_2714,N_2389,N_2468);
and U2715 (N_2715,N_2263,N_2261);
xor U2716 (N_2716,N_2462,N_2281);
xnor U2717 (N_2717,N_2492,N_2302);
nor U2718 (N_2718,N_2447,N_2488);
nand U2719 (N_2719,N_2426,N_2404);
nor U2720 (N_2720,N_2321,N_2299);
or U2721 (N_2721,N_2384,N_2440);
nand U2722 (N_2722,N_2427,N_2374);
and U2723 (N_2723,N_2393,N_2368);
and U2724 (N_2724,N_2313,N_2382);
or U2725 (N_2725,N_2273,N_2280);
nand U2726 (N_2726,N_2427,N_2293);
and U2727 (N_2727,N_2406,N_2271);
xor U2728 (N_2728,N_2335,N_2395);
xnor U2729 (N_2729,N_2353,N_2488);
xor U2730 (N_2730,N_2496,N_2310);
or U2731 (N_2731,N_2376,N_2396);
or U2732 (N_2732,N_2269,N_2337);
and U2733 (N_2733,N_2409,N_2288);
nand U2734 (N_2734,N_2317,N_2424);
xor U2735 (N_2735,N_2339,N_2253);
nand U2736 (N_2736,N_2358,N_2300);
xnor U2737 (N_2737,N_2465,N_2421);
and U2738 (N_2738,N_2468,N_2280);
nand U2739 (N_2739,N_2291,N_2313);
xor U2740 (N_2740,N_2376,N_2451);
or U2741 (N_2741,N_2296,N_2337);
or U2742 (N_2742,N_2388,N_2270);
or U2743 (N_2743,N_2447,N_2459);
nor U2744 (N_2744,N_2462,N_2383);
or U2745 (N_2745,N_2251,N_2359);
or U2746 (N_2746,N_2270,N_2333);
and U2747 (N_2747,N_2472,N_2412);
xnor U2748 (N_2748,N_2451,N_2363);
and U2749 (N_2749,N_2277,N_2253);
xor U2750 (N_2750,N_2673,N_2636);
or U2751 (N_2751,N_2660,N_2588);
and U2752 (N_2752,N_2732,N_2570);
or U2753 (N_2753,N_2736,N_2670);
xnor U2754 (N_2754,N_2669,N_2652);
or U2755 (N_2755,N_2663,N_2556);
or U2756 (N_2756,N_2526,N_2508);
and U2757 (N_2757,N_2701,N_2714);
and U2758 (N_2758,N_2733,N_2579);
and U2759 (N_2759,N_2541,N_2706);
nand U2760 (N_2760,N_2597,N_2598);
xor U2761 (N_2761,N_2726,N_2716);
or U2762 (N_2762,N_2645,N_2688);
and U2763 (N_2763,N_2538,N_2662);
xor U2764 (N_2764,N_2523,N_2692);
nand U2765 (N_2765,N_2703,N_2517);
and U2766 (N_2766,N_2728,N_2513);
nor U2767 (N_2767,N_2537,N_2699);
xor U2768 (N_2768,N_2543,N_2568);
and U2769 (N_2769,N_2525,N_2615);
and U2770 (N_2770,N_2519,N_2740);
or U2771 (N_2771,N_2647,N_2544);
or U2772 (N_2772,N_2718,N_2531);
xor U2773 (N_2773,N_2571,N_2631);
and U2774 (N_2774,N_2607,N_2576);
and U2775 (N_2775,N_2661,N_2533);
xnor U2776 (N_2776,N_2727,N_2539);
nand U2777 (N_2777,N_2651,N_2514);
or U2778 (N_2778,N_2616,N_2697);
or U2779 (N_2779,N_2634,N_2593);
nor U2780 (N_2780,N_2749,N_2618);
nand U2781 (N_2781,N_2656,N_2730);
and U2782 (N_2782,N_2552,N_2602);
and U2783 (N_2783,N_2545,N_2599);
or U2784 (N_2784,N_2592,N_2553);
xnor U2785 (N_2785,N_2562,N_2502);
nand U2786 (N_2786,N_2509,N_2698);
nand U2787 (N_2787,N_2725,N_2512);
nor U2788 (N_2788,N_2594,N_2516);
or U2789 (N_2789,N_2683,N_2561);
and U2790 (N_2790,N_2624,N_2610);
or U2791 (N_2791,N_2695,N_2528);
and U2792 (N_2792,N_2671,N_2687);
or U2793 (N_2793,N_2569,N_2711);
and U2794 (N_2794,N_2705,N_2685);
and U2795 (N_2795,N_2664,N_2518);
xnor U2796 (N_2796,N_2555,N_2583);
and U2797 (N_2797,N_2667,N_2551);
and U2798 (N_2798,N_2560,N_2620);
nor U2799 (N_2799,N_2735,N_2715);
nor U2800 (N_2800,N_2527,N_2748);
or U2801 (N_2801,N_2691,N_2680);
or U2802 (N_2802,N_2694,N_2710);
or U2803 (N_2803,N_2549,N_2621);
or U2804 (N_2804,N_2505,N_2741);
nor U2805 (N_2805,N_2632,N_2573);
nor U2806 (N_2806,N_2596,N_2734);
xor U2807 (N_2807,N_2613,N_2581);
or U2808 (N_2808,N_2640,N_2679);
xor U2809 (N_2809,N_2604,N_2693);
nand U2810 (N_2810,N_2739,N_2729);
nor U2811 (N_2811,N_2682,N_2511);
and U2812 (N_2812,N_2666,N_2582);
and U2813 (N_2813,N_2720,N_2665);
nand U2814 (N_2814,N_2707,N_2677);
and U2815 (N_2815,N_2678,N_2704);
and U2816 (N_2816,N_2719,N_2623);
xor U2817 (N_2817,N_2668,N_2619);
nand U2818 (N_2818,N_2737,N_2724);
nor U2819 (N_2819,N_2563,N_2622);
or U2820 (N_2820,N_2627,N_2655);
or U2821 (N_2821,N_2501,N_2689);
or U2822 (N_2822,N_2690,N_2743);
xor U2823 (N_2823,N_2535,N_2684);
nand U2824 (N_2824,N_2591,N_2589);
or U2825 (N_2825,N_2674,N_2595);
and U2826 (N_2826,N_2630,N_2547);
nor U2827 (N_2827,N_2575,N_2534);
xor U2828 (N_2828,N_2738,N_2530);
xor U2829 (N_2829,N_2565,N_2717);
and U2830 (N_2830,N_2574,N_2658);
or U2831 (N_2831,N_2659,N_2510);
or U2832 (N_2832,N_2567,N_2731);
or U2833 (N_2833,N_2587,N_2605);
nand U2834 (N_2834,N_2648,N_2586);
nand U2835 (N_2835,N_2612,N_2542);
nor U2836 (N_2836,N_2686,N_2629);
nor U2837 (N_2837,N_2696,N_2548);
xor U2838 (N_2838,N_2559,N_2637);
or U2839 (N_2839,N_2722,N_2600);
xor U2840 (N_2840,N_2676,N_2500);
or U2841 (N_2841,N_2708,N_2590);
xnor U2842 (N_2842,N_2601,N_2649);
or U2843 (N_2843,N_2520,N_2747);
nand U2844 (N_2844,N_2611,N_2578);
and U2845 (N_2845,N_2635,N_2625);
xor U2846 (N_2846,N_2745,N_2709);
and U2847 (N_2847,N_2529,N_2558);
xnor U2848 (N_2848,N_2580,N_2522);
or U2849 (N_2849,N_2723,N_2638);
xnor U2850 (N_2850,N_2700,N_2550);
nand U2851 (N_2851,N_2557,N_2577);
nand U2852 (N_2852,N_2643,N_2675);
or U2853 (N_2853,N_2650,N_2653);
nor U2854 (N_2854,N_2606,N_2546);
or U2855 (N_2855,N_2614,N_2503);
or U2856 (N_2856,N_2746,N_2744);
nand U2857 (N_2857,N_2584,N_2524);
nand U2858 (N_2858,N_2672,N_2639);
xnor U2859 (N_2859,N_2713,N_2515);
and U2860 (N_2860,N_2628,N_2642);
nor U2861 (N_2861,N_2702,N_2654);
nand U2862 (N_2862,N_2633,N_2609);
nand U2863 (N_2863,N_2681,N_2540);
and U2864 (N_2864,N_2504,N_2657);
xor U2865 (N_2865,N_2521,N_2507);
nand U2866 (N_2866,N_2564,N_2712);
or U2867 (N_2867,N_2536,N_2644);
and U2868 (N_2868,N_2617,N_2626);
nand U2869 (N_2869,N_2572,N_2641);
and U2870 (N_2870,N_2608,N_2506);
and U2871 (N_2871,N_2646,N_2554);
nand U2872 (N_2872,N_2585,N_2742);
xor U2873 (N_2873,N_2566,N_2532);
and U2874 (N_2874,N_2603,N_2721);
nand U2875 (N_2875,N_2624,N_2718);
nor U2876 (N_2876,N_2690,N_2575);
xnor U2877 (N_2877,N_2646,N_2703);
and U2878 (N_2878,N_2570,N_2718);
nand U2879 (N_2879,N_2638,N_2570);
and U2880 (N_2880,N_2677,N_2567);
or U2881 (N_2881,N_2689,N_2638);
xnor U2882 (N_2882,N_2583,N_2681);
or U2883 (N_2883,N_2542,N_2544);
and U2884 (N_2884,N_2563,N_2703);
or U2885 (N_2885,N_2605,N_2651);
xor U2886 (N_2886,N_2649,N_2605);
nor U2887 (N_2887,N_2608,N_2716);
xnor U2888 (N_2888,N_2574,N_2737);
and U2889 (N_2889,N_2711,N_2723);
nand U2890 (N_2890,N_2635,N_2641);
xnor U2891 (N_2891,N_2611,N_2597);
xor U2892 (N_2892,N_2500,N_2585);
or U2893 (N_2893,N_2594,N_2581);
xnor U2894 (N_2894,N_2739,N_2556);
and U2895 (N_2895,N_2738,N_2596);
nand U2896 (N_2896,N_2550,N_2585);
and U2897 (N_2897,N_2748,N_2513);
and U2898 (N_2898,N_2508,N_2666);
and U2899 (N_2899,N_2579,N_2700);
and U2900 (N_2900,N_2610,N_2508);
or U2901 (N_2901,N_2570,N_2657);
and U2902 (N_2902,N_2698,N_2512);
nor U2903 (N_2903,N_2589,N_2614);
or U2904 (N_2904,N_2716,N_2649);
or U2905 (N_2905,N_2553,N_2546);
nand U2906 (N_2906,N_2644,N_2531);
xor U2907 (N_2907,N_2692,N_2505);
nor U2908 (N_2908,N_2598,N_2629);
nand U2909 (N_2909,N_2726,N_2578);
and U2910 (N_2910,N_2682,N_2565);
or U2911 (N_2911,N_2711,N_2566);
or U2912 (N_2912,N_2515,N_2706);
nor U2913 (N_2913,N_2513,N_2691);
nor U2914 (N_2914,N_2706,N_2576);
nor U2915 (N_2915,N_2741,N_2514);
and U2916 (N_2916,N_2694,N_2605);
and U2917 (N_2917,N_2563,N_2560);
nand U2918 (N_2918,N_2675,N_2627);
nand U2919 (N_2919,N_2639,N_2633);
xor U2920 (N_2920,N_2613,N_2542);
and U2921 (N_2921,N_2709,N_2626);
nor U2922 (N_2922,N_2597,N_2548);
or U2923 (N_2923,N_2545,N_2523);
nor U2924 (N_2924,N_2587,N_2599);
and U2925 (N_2925,N_2522,N_2681);
or U2926 (N_2926,N_2563,N_2646);
xor U2927 (N_2927,N_2696,N_2672);
nor U2928 (N_2928,N_2613,N_2643);
nor U2929 (N_2929,N_2685,N_2655);
or U2930 (N_2930,N_2501,N_2552);
nor U2931 (N_2931,N_2562,N_2581);
or U2932 (N_2932,N_2553,N_2540);
and U2933 (N_2933,N_2707,N_2688);
nor U2934 (N_2934,N_2515,N_2719);
and U2935 (N_2935,N_2616,N_2640);
xnor U2936 (N_2936,N_2500,N_2739);
nand U2937 (N_2937,N_2692,N_2597);
nand U2938 (N_2938,N_2535,N_2616);
xor U2939 (N_2939,N_2609,N_2736);
xor U2940 (N_2940,N_2667,N_2568);
nor U2941 (N_2941,N_2737,N_2659);
nor U2942 (N_2942,N_2686,N_2709);
xor U2943 (N_2943,N_2695,N_2568);
nand U2944 (N_2944,N_2660,N_2542);
xnor U2945 (N_2945,N_2593,N_2646);
nand U2946 (N_2946,N_2643,N_2697);
or U2947 (N_2947,N_2657,N_2597);
nand U2948 (N_2948,N_2665,N_2529);
nor U2949 (N_2949,N_2683,N_2746);
nand U2950 (N_2950,N_2618,N_2572);
nor U2951 (N_2951,N_2696,N_2627);
and U2952 (N_2952,N_2605,N_2724);
and U2953 (N_2953,N_2520,N_2564);
nor U2954 (N_2954,N_2655,N_2738);
nand U2955 (N_2955,N_2506,N_2604);
xor U2956 (N_2956,N_2693,N_2631);
or U2957 (N_2957,N_2689,N_2661);
nor U2958 (N_2958,N_2676,N_2709);
xnor U2959 (N_2959,N_2672,N_2586);
nand U2960 (N_2960,N_2712,N_2681);
nor U2961 (N_2961,N_2500,N_2621);
nor U2962 (N_2962,N_2584,N_2708);
or U2963 (N_2963,N_2708,N_2654);
and U2964 (N_2964,N_2545,N_2515);
xor U2965 (N_2965,N_2690,N_2542);
nor U2966 (N_2966,N_2717,N_2683);
nand U2967 (N_2967,N_2557,N_2566);
nor U2968 (N_2968,N_2660,N_2731);
or U2969 (N_2969,N_2641,N_2593);
nor U2970 (N_2970,N_2509,N_2654);
and U2971 (N_2971,N_2642,N_2516);
nand U2972 (N_2972,N_2736,N_2553);
nor U2973 (N_2973,N_2602,N_2714);
nand U2974 (N_2974,N_2564,N_2546);
and U2975 (N_2975,N_2736,N_2730);
and U2976 (N_2976,N_2747,N_2514);
or U2977 (N_2977,N_2597,N_2616);
and U2978 (N_2978,N_2541,N_2620);
nor U2979 (N_2979,N_2579,N_2726);
nand U2980 (N_2980,N_2711,N_2526);
or U2981 (N_2981,N_2685,N_2538);
xnor U2982 (N_2982,N_2558,N_2553);
xor U2983 (N_2983,N_2561,N_2596);
nor U2984 (N_2984,N_2748,N_2720);
nor U2985 (N_2985,N_2549,N_2503);
nand U2986 (N_2986,N_2676,N_2526);
and U2987 (N_2987,N_2634,N_2529);
or U2988 (N_2988,N_2650,N_2557);
nand U2989 (N_2989,N_2668,N_2714);
or U2990 (N_2990,N_2601,N_2623);
xnor U2991 (N_2991,N_2672,N_2526);
nand U2992 (N_2992,N_2507,N_2684);
xor U2993 (N_2993,N_2709,N_2590);
nand U2994 (N_2994,N_2654,N_2731);
xnor U2995 (N_2995,N_2545,N_2650);
nor U2996 (N_2996,N_2509,N_2730);
xor U2997 (N_2997,N_2596,N_2531);
and U2998 (N_2998,N_2675,N_2629);
and U2999 (N_2999,N_2670,N_2539);
nor U3000 (N_3000,N_2944,N_2918);
and U3001 (N_3001,N_2956,N_2910);
nor U3002 (N_3002,N_2809,N_2883);
xnor U3003 (N_3003,N_2840,N_2777);
and U3004 (N_3004,N_2926,N_2999);
and U3005 (N_3005,N_2933,N_2882);
or U3006 (N_3006,N_2990,N_2808);
nand U3007 (N_3007,N_2753,N_2997);
xnor U3008 (N_3008,N_2906,N_2874);
xnor U3009 (N_3009,N_2811,N_2837);
or U3010 (N_3010,N_2820,N_2986);
nor U3011 (N_3011,N_2915,N_2920);
xor U3012 (N_3012,N_2832,N_2873);
nor U3013 (N_3013,N_2781,N_2785);
nand U3014 (N_3014,N_2912,N_2767);
nor U3015 (N_3015,N_2876,N_2869);
and U3016 (N_3016,N_2831,N_2967);
and U3017 (N_3017,N_2804,N_2846);
and U3018 (N_3018,N_2935,N_2870);
and U3019 (N_3019,N_2819,N_2988);
nand U3020 (N_3020,N_2973,N_2851);
or U3021 (N_3021,N_2864,N_2858);
xnor U3022 (N_3022,N_2798,N_2843);
xor U3023 (N_3023,N_2818,N_2927);
or U3024 (N_3024,N_2959,N_2860);
and U3025 (N_3025,N_2760,N_2756);
nand U3026 (N_3026,N_2751,N_2937);
or U3027 (N_3027,N_2904,N_2932);
nor U3028 (N_3028,N_2847,N_2752);
nand U3029 (N_3029,N_2815,N_2881);
xor U3030 (N_3030,N_2963,N_2845);
or U3031 (N_3031,N_2946,N_2909);
xor U3032 (N_3032,N_2816,N_2795);
nand U3033 (N_3033,N_2784,N_2992);
nor U3034 (N_3034,N_2991,N_2902);
or U3035 (N_3035,N_2953,N_2897);
or U3036 (N_3036,N_2850,N_2810);
and U3037 (N_3037,N_2805,N_2993);
or U3038 (N_3038,N_2759,N_2768);
nor U3039 (N_3039,N_2916,N_2769);
and U3040 (N_3040,N_2930,N_2823);
or U3041 (N_3041,N_2822,N_2940);
nor U3042 (N_3042,N_2981,N_2901);
xnor U3043 (N_3043,N_2828,N_2865);
and U3044 (N_3044,N_2826,N_2825);
and U3045 (N_3045,N_2779,N_2880);
nor U3046 (N_3046,N_2895,N_2894);
nand U3047 (N_3047,N_2834,N_2854);
nor U3048 (N_3048,N_2970,N_2939);
xor U3049 (N_3049,N_2841,N_2955);
and U3050 (N_3050,N_2766,N_2971);
and U3051 (N_3051,N_2855,N_2764);
nor U3052 (N_3052,N_2821,N_2985);
nand U3053 (N_3053,N_2977,N_2788);
nor U3054 (N_3054,N_2879,N_2774);
or U3055 (N_3055,N_2789,N_2799);
or U3056 (N_3056,N_2833,N_2857);
nand U3057 (N_3057,N_2903,N_2979);
nand U3058 (N_3058,N_2758,N_2787);
xor U3059 (N_3059,N_2954,N_2907);
xnor U3060 (N_3060,N_2890,N_2972);
and U3061 (N_3061,N_2908,N_2861);
nand U3062 (N_3062,N_2797,N_2807);
nor U3063 (N_3063,N_2998,N_2950);
and U3064 (N_3064,N_2987,N_2800);
and U3065 (N_3065,N_2934,N_2975);
and U3066 (N_3066,N_2887,N_2806);
and U3067 (N_3067,N_2761,N_2824);
nand U3068 (N_3068,N_2814,N_2817);
nor U3069 (N_3069,N_2771,N_2938);
nor U3070 (N_3070,N_2871,N_2849);
nor U3071 (N_3071,N_2796,N_2856);
and U3072 (N_3072,N_2965,N_2786);
or U3073 (N_3073,N_2896,N_2919);
nor U3074 (N_3074,N_2866,N_2958);
nand U3075 (N_3075,N_2925,N_2936);
nor U3076 (N_3076,N_2862,N_2829);
nand U3077 (N_3077,N_2772,N_2921);
nor U3078 (N_3078,N_2966,N_2877);
nand U3079 (N_3079,N_2917,N_2852);
and U3080 (N_3080,N_2983,N_2848);
and U3081 (N_3081,N_2949,N_2969);
nor U3082 (N_3082,N_2948,N_2941);
and U3083 (N_3083,N_2863,N_2951);
or U3084 (N_3084,N_2780,N_2929);
nor U3085 (N_3085,N_2775,N_2762);
or U3086 (N_3086,N_2754,N_2844);
xor U3087 (N_3087,N_2773,N_2962);
nor U3088 (N_3088,N_2812,N_2928);
or U3089 (N_3089,N_2889,N_2763);
xor U3090 (N_3090,N_2984,N_2899);
nand U3091 (N_3091,N_2924,N_2922);
xnor U3092 (N_3092,N_2978,N_2960);
or U3093 (N_3093,N_2947,N_2957);
or U3094 (N_3094,N_2867,N_2982);
and U3095 (N_3095,N_2842,N_2980);
or U3096 (N_3096,N_2838,N_2770);
and U3097 (N_3097,N_2790,N_2835);
nand U3098 (N_3098,N_2778,N_2923);
xor U3099 (N_3099,N_2961,N_2859);
nor U3100 (N_3100,N_2943,N_2827);
or U3101 (N_3101,N_2803,N_2911);
nor U3102 (N_3102,N_2885,N_2952);
xor U3103 (N_3103,N_2898,N_2996);
or U3104 (N_3104,N_2776,N_2878);
nand U3105 (N_3105,N_2931,N_2868);
or U3106 (N_3106,N_2791,N_2989);
nor U3107 (N_3107,N_2765,N_2976);
xor U3108 (N_3108,N_2994,N_2892);
and U3109 (N_3109,N_2830,N_2801);
nand U3110 (N_3110,N_2793,N_2802);
nand U3111 (N_3111,N_2893,N_2872);
and U3112 (N_3112,N_2968,N_2839);
xnor U3113 (N_3113,N_2792,N_2886);
nor U3114 (N_3114,N_2813,N_2884);
nor U3115 (N_3115,N_2853,N_2794);
nand U3116 (N_3116,N_2945,N_2888);
nor U3117 (N_3117,N_2914,N_2836);
xor U3118 (N_3118,N_2913,N_2905);
and U3119 (N_3119,N_2782,N_2875);
or U3120 (N_3120,N_2750,N_2900);
xnor U3121 (N_3121,N_2783,N_2995);
or U3122 (N_3122,N_2757,N_2974);
xor U3123 (N_3123,N_2755,N_2891);
and U3124 (N_3124,N_2942,N_2964);
or U3125 (N_3125,N_2833,N_2977);
nand U3126 (N_3126,N_2837,N_2874);
nand U3127 (N_3127,N_2856,N_2842);
and U3128 (N_3128,N_2819,N_2773);
and U3129 (N_3129,N_2957,N_2803);
or U3130 (N_3130,N_2957,N_2905);
nand U3131 (N_3131,N_2976,N_2851);
nand U3132 (N_3132,N_2891,N_2947);
or U3133 (N_3133,N_2977,N_2925);
or U3134 (N_3134,N_2849,N_2901);
nand U3135 (N_3135,N_2798,N_2763);
or U3136 (N_3136,N_2956,N_2760);
or U3137 (N_3137,N_2937,N_2805);
nor U3138 (N_3138,N_2783,N_2872);
or U3139 (N_3139,N_2807,N_2831);
nand U3140 (N_3140,N_2767,N_2854);
and U3141 (N_3141,N_2923,N_2898);
or U3142 (N_3142,N_2937,N_2840);
xnor U3143 (N_3143,N_2834,N_2764);
and U3144 (N_3144,N_2885,N_2916);
and U3145 (N_3145,N_2968,N_2766);
nor U3146 (N_3146,N_2883,N_2829);
and U3147 (N_3147,N_2912,N_2808);
nand U3148 (N_3148,N_2825,N_2818);
and U3149 (N_3149,N_2913,N_2976);
xnor U3150 (N_3150,N_2875,N_2994);
and U3151 (N_3151,N_2807,N_2762);
nor U3152 (N_3152,N_2899,N_2895);
and U3153 (N_3153,N_2944,N_2860);
nand U3154 (N_3154,N_2947,N_2895);
xnor U3155 (N_3155,N_2849,N_2757);
or U3156 (N_3156,N_2830,N_2817);
nand U3157 (N_3157,N_2919,N_2790);
xor U3158 (N_3158,N_2875,N_2925);
nand U3159 (N_3159,N_2845,N_2971);
nand U3160 (N_3160,N_2947,N_2795);
and U3161 (N_3161,N_2942,N_2882);
and U3162 (N_3162,N_2890,N_2852);
nor U3163 (N_3163,N_2858,N_2802);
xnor U3164 (N_3164,N_2849,N_2872);
or U3165 (N_3165,N_2915,N_2926);
xnor U3166 (N_3166,N_2862,N_2784);
or U3167 (N_3167,N_2787,N_2851);
or U3168 (N_3168,N_2995,N_2957);
nand U3169 (N_3169,N_2858,N_2842);
and U3170 (N_3170,N_2974,N_2815);
nor U3171 (N_3171,N_2857,N_2928);
and U3172 (N_3172,N_2833,N_2981);
and U3173 (N_3173,N_2908,N_2979);
nand U3174 (N_3174,N_2925,N_2818);
nand U3175 (N_3175,N_2758,N_2850);
or U3176 (N_3176,N_2876,N_2838);
and U3177 (N_3177,N_2905,N_2791);
nand U3178 (N_3178,N_2803,N_2980);
and U3179 (N_3179,N_2955,N_2975);
or U3180 (N_3180,N_2766,N_2819);
nor U3181 (N_3181,N_2912,N_2795);
or U3182 (N_3182,N_2899,N_2858);
nand U3183 (N_3183,N_2939,N_2783);
and U3184 (N_3184,N_2932,N_2830);
nor U3185 (N_3185,N_2895,N_2962);
nand U3186 (N_3186,N_2816,N_2885);
and U3187 (N_3187,N_2931,N_2887);
nor U3188 (N_3188,N_2850,N_2845);
nand U3189 (N_3189,N_2846,N_2976);
nor U3190 (N_3190,N_2775,N_2996);
xnor U3191 (N_3191,N_2965,N_2901);
nand U3192 (N_3192,N_2839,N_2960);
nand U3193 (N_3193,N_2758,N_2910);
and U3194 (N_3194,N_2978,N_2820);
or U3195 (N_3195,N_2833,N_2914);
xor U3196 (N_3196,N_2784,N_2954);
and U3197 (N_3197,N_2823,N_2819);
and U3198 (N_3198,N_2996,N_2941);
or U3199 (N_3199,N_2955,N_2875);
xnor U3200 (N_3200,N_2805,N_2816);
nand U3201 (N_3201,N_2907,N_2823);
nor U3202 (N_3202,N_2839,N_2976);
nor U3203 (N_3203,N_2949,N_2815);
nor U3204 (N_3204,N_2796,N_2941);
nor U3205 (N_3205,N_2954,N_2860);
and U3206 (N_3206,N_2877,N_2967);
and U3207 (N_3207,N_2808,N_2814);
and U3208 (N_3208,N_2822,N_2814);
nand U3209 (N_3209,N_2778,N_2753);
nor U3210 (N_3210,N_2848,N_2951);
or U3211 (N_3211,N_2956,N_2811);
xnor U3212 (N_3212,N_2783,N_2787);
nor U3213 (N_3213,N_2998,N_2776);
or U3214 (N_3214,N_2785,N_2824);
or U3215 (N_3215,N_2865,N_2795);
nor U3216 (N_3216,N_2844,N_2762);
and U3217 (N_3217,N_2878,N_2966);
or U3218 (N_3218,N_2955,N_2797);
or U3219 (N_3219,N_2969,N_2815);
xor U3220 (N_3220,N_2910,N_2864);
and U3221 (N_3221,N_2842,N_2757);
nand U3222 (N_3222,N_2880,N_2960);
or U3223 (N_3223,N_2864,N_2950);
nor U3224 (N_3224,N_2851,N_2790);
nor U3225 (N_3225,N_2959,N_2839);
or U3226 (N_3226,N_2837,N_2877);
xnor U3227 (N_3227,N_2872,N_2944);
xor U3228 (N_3228,N_2770,N_2882);
nor U3229 (N_3229,N_2774,N_2932);
and U3230 (N_3230,N_2950,N_2824);
xor U3231 (N_3231,N_2989,N_2894);
xor U3232 (N_3232,N_2965,N_2959);
or U3233 (N_3233,N_2989,N_2754);
nand U3234 (N_3234,N_2899,N_2910);
or U3235 (N_3235,N_2800,N_2871);
xor U3236 (N_3236,N_2906,N_2796);
and U3237 (N_3237,N_2974,N_2837);
and U3238 (N_3238,N_2780,N_2890);
nand U3239 (N_3239,N_2982,N_2878);
or U3240 (N_3240,N_2942,N_2892);
and U3241 (N_3241,N_2872,N_2850);
and U3242 (N_3242,N_2981,N_2906);
or U3243 (N_3243,N_2990,N_2769);
nand U3244 (N_3244,N_2990,N_2824);
nand U3245 (N_3245,N_2989,N_2801);
or U3246 (N_3246,N_2882,N_2983);
nand U3247 (N_3247,N_2769,N_2859);
nand U3248 (N_3248,N_2807,N_2863);
nor U3249 (N_3249,N_2842,N_2996);
xnor U3250 (N_3250,N_3232,N_3068);
or U3251 (N_3251,N_3092,N_3146);
nor U3252 (N_3252,N_3094,N_3016);
or U3253 (N_3253,N_3187,N_3162);
nor U3254 (N_3254,N_3130,N_3243);
and U3255 (N_3255,N_3037,N_3085);
and U3256 (N_3256,N_3116,N_3181);
nor U3257 (N_3257,N_3239,N_3125);
xnor U3258 (N_3258,N_3129,N_3168);
or U3259 (N_3259,N_3020,N_3179);
and U3260 (N_3260,N_3060,N_3190);
nor U3261 (N_3261,N_3107,N_3026);
nor U3262 (N_3262,N_3200,N_3199);
and U3263 (N_3263,N_3046,N_3227);
or U3264 (N_3264,N_3230,N_3045);
nand U3265 (N_3265,N_3233,N_3214);
or U3266 (N_3266,N_3089,N_3196);
xor U3267 (N_3267,N_3122,N_3029);
nor U3268 (N_3268,N_3154,N_3110);
nor U3269 (N_3269,N_3184,N_3015);
nor U3270 (N_3270,N_3101,N_3215);
or U3271 (N_3271,N_3198,N_3071);
and U3272 (N_3272,N_3013,N_3160);
nand U3273 (N_3273,N_3035,N_3242);
nand U3274 (N_3274,N_3102,N_3176);
or U3275 (N_3275,N_3072,N_3065);
nor U3276 (N_3276,N_3147,N_3103);
or U3277 (N_3277,N_3053,N_3202);
and U3278 (N_3278,N_3174,N_3024);
and U3279 (N_3279,N_3106,N_3022);
and U3280 (N_3280,N_3100,N_3134);
nor U3281 (N_3281,N_3157,N_3010);
or U3282 (N_3282,N_3124,N_3237);
nand U3283 (N_3283,N_3007,N_3169);
nand U3284 (N_3284,N_3098,N_3170);
nor U3285 (N_3285,N_3021,N_3240);
and U3286 (N_3286,N_3248,N_3104);
xor U3287 (N_3287,N_3244,N_3178);
xor U3288 (N_3288,N_3114,N_3152);
or U3289 (N_3289,N_3051,N_3220);
and U3290 (N_3290,N_3188,N_3058);
and U3291 (N_3291,N_3142,N_3027);
nor U3292 (N_3292,N_3088,N_3025);
xnor U3293 (N_3293,N_3002,N_3245);
and U3294 (N_3294,N_3216,N_3062);
and U3295 (N_3295,N_3135,N_3166);
nor U3296 (N_3296,N_3090,N_3226);
nand U3297 (N_3297,N_3086,N_3042);
nor U3298 (N_3298,N_3039,N_3212);
nor U3299 (N_3299,N_3224,N_3066);
nand U3300 (N_3300,N_3077,N_3004);
nor U3301 (N_3301,N_3121,N_3141);
or U3302 (N_3302,N_3186,N_3052);
xor U3303 (N_3303,N_3145,N_3011);
or U3304 (N_3304,N_3050,N_3218);
nor U3305 (N_3305,N_3209,N_3204);
nor U3306 (N_3306,N_3189,N_3056);
and U3307 (N_3307,N_3126,N_3097);
nand U3308 (N_3308,N_3222,N_3017);
xor U3309 (N_3309,N_3109,N_3192);
or U3310 (N_3310,N_3070,N_3185);
nor U3311 (N_3311,N_3118,N_3000);
nor U3312 (N_3312,N_3005,N_3207);
nand U3313 (N_3313,N_3069,N_3064);
or U3314 (N_3314,N_3193,N_3028);
nor U3315 (N_3315,N_3228,N_3213);
xnor U3316 (N_3316,N_3140,N_3123);
nor U3317 (N_3317,N_3177,N_3009);
nand U3318 (N_3318,N_3210,N_3076);
nor U3319 (N_3319,N_3012,N_3034);
nor U3320 (N_3320,N_3083,N_3019);
or U3321 (N_3321,N_3164,N_3229);
nand U3322 (N_3322,N_3084,N_3172);
and U3323 (N_3323,N_3074,N_3047);
nor U3324 (N_3324,N_3105,N_3238);
or U3325 (N_3325,N_3055,N_3151);
nand U3326 (N_3326,N_3115,N_3246);
or U3327 (N_3327,N_3119,N_3030);
nor U3328 (N_3328,N_3149,N_3175);
and U3329 (N_3329,N_3113,N_3099);
nor U3330 (N_3330,N_3137,N_3194);
or U3331 (N_3331,N_3111,N_3023);
nor U3332 (N_3332,N_3096,N_3225);
nand U3333 (N_3333,N_3031,N_3082);
or U3334 (N_3334,N_3195,N_3234);
xnor U3335 (N_3335,N_3033,N_3048);
nor U3336 (N_3336,N_3041,N_3078);
nor U3337 (N_3337,N_3138,N_3156);
xor U3338 (N_3338,N_3143,N_3075);
or U3339 (N_3339,N_3127,N_3036);
or U3340 (N_3340,N_3003,N_3095);
or U3341 (N_3341,N_3159,N_3108);
xnor U3342 (N_3342,N_3236,N_3008);
and U3343 (N_3343,N_3014,N_3206);
xnor U3344 (N_3344,N_3038,N_3093);
nand U3345 (N_3345,N_3128,N_3067);
or U3346 (N_3346,N_3201,N_3136);
or U3347 (N_3347,N_3120,N_3191);
or U3348 (N_3348,N_3081,N_3043);
or U3349 (N_3349,N_3054,N_3148);
and U3350 (N_3350,N_3219,N_3247);
xnor U3351 (N_3351,N_3079,N_3049);
or U3352 (N_3352,N_3063,N_3167);
xor U3353 (N_3353,N_3180,N_3006);
and U3354 (N_3354,N_3150,N_3087);
xor U3355 (N_3355,N_3018,N_3158);
nor U3356 (N_3356,N_3155,N_3211);
nand U3357 (N_3357,N_3059,N_3040);
or U3358 (N_3358,N_3032,N_3205);
nand U3359 (N_3359,N_3112,N_3163);
or U3360 (N_3360,N_3182,N_3249);
nor U3361 (N_3361,N_3001,N_3165);
xnor U3362 (N_3362,N_3153,N_3132);
nand U3363 (N_3363,N_3171,N_3131);
nand U3364 (N_3364,N_3080,N_3203);
or U3365 (N_3365,N_3217,N_3173);
nand U3366 (N_3366,N_3117,N_3061);
or U3367 (N_3367,N_3241,N_3161);
xnor U3368 (N_3368,N_3073,N_3044);
xnor U3369 (N_3369,N_3091,N_3057);
nor U3370 (N_3370,N_3208,N_3235);
or U3371 (N_3371,N_3221,N_3139);
nor U3372 (N_3372,N_3133,N_3197);
nand U3373 (N_3373,N_3223,N_3231);
nand U3374 (N_3374,N_3144,N_3183);
xor U3375 (N_3375,N_3138,N_3172);
and U3376 (N_3376,N_3046,N_3140);
nor U3377 (N_3377,N_3214,N_3195);
or U3378 (N_3378,N_3239,N_3080);
or U3379 (N_3379,N_3100,N_3198);
and U3380 (N_3380,N_3221,N_3069);
nor U3381 (N_3381,N_3185,N_3170);
nor U3382 (N_3382,N_3020,N_3125);
or U3383 (N_3383,N_3057,N_3061);
nand U3384 (N_3384,N_3236,N_3048);
or U3385 (N_3385,N_3055,N_3196);
xor U3386 (N_3386,N_3093,N_3067);
xnor U3387 (N_3387,N_3106,N_3118);
nor U3388 (N_3388,N_3235,N_3070);
nand U3389 (N_3389,N_3173,N_3153);
and U3390 (N_3390,N_3000,N_3154);
and U3391 (N_3391,N_3025,N_3170);
xor U3392 (N_3392,N_3151,N_3105);
xnor U3393 (N_3393,N_3229,N_3198);
or U3394 (N_3394,N_3073,N_3011);
nor U3395 (N_3395,N_3113,N_3244);
nand U3396 (N_3396,N_3172,N_3249);
xnor U3397 (N_3397,N_3033,N_3246);
xor U3398 (N_3398,N_3239,N_3174);
nand U3399 (N_3399,N_3243,N_3242);
nor U3400 (N_3400,N_3013,N_3190);
nand U3401 (N_3401,N_3193,N_3032);
xor U3402 (N_3402,N_3077,N_3222);
and U3403 (N_3403,N_3164,N_3134);
nand U3404 (N_3404,N_3215,N_3097);
nand U3405 (N_3405,N_3071,N_3145);
or U3406 (N_3406,N_3125,N_3150);
nand U3407 (N_3407,N_3022,N_3023);
nand U3408 (N_3408,N_3140,N_3168);
nand U3409 (N_3409,N_3189,N_3238);
xnor U3410 (N_3410,N_3181,N_3008);
xor U3411 (N_3411,N_3211,N_3036);
and U3412 (N_3412,N_3053,N_3013);
xor U3413 (N_3413,N_3185,N_3080);
xor U3414 (N_3414,N_3025,N_3205);
nor U3415 (N_3415,N_3178,N_3029);
xnor U3416 (N_3416,N_3180,N_3244);
xor U3417 (N_3417,N_3124,N_3139);
nor U3418 (N_3418,N_3092,N_3175);
xor U3419 (N_3419,N_3176,N_3239);
xor U3420 (N_3420,N_3043,N_3229);
nor U3421 (N_3421,N_3226,N_3118);
xnor U3422 (N_3422,N_3179,N_3248);
xnor U3423 (N_3423,N_3190,N_3147);
nand U3424 (N_3424,N_3235,N_3047);
nand U3425 (N_3425,N_3246,N_3176);
nor U3426 (N_3426,N_3154,N_3218);
nand U3427 (N_3427,N_3060,N_3077);
and U3428 (N_3428,N_3242,N_3227);
xnor U3429 (N_3429,N_3041,N_3163);
or U3430 (N_3430,N_3071,N_3245);
nand U3431 (N_3431,N_3100,N_3168);
nand U3432 (N_3432,N_3129,N_3131);
nor U3433 (N_3433,N_3156,N_3152);
or U3434 (N_3434,N_3141,N_3166);
nand U3435 (N_3435,N_3055,N_3197);
nor U3436 (N_3436,N_3102,N_3198);
nor U3437 (N_3437,N_3159,N_3002);
nor U3438 (N_3438,N_3226,N_3015);
xnor U3439 (N_3439,N_3063,N_3117);
or U3440 (N_3440,N_3240,N_3029);
or U3441 (N_3441,N_3137,N_3161);
nor U3442 (N_3442,N_3199,N_3078);
nor U3443 (N_3443,N_3006,N_3172);
xnor U3444 (N_3444,N_3100,N_3060);
and U3445 (N_3445,N_3224,N_3182);
and U3446 (N_3446,N_3008,N_3095);
nand U3447 (N_3447,N_3050,N_3097);
and U3448 (N_3448,N_3060,N_3019);
nand U3449 (N_3449,N_3094,N_3042);
or U3450 (N_3450,N_3234,N_3184);
xor U3451 (N_3451,N_3232,N_3082);
or U3452 (N_3452,N_3039,N_3037);
xnor U3453 (N_3453,N_3088,N_3154);
xnor U3454 (N_3454,N_3049,N_3102);
nand U3455 (N_3455,N_3030,N_3146);
or U3456 (N_3456,N_3218,N_3011);
nand U3457 (N_3457,N_3065,N_3122);
and U3458 (N_3458,N_3178,N_3184);
and U3459 (N_3459,N_3001,N_3063);
nor U3460 (N_3460,N_3150,N_3037);
nand U3461 (N_3461,N_3224,N_3188);
and U3462 (N_3462,N_3097,N_3018);
nor U3463 (N_3463,N_3179,N_3225);
xor U3464 (N_3464,N_3160,N_3204);
xnor U3465 (N_3465,N_3241,N_3090);
nand U3466 (N_3466,N_3016,N_3050);
nor U3467 (N_3467,N_3016,N_3198);
or U3468 (N_3468,N_3026,N_3061);
xnor U3469 (N_3469,N_3195,N_3156);
nand U3470 (N_3470,N_3183,N_3193);
or U3471 (N_3471,N_3106,N_3197);
xor U3472 (N_3472,N_3249,N_3020);
or U3473 (N_3473,N_3021,N_3131);
or U3474 (N_3474,N_3116,N_3138);
or U3475 (N_3475,N_3238,N_3201);
nor U3476 (N_3476,N_3066,N_3109);
and U3477 (N_3477,N_3185,N_3050);
nor U3478 (N_3478,N_3193,N_3194);
xnor U3479 (N_3479,N_3140,N_3047);
nand U3480 (N_3480,N_3086,N_3049);
nor U3481 (N_3481,N_3089,N_3221);
nor U3482 (N_3482,N_3128,N_3003);
and U3483 (N_3483,N_3167,N_3124);
nand U3484 (N_3484,N_3193,N_3085);
or U3485 (N_3485,N_3051,N_3224);
xor U3486 (N_3486,N_3080,N_3044);
xnor U3487 (N_3487,N_3126,N_3069);
xnor U3488 (N_3488,N_3183,N_3168);
nand U3489 (N_3489,N_3213,N_3081);
and U3490 (N_3490,N_3113,N_3163);
or U3491 (N_3491,N_3014,N_3136);
and U3492 (N_3492,N_3072,N_3157);
nor U3493 (N_3493,N_3003,N_3245);
nor U3494 (N_3494,N_3082,N_3074);
xor U3495 (N_3495,N_3191,N_3065);
or U3496 (N_3496,N_3177,N_3011);
xor U3497 (N_3497,N_3128,N_3219);
nand U3498 (N_3498,N_3012,N_3021);
or U3499 (N_3499,N_3055,N_3165);
nor U3500 (N_3500,N_3491,N_3397);
nand U3501 (N_3501,N_3366,N_3436);
nand U3502 (N_3502,N_3254,N_3403);
xnor U3503 (N_3503,N_3431,N_3466);
xor U3504 (N_3504,N_3418,N_3396);
and U3505 (N_3505,N_3393,N_3359);
and U3506 (N_3506,N_3377,N_3442);
nand U3507 (N_3507,N_3482,N_3262);
or U3508 (N_3508,N_3319,N_3405);
xor U3509 (N_3509,N_3429,N_3352);
and U3510 (N_3510,N_3361,N_3327);
and U3511 (N_3511,N_3392,N_3499);
nor U3512 (N_3512,N_3363,N_3287);
nor U3513 (N_3513,N_3350,N_3326);
or U3514 (N_3514,N_3268,N_3416);
nor U3515 (N_3515,N_3400,N_3290);
nor U3516 (N_3516,N_3465,N_3496);
or U3517 (N_3517,N_3401,N_3269);
or U3518 (N_3518,N_3395,N_3309);
xnor U3519 (N_3519,N_3272,N_3425);
or U3520 (N_3520,N_3468,N_3479);
nor U3521 (N_3521,N_3320,N_3369);
nand U3522 (N_3522,N_3475,N_3489);
nand U3523 (N_3523,N_3376,N_3312);
and U3524 (N_3524,N_3478,N_3256);
nand U3525 (N_3525,N_3346,N_3306);
nor U3526 (N_3526,N_3286,N_3345);
or U3527 (N_3527,N_3329,N_3297);
or U3528 (N_3528,N_3318,N_3258);
or U3529 (N_3529,N_3337,N_3427);
nor U3530 (N_3530,N_3263,N_3411);
and U3531 (N_3531,N_3467,N_3276);
and U3532 (N_3532,N_3282,N_3448);
nor U3533 (N_3533,N_3494,N_3382);
xor U3534 (N_3534,N_3351,N_3455);
nor U3535 (N_3535,N_3460,N_3347);
or U3536 (N_3536,N_3307,N_3449);
nor U3537 (N_3537,N_3445,N_3493);
or U3538 (N_3538,N_3324,N_3378);
nand U3539 (N_3539,N_3295,N_3332);
or U3540 (N_3540,N_3275,N_3355);
nor U3541 (N_3541,N_3298,N_3338);
or U3542 (N_3542,N_3349,N_3438);
and U3543 (N_3543,N_3474,N_3291);
nor U3544 (N_3544,N_3495,N_3278);
or U3545 (N_3545,N_3390,N_3341);
or U3546 (N_3546,N_3348,N_3267);
xor U3547 (N_3547,N_3296,N_3308);
nor U3548 (N_3548,N_3457,N_3339);
and U3549 (N_3549,N_3261,N_3406);
nor U3550 (N_3550,N_3492,N_3409);
and U3551 (N_3551,N_3452,N_3367);
nand U3552 (N_3552,N_3321,N_3333);
or U3553 (N_3553,N_3381,N_3335);
or U3554 (N_3554,N_3444,N_3266);
or U3555 (N_3555,N_3440,N_3432);
xor U3556 (N_3556,N_3292,N_3343);
nor U3557 (N_3557,N_3370,N_3404);
or U3558 (N_3558,N_3463,N_3430);
xor U3559 (N_3559,N_3328,N_3402);
and U3560 (N_3560,N_3435,N_3316);
nor U3561 (N_3561,N_3477,N_3446);
xnor U3562 (N_3562,N_3487,N_3357);
or U3563 (N_3563,N_3423,N_3305);
xor U3564 (N_3564,N_3301,N_3277);
xnor U3565 (N_3565,N_3399,N_3454);
xor U3566 (N_3566,N_3451,N_3274);
nor U3567 (N_3567,N_3424,N_3322);
and U3568 (N_3568,N_3310,N_3375);
nor U3569 (N_3569,N_3471,N_3385);
nand U3570 (N_3570,N_3304,N_3336);
nor U3571 (N_3571,N_3250,N_3302);
or U3572 (N_3572,N_3437,N_3255);
nor U3573 (N_3573,N_3314,N_3472);
or U3574 (N_3574,N_3365,N_3284);
nand U3575 (N_3575,N_3421,N_3485);
or U3576 (N_3576,N_3371,N_3426);
xor U3577 (N_3577,N_3453,N_3265);
nand U3578 (N_3578,N_3356,N_3360);
xor U3579 (N_3579,N_3389,N_3353);
nor U3580 (N_3580,N_3280,N_3270);
or U3581 (N_3581,N_3422,N_3264);
nor U3582 (N_3582,N_3315,N_3481);
and U3583 (N_3583,N_3374,N_3368);
and U3584 (N_3584,N_3384,N_3317);
nor U3585 (N_3585,N_3344,N_3294);
and U3586 (N_3586,N_3461,N_3259);
xor U3587 (N_3587,N_3413,N_3383);
nor U3588 (N_3588,N_3407,N_3412);
nor U3589 (N_3589,N_3260,N_3470);
xor U3590 (N_3590,N_3334,N_3289);
and U3591 (N_3591,N_3288,N_3380);
xnor U3592 (N_3592,N_3462,N_3490);
and U3593 (N_3593,N_3379,N_3441);
nor U3594 (N_3594,N_3443,N_3313);
or U3595 (N_3595,N_3498,N_3303);
and U3596 (N_3596,N_3299,N_3386);
xor U3597 (N_3597,N_3387,N_3331);
xor U3598 (N_3598,N_3464,N_3257);
or U3599 (N_3599,N_3330,N_3293);
nand U3600 (N_3600,N_3388,N_3279);
and U3601 (N_3601,N_3372,N_3488);
nand U3602 (N_3602,N_3325,N_3285);
nand U3603 (N_3603,N_3476,N_3251);
and U3604 (N_3604,N_3323,N_3458);
nand U3605 (N_3605,N_3300,N_3354);
nor U3606 (N_3606,N_3450,N_3311);
nor U3607 (N_3607,N_3364,N_3391);
and U3608 (N_3608,N_3340,N_3281);
nor U3609 (N_3609,N_3253,N_3486);
or U3610 (N_3610,N_3469,N_3271);
nand U3611 (N_3611,N_3497,N_3408);
and U3612 (N_3612,N_3428,N_3252);
nor U3613 (N_3613,N_3439,N_3420);
nand U3614 (N_3614,N_3484,N_3447);
nor U3615 (N_3615,N_3373,N_3394);
and U3616 (N_3616,N_3419,N_3283);
nor U3617 (N_3617,N_3414,N_3410);
nor U3618 (N_3618,N_3459,N_3456);
and U3619 (N_3619,N_3415,N_3480);
nor U3620 (N_3620,N_3362,N_3483);
nand U3621 (N_3621,N_3417,N_3433);
nor U3622 (N_3622,N_3358,N_3273);
nand U3623 (N_3623,N_3473,N_3434);
xnor U3624 (N_3624,N_3342,N_3398);
or U3625 (N_3625,N_3386,N_3360);
nor U3626 (N_3626,N_3321,N_3308);
or U3627 (N_3627,N_3390,N_3489);
nor U3628 (N_3628,N_3441,N_3389);
xnor U3629 (N_3629,N_3428,N_3387);
or U3630 (N_3630,N_3317,N_3329);
or U3631 (N_3631,N_3467,N_3457);
or U3632 (N_3632,N_3448,N_3313);
and U3633 (N_3633,N_3264,N_3312);
nand U3634 (N_3634,N_3280,N_3493);
nor U3635 (N_3635,N_3453,N_3251);
nor U3636 (N_3636,N_3299,N_3402);
xor U3637 (N_3637,N_3284,N_3374);
nand U3638 (N_3638,N_3433,N_3399);
nand U3639 (N_3639,N_3456,N_3253);
nand U3640 (N_3640,N_3381,N_3471);
and U3641 (N_3641,N_3454,N_3357);
xnor U3642 (N_3642,N_3478,N_3366);
nor U3643 (N_3643,N_3319,N_3371);
or U3644 (N_3644,N_3423,N_3425);
nor U3645 (N_3645,N_3406,N_3336);
xnor U3646 (N_3646,N_3413,N_3338);
nand U3647 (N_3647,N_3352,N_3338);
or U3648 (N_3648,N_3448,N_3260);
or U3649 (N_3649,N_3389,N_3341);
xnor U3650 (N_3650,N_3323,N_3282);
or U3651 (N_3651,N_3466,N_3420);
xnor U3652 (N_3652,N_3475,N_3324);
nor U3653 (N_3653,N_3448,N_3478);
and U3654 (N_3654,N_3348,N_3289);
xnor U3655 (N_3655,N_3310,N_3305);
xor U3656 (N_3656,N_3487,N_3347);
nor U3657 (N_3657,N_3416,N_3289);
nand U3658 (N_3658,N_3303,N_3400);
xor U3659 (N_3659,N_3255,N_3271);
xnor U3660 (N_3660,N_3384,N_3329);
xor U3661 (N_3661,N_3472,N_3392);
and U3662 (N_3662,N_3311,N_3431);
and U3663 (N_3663,N_3345,N_3259);
nor U3664 (N_3664,N_3273,N_3330);
or U3665 (N_3665,N_3311,N_3366);
nor U3666 (N_3666,N_3362,N_3400);
or U3667 (N_3667,N_3417,N_3261);
and U3668 (N_3668,N_3413,N_3378);
xnor U3669 (N_3669,N_3301,N_3360);
or U3670 (N_3670,N_3359,N_3312);
xor U3671 (N_3671,N_3371,N_3254);
nor U3672 (N_3672,N_3304,N_3480);
or U3673 (N_3673,N_3324,N_3369);
xor U3674 (N_3674,N_3328,N_3488);
xor U3675 (N_3675,N_3349,N_3472);
or U3676 (N_3676,N_3448,N_3284);
and U3677 (N_3677,N_3480,N_3402);
or U3678 (N_3678,N_3351,N_3472);
and U3679 (N_3679,N_3341,N_3374);
xor U3680 (N_3680,N_3367,N_3322);
and U3681 (N_3681,N_3290,N_3433);
nand U3682 (N_3682,N_3446,N_3259);
nor U3683 (N_3683,N_3496,N_3395);
and U3684 (N_3684,N_3450,N_3422);
xor U3685 (N_3685,N_3438,N_3277);
and U3686 (N_3686,N_3316,N_3298);
and U3687 (N_3687,N_3251,N_3429);
or U3688 (N_3688,N_3442,N_3457);
xor U3689 (N_3689,N_3384,N_3318);
or U3690 (N_3690,N_3480,N_3498);
nor U3691 (N_3691,N_3488,N_3423);
xor U3692 (N_3692,N_3400,N_3413);
nand U3693 (N_3693,N_3296,N_3343);
nand U3694 (N_3694,N_3429,N_3303);
and U3695 (N_3695,N_3400,N_3274);
nor U3696 (N_3696,N_3392,N_3387);
or U3697 (N_3697,N_3275,N_3438);
nand U3698 (N_3698,N_3278,N_3465);
or U3699 (N_3699,N_3427,N_3409);
nor U3700 (N_3700,N_3474,N_3396);
and U3701 (N_3701,N_3457,N_3316);
xnor U3702 (N_3702,N_3301,N_3365);
or U3703 (N_3703,N_3382,N_3418);
xnor U3704 (N_3704,N_3327,N_3291);
or U3705 (N_3705,N_3449,N_3468);
and U3706 (N_3706,N_3375,N_3377);
nor U3707 (N_3707,N_3476,N_3433);
or U3708 (N_3708,N_3418,N_3370);
nor U3709 (N_3709,N_3443,N_3463);
nand U3710 (N_3710,N_3361,N_3316);
xor U3711 (N_3711,N_3260,N_3353);
nand U3712 (N_3712,N_3355,N_3390);
or U3713 (N_3713,N_3345,N_3292);
nor U3714 (N_3714,N_3350,N_3292);
and U3715 (N_3715,N_3344,N_3452);
or U3716 (N_3716,N_3448,N_3343);
and U3717 (N_3717,N_3428,N_3276);
nand U3718 (N_3718,N_3437,N_3335);
nor U3719 (N_3719,N_3409,N_3414);
and U3720 (N_3720,N_3495,N_3306);
or U3721 (N_3721,N_3329,N_3350);
nand U3722 (N_3722,N_3289,N_3325);
nor U3723 (N_3723,N_3415,N_3458);
xnor U3724 (N_3724,N_3442,N_3428);
xor U3725 (N_3725,N_3446,N_3400);
nand U3726 (N_3726,N_3423,N_3445);
or U3727 (N_3727,N_3336,N_3369);
xor U3728 (N_3728,N_3455,N_3272);
nand U3729 (N_3729,N_3453,N_3318);
and U3730 (N_3730,N_3258,N_3410);
nand U3731 (N_3731,N_3487,N_3419);
xor U3732 (N_3732,N_3368,N_3286);
nor U3733 (N_3733,N_3301,N_3495);
nor U3734 (N_3734,N_3429,N_3445);
nor U3735 (N_3735,N_3305,N_3455);
nand U3736 (N_3736,N_3409,N_3257);
nand U3737 (N_3737,N_3286,N_3252);
xor U3738 (N_3738,N_3416,N_3365);
or U3739 (N_3739,N_3493,N_3258);
or U3740 (N_3740,N_3447,N_3481);
xnor U3741 (N_3741,N_3365,N_3392);
and U3742 (N_3742,N_3489,N_3494);
or U3743 (N_3743,N_3473,N_3297);
nand U3744 (N_3744,N_3291,N_3315);
and U3745 (N_3745,N_3347,N_3386);
and U3746 (N_3746,N_3390,N_3441);
xnor U3747 (N_3747,N_3421,N_3338);
nand U3748 (N_3748,N_3486,N_3414);
nor U3749 (N_3749,N_3281,N_3375);
nand U3750 (N_3750,N_3599,N_3705);
or U3751 (N_3751,N_3540,N_3575);
xor U3752 (N_3752,N_3632,N_3678);
nor U3753 (N_3753,N_3604,N_3512);
or U3754 (N_3754,N_3694,N_3552);
nand U3755 (N_3755,N_3697,N_3610);
or U3756 (N_3756,N_3631,N_3740);
nand U3757 (N_3757,N_3651,N_3531);
nand U3758 (N_3758,N_3502,N_3505);
nor U3759 (N_3759,N_3749,N_3707);
nand U3760 (N_3760,N_3623,N_3588);
xor U3761 (N_3761,N_3544,N_3656);
xnor U3762 (N_3762,N_3548,N_3523);
nand U3763 (N_3763,N_3521,N_3676);
nor U3764 (N_3764,N_3723,N_3695);
nor U3765 (N_3765,N_3519,N_3533);
nor U3766 (N_3766,N_3539,N_3731);
and U3767 (N_3767,N_3592,N_3681);
xnor U3768 (N_3768,N_3609,N_3672);
nor U3769 (N_3769,N_3606,N_3549);
nand U3770 (N_3770,N_3598,N_3503);
and U3771 (N_3771,N_3542,N_3581);
and U3772 (N_3772,N_3657,N_3641);
xor U3773 (N_3773,N_3711,N_3737);
or U3774 (N_3774,N_3579,N_3665);
nor U3775 (N_3775,N_3600,N_3666);
or U3776 (N_3776,N_3674,N_3617);
or U3777 (N_3777,N_3593,N_3710);
or U3778 (N_3778,N_3667,N_3659);
and U3779 (N_3779,N_3650,N_3625);
or U3780 (N_3780,N_3716,N_3547);
xor U3781 (N_3781,N_3508,N_3722);
nor U3782 (N_3782,N_3560,N_3693);
xor U3783 (N_3783,N_3607,N_3529);
nand U3784 (N_3784,N_3597,N_3574);
and U3785 (N_3785,N_3639,N_3712);
xnor U3786 (N_3786,N_3648,N_3511);
nor U3787 (N_3787,N_3743,N_3701);
nand U3788 (N_3788,N_3534,N_3562);
and U3789 (N_3789,N_3718,N_3526);
and U3790 (N_3790,N_3727,N_3500);
nand U3791 (N_3791,N_3515,N_3528);
nor U3792 (N_3792,N_3668,N_3611);
xor U3793 (N_3793,N_3742,N_3570);
nand U3794 (N_3794,N_3647,N_3628);
nor U3795 (N_3795,N_3567,N_3514);
nand U3796 (N_3796,N_3585,N_3596);
or U3797 (N_3797,N_3662,N_3688);
nor U3798 (N_3798,N_3522,N_3642);
nand U3799 (N_3799,N_3565,N_3527);
xnor U3800 (N_3800,N_3538,N_3590);
nor U3801 (N_3801,N_3714,N_3734);
and U3802 (N_3802,N_3653,N_3728);
xnor U3803 (N_3803,N_3564,N_3633);
or U3804 (N_3804,N_3645,N_3739);
nor U3805 (N_3805,N_3556,N_3660);
xor U3806 (N_3806,N_3735,N_3664);
and U3807 (N_3807,N_3572,N_3715);
nand U3808 (N_3808,N_3510,N_3725);
or U3809 (N_3809,N_3732,N_3525);
xnor U3810 (N_3810,N_3577,N_3551);
xor U3811 (N_3811,N_3680,N_3702);
nand U3812 (N_3812,N_3569,N_3613);
xor U3813 (N_3813,N_3608,N_3685);
xnor U3814 (N_3814,N_3677,N_3586);
or U3815 (N_3815,N_3626,N_3741);
nor U3816 (N_3816,N_3594,N_3669);
nor U3817 (N_3817,N_3602,N_3524);
xor U3818 (N_3818,N_3584,N_3673);
nor U3819 (N_3819,N_3566,N_3646);
or U3820 (N_3820,N_3640,N_3553);
or U3821 (N_3821,N_3615,N_3605);
nor U3822 (N_3822,N_3699,N_3745);
or U3823 (N_3823,N_3720,N_3627);
or U3824 (N_3824,N_3535,N_3516);
nand U3825 (N_3825,N_3689,N_3638);
xor U3826 (N_3826,N_3679,N_3671);
xor U3827 (N_3827,N_3541,N_3643);
or U3828 (N_3828,N_3675,N_3746);
xnor U3829 (N_3829,N_3655,N_3603);
xnor U3830 (N_3830,N_3618,N_3545);
nor U3831 (N_3831,N_3644,N_3621);
and U3832 (N_3832,N_3687,N_3703);
and U3833 (N_3833,N_3736,N_3558);
and U3834 (N_3834,N_3690,N_3612);
nand U3835 (N_3835,N_3559,N_3520);
nor U3836 (N_3836,N_3563,N_3738);
or U3837 (N_3837,N_3748,N_3698);
or U3838 (N_3838,N_3747,N_3561);
or U3839 (N_3839,N_3704,N_3652);
and U3840 (N_3840,N_3719,N_3637);
nand U3841 (N_3841,N_3724,N_3580);
or U3842 (N_3842,N_3717,N_3587);
or U3843 (N_3843,N_3730,N_3616);
nor U3844 (N_3844,N_3543,N_3663);
nand U3845 (N_3845,N_3635,N_3591);
nor U3846 (N_3846,N_3634,N_3557);
nor U3847 (N_3847,N_3683,N_3509);
or U3848 (N_3848,N_3729,N_3555);
nor U3849 (N_3849,N_3582,N_3532);
and U3850 (N_3850,N_3501,N_3589);
nor U3851 (N_3851,N_3622,N_3517);
and U3852 (N_3852,N_3661,N_3571);
nand U3853 (N_3853,N_3658,N_3709);
or U3854 (N_3854,N_3682,N_3696);
and U3855 (N_3855,N_3504,N_3726);
xor U3856 (N_3856,N_3654,N_3583);
or U3857 (N_3857,N_3686,N_3624);
nor U3858 (N_3858,N_3629,N_3636);
or U3859 (N_3859,N_3700,N_3513);
or U3860 (N_3860,N_3573,N_3713);
or U3861 (N_3861,N_3530,N_3578);
nand U3862 (N_3862,N_3550,N_3630);
nand U3863 (N_3863,N_3536,N_3649);
nand U3864 (N_3864,N_3733,N_3620);
nor U3865 (N_3865,N_3706,N_3684);
and U3866 (N_3866,N_3744,N_3601);
and U3867 (N_3867,N_3568,N_3692);
nor U3868 (N_3868,N_3576,N_3670);
and U3869 (N_3869,N_3595,N_3619);
and U3870 (N_3870,N_3506,N_3507);
xnor U3871 (N_3871,N_3614,N_3537);
and U3872 (N_3872,N_3721,N_3708);
nor U3873 (N_3873,N_3546,N_3691);
nand U3874 (N_3874,N_3554,N_3518);
nand U3875 (N_3875,N_3684,N_3511);
or U3876 (N_3876,N_3539,N_3621);
and U3877 (N_3877,N_3566,N_3553);
nand U3878 (N_3878,N_3723,N_3670);
xor U3879 (N_3879,N_3607,N_3543);
and U3880 (N_3880,N_3747,N_3683);
or U3881 (N_3881,N_3511,N_3537);
or U3882 (N_3882,N_3629,N_3706);
and U3883 (N_3883,N_3509,N_3679);
or U3884 (N_3884,N_3525,N_3541);
or U3885 (N_3885,N_3633,N_3551);
nor U3886 (N_3886,N_3646,N_3677);
and U3887 (N_3887,N_3610,N_3578);
nor U3888 (N_3888,N_3560,N_3679);
nor U3889 (N_3889,N_3604,N_3736);
and U3890 (N_3890,N_3641,N_3610);
or U3891 (N_3891,N_3645,N_3713);
and U3892 (N_3892,N_3747,N_3529);
or U3893 (N_3893,N_3511,N_3524);
nand U3894 (N_3894,N_3537,N_3562);
or U3895 (N_3895,N_3636,N_3646);
and U3896 (N_3896,N_3594,N_3619);
nor U3897 (N_3897,N_3679,N_3506);
xor U3898 (N_3898,N_3543,N_3684);
and U3899 (N_3899,N_3513,N_3721);
nand U3900 (N_3900,N_3536,N_3553);
nand U3901 (N_3901,N_3521,N_3715);
xor U3902 (N_3902,N_3640,N_3720);
and U3903 (N_3903,N_3690,N_3501);
xor U3904 (N_3904,N_3639,N_3692);
nand U3905 (N_3905,N_3561,N_3501);
and U3906 (N_3906,N_3568,N_3506);
nand U3907 (N_3907,N_3646,N_3569);
or U3908 (N_3908,N_3663,N_3590);
nor U3909 (N_3909,N_3659,N_3742);
xor U3910 (N_3910,N_3670,N_3583);
nor U3911 (N_3911,N_3582,N_3655);
nor U3912 (N_3912,N_3556,N_3662);
and U3913 (N_3913,N_3504,N_3558);
nor U3914 (N_3914,N_3531,N_3594);
xnor U3915 (N_3915,N_3732,N_3579);
or U3916 (N_3916,N_3587,N_3652);
nand U3917 (N_3917,N_3555,N_3504);
nor U3918 (N_3918,N_3676,N_3523);
nor U3919 (N_3919,N_3672,N_3528);
and U3920 (N_3920,N_3523,N_3738);
and U3921 (N_3921,N_3673,N_3724);
and U3922 (N_3922,N_3736,N_3667);
nor U3923 (N_3923,N_3572,N_3622);
nor U3924 (N_3924,N_3609,N_3547);
and U3925 (N_3925,N_3539,N_3597);
nor U3926 (N_3926,N_3559,N_3731);
or U3927 (N_3927,N_3514,N_3579);
and U3928 (N_3928,N_3682,N_3735);
or U3929 (N_3929,N_3501,N_3697);
nor U3930 (N_3930,N_3650,N_3532);
or U3931 (N_3931,N_3526,N_3512);
and U3932 (N_3932,N_3510,N_3500);
nor U3933 (N_3933,N_3631,N_3587);
xor U3934 (N_3934,N_3730,N_3635);
nand U3935 (N_3935,N_3572,N_3671);
or U3936 (N_3936,N_3697,N_3504);
nand U3937 (N_3937,N_3713,N_3620);
and U3938 (N_3938,N_3641,N_3704);
xnor U3939 (N_3939,N_3548,N_3570);
and U3940 (N_3940,N_3726,N_3526);
xnor U3941 (N_3941,N_3721,N_3537);
or U3942 (N_3942,N_3672,N_3682);
or U3943 (N_3943,N_3563,N_3548);
or U3944 (N_3944,N_3540,N_3598);
or U3945 (N_3945,N_3576,N_3683);
nand U3946 (N_3946,N_3674,N_3549);
nor U3947 (N_3947,N_3589,N_3648);
or U3948 (N_3948,N_3546,N_3526);
and U3949 (N_3949,N_3641,N_3656);
xnor U3950 (N_3950,N_3565,N_3593);
nand U3951 (N_3951,N_3632,N_3644);
nor U3952 (N_3952,N_3731,N_3729);
nor U3953 (N_3953,N_3738,N_3604);
or U3954 (N_3954,N_3744,N_3618);
nor U3955 (N_3955,N_3584,N_3655);
nor U3956 (N_3956,N_3699,N_3712);
and U3957 (N_3957,N_3745,N_3683);
nor U3958 (N_3958,N_3516,N_3650);
or U3959 (N_3959,N_3502,N_3582);
or U3960 (N_3960,N_3622,N_3710);
nor U3961 (N_3961,N_3632,N_3600);
and U3962 (N_3962,N_3602,N_3688);
and U3963 (N_3963,N_3594,N_3647);
nand U3964 (N_3964,N_3594,N_3641);
xor U3965 (N_3965,N_3748,N_3528);
and U3966 (N_3966,N_3611,N_3650);
nand U3967 (N_3967,N_3607,N_3600);
xnor U3968 (N_3968,N_3523,N_3590);
nor U3969 (N_3969,N_3748,N_3518);
nor U3970 (N_3970,N_3749,N_3515);
xor U3971 (N_3971,N_3635,N_3512);
or U3972 (N_3972,N_3607,N_3620);
nor U3973 (N_3973,N_3570,N_3623);
or U3974 (N_3974,N_3655,N_3548);
or U3975 (N_3975,N_3728,N_3678);
nand U3976 (N_3976,N_3604,N_3567);
nand U3977 (N_3977,N_3683,N_3620);
nand U3978 (N_3978,N_3682,N_3741);
nor U3979 (N_3979,N_3612,N_3641);
or U3980 (N_3980,N_3728,N_3594);
nor U3981 (N_3981,N_3613,N_3654);
xor U3982 (N_3982,N_3702,N_3694);
xnor U3983 (N_3983,N_3563,N_3657);
nor U3984 (N_3984,N_3672,N_3642);
or U3985 (N_3985,N_3534,N_3738);
nand U3986 (N_3986,N_3660,N_3746);
nor U3987 (N_3987,N_3632,N_3597);
and U3988 (N_3988,N_3664,N_3592);
or U3989 (N_3989,N_3697,N_3575);
or U3990 (N_3990,N_3502,N_3536);
and U3991 (N_3991,N_3591,N_3564);
and U3992 (N_3992,N_3513,N_3522);
or U3993 (N_3993,N_3612,N_3608);
nor U3994 (N_3994,N_3572,N_3568);
nor U3995 (N_3995,N_3670,N_3569);
xnor U3996 (N_3996,N_3525,N_3736);
and U3997 (N_3997,N_3705,N_3570);
nand U3998 (N_3998,N_3740,N_3512);
xnor U3999 (N_3999,N_3727,N_3533);
nand U4000 (N_4000,N_3990,N_3941);
and U4001 (N_4001,N_3755,N_3782);
xor U4002 (N_4002,N_3917,N_3750);
xor U4003 (N_4003,N_3790,N_3769);
nand U4004 (N_4004,N_3845,N_3882);
and U4005 (N_4005,N_3835,N_3777);
xnor U4006 (N_4006,N_3817,N_3818);
nand U4007 (N_4007,N_3809,N_3810);
nand U4008 (N_4008,N_3972,N_3890);
nor U4009 (N_4009,N_3821,N_3836);
nor U4010 (N_4010,N_3898,N_3988);
xor U4011 (N_4011,N_3993,N_3914);
and U4012 (N_4012,N_3760,N_3780);
nand U4013 (N_4013,N_3753,N_3830);
xor U4014 (N_4014,N_3979,N_3932);
nand U4015 (N_4015,N_3975,N_3969);
and U4016 (N_4016,N_3935,N_3920);
and U4017 (N_4017,N_3874,N_3791);
or U4018 (N_4018,N_3759,N_3970);
nor U4019 (N_4019,N_3994,N_3913);
nand U4020 (N_4020,N_3858,N_3971);
or U4021 (N_4021,N_3880,N_3794);
xnor U4022 (N_4022,N_3894,N_3752);
nand U4023 (N_4023,N_3905,N_3856);
or U4024 (N_4024,N_3842,N_3866);
xnor U4025 (N_4025,N_3813,N_3958);
or U4026 (N_4026,N_3981,N_3837);
and U4027 (N_4027,N_3807,N_3977);
xnor U4028 (N_4028,N_3846,N_3860);
xnor U4029 (N_4029,N_3829,N_3862);
nor U4030 (N_4030,N_3937,N_3801);
or U4031 (N_4031,N_3853,N_3827);
nand U4032 (N_4032,N_3916,N_3924);
nor U4033 (N_4033,N_3840,N_3919);
nand U4034 (N_4034,N_3915,N_3761);
xnor U4035 (N_4035,N_3923,N_3831);
or U4036 (N_4036,N_3844,N_3768);
or U4037 (N_4037,N_3756,N_3870);
and U4038 (N_4038,N_3887,N_3978);
and U4039 (N_4039,N_3863,N_3798);
and U4040 (N_4040,N_3814,N_3852);
nand U4041 (N_4041,N_3825,N_3968);
nor U4042 (N_4042,N_3795,N_3967);
xnor U4043 (N_4043,N_3921,N_3767);
nor U4044 (N_4044,N_3765,N_3980);
xnor U4045 (N_4045,N_3816,N_3966);
and U4046 (N_4046,N_3877,N_3878);
or U4047 (N_4047,N_3951,N_3948);
xnor U4048 (N_4048,N_3773,N_3945);
and U4049 (N_4049,N_3823,N_3824);
nor U4050 (N_4050,N_3995,N_3869);
and U4051 (N_4051,N_3886,N_3800);
nand U4052 (N_4052,N_3875,N_3786);
and U4053 (N_4053,N_3751,N_3854);
and U4054 (N_4054,N_3868,N_3901);
or U4055 (N_4055,N_3865,N_3763);
nor U4056 (N_4056,N_3984,N_3892);
nor U4057 (N_4057,N_3778,N_3888);
nor U4058 (N_4058,N_3954,N_3986);
nand U4059 (N_4059,N_3762,N_3922);
nor U4060 (N_4060,N_3891,N_3861);
nand U4061 (N_4061,N_3959,N_3999);
nor U4062 (N_4062,N_3797,N_3904);
nor U4063 (N_4063,N_3847,N_3871);
nand U4064 (N_4064,N_3893,N_3873);
nor U4065 (N_4065,N_3787,N_3872);
xnor U4066 (N_4066,N_3938,N_3973);
xor U4067 (N_4067,N_3952,N_3855);
and U4068 (N_4068,N_3931,N_3802);
nand U4069 (N_4069,N_3895,N_3851);
xor U4070 (N_4070,N_3960,N_3947);
nand U4071 (N_4071,N_3838,N_3939);
nor U4072 (N_4072,N_3930,N_3883);
nand U4073 (N_4073,N_3857,N_3754);
xnor U4074 (N_4074,N_3841,N_3820);
nor U4075 (N_4075,N_3811,N_3849);
nand U4076 (N_4076,N_3771,N_3911);
nor U4077 (N_4077,N_3757,N_3889);
nor U4078 (N_4078,N_3964,N_3942);
or U4079 (N_4079,N_3758,N_3864);
or U4080 (N_4080,N_3806,N_3955);
xnor U4081 (N_4081,N_3792,N_3876);
or U4082 (N_4082,N_3772,N_3962);
and U4083 (N_4083,N_3929,N_3910);
nor U4084 (N_4084,N_3991,N_3940);
nand U4085 (N_4085,N_3900,N_3828);
nand U4086 (N_4086,N_3996,N_3925);
and U4087 (N_4087,N_3804,N_3957);
xnor U4088 (N_4088,N_3928,N_3982);
nand U4089 (N_4089,N_3805,N_3946);
or U4090 (N_4090,N_3956,N_3974);
and U4091 (N_4091,N_3985,N_3976);
nor U4092 (N_4092,N_3812,N_3788);
or U4093 (N_4093,N_3867,N_3764);
and U4094 (N_4094,N_3949,N_3781);
or U4095 (N_4095,N_3987,N_3850);
xor U4096 (N_4096,N_3897,N_3783);
and U4097 (N_4097,N_3785,N_3992);
nand U4098 (N_4098,N_3983,N_3950);
nand U4099 (N_4099,N_3848,N_3907);
nand U4100 (N_4100,N_3815,N_3903);
or U4101 (N_4101,N_3918,N_3953);
and U4102 (N_4102,N_3774,N_3927);
or U4103 (N_4103,N_3933,N_3944);
or U4104 (N_4104,N_3908,N_3896);
nor U4105 (N_4105,N_3997,N_3834);
nand U4106 (N_4106,N_3776,N_3799);
nor U4107 (N_4107,N_3989,N_3770);
nor U4108 (N_4108,N_3803,N_3902);
or U4109 (N_4109,N_3998,N_3859);
nand U4110 (N_4110,N_3839,N_3833);
and U4111 (N_4111,N_3808,N_3965);
xor U4112 (N_4112,N_3775,N_3832);
and U4113 (N_4113,N_3879,N_3884);
or U4114 (N_4114,N_3796,N_3934);
xor U4115 (N_4115,N_3843,N_3779);
xor U4116 (N_4116,N_3822,N_3906);
nor U4117 (N_4117,N_3926,N_3881);
or U4118 (N_4118,N_3909,N_3912);
and U4119 (N_4119,N_3943,N_3936);
xnor U4120 (N_4120,N_3784,N_3961);
or U4121 (N_4121,N_3963,N_3826);
nor U4122 (N_4122,N_3819,N_3766);
nor U4123 (N_4123,N_3793,N_3899);
or U4124 (N_4124,N_3885,N_3789);
and U4125 (N_4125,N_3903,N_3757);
nand U4126 (N_4126,N_3893,N_3808);
and U4127 (N_4127,N_3778,N_3921);
xor U4128 (N_4128,N_3950,N_3937);
and U4129 (N_4129,N_3792,N_3932);
and U4130 (N_4130,N_3873,N_3996);
xor U4131 (N_4131,N_3886,N_3789);
or U4132 (N_4132,N_3933,N_3753);
nor U4133 (N_4133,N_3880,N_3816);
or U4134 (N_4134,N_3955,N_3892);
or U4135 (N_4135,N_3967,N_3777);
nor U4136 (N_4136,N_3778,N_3874);
nor U4137 (N_4137,N_3981,N_3991);
nand U4138 (N_4138,N_3882,N_3978);
nor U4139 (N_4139,N_3906,N_3824);
xnor U4140 (N_4140,N_3873,N_3892);
xor U4141 (N_4141,N_3930,N_3893);
nand U4142 (N_4142,N_3840,N_3825);
nand U4143 (N_4143,N_3804,N_3768);
or U4144 (N_4144,N_3861,N_3850);
xor U4145 (N_4145,N_3930,N_3894);
xor U4146 (N_4146,N_3969,N_3806);
nor U4147 (N_4147,N_3981,N_3953);
or U4148 (N_4148,N_3992,N_3820);
xor U4149 (N_4149,N_3957,N_3861);
or U4150 (N_4150,N_3784,N_3894);
nor U4151 (N_4151,N_3788,N_3882);
nand U4152 (N_4152,N_3764,N_3904);
xnor U4153 (N_4153,N_3864,N_3881);
nand U4154 (N_4154,N_3930,N_3960);
nor U4155 (N_4155,N_3855,N_3884);
nor U4156 (N_4156,N_3783,N_3938);
nand U4157 (N_4157,N_3867,N_3998);
or U4158 (N_4158,N_3882,N_3796);
nor U4159 (N_4159,N_3966,N_3993);
xor U4160 (N_4160,N_3967,N_3771);
or U4161 (N_4161,N_3768,N_3772);
and U4162 (N_4162,N_3945,N_3785);
and U4163 (N_4163,N_3982,N_3944);
nand U4164 (N_4164,N_3880,N_3751);
xnor U4165 (N_4165,N_3759,N_3823);
nand U4166 (N_4166,N_3925,N_3884);
or U4167 (N_4167,N_3880,N_3915);
and U4168 (N_4168,N_3876,N_3959);
nor U4169 (N_4169,N_3765,N_3944);
nor U4170 (N_4170,N_3903,N_3912);
nor U4171 (N_4171,N_3866,N_3981);
and U4172 (N_4172,N_3774,N_3901);
or U4173 (N_4173,N_3767,N_3797);
and U4174 (N_4174,N_3841,N_3923);
xnor U4175 (N_4175,N_3977,N_3901);
or U4176 (N_4176,N_3840,N_3838);
or U4177 (N_4177,N_3928,N_3988);
or U4178 (N_4178,N_3769,N_3787);
and U4179 (N_4179,N_3772,N_3893);
xor U4180 (N_4180,N_3774,N_3805);
nand U4181 (N_4181,N_3776,N_3895);
xnor U4182 (N_4182,N_3977,N_3752);
or U4183 (N_4183,N_3898,N_3803);
and U4184 (N_4184,N_3897,N_3991);
nand U4185 (N_4185,N_3805,N_3881);
and U4186 (N_4186,N_3771,N_3921);
and U4187 (N_4187,N_3925,N_3972);
or U4188 (N_4188,N_3932,N_3884);
nand U4189 (N_4189,N_3954,N_3918);
and U4190 (N_4190,N_3894,N_3781);
xnor U4191 (N_4191,N_3872,N_3875);
nand U4192 (N_4192,N_3859,N_3794);
or U4193 (N_4193,N_3829,N_3920);
xnor U4194 (N_4194,N_3947,N_3887);
or U4195 (N_4195,N_3822,N_3966);
or U4196 (N_4196,N_3870,N_3809);
and U4197 (N_4197,N_3803,N_3926);
or U4198 (N_4198,N_3953,N_3926);
xor U4199 (N_4199,N_3935,N_3933);
or U4200 (N_4200,N_3916,N_3907);
or U4201 (N_4201,N_3799,N_3919);
nor U4202 (N_4202,N_3930,N_3785);
or U4203 (N_4203,N_3900,N_3824);
or U4204 (N_4204,N_3799,N_3831);
nor U4205 (N_4205,N_3849,N_3922);
nor U4206 (N_4206,N_3814,N_3963);
or U4207 (N_4207,N_3917,N_3784);
nor U4208 (N_4208,N_3912,N_3992);
and U4209 (N_4209,N_3962,N_3764);
or U4210 (N_4210,N_3752,N_3863);
nor U4211 (N_4211,N_3904,N_3906);
nand U4212 (N_4212,N_3891,N_3901);
nor U4213 (N_4213,N_3834,N_3863);
xor U4214 (N_4214,N_3785,N_3929);
xnor U4215 (N_4215,N_3989,N_3984);
and U4216 (N_4216,N_3894,N_3932);
xnor U4217 (N_4217,N_3927,N_3919);
and U4218 (N_4218,N_3900,N_3812);
or U4219 (N_4219,N_3940,N_3782);
and U4220 (N_4220,N_3757,N_3797);
xor U4221 (N_4221,N_3980,N_3942);
nor U4222 (N_4222,N_3862,N_3857);
or U4223 (N_4223,N_3919,N_3852);
or U4224 (N_4224,N_3833,N_3925);
nor U4225 (N_4225,N_3760,N_3840);
xor U4226 (N_4226,N_3860,N_3793);
xor U4227 (N_4227,N_3871,N_3868);
nand U4228 (N_4228,N_3970,N_3795);
xnor U4229 (N_4229,N_3923,N_3974);
nand U4230 (N_4230,N_3963,N_3953);
nand U4231 (N_4231,N_3800,N_3881);
xor U4232 (N_4232,N_3814,N_3949);
nor U4233 (N_4233,N_3888,N_3838);
and U4234 (N_4234,N_3980,N_3880);
xnor U4235 (N_4235,N_3871,N_3839);
nand U4236 (N_4236,N_3875,N_3967);
or U4237 (N_4237,N_3794,N_3951);
or U4238 (N_4238,N_3939,N_3859);
and U4239 (N_4239,N_3840,N_3866);
or U4240 (N_4240,N_3856,N_3978);
nand U4241 (N_4241,N_3776,N_3839);
or U4242 (N_4242,N_3823,N_3788);
nor U4243 (N_4243,N_3972,N_3812);
or U4244 (N_4244,N_3928,N_3977);
or U4245 (N_4245,N_3817,N_3936);
xor U4246 (N_4246,N_3914,N_3983);
nor U4247 (N_4247,N_3840,N_3953);
nor U4248 (N_4248,N_3983,N_3951);
or U4249 (N_4249,N_3770,N_3852);
nor U4250 (N_4250,N_4168,N_4199);
or U4251 (N_4251,N_4071,N_4183);
nor U4252 (N_4252,N_4160,N_4220);
nor U4253 (N_4253,N_4149,N_4127);
nand U4254 (N_4254,N_4205,N_4050);
xnor U4255 (N_4255,N_4120,N_4113);
nand U4256 (N_4256,N_4118,N_4147);
or U4257 (N_4257,N_4055,N_4212);
nor U4258 (N_4258,N_4176,N_4235);
and U4259 (N_4259,N_4049,N_4066);
and U4260 (N_4260,N_4027,N_4013);
or U4261 (N_4261,N_4022,N_4141);
and U4262 (N_4262,N_4069,N_4230);
or U4263 (N_4263,N_4023,N_4005);
and U4264 (N_4264,N_4241,N_4107);
xor U4265 (N_4265,N_4133,N_4000);
and U4266 (N_4266,N_4053,N_4126);
nand U4267 (N_4267,N_4248,N_4209);
xor U4268 (N_4268,N_4232,N_4096);
nor U4269 (N_4269,N_4078,N_4076);
xor U4270 (N_4270,N_4070,N_4009);
xnor U4271 (N_4271,N_4156,N_4181);
xor U4272 (N_4272,N_4024,N_4187);
nand U4273 (N_4273,N_4144,N_4136);
and U4274 (N_4274,N_4048,N_4082);
and U4275 (N_4275,N_4179,N_4128);
and U4276 (N_4276,N_4152,N_4017);
or U4277 (N_4277,N_4042,N_4065);
xor U4278 (N_4278,N_4134,N_4083);
nor U4279 (N_4279,N_4135,N_4240);
and U4280 (N_4280,N_4057,N_4154);
xnor U4281 (N_4281,N_4196,N_4067);
nand U4282 (N_4282,N_4226,N_4040);
xnor U4283 (N_4283,N_4056,N_4112);
and U4284 (N_4284,N_4225,N_4245);
and U4285 (N_4285,N_4170,N_4234);
xor U4286 (N_4286,N_4028,N_4215);
or U4287 (N_4287,N_4195,N_4249);
nor U4288 (N_4288,N_4124,N_4011);
xor U4289 (N_4289,N_4025,N_4063);
xor U4290 (N_4290,N_4004,N_4015);
and U4291 (N_4291,N_4123,N_4242);
or U4292 (N_4292,N_4158,N_4090);
xor U4293 (N_4293,N_4148,N_4210);
xor U4294 (N_4294,N_4142,N_4041);
nor U4295 (N_4295,N_4099,N_4091);
or U4296 (N_4296,N_4021,N_4044);
and U4297 (N_4297,N_4052,N_4084);
nor U4298 (N_4298,N_4102,N_4054);
nor U4299 (N_4299,N_4244,N_4008);
and U4300 (N_4300,N_4138,N_4109);
nand U4301 (N_4301,N_4060,N_4026);
or U4302 (N_4302,N_4197,N_4012);
nand U4303 (N_4303,N_4016,N_4033);
or U4304 (N_4304,N_4150,N_4191);
and U4305 (N_4305,N_4064,N_4051);
nor U4306 (N_4306,N_4146,N_4037);
nor U4307 (N_4307,N_4182,N_4121);
and U4308 (N_4308,N_4175,N_4098);
or U4309 (N_4309,N_4155,N_4130);
and U4310 (N_4310,N_4074,N_4122);
and U4311 (N_4311,N_4014,N_4189);
nor U4312 (N_4312,N_4247,N_4081);
nand U4313 (N_4313,N_4218,N_4031);
xor U4314 (N_4314,N_4072,N_4105);
or U4315 (N_4315,N_4001,N_4110);
or U4316 (N_4316,N_4172,N_4139);
or U4317 (N_4317,N_4068,N_4193);
and U4318 (N_4318,N_4007,N_4213);
nor U4319 (N_4319,N_4207,N_4204);
and U4320 (N_4320,N_4173,N_4020);
xor U4321 (N_4321,N_4058,N_4219);
or U4322 (N_4322,N_4104,N_4117);
or U4323 (N_4323,N_4243,N_4062);
nor U4324 (N_4324,N_4184,N_4237);
nand U4325 (N_4325,N_4200,N_4227);
xnor U4326 (N_4326,N_4002,N_4140);
xnor U4327 (N_4327,N_4029,N_4223);
or U4328 (N_4328,N_4178,N_4162);
nand U4329 (N_4329,N_4239,N_4194);
xor U4330 (N_4330,N_4228,N_4171);
nor U4331 (N_4331,N_4151,N_4224);
xnor U4332 (N_4332,N_4116,N_4131);
or U4333 (N_4333,N_4019,N_4103);
nand U4334 (N_4334,N_4093,N_4153);
and U4335 (N_4335,N_4087,N_4161);
xnor U4336 (N_4336,N_4108,N_4164);
and U4337 (N_4337,N_4114,N_4165);
and U4338 (N_4338,N_4129,N_4180);
and U4339 (N_4339,N_4079,N_4073);
xnor U4340 (N_4340,N_4174,N_4075);
or U4341 (N_4341,N_4167,N_4169);
xor U4342 (N_4342,N_4203,N_4003);
and U4343 (N_4343,N_4166,N_4080);
or U4344 (N_4344,N_4125,N_4163);
or U4345 (N_4345,N_4132,N_4097);
xor U4346 (N_4346,N_4192,N_4010);
nor U4347 (N_4347,N_4201,N_4119);
nor U4348 (N_4348,N_4143,N_4092);
nor U4349 (N_4349,N_4094,N_4035);
or U4350 (N_4350,N_4202,N_4032);
nor U4351 (N_4351,N_4036,N_4231);
and U4352 (N_4352,N_4186,N_4157);
or U4353 (N_4353,N_4177,N_4045);
nand U4354 (N_4354,N_4211,N_4030);
nor U4355 (N_4355,N_4216,N_4086);
and U4356 (N_4356,N_4190,N_4229);
nand U4357 (N_4357,N_4089,N_4214);
nor U4358 (N_4358,N_4034,N_4198);
and U4359 (N_4359,N_4208,N_4006);
and U4360 (N_4360,N_4236,N_4059);
or U4361 (N_4361,N_4188,N_4095);
nor U4362 (N_4362,N_4039,N_4085);
nand U4363 (N_4363,N_4043,N_4206);
nand U4364 (N_4364,N_4046,N_4088);
and U4365 (N_4365,N_4159,N_4238);
xor U4366 (N_4366,N_4077,N_4101);
nand U4367 (N_4367,N_4100,N_4145);
nand U4368 (N_4368,N_4047,N_4137);
or U4369 (N_4369,N_4222,N_4111);
xor U4370 (N_4370,N_4106,N_4038);
and U4371 (N_4371,N_4115,N_4217);
nand U4372 (N_4372,N_4018,N_4185);
xnor U4373 (N_4373,N_4221,N_4233);
and U4374 (N_4374,N_4246,N_4061);
nand U4375 (N_4375,N_4021,N_4004);
xnor U4376 (N_4376,N_4196,N_4123);
xnor U4377 (N_4377,N_4071,N_4080);
xor U4378 (N_4378,N_4216,N_4104);
or U4379 (N_4379,N_4075,N_4211);
or U4380 (N_4380,N_4051,N_4045);
nor U4381 (N_4381,N_4245,N_4215);
nor U4382 (N_4382,N_4127,N_4122);
xnor U4383 (N_4383,N_4100,N_4162);
and U4384 (N_4384,N_4009,N_4231);
xor U4385 (N_4385,N_4177,N_4092);
or U4386 (N_4386,N_4138,N_4065);
xnor U4387 (N_4387,N_4211,N_4069);
xnor U4388 (N_4388,N_4092,N_4116);
and U4389 (N_4389,N_4129,N_4242);
nor U4390 (N_4390,N_4233,N_4222);
and U4391 (N_4391,N_4057,N_4205);
or U4392 (N_4392,N_4039,N_4186);
nor U4393 (N_4393,N_4076,N_4214);
xnor U4394 (N_4394,N_4037,N_4132);
or U4395 (N_4395,N_4081,N_4070);
nor U4396 (N_4396,N_4158,N_4157);
and U4397 (N_4397,N_4078,N_4202);
or U4398 (N_4398,N_4076,N_4084);
nor U4399 (N_4399,N_4210,N_4089);
nand U4400 (N_4400,N_4247,N_4003);
xor U4401 (N_4401,N_4161,N_4241);
and U4402 (N_4402,N_4068,N_4186);
nand U4403 (N_4403,N_4143,N_4228);
or U4404 (N_4404,N_4039,N_4023);
or U4405 (N_4405,N_4075,N_4046);
xnor U4406 (N_4406,N_4157,N_4200);
and U4407 (N_4407,N_4154,N_4217);
nor U4408 (N_4408,N_4052,N_4160);
and U4409 (N_4409,N_4071,N_4124);
nor U4410 (N_4410,N_4187,N_4005);
nand U4411 (N_4411,N_4002,N_4116);
nor U4412 (N_4412,N_4101,N_4084);
and U4413 (N_4413,N_4053,N_4164);
nand U4414 (N_4414,N_4211,N_4088);
and U4415 (N_4415,N_4220,N_4148);
and U4416 (N_4416,N_4127,N_4001);
nor U4417 (N_4417,N_4158,N_4222);
and U4418 (N_4418,N_4062,N_4158);
xor U4419 (N_4419,N_4139,N_4081);
or U4420 (N_4420,N_4203,N_4205);
xor U4421 (N_4421,N_4074,N_4079);
nand U4422 (N_4422,N_4058,N_4080);
and U4423 (N_4423,N_4186,N_4154);
xnor U4424 (N_4424,N_4095,N_4109);
or U4425 (N_4425,N_4221,N_4075);
xor U4426 (N_4426,N_4051,N_4242);
nand U4427 (N_4427,N_4056,N_4097);
nand U4428 (N_4428,N_4134,N_4165);
nor U4429 (N_4429,N_4244,N_4087);
or U4430 (N_4430,N_4035,N_4089);
nand U4431 (N_4431,N_4033,N_4061);
nor U4432 (N_4432,N_4171,N_4195);
nor U4433 (N_4433,N_4180,N_4031);
nor U4434 (N_4434,N_4243,N_4198);
or U4435 (N_4435,N_4075,N_4067);
or U4436 (N_4436,N_4129,N_4184);
and U4437 (N_4437,N_4197,N_4133);
nand U4438 (N_4438,N_4169,N_4008);
nor U4439 (N_4439,N_4145,N_4229);
nor U4440 (N_4440,N_4003,N_4152);
nand U4441 (N_4441,N_4193,N_4082);
or U4442 (N_4442,N_4150,N_4116);
nor U4443 (N_4443,N_4151,N_4230);
xnor U4444 (N_4444,N_4019,N_4127);
xor U4445 (N_4445,N_4173,N_4167);
nand U4446 (N_4446,N_4100,N_4206);
and U4447 (N_4447,N_4076,N_4168);
xor U4448 (N_4448,N_4240,N_4044);
nand U4449 (N_4449,N_4069,N_4196);
xnor U4450 (N_4450,N_4198,N_4109);
xnor U4451 (N_4451,N_4112,N_4103);
and U4452 (N_4452,N_4204,N_4034);
nor U4453 (N_4453,N_4170,N_4161);
or U4454 (N_4454,N_4007,N_4003);
nand U4455 (N_4455,N_4063,N_4079);
and U4456 (N_4456,N_4081,N_4137);
nor U4457 (N_4457,N_4078,N_4148);
or U4458 (N_4458,N_4178,N_4017);
and U4459 (N_4459,N_4137,N_4009);
nor U4460 (N_4460,N_4236,N_4046);
and U4461 (N_4461,N_4013,N_4009);
xor U4462 (N_4462,N_4218,N_4220);
or U4463 (N_4463,N_4134,N_4125);
and U4464 (N_4464,N_4188,N_4109);
or U4465 (N_4465,N_4216,N_4094);
and U4466 (N_4466,N_4187,N_4101);
xor U4467 (N_4467,N_4218,N_4034);
and U4468 (N_4468,N_4195,N_4071);
nand U4469 (N_4469,N_4069,N_4146);
xor U4470 (N_4470,N_4169,N_4223);
nor U4471 (N_4471,N_4086,N_4038);
nand U4472 (N_4472,N_4203,N_4139);
nand U4473 (N_4473,N_4117,N_4047);
and U4474 (N_4474,N_4208,N_4097);
or U4475 (N_4475,N_4055,N_4087);
nor U4476 (N_4476,N_4200,N_4202);
or U4477 (N_4477,N_4092,N_4149);
and U4478 (N_4478,N_4220,N_4216);
and U4479 (N_4479,N_4021,N_4064);
xor U4480 (N_4480,N_4142,N_4013);
nor U4481 (N_4481,N_4040,N_4091);
or U4482 (N_4482,N_4079,N_4044);
or U4483 (N_4483,N_4062,N_4054);
nand U4484 (N_4484,N_4197,N_4207);
and U4485 (N_4485,N_4150,N_4141);
xnor U4486 (N_4486,N_4092,N_4118);
nand U4487 (N_4487,N_4121,N_4064);
nor U4488 (N_4488,N_4146,N_4111);
or U4489 (N_4489,N_4156,N_4073);
xor U4490 (N_4490,N_4233,N_4121);
or U4491 (N_4491,N_4071,N_4193);
or U4492 (N_4492,N_4107,N_4144);
nand U4493 (N_4493,N_4193,N_4059);
and U4494 (N_4494,N_4108,N_4033);
or U4495 (N_4495,N_4156,N_4057);
and U4496 (N_4496,N_4039,N_4107);
nand U4497 (N_4497,N_4248,N_4040);
nand U4498 (N_4498,N_4185,N_4017);
nor U4499 (N_4499,N_4069,N_4138);
or U4500 (N_4500,N_4295,N_4491);
nor U4501 (N_4501,N_4444,N_4268);
nor U4502 (N_4502,N_4496,N_4470);
nor U4503 (N_4503,N_4480,N_4395);
nand U4504 (N_4504,N_4429,N_4372);
xnor U4505 (N_4505,N_4456,N_4296);
or U4506 (N_4506,N_4399,N_4432);
or U4507 (N_4507,N_4400,N_4393);
nor U4508 (N_4508,N_4412,N_4466);
or U4509 (N_4509,N_4443,N_4338);
nor U4510 (N_4510,N_4390,N_4379);
or U4511 (N_4511,N_4333,N_4281);
xnor U4512 (N_4512,N_4357,N_4273);
nand U4513 (N_4513,N_4384,N_4417);
and U4514 (N_4514,N_4300,N_4326);
nor U4515 (N_4515,N_4292,N_4301);
or U4516 (N_4516,N_4499,N_4262);
or U4517 (N_4517,N_4469,N_4436);
xnor U4518 (N_4518,N_4284,N_4286);
nand U4519 (N_4519,N_4465,N_4360);
xnor U4520 (N_4520,N_4265,N_4314);
or U4521 (N_4521,N_4477,N_4373);
and U4522 (N_4522,N_4317,N_4342);
nor U4523 (N_4523,N_4433,N_4327);
and U4524 (N_4524,N_4340,N_4358);
nor U4525 (N_4525,N_4413,N_4462);
or U4526 (N_4526,N_4405,N_4370);
xnor U4527 (N_4527,N_4359,N_4403);
nand U4528 (N_4528,N_4282,N_4454);
or U4529 (N_4529,N_4485,N_4332);
nand U4530 (N_4530,N_4345,N_4419);
nor U4531 (N_4531,N_4442,N_4483);
nor U4532 (N_4532,N_4479,N_4427);
or U4533 (N_4533,N_4337,N_4418);
nand U4534 (N_4534,N_4294,N_4478);
or U4535 (N_4535,N_4458,N_4492);
nand U4536 (N_4536,N_4283,N_4375);
xnor U4537 (N_4537,N_4398,N_4253);
nor U4538 (N_4538,N_4488,N_4409);
nand U4539 (N_4539,N_4394,N_4331);
nand U4540 (N_4540,N_4315,N_4285);
and U4541 (N_4541,N_4451,N_4290);
nand U4542 (N_4542,N_4303,N_4252);
nand U4543 (N_4543,N_4309,N_4426);
and U4544 (N_4544,N_4264,N_4307);
and U4545 (N_4545,N_4457,N_4366);
nand U4546 (N_4546,N_4328,N_4420);
and U4547 (N_4547,N_4353,N_4453);
nand U4548 (N_4548,N_4494,N_4310);
nor U4549 (N_4549,N_4385,N_4367);
nand U4550 (N_4550,N_4259,N_4441);
and U4551 (N_4551,N_4493,N_4424);
or U4552 (N_4552,N_4377,N_4274);
and U4553 (N_4553,N_4455,N_4439);
and U4554 (N_4554,N_4411,N_4322);
nor U4555 (N_4555,N_4316,N_4334);
nand U4556 (N_4556,N_4490,N_4404);
nor U4557 (N_4557,N_4430,N_4425);
xnor U4558 (N_4558,N_4497,N_4368);
xor U4559 (N_4559,N_4335,N_4459);
xnor U4560 (N_4560,N_4389,N_4304);
or U4561 (N_4561,N_4448,N_4461);
and U4562 (N_4562,N_4329,N_4287);
or U4563 (N_4563,N_4380,N_4408);
and U4564 (N_4564,N_4346,N_4392);
or U4565 (N_4565,N_4431,N_4422);
and U4566 (N_4566,N_4498,N_4481);
xor U4567 (N_4567,N_4364,N_4361);
nor U4568 (N_4568,N_4387,N_4415);
xnor U4569 (N_4569,N_4365,N_4257);
and U4570 (N_4570,N_4449,N_4347);
or U4571 (N_4571,N_4330,N_4371);
and U4572 (N_4572,N_4348,N_4401);
nor U4573 (N_4573,N_4320,N_4382);
and U4574 (N_4574,N_4277,N_4402);
nor U4575 (N_4575,N_4339,N_4450);
xor U4576 (N_4576,N_4421,N_4298);
nor U4577 (N_4577,N_4258,N_4474);
xnor U4578 (N_4578,N_4473,N_4471);
nand U4579 (N_4579,N_4369,N_4278);
or U4580 (N_4580,N_4434,N_4476);
nor U4581 (N_4581,N_4468,N_4279);
and U4582 (N_4582,N_4318,N_4374);
nor U4583 (N_4583,N_4410,N_4349);
or U4584 (N_4584,N_4355,N_4437);
or U4585 (N_4585,N_4291,N_4251);
or U4586 (N_4586,N_4363,N_4495);
nand U4587 (N_4587,N_4452,N_4325);
or U4588 (N_4588,N_4313,N_4306);
or U4589 (N_4589,N_4486,N_4312);
and U4590 (N_4590,N_4299,N_4487);
or U4591 (N_4591,N_4383,N_4271);
and U4592 (N_4592,N_4447,N_4269);
xnor U4593 (N_4593,N_4446,N_4397);
nand U4594 (N_4594,N_4416,N_4352);
nand U4595 (N_4595,N_4438,N_4344);
nand U4596 (N_4596,N_4435,N_4256);
nor U4597 (N_4597,N_4263,N_4275);
nor U4598 (N_4598,N_4464,N_4311);
or U4599 (N_4599,N_4305,N_4319);
or U4600 (N_4600,N_4472,N_4280);
and U4601 (N_4601,N_4321,N_4423);
or U4602 (N_4602,N_4260,N_4276);
and U4603 (N_4603,N_4386,N_4302);
or U4604 (N_4604,N_4288,N_4354);
and U4605 (N_4605,N_4484,N_4343);
or U4606 (N_4606,N_4308,N_4270);
xnor U4607 (N_4607,N_4250,N_4350);
and U4608 (N_4608,N_4414,N_4463);
and U4609 (N_4609,N_4254,N_4356);
nand U4610 (N_4610,N_4407,N_4406);
nor U4611 (N_4611,N_4297,N_4396);
or U4612 (N_4612,N_4362,N_4289);
and U4613 (N_4613,N_4266,N_4378);
nor U4614 (N_4614,N_4351,N_4267);
and U4615 (N_4615,N_4261,N_4336);
nor U4616 (N_4616,N_4381,N_4391);
and U4617 (N_4617,N_4475,N_4376);
xor U4618 (N_4618,N_4489,N_4467);
or U4619 (N_4619,N_4460,N_4482);
nor U4620 (N_4620,N_4324,N_4323);
nand U4621 (N_4621,N_4388,N_4440);
nand U4622 (N_4622,N_4341,N_4428);
nor U4623 (N_4623,N_4445,N_4272);
or U4624 (N_4624,N_4255,N_4293);
or U4625 (N_4625,N_4289,N_4442);
xor U4626 (N_4626,N_4268,N_4462);
nand U4627 (N_4627,N_4459,N_4358);
nand U4628 (N_4628,N_4331,N_4442);
xor U4629 (N_4629,N_4475,N_4457);
and U4630 (N_4630,N_4271,N_4475);
nand U4631 (N_4631,N_4253,N_4455);
or U4632 (N_4632,N_4260,N_4478);
xor U4633 (N_4633,N_4258,N_4283);
xor U4634 (N_4634,N_4452,N_4390);
nor U4635 (N_4635,N_4496,N_4489);
nand U4636 (N_4636,N_4339,N_4372);
and U4637 (N_4637,N_4343,N_4271);
nor U4638 (N_4638,N_4398,N_4423);
nor U4639 (N_4639,N_4381,N_4332);
xor U4640 (N_4640,N_4337,N_4490);
xor U4641 (N_4641,N_4422,N_4260);
and U4642 (N_4642,N_4399,N_4272);
nor U4643 (N_4643,N_4433,N_4321);
nand U4644 (N_4644,N_4304,N_4453);
and U4645 (N_4645,N_4495,N_4329);
or U4646 (N_4646,N_4474,N_4385);
xnor U4647 (N_4647,N_4488,N_4492);
and U4648 (N_4648,N_4419,N_4361);
nand U4649 (N_4649,N_4274,N_4491);
nand U4650 (N_4650,N_4363,N_4367);
nand U4651 (N_4651,N_4251,N_4303);
and U4652 (N_4652,N_4423,N_4498);
or U4653 (N_4653,N_4283,N_4253);
nand U4654 (N_4654,N_4322,N_4496);
or U4655 (N_4655,N_4418,N_4328);
and U4656 (N_4656,N_4317,N_4302);
and U4657 (N_4657,N_4384,N_4458);
nand U4658 (N_4658,N_4422,N_4383);
nand U4659 (N_4659,N_4275,N_4293);
and U4660 (N_4660,N_4479,N_4463);
nand U4661 (N_4661,N_4423,N_4356);
and U4662 (N_4662,N_4319,N_4314);
nor U4663 (N_4663,N_4473,N_4375);
and U4664 (N_4664,N_4383,N_4333);
nor U4665 (N_4665,N_4405,N_4292);
nand U4666 (N_4666,N_4324,N_4294);
or U4667 (N_4667,N_4266,N_4403);
nor U4668 (N_4668,N_4419,N_4250);
nand U4669 (N_4669,N_4327,N_4456);
or U4670 (N_4670,N_4423,N_4357);
nor U4671 (N_4671,N_4409,N_4492);
nand U4672 (N_4672,N_4433,N_4310);
nand U4673 (N_4673,N_4344,N_4281);
or U4674 (N_4674,N_4342,N_4462);
nand U4675 (N_4675,N_4452,N_4324);
nand U4676 (N_4676,N_4443,N_4302);
and U4677 (N_4677,N_4479,N_4456);
nor U4678 (N_4678,N_4413,N_4304);
nand U4679 (N_4679,N_4372,N_4392);
nand U4680 (N_4680,N_4426,N_4308);
xor U4681 (N_4681,N_4313,N_4423);
nand U4682 (N_4682,N_4400,N_4488);
or U4683 (N_4683,N_4497,N_4323);
nor U4684 (N_4684,N_4470,N_4327);
and U4685 (N_4685,N_4313,N_4298);
nor U4686 (N_4686,N_4348,N_4459);
xor U4687 (N_4687,N_4304,N_4423);
xor U4688 (N_4688,N_4409,N_4420);
xor U4689 (N_4689,N_4456,N_4453);
and U4690 (N_4690,N_4255,N_4430);
nand U4691 (N_4691,N_4382,N_4453);
xnor U4692 (N_4692,N_4271,N_4319);
nor U4693 (N_4693,N_4391,N_4346);
xnor U4694 (N_4694,N_4313,N_4394);
or U4695 (N_4695,N_4317,N_4481);
nand U4696 (N_4696,N_4489,N_4402);
and U4697 (N_4697,N_4339,N_4430);
nor U4698 (N_4698,N_4400,N_4264);
or U4699 (N_4699,N_4270,N_4252);
nand U4700 (N_4700,N_4344,N_4280);
nand U4701 (N_4701,N_4329,N_4320);
xor U4702 (N_4702,N_4402,N_4463);
nor U4703 (N_4703,N_4260,N_4307);
or U4704 (N_4704,N_4406,N_4378);
nor U4705 (N_4705,N_4275,N_4364);
nand U4706 (N_4706,N_4473,N_4489);
and U4707 (N_4707,N_4378,N_4433);
nand U4708 (N_4708,N_4298,N_4397);
xnor U4709 (N_4709,N_4344,N_4277);
or U4710 (N_4710,N_4326,N_4446);
xor U4711 (N_4711,N_4408,N_4270);
nor U4712 (N_4712,N_4363,N_4303);
and U4713 (N_4713,N_4485,N_4441);
nand U4714 (N_4714,N_4444,N_4386);
or U4715 (N_4715,N_4479,N_4470);
nand U4716 (N_4716,N_4466,N_4321);
and U4717 (N_4717,N_4395,N_4406);
and U4718 (N_4718,N_4363,N_4355);
xnor U4719 (N_4719,N_4318,N_4322);
nor U4720 (N_4720,N_4267,N_4304);
nand U4721 (N_4721,N_4328,N_4443);
nand U4722 (N_4722,N_4273,N_4299);
and U4723 (N_4723,N_4430,N_4348);
nand U4724 (N_4724,N_4371,N_4436);
nor U4725 (N_4725,N_4413,N_4375);
nand U4726 (N_4726,N_4362,N_4250);
and U4727 (N_4727,N_4420,N_4405);
nor U4728 (N_4728,N_4329,N_4400);
or U4729 (N_4729,N_4359,N_4283);
and U4730 (N_4730,N_4477,N_4272);
xnor U4731 (N_4731,N_4446,N_4342);
nor U4732 (N_4732,N_4318,N_4440);
nand U4733 (N_4733,N_4401,N_4271);
nand U4734 (N_4734,N_4462,N_4335);
nand U4735 (N_4735,N_4341,N_4290);
xnor U4736 (N_4736,N_4294,N_4474);
and U4737 (N_4737,N_4388,N_4304);
nand U4738 (N_4738,N_4276,N_4395);
and U4739 (N_4739,N_4442,N_4459);
and U4740 (N_4740,N_4267,N_4498);
xnor U4741 (N_4741,N_4419,N_4433);
or U4742 (N_4742,N_4261,N_4389);
xor U4743 (N_4743,N_4386,N_4369);
nor U4744 (N_4744,N_4304,N_4457);
xnor U4745 (N_4745,N_4324,N_4314);
and U4746 (N_4746,N_4291,N_4297);
xnor U4747 (N_4747,N_4283,N_4328);
and U4748 (N_4748,N_4319,N_4391);
and U4749 (N_4749,N_4476,N_4266);
nor U4750 (N_4750,N_4603,N_4703);
nor U4751 (N_4751,N_4690,N_4674);
and U4752 (N_4752,N_4546,N_4553);
xnor U4753 (N_4753,N_4728,N_4695);
and U4754 (N_4754,N_4713,N_4622);
nand U4755 (N_4755,N_4542,N_4643);
nand U4756 (N_4756,N_4531,N_4733);
xnor U4757 (N_4757,N_4620,N_4694);
nor U4758 (N_4758,N_4502,N_4641);
nor U4759 (N_4759,N_4572,N_4618);
or U4760 (N_4760,N_4732,N_4574);
xnor U4761 (N_4761,N_4719,N_4688);
xor U4762 (N_4762,N_4636,N_4539);
and U4763 (N_4763,N_4563,N_4665);
and U4764 (N_4764,N_4693,N_4509);
nand U4765 (N_4765,N_4734,N_4692);
or U4766 (N_4766,N_4746,N_4651);
xor U4767 (N_4767,N_4710,N_4528);
nor U4768 (N_4768,N_4564,N_4549);
and U4769 (N_4769,N_4616,N_4601);
or U4770 (N_4770,N_4701,N_4555);
nand U4771 (N_4771,N_4657,N_4606);
xnor U4772 (N_4772,N_4738,N_4550);
and U4773 (N_4773,N_4681,N_4634);
nor U4774 (N_4774,N_4679,N_4672);
xnor U4775 (N_4775,N_4716,N_4554);
and U4776 (N_4776,N_4538,N_4698);
nand U4777 (N_4777,N_4658,N_4562);
nand U4778 (N_4778,N_4578,N_4610);
nand U4779 (N_4779,N_4630,N_4737);
or U4780 (N_4780,N_4519,N_4534);
nand U4781 (N_4781,N_4584,N_4678);
and U4782 (N_4782,N_4525,N_4743);
and U4783 (N_4783,N_4704,N_4541);
nor U4784 (N_4784,N_4640,N_4548);
nor U4785 (N_4785,N_4614,N_4506);
nor U4786 (N_4786,N_4712,N_4514);
nor U4787 (N_4787,N_4568,N_4510);
and U4788 (N_4788,N_4705,N_4575);
and U4789 (N_4789,N_4512,N_4567);
or U4790 (N_4790,N_4645,N_4729);
and U4791 (N_4791,N_4566,N_4544);
nand U4792 (N_4792,N_4588,N_4505);
nor U4793 (N_4793,N_4726,N_4589);
xnor U4794 (N_4794,N_4676,N_4646);
nor U4795 (N_4795,N_4604,N_4659);
and U4796 (N_4796,N_4523,N_4532);
nor U4797 (N_4797,N_4661,N_4748);
or U4798 (N_4798,N_4552,N_4526);
and U4799 (N_4799,N_4558,N_4656);
or U4800 (N_4800,N_4621,N_4536);
and U4801 (N_4801,N_4708,N_4613);
nand U4802 (N_4802,N_4721,N_4709);
nor U4803 (N_4803,N_4520,N_4740);
or U4804 (N_4804,N_4675,N_4594);
or U4805 (N_4805,N_4591,N_4670);
nor U4806 (N_4806,N_4625,N_4633);
or U4807 (N_4807,N_4668,N_4624);
or U4808 (N_4808,N_4663,N_4569);
or U4809 (N_4809,N_4653,N_4654);
nor U4810 (N_4810,N_4682,N_4596);
nor U4811 (N_4811,N_4718,N_4608);
xnor U4812 (N_4812,N_4581,N_4673);
xnor U4813 (N_4813,N_4714,N_4619);
or U4814 (N_4814,N_4623,N_4609);
nand U4815 (N_4815,N_4725,N_4745);
xnor U4816 (N_4816,N_4628,N_4667);
nand U4817 (N_4817,N_4583,N_4741);
and U4818 (N_4818,N_4611,N_4617);
xor U4819 (N_4819,N_4739,N_4530);
or U4820 (N_4820,N_4504,N_4664);
or U4821 (N_4821,N_4561,N_4626);
nand U4822 (N_4822,N_4730,N_4685);
xor U4823 (N_4823,N_4501,N_4707);
nor U4824 (N_4824,N_4691,N_4533);
nand U4825 (N_4825,N_4735,N_4631);
or U4826 (N_4826,N_4590,N_4602);
nor U4827 (N_4827,N_4724,N_4699);
xor U4828 (N_4828,N_4700,N_4749);
or U4829 (N_4829,N_4545,N_4577);
nor U4830 (N_4830,N_4731,N_4727);
or U4831 (N_4831,N_4650,N_4747);
nand U4832 (N_4832,N_4711,N_4521);
or U4833 (N_4833,N_4696,N_4706);
nor U4834 (N_4834,N_4652,N_4587);
or U4835 (N_4835,N_4689,N_4686);
or U4836 (N_4836,N_4511,N_4615);
and U4837 (N_4837,N_4744,N_4715);
nand U4838 (N_4838,N_4559,N_4669);
or U4839 (N_4839,N_4666,N_4522);
or U4840 (N_4840,N_4736,N_4671);
nand U4841 (N_4841,N_4638,N_4579);
nor U4842 (N_4842,N_4647,N_4649);
xnor U4843 (N_4843,N_4597,N_4723);
xnor U4844 (N_4844,N_4598,N_4607);
nand U4845 (N_4845,N_4605,N_4529);
nor U4846 (N_4846,N_4503,N_4500);
nand U4847 (N_4847,N_4600,N_4644);
xnor U4848 (N_4848,N_4516,N_4639);
nand U4849 (N_4849,N_4680,N_4629);
or U4850 (N_4850,N_4717,N_4655);
xnor U4851 (N_4851,N_4576,N_4632);
and U4852 (N_4852,N_4627,N_4551);
xor U4853 (N_4853,N_4684,N_4599);
or U4854 (N_4854,N_4593,N_4515);
xor U4855 (N_4855,N_4556,N_4585);
xnor U4856 (N_4856,N_4507,N_4677);
and U4857 (N_4857,N_4697,N_4720);
nand U4858 (N_4858,N_4508,N_4565);
nor U4859 (N_4859,N_4592,N_4537);
nor U4860 (N_4860,N_4518,N_4702);
nor U4861 (N_4861,N_4648,N_4535);
xnor U4862 (N_4862,N_4660,N_4524);
nor U4863 (N_4863,N_4571,N_4683);
or U4864 (N_4864,N_4513,N_4595);
nand U4865 (N_4865,N_4582,N_4560);
or U4866 (N_4866,N_4517,N_4742);
nand U4867 (N_4867,N_4635,N_4557);
or U4868 (N_4868,N_4637,N_4527);
nand U4869 (N_4869,N_4722,N_4642);
xor U4870 (N_4870,N_4543,N_4580);
and U4871 (N_4871,N_4540,N_4612);
or U4872 (N_4872,N_4570,N_4586);
xor U4873 (N_4873,N_4687,N_4573);
nand U4874 (N_4874,N_4547,N_4662);
nor U4875 (N_4875,N_4618,N_4684);
xnor U4876 (N_4876,N_4571,N_4687);
nor U4877 (N_4877,N_4559,N_4611);
nand U4878 (N_4878,N_4745,N_4694);
nand U4879 (N_4879,N_4515,N_4701);
nor U4880 (N_4880,N_4627,N_4521);
and U4881 (N_4881,N_4700,N_4585);
nand U4882 (N_4882,N_4560,N_4625);
nand U4883 (N_4883,N_4632,N_4687);
and U4884 (N_4884,N_4746,N_4698);
or U4885 (N_4885,N_4660,N_4507);
nand U4886 (N_4886,N_4516,N_4564);
and U4887 (N_4887,N_4740,N_4523);
nor U4888 (N_4888,N_4731,N_4526);
and U4889 (N_4889,N_4543,N_4522);
nand U4890 (N_4890,N_4636,N_4653);
nor U4891 (N_4891,N_4518,N_4515);
nor U4892 (N_4892,N_4545,N_4510);
nor U4893 (N_4893,N_4692,N_4594);
xnor U4894 (N_4894,N_4525,N_4523);
or U4895 (N_4895,N_4692,N_4588);
and U4896 (N_4896,N_4703,N_4588);
nor U4897 (N_4897,N_4509,N_4566);
and U4898 (N_4898,N_4632,N_4726);
and U4899 (N_4899,N_4570,N_4600);
nor U4900 (N_4900,N_4638,N_4680);
or U4901 (N_4901,N_4525,N_4713);
and U4902 (N_4902,N_4624,N_4636);
xor U4903 (N_4903,N_4501,N_4656);
nand U4904 (N_4904,N_4581,N_4515);
xor U4905 (N_4905,N_4546,N_4634);
nor U4906 (N_4906,N_4547,N_4659);
and U4907 (N_4907,N_4668,N_4609);
and U4908 (N_4908,N_4722,N_4713);
and U4909 (N_4909,N_4600,N_4568);
or U4910 (N_4910,N_4720,N_4721);
nor U4911 (N_4911,N_4617,N_4694);
nand U4912 (N_4912,N_4602,N_4566);
nand U4913 (N_4913,N_4641,N_4628);
nor U4914 (N_4914,N_4586,N_4672);
nand U4915 (N_4915,N_4742,N_4705);
nand U4916 (N_4916,N_4574,N_4682);
xor U4917 (N_4917,N_4595,N_4623);
nor U4918 (N_4918,N_4528,N_4545);
nor U4919 (N_4919,N_4646,N_4722);
or U4920 (N_4920,N_4561,N_4547);
nor U4921 (N_4921,N_4748,N_4703);
or U4922 (N_4922,N_4688,N_4747);
or U4923 (N_4923,N_4594,N_4569);
or U4924 (N_4924,N_4681,N_4607);
nor U4925 (N_4925,N_4674,N_4519);
or U4926 (N_4926,N_4717,N_4691);
or U4927 (N_4927,N_4563,N_4662);
nand U4928 (N_4928,N_4574,N_4570);
nand U4929 (N_4929,N_4691,N_4636);
xor U4930 (N_4930,N_4652,N_4546);
or U4931 (N_4931,N_4748,N_4576);
or U4932 (N_4932,N_4633,N_4699);
nor U4933 (N_4933,N_4606,N_4596);
nor U4934 (N_4934,N_4669,N_4501);
nor U4935 (N_4935,N_4661,N_4581);
nand U4936 (N_4936,N_4740,N_4627);
nor U4937 (N_4937,N_4563,N_4527);
or U4938 (N_4938,N_4703,N_4596);
or U4939 (N_4939,N_4596,N_4665);
nand U4940 (N_4940,N_4734,N_4502);
nand U4941 (N_4941,N_4698,N_4545);
and U4942 (N_4942,N_4660,N_4560);
xor U4943 (N_4943,N_4693,N_4679);
nor U4944 (N_4944,N_4567,N_4681);
or U4945 (N_4945,N_4546,N_4683);
xor U4946 (N_4946,N_4573,N_4506);
nand U4947 (N_4947,N_4663,N_4608);
nor U4948 (N_4948,N_4574,N_4698);
nand U4949 (N_4949,N_4680,N_4627);
and U4950 (N_4950,N_4713,N_4569);
xnor U4951 (N_4951,N_4572,N_4570);
and U4952 (N_4952,N_4666,N_4686);
xor U4953 (N_4953,N_4736,N_4597);
and U4954 (N_4954,N_4559,N_4518);
nand U4955 (N_4955,N_4699,N_4741);
xnor U4956 (N_4956,N_4512,N_4597);
or U4957 (N_4957,N_4509,N_4746);
and U4958 (N_4958,N_4621,N_4624);
nor U4959 (N_4959,N_4599,N_4534);
xnor U4960 (N_4960,N_4741,N_4619);
and U4961 (N_4961,N_4584,N_4587);
nor U4962 (N_4962,N_4698,N_4627);
xnor U4963 (N_4963,N_4716,N_4504);
xnor U4964 (N_4964,N_4569,N_4667);
nor U4965 (N_4965,N_4724,N_4621);
nand U4966 (N_4966,N_4701,N_4593);
nor U4967 (N_4967,N_4683,N_4558);
nor U4968 (N_4968,N_4630,N_4508);
or U4969 (N_4969,N_4648,N_4579);
xor U4970 (N_4970,N_4730,N_4640);
nand U4971 (N_4971,N_4636,N_4502);
and U4972 (N_4972,N_4704,N_4688);
nor U4973 (N_4973,N_4518,N_4543);
nor U4974 (N_4974,N_4733,N_4713);
nor U4975 (N_4975,N_4561,N_4514);
xor U4976 (N_4976,N_4658,N_4508);
nand U4977 (N_4977,N_4628,N_4736);
or U4978 (N_4978,N_4675,N_4726);
nand U4979 (N_4979,N_4611,N_4581);
xnor U4980 (N_4980,N_4744,N_4599);
xnor U4981 (N_4981,N_4667,N_4613);
and U4982 (N_4982,N_4614,N_4572);
xor U4983 (N_4983,N_4567,N_4613);
or U4984 (N_4984,N_4619,N_4649);
nand U4985 (N_4985,N_4527,N_4662);
or U4986 (N_4986,N_4609,N_4578);
nand U4987 (N_4987,N_4664,N_4604);
nor U4988 (N_4988,N_4749,N_4524);
xnor U4989 (N_4989,N_4581,N_4679);
nor U4990 (N_4990,N_4554,N_4746);
xnor U4991 (N_4991,N_4551,N_4523);
or U4992 (N_4992,N_4620,N_4642);
xnor U4993 (N_4993,N_4577,N_4536);
xnor U4994 (N_4994,N_4745,N_4743);
xor U4995 (N_4995,N_4632,N_4552);
nand U4996 (N_4996,N_4665,N_4606);
nand U4997 (N_4997,N_4646,N_4618);
nand U4998 (N_4998,N_4544,N_4585);
nor U4999 (N_4999,N_4641,N_4706);
and U5000 (N_5000,N_4810,N_4803);
xor U5001 (N_5001,N_4912,N_4991);
xor U5002 (N_5002,N_4949,N_4986);
nor U5003 (N_5003,N_4799,N_4885);
xnor U5004 (N_5004,N_4752,N_4941);
nand U5005 (N_5005,N_4998,N_4893);
xnor U5006 (N_5006,N_4953,N_4851);
or U5007 (N_5007,N_4963,N_4878);
nor U5008 (N_5008,N_4853,N_4890);
and U5009 (N_5009,N_4967,N_4789);
xor U5010 (N_5010,N_4757,N_4806);
nand U5011 (N_5011,N_4954,N_4892);
nand U5012 (N_5012,N_4999,N_4914);
nand U5013 (N_5013,N_4997,N_4867);
nor U5014 (N_5014,N_4881,N_4966);
xor U5015 (N_5015,N_4942,N_4809);
xnor U5016 (N_5016,N_4819,N_4968);
nor U5017 (N_5017,N_4877,N_4945);
or U5018 (N_5018,N_4759,N_4830);
nor U5019 (N_5019,N_4797,N_4965);
or U5020 (N_5020,N_4792,N_4925);
and U5021 (N_5021,N_4932,N_4811);
and U5022 (N_5022,N_4871,N_4842);
and U5023 (N_5023,N_4971,N_4838);
and U5024 (N_5024,N_4787,N_4921);
and U5025 (N_5025,N_4850,N_4899);
or U5026 (N_5026,N_4961,N_4758);
nor U5027 (N_5027,N_4984,N_4785);
and U5028 (N_5028,N_4959,N_4858);
xor U5029 (N_5029,N_4772,N_4798);
nand U5030 (N_5030,N_4768,N_4948);
and U5031 (N_5031,N_4995,N_4927);
xor U5032 (N_5032,N_4822,N_4989);
xor U5033 (N_5033,N_4766,N_4859);
nor U5034 (N_5034,N_4911,N_4919);
xnor U5035 (N_5035,N_4751,N_4831);
nor U5036 (N_5036,N_4760,N_4804);
nand U5037 (N_5037,N_4754,N_4990);
nor U5038 (N_5038,N_4753,N_4970);
or U5039 (N_5039,N_4764,N_4889);
nor U5040 (N_5040,N_4902,N_4796);
or U5041 (N_5041,N_4983,N_4863);
nand U5042 (N_5042,N_4905,N_4762);
and U5043 (N_5043,N_4770,N_4765);
or U5044 (N_5044,N_4940,N_4982);
and U5045 (N_5045,N_4891,N_4866);
nand U5046 (N_5046,N_4956,N_4993);
xnor U5047 (N_5047,N_4779,N_4898);
nor U5048 (N_5048,N_4778,N_4934);
nand U5049 (N_5049,N_4864,N_4782);
and U5050 (N_5050,N_4832,N_4775);
nand U5051 (N_5051,N_4923,N_4801);
and U5052 (N_5052,N_4848,N_4937);
xor U5053 (N_5053,N_4916,N_4788);
nand U5054 (N_5054,N_4821,N_4996);
nor U5055 (N_5055,N_4888,N_4973);
and U5056 (N_5056,N_4976,N_4913);
and U5057 (N_5057,N_4897,N_4774);
nor U5058 (N_5058,N_4975,N_4992);
or U5059 (N_5059,N_4988,N_4755);
or U5060 (N_5060,N_4761,N_4869);
nor U5061 (N_5061,N_4813,N_4929);
and U5062 (N_5062,N_4946,N_4872);
nand U5063 (N_5063,N_4987,N_4835);
xor U5064 (N_5064,N_4763,N_4794);
nor U5065 (N_5065,N_4880,N_4933);
or U5066 (N_5066,N_4960,N_4874);
nor U5067 (N_5067,N_4786,N_4854);
and U5068 (N_5068,N_4833,N_4756);
or U5069 (N_5069,N_4834,N_4868);
xnor U5070 (N_5070,N_4994,N_4847);
nand U5071 (N_5071,N_4839,N_4817);
nor U5072 (N_5072,N_4780,N_4777);
xnor U5073 (N_5073,N_4807,N_4951);
xor U5074 (N_5074,N_4865,N_4906);
nor U5075 (N_5075,N_4922,N_4828);
nor U5076 (N_5076,N_4950,N_4978);
nor U5077 (N_5077,N_4860,N_4886);
or U5078 (N_5078,N_4955,N_4882);
nor U5079 (N_5079,N_4800,N_4875);
and U5080 (N_5080,N_4856,N_4944);
nor U5081 (N_5081,N_4790,N_4861);
xnor U5082 (N_5082,N_4802,N_4845);
nor U5083 (N_5083,N_4805,N_4849);
nor U5084 (N_5084,N_4964,N_4939);
nor U5085 (N_5085,N_4781,N_4795);
and U5086 (N_5086,N_4776,N_4894);
and U5087 (N_5087,N_4972,N_4767);
nand U5088 (N_5088,N_4930,N_4926);
and U5089 (N_5089,N_4903,N_4783);
nor U5090 (N_5090,N_4901,N_4876);
or U5091 (N_5091,N_4829,N_4826);
nor U5092 (N_5092,N_4895,N_4814);
nand U5093 (N_5093,N_4924,N_4977);
and U5094 (N_5094,N_4900,N_4947);
nor U5095 (N_5095,N_4985,N_4840);
nand U5096 (N_5096,N_4896,N_4815);
or U5097 (N_5097,N_4862,N_4943);
or U5098 (N_5098,N_4816,N_4846);
nor U5099 (N_5099,N_4907,N_4818);
nor U5100 (N_5100,N_4857,N_4773);
nor U5101 (N_5101,N_4824,N_4909);
and U5102 (N_5102,N_4962,N_4928);
xor U5103 (N_5103,N_4836,N_4883);
xor U5104 (N_5104,N_4957,N_4980);
xnor U5105 (N_5105,N_4750,N_4974);
xnor U5106 (N_5106,N_4910,N_4969);
or U5107 (N_5107,N_4958,N_4884);
nand U5108 (N_5108,N_4908,N_4841);
or U5109 (N_5109,N_4825,N_4920);
and U5110 (N_5110,N_4917,N_4981);
and U5111 (N_5111,N_4918,N_4935);
nand U5112 (N_5112,N_4936,N_4837);
nor U5113 (N_5113,N_4931,N_4844);
nor U5114 (N_5114,N_4855,N_4979);
nand U5115 (N_5115,N_4771,N_4879);
and U5116 (N_5116,N_4784,N_4870);
nor U5117 (N_5117,N_4812,N_4915);
xnor U5118 (N_5118,N_4808,N_4791);
and U5119 (N_5119,N_4769,N_4823);
nand U5120 (N_5120,N_4904,N_4952);
xor U5121 (N_5121,N_4873,N_4843);
xor U5122 (N_5122,N_4793,N_4938);
nor U5123 (N_5123,N_4852,N_4827);
or U5124 (N_5124,N_4820,N_4887);
and U5125 (N_5125,N_4868,N_4995);
and U5126 (N_5126,N_4863,N_4931);
nand U5127 (N_5127,N_4831,N_4960);
and U5128 (N_5128,N_4894,N_4962);
or U5129 (N_5129,N_4865,N_4940);
xor U5130 (N_5130,N_4880,N_4918);
xor U5131 (N_5131,N_4975,N_4788);
and U5132 (N_5132,N_4802,N_4865);
and U5133 (N_5133,N_4950,N_4848);
and U5134 (N_5134,N_4901,N_4837);
or U5135 (N_5135,N_4816,N_4889);
nand U5136 (N_5136,N_4902,N_4820);
nor U5137 (N_5137,N_4851,N_4988);
xnor U5138 (N_5138,N_4917,N_4833);
nor U5139 (N_5139,N_4788,N_4844);
xnor U5140 (N_5140,N_4852,N_4824);
xnor U5141 (N_5141,N_4792,N_4918);
nor U5142 (N_5142,N_4990,N_4825);
nor U5143 (N_5143,N_4815,N_4792);
or U5144 (N_5144,N_4942,N_4943);
xor U5145 (N_5145,N_4883,N_4978);
or U5146 (N_5146,N_4876,N_4986);
nor U5147 (N_5147,N_4856,N_4867);
xor U5148 (N_5148,N_4924,N_4846);
nor U5149 (N_5149,N_4837,N_4942);
nor U5150 (N_5150,N_4843,N_4865);
xnor U5151 (N_5151,N_4795,N_4875);
xor U5152 (N_5152,N_4827,N_4782);
or U5153 (N_5153,N_4909,N_4914);
and U5154 (N_5154,N_4855,N_4859);
xor U5155 (N_5155,N_4870,N_4885);
nor U5156 (N_5156,N_4890,N_4847);
nand U5157 (N_5157,N_4829,N_4760);
nand U5158 (N_5158,N_4795,N_4761);
nand U5159 (N_5159,N_4953,N_4758);
xnor U5160 (N_5160,N_4950,N_4835);
nand U5161 (N_5161,N_4853,N_4792);
xor U5162 (N_5162,N_4803,N_4871);
or U5163 (N_5163,N_4798,N_4827);
and U5164 (N_5164,N_4759,N_4851);
nor U5165 (N_5165,N_4976,N_4930);
nand U5166 (N_5166,N_4981,N_4914);
and U5167 (N_5167,N_4838,N_4931);
and U5168 (N_5168,N_4909,N_4893);
nand U5169 (N_5169,N_4862,N_4917);
nor U5170 (N_5170,N_4786,N_4879);
xnor U5171 (N_5171,N_4981,N_4951);
or U5172 (N_5172,N_4949,N_4980);
xnor U5173 (N_5173,N_4931,N_4829);
and U5174 (N_5174,N_4890,N_4858);
xor U5175 (N_5175,N_4862,N_4763);
and U5176 (N_5176,N_4987,N_4781);
nand U5177 (N_5177,N_4869,N_4891);
xor U5178 (N_5178,N_4987,N_4919);
or U5179 (N_5179,N_4825,N_4950);
nor U5180 (N_5180,N_4999,N_4863);
nand U5181 (N_5181,N_4767,N_4992);
nand U5182 (N_5182,N_4852,N_4785);
nand U5183 (N_5183,N_4988,N_4872);
nor U5184 (N_5184,N_4825,N_4805);
nand U5185 (N_5185,N_4816,N_4989);
xnor U5186 (N_5186,N_4974,N_4924);
nor U5187 (N_5187,N_4903,N_4994);
and U5188 (N_5188,N_4877,N_4872);
and U5189 (N_5189,N_4776,N_4931);
nand U5190 (N_5190,N_4946,N_4932);
nand U5191 (N_5191,N_4955,N_4784);
or U5192 (N_5192,N_4884,N_4776);
nor U5193 (N_5193,N_4901,N_4886);
nor U5194 (N_5194,N_4898,N_4885);
or U5195 (N_5195,N_4944,N_4910);
nor U5196 (N_5196,N_4760,N_4777);
xor U5197 (N_5197,N_4978,N_4809);
and U5198 (N_5198,N_4816,N_4949);
or U5199 (N_5199,N_4896,N_4765);
xnor U5200 (N_5200,N_4952,N_4784);
xor U5201 (N_5201,N_4766,N_4967);
xnor U5202 (N_5202,N_4923,N_4947);
and U5203 (N_5203,N_4898,N_4858);
nor U5204 (N_5204,N_4951,N_4814);
or U5205 (N_5205,N_4986,N_4851);
nor U5206 (N_5206,N_4893,N_4864);
nor U5207 (N_5207,N_4896,N_4934);
and U5208 (N_5208,N_4891,N_4879);
and U5209 (N_5209,N_4859,N_4981);
nand U5210 (N_5210,N_4889,N_4830);
or U5211 (N_5211,N_4939,N_4893);
xnor U5212 (N_5212,N_4893,N_4943);
nand U5213 (N_5213,N_4942,N_4939);
or U5214 (N_5214,N_4779,N_4895);
and U5215 (N_5215,N_4950,N_4814);
and U5216 (N_5216,N_4914,N_4915);
nand U5217 (N_5217,N_4782,N_4973);
nand U5218 (N_5218,N_4947,N_4798);
nand U5219 (N_5219,N_4812,N_4897);
and U5220 (N_5220,N_4827,N_4972);
or U5221 (N_5221,N_4904,N_4801);
nor U5222 (N_5222,N_4881,N_4807);
xnor U5223 (N_5223,N_4848,N_4930);
and U5224 (N_5224,N_4924,N_4799);
or U5225 (N_5225,N_4870,N_4750);
and U5226 (N_5226,N_4946,N_4897);
nor U5227 (N_5227,N_4762,N_4878);
nand U5228 (N_5228,N_4856,N_4910);
and U5229 (N_5229,N_4888,N_4754);
nor U5230 (N_5230,N_4958,N_4963);
xnor U5231 (N_5231,N_4955,N_4976);
nand U5232 (N_5232,N_4822,N_4795);
and U5233 (N_5233,N_4791,N_4937);
nand U5234 (N_5234,N_4908,N_4986);
nor U5235 (N_5235,N_4999,N_4806);
nand U5236 (N_5236,N_4901,N_4894);
nor U5237 (N_5237,N_4974,N_4836);
xnor U5238 (N_5238,N_4793,N_4800);
and U5239 (N_5239,N_4906,N_4919);
nand U5240 (N_5240,N_4847,N_4996);
nand U5241 (N_5241,N_4786,N_4763);
or U5242 (N_5242,N_4847,N_4910);
nor U5243 (N_5243,N_4893,N_4908);
and U5244 (N_5244,N_4987,N_4933);
xnor U5245 (N_5245,N_4912,N_4795);
xor U5246 (N_5246,N_4916,N_4975);
xnor U5247 (N_5247,N_4849,N_4881);
or U5248 (N_5248,N_4791,N_4974);
or U5249 (N_5249,N_4953,N_4817);
nand U5250 (N_5250,N_5137,N_5227);
nand U5251 (N_5251,N_5090,N_5014);
or U5252 (N_5252,N_5145,N_5178);
nor U5253 (N_5253,N_5111,N_5007);
nor U5254 (N_5254,N_5146,N_5105);
and U5255 (N_5255,N_5051,N_5098);
xor U5256 (N_5256,N_5058,N_5107);
nand U5257 (N_5257,N_5008,N_5134);
nor U5258 (N_5258,N_5237,N_5205);
nand U5259 (N_5259,N_5156,N_5119);
nor U5260 (N_5260,N_5140,N_5034);
xnor U5261 (N_5261,N_5240,N_5194);
nand U5262 (N_5262,N_5077,N_5039);
xor U5263 (N_5263,N_5023,N_5061);
nand U5264 (N_5264,N_5201,N_5216);
nor U5265 (N_5265,N_5215,N_5168);
or U5266 (N_5266,N_5018,N_5091);
and U5267 (N_5267,N_5095,N_5085);
nand U5268 (N_5268,N_5028,N_5226);
nor U5269 (N_5269,N_5245,N_5167);
nor U5270 (N_5270,N_5116,N_5186);
or U5271 (N_5271,N_5157,N_5093);
or U5272 (N_5272,N_5069,N_5219);
or U5273 (N_5273,N_5197,N_5059);
and U5274 (N_5274,N_5015,N_5249);
and U5275 (N_5275,N_5055,N_5114);
and U5276 (N_5276,N_5068,N_5244);
xnor U5277 (N_5277,N_5043,N_5211);
and U5278 (N_5278,N_5092,N_5212);
nor U5279 (N_5279,N_5173,N_5135);
xor U5280 (N_5280,N_5049,N_5081);
nand U5281 (N_5281,N_5172,N_5158);
nor U5282 (N_5282,N_5248,N_5188);
xor U5283 (N_5283,N_5047,N_5064);
nor U5284 (N_5284,N_5118,N_5189);
and U5285 (N_5285,N_5208,N_5067);
xor U5286 (N_5286,N_5224,N_5196);
and U5287 (N_5287,N_5121,N_5094);
nand U5288 (N_5288,N_5027,N_5080);
nand U5289 (N_5289,N_5239,N_5152);
or U5290 (N_5290,N_5083,N_5013);
or U5291 (N_5291,N_5163,N_5171);
nor U5292 (N_5292,N_5183,N_5184);
nor U5293 (N_5293,N_5225,N_5231);
nor U5294 (N_5294,N_5048,N_5151);
and U5295 (N_5295,N_5228,N_5076);
xor U5296 (N_5296,N_5170,N_5053);
or U5297 (N_5297,N_5030,N_5072);
xnor U5298 (N_5298,N_5056,N_5180);
nand U5299 (N_5299,N_5133,N_5210);
nand U5300 (N_5300,N_5169,N_5035);
and U5301 (N_5301,N_5160,N_5032);
xnor U5302 (N_5302,N_5022,N_5036);
or U5303 (N_5303,N_5166,N_5187);
and U5304 (N_5304,N_5129,N_5001);
or U5305 (N_5305,N_5123,N_5154);
nor U5306 (N_5306,N_5042,N_5016);
and U5307 (N_5307,N_5220,N_5086);
xor U5308 (N_5308,N_5079,N_5041);
nand U5309 (N_5309,N_5117,N_5174);
xor U5310 (N_5310,N_5143,N_5024);
xnor U5311 (N_5311,N_5177,N_5192);
xnor U5312 (N_5312,N_5142,N_5110);
nor U5313 (N_5313,N_5153,N_5103);
xor U5314 (N_5314,N_5207,N_5221);
nor U5315 (N_5315,N_5078,N_5162);
xor U5316 (N_5316,N_5235,N_5230);
xnor U5317 (N_5317,N_5089,N_5234);
xor U5318 (N_5318,N_5029,N_5124);
and U5319 (N_5319,N_5054,N_5071);
xor U5320 (N_5320,N_5199,N_5075);
nor U5321 (N_5321,N_5006,N_5179);
or U5322 (N_5322,N_5099,N_5217);
or U5323 (N_5323,N_5149,N_5181);
and U5324 (N_5324,N_5082,N_5011);
or U5325 (N_5325,N_5144,N_5052);
or U5326 (N_5326,N_5109,N_5131);
and U5327 (N_5327,N_5070,N_5044);
or U5328 (N_5328,N_5159,N_5038);
nand U5329 (N_5329,N_5242,N_5010);
and U5330 (N_5330,N_5074,N_5204);
or U5331 (N_5331,N_5198,N_5040);
xor U5332 (N_5332,N_5191,N_5246);
xnor U5333 (N_5333,N_5012,N_5087);
nor U5334 (N_5334,N_5065,N_5136);
nand U5335 (N_5335,N_5003,N_5057);
xnor U5336 (N_5336,N_5097,N_5031);
nor U5337 (N_5337,N_5127,N_5164);
nand U5338 (N_5338,N_5165,N_5120);
nor U5339 (N_5339,N_5132,N_5126);
and U5340 (N_5340,N_5002,N_5102);
nand U5341 (N_5341,N_5026,N_5190);
and U5342 (N_5342,N_5020,N_5236);
nor U5343 (N_5343,N_5004,N_5241);
and U5344 (N_5344,N_5009,N_5209);
nand U5345 (N_5345,N_5161,N_5213);
xnor U5346 (N_5346,N_5000,N_5243);
or U5347 (N_5347,N_5222,N_5150);
nand U5348 (N_5348,N_5193,N_5017);
xnor U5349 (N_5349,N_5148,N_5050);
xnor U5350 (N_5350,N_5084,N_5019);
xor U5351 (N_5351,N_5088,N_5125);
nor U5352 (N_5352,N_5233,N_5176);
or U5353 (N_5353,N_5223,N_5138);
or U5354 (N_5354,N_5115,N_5113);
or U5355 (N_5355,N_5066,N_5112);
xnor U5356 (N_5356,N_5200,N_5100);
or U5357 (N_5357,N_5122,N_5232);
and U5358 (N_5358,N_5060,N_5037);
and U5359 (N_5359,N_5182,N_5247);
nand U5360 (N_5360,N_5021,N_5195);
and U5361 (N_5361,N_5175,N_5101);
nand U5362 (N_5362,N_5108,N_5139);
nand U5363 (N_5363,N_5045,N_5206);
or U5364 (N_5364,N_5025,N_5155);
nor U5365 (N_5365,N_5130,N_5096);
nor U5366 (N_5366,N_5033,N_5147);
nor U5367 (N_5367,N_5073,N_5106);
nor U5368 (N_5368,N_5141,N_5046);
and U5369 (N_5369,N_5005,N_5238);
nand U5370 (N_5370,N_5062,N_5104);
and U5371 (N_5371,N_5218,N_5202);
nor U5372 (N_5372,N_5229,N_5128);
and U5373 (N_5373,N_5185,N_5203);
xor U5374 (N_5374,N_5214,N_5063);
nor U5375 (N_5375,N_5059,N_5116);
nand U5376 (N_5376,N_5155,N_5231);
xnor U5377 (N_5377,N_5018,N_5176);
nor U5378 (N_5378,N_5106,N_5239);
and U5379 (N_5379,N_5082,N_5009);
and U5380 (N_5380,N_5227,N_5161);
nand U5381 (N_5381,N_5033,N_5091);
or U5382 (N_5382,N_5209,N_5102);
or U5383 (N_5383,N_5226,N_5022);
nand U5384 (N_5384,N_5193,N_5091);
nand U5385 (N_5385,N_5043,N_5121);
xnor U5386 (N_5386,N_5147,N_5171);
and U5387 (N_5387,N_5019,N_5248);
xnor U5388 (N_5388,N_5045,N_5010);
nor U5389 (N_5389,N_5074,N_5249);
xor U5390 (N_5390,N_5193,N_5014);
xnor U5391 (N_5391,N_5193,N_5043);
xnor U5392 (N_5392,N_5145,N_5137);
nand U5393 (N_5393,N_5041,N_5145);
xnor U5394 (N_5394,N_5012,N_5223);
nand U5395 (N_5395,N_5136,N_5033);
or U5396 (N_5396,N_5020,N_5003);
nor U5397 (N_5397,N_5039,N_5194);
or U5398 (N_5398,N_5076,N_5018);
and U5399 (N_5399,N_5026,N_5052);
or U5400 (N_5400,N_5102,N_5242);
or U5401 (N_5401,N_5074,N_5156);
and U5402 (N_5402,N_5074,N_5199);
nand U5403 (N_5403,N_5061,N_5239);
xnor U5404 (N_5404,N_5242,N_5019);
nor U5405 (N_5405,N_5001,N_5088);
nand U5406 (N_5406,N_5199,N_5191);
xnor U5407 (N_5407,N_5175,N_5204);
xnor U5408 (N_5408,N_5094,N_5222);
or U5409 (N_5409,N_5147,N_5208);
or U5410 (N_5410,N_5088,N_5233);
nand U5411 (N_5411,N_5202,N_5174);
xor U5412 (N_5412,N_5018,N_5055);
or U5413 (N_5413,N_5211,N_5047);
and U5414 (N_5414,N_5214,N_5172);
and U5415 (N_5415,N_5165,N_5241);
and U5416 (N_5416,N_5164,N_5191);
or U5417 (N_5417,N_5198,N_5023);
xor U5418 (N_5418,N_5157,N_5218);
nor U5419 (N_5419,N_5249,N_5181);
nor U5420 (N_5420,N_5241,N_5208);
nor U5421 (N_5421,N_5104,N_5029);
and U5422 (N_5422,N_5154,N_5096);
or U5423 (N_5423,N_5191,N_5236);
nor U5424 (N_5424,N_5237,N_5147);
or U5425 (N_5425,N_5166,N_5189);
and U5426 (N_5426,N_5114,N_5185);
and U5427 (N_5427,N_5054,N_5072);
and U5428 (N_5428,N_5046,N_5055);
nor U5429 (N_5429,N_5213,N_5170);
and U5430 (N_5430,N_5093,N_5115);
or U5431 (N_5431,N_5248,N_5247);
or U5432 (N_5432,N_5082,N_5068);
or U5433 (N_5433,N_5034,N_5144);
xor U5434 (N_5434,N_5141,N_5138);
nand U5435 (N_5435,N_5165,N_5217);
xor U5436 (N_5436,N_5231,N_5235);
nand U5437 (N_5437,N_5142,N_5239);
nand U5438 (N_5438,N_5184,N_5022);
nor U5439 (N_5439,N_5008,N_5208);
nand U5440 (N_5440,N_5176,N_5210);
and U5441 (N_5441,N_5015,N_5184);
xnor U5442 (N_5442,N_5212,N_5022);
nand U5443 (N_5443,N_5241,N_5230);
nor U5444 (N_5444,N_5103,N_5205);
nor U5445 (N_5445,N_5226,N_5149);
xor U5446 (N_5446,N_5208,N_5075);
nor U5447 (N_5447,N_5083,N_5116);
xnor U5448 (N_5448,N_5219,N_5092);
nand U5449 (N_5449,N_5174,N_5126);
and U5450 (N_5450,N_5091,N_5224);
and U5451 (N_5451,N_5146,N_5207);
xnor U5452 (N_5452,N_5154,N_5204);
nand U5453 (N_5453,N_5084,N_5000);
nor U5454 (N_5454,N_5126,N_5153);
and U5455 (N_5455,N_5067,N_5197);
or U5456 (N_5456,N_5097,N_5092);
or U5457 (N_5457,N_5045,N_5221);
nor U5458 (N_5458,N_5053,N_5018);
nor U5459 (N_5459,N_5234,N_5041);
nand U5460 (N_5460,N_5110,N_5124);
nor U5461 (N_5461,N_5058,N_5234);
or U5462 (N_5462,N_5156,N_5054);
nor U5463 (N_5463,N_5237,N_5167);
nor U5464 (N_5464,N_5096,N_5080);
nor U5465 (N_5465,N_5228,N_5200);
and U5466 (N_5466,N_5222,N_5247);
and U5467 (N_5467,N_5191,N_5046);
xnor U5468 (N_5468,N_5225,N_5228);
xor U5469 (N_5469,N_5150,N_5001);
nor U5470 (N_5470,N_5054,N_5207);
nand U5471 (N_5471,N_5186,N_5233);
xor U5472 (N_5472,N_5164,N_5113);
nor U5473 (N_5473,N_5203,N_5167);
nor U5474 (N_5474,N_5209,N_5224);
nand U5475 (N_5475,N_5029,N_5122);
xnor U5476 (N_5476,N_5143,N_5003);
nand U5477 (N_5477,N_5032,N_5064);
nand U5478 (N_5478,N_5198,N_5190);
and U5479 (N_5479,N_5079,N_5068);
nand U5480 (N_5480,N_5153,N_5059);
or U5481 (N_5481,N_5098,N_5167);
nor U5482 (N_5482,N_5156,N_5053);
or U5483 (N_5483,N_5082,N_5003);
nor U5484 (N_5484,N_5202,N_5091);
and U5485 (N_5485,N_5234,N_5161);
and U5486 (N_5486,N_5049,N_5224);
xnor U5487 (N_5487,N_5096,N_5206);
nor U5488 (N_5488,N_5009,N_5191);
and U5489 (N_5489,N_5208,N_5090);
nor U5490 (N_5490,N_5190,N_5034);
xnor U5491 (N_5491,N_5079,N_5179);
and U5492 (N_5492,N_5233,N_5164);
xor U5493 (N_5493,N_5160,N_5210);
xor U5494 (N_5494,N_5228,N_5207);
and U5495 (N_5495,N_5021,N_5027);
nand U5496 (N_5496,N_5194,N_5007);
and U5497 (N_5497,N_5085,N_5079);
and U5498 (N_5498,N_5126,N_5245);
nor U5499 (N_5499,N_5020,N_5141);
and U5500 (N_5500,N_5367,N_5437);
nand U5501 (N_5501,N_5431,N_5327);
xor U5502 (N_5502,N_5386,N_5392);
nand U5503 (N_5503,N_5472,N_5433);
or U5504 (N_5504,N_5255,N_5494);
or U5505 (N_5505,N_5400,N_5273);
and U5506 (N_5506,N_5389,N_5432);
or U5507 (N_5507,N_5287,N_5463);
nand U5508 (N_5508,N_5436,N_5484);
xnor U5509 (N_5509,N_5440,N_5364);
and U5510 (N_5510,N_5260,N_5333);
xor U5511 (N_5511,N_5474,N_5279);
nor U5512 (N_5512,N_5483,N_5261);
nand U5513 (N_5513,N_5376,N_5290);
nor U5514 (N_5514,N_5286,N_5485);
or U5515 (N_5515,N_5357,N_5384);
nor U5516 (N_5516,N_5407,N_5331);
and U5517 (N_5517,N_5382,N_5465);
xnor U5518 (N_5518,N_5319,N_5322);
nor U5519 (N_5519,N_5309,N_5481);
nand U5520 (N_5520,N_5269,N_5341);
xor U5521 (N_5521,N_5305,N_5476);
nor U5522 (N_5522,N_5359,N_5324);
xor U5523 (N_5523,N_5443,N_5438);
nand U5524 (N_5524,N_5492,N_5416);
and U5525 (N_5525,N_5499,N_5434);
nand U5526 (N_5526,N_5394,N_5366);
nand U5527 (N_5527,N_5401,N_5352);
nor U5528 (N_5528,N_5450,N_5423);
and U5529 (N_5529,N_5312,N_5455);
nor U5530 (N_5530,N_5398,N_5390);
and U5531 (N_5531,N_5425,N_5314);
xor U5532 (N_5532,N_5428,N_5466);
nand U5533 (N_5533,N_5262,N_5265);
and U5534 (N_5534,N_5289,N_5393);
xor U5535 (N_5535,N_5297,N_5325);
nor U5536 (N_5536,N_5372,N_5422);
or U5537 (N_5537,N_5361,N_5329);
and U5538 (N_5538,N_5449,N_5301);
or U5539 (N_5539,N_5315,N_5412);
nand U5540 (N_5540,N_5275,N_5468);
and U5541 (N_5541,N_5293,N_5282);
xnor U5542 (N_5542,N_5411,N_5452);
nand U5543 (N_5543,N_5439,N_5459);
and U5544 (N_5544,N_5444,N_5285);
or U5545 (N_5545,N_5469,N_5473);
xnor U5546 (N_5546,N_5300,N_5413);
or U5547 (N_5547,N_5471,N_5259);
and U5548 (N_5548,N_5424,N_5368);
or U5549 (N_5549,N_5462,N_5385);
or U5550 (N_5550,N_5334,N_5266);
nand U5551 (N_5551,N_5447,N_5295);
and U5552 (N_5552,N_5490,N_5268);
and U5553 (N_5553,N_5464,N_5267);
and U5554 (N_5554,N_5427,N_5362);
and U5555 (N_5555,N_5256,N_5426);
and U5556 (N_5556,N_5283,N_5391);
or U5557 (N_5557,N_5350,N_5363);
or U5558 (N_5558,N_5461,N_5253);
nand U5559 (N_5559,N_5467,N_5373);
and U5560 (N_5560,N_5403,N_5277);
nand U5561 (N_5561,N_5264,N_5291);
or U5562 (N_5562,N_5370,N_5257);
and U5563 (N_5563,N_5272,N_5351);
xnor U5564 (N_5564,N_5396,N_5345);
nor U5565 (N_5565,N_5489,N_5454);
nand U5566 (N_5566,N_5408,N_5251);
and U5567 (N_5567,N_5343,N_5446);
xor U5568 (N_5568,N_5418,N_5288);
nor U5569 (N_5569,N_5380,N_5337);
xnor U5570 (N_5570,N_5338,N_5441);
and U5571 (N_5571,N_5284,N_5296);
or U5572 (N_5572,N_5419,N_5460);
nor U5573 (N_5573,N_5307,N_5375);
nor U5574 (N_5574,N_5310,N_5303);
xnor U5575 (N_5575,N_5326,N_5317);
and U5576 (N_5576,N_5371,N_5347);
nor U5577 (N_5577,N_5448,N_5365);
nand U5578 (N_5578,N_5276,N_5360);
nor U5579 (N_5579,N_5404,N_5453);
xor U5580 (N_5580,N_5335,N_5344);
xnor U5581 (N_5581,N_5294,N_5496);
nand U5582 (N_5582,N_5387,N_5498);
nand U5583 (N_5583,N_5281,N_5379);
xor U5584 (N_5584,N_5479,N_5429);
and U5585 (N_5585,N_5487,N_5313);
nand U5586 (N_5586,N_5417,N_5480);
and U5587 (N_5587,N_5470,N_5377);
and U5588 (N_5588,N_5406,N_5442);
nor U5589 (N_5589,N_5250,N_5478);
nand U5590 (N_5590,N_5270,N_5302);
and U5591 (N_5591,N_5356,N_5409);
and U5592 (N_5592,N_5488,N_5321);
and U5593 (N_5593,N_5482,N_5491);
or U5594 (N_5594,N_5320,N_5497);
and U5595 (N_5595,N_5292,N_5304);
nor U5596 (N_5596,N_5323,N_5405);
or U5597 (N_5597,N_5381,N_5388);
or U5598 (N_5598,N_5349,N_5311);
or U5599 (N_5599,N_5456,N_5475);
nand U5600 (N_5600,N_5355,N_5397);
xnor U5601 (N_5601,N_5358,N_5410);
xor U5602 (N_5602,N_5420,N_5340);
and U5603 (N_5603,N_5252,N_5414);
and U5604 (N_5604,N_5328,N_5332);
nor U5605 (N_5605,N_5348,N_5308);
or U5606 (N_5606,N_5495,N_5458);
nor U5607 (N_5607,N_5278,N_5399);
and U5608 (N_5608,N_5477,N_5451);
or U5609 (N_5609,N_5378,N_5336);
nor U5610 (N_5610,N_5306,N_5445);
nor U5611 (N_5611,N_5339,N_5493);
nand U5612 (N_5612,N_5421,N_5457);
nor U5613 (N_5613,N_5353,N_5402);
nand U5614 (N_5614,N_5486,N_5258);
nand U5615 (N_5615,N_5342,N_5430);
or U5616 (N_5616,N_5280,N_5383);
and U5617 (N_5617,N_5254,N_5299);
xor U5618 (N_5618,N_5263,N_5369);
nand U5619 (N_5619,N_5346,N_5316);
xnor U5620 (N_5620,N_5330,N_5271);
and U5621 (N_5621,N_5435,N_5374);
and U5622 (N_5622,N_5354,N_5395);
and U5623 (N_5623,N_5274,N_5415);
nand U5624 (N_5624,N_5298,N_5318);
xor U5625 (N_5625,N_5417,N_5406);
nand U5626 (N_5626,N_5264,N_5412);
nor U5627 (N_5627,N_5477,N_5273);
xnor U5628 (N_5628,N_5285,N_5434);
or U5629 (N_5629,N_5430,N_5373);
or U5630 (N_5630,N_5349,N_5401);
nor U5631 (N_5631,N_5255,N_5357);
xnor U5632 (N_5632,N_5460,N_5295);
nand U5633 (N_5633,N_5295,N_5475);
or U5634 (N_5634,N_5397,N_5499);
nand U5635 (N_5635,N_5401,N_5420);
or U5636 (N_5636,N_5457,N_5365);
nand U5637 (N_5637,N_5375,N_5412);
or U5638 (N_5638,N_5475,N_5498);
xor U5639 (N_5639,N_5329,N_5255);
or U5640 (N_5640,N_5387,N_5354);
nand U5641 (N_5641,N_5329,N_5424);
xnor U5642 (N_5642,N_5498,N_5453);
or U5643 (N_5643,N_5281,N_5265);
and U5644 (N_5644,N_5498,N_5269);
nand U5645 (N_5645,N_5414,N_5347);
nand U5646 (N_5646,N_5308,N_5354);
xnor U5647 (N_5647,N_5264,N_5369);
and U5648 (N_5648,N_5370,N_5340);
xor U5649 (N_5649,N_5292,N_5324);
nand U5650 (N_5650,N_5293,N_5278);
or U5651 (N_5651,N_5407,N_5433);
and U5652 (N_5652,N_5271,N_5496);
and U5653 (N_5653,N_5442,N_5346);
xnor U5654 (N_5654,N_5364,N_5456);
xor U5655 (N_5655,N_5391,N_5302);
nand U5656 (N_5656,N_5296,N_5472);
xor U5657 (N_5657,N_5459,N_5334);
or U5658 (N_5658,N_5250,N_5337);
and U5659 (N_5659,N_5378,N_5315);
xor U5660 (N_5660,N_5460,N_5337);
xnor U5661 (N_5661,N_5335,N_5261);
nand U5662 (N_5662,N_5266,N_5264);
xor U5663 (N_5663,N_5491,N_5347);
and U5664 (N_5664,N_5398,N_5465);
xnor U5665 (N_5665,N_5398,N_5328);
and U5666 (N_5666,N_5258,N_5277);
xnor U5667 (N_5667,N_5437,N_5481);
nor U5668 (N_5668,N_5313,N_5254);
nand U5669 (N_5669,N_5365,N_5285);
nor U5670 (N_5670,N_5284,N_5405);
nand U5671 (N_5671,N_5318,N_5371);
nor U5672 (N_5672,N_5344,N_5461);
or U5673 (N_5673,N_5445,N_5352);
xor U5674 (N_5674,N_5498,N_5429);
xor U5675 (N_5675,N_5444,N_5473);
nor U5676 (N_5676,N_5312,N_5494);
or U5677 (N_5677,N_5403,N_5460);
xor U5678 (N_5678,N_5481,N_5293);
and U5679 (N_5679,N_5459,N_5348);
and U5680 (N_5680,N_5350,N_5464);
xor U5681 (N_5681,N_5442,N_5417);
nand U5682 (N_5682,N_5369,N_5279);
xnor U5683 (N_5683,N_5462,N_5472);
nor U5684 (N_5684,N_5471,N_5491);
nand U5685 (N_5685,N_5445,N_5386);
and U5686 (N_5686,N_5376,N_5273);
and U5687 (N_5687,N_5393,N_5318);
and U5688 (N_5688,N_5463,N_5425);
or U5689 (N_5689,N_5287,N_5339);
nor U5690 (N_5690,N_5344,N_5339);
and U5691 (N_5691,N_5292,N_5405);
and U5692 (N_5692,N_5336,N_5298);
xnor U5693 (N_5693,N_5374,N_5490);
nor U5694 (N_5694,N_5425,N_5365);
nand U5695 (N_5695,N_5428,N_5440);
or U5696 (N_5696,N_5282,N_5419);
xor U5697 (N_5697,N_5451,N_5434);
nor U5698 (N_5698,N_5400,N_5360);
nand U5699 (N_5699,N_5266,N_5391);
xor U5700 (N_5700,N_5439,N_5454);
nand U5701 (N_5701,N_5255,N_5424);
nor U5702 (N_5702,N_5287,N_5369);
and U5703 (N_5703,N_5421,N_5343);
or U5704 (N_5704,N_5298,N_5296);
xor U5705 (N_5705,N_5398,N_5479);
nand U5706 (N_5706,N_5441,N_5452);
nand U5707 (N_5707,N_5267,N_5447);
nand U5708 (N_5708,N_5338,N_5481);
and U5709 (N_5709,N_5302,N_5465);
and U5710 (N_5710,N_5454,N_5318);
nand U5711 (N_5711,N_5413,N_5285);
or U5712 (N_5712,N_5462,N_5288);
nor U5713 (N_5713,N_5284,N_5332);
and U5714 (N_5714,N_5338,N_5344);
or U5715 (N_5715,N_5283,N_5409);
and U5716 (N_5716,N_5404,N_5492);
xor U5717 (N_5717,N_5346,N_5272);
or U5718 (N_5718,N_5281,N_5302);
and U5719 (N_5719,N_5260,N_5474);
or U5720 (N_5720,N_5273,N_5371);
or U5721 (N_5721,N_5413,N_5416);
nor U5722 (N_5722,N_5313,N_5466);
xor U5723 (N_5723,N_5484,N_5341);
and U5724 (N_5724,N_5460,N_5331);
nor U5725 (N_5725,N_5468,N_5456);
and U5726 (N_5726,N_5428,N_5472);
and U5727 (N_5727,N_5346,N_5414);
or U5728 (N_5728,N_5277,N_5450);
or U5729 (N_5729,N_5274,N_5300);
or U5730 (N_5730,N_5387,N_5425);
or U5731 (N_5731,N_5497,N_5493);
and U5732 (N_5732,N_5330,N_5489);
xnor U5733 (N_5733,N_5410,N_5267);
nand U5734 (N_5734,N_5472,N_5385);
or U5735 (N_5735,N_5335,N_5255);
nand U5736 (N_5736,N_5465,N_5437);
nor U5737 (N_5737,N_5400,N_5282);
or U5738 (N_5738,N_5305,N_5265);
nor U5739 (N_5739,N_5382,N_5473);
and U5740 (N_5740,N_5343,N_5443);
and U5741 (N_5741,N_5330,N_5255);
nand U5742 (N_5742,N_5440,N_5266);
nand U5743 (N_5743,N_5309,N_5290);
nor U5744 (N_5744,N_5341,N_5271);
nor U5745 (N_5745,N_5462,N_5281);
and U5746 (N_5746,N_5275,N_5459);
xnor U5747 (N_5747,N_5482,N_5330);
and U5748 (N_5748,N_5492,N_5427);
or U5749 (N_5749,N_5437,N_5487);
nor U5750 (N_5750,N_5738,N_5519);
or U5751 (N_5751,N_5695,N_5588);
nand U5752 (N_5752,N_5554,N_5606);
nor U5753 (N_5753,N_5691,N_5569);
or U5754 (N_5754,N_5715,N_5581);
nor U5755 (N_5755,N_5642,N_5627);
or U5756 (N_5756,N_5673,N_5589);
or U5757 (N_5757,N_5726,N_5528);
or U5758 (N_5758,N_5643,N_5530);
nand U5759 (N_5759,N_5578,N_5582);
or U5760 (N_5760,N_5712,N_5565);
or U5761 (N_5761,N_5711,N_5682);
and U5762 (N_5762,N_5584,N_5508);
or U5763 (N_5763,N_5634,N_5677);
xor U5764 (N_5764,N_5723,N_5628);
nor U5765 (N_5765,N_5720,N_5592);
xor U5766 (N_5766,N_5529,N_5690);
nand U5767 (N_5767,N_5646,N_5551);
and U5768 (N_5768,N_5559,N_5647);
or U5769 (N_5769,N_5524,N_5610);
xor U5770 (N_5770,N_5639,N_5618);
xor U5771 (N_5771,N_5629,N_5697);
and U5772 (N_5772,N_5544,N_5686);
and U5773 (N_5773,N_5567,N_5600);
or U5774 (N_5774,N_5687,N_5611);
or U5775 (N_5775,N_5648,N_5607);
nor U5776 (N_5776,N_5709,N_5616);
xor U5777 (N_5777,N_5652,N_5573);
nor U5778 (N_5778,N_5729,N_5692);
or U5779 (N_5779,N_5568,N_5742);
and U5780 (N_5780,N_5710,N_5527);
nand U5781 (N_5781,N_5502,N_5603);
nor U5782 (N_5782,N_5670,N_5577);
xor U5783 (N_5783,N_5556,N_5659);
nand U5784 (N_5784,N_5698,N_5651);
xor U5785 (N_5785,N_5717,N_5641);
nor U5786 (N_5786,N_5552,N_5721);
nor U5787 (N_5787,N_5625,N_5674);
nand U5788 (N_5788,N_5623,N_5526);
nand U5789 (N_5789,N_5617,N_5521);
xnor U5790 (N_5790,N_5566,N_5596);
nor U5791 (N_5791,N_5671,N_5683);
and U5792 (N_5792,N_5580,N_5702);
xnor U5793 (N_5793,N_5681,N_5658);
nor U5794 (N_5794,N_5550,N_5736);
nor U5795 (N_5795,N_5672,N_5700);
and U5796 (N_5796,N_5733,N_5540);
nand U5797 (N_5797,N_5707,N_5590);
xnor U5798 (N_5798,N_5587,N_5688);
xnor U5799 (N_5799,N_5562,N_5727);
nor U5800 (N_5800,N_5663,N_5680);
nor U5801 (N_5801,N_5539,N_5598);
nand U5802 (N_5802,N_5509,N_5503);
or U5803 (N_5803,N_5576,N_5746);
or U5804 (N_5804,N_5655,N_5553);
xnor U5805 (N_5805,N_5696,N_5511);
or U5806 (N_5806,N_5693,N_5701);
and U5807 (N_5807,N_5579,N_5522);
xor U5808 (N_5808,N_5520,N_5694);
or U5809 (N_5809,N_5593,N_5548);
xor U5810 (N_5810,N_5708,N_5513);
nor U5811 (N_5811,N_5608,N_5679);
nand U5812 (N_5812,N_5512,N_5541);
nand U5813 (N_5813,N_5704,N_5633);
nor U5814 (N_5814,N_5745,N_5668);
nor U5815 (N_5815,N_5725,N_5716);
and U5816 (N_5816,N_5730,N_5703);
or U5817 (N_5817,N_5735,N_5574);
nand U5818 (N_5818,N_5615,N_5661);
nand U5819 (N_5819,N_5741,N_5514);
nor U5820 (N_5820,N_5583,N_5505);
and U5821 (N_5821,N_5619,N_5501);
nor U5822 (N_5822,N_5523,N_5635);
xnor U5823 (N_5823,N_5605,N_5506);
nand U5824 (N_5824,N_5561,N_5743);
and U5825 (N_5825,N_5620,N_5713);
or U5826 (N_5826,N_5599,N_5557);
xnor U5827 (N_5827,N_5739,N_5591);
nand U5828 (N_5828,N_5585,N_5549);
nor U5829 (N_5829,N_5586,N_5676);
and U5830 (N_5830,N_5689,N_5664);
nand U5831 (N_5831,N_5678,N_5645);
nor U5832 (N_5832,N_5604,N_5669);
nand U5833 (N_5833,N_5719,N_5560);
xnor U5834 (N_5834,N_5660,N_5546);
and U5835 (N_5835,N_5657,N_5699);
or U5836 (N_5836,N_5644,N_5609);
or U5837 (N_5837,N_5517,N_5500);
nand U5838 (N_5838,N_5525,N_5649);
and U5839 (N_5839,N_5737,N_5722);
nand U5840 (N_5840,N_5515,N_5631);
and U5841 (N_5841,N_5705,N_5747);
and U5842 (N_5842,N_5595,N_5516);
nand U5843 (N_5843,N_5653,N_5572);
and U5844 (N_5844,N_5638,N_5732);
or U5845 (N_5845,N_5636,N_5613);
nor U5846 (N_5846,N_5534,N_5675);
and U5847 (N_5847,N_5667,N_5594);
xnor U5848 (N_5848,N_5734,N_5563);
or U5849 (N_5849,N_5601,N_5622);
xnor U5850 (N_5850,N_5612,N_5538);
nor U5851 (N_5851,N_5685,N_5518);
nand U5852 (N_5852,N_5662,N_5731);
nand U5853 (N_5853,N_5531,N_5632);
and U5854 (N_5854,N_5537,N_5724);
xor U5855 (N_5855,N_5543,N_5656);
xor U5856 (N_5856,N_5666,N_5571);
xnor U5857 (N_5857,N_5507,N_5740);
and U5858 (N_5858,N_5558,N_5535);
nand U5859 (N_5859,N_5718,N_5510);
xor U5860 (N_5860,N_5564,N_5728);
nor U5861 (N_5861,N_5654,N_5614);
or U5862 (N_5862,N_5504,N_5624);
and U5863 (N_5863,N_5684,N_5536);
nor U5864 (N_5864,N_5665,N_5748);
or U5865 (N_5865,N_5547,N_5621);
nor U5866 (N_5866,N_5555,N_5545);
nor U5867 (N_5867,N_5533,N_5602);
nand U5868 (N_5868,N_5714,N_5706);
nor U5869 (N_5869,N_5650,N_5570);
and U5870 (N_5870,N_5637,N_5630);
nor U5871 (N_5871,N_5749,N_5626);
or U5872 (N_5872,N_5597,N_5575);
and U5873 (N_5873,N_5640,N_5744);
xnor U5874 (N_5874,N_5532,N_5542);
or U5875 (N_5875,N_5522,N_5625);
nor U5876 (N_5876,N_5735,N_5621);
or U5877 (N_5877,N_5645,N_5672);
nand U5878 (N_5878,N_5688,N_5731);
or U5879 (N_5879,N_5622,N_5547);
nor U5880 (N_5880,N_5719,N_5746);
nand U5881 (N_5881,N_5554,N_5747);
or U5882 (N_5882,N_5642,N_5543);
nand U5883 (N_5883,N_5618,N_5517);
xor U5884 (N_5884,N_5692,N_5560);
or U5885 (N_5885,N_5731,N_5666);
nand U5886 (N_5886,N_5693,N_5508);
xor U5887 (N_5887,N_5578,N_5677);
nand U5888 (N_5888,N_5524,N_5746);
or U5889 (N_5889,N_5690,N_5646);
nand U5890 (N_5890,N_5665,N_5667);
and U5891 (N_5891,N_5627,N_5653);
or U5892 (N_5892,N_5729,N_5633);
xnor U5893 (N_5893,N_5646,N_5653);
and U5894 (N_5894,N_5697,N_5701);
or U5895 (N_5895,N_5621,N_5633);
or U5896 (N_5896,N_5568,N_5736);
nand U5897 (N_5897,N_5567,N_5627);
xnor U5898 (N_5898,N_5604,N_5696);
or U5899 (N_5899,N_5745,N_5689);
xnor U5900 (N_5900,N_5612,N_5676);
xor U5901 (N_5901,N_5506,N_5501);
or U5902 (N_5902,N_5558,N_5692);
xor U5903 (N_5903,N_5538,N_5524);
xor U5904 (N_5904,N_5709,N_5578);
nor U5905 (N_5905,N_5658,N_5675);
nor U5906 (N_5906,N_5625,N_5501);
xnor U5907 (N_5907,N_5723,N_5504);
nand U5908 (N_5908,N_5603,N_5665);
nor U5909 (N_5909,N_5674,N_5671);
and U5910 (N_5910,N_5665,N_5672);
xor U5911 (N_5911,N_5633,N_5705);
xor U5912 (N_5912,N_5547,N_5594);
and U5913 (N_5913,N_5583,N_5711);
nand U5914 (N_5914,N_5510,N_5658);
and U5915 (N_5915,N_5587,N_5502);
or U5916 (N_5916,N_5682,N_5523);
nor U5917 (N_5917,N_5681,N_5620);
nand U5918 (N_5918,N_5633,N_5569);
nor U5919 (N_5919,N_5627,N_5704);
nand U5920 (N_5920,N_5634,N_5507);
nand U5921 (N_5921,N_5512,N_5653);
nand U5922 (N_5922,N_5542,N_5572);
nand U5923 (N_5923,N_5733,N_5720);
xor U5924 (N_5924,N_5699,N_5614);
and U5925 (N_5925,N_5613,N_5594);
xor U5926 (N_5926,N_5555,N_5546);
or U5927 (N_5927,N_5650,N_5577);
and U5928 (N_5928,N_5645,N_5694);
and U5929 (N_5929,N_5679,N_5536);
or U5930 (N_5930,N_5574,N_5532);
nor U5931 (N_5931,N_5598,N_5649);
xnor U5932 (N_5932,N_5572,N_5538);
xor U5933 (N_5933,N_5552,N_5644);
nand U5934 (N_5934,N_5638,N_5658);
nor U5935 (N_5935,N_5504,N_5575);
or U5936 (N_5936,N_5602,N_5574);
and U5937 (N_5937,N_5740,N_5584);
xor U5938 (N_5938,N_5630,N_5726);
nand U5939 (N_5939,N_5522,N_5583);
xor U5940 (N_5940,N_5535,N_5719);
or U5941 (N_5941,N_5690,N_5689);
xnor U5942 (N_5942,N_5551,N_5686);
or U5943 (N_5943,N_5681,N_5639);
nor U5944 (N_5944,N_5680,N_5563);
and U5945 (N_5945,N_5634,N_5558);
xnor U5946 (N_5946,N_5549,N_5559);
nor U5947 (N_5947,N_5511,N_5626);
xnor U5948 (N_5948,N_5617,N_5545);
xor U5949 (N_5949,N_5527,N_5600);
nor U5950 (N_5950,N_5747,N_5697);
xor U5951 (N_5951,N_5561,N_5585);
and U5952 (N_5952,N_5592,N_5648);
or U5953 (N_5953,N_5576,N_5683);
or U5954 (N_5954,N_5727,N_5552);
or U5955 (N_5955,N_5695,N_5619);
and U5956 (N_5956,N_5540,N_5545);
nor U5957 (N_5957,N_5698,N_5700);
and U5958 (N_5958,N_5739,N_5611);
nand U5959 (N_5959,N_5626,N_5510);
nand U5960 (N_5960,N_5699,N_5645);
and U5961 (N_5961,N_5700,N_5656);
xor U5962 (N_5962,N_5667,N_5692);
and U5963 (N_5963,N_5526,N_5628);
xor U5964 (N_5964,N_5549,N_5675);
or U5965 (N_5965,N_5743,N_5660);
nand U5966 (N_5966,N_5538,N_5723);
xnor U5967 (N_5967,N_5501,N_5640);
nand U5968 (N_5968,N_5525,N_5573);
nor U5969 (N_5969,N_5607,N_5746);
nand U5970 (N_5970,N_5735,N_5639);
or U5971 (N_5971,N_5729,N_5565);
xor U5972 (N_5972,N_5519,N_5698);
or U5973 (N_5973,N_5573,N_5513);
xor U5974 (N_5974,N_5653,N_5579);
nor U5975 (N_5975,N_5605,N_5576);
or U5976 (N_5976,N_5685,N_5596);
xor U5977 (N_5977,N_5536,N_5711);
nor U5978 (N_5978,N_5500,N_5583);
xnor U5979 (N_5979,N_5508,N_5522);
nor U5980 (N_5980,N_5654,N_5554);
and U5981 (N_5981,N_5604,N_5727);
and U5982 (N_5982,N_5586,N_5652);
or U5983 (N_5983,N_5719,N_5591);
or U5984 (N_5984,N_5724,N_5627);
xnor U5985 (N_5985,N_5547,N_5522);
nor U5986 (N_5986,N_5727,N_5633);
nand U5987 (N_5987,N_5574,N_5648);
and U5988 (N_5988,N_5519,N_5684);
and U5989 (N_5989,N_5647,N_5517);
and U5990 (N_5990,N_5630,N_5683);
nand U5991 (N_5991,N_5543,N_5665);
xnor U5992 (N_5992,N_5651,N_5636);
nor U5993 (N_5993,N_5558,N_5530);
nand U5994 (N_5994,N_5716,N_5607);
nand U5995 (N_5995,N_5606,N_5539);
or U5996 (N_5996,N_5704,N_5588);
and U5997 (N_5997,N_5550,N_5746);
or U5998 (N_5998,N_5696,N_5503);
nor U5999 (N_5999,N_5725,N_5623);
and U6000 (N_6000,N_5801,N_5997);
or U6001 (N_6001,N_5768,N_5931);
or U6002 (N_6002,N_5813,N_5962);
nor U6003 (N_6003,N_5818,N_5804);
nand U6004 (N_6004,N_5845,N_5900);
nand U6005 (N_6005,N_5917,N_5950);
nand U6006 (N_6006,N_5980,N_5988);
and U6007 (N_6007,N_5874,N_5972);
and U6008 (N_6008,N_5883,N_5762);
nand U6009 (N_6009,N_5771,N_5852);
nor U6010 (N_6010,N_5807,N_5864);
nand U6011 (N_6011,N_5919,N_5822);
nand U6012 (N_6012,N_5786,N_5834);
nand U6013 (N_6013,N_5871,N_5985);
nor U6014 (N_6014,N_5947,N_5821);
nor U6015 (N_6015,N_5894,N_5909);
and U6016 (N_6016,N_5964,N_5974);
nand U6017 (N_6017,N_5904,N_5925);
xnor U6018 (N_6018,N_5986,N_5893);
nand U6019 (N_6019,N_5884,N_5803);
nor U6020 (N_6020,N_5857,N_5926);
and U6021 (N_6021,N_5844,N_5906);
nor U6022 (N_6022,N_5887,N_5969);
nand U6023 (N_6023,N_5814,N_5794);
nand U6024 (N_6024,N_5903,N_5775);
nand U6025 (N_6025,N_5832,N_5809);
nor U6026 (N_6026,N_5790,N_5802);
xnor U6027 (N_6027,N_5949,N_5895);
nand U6028 (N_6028,N_5930,N_5867);
nor U6029 (N_6029,N_5922,N_5860);
and U6030 (N_6030,N_5849,N_5779);
and U6031 (N_6031,N_5861,N_5838);
xnor U6032 (N_6032,N_5777,N_5853);
and U6033 (N_6033,N_5940,N_5916);
xnor U6034 (N_6034,N_5851,N_5820);
or U6035 (N_6035,N_5817,N_5939);
nor U6036 (N_6036,N_5907,N_5810);
nand U6037 (N_6037,N_5758,N_5911);
or U6038 (N_6038,N_5889,N_5761);
nor U6039 (N_6039,N_5798,N_5928);
xnor U6040 (N_6040,N_5766,N_5971);
or U6041 (N_6041,N_5836,N_5800);
nand U6042 (N_6042,N_5875,N_5825);
xnor U6043 (N_6043,N_5858,N_5862);
nand U6044 (N_6044,N_5990,N_5989);
xnor U6045 (N_6045,N_5885,N_5993);
xnor U6046 (N_6046,N_5886,N_5929);
and U6047 (N_6047,N_5856,N_5827);
xnor U6048 (N_6048,N_5952,N_5995);
nor U6049 (N_6049,N_5973,N_5991);
nor U6050 (N_6050,N_5773,N_5927);
nor U6051 (N_6051,N_5908,N_5815);
xnor U6052 (N_6052,N_5846,N_5979);
and U6053 (N_6053,N_5776,N_5982);
nor U6054 (N_6054,N_5759,N_5921);
nand U6055 (N_6055,N_5924,N_5863);
or U6056 (N_6056,N_5787,N_5797);
nand U6057 (N_6057,N_5869,N_5914);
or U6058 (N_6058,N_5769,N_5840);
nor U6059 (N_6059,N_5806,N_5850);
or U6060 (N_6060,N_5937,N_5896);
and U6061 (N_6061,N_5942,N_5953);
and U6062 (N_6062,N_5932,N_5913);
and U6063 (N_6063,N_5783,N_5791);
xnor U6064 (N_6064,N_5841,N_5782);
xor U6065 (N_6065,N_5890,N_5915);
or U6066 (N_6066,N_5912,N_5774);
nor U6067 (N_6067,N_5918,N_5981);
or U6068 (N_6068,N_5765,N_5984);
nand U6069 (N_6069,N_5785,N_5975);
or U6070 (N_6070,N_5870,N_5837);
or U6071 (N_6071,N_5760,N_5999);
and U6072 (N_6072,N_5868,N_5954);
and U6073 (N_6073,N_5811,N_5966);
nor U6074 (N_6074,N_5823,N_5866);
and U6075 (N_6075,N_5750,N_5835);
nand U6076 (N_6076,N_5828,N_5754);
or U6077 (N_6077,N_5910,N_5812);
nor U6078 (N_6078,N_5959,N_5843);
xnor U6079 (N_6079,N_5781,N_5830);
nor U6080 (N_6080,N_5957,N_5756);
or U6081 (N_6081,N_5876,N_5902);
or U6082 (N_6082,N_5805,N_5880);
and U6083 (N_6083,N_5934,N_5978);
nor U6084 (N_6084,N_5970,N_5784);
nor U6085 (N_6085,N_5994,N_5795);
nand U6086 (N_6086,N_5882,N_5751);
or U6087 (N_6087,N_5796,N_5819);
nand U6088 (N_6088,N_5764,N_5848);
and U6089 (N_6089,N_5945,N_5799);
or U6090 (N_6090,N_5833,N_5808);
xor U6091 (N_6091,N_5998,N_5770);
nor U6092 (N_6092,N_5923,N_5996);
or U6093 (N_6093,N_5977,N_5892);
and U6094 (N_6094,N_5965,N_5873);
or U6095 (N_6095,N_5767,N_5872);
xor U6096 (N_6096,N_5792,N_5935);
xnor U6097 (N_6097,N_5772,N_5897);
or U6098 (N_6098,N_5891,N_5943);
or U6099 (N_6099,N_5967,N_5992);
nor U6100 (N_6100,N_5855,N_5878);
nor U6101 (N_6101,N_5859,N_5968);
nand U6102 (N_6102,N_5956,N_5933);
nor U6103 (N_6103,N_5829,N_5816);
and U6104 (N_6104,N_5901,N_5958);
or U6105 (N_6105,N_5936,N_5752);
nor U6106 (N_6106,N_5888,N_5987);
nor U6107 (N_6107,N_5955,N_5824);
nand U6108 (N_6108,N_5753,N_5963);
xor U6109 (N_6109,N_5839,N_5842);
xor U6110 (N_6110,N_5831,N_5788);
nor U6111 (N_6111,N_5976,N_5793);
and U6112 (N_6112,N_5879,N_5865);
nand U6113 (N_6113,N_5881,N_5944);
nand U6114 (N_6114,N_5920,N_5763);
xnor U6115 (N_6115,N_5960,N_5938);
and U6116 (N_6116,N_5778,N_5946);
or U6117 (N_6117,N_5948,N_5961);
and U6118 (N_6118,N_5983,N_5898);
xor U6119 (N_6119,N_5780,N_5847);
nor U6120 (N_6120,N_5757,N_5789);
nor U6121 (N_6121,N_5755,N_5854);
nor U6122 (N_6122,N_5941,N_5951);
and U6123 (N_6123,N_5877,N_5826);
xor U6124 (N_6124,N_5899,N_5905);
nor U6125 (N_6125,N_5945,N_5810);
nand U6126 (N_6126,N_5894,N_5843);
nor U6127 (N_6127,N_5775,N_5998);
xnor U6128 (N_6128,N_5982,N_5794);
and U6129 (N_6129,N_5773,N_5983);
and U6130 (N_6130,N_5799,N_5997);
nand U6131 (N_6131,N_5905,N_5816);
and U6132 (N_6132,N_5996,N_5910);
nor U6133 (N_6133,N_5940,N_5915);
nand U6134 (N_6134,N_5848,N_5909);
and U6135 (N_6135,N_5833,N_5820);
xnor U6136 (N_6136,N_5877,N_5979);
nor U6137 (N_6137,N_5874,N_5754);
xor U6138 (N_6138,N_5826,N_5854);
nand U6139 (N_6139,N_5764,N_5825);
nor U6140 (N_6140,N_5895,N_5858);
and U6141 (N_6141,N_5841,N_5868);
nor U6142 (N_6142,N_5759,N_5832);
xor U6143 (N_6143,N_5777,N_5961);
nand U6144 (N_6144,N_5857,N_5764);
nor U6145 (N_6145,N_5845,N_5964);
nand U6146 (N_6146,N_5803,N_5762);
and U6147 (N_6147,N_5928,N_5818);
xor U6148 (N_6148,N_5898,N_5955);
or U6149 (N_6149,N_5788,N_5980);
xnor U6150 (N_6150,N_5790,N_5980);
xor U6151 (N_6151,N_5983,N_5850);
and U6152 (N_6152,N_5924,N_5947);
nand U6153 (N_6153,N_5804,N_5759);
and U6154 (N_6154,N_5945,N_5750);
or U6155 (N_6155,N_5934,N_5803);
nand U6156 (N_6156,N_5913,N_5940);
and U6157 (N_6157,N_5936,N_5930);
nand U6158 (N_6158,N_5863,N_5784);
nor U6159 (N_6159,N_5927,N_5969);
xor U6160 (N_6160,N_5922,N_5942);
xnor U6161 (N_6161,N_5783,N_5805);
xnor U6162 (N_6162,N_5822,N_5984);
and U6163 (N_6163,N_5845,N_5823);
xnor U6164 (N_6164,N_5785,N_5868);
or U6165 (N_6165,N_5897,N_5773);
or U6166 (N_6166,N_5941,N_5829);
nand U6167 (N_6167,N_5838,N_5957);
nand U6168 (N_6168,N_5980,N_5875);
xor U6169 (N_6169,N_5826,N_5770);
nor U6170 (N_6170,N_5886,N_5857);
or U6171 (N_6171,N_5989,N_5769);
nor U6172 (N_6172,N_5971,N_5868);
or U6173 (N_6173,N_5776,N_5847);
and U6174 (N_6174,N_5877,N_5794);
nor U6175 (N_6175,N_5811,N_5792);
nor U6176 (N_6176,N_5857,N_5953);
nor U6177 (N_6177,N_5841,N_5999);
nand U6178 (N_6178,N_5931,N_5880);
xnor U6179 (N_6179,N_5824,N_5809);
xnor U6180 (N_6180,N_5875,N_5977);
and U6181 (N_6181,N_5788,N_5778);
and U6182 (N_6182,N_5905,N_5882);
nand U6183 (N_6183,N_5793,N_5980);
and U6184 (N_6184,N_5994,N_5900);
nand U6185 (N_6185,N_5900,N_5834);
and U6186 (N_6186,N_5866,N_5945);
nand U6187 (N_6187,N_5913,N_5871);
and U6188 (N_6188,N_5976,N_5958);
nand U6189 (N_6189,N_5823,N_5834);
nor U6190 (N_6190,N_5952,N_5853);
nor U6191 (N_6191,N_5845,N_5768);
and U6192 (N_6192,N_5903,N_5755);
and U6193 (N_6193,N_5780,N_5779);
or U6194 (N_6194,N_5822,N_5917);
nor U6195 (N_6195,N_5941,N_5933);
nand U6196 (N_6196,N_5969,N_5870);
or U6197 (N_6197,N_5772,N_5878);
and U6198 (N_6198,N_5979,N_5911);
or U6199 (N_6199,N_5751,N_5766);
and U6200 (N_6200,N_5839,N_5954);
or U6201 (N_6201,N_5831,N_5884);
nand U6202 (N_6202,N_5777,N_5974);
and U6203 (N_6203,N_5908,N_5858);
nand U6204 (N_6204,N_5934,N_5880);
xnor U6205 (N_6205,N_5932,N_5844);
nor U6206 (N_6206,N_5868,N_5952);
and U6207 (N_6207,N_5907,N_5948);
xor U6208 (N_6208,N_5858,N_5874);
nor U6209 (N_6209,N_5949,N_5752);
xor U6210 (N_6210,N_5763,N_5960);
and U6211 (N_6211,N_5859,N_5907);
or U6212 (N_6212,N_5936,N_5890);
and U6213 (N_6213,N_5996,N_5887);
and U6214 (N_6214,N_5860,N_5943);
xor U6215 (N_6215,N_5829,N_5971);
and U6216 (N_6216,N_5775,N_5884);
and U6217 (N_6217,N_5770,N_5888);
or U6218 (N_6218,N_5946,N_5949);
or U6219 (N_6219,N_5985,N_5849);
nor U6220 (N_6220,N_5912,N_5918);
nor U6221 (N_6221,N_5802,N_5918);
and U6222 (N_6222,N_5848,N_5806);
xor U6223 (N_6223,N_5971,N_5779);
nand U6224 (N_6224,N_5956,N_5986);
and U6225 (N_6225,N_5989,N_5795);
or U6226 (N_6226,N_5899,N_5929);
or U6227 (N_6227,N_5796,N_5974);
nor U6228 (N_6228,N_5847,N_5898);
xor U6229 (N_6229,N_5824,N_5790);
nand U6230 (N_6230,N_5995,N_5933);
xnor U6231 (N_6231,N_5768,N_5919);
nand U6232 (N_6232,N_5927,N_5953);
and U6233 (N_6233,N_5876,N_5868);
or U6234 (N_6234,N_5789,N_5849);
xor U6235 (N_6235,N_5801,N_5914);
and U6236 (N_6236,N_5926,N_5859);
or U6237 (N_6237,N_5995,N_5885);
xnor U6238 (N_6238,N_5952,N_5811);
nand U6239 (N_6239,N_5766,N_5890);
nor U6240 (N_6240,N_5980,N_5797);
nor U6241 (N_6241,N_5839,N_5805);
nor U6242 (N_6242,N_5752,N_5887);
nor U6243 (N_6243,N_5815,N_5833);
nand U6244 (N_6244,N_5926,N_5896);
nor U6245 (N_6245,N_5785,N_5789);
nor U6246 (N_6246,N_5845,N_5852);
xor U6247 (N_6247,N_5855,N_5834);
and U6248 (N_6248,N_5864,N_5760);
nor U6249 (N_6249,N_5911,N_5803);
and U6250 (N_6250,N_6101,N_6233);
and U6251 (N_6251,N_6016,N_6196);
xnor U6252 (N_6252,N_6045,N_6070);
nor U6253 (N_6253,N_6083,N_6041);
or U6254 (N_6254,N_6166,N_6159);
nand U6255 (N_6255,N_6200,N_6248);
and U6256 (N_6256,N_6210,N_6240);
nor U6257 (N_6257,N_6192,N_6181);
nand U6258 (N_6258,N_6130,N_6216);
xor U6259 (N_6259,N_6162,N_6209);
xor U6260 (N_6260,N_6220,N_6241);
nor U6261 (N_6261,N_6002,N_6039);
xor U6262 (N_6262,N_6054,N_6182);
nand U6263 (N_6263,N_6029,N_6112);
or U6264 (N_6264,N_6138,N_6154);
nand U6265 (N_6265,N_6214,N_6089);
nor U6266 (N_6266,N_6079,N_6151);
nand U6267 (N_6267,N_6064,N_6003);
and U6268 (N_6268,N_6051,N_6027);
or U6269 (N_6269,N_6219,N_6245);
and U6270 (N_6270,N_6174,N_6204);
nand U6271 (N_6271,N_6177,N_6131);
or U6272 (N_6272,N_6038,N_6024);
or U6273 (N_6273,N_6232,N_6031);
or U6274 (N_6274,N_6048,N_6156);
nand U6275 (N_6275,N_6008,N_6099);
and U6276 (N_6276,N_6218,N_6078);
nor U6277 (N_6277,N_6042,N_6132);
and U6278 (N_6278,N_6100,N_6224);
nor U6279 (N_6279,N_6212,N_6145);
nand U6280 (N_6280,N_6134,N_6186);
nand U6281 (N_6281,N_6060,N_6021);
xor U6282 (N_6282,N_6180,N_6193);
xor U6283 (N_6283,N_6116,N_6128);
xnor U6284 (N_6284,N_6102,N_6142);
and U6285 (N_6285,N_6197,N_6084);
xor U6286 (N_6286,N_6153,N_6006);
nor U6287 (N_6287,N_6032,N_6201);
nor U6288 (N_6288,N_6030,N_6000);
nand U6289 (N_6289,N_6242,N_6085);
nor U6290 (N_6290,N_6015,N_6103);
xor U6291 (N_6291,N_6081,N_6143);
and U6292 (N_6292,N_6184,N_6217);
and U6293 (N_6293,N_6043,N_6080);
nor U6294 (N_6294,N_6092,N_6237);
and U6295 (N_6295,N_6194,N_6234);
or U6296 (N_6296,N_6026,N_6111);
or U6297 (N_6297,N_6236,N_6071);
or U6298 (N_6298,N_6191,N_6185);
nor U6299 (N_6299,N_6033,N_6028);
nor U6300 (N_6300,N_6249,N_6239);
and U6301 (N_6301,N_6188,N_6001);
xnor U6302 (N_6302,N_6059,N_6198);
xnor U6303 (N_6303,N_6011,N_6175);
and U6304 (N_6304,N_6072,N_6222);
nor U6305 (N_6305,N_6007,N_6161);
xnor U6306 (N_6306,N_6140,N_6055);
and U6307 (N_6307,N_6195,N_6208);
nor U6308 (N_6308,N_6144,N_6058);
or U6309 (N_6309,N_6179,N_6020);
nand U6310 (N_6310,N_6004,N_6173);
xnor U6311 (N_6311,N_6109,N_6164);
and U6312 (N_6312,N_6090,N_6123);
xnor U6313 (N_6313,N_6013,N_6023);
and U6314 (N_6314,N_6129,N_6225);
or U6315 (N_6315,N_6235,N_6040);
nor U6316 (N_6316,N_6148,N_6057);
nor U6317 (N_6317,N_6095,N_6034);
nand U6318 (N_6318,N_6005,N_6213);
nor U6319 (N_6319,N_6127,N_6025);
nor U6320 (N_6320,N_6167,N_6187);
xor U6321 (N_6321,N_6049,N_6091);
nor U6322 (N_6322,N_6183,N_6066);
or U6323 (N_6323,N_6098,N_6076);
nor U6324 (N_6324,N_6247,N_6061);
nand U6325 (N_6325,N_6121,N_6065);
and U6326 (N_6326,N_6229,N_6152);
and U6327 (N_6327,N_6113,N_6238);
nand U6328 (N_6328,N_6178,N_6010);
xor U6329 (N_6329,N_6137,N_6149);
or U6330 (N_6330,N_6110,N_6163);
and U6331 (N_6331,N_6035,N_6115);
xor U6332 (N_6332,N_6014,N_6018);
xnor U6333 (N_6333,N_6075,N_6107);
or U6334 (N_6334,N_6108,N_6105);
nand U6335 (N_6335,N_6160,N_6147);
or U6336 (N_6336,N_6122,N_6125);
or U6337 (N_6337,N_6047,N_6221);
nor U6338 (N_6338,N_6022,N_6093);
or U6339 (N_6339,N_6136,N_6243);
nand U6340 (N_6340,N_6086,N_6189);
xnor U6341 (N_6341,N_6139,N_6087);
xnor U6342 (N_6342,N_6009,N_6052);
and U6343 (N_6343,N_6056,N_6176);
nor U6344 (N_6344,N_6206,N_6017);
and U6345 (N_6345,N_6228,N_6117);
nand U6346 (N_6346,N_6114,N_6157);
nand U6347 (N_6347,N_6012,N_6063);
xnor U6348 (N_6348,N_6202,N_6155);
xnor U6349 (N_6349,N_6133,N_6227);
nand U6350 (N_6350,N_6171,N_6207);
xnor U6351 (N_6351,N_6050,N_6062);
nor U6352 (N_6352,N_6074,N_6119);
and U6353 (N_6353,N_6126,N_6069);
nor U6354 (N_6354,N_6096,N_6068);
or U6355 (N_6355,N_6172,N_6077);
and U6356 (N_6356,N_6104,N_6044);
and U6357 (N_6357,N_6223,N_6141);
nor U6358 (N_6358,N_6168,N_6205);
nand U6359 (N_6359,N_6146,N_6037);
xnor U6360 (N_6360,N_6231,N_6199);
nand U6361 (N_6361,N_6124,N_6082);
xor U6362 (N_6362,N_6106,N_6203);
nand U6363 (N_6363,N_6019,N_6097);
or U6364 (N_6364,N_6158,N_6244);
or U6365 (N_6365,N_6046,N_6135);
nand U6366 (N_6366,N_6226,N_6190);
and U6367 (N_6367,N_6215,N_6211);
xor U6368 (N_6368,N_6165,N_6036);
xor U6369 (N_6369,N_6067,N_6169);
nand U6370 (N_6370,N_6230,N_6088);
or U6371 (N_6371,N_6053,N_6094);
xnor U6372 (N_6372,N_6073,N_6118);
nand U6373 (N_6373,N_6170,N_6246);
nor U6374 (N_6374,N_6150,N_6120);
nand U6375 (N_6375,N_6145,N_6178);
nand U6376 (N_6376,N_6236,N_6189);
or U6377 (N_6377,N_6040,N_6046);
nand U6378 (N_6378,N_6104,N_6015);
xor U6379 (N_6379,N_6063,N_6019);
nor U6380 (N_6380,N_6048,N_6164);
or U6381 (N_6381,N_6123,N_6155);
or U6382 (N_6382,N_6009,N_6158);
nor U6383 (N_6383,N_6040,N_6160);
nand U6384 (N_6384,N_6127,N_6012);
or U6385 (N_6385,N_6182,N_6142);
and U6386 (N_6386,N_6239,N_6233);
nand U6387 (N_6387,N_6194,N_6176);
or U6388 (N_6388,N_6053,N_6036);
nor U6389 (N_6389,N_6211,N_6182);
nor U6390 (N_6390,N_6231,N_6000);
and U6391 (N_6391,N_6035,N_6170);
nor U6392 (N_6392,N_6106,N_6144);
nand U6393 (N_6393,N_6050,N_6120);
and U6394 (N_6394,N_6108,N_6125);
nor U6395 (N_6395,N_6223,N_6069);
nor U6396 (N_6396,N_6049,N_6175);
or U6397 (N_6397,N_6111,N_6032);
or U6398 (N_6398,N_6038,N_6175);
xnor U6399 (N_6399,N_6246,N_6185);
nor U6400 (N_6400,N_6144,N_6127);
xnor U6401 (N_6401,N_6222,N_6106);
nand U6402 (N_6402,N_6019,N_6181);
and U6403 (N_6403,N_6238,N_6217);
nor U6404 (N_6404,N_6218,N_6195);
nand U6405 (N_6405,N_6021,N_6194);
or U6406 (N_6406,N_6010,N_6243);
nand U6407 (N_6407,N_6024,N_6169);
xnor U6408 (N_6408,N_6216,N_6220);
xor U6409 (N_6409,N_6189,N_6068);
or U6410 (N_6410,N_6080,N_6155);
xor U6411 (N_6411,N_6248,N_6023);
and U6412 (N_6412,N_6052,N_6174);
nor U6413 (N_6413,N_6029,N_6198);
nor U6414 (N_6414,N_6230,N_6212);
or U6415 (N_6415,N_6127,N_6219);
nor U6416 (N_6416,N_6087,N_6000);
or U6417 (N_6417,N_6067,N_6021);
xor U6418 (N_6418,N_6004,N_6082);
nand U6419 (N_6419,N_6059,N_6165);
or U6420 (N_6420,N_6030,N_6141);
nor U6421 (N_6421,N_6017,N_6166);
xor U6422 (N_6422,N_6245,N_6120);
and U6423 (N_6423,N_6016,N_6080);
and U6424 (N_6424,N_6155,N_6199);
xor U6425 (N_6425,N_6195,N_6153);
and U6426 (N_6426,N_6221,N_6110);
and U6427 (N_6427,N_6124,N_6237);
nor U6428 (N_6428,N_6129,N_6087);
xor U6429 (N_6429,N_6010,N_6097);
and U6430 (N_6430,N_6032,N_6090);
nand U6431 (N_6431,N_6038,N_6142);
and U6432 (N_6432,N_6090,N_6031);
xor U6433 (N_6433,N_6131,N_6135);
and U6434 (N_6434,N_6084,N_6072);
or U6435 (N_6435,N_6104,N_6230);
nand U6436 (N_6436,N_6068,N_6046);
and U6437 (N_6437,N_6062,N_6212);
nand U6438 (N_6438,N_6246,N_6119);
xor U6439 (N_6439,N_6142,N_6219);
nand U6440 (N_6440,N_6024,N_6166);
nor U6441 (N_6441,N_6068,N_6007);
nand U6442 (N_6442,N_6137,N_6100);
xor U6443 (N_6443,N_6231,N_6239);
xnor U6444 (N_6444,N_6060,N_6172);
nor U6445 (N_6445,N_6211,N_6069);
xnor U6446 (N_6446,N_6127,N_6236);
and U6447 (N_6447,N_6216,N_6132);
nor U6448 (N_6448,N_6010,N_6105);
nand U6449 (N_6449,N_6166,N_6011);
and U6450 (N_6450,N_6141,N_6064);
xor U6451 (N_6451,N_6087,N_6033);
xor U6452 (N_6452,N_6041,N_6230);
xnor U6453 (N_6453,N_6121,N_6199);
nand U6454 (N_6454,N_6049,N_6120);
nand U6455 (N_6455,N_6213,N_6241);
and U6456 (N_6456,N_6086,N_6019);
and U6457 (N_6457,N_6160,N_6158);
nor U6458 (N_6458,N_6013,N_6221);
nand U6459 (N_6459,N_6144,N_6143);
and U6460 (N_6460,N_6244,N_6066);
nor U6461 (N_6461,N_6041,N_6093);
and U6462 (N_6462,N_6173,N_6208);
nand U6463 (N_6463,N_6216,N_6078);
xor U6464 (N_6464,N_6037,N_6090);
nand U6465 (N_6465,N_6039,N_6166);
nand U6466 (N_6466,N_6122,N_6014);
nor U6467 (N_6467,N_6060,N_6034);
or U6468 (N_6468,N_6234,N_6212);
xnor U6469 (N_6469,N_6182,N_6013);
nor U6470 (N_6470,N_6084,N_6153);
or U6471 (N_6471,N_6158,N_6084);
or U6472 (N_6472,N_6168,N_6178);
nor U6473 (N_6473,N_6165,N_6157);
and U6474 (N_6474,N_6033,N_6052);
and U6475 (N_6475,N_6243,N_6069);
and U6476 (N_6476,N_6047,N_6026);
or U6477 (N_6477,N_6162,N_6082);
xor U6478 (N_6478,N_6039,N_6007);
nand U6479 (N_6479,N_6024,N_6093);
xnor U6480 (N_6480,N_6197,N_6179);
nand U6481 (N_6481,N_6080,N_6132);
nand U6482 (N_6482,N_6012,N_6100);
or U6483 (N_6483,N_6081,N_6065);
nor U6484 (N_6484,N_6213,N_6155);
nand U6485 (N_6485,N_6236,N_6058);
xor U6486 (N_6486,N_6069,N_6204);
nor U6487 (N_6487,N_6196,N_6092);
nand U6488 (N_6488,N_6198,N_6222);
xor U6489 (N_6489,N_6060,N_6152);
and U6490 (N_6490,N_6023,N_6171);
and U6491 (N_6491,N_6135,N_6114);
and U6492 (N_6492,N_6137,N_6199);
nor U6493 (N_6493,N_6131,N_6215);
nor U6494 (N_6494,N_6099,N_6145);
and U6495 (N_6495,N_6180,N_6086);
and U6496 (N_6496,N_6005,N_6063);
nand U6497 (N_6497,N_6106,N_6052);
and U6498 (N_6498,N_6068,N_6162);
xor U6499 (N_6499,N_6033,N_6036);
and U6500 (N_6500,N_6367,N_6369);
nor U6501 (N_6501,N_6265,N_6379);
and U6502 (N_6502,N_6330,N_6373);
nor U6503 (N_6503,N_6336,N_6411);
nor U6504 (N_6504,N_6387,N_6442);
xnor U6505 (N_6505,N_6472,N_6278);
or U6506 (N_6506,N_6497,N_6337);
xor U6507 (N_6507,N_6291,N_6466);
xnor U6508 (N_6508,N_6272,N_6421);
nor U6509 (N_6509,N_6434,N_6485);
nor U6510 (N_6510,N_6276,N_6308);
or U6511 (N_6511,N_6455,N_6293);
nand U6512 (N_6512,N_6295,N_6359);
nand U6513 (N_6513,N_6393,N_6462);
and U6514 (N_6514,N_6323,N_6324);
nor U6515 (N_6515,N_6381,N_6436);
nor U6516 (N_6516,N_6329,N_6396);
or U6517 (N_6517,N_6408,N_6332);
xnor U6518 (N_6518,N_6374,N_6261);
nand U6519 (N_6519,N_6481,N_6377);
nand U6520 (N_6520,N_6437,N_6496);
nand U6521 (N_6521,N_6457,N_6270);
xnor U6522 (N_6522,N_6380,N_6451);
xor U6523 (N_6523,N_6264,N_6383);
nor U6524 (N_6524,N_6486,N_6358);
and U6525 (N_6525,N_6288,N_6403);
and U6526 (N_6526,N_6334,N_6287);
or U6527 (N_6527,N_6430,N_6465);
and U6528 (N_6528,N_6453,N_6348);
nor U6529 (N_6529,N_6355,N_6290);
or U6530 (N_6530,N_6433,N_6494);
nor U6531 (N_6531,N_6353,N_6467);
or U6532 (N_6532,N_6346,N_6417);
xnor U6533 (N_6533,N_6476,N_6303);
or U6534 (N_6534,N_6309,N_6474);
xnor U6535 (N_6535,N_6452,N_6427);
nand U6536 (N_6536,N_6438,N_6252);
nor U6537 (N_6537,N_6286,N_6487);
nand U6538 (N_6538,N_6413,N_6370);
or U6539 (N_6539,N_6406,N_6328);
nor U6540 (N_6540,N_6274,N_6285);
xnor U6541 (N_6541,N_6339,N_6493);
and U6542 (N_6542,N_6464,N_6416);
or U6543 (N_6543,N_6304,N_6354);
or U6544 (N_6544,N_6326,N_6311);
nand U6545 (N_6545,N_6420,N_6371);
or U6546 (N_6546,N_6410,N_6356);
nand U6547 (N_6547,N_6297,N_6458);
nand U6548 (N_6548,N_6447,N_6492);
nand U6549 (N_6549,N_6321,N_6426);
or U6550 (N_6550,N_6357,N_6405);
and U6551 (N_6551,N_6267,N_6366);
nor U6552 (N_6552,N_6491,N_6350);
or U6553 (N_6553,N_6251,N_6402);
or U6554 (N_6554,N_6418,N_6269);
nor U6555 (N_6555,N_6386,N_6432);
nand U6556 (N_6556,N_6327,N_6266);
or U6557 (N_6557,N_6482,N_6384);
xnor U6558 (N_6558,N_6262,N_6435);
and U6559 (N_6559,N_6372,N_6347);
nor U6560 (N_6560,N_6407,N_6382);
nor U6561 (N_6561,N_6422,N_6448);
nand U6562 (N_6562,N_6463,N_6443);
or U6563 (N_6563,N_6250,N_6376);
nand U6564 (N_6564,N_6343,N_6282);
nor U6565 (N_6565,N_6310,N_6361);
xor U6566 (N_6566,N_6306,N_6419);
and U6567 (N_6567,N_6449,N_6341);
nand U6568 (N_6568,N_6268,N_6389);
or U6569 (N_6569,N_6319,N_6298);
nand U6570 (N_6570,N_6483,N_6456);
and U6571 (N_6571,N_6469,N_6489);
or U6572 (N_6572,N_6445,N_6320);
xor U6573 (N_6573,N_6335,N_6484);
and U6574 (N_6574,N_6409,N_6260);
xor U6575 (N_6575,N_6375,N_6385);
nand U6576 (N_6576,N_6314,N_6351);
nor U6577 (N_6577,N_6271,N_6255);
or U6578 (N_6578,N_6280,N_6400);
xor U6579 (N_6579,N_6461,N_6344);
or U6580 (N_6580,N_6399,N_6296);
nand U6581 (N_6581,N_6460,N_6360);
and U6582 (N_6582,N_6284,N_6391);
and U6583 (N_6583,N_6352,N_6440);
xor U6584 (N_6584,N_6257,N_6302);
and U6585 (N_6585,N_6490,N_6412);
or U6586 (N_6586,N_6301,N_6363);
or U6587 (N_6587,N_6470,N_6283);
nor U6588 (N_6588,N_6415,N_6459);
xor U6589 (N_6589,N_6256,N_6258);
xnor U6590 (N_6590,N_6368,N_6477);
nand U6591 (N_6591,N_6475,N_6404);
and U6592 (N_6592,N_6431,N_6499);
and U6593 (N_6593,N_6479,N_6253);
and U6594 (N_6594,N_6279,N_6349);
xor U6595 (N_6595,N_6277,N_6392);
or U6596 (N_6596,N_6313,N_6345);
or U6597 (N_6597,N_6300,N_6468);
xnor U6598 (N_6598,N_6441,N_6444);
and U6599 (N_6599,N_6331,N_6325);
nor U6600 (N_6600,N_6281,N_6378);
nor U6601 (N_6601,N_6273,N_6401);
xor U6602 (N_6602,N_6394,N_6340);
and U6603 (N_6603,N_6388,N_6275);
and U6604 (N_6604,N_6307,N_6471);
nor U6605 (N_6605,N_6424,N_6259);
or U6606 (N_6606,N_6450,N_6478);
or U6607 (N_6607,N_6473,N_6254);
xor U6608 (N_6608,N_6398,N_6480);
nor U6609 (N_6609,N_6312,N_6390);
nor U6610 (N_6610,N_6498,N_6425);
nand U6611 (N_6611,N_6263,N_6305);
nand U6612 (N_6612,N_6362,N_6364);
xnor U6613 (N_6613,N_6316,N_6322);
nor U6614 (N_6614,N_6318,N_6439);
xnor U6615 (N_6615,N_6289,N_6299);
and U6616 (N_6616,N_6342,N_6338);
and U6617 (N_6617,N_6429,N_6333);
xnor U6618 (N_6618,N_6495,N_6428);
or U6619 (N_6619,N_6294,N_6414);
or U6620 (N_6620,N_6292,N_6454);
and U6621 (N_6621,N_6423,N_6488);
nand U6622 (N_6622,N_6446,N_6315);
xnor U6623 (N_6623,N_6365,N_6317);
xnor U6624 (N_6624,N_6397,N_6395);
or U6625 (N_6625,N_6476,N_6403);
nand U6626 (N_6626,N_6364,N_6304);
and U6627 (N_6627,N_6252,N_6424);
and U6628 (N_6628,N_6260,N_6476);
or U6629 (N_6629,N_6398,N_6470);
and U6630 (N_6630,N_6278,N_6347);
or U6631 (N_6631,N_6301,N_6457);
xnor U6632 (N_6632,N_6401,N_6390);
nor U6633 (N_6633,N_6321,N_6303);
and U6634 (N_6634,N_6435,N_6271);
nand U6635 (N_6635,N_6294,N_6311);
or U6636 (N_6636,N_6252,N_6327);
xnor U6637 (N_6637,N_6267,N_6462);
and U6638 (N_6638,N_6378,N_6250);
or U6639 (N_6639,N_6436,N_6489);
xor U6640 (N_6640,N_6291,N_6289);
xnor U6641 (N_6641,N_6253,N_6427);
or U6642 (N_6642,N_6475,N_6465);
nand U6643 (N_6643,N_6494,N_6270);
and U6644 (N_6644,N_6390,N_6480);
nand U6645 (N_6645,N_6459,N_6330);
or U6646 (N_6646,N_6360,N_6338);
nor U6647 (N_6647,N_6498,N_6364);
nand U6648 (N_6648,N_6460,N_6318);
nor U6649 (N_6649,N_6272,N_6357);
nand U6650 (N_6650,N_6324,N_6477);
nand U6651 (N_6651,N_6325,N_6316);
nand U6652 (N_6652,N_6381,N_6368);
nand U6653 (N_6653,N_6365,N_6492);
or U6654 (N_6654,N_6370,N_6353);
xnor U6655 (N_6655,N_6294,N_6438);
or U6656 (N_6656,N_6370,N_6489);
nor U6657 (N_6657,N_6273,N_6355);
nor U6658 (N_6658,N_6311,N_6340);
xnor U6659 (N_6659,N_6468,N_6333);
nand U6660 (N_6660,N_6456,N_6448);
or U6661 (N_6661,N_6371,N_6277);
nand U6662 (N_6662,N_6480,N_6300);
nor U6663 (N_6663,N_6334,N_6262);
or U6664 (N_6664,N_6340,N_6427);
or U6665 (N_6665,N_6468,N_6295);
and U6666 (N_6666,N_6476,N_6394);
xnor U6667 (N_6667,N_6321,N_6414);
and U6668 (N_6668,N_6268,N_6274);
and U6669 (N_6669,N_6415,N_6255);
nor U6670 (N_6670,N_6425,N_6354);
and U6671 (N_6671,N_6413,N_6405);
or U6672 (N_6672,N_6391,N_6271);
and U6673 (N_6673,N_6353,N_6333);
or U6674 (N_6674,N_6305,N_6402);
or U6675 (N_6675,N_6252,N_6362);
nor U6676 (N_6676,N_6420,N_6428);
or U6677 (N_6677,N_6280,N_6389);
and U6678 (N_6678,N_6350,N_6402);
or U6679 (N_6679,N_6285,N_6253);
and U6680 (N_6680,N_6386,N_6370);
nor U6681 (N_6681,N_6384,N_6348);
and U6682 (N_6682,N_6438,N_6264);
xor U6683 (N_6683,N_6415,N_6315);
and U6684 (N_6684,N_6267,N_6384);
nor U6685 (N_6685,N_6376,N_6261);
or U6686 (N_6686,N_6287,N_6488);
and U6687 (N_6687,N_6466,N_6253);
and U6688 (N_6688,N_6357,N_6397);
or U6689 (N_6689,N_6316,N_6410);
nand U6690 (N_6690,N_6366,N_6405);
xnor U6691 (N_6691,N_6391,N_6396);
and U6692 (N_6692,N_6383,N_6470);
nand U6693 (N_6693,N_6344,N_6445);
nand U6694 (N_6694,N_6440,N_6433);
nor U6695 (N_6695,N_6410,N_6470);
nor U6696 (N_6696,N_6265,N_6253);
nand U6697 (N_6697,N_6415,N_6445);
nand U6698 (N_6698,N_6305,N_6401);
and U6699 (N_6699,N_6446,N_6403);
xnor U6700 (N_6700,N_6324,N_6316);
or U6701 (N_6701,N_6420,N_6400);
nor U6702 (N_6702,N_6375,N_6329);
nor U6703 (N_6703,N_6434,N_6424);
xor U6704 (N_6704,N_6462,N_6381);
xor U6705 (N_6705,N_6386,N_6385);
nor U6706 (N_6706,N_6289,N_6265);
or U6707 (N_6707,N_6326,N_6377);
and U6708 (N_6708,N_6319,N_6281);
nand U6709 (N_6709,N_6390,N_6363);
xnor U6710 (N_6710,N_6281,N_6458);
or U6711 (N_6711,N_6427,N_6321);
nand U6712 (N_6712,N_6370,N_6267);
nand U6713 (N_6713,N_6438,N_6285);
nor U6714 (N_6714,N_6266,N_6350);
and U6715 (N_6715,N_6276,N_6368);
and U6716 (N_6716,N_6305,N_6350);
or U6717 (N_6717,N_6392,N_6309);
xor U6718 (N_6718,N_6479,N_6334);
xnor U6719 (N_6719,N_6291,N_6412);
xor U6720 (N_6720,N_6383,N_6445);
nor U6721 (N_6721,N_6444,N_6330);
nor U6722 (N_6722,N_6313,N_6402);
xnor U6723 (N_6723,N_6492,N_6499);
and U6724 (N_6724,N_6437,N_6386);
xor U6725 (N_6725,N_6453,N_6309);
nand U6726 (N_6726,N_6275,N_6329);
nand U6727 (N_6727,N_6341,N_6390);
or U6728 (N_6728,N_6472,N_6418);
nand U6729 (N_6729,N_6290,N_6422);
or U6730 (N_6730,N_6252,N_6444);
or U6731 (N_6731,N_6420,N_6397);
xor U6732 (N_6732,N_6263,N_6428);
or U6733 (N_6733,N_6440,N_6473);
nor U6734 (N_6734,N_6279,N_6312);
and U6735 (N_6735,N_6362,N_6418);
nor U6736 (N_6736,N_6485,N_6320);
nor U6737 (N_6737,N_6457,N_6267);
and U6738 (N_6738,N_6383,N_6354);
or U6739 (N_6739,N_6417,N_6320);
and U6740 (N_6740,N_6271,N_6329);
nand U6741 (N_6741,N_6308,N_6427);
xor U6742 (N_6742,N_6424,N_6354);
and U6743 (N_6743,N_6300,N_6497);
and U6744 (N_6744,N_6377,N_6395);
xor U6745 (N_6745,N_6262,N_6278);
xnor U6746 (N_6746,N_6341,N_6434);
and U6747 (N_6747,N_6264,N_6447);
nor U6748 (N_6748,N_6316,N_6398);
or U6749 (N_6749,N_6498,N_6450);
nand U6750 (N_6750,N_6549,N_6628);
and U6751 (N_6751,N_6603,N_6523);
xnor U6752 (N_6752,N_6653,N_6596);
xnor U6753 (N_6753,N_6651,N_6577);
or U6754 (N_6754,N_6691,N_6660);
nor U6755 (N_6755,N_6693,N_6630);
and U6756 (N_6756,N_6624,N_6532);
or U6757 (N_6757,N_6568,N_6696);
nor U6758 (N_6758,N_6530,N_6527);
nand U6759 (N_6759,N_6519,N_6698);
xnor U6760 (N_6760,N_6725,N_6697);
nor U6761 (N_6761,N_6548,N_6672);
or U6762 (N_6762,N_6609,N_6613);
or U6763 (N_6763,N_6553,N_6644);
nand U6764 (N_6764,N_6719,N_6614);
xor U6765 (N_6765,N_6703,N_6610);
or U6766 (N_6766,N_6734,N_6701);
nand U6767 (N_6767,N_6678,N_6506);
nand U6768 (N_6768,N_6726,N_6745);
nand U6769 (N_6769,N_6522,N_6733);
or U6770 (N_6770,N_6702,N_6547);
nand U6771 (N_6771,N_6720,N_6704);
and U6772 (N_6772,N_6747,N_6552);
nor U6773 (N_6773,N_6604,N_6543);
xor U6774 (N_6774,N_6668,N_6667);
nand U6775 (N_6775,N_6625,N_6557);
nand U6776 (N_6776,N_6588,N_6615);
or U6777 (N_6777,N_6652,N_6544);
nand U6778 (N_6778,N_6599,N_6714);
xor U6779 (N_6779,N_6744,N_6647);
and U6780 (N_6780,N_6605,N_6677);
or U6781 (N_6781,N_6535,N_6724);
or U6782 (N_6782,N_6546,N_6616);
and U6783 (N_6783,N_6511,N_6641);
nand U6784 (N_6784,N_6593,N_6686);
nand U6785 (N_6785,N_6526,N_6556);
nand U6786 (N_6786,N_6607,N_6512);
nor U6787 (N_6787,N_6654,N_6658);
xor U6788 (N_6788,N_6514,N_6537);
nor U6789 (N_6789,N_6580,N_6534);
xor U6790 (N_6790,N_6674,N_6595);
and U6791 (N_6791,N_6562,N_6579);
and U6792 (N_6792,N_6505,N_6611);
and U6793 (N_6793,N_6706,N_6554);
or U6794 (N_6794,N_6594,N_6707);
or U6795 (N_6795,N_6575,N_6578);
nand U6796 (N_6796,N_6673,N_6528);
and U6797 (N_6797,N_6560,N_6656);
or U6798 (N_6798,N_6550,N_6619);
nor U6799 (N_6799,N_6541,N_6558);
or U6800 (N_6800,N_6569,N_6705);
or U6801 (N_6801,N_6680,N_6679);
nor U6802 (N_6802,N_6529,N_6748);
nor U6803 (N_6803,N_6640,N_6638);
nand U6804 (N_6804,N_6617,N_6730);
and U6805 (N_6805,N_6699,N_6570);
nand U6806 (N_6806,N_6684,N_6713);
and U6807 (N_6807,N_6631,N_6539);
xor U6808 (N_6808,N_6695,N_6500);
or U6809 (N_6809,N_6700,N_6559);
and U6810 (N_6810,N_6520,N_6587);
and U6811 (N_6811,N_6662,N_6735);
nor U6812 (N_6812,N_6676,N_6510);
nand U6813 (N_6813,N_6710,N_6592);
or U6814 (N_6814,N_6589,N_6634);
and U6815 (N_6815,N_6643,N_6565);
and U6816 (N_6816,N_6716,N_6688);
nand U6817 (N_6817,N_6708,N_6622);
nand U6818 (N_6818,N_6712,N_6533);
nand U6819 (N_6819,N_6682,N_6685);
xnor U6820 (N_6820,N_6524,N_6602);
and U6821 (N_6821,N_6642,N_6737);
nand U6822 (N_6822,N_6635,N_6743);
or U6823 (N_6823,N_6501,N_6612);
or U6824 (N_6824,N_6671,N_6650);
nor U6825 (N_6825,N_6591,N_6606);
xnor U6826 (N_6826,N_6709,N_6563);
nand U6827 (N_6827,N_6664,N_6632);
and U6828 (N_6828,N_6749,N_6681);
or U6829 (N_6829,N_6627,N_6608);
or U6830 (N_6830,N_6503,N_6525);
nand U6831 (N_6831,N_6620,N_6732);
xnor U6832 (N_6832,N_6618,N_6661);
and U6833 (N_6833,N_6600,N_6740);
nand U6834 (N_6834,N_6584,N_6746);
or U6835 (N_6835,N_6741,N_6645);
or U6836 (N_6836,N_6646,N_6637);
or U6837 (N_6837,N_6648,N_6542);
and U6838 (N_6838,N_6742,N_6728);
xnor U6839 (N_6839,N_6518,N_6517);
nand U6840 (N_6840,N_6736,N_6683);
nor U6841 (N_6841,N_6636,N_6626);
xnor U6842 (N_6842,N_6540,N_6586);
xnor U6843 (N_6843,N_6576,N_6687);
and U6844 (N_6844,N_6555,N_6536);
nor U6845 (N_6845,N_6690,N_6582);
xor U6846 (N_6846,N_6561,N_6598);
and U6847 (N_6847,N_6567,N_6675);
and U6848 (N_6848,N_6739,N_6574);
xnor U6849 (N_6849,N_6572,N_6721);
nor U6850 (N_6850,N_6649,N_6692);
and U6851 (N_6851,N_6513,N_6669);
nand U6852 (N_6852,N_6666,N_6718);
or U6853 (N_6853,N_6723,N_6502);
xor U6854 (N_6854,N_6665,N_6639);
nor U6855 (N_6855,N_6621,N_6581);
and U6856 (N_6856,N_6657,N_6689);
and U6857 (N_6857,N_6545,N_6623);
or U6858 (N_6858,N_6515,N_6715);
xnor U6859 (N_6859,N_6585,N_6711);
xnor U6860 (N_6860,N_6727,N_6504);
and U6861 (N_6861,N_6722,N_6531);
nand U6862 (N_6862,N_6566,N_6508);
and U6863 (N_6863,N_6633,N_6694);
or U6864 (N_6864,N_6571,N_6729);
nand U6865 (N_6865,N_6509,N_6516);
nand U6866 (N_6866,N_6670,N_6717);
xor U6867 (N_6867,N_6564,N_6507);
or U6868 (N_6868,N_6583,N_6521);
or U6869 (N_6869,N_6590,N_6629);
nand U6870 (N_6870,N_6601,N_6659);
nor U6871 (N_6871,N_6731,N_6663);
nor U6872 (N_6872,N_6573,N_6551);
nor U6873 (N_6873,N_6738,N_6655);
and U6874 (N_6874,N_6597,N_6538);
nand U6875 (N_6875,N_6598,N_6503);
and U6876 (N_6876,N_6595,N_6575);
nand U6877 (N_6877,N_6552,N_6545);
nor U6878 (N_6878,N_6569,N_6591);
nor U6879 (N_6879,N_6684,N_6716);
and U6880 (N_6880,N_6537,N_6558);
nand U6881 (N_6881,N_6545,N_6686);
nor U6882 (N_6882,N_6555,N_6503);
and U6883 (N_6883,N_6592,N_6573);
or U6884 (N_6884,N_6611,N_6603);
nor U6885 (N_6885,N_6721,N_6682);
xor U6886 (N_6886,N_6743,N_6592);
nor U6887 (N_6887,N_6746,N_6656);
xor U6888 (N_6888,N_6748,N_6570);
and U6889 (N_6889,N_6612,N_6744);
nand U6890 (N_6890,N_6733,N_6676);
and U6891 (N_6891,N_6623,N_6647);
xnor U6892 (N_6892,N_6608,N_6587);
xnor U6893 (N_6893,N_6575,N_6586);
and U6894 (N_6894,N_6616,N_6698);
or U6895 (N_6895,N_6551,N_6642);
nand U6896 (N_6896,N_6706,N_6700);
and U6897 (N_6897,N_6733,N_6509);
xor U6898 (N_6898,N_6716,N_6678);
nor U6899 (N_6899,N_6610,N_6548);
nand U6900 (N_6900,N_6695,N_6685);
nor U6901 (N_6901,N_6527,N_6656);
xnor U6902 (N_6902,N_6620,N_6624);
nor U6903 (N_6903,N_6651,N_6687);
xnor U6904 (N_6904,N_6740,N_6641);
nand U6905 (N_6905,N_6611,N_6598);
nor U6906 (N_6906,N_6736,N_6739);
or U6907 (N_6907,N_6656,N_6566);
or U6908 (N_6908,N_6570,N_6561);
or U6909 (N_6909,N_6563,N_6560);
xnor U6910 (N_6910,N_6531,N_6525);
nor U6911 (N_6911,N_6556,N_6651);
nor U6912 (N_6912,N_6567,N_6550);
or U6913 (N_6913,N_6586,N_6517);
xnor U6914 (N_6914,N_6688,N_6690);
nand U6915 (N_6915,N_6579,N_6686);
nor U6916 (N_6916,N_6719,N_6535);
or U6917 (N_6917,N_6674,N_6687);
nand U6918 (N_6918,N_6735,N_6669);
nor U6919 (N_6919,N_6729,N_6623);
nand U6920 (N_6920,N_6691,N_6653);
and U6921 (N_6921,N_6655,N_6745);
xnor U6922 (N_6922,N_6749,N_6525);
nor U6923 (N_6923,N_6500,N_6744);
nand U6924 (N_6924,N_6582,N_6627);
nor U6925 (N_6925,N_6508,N_6730);
or U6926 (N_6926,N_6522,N_6655);
and U6927 (N_6927,N_6742,N_6724);
nand U6928 (N_6928,N_6723,N_6710);
nor U6929 (N_6929,N_6560,N_6582);
nor U6930 (N_6930,N_6651,N_6692);
nand U6931 (N_6931,N_6621,N_6730);
and U6932 (N_6932,N_6639,N_6508);
or U6933 (N_6933,N_6701,N_6726);
nor U6934 (N_6934,N_6709,N_6686);
and U6935 (N_6935,N_6564,N_6734);
or U6936 (N_6936,N_6577,N_6713);
and U6937 (N_6937,N_6547,N_6662);
and U6938 (N_6938,N_6578,N_6531);
and U6939 (N_6939,N_6679,N_6550);
nand U6940 (N_6940,N_6600,N_6565);
and U6941 (N_6941,N_6597,N_6637);
nand U6942 (N_6942,N_6679,N_6729);
and U6943 (N_6943,N_6620,N_6576);
xor U6944 (N_6944,N_6564,N_6672);
xnor U6945 (N_6945,N_6681,N_6610);
nor U6946 (N_6946,N_6638,N_6623);
xnor U6947 (N_6947,N_6532,N_6674);
or U6948 (N_6948,N_6562,N_6647);
nand U6949 (N_6949,N_6530,N_6649);
and U6950 (N_6950,N_6651,N_6581);
and U6951 (N_6951,N_6679,N_6699);
and U6952 (N_6952,N_6634,N_6618);
or U6953 (N_6953,N_6708,N_6569);
xnor U6954 (N_6954,N_6573,N_6553);
xnor U6955 (N_6955,N_6521,N_6723);
nand U6956 (N_6956,N_6721,N_6510);
xnor U6957 (N_6957,N_6724,N_6735);
xor U6958 (N_6958,N_6547,N_6524);
or U6959 (N_6959,N_6673,N_6720);
and U6960 (N_6960,N_6547,N_6533);
xor U6961 (N_6961,N_6590,N_6632);
xnor U6962 (N_6962,N_6613,N_6626);
or U6963 (N_6963,N_6635,N_6705);
nor U6964 (N_6964,N_6745,N_6669);
and U6965 (N_6965,N_6735,N_6616);
or U6966 (N_6966,N_6658,N_6704);
or U6967 (N_6967,N_6697,N_6683);
or U6968 (N_6968,N_6736,N_6664);
or U6969 (N_6969,N_6575,N_6727);
xnor U6970 (N_6970,N_6622,N_6641);
nor U6971 (N_6971,N_6710,N_6588);
nand U6972 (N_6972,N_6552,N_6521);
nor U6973 (N_6973,N_6563,N_6545);
xnor U6974 (N_6974,N_6621,N_6671);
nand U6975 (N_6975,N_6542,N_6588);
and U6976 (N_6976,N_6546,N_6568);
xnor U6977 (N_6977,N_6520,N_6509);
xnor U6978 (N_6978,N_6502,N_6540);
nand U6979 (N_6979,N_6692,N_6606);
and U6980 (N_6980,N_6593,N_6573);
and U6981 (N_6981,N_6507,N_6666);
or U6982 (N_6982,N_6650,N_6590);
xor U6983 (N_6983,N_6741,N_6561);
nand U6984 (N_6984,N_6586,N_6557);
and U6985 (N_6985,N_6696,N_6529);
nand U6986 (N_6986,N_6739,N_6577);
nand U6987 (N_6987,N_6593,N_6669);
xor U6988 (N_6988,N_6638,N_6694);
and U6989 (N_6989,N_6714,N_6575);
nor U6990 (N_6990,N_6542,N_6742);
or U6991 (N_6991,N_6716,N_6665);
and U6992 (N_6992,N_6542,N_6509);
and U6993 (N_6993,N_6644,N_6544);
nand U6994 (N_6994,N_6594,N_6549);
xor U6995 (N_6995,N_6552,N_6587);
nor U6996 (N_6996,N_6617,N_6675);
and U6997 (N_6997,N_6706,N_6720);
or U6998 (N_6998,N_6711,N_6643);
xor U6999 (N_6999,N_6681,N_6746);
nand U7000 (N_7000,N_6816,N_6894);
or U7001 (N_7001,N_6952,N_6792);
or U7002 (N_7002,N_6796,N_6785);
or U7003 (N_7003,N_6804,N_6780);
nand U7004 (N_7004,N_6766,N_6859);
and U7005 (N_7005,N_6784,N_6813);
and U7006 (N_7006,N_6931,N_6820);
xnor U7007 (N_7007,N_6982,N_6830);
or U7008 (N_7008,N_6840,N_6868);
and U7009 (N_7009,N_6790,N_6872);
nor U7010 (N_7010,N_6918,N_6976);
and U7011 (N_7011,N_6902,N_6835);
and U7012 (N_7012,N_6980,N_6922);
nand U7013 (N_7013,N_6923,N_6850);
nand U7014 (N_7014,N_6983,N_6912);
nand U7015 (N_7015,N_6809,N_6885);
and U7016 (N_7016,N_6782,N_6936);
xnor U7017 (N_7017,N_6765,N_6843);
xor U7018 (N_7018,N_6966,N_6846);
nor U7019 (N_7019,N_6951,N_6934);
xor U7020 (N_7020,N_6879,N_6803);
nor U7021 (N_7021,N_6751,N_6960);
or U7022 (N_7022,N_6888,N_6834);
and U7023 (N_7023,N_6783,N_6896);
nand U7024 (N_7024,N_6778,N_6866);
nor U7025 (N_7025,N_6979,N_6787);
xor U7026 (N_7026,N_6965,N_6895);
nor U7027 (N_7027,N_6821,N_6818);
xor U7028 (N_7028,N_6822,N_6954);
nand U7029 (N_7029,N_6793,N_6768);
and U7030 (N_7030,N_6975,N_6777);
xor U7031 (N_7031,N_6985,N_6926);
xor U7032 (N_7032,N_6769,N_6761);
nor U7033 (N_7033,N_6984,N_6958);
and U7034 (N_7034,N_6771,N_6986);
xnor U7035 (N_7035,N_6935,N_6759);
and U7036 (N_7036,N_6797,N_6849);
nand U7037 (N_7037,N_6915,N_6947);
nand U7038 (N_7038,N_6824,N_6832);
nand U7039 (N_7039,N_6950,N_6837);
and U7040 (N_7040,N_6946,N_6869);
xnor U7041 (N_7041,N_6973,N_6924);
or U7042 (N_7042,N_6997,N_6929);
or U7043 (N_7043,N_6981,N_6779);
nand U7044 (N_7044,N_6905,N_6842);
xnor U7045 (N_7045,N_6776,N_6827);
nand U7046 (N_7046,N_6774,N_6959);
nand U7047 (N_7047,N_6961,N_6917);
nor U7048 (N_7048,N_6970,N_6874);
or U7049 (N_7049,N_6811,N_6755);
nand U7050 (N_7050,N_6999,N_6773);
xnor U7051 (N_7051,N_6848,N_6826);
xnor U7052 (N_7052,N_6873,N_6753);
xor U7053 (N_7053,N_6889,N_6855);
or U7054 (N_7054,N_6943,N_6908);
and U7055 (N_7055,N_6756,N_6991);
and U7056 (N_7056,N_6786,N_6993);
nand U7057 (N_7057,N_6948,N_6847);
nand U7058 (N_7058,N_6857,N_6863);
or U7059 (N_7059,N_6938,N_6928);
or U7060 (N_7060,N_6914,N_6978);
nor U7061 (N_7061,N_6812,N_6994);
nand U7062 (N_7062,N_6845,N_6899);
xor U7063 (N_7063,N_6844,N_6903);
and U7064 (N_7064,N_6957,N_6897);
or U7065 (N_7065,N_6906,N_6831);
nor U7066 (N_7066,N_6937,N_6758);
and U7067 (N_7067,N_6875,N_6851);
or U7068 (N_7068,N_6987,N_6815);
nand U7069 (N_7069,N_6968,N_6838);
nand U7070 (N_7070,N_6916,N_6825);
nor U7071 (N_7071,N_6884,N_6932);
nand U7072 (N_7072,N_6967,N_6750);
and U7073 (N_7073,N_6963,N_6865);
or U7074 (N_7074,N_6799,N_6883);
nor U7075 (N_7075,N_6805,N_6921);
and U7076 (N_7076,N_6760,N_6870);
nand U7077 (N_7077,N_6964,N_6864);
or U7078 (N_7078,N_6819,N_6904);
nand U7079 (N_7079,N_6886,N_6828);
nor U7080 (N_7080,N_6925,N_6881);
and U7081 (N_7081,N_6930,N_6798);
nand U7082 (N_7082,N_6927,N_6996);
nand U7083 (N_7083,N_6953,N_6789);
and U7084 (N_7084,N_6992,N_6770);
or U7085 (N_7085,N_6969,N_6808);
nor U7086 (N_7086,N_6945,N_6757);
xnor U7087 (N_7087,N_6882,N_6802);
xor U7088 (N_7088,N_6763,N_6907);
and U7089 (N_7089,N_6949,N_6762);
and U7090 (N_7090,N_6829,N_6781);
or U7091 (N_7091,N_6800,N_6910);
or U7092 (N_7092,N_6988,N_6880);
and U7093 (N_7093,N_6795,N_6841);
or U7094 (N_7094,N_6807,N_6887);
or U7095 (N_7095,N_6767,N_6913);
nor U7096 (N_7096,N_6764,N_6911);
or U7097 (N_7097,N_6977,N_6974);
nor U7098 (N_7098,N_6775,N_6867);
and U7099 (N_7099,N_6971,N_6933);
xor U7100 (N_7100,N_6939,N_6853);
nand U7101 (N_7101,N_6754,N_6989);
and U7102 (N_7102,N_6944,N_6920);
xnor U7103 (N_7103,N_6852,N_6810);
and U7104 (N_7104,N_6876,N_6891);
or U7105 (N_7105,N_6955,N_6801);
or U7106 (N_7106,N_6909,N_6814);
xnor U7107 (N_7107,N_6890,N_6854);
xnor U7108 (N_7108,N_6878,N_6861);
nand U7109 (N_7109,N_6900,N_6839);
nand U7110 (N_7110,N_6788,N_6871);
or U7111 (N_7111,N_6901,N_6856);
nor U7112 (N_7112,N_6877,N_6962);
nand U7113 (N_7113,N_6998,N_6858);
nor U7114 (N_7114,N_6862,N_6990);
or U7115 (N_7115,N_6972,N_6823);
or U7116 (N_7116,N_6772,N_6898);
nand U7117 (N_7117,N_6836,N_6817);
nor U7118 (N_7118,N_6941,N_6791);
xor U7119 (N_7119,N_6806,N_6995);
xnor U7120 (N_7120,N_6942,N_6940);
or U7121 (N_7121,N_6919,N_6752);
or U7122 (N_7122,N_6833,N_6956);
and U7123 (N_7123,N_6893,N_6794);
and U7124 (N_7124,N_6860,N_6892);
or U7125 (N_7125,N_6755,N_6775);
nand U7126 (N_7126,N_6908,N_6927);
xor U7127 (N_7127,N_6784,N_6891);
or U7128 (N_7128,N_6891,N_6774);
and U7129 (N_7129,N_6977,N_6900);
xnor U7130 (N_7130,N_6934,N_6857);
nor U7131 (N_7131,N_6758,N_6872);
nor U7132 (N_7132,N_6920,N_6924);
nand U7133 (N_7133,N_6777,N_6917);
nor U7134 (N_7134,N_6963,N_6868);
and U7135 (N_7135,N_6892,N_6990);
and U7136 (N_7136,N_6840,N_6878);
nor U7137 (N_7137,N_6861,N_6852);
or U7138 (N_7138,N_6886,N_6814);
nand U7139 (N_7139,N_6893,N_6928);
nand U7140 (N_7140,N_6943,N_6942);
or U7141 (N_7141,N_6782,N_6813);
or U7142 (N_7142,N_6820,N_6989);
and U7143 (N_7143,N_6942,N_6852);
or U7144 (N_7144,N_6820,N_6861);
xnor U7145 (N_7145,N_6986,N_6922);
nand U7146 (N_7146,N_6812,N_6881);
xnor U7147 (N_7147,N_6793,N_6896);
or U7148 (N_7148,N_6841,N_6970);
or U7149 (N_7149,N_6988,N_6912);
nand U7150 (N_7150,N_6933,N_6928);
nor U7151 (N_7151,N_6816,N_6851);
nor U7152 (N_7152,N_6919,N_6757);
or U7153 (N_7153,N_6887,N_6952);
xnor U7154 (N_7154,N_6947,N_6861);
xnor U7155 (N_7155,N_6804,N_6826);
nor U7156 (N_7156,N_6867,N_6931);
nor U7157 (N_7157,N_6789,N_6970);
or U7158 (N_7158,N_6991,N_6909);
xor U7159 (N_7159,N_6767,N_6754);
nor U7160 (N_7160,N_6898,N_6967);
xnor U7161 (N_7161,N_6791,N_6768);
nor U7162 (N_7162,N_6828,N_6981);
xnor U7163 (N_7163,N_6972,N_6967);
nand U7164 (N_7164,N_6809,N_6978);
nor U7165 (N_7165,N_6873,N_6843);
xnor U7166 (N_7166,N_6887,N_6913);
or U7167 (N_7167,N_6828,N_6941);
nor U7168 (N_7168,N_6966,N_6989);
xnor U7169 (N_7169,N_6857,N_6891);
xor U7170 (N_7170,N_6951,N_6883);
or U7171 (N_7171,N_6822,N_6827);
or U7172 (N_7172,N_6821,N_6801);
and U7173 (N_7173,N_6982,N_6987);
nand U7174 (N_7174,N_6770,N_6819);
nand U7175 (N_7175,N_6981,N_6989);
nand U7176 (N_7176,N_6797,N_6795);
or U7177 (N_7177,N_6820,N_6926);
or U7178 (N_7178,N_6750,N_6859);
nor U7179 (N_7179,N_6762,N_6890);
nand U7180 (N_7180,N_6968,N_6982);
nand U7181 (N_7181,N_6767,N_6780);
nand U7182 (N_7182,N_6865,N_6774);
or U7183 (N_7183,N_6860,N_6883);
xor U7184 (N_7184,N_6786,N_6828);
nor U7185 (N_7185,N_6839,N_6965);
or U7186 (N_7186,N_6936,N_6808);
nand U7187 (N_7187,N_6971,N_6886);
xnor U7188 (N_7188,N_6750,N_6959);
and U7189 (N_7189,N_6912,N_6787);
or U7190 (N_7190,N_6847,N_6766);
nor U7191 (N_7191,N_6868,N_6756);
or U7192 (N_7192,N_6810,N_6774);
nor U7193 (N_7193,N_6942,N_6975);
or U7194 (N_7194,N_6848,N_6946);
xor U7195 (N_7195,N_6810,N_6776);
nand U7196 (N_7196,N_6964,N_6865);
nand U7197 (N_7197,N_6923,N_6778);
nor U7198 (N_7198,N_6870,N_6890);
and U7199 (N_7199,N_6870,N_6837);
nand U7200 (N_7200,N_6897,N_6934);
or U7201 (N_7201,N_6987,N_6757);
xnor U7202 (N_7202,N_6981,N_6987);
xor U7203 (N_7203,N_6805,N_6781);
nor U7204 (N_7204,N_6800,N_6913);
nor U7205 (N_7205,N_6788,N_6948);
nor U7206 (N_7206,N_6889,N_6958);
nor U7207 (N_7207,N_6924,N_6758);
xnor U7208 (N_7208,N_6753,N_6976);
and U7209 (N_7209,N_6859,N_6978);
xnor U7210 (N_7210,N_6990,N_6802);
xnor U7211 (N_7211,N_6829,N_6977);
nand U7212 (N_7212,N_6775,N_6843);
nor U7213 (N_7213,N_6789,N_6813);
nand U7214 (N_7214,N_6768,N_6921);
nor U7215 (N_7215,N_6871,N_6762);
xnor U7216 (N_7216,N_6769,N_6908);
xor U7217 (N_7217,N_6825,N_6817);
nand U7218 (N_7218,N_6871,N_6988);
nand U7219 (N_7219,N_6782,N_6867);
and U7220 (N_7220,N_6964,N_6954);
or U7221 (N_7221,N_6901,N_6805);
xnor U7222 (N_7222,N_6762,N_6885);
nor U7223 (N_7223,N_6768,N_6758);
nand U7224 (N_7224,N_6890,N_6817);
and U7225 (N_7225,N_6817,N_6863);
nor U7226 (N_7226,N_6782,N_6847);
nand U7227 (N_7227,N_6973,N_6987);
nor U7228 (N_7228,N_6768,N_6888);
and U7229 (N_7229,N_6979,N_6806);
or U7230 (N_7230,N_6860,N_6931);
nand U7231 (N_7231,N_6820,N_6811);
nand U7232 (N_7232,N_6908,N_6795);
or U7233 (N_7233,N_6845,N_6831);
nor U7234 (N_7234,N_6931,N_6872);
nor U7235 (N_7235,N_6973,N_6813);
or U7236 (N_7236,N_6789,N_6978);
or U7237 (N_7237,N_6848,N_6799);
nand U7238 (N_7238,N_6800,N_6915);
or U7239 (N_7239,N_6960,N_6943);
xor U7240 (N_7240,N_6904,N_6810);
and U7241 (N_7241,N_6921,N_6974);
xor U7242 (N_7242,N_6809,N_6774);
xor U7243 (N_7243,N_6873,N_6967);
xnor U7244 (N_7244,N_6763,N_6817);
and U7245 (N_7245,N_6858,N_6755);
nand U7246 (N_7246,N_6903,N_6816);
nand U7247 (N_7247,N_6936,N_6840);
xor U7248 (N_7248,N_6978,N_6824);
xor U7249 (N_7249,N_6808,N_6819);
or U7250 (N_7250,N_7055,N_7119);
nor U7251 (N_7251,N_7016,N_7096);
or U7252 (N_7252,N_7073,N_7037);
xnor U7253 (N_7253,N_7174,N_7061);
or U7254 (N_7254,N_7018,N_7023);
or U7255 (N_7255,N_7208,N_7186);
nor U7256 (N_7256,N_7101,N_7029);
and U7257 (N_7257,N_7241,N_7113);
nor U7258 (N_7258,N_7194,N_7158);
nand U7259 (N_7259,N_7027,N_7100);
and U7260 (N_7260,N_7078,N_7072);
nand U7261 (N_7261,N_7170,N_7065);
or U7262 (N_7262,N_7229,N_7058);
and U7263 (N_7263,N_7070,N_7026);
and U7264 (N_7264,N_7031,N_7084);
and U7265 (N_7265,N_7021,N_7011);
xnor U7266 (N_7266,N_7066,N_7187);
nand U7267 (N_7267,N_7122,N_7039);
and U7268 (N_7268,N_7231,N_7213);
xor U7269 (N_7269,N_7198,N_7017);
nor U7270 (N_7270,N_7243,N_7233);
nand U7271 (N_7271,N_7242,N_7059);
xor U7272 (N_7272,N_7206,N_7125);
nand U7273 (N_7273,N_7034,N_7077);
and U7274 (N_7274,N_7162,N_7166);
xor U7275 (N_7275,N_7133,N_7216);
and U7276 (N_7276,N_7212,N_7217);
nand U7277 (N_7277,N_7050,N_7107);
nor U7278 (N_7278,N_7130,N_7144);
nor U7279 (N_7279,N_7067,N_7049);
xor U7280 (N_7280,N_7115,N_7041);
nand U7281 (N_7281,N_7117,N_7136);
nand U7282 (N_7282,N_7160,N_7134);
and U7283 (N_7283,N_7188,N_7168);
and U7284 (N_7284,N_7190,N_7135);
or U7285 (N_7285,N_7056,N_7218);
xnor U7286 (N_7286,N_7116,N_7121);
and U7287 (N_7287,N_7112,N_7140);
and U7288 (N_7288,N_7129,N_7114);
nand U7289 (N_7289,N_7087,N_7045);
xnor U7290 (N_7290,N_7109,N_7146);
and U7291 (N_7291,N_7075,N_7161);
or U7292 (N_7292,N_7009,N_7060);
xor U7293 (N_7293,N_7030,N_7052);
nand U7294 (N_7294,N_7015,N_7230);
nor U7295 (N_7295,N_7238,N_7197);
nand U7296 (N_7296,N_7203,N_7032);
and U7297 (N_7297,N_7148,N_7110);
or U7298 (N_7298,N_7155,N_7089);
xnor U7299 (N_7299,N_7182,N_7120);
nor U7300 (N_7300,N_7071,N_7178);
and U7301 (N_7301,N_7085,N_7132);
nand U7302 (N_7302,N_7074,N_7046);
or U7303 (N_7303,N_7051,N_7036);
xor U7304 (N_7304,N_7228,N_7022);
and U7305 (N_7305,N_7124,N_7137);
nand U7306 (N_7306,N_7200,N_7076);
nand U7307 (N_7307,N_7092,N_7042);
or U7308 (N_7308,N_7008,N_7010);
xnor U7309 (N_7309,N_7245,N_7111);
and U7310 (N_7310,N_7081,N_7196);
and U7311 (N_7311,N_7012,N_7005);
xor U7312 (N_7312,N_7159,N_7035);
xnor U7313 (N_7313,N_7079,N_7225);
nand U7314 (N_7314,N_7099,N_7183);
nor U7315 (N_7315,N_7240,N_7098);
and U7316 (N_7316,N_7167,N_7176);
nor U7317 (N_7317,N_7063,N_7207);
or U7318 (N_7318,N_7103,N_7088);
nor U7319 (N_7319,N_7033,N_7173);
nand U7320 (N_7320,N_7097,N_7222);
nand U7321 (N_7321,N_7142,N_7249);
nor U7322 (N_7322,N_7086,N_7083);
xnor U7323 (N_7323,N_7062,N_7210);
xor U7324 (N_7324,N_7091,N_7028);
nand U7325 (N_7325,N_7165,N_7195);
or U7326 (N_7326,N_7152,N_7118);
xor U7327 (N_7327,N_7239,N_7246);
nor U7328 (N_7328,N_7095,N_7043);
nor U7329 (N_7329,N_7247,N_7007);
xnor U7330 (N_7330,N_7201,N_7224);
or U7331 (N_7331,N_7164,N_7053);
nand U7332 (N_7332,N_7127,N_7038);
nor U7333 (N_7333,N_7184,N_7221);
nand U7334 (N_7334,N_7054,N_7226);
nor U7335 (N_7335,N_7189,N_7094);
or U7336 (N_7336,N_7232,N_7002);
and U7337 (N_7337,N_7145,N_7082);
nand U7338 (N_7338,N_7205,N_7234);
nor U7339 (N_7339,N_7047,N_7181);
nand U7340 (N_7340,N_7211,N_7235);
xor U7341 (N_7341,N_7003,N_7215);
or U7342 (N_7342,N_7169,N_7179);
or U7343 (N_7343,N_7202,N_7068);
or U7344 (N_7344,N_7172,N_7044);
or U7345 (N_7345,N_7147,N_7223);
or U7346 (N_7346,N_7151,N_7141);
nor U7347 (N_7347,N_7143,N_7126);
xnor U7348 (N_7348,N_7149,N_7093);
xor U7349 (N_7349,N_7013,N_7192);
nor U7350 (N_7350,N_7080,N_7020);
or U7351 (N_7351,N_7069,N_7191);
and U7352 (N_7352,N_7014,N_7104);
xnor U7353 (N_7353,N_7057,N_7024);
or U7354 (N_7354,N_7244,N_7108);
xor U7355 (N_7355,N_7180,N_7128);
and U7356 (N_7356,N_7139,N_7236);
or U7357 (N_7357,N_7204,N_7004);
or U7358 (N_7358,N_7105,N_7163);
nand U7359 (N_7359,N_7019,N_7185);
and U7360 (N_7360,N_7025,N_7220);
nand U7361 (N_7361,N_7154,N_7000);
and U7362 (N_7362,N_7153,N_7248);
xnor U7363 (N_7363,N_7006,N_7106);
or U7364 (N_7364,N_7171,N_7199);
or U7365 (N_7365,N_7001,N_7090);
nand U7366 (N_7366,N_7193,N_7123);
xnor U7367 (N_7367,N_7237,N_7131);
xor U7368 (N_7368,N_7209,N_7157);
nor U7369 (N_7369,N_7040,N_7150);
nand U7370 (N_7370,N_7214,N_7138);
nand U7371 (N_7371,N_7177,N_7064);
or U7372 (N_7372,N_7156,N_7175);
or U7373 (N_7373,N_7219,N_7048);
or U7374 (N_7374,N_7102,N_7227);
and U7375 (N_7375,N_7246,N_7144);
nand U7376 (N_7376,N_7225,N_7165);
or U7377 (N_7377,N_7017,N_7108);
or U7378 (N_7378,N_7225,N_7128);
nor U7379 (N_7379,N_7207,N_7121);
xnor U7380 (N_7380,N_7198,N_7168);
nor U7381 (N_7381,N_7204,N_7146);
nand U7382 (N_7382,N_7207,N_7150);
nor U7383 (N_7383,N_7135,N_7151);
nand U7384 (N_7384,N_7098,N_7045);
or U7385 (N_7385,N_7023,N_7077);
and U7386 (N_7386,N_7064,N_7203);
and U7387 (N_7387,N_7012,N_7032);
nand U7388 (N_7388,N_7095,N_7081);
nor U7389 (N_7389,N_7063,N_7043);
and U7390 (N_7390,N_7160,N_7111);
and U7391 (N_7391,N_7167,N_7070);
nor U7392 (N_7392,N_7202,N_7101);
or U7393 (N_7393,N_7046,N_7037);
or U7394 (N_7394,N_7246,N_7121);
nor U7395 (N_7395,N_7237,N_7029);
nor U7396 (N_7396,N_7208,N_7146);
xnor U7397 (N_7397,N_7222,N_7016);
nor U7398 (N_7398,N_7058,N_7148);
nand U7399 (N_7399,N_7034,N_7065);
nand U7400 (N_7400,N_7195,N_7090);
nand U7401 (N_7401,N_7070,N_7007);
and U7402 (N_7402,N_7179,N_7233);
and U7403 (N_7403,N_7140,N_7111);
and U7404 (N_7404,N_7008,N_7221);
and U7405 (N_7405,N_7048,N_7083);
nor U7406 (N_7406,N_7191,N_7217);
nor U7407 (N_7407,N_7032,N_7149);
and U7408 (N_7408,N_7087,N_7225);
xnor U7409 (N_7409,N_7230,N_7073);
nand U7410 (N_7410,N_7136,N_7113);
nand U7411 (N_7411,N_7171,N_7008);
and U7412 (N_7412,N_7036,N_7073);
nor U7413 (N_7413,N_7243,N_7238);
nand U7414 (N_7414,N_7047,N_7186);
xnor U7415 (N_7415,N_7063,N_7219);
nand U7416 (N_7416,N_7146,N_7107);
nand U7417 (N_7417,N_7176,N_7227);
nor U7418 (N_7418,N_7057,N_7134);
nand U7419 (N_7419,N_7232,N_7059);
or U7420 (N_7420,N_7131,N_7116);
nor U7421 (N_7421,N_7014,N_7230);
nand U7422 (N_7422,N_7085,N_7177);
and U7423 (N_7423,N_7086,N_7160);
and U7424 (N_7424,N_7216,N_7238);
or U7425 (N_7425,N_7032,N_7207);
and U7426 (N_7426,N_7108,N_7239);
nand U7427 (N_7427,N_7108,N_7133);
or U7428 (N_7428,N_7135,N_7178);
and U7429 (N_7429,N_7230,N_7086);
xnor U7430 (N_7430,N_7139,N_7171);
nor U7431 (N_7431,N_7242,N_7109);
xor U7432 (N_7432,N_7185,N_7174);
nor U7433 (N_7433,N_7083,N_7204);
xnor U7434 (N_7434,N_7192,N_7042);
xor U7435 (N_7435,N_7076,N_7248);
and U7436 (N_7436,N_7061,N_7077);
nor U7437 (N_7437,N_7130,N_7105);
or U7438 (N_7438,N_7037,N_7143);
or U7439 (N_7439,N_7167,N_7243);
and U7440 (N_7440,N_7159,N_7172);
xor U7441 (N_7441,N_7005,N_7185);
xor U7442 (N_7442,N_7172,N_7204);
or U7443 (N_7443,N_7059,N_7014);
or U7444 (N_7444,N_7007,N_7234);
or U7445 (N_7445,N_7106,N_7120);
or U7446 (N_7446,N_7128,N_7091);
xnor U7447 (N_7447,N_7064,N_7048);
xnor U7448 (N_7448,N_7109,N_7047);
nor U7449 (N_7449,N_7167,N_7153);
nor U7450 (N_7450,N_7174,N_7184);
nor U7451 (N_7451,N_7061,N_7228);
nor U7452 (N_7452,N_7040,N_7211);
or U7453 (N_7453,N_7024,N_7228);
or U7454 (N_7454,N_7048,N_7046);
xnor U7455 (N_7455,N_7099,N_7176);
nand U7456 (N_7456,N_7095,N_7231);
xor U7457 (N_7457,N_7178,N_7052);
nor U7458 (N_7458,N_7103,N_7169);
nor U7459 (N_7459,N_7243,N_7069);
xor U7460 (N_7460,N_7037,N_7242);
nor U7461 (N_7461,N_7088,N_7038);
or U7462 (N_7462,N_7202,N_7188);
nand U7463 (N_7463,N_7135,N_7171);
nand U7464 (N_7464,N_7194,N_7084);
nor U7465 (N_7465,N_7206,N_7084);
nor U7466 (N_7466,N_7215,N_7026);
nand U7467 (N_7467,N_7210,N_7006);
nand U7468 (N_7468,N_7235,N_7010);
and U7469 (N_7469,N_7010,N_7203);
or U7470 (N_7470,N_7040,N_7006);
nand U7471 (N_7471,N_7031,N_7045);
and U7472 (N_7472,N_7161,N_7100);
and U7473 (N_7473,N_7028,N_7093);
and U7474 (N_7474,N_7241,N_7150);
nor U7475 (N_7475,N_7041,N_7197);
nor U7476 (N_7476,N_7016,N_7042);
or U7477 (N_7477,N_7157,N_7183);
or U7478 (N_7478,N_7178,N_7068);
or U7479 (N_7479,N_7109,N_7007);
nor U7480 (N_7480,N_7135,N_7207);
nand U7481 (N_7481,N_7124,N_7246);
and U7482 (N_7482,N_7076,N_7134);
nor U7483 (N_7483,N_7158,N_7064);
and U7484 (N_7484,N_7159,N_7185);
nor U7485 (N_7485,N_7128,N_7085);
nor U7486 (N_7486,N_7113,N_7141);
nand U7487 (N_7487,N_7189,N_7155);
or U7488 (N_7488,N_7177,N_7073);
nand U7489 (N_7489,N_7087,N_7122);
nand U7490 (N_7490,N_7074,N_7070);
nor U7491 (N_7491,N_7132,N_7056);
nor U7492 (N_7492,N_7119,N_7161);
or U7493 (N_7493,N_7028,N_7224);
nand U7494 (N_7494,N_7122,N_7232);
and U7495 (N_7495,N_7059,N_7096);
or U7496 (N_7496,N_7101,N_7195);
and U7497 (N_7497,N_7081,N_7093);
and U7498 (N_7498,N_7195,N_7021);
nor U7499 (N_7499,N_7238,N_7160);
nand U7500 (N_7500,N_7373,N_7432);
or U7501 (N_7501,N_7485,N_7317);
nor U7502 (N_7502,N_7271,N_7437);
nand U7503 (N_7503,N_7475,N_7496);
nor U7504 (N_7504,N_7285,N_7277);
nand U7505 (N_7505,N_7387,N_7328);
and U7506 (N_7506,N_7431,N_7260);
or U7507 (N_7507,N_7411,N_7428);
and U7508 (N_7508,N_7350,N_7310);
nand U7509 (N_7509,N_7474,N_7423);
and U7510 (N_7510,N_7446,N_7283);
nand U7511 (N_7511,N_7424,N_7326);
nand U7512 (N_7512,N_7347,N_7440);
xnor U7513 (N_7513,N_7395,N_7419);
and U7514 (N_7514,N_7416,N_7267);
nor U7515 (N_7515,N_7262,N_7315);
or U7516 (N_7516,N_7459,N_7489);
nor U7517 (N_7517,N_7257,N_7451);
xnor U7518 (N_7518,N_7327,N_7417);
xor U7519 (N_7519,N_7392,N_7410);
xnor U7520 (N_7520,N_7358,N_7284);
or U7521 (N_7521,N_7287,N_7320);
nor U7522 (N_7522,N_7425,N_7385);
and U7523 (N_7523,N_7409,N_7281);
nor U7524 (N_7524,N_7445,N_7407);
nand U7525 (N_7525,N_7361,N_7458);
nor U7526 (N_7526,N_7273,N_7453);
and U7527 (N_7527,N_7369,N_7316);
nand U7528 (N_7528,N_7389,N_7405);
nand U7529 (N_7529,N_7280,N_7335);
nand U7530 (N_7530,N_7343,N_7483);
xnor U7531 (N_7531,N_7379,N_7270);
nand U7532 (N_7532,N_7377,N_7415);
or U7533 (N_7533,N_7430,N_7336);
nor U7534 (N_7534,N_7418,N_7408);
nor U7535 (N_7535,N_7490,N_7339);
or U7536 (N_7536,N_7355,N_7472);
nor U7537 (N_7537,N_7384,N_7290);
and U7538 (N_7538,N_7365,N_7497);
nor U7539 (N_7539,N_7380,N_7396);
or U7540 (N_7540,N_7482,N_7499);
and U7541 (N_7541,N_7442,N_7289);
and U7542 (N_7542,N_7253,N_7266);
xor U7543 (N_7543,N_7341,N_7264);
and U7544 (N_7544,N_7414,N_7330);
nand U7545 (N_7545,N_7397,N_7332);
xor U7546 (N_7546,N_7466,N_7311);
or U7547 (N_7547,N_7307,N_7299);
xnor U7548 (N_7548,N_7366,N_7457);
nand U7549 (N_7549,N_7353,N_7469);
and U7550 (N_7550,N_7337,N_7346);
and U7551 (N_7551,N_7374,N_7439);
nand U7552 (N_7552,N_7376,N_7463);
and U7553 (N_7553,N_7433,N_7404);
or U7554 (N_7554,N_7268,N_7256);
nor U7555 (N_7555,N_7441,N_7252);
and U7556 (N_7556,N_7406,N_7486);
and U7557 (N_7557,N_7470,N_7494);
nor U7558 (N_7558,N_7449,N_7308);
nor U7559 (N_7559,N_7455,N_7434);
or U7560 (N_7560,N_7293,N_7325);
or U7561 (N_7561,N_7334,N_7388);
nand U7562 (N_7562,N_7381,N_7322);
or U7563 (N_7563,N_7342,N_7471);
nor U7564 (N_7564,N_7261,N_7464);
nand U7565 (N_7565,N_7391,N_7421);
xnor U7566 (N_7566,N_7359,N_7420);
and U7567 (N_7567,N_7398,N_7286);
xor U7568 (N_7568,N_7498,N_7321);
xnor U7569 (N_7569,N_7495,N_7371);
nand U7570 (N_7570,N_7324,N_7447);
nor U7571 (N_7571,N_7477,N_7300);
nor U7572 (N_7572,N_7468,N_7305);
or U7573 (N_7573,N_7360,N_7402);
xnor U7574 (N_7574,N_7295,N_7333);
or U7575 (N_7575,N_7390,N_7329);
and U7576 (N_7576,N_7383,N_7488);
and U7577 (N_7577,N_7427,N_7296);
nand U7578 (N_7578,N_7476,N_7484);
xnor U7579 (N_7579,N_7251,N_7375);
nor U7580 (N_7580,N_7399,N_7344);
nor U7581 (N_7581,N_7259,N_7368);
and U7582 (N_7582,N_7288,N_7378);
nand U7583 (N_7583,N_7255,N_7479);
or U7584 (N_7584,N_7370,N_7318);
xnor U7585 (N_7585,N_7429,N_7302);
and U7586 (N_7586,N_7276,N_7436);
or U7587 (N_7587,N_7362,N_7291);
and U7588 (N_7588,N_7491,N_7400);
nand U7589 (N_7589,N_7356,N_7292);
nand U7590 (N_7590,N_7403,N_7493);
nor U7591 (N_7591,N_7275,N_7367);
and U7592 (N_7592,N_7443,N_7372);
nor U7593 (N_7593,N_7274,N_7345);
xor U7594 (N_7594,N_7279,N_7487);
nor U7595 (N_7595,N_7386,N_7444);
xor U7596 (N_7596,N_7461,N_7454);
nor U7597 (N_7597,N_7269,N_7467);
xnor U7598 (N_7598,N_7462,N_7323);
nor U7599 (N_7599,N_7309,N_7422);
or U7600 (N_7600,N_7278,N_7357);
and U7601 (N_7601,N_7478,N_7393);
nand U7602 (N_7602,N_7412,N_7456);
nor U7603 (N_7603,N_7382,N_7331);
and U7604 (N_7604,N_7450,N_7435);
nand U7605 (N_7605,N_7340,N_7413);
xor U7606 (N_7606,N_7314,N_7351);
xor U7607 (N_7607,N_7250,N_7401);
or U7608 (N_7608,N_7254,N_7263);
xnor U7609 (N_7609,N_7304,N_7473);
or U7610 (N_7610,N_7282,N_7352);
and U7611 (N_7611,N_7448,N_7306);
and U7612 (N_7612,N_7294,N_7426);
and U7613 (N_7613,N_7348,N_7258);
xor U7614 (N_7614,N_7272,N_7481);
nand U7615 (N_7615,N_7354,N_7364);
and U7616 (N_7616,N_7394,N_7363);
nor U7617 (N_7617,N_7349,N_7312);
nand U7618 (N_7618,N_7303,N_7265);
nor U7619 (N_7619,N_7465,N_7338);
nor U7620 (N_7620,N_7297,N_7298);
nand U7621 (N_7621,N_7319,N_7452);
or U7622 (N_7622,N_7438,N_7480);
and U7623 (N_7623,N_7313,N_7301);
xnor U7624 (N_7624,N_7460,N_7492);
nor U7625 (N_7625,N_7350,N_7464);
nand U7626 (N_7626,N_7360,N_7391);
nor U7627 (N_7627,N_7418,N_7250);
and U7628 (N_7628,N_7414,N_7456);
or U7629 (N_7629,N_7295,N_7391);
xor U7630 (N_7630,N_7364,N_7376);
or U7631 (N_7631,N_7392,N_7332);
nor U7632 (N_7632,N_7424,N_7383);
nand U7633 (N_7633,N_7291,N_7420);
nor U7634 (N_7634,N_7457,N_7396);
xor U7635 (N_7635,N_7394,N_7386);
or U7636 (N_7636,N_7320,N_7351);
xnor U7637 (N_7637,N_7476,N_7424);
xor U7638 (N_7638,N_7470,N_7371);
xnor U7639 (N_7639,N_7371,N_7390);
xnor U7640 (N_7640,N_7335,N_7295);
or U7641 (N_7641,N_7465,N_7420);
nand U7642 (N_7642,N_7490,N_7282);
or U7643 (N_7643,N_7251,N_7380);
xor U7644 (N_7644,N_7417,N_7351);
xnor U7645 (N_7645,N_7412,N_7403);
or U7646 (N_7646,N_7469,N_7267);
or U7647 (N_7647,N_7311,N_7387);
nor U7648 (N_7648,N_7289,N_7339);
or U7649 (N_7649,N_7479,N_7397);
or U7650 (N_7650,N_7424,N_7282);
and U7651 (N_7651,N_7299,N_7266);
or U7652 (N_7652,N_7301,N_7464);
xor U7653 (N_7653,N_7487,N_7330);
nor U7654 (N_7654,N_7498,N_7312);
and U7655 (N_7655,N_7443,N_7251);
nor U7656 (N_7656,N_7362,N_7479);
or U7657 (N_7657,N_7417,N_7446);
xnor U7658 (N_7658,N_7341,N_7482);
xor U7659 (N_7659,N_7416,N_7255);
nor U7660 (N_7660,N_7394,N_7426);
nor U7661 (N_7661,N_7258,N_7361);
nor U7662 (N_7662,N_7340,N_7301);
nor U7663 (N_7663,N_7264,N_7343);
and U7664 (N_7664,N_7465,N_7257);
nor U7665 (N_7665,N_7464,N_7348);
or U7666 (N_7666,N_7259,N_7369);
or U7667 (N_7667,N_7415,N_7301);
or U7668 (N_7668,N_7275,N_7422);
xor U7669 (N_7669,N_7395,N_7354);
nand U7670 (N_7670,N_7354,N_7437);
xor U7671 (N_7671,N_7304,N_7480);
nor U7672 (N_7672,N_7459,N_7292);
or U7673 (N_7673,N_7446,N_7269);
or U7674 (N_7674,N_7388,N_7405);
or U7675 (N_7675,N_7417,N_7360);
nand U7676 (N_7676,N_7383,N_7436);
and U7677 (N_7677,N_7276,N_7354);
nor U7678 (N_7678,N_7268,N_7266);
xor U7679 (N_7679,N_7416,N_7397);
nor U7680 (N_7680,N_7407,N_7414);
nand U7681 (N_7681,N_7365,N_7273);
nor U7682 (N_7682,N_7414,N_7265);
xnor U7683 (N_7683,N_7463,N_7427);
xnor U7684 (N_7684,N_7288,N_7336);
nand U7685 (N_7685,N_7465,N_7459);
and U7686 (N_7686,N_7438,N_7366);
nand U7687 (N_7687,N_7252,N_7485);
nor U7688 (N_7688,N_7407,N_7468);
and U7689 (N_7689,N_7444,N_7327);
and U7690 (N_7690,N_7441,N_7396);
xnor U7691 (N_7691,N_7481,N_7365);
and U7692 (N_7692,N_7259,N_7313);
xnor U7693 (N_7693,N_7400,N_7376);
xnor U7694 (N_7694,N_7442,N_7346);
xnor U7695 (N_7695,N_7325,N_7277);
and U7696 (N_7696,N_7459,N_7477);
xnor U7697 (N_7697,N_7282,N_7474);
nand U7698 (N_7698,N_7411,N_7439);
xor U7699 (N_7699,N_7439,N_7310);
nor U7700 (N_7700,N_7460,N_7356);
or U7701 (N_7701,N_7427,N_7451);
nand U7702 (N_7702,N_7302,N_7280);
xnor U7703 (N_7703,N_7370,N_7489);
xnor U7704 (N_7704,N_7468,N_7430);
and U7705 (N_7705,N_7412,N_7427);
nor U7706 (N_7706,N_7326,N_7283);
nand U7707 (N_7707,N_7397,N_7499);
or U7708 (N_7708,N_7374,N_7466);
nand U7709 (N_7709,N_7422,N_7297);
or U7710 (N_7710,N_7315,N_7493);
or U7711 (N_7711,N_7346,N_7340);
or U7712 (N_7712,N_7357,N_7477);
or U7713 (N_7713,N_7417,N_7423);
and U7714 (N_7714,N_7413,N_7287);
nor U7715 (N_7715,N_7288,N_7312);
and U7716 (N_7716,N_7482,N_7471);
nand U7717 (N_7717,N_7399,N_7461);
and U7718 (N_7718,N_7405,N_7339);
or U7719 (N_7719,N_7309,N_7364);
nor U7720 (N_7720,N_7437,N_7359);
and U7721 (N_7721,N_7309,N_7443);
xnor U7722 (N_7722,N_7338,N_7480);
nand U7723 (N_7723,N_7310,N_7427);
and U7724 (N_7724,N_7406,N_7301);
nand U7725 (N_7725,N_7251,N_7397);
nand U7726 (N_7726,N_7274,N_7454);
nand U7727 (N_7727,N_7321,N_7274);
or U7728 (N_7728,N_7353,N_7463);
and U7729 (N_7729,N_7251,N_7485);
xnor U7730 (N_7730,N_7417,N_7253);
xor U7731 (N_7731,N_7454,N_7371);
nor U7732 (N_7732,N_7398,N_7415);
nor U7733 (N_7733,N_7450,N_7418);
xor U7734 (N_7734,N_7395,N_7310);
xor U7735 (N_7735,N_7391,N_7470);
xor U7736 (N_7736,N_7260,N_7466);
nand U7737 (N_7737,N_7423,N_7457);
or U7738 (N_7738,N_7496,N_7398);
or U7739 (N_7739,N_7332,N_7450);
and U7740 (N_7740,N_7265,N_7257);
nor U7741 (N_7741,N_7380,N_7456);
and U7742 (N_7742,N_7426,N_7461);
xnor U7743 (N_7743,N_7255,N_7351);
nor U7744 (N_7744,N_7386,N_7307);
or U7745 (N_7745,N_7284,N_7450);
nor U7746 (N_7746,N_7307,N_7458);
nand U7747 (N_7747,N_7396,N_7285);
nand U7748 (N_7748,N_7482,N_7445);
nor U7749 (N_7749,N_7460,N_7365);
and U7750 (N_7750,N_7552,N_7514);
nand U7751 (N_7751,N_7540,N_7594);
nand U7752 (N_7752,N_7666,N_7685);
nor U7753 (N_7753,N_7523,N_7601);
xnor U7754 (N_7754,N_7574,N_7597);
or U7755 (N_7755,N_7660,N_7647);
xnor U7756 (N_7756,N_7578,N_7687);
xor U7757 (N_7757,N_7588,N_7630);
xor U7758 (N_7758,N_7712,N_7681);
nor U7759 (N_7759,N_7707,N_7701);
and U7760 (N_7760,N_7742,N_7605);
nand U7761 (N_7761,N_7589,N_7662);
nor U7762 (N_7762,N_7583,N_7725);
nand U7763 (N_7763,N_7646,N_7537);
xor U7764 (N_7764,N_7546,N_7746);
xnor U7765 (N_7765,N_7658,N_7694);
nor U7766 (N_7766,N_7555,N_7545);
nand U7767 (N_7767,N_7517,N_7645);
nand U7768 (N_7768,N_7745,N_7604);
or U7769 (N_7769,N_7634,N_7683);
and U7770 (N_7770,N_7679,N_7542);
nand U7771 (N_7771,N_7623,N_7573);
nor U7772 (N_7772,N_7511,N_7611);
nor U7773 (N_7773,N_7561,N_7501);
nor U7774 (N_7774,N_7619,N_7717);
nor U7775 (N_7775,N_7529,N_7600);
or U7776 (N_7776,N_7720,N_7535);
and U7777 (N_7777,N_7741,N_7509);
and U7778 (N_7778,N_7560,N_7699);
or U7779 (N_7779,N_7677,N_7722);
or U7780 (N_7780,N_7569,N_7633);
nand U7781 (N_7781,N_7676,N_7715);
nor U7782 (N_7782,N_7650,N_7591);
nor U7783 (N_7783,N_7515,N_7644);
nand U7784 (N_7784,N_7642,N_7695);
nor U7785 (N_7785,N_7705,N_7626);
xor U7786 (N_7786,N_7627,N_7661);
and U7787 (N_7787,N_7628,N_7549);
or U7788 (N_7788,N_7551,N_7575);
xor U7789 (N_7789,N_7587,N_7708);
xnor U7790 (N_7790,N_7543,N_7553);
nand U7791 (N_7791,N_7706,N_7731);
nor U7792 (N_7792,N_7547,N_7688);
or U7793 (N_7793,N_7632,N_7723);
xnor U7794 (N_7794,N_7516,N_7652);
xor U7795 (N_7795,N_7500,N_7593);
nor U7796 (N_7796,N_7518,N_7590);
or U7797 (N_7797,N_7592,N_7709);
xnor U7798 (N_7798,N_7564,N_7513);
xnor U7799 (N_7799,N_7739,N_7544);
nor U7800 (N_7800,N_7669,N_7654);
nand U7801 (N_7801,N_7572,N_7571);
and U7802 (N_7802,N_7610,N_7530);
nor U7803 (N_7803,N_7638,N_7657);
and U7804 (N_7804,N_7702,N_7556);
nor U7805 (N_7805,N_7686,N_7749);
or U7806 (N_7806,N_7736,N_7651);
nor U7807 (N_7807,N_7629,N_7625);
xor U7808 (N_7808,N_7733,N_7748);
nand U7809 (N_7809,N_7538,N_7693);
nor U7810 (N_7810,N_7643,N_7502);
nor U7811 (N_7811,N_7562,N_7570);
nand U7812 (N_7812,N_7678,N_7698);
xor U7813 (N_7813,N_7747,N_7729);
nand U7814 (N_7814,N_7621,N_7528);
xnor U7815 (N_7815,N_7531,N_7711);
xor U7816 (N_7816,N_7503,N_7690);
xnor U7817 (N_7817,N_7636,N_7639);
or U7818 (N_7818,N_7635,N_7691);
and U7819 (N_7819,N_7567,N_7704);
nor U7820 (N_7820,N_7668,N_7671);
and U7821 (N_7821,N_7697,N_7684);
nor U7822 (N_7822,N_7525,N_7527);
nand U7823 (N_7823,N_7738,N_7582);
or U7824 (N_7824,N_7504,N_7519);
nand U7825 (N_7825,N_7512,N_7724);
and U7826 (N_7826,N_7655,N_7648);
xnor U7827 (N_7827,N_7732,N_7599);
or U7828 (N_7828,N_7550,N_7656);
and U7829 (N_7829,N_7670,N_7584);
or U7830 (N_7830,N_7674,N_7539);
nand U7831 (N_7831,N_7737,N_7609);
xnor U7832 (N_7832,N_7653,N_7734);
or U7833 (N_7833,N_7521,N_7579);
nand U7834 (N_7834,N_7682,N_7603);
nand U7835 (N_7835,N_7596,N_7522);
and U7836 (N_7836,N_7728,N_7719);
xor U7837 (N_7837,N_7641,N_7718);
nand U7838 (N_7838,N_7507,N_7526);
nand U7839 (N_7839,N_7602,N_7508);
xnor U7840 (N_7840,N_7563,N_7580);
and U7841 (N_7841,N_7700,N_7505);
or U7842 (N_7842,N_7689,N_7620);
and U7843 (N_7843,N_7536,N_7692);
nor U7844 (N_7844,N_7640,N_7606);
nand U7845 (N_7845,N_7649,N_7675);
xor U7846 (N_7846,N_7532,N_7624);
xnor U7847 (N_7847,N_7506,N_7714);
and U7848 (N_7848,N_7622,N_7617);
and U7849 (N_7849,N_7659,N_7735);
xor U7850 (N_7850,N_7559,N_7557);
nand U7851 (N_7851,N_7585,N_7566);
nor U7852 (N_7852,N_7595,N_7607);
or U7853 (N_7853,N_7730,N_7581);
nor U7854 (N_7854,N_7613,N_7586);
nor U7855 (N_7855,N_7565,N_7713);
nor U7856 (N_7856,N_7664,N_7716);
and U7857 (N_7857,N_7554,N_7703);
nor U7858 (N_7858,N_7637,N_7576);
nor U7859 (N_7859,N_7726,N_7533);
or U7860 (N_7860,N_7696,N_7680);
or U7861 (N_7861,N_7568,N_7667);
and U7862 (N_7862,N_7534,N_7520);
nand U7863 (N_7863,N_7618,N_7541);
and U7864 (N_7864,N_7524,N_7614);
xor U7865 (N_7865,N_7548,N_7577);
nand U7866 (N_7866,N_7612,N_7744);
nor U7867 (N_7867,N_7727,N_7510);
xor U7868 (N_7868,N_7743,N_7740);
xor U7869 (N_7869,N_7598,N_7663);
nor U7870 (N_7870,N_7608,N_7616);
and U7871 (N_7871,N_7721,N_7615);
and U7872 (N_7872,N_7672,N_7673);
xnor U7873 (N_7873,N_7665,N_7631);
xor U7874 (N_7874,N_7558,N_7710);
nand U7875 (N_7875,N_7594,N_7667);
xnor U7876 (N_7876,N_7517,N_7736);
and U7877 (N_7877,N_7503,N_7643);
nand U7878 (N_7878,N_7662,N_7618);
nand U7879 (N_7879,N_7547,N_7574);
and U7880 (N_7880,N_7542,N_7639);
xnor U7881 (N_7881,N_7527,N_7522);
or U7882 (N_7882,N_7656,N_7647);
and U7883 (N_7883,N_7656,N_7739);
nand U7884 (N_7884,N_7556,N_7542);
nor U7885 (N_7885,N_7694,N_7738);
or U7886 (N_7886,N_7721,N_7592);
xnor U7887 (N_7887,N_7710,N_7533);
or U7888 (N_7888,N_7683,N_7741);
or U7889 (N_7889,N_7639,N_7605);
nand U7890 (N_7890,N_7537,N_7671);
nand U7891 (N_7891,N_7678,N_7660);
nor U7892 (N_7892,N_7568,N_7511);
and U7893 (N_7893,N_7677,N_7613);
xnor U7894 (N_7894,N_7708,N_7615);
xor U7895 (N_7895,N_7622,N_7744);
or U7896 (N_7896,N_7668,N_7662);
nand U7897 (N_7897,N_7569,N_7714);
xor U7898 (N_7898,N_7609,N_7548);
xnor U7899 (N_7899,N_7697,N_7681);
or U7900 (N_7900,N_7628,N_7531);
or U7901 (N_7901,N_7507,N_7741);
xor U7902 (N_7902,N_7645,N_7506);
or U7903 (N_7903,N_7705,N_7704);
or U7904 (N_7904,N_7576,N_7592);
nor U7905 (N_7905,N_7625,N_7607);
xor U7906 (N_7906,N_7710,N_7501);
and U7907 (N_7907,N_7697,N_7587);
or U7908 (N_7908,N_7693,N_7584);
or U7909 (N_7909,N_7719,N_7532);
or U7910 (N_7910,N_7568,N_7529);
nand U7911 (N_7911,N_7656,N_7540);
nor U7912 (N_7912,N_7651,N_7503);
xor U7913 (N_7913,N_7681,N_7608);
xor U7914 (N_7914,N_7740,N_7613);
and U7915 (N_7915,N_7697,N_7621);
or U7916 (N_7916,N_7699,N_7710);
and U7917 (N_7917,N_7739,N_7686);
or U7918 (N_7918,N_7749,N_7595);
xor U7919 (N_7919,N_7657,N_7738);
and U7920 (N_7920,N_7605,N_7665);
and U7921 (N_7921,N_7577,N_7638);
xnor U7922 (N_7922,N_7533,N_7667);
xnor U7923 (N_7923,N_7679,N_7716);
nor U7924 (N_7924,N_7602,N_7570);
nor U7925 (N_7925,N_7643,N_7682);
xnor U7926 (N_7926,N_7660,N_7595);
xor U7927 (N_7927,N_7544,N_7741);
nand U7928 (N_7928,N_7658,N_7741);
or U7929 (N_7929,N_7627,N_7616);
or U7930 (N_7930,N_7682,N_7515);
nand U7931 (N_7931,N_7636,N_7744);
nor U7932 (N_7932,N_7691,N_7670);
nand U7933 (N_7933,N_7525,N_7507);
nor U7934 (N_7934,N_7573,N_7642);
nand U7935 (N_7935,N_7552,N_7693);
xor U7936 (N_7936,N_7539,N_7685);
and U7937 (N_7937,N_7569,N_7543);
xor U7938 (N_7938,N_7710,N_7559);
nand U7939 (N_7939,N_7721,N_7535);
and U7940 (N_7940,N_7523,N_7729);
and U7941 (N_7941,N_7746,N_7607);
or U7942 (N_7942,N_7639,N_7693);
or U7943 (N_7943,N_7651,N_7712);
or U7944 (N_7944,N_7645,N_7569);
and U7945 (N_7945,N_7745,N_7664);
nor U7946 (N_7946,N_7696,N_7665);
or U7947 (N_7947,N_7596,N_7681);
xnor U7948 (N_7948,N_7567,N_7691);
nand U7949 (N_7949,N_7587,N_7622);
nand U7950 (N_7950,N_7662,N_7583);
xor U7951 (N_7951,N_7640,N_7660);
nand U7952 (N_7952,N_7654,N_7550);
nor U7953 (N_7953,N_7591,N_7690);
nand U7954 (N_7954,N_7586,N_7592);
or U7955 (N_7955,N_7735,N_7715);
and U7956 (N_7956,N_7541,N_7548);
or U7957 (N_7957,N_7500,N_7566);
nor U7958 (N_7958,N_7625,N_7544);
nor U7959 (N_7959,N_7684,N_7578);
and U7960 (N_7960,N_7704,N_7677);
nor U7961 (N_7961,N_7723,N_7519);
or U7962 (N_7962,N_7512,N_7639);
nand U7963 (N_7963,N_7623,N_7613);
xnor U7964 (N_7964,N_7509,N_7594);
xnor U7965 (N_7965,N_7580,N_7711);
nand U7966 (N_7966,N_7582,N_7553);
and U7967 (N_7967,N_7682,N_7628);
or U7968 (N_7968,N_7727,N_7611);
nor U7969 (N_7969,N_7612,N_7645);
nor U7970 (N_7970,N_7630,N_7685);
nand U7971 (N_7971,N_7551,N_7635);
xnor U7972 (N_7972,N_7745,N_7658);
nand U7973 (N_7973,N_7683,N_7509);
xor U7974 (N_7974,N_7567,N_7666);
or U7975 (N_7975,N_7517,N_7592);
xor U7976 (N_7976,N_7623,N_7690);
and U7977 (N_7977,N_7521,N_7604);
or U7978 (N_7978,N_7652,N_7691);
nor U7979 (N_7979,N_7551,N_7618);
or U7980 (N_7980,N_7749,N_7667);
xor U7981 (N_7981,N_7540,N_7639);
and U7982 (N_7982,N_7536,N_7678);
and U7983 (N_7983,N_7706,N_7691);
nor U7984 (N_7984,N_7536,N_7673);
nor U7985 (N_7985,N_7529,N_7582);
nor U7986 (N_7986,N_7731,N_7745);
and U7987 (N_7987,N_7544,N_7650);
or U7988 (N_7988,N_7603,N_7669);
nor U7989 (N_7989,N_7715,N_7600);
nand U7990 (N_7990,N_7736,N_7639);
nand U7991 (N_7991,N_7589,N_7632);
nor U7992 (N_7992,N_7583,N_7726);
nand U7993 (N_7993,N_7572,N_7629);
xor U7994 (N_7994,N_7509,N_7615);
nand U7995 (N_7995,N_7533,N_7747);
xnor U7996 (N_7996,N_7530,N_7508);
nor U7997 (N_7997,N_7720,N_7737);
nor U7998 (N_7998,N_7646,N_7507);
nand U7999 (N_7999,N_7608,N_7584);
and U8000 (N_8000,N_7933,N_7945);
xor U8001 (N_8001,N_7861,N_7938);
and U8002 (N_8002,N_7809,N_7999);
nand U8003 (N_8003,N_7786,N_7842);
xor U8004 (N_8004,N_7814,N_7890);
xnor U8005 (N_8005,N_7979,N_7867);
or U8006 (N_8006,N_7960,N_7758);
or U8007 (N_8007,N_7771,N_7953);
xor U8008 (N_8008,N_7971,N_7828);
xor U8009 (N_8009,N_7893,N_7839);
nor U8010 (N_8010,N_7838,N_7898);
or U8011 (N_8011,N_7783,N_7928);
nand U8012 (N_8012,N_7860,N_7954);
nor U8013 (N_8013,N_7991,N_7874);
or U8014 (N_8014,N_7869,N_7910);
nand U8015 (N_8015,N_7832,N_7961);
xnor U8016 (N_8016,N_7858,N_7949);
nor U8017 (N_8017,N_7926,N_7957);
nor U8018 (N_8018,N_7816,N_7851);
nand U8019 (N_8019,N_7752,N_7792);
xnor U8020 (N_8020,N_7947,N_7856);
xor U8021 (N_8021,N_7889,N_7985);
and U8022 (N_8022,N_7925,N_7956);
or U8023 (N_8023,N_7941,N_7766);
nand U8024 (N_8024,N_7849,N_7976);
nand U8025 (N_8025,N_7875,N_7944);
and U8026 (N_8026,N_7914,N_7996);
and U8027 (N_8027,N_7797,N_7895);
nand U8028 (N_8028,N_7845,N_7772);
or U8029 (N_8029,N_7800,N_7930);
or U8030 (N_8030,N_7884,N_7959);
xnor U8031 (N_8031,N_7826,N_7769);
or U8032 (N_8032,N_7862,N_7866);
or U8033 (N_8033,N_7810,N_7970);
nand U8034 (N_8034,N_7919,N_7847);
or U8035 (N_8035,N_7878,N_7812);
and U8036 (N_8036,N_7865,N_7894);
xor U8037 (N_8037,N_7972,N_7750);
nor U8038 (N_8038,N_7940,N_7964);
and U8039 (N_8039,N_7929,N_7921);
or U8040 (N_8040,N_7932,N_7904);
or U8041 (N_8041,N_7844,N_7891);
nor U8042 (N_8042,N_7807,N_7936);
or U8043 (N_8043,N_7831,N_7794);
nor U8044 (N_8044,N_7883,N_7984);
xnor U8045 (N_8045,N_7859,N_7871);
nand U8046 (N_8046,N_7784,N_7753);
and U8047 (N_8047,N_7983,N_7882);
xor U8048 (N_8048,N_7791,N_7974);
nand U8049 (N_8049,N_7751,N_7775);
or U8050 (N_8050,N_7823,N_7967);
and U8051 (N_8051,N_7853,N_7975);
nand U8052 (N_8052,N_7924,N_7789);
and U8053 (N_8053,N_7958,N_7969);
xor U8054 (N_8054,N_7988,N_7808);
nand U8055 (N_8055,N_7760,N_7824);
and U8056 (N_8056,N_7913,N_7879);
or U8057 (N_8057,N_7822,N_7880);
or U8058 (N_8058,N_7833,N_7781);
nor U8059 (N_8059,N_7780,N_7804);
nand U8060 (N_8060,N_7905,N_7778);
nor U8061 (N_8061,N_7992,N_7835);
nand U8062 (N_8062,N_7907,N_7903);
nand U8063 (N_8063,N_7952,N_7908);
nor U8064 (N_8064,N_7801,N_7899);
xnor U8065 (N_8065,N_7798,N_7968);
nand U8066 (N_8066,N_7790,N_7888);
xnor U8067 (N_8067,N_7872,N_7868);
and U8068 (N_8068,N_7916,N_7840);
nor U8069 (N_8069,N_7762,N_7955);
nand U8070 (N_8070,N_7942,N_7962);
nand U8071 (N_8071,N_7793,N_7855);
nor U8072 (N_8072,N_7806,N_7788);
nor U8073 (N_8073,N_7857,N_7843);
nor U8074 (N_8074,N_7764,N_7963);
and U8075 (N_8075,N_7796,N_7900);
xor U8076 (N_8076,N_7761,N_7795);
and U8077 (N_8077,N_7852,N_7821);
nand U8078 (N_8078,N_7773,N_7965);
or U8079 (N_8079,N_7763,N_7837);
xor U8080 (N_8080,N_7931,N_7981);
and U8081 (N_8081,N_7811,N_7876);
nand U8082 (N_8082,N_7922,N_7864);
or U8083 (N_8083,N_7841,N_7966);
nand U8084 (N_8084,N_7887,N_7848);
and U8085 (N_8085,N_7825,N_7918);
or U8086 (N_8086,N_7896,N_7820);
or U8087 (N_8087,N_7989,N_7998);
and U8088 (N_8088,N_7756,N_7846);
nor U8089 (N_8089,N_7755,N_7920);
and U8090 (N_8090,N_7815,N_7829);
or U8091 (N_8091,N_7906,N_7870);
nor U8092 (N_8092,N_7877,N_7863);
and U8093 (N_8093,N_7767,N_7997);
and U8094 (N_8094,N_7946,N_7782);
nor U8095 (N_8095,N_7834,N_7917);
or U8096 (N_8096,N_7977,N_7776);
nor U8097 (N_8097,N_7927,N_7802);
nor U8098 (N_8098,N_7951,N_7787);
nor U8099 (N_8099,N_7805,N_7911);
and U8100 (N_8100,N_7765,N_7799);
or U8101 (N_8101,N_7915,N_7754);
nand U8102 (N_8102,N_7909,N_7897);
nand U8103 (N_8103,N_7768,N_7779);
and U8104 (N_8104,N_7934,N_7813);
xnor U8105 (N_8105,N_7757,N_7902);
nand U8106 (N_8106,N_7982,N_7912);
and U8107 (N_8107,N_7818,N_7817);
nor U8108 (N_8108,N_7980,N_7987);
xor U8109 (N_8109,N_7836,N_7994);
nand U8110 (N_8110,N_7939,N_7850);
nand U8111 (N_8111,N_7759,N_7892);
nand U8112 (N_8112,N_7948,N_7803);
nor U8113 (N_8113,N_7990,N_7973);
or U8114 (N_8114,N_7854,N_7774);
xor U8115 (N_8115,N_7937,N_7950);
xnor U8116 (N_8116,N_7978,N_7830);
xnor U8117 (N_8117,N_7993,N_7995);
or U8118 (N_8118,N_7785,N_7873);
nor U8119 (N_8119,N_7881,N_7986);
and U8120 (N_8120,N_7935,N_7943);
nor U8121 (N_8121,N_7885,N_7827);
and U8122 (N_8122,N_7901,N_7886);
nand U8123 (N_8123,N_7819,N_7777);
nand U8124 (N_8124,N_7770,N_7923);
or U8125 (N_8125,N_7859,N_7776);
or U8126 (N_8126,N_7936,N_7835);
nor U8127 (N_8127,N_7787,N_7761);
nor U8128 (N_8128,N_7906,N_7919);
or U8129 (N_8129,N_7892,N_7815);
nand U8130 (N_8130,N_7882,N_7779);
nand U8131 (N_8131,N_7904,N_7872);
and U8132 (N_8132,N_7959,N_7764);
xor U8133 (N_8133,N_7766,N_7838);
xor U8134 (N_8134,N_7890,N_7802);
xor U8135 (N_8135,N_7972,N_7852);
nor U8136 (N_8136,N_7946,N_7794);
and U8137 (N_8137,N_7928,N_7912);
nor U8138 (N_8138,N_7854,N_7910);
nor U8139 (N_8139,N_7774,N_7879);
nand U8140 (N_8140,N_7871,N_7953);
nand U8141 (N_8141,N_7861,N_7891);
nand U8142 (N_8142,N_7810,N_7844);
or U8143 (N_8143,N_7790,N_7951);
and U8144 (N_8144,N_7775,N_7893);
or U8145 (N_8145,N_7941,N_7875);
or U8146 (N_8146,N_7872,N_7927);
nor U8147 (N_8147,N_7803,N_7784);
nand U8148 (N_8148,N_7975,N_7828);
xor U8149 (N_8149,N_7978,N_7800);
nand U8150 (N_8150,N_7840,N_7773);
nand U8151 (N_8151,N_7919,N_7956);
nand U8152 (N_8152,N_7931,N_7775);
xnor U8153 (N_8153,N_7909,N_7751);
nor U8154 (N_8154,N_7893,N_7753);
nor U8155 (N_8155,N_7808,N_7804);
xor U8156 (N_8156,N_7900,N_7938);
nor U8157 (N_8157,N_7902,N_7924);
or U8158 (N_8158,N_7896,N_7956);
xnor U8159 (N_8159,N_7967,N_7820);
or U8160 (N_8160,N_7855,N_7854);
and U8161 (N_8161,N_7962,N_7771);
nor U8162 (N_8162,N_7829,N_7856);
nor U8163 (N_8163,N_7928,N_7763);
and U8164 (N_8164,N_7951,N_7777);
nor U8165 (N_8165,N_7972,N_7915);
xnor U8166 (N_8166,N_7941,N_7983);
nor U8167 (N_8167,N_7895,N_7904);
nand U8168 (N_8168,N_7831,N_7891);
and U8169 (N_8169,N_7879,N_7819);
nor U8170 (N_8170,N_7795,N_7837);
or U8171 (N_8171,N_7750,N_7767);
nor U8172 (N_8172,N_7827,N_7840);
nand U8173 (N_8173,N_7866,N_7804);
nor U8174 (N_8174,N_7776,N_7775);
xor U8175 (N_8175,N_7776,N_7935);
nand U8176 (N_8176,N_7904,N_7995);
xor U8177 (N_8177,N_7838,N_7955);
nand U8178 (N_8178,N_7936,N_7868);
nor U8179 (N_8179,N_7885,N_7975);
and U8180 (N_8180,N_7912,N_7966);
nand U8181 (N_8181,N_7995,N_7833);
and U8182 (N_8182,N_7936,N_7922);
and U8183 (N_8183,N_7849,N_7927);
nor U8184 (N_8184,N_7815,N_7789);
nand U8185 (N_8185,N_7916,N_7819);
nand U8186 (N_8186,N_7817,N_7879);
nor U8187 (N_8187,N_7891,N_7906);
and U8188 (N_8188,N_7888,N_7859);
xor U8189 (N_8189,N_7900,N_7760);
or U8190 (N_8190,N_7967,N_7930);
nor U8191 (N_8191,N_7936,N_7826);
xnor U8192 (N_8192,N_7989,N_7943);
xnor U8193 (N_8193,N_7834,N_7929);
nor U8194 (N_8194,N_7794,N_7760);
or U8195 (N_8195,N_7799,N_7801);
xor U8196 (N_8196,N_7970,N_7843);
or U8197 (N_8197,N_7934,N_7883);
nand U8198 (N_8198,N_7935,N_7929);
nand U8199 (N_8199,N_7942,N_7973);
nor U8200 (N_8200,N_7862,N_7846);
or U8201 (N_8201,N_7919,N_7988);
nor U8202 (N_8202,N_7759,N_7938);
or U8203 (N_8203,N_7939,N_7995);
and U8204 (N_8204,N_7893,N_7957);
and U8205 (N_8205,N_7983,N_7944);
xnor U8206 (N_8206,N_7867,N_7804);
nor U8207 (N_8207,N_7904,N_7896);
xnor U8208 (N_8208,N_7880,N_7796);
xnor U8209 (N_8209,N_7820,N_7785);
and U8210 (N_8210,N_7791,N_7852);
and U8211 (N_8211,N_7982,N_7913);
nor U8212 (N_8212,N_7908,N_7903);
or U8213 (N_8213,N_7942,N_7981);
or U8214 (N_8214,N_7875,N_7945);
and U8215 (N_8215,N_7835,N_7996);
and U8216 (N_8216,N_7920,N_7974);
or U8217 (N_8217,N_7933,N_7912);
and U8218 (N_8218,N_7868,N_7808);
nand U8219 (N_8219,N_7959,N_7773);
nor U8220 (N_8220,N_7973,N_7874);
nor U8221 (N_8221,N_7821,N_7917);
nand U8222 (N_8222,N_7827,N_7900);
and U8223 (N_8223,N_7783,N_7987);
nor U8224 (N_8224,N_7758,N_7988);
or U8225 (N_8225,N_7859,N_7842);
nand U8226 (N_8226,N_7976,N_7912);
and U8227 (N_8227,N_7945,N_7952);
and U8228 (N_8228,N_7971,N_7976);
and U8229 (N_8229,N_7755,N_7787);
or U8230 (N_8230,N_7762,N_7973);
or U8231 (N_8231,N_7968,N_7916);
xnor U8232 (N_8232,N_7919,N_7889);
or U8233 (N_8233,N_7999,N_7871);
or U8234 (N_8234,N_7902,N_7955);
nand U8235 (N_8235,N_7982,N_7879);
nor U8236 (N_8236,N_7989,N_7783);
nor U8237 (N_8237,N_7750,N_7944);
nand U8238 (N_8238,N_7886,N_7813);
or U8239 (N_8239,N_7921,N_7922);
nor U8240 (N_8240,N_7969,N_7980);
or U8241 (N_8241,N_7965,N_7945);
nand U8242 (N_8242,N_7774,N_7767);
nor U8243 (N_8243,N_7779,N_7807);
and U8244 (N_8244,N_7882,N_7818);
or U8245 (N_8245,N_7853,N_7916);
or U8246 (N_8246,N_7949,N_7818);
nor U8247 (N_8247,N_7788,N_7877);
nand U8248 (N_8248,N_7835,N_7856);
or U8249 (N_8249,N_7775,N_7985);
or U8250 (N_8250,N_8127,N_8199);
nor U8251 (N_8251,N_8064,N_8108);
nor U8252 (N_8252,N_8090,N_8116);
xor U8253 (N_8253,N_8224,N_8153);
and U8254 (N_8254,N_8117,N_8088);
xnor U8255 (N_8255,N_8119,N_8019);
xor U8256 (N_8256,N_8042,N_8076);
and U8257 (N_8257,N_8248,N_8078);
and U8258 (N_8258,N_8187,N_8202);
xor U8259 (N_8259,N_8073,N_8188);
or U8260 (N_8260,N_8156,N_8138);
nor U8261 (N_8261,N_8045,N_8154);
xor U8262 (N_8262,N_8104,N_8130);
or U8263 (N_8263,N_8174,N_8067);
nor U8264 (N_8264,N_8150,N_8161);
and U8265 (N_8265,N_8216,N_8121);
nor U8266 (N_8266,N_8231,N_8068);
and U8267 (N_8267,N_8179,N_8097);
nor U8268 (N_8268,N_8144,N_8075);
nor U8269 (N_8269,N_8194,N_8024);
nand U8270 (N_8270,N_8186,N_8203);
and U8271 (N_8271,N_8167,N_8109);
xnor U8272 (N_8272,N_8103,N_8239);
nand U8273 (N_8273,N_8141,N_8027);
nor U8274 (N_8274,N_8034,N_8219);
nor U8275 (N_8275,N_8227,N_8062);
and U8276 (N_8276,N_8147,N_8018);
and U8277 (N_8277,N_8053,N_8046);
xnor U8278 (N_8278,N_8201,N_8180);
and U8279 (N_8279,N_8206,N_8099);
nor U8280 (N_8280,N_8001,N_8181);
and U8281 (N_8281,N_8012,N_8168);
nor U8282 (N_8282,N_8157,N_8217);
xnor U8283 (N_8283,N_8094,N_8237);
nand U8284 (N_8284,N_8101,N_8006);
nor U8285 (N_8285,N_8165,N_8115);
nor U8286 (N_8286,N_8079,N_8095);
nor U8287 (N_8287,N_8143,N_8074);
and U8288 (N_8288,N_8210,N_8124);
and U8289 (N_8289,N_8120,N_8133);
nand U8290 (N_8290,N_8085,N_8035);
or U8291 (N_8291,N_8171,N_8063);
and U8292 (N_8292,N_8032,N_8069);
and U8293 (N_8293,N_8198,N_8049);
nor U8294 (N_8294,N_8057,N_8240);
nand U8295 (N_8295,N_8122,N_8055);
and U8296 (N_8296,N_8244,N_8111);
nor U8297 (N_8297,N_8233,N_8234);
nand U8298 (N_8298,N_8070,N_8195);
xnor U8299 (N_8299,N_8232,N_8005);
nor U8300 (N_8300,N_8030,N_8044);
xor U8301 (N_8301,N_8082,N_8148);
or U8302 (N_8302,N_8176,N_8092);
and U8303 (N_8303,N_8016,N_8196);
nand U8304 (N_8304,N_8158,N_8118);
nor U8305 (N_8305,N_8028,N_8169);
and U8306 (N_8306,N_8081,N_8087);
xor U8307 (N_8307,N_8086,N_8205);
nand U8308 (N_8308,N_8007,N_8096);
nor U8309 (N_8309,N_8222,N_8243);
nor U8310 (N_8310,N_8235,N_8223);
or U8311 (N_8311,N_8000,N_8015);
or U8312 (N_8312,N_8043,N_8060);
or U8313 (N_8313,N_8139,N_8066);
or U8314 (N_8314,N_8008,N_8056);
nand U8315 (N_8315,N_8136,N_8159);
nand U8316 (N_8316,N_8191,N_8160);
xnor U8317 (N_8317,N_8149,N_8110);
or U8318 (N_8318,N_8215,N_8221);
nor U8319 (N_8319,N_8129,N_8184);
or U8320 (N_8320,N_8189,N_8170);
nand U8321 (N_8321,N_8151,N_8175);
and U8322 (N_8322,N_8083,N_8051);
nor U8323 (N_8323,N_8236,N_8178);
and U8324 (N_8324,N_8212,N_8023);
xnor U8325 (N_8325,N_8220,N_8214);
or U8326 (N_8326,N_8065,N_8100);
nand U8327 (N_8327,N_8190,N_8113);
nand U8328 (N_8328,N_8052,N_8142);
nand U8329 (N_8329,N_8192,N_8172);
or U8330 (N_8330,N_8197,N_8207);
xnor U8331 (N_8331,N_8166,N_8047);
nand U8332 (N_8332,N_8228,N_8246);
nand U8333 (N_8333,N_8245,N_8020);
xnor U8334 (N_8334,N_8218,N_8013);
nor U8335 (N_8335,N_8021,N_8112);
or U8336 (N_8336,N_8107,N_8004);
and U8337 (N_8337,N_8128,N_8132);
nor U8338 (N_8338,N_8152,N_8054);
nor U8339 (N_8339,N_8230,N_8077);
xor U8340 (N_8340,N_8080,N_8105);
nor U8341 (N_8341,N_8039,N_8238);
xor U8342 (N_8342,N_8071,N_8089);
nand U8343 (N_8343,N_8098,N_8058);
and U8344 (N_8344,N_8226,N_8040);
nand U8345 (N_8345,N_8155,N_8091);
nor U8346 (N_8346,N_8137,N_8010);
or U8347 (N_8347,N_8126,N_8182);
nor U8348 (N_8348,N_8048,N_8106);
nor U8349 (N_8349,N_8037,N_8249);
or U8350 (N_8350,N_8213,N_8185);
or U8351 (N_8351,N_8061,N_8229);
or U8352 (N_8352,N_8183,N_8200);
or U8353 (N_8353,N_8247,N_8022);
nand U8354 (N_8354,N_8036,N_8177);
xnor U8355 (N_8355,N_8026,N_8193);
xnor U8356 (N_8356,N_8163,N_8014);
and U8357 (N_8357,N_8031,N_8084);
or U8358 (N_8358,N_8164,N_8029);
nor U8359 (N_8359,N_8241,N_8131);
nor U8360 (N_8360,N_8009,N_8242);
xnor U8361 (N_8361,N_8072,N_8025);
and U8362 (N_8362,N_8114,N_8003);
nand U8363 (N_8363,N_8209,N_8002);
nand U8364 (N_8364,N_8211,N_8033);
xor U8365 (N_8365,N_8125,N_8134);
nor U8366 (N_8366,N_8204,N_8102);
nand U8367 (N_8367,N_8059,N_8038);
nor U8368 (N_8368,N_8208,N_8093);
and U8369 (N_8369,N_8225,N_8050);
or U8370 (N_8370,N_8041,N_8140);
xor U8371 (N_8371,N_8011,N_8173);
nor U8372 (N_8372,N_8135,N_8123);
and U8373 (N_8373,N_8145,N_8146);
nor U8374 (N_8374,N_8017,N_8162);
or U8375 (N_8375,N_8089,N_8195);
nand U8376 (N_8376,N_8013,N_8221);
xnor U8377 (N_8377,N_8166,N_8084);
xnor U8378 (N_8378,N_8122,N_8039);
xnor U8379 (N_8379,N_8057,N_8204);
or U8380 (N_8380,N_8108,N_8248);
xor U8381 (N_8381,N_8039,N_8218);
nor U8382 (N_8382,N_8174,N_8107);
and U8383 (N_8383,N_8067,N_8224);
or U8384 (N_8384,N_8169,N_8086);
or U8385 (N_8385,N_8074,N_8036);
nand U8386 (N_8386,N_8125,N_8234);
and U8387 (N_8387,N_8104,N_8197);
nand U8388 (N_8388,N_8077,N_8124);
nand U8389 (N_8389,N_8083,N_8038);
nand U8390 (N_8390,N_8203,N_8196);
nand U8391 (N_8391,N_8169,N_8083);
and U8392 (N_8392,N_8234,N_8220);
xnor U8393 (N_8393,N_8061,N_8224);
or U8394 (N_8394,N_8212,N_8169);
and U8395 (N_8395,N_8247,N_8177);
xor U8396 (N_8396,N_8082,N_8053);
and U8397 (N_8397,N_8147,N_8192);
and U8398 (N_8398,N_8115,N_8169);
or U8399 (N_8399,N_8234,N_8059);
xnor U8400 (N_8400,N_8243,N_8117);
and U8401 (N_8401,N_8199,N_8131);
and U8402 (N_8402,N_8190,N_8202);
xnor U8403 (N_8403,N_8159,N_8079);
nand U8404 (N_8404,N_8122,N_8051);
nor U8405 (N_8405,N_8094,N_8080);
or U8406 (N_8406,N_8059,N_8204);
and U8407 (N_8407,N_8223,N_8249);
nand U8408 (N_8408,N_8146,N_8091);
and U8409 (N_8409,N_8141,N_8082);
or U8410 (N_8410,N_8180,N_8053);
and U8411 (N_8411,N_8039,N_8028);
or U8412 (N_8412,N_8149,N_8132);
nor U8413 (N_8413,N_8177,N_8134);
nand U8414 (N_8414,N_8157,N_8012);
or U8415 (N_8415,N_8057,N_8247);
nor U8416 (N_8416,N_8045,N_8095);
xor U8417 (N_8417,N_8095,N_8013);
or U8418 (N_8418,N_8188,N_8208);
and U8419 (N_8419,N_8048,N_8236);
nand U8420 (N_8420,N_8148,N_8064);
nand U8421 (N_8421,N_8212,N_8175);
xor U8422 (N_8422,N_8021,N_8142);
nor U8423 (N_8423,N_8065,N_8142);
or U8424 (N_8424,N_8111,N_8159);
xnor U8425 (N_8425,N_8057,N_8092);
and U8426 (N_8426,N_8182,N_8128);
nand U8427 (N_8427,N_8131,N_8205);
or U8428 (N_8428,N_8145,N_8196);
and U8429 (N_8429,N_8246,N_8140);
nand U8430 (N_8430,N_8033,N_8169);
or U8431 (N_8431,N_8102,N_8239);
or U8432 (N_8432,N_8161,N_8044);
nand U8433 (N_8433,N_8146,N_8063);
nor U8434 (N_8434,N_8228,N_8010);
nand U8435 (N_8435,N_8089,N_8050);
or U8436 (N_8436,N_8012,N_8233);
nand U8437 (N_8437,N_8107,N_8038);
nand U8438 (N_8438,N_8036,N_8208);
or U8439 (N_8439,N_8090,N_8237);
or U8440 (N_8440,N_8124,N_8164);
xor U8441 (N_8441,N_8016,N_8129);
nand U8442 (N_8442,N_8133,N_8160);
nor U8443 (N_8443,N_8201,N_8133);
xor U8444 (N_8444,N_8084,N_8239);
nor U8445 (N_8445,N_8010,N_8123);
or U8446 (N_8446,N_8120,N_8238);
nor U8447 (N_8447,N_8041,N_8076);
or U8448 (N_8448,N_8174,N_8034);
xnor U8449 (N_8449,N_8234,N_8175);
and U8450 (N_8450,N_8053,N_8006);
nor U8451 (N_8451,N_8025,N_8112);
nor U8452 (N_8452,N_8202,N_8230);
xor U8453 (N_8453,N_8245,N_8233);
xor U8454 (N_8454,N_8159,N_8004);
nor U8455 (N_8455,N_8076,N_8108);
nand U8456 (N_8456,N_8060,N_8040);
and U8457 (N_8457,N_8160,N_8012);
nand U8458 (N_8458,N_8160,N_8094);
nand U8459 (N_8459,N_8241,N_8003);
nand U8460 (N_8460,N_8068,N_8085);
and U8461 (N_8461,N_8096,N_8112);
nand U8462 (N_8462,N_8138,N_8134);
nand U8463 (N_8463,N_8165,N_8218);
xnor U8464 (N_8464,N_8083,N_8087);
or U8465 (N_8465,N_8150,N_8111);
nand U8466 (N_8466,N_8026,N_8126);
xnor U8467 (N_8467,N_8075,N_8203);
or U8468 (N_8468,N_8153,N_8060);
nor U8469 (N_8469,N_8170,N_8126);
xnor U8470 (N_8470,N_8246,N_8141);
or U8471 (N_8471,N_8013,N_8155);
and U8472 (N_8472,N_8226,N_8202);
and U8473 (N_8473,N_8218,N_8079);
and U8474 (N_8474,N_8127,N_8217);
nand U8475 (N_8475,N_8103,N_8119);
or U8476 (N_8476,N_8214,N_8063);
and U8477 (N_8477,N_8215,N_8245);
nor U8478 (N_8478,N_8221,N_8151);
nor U8479 (N_8479,N_8184,N_8187);
and U8480 (N_8480,N_8186,N_8126);
or U8481 (N_8481,N_8104,N_8160);
or U8482 (N_8482,N_8127,N_8022);
xor U8483 (N_8483,N_8142,N_8233);
and U8484 (N_8484,N_8022,N_8097);
xnor U8485 (N_8485,N_8039,N_8029);
or U8486 (N_8486,N_8152,N_8134);
and U8487 (N_8487,N_8079,N_8220);
or U8488 (N_8488,N_8019,N_8242);
or U8489 (N_8489,N_8077,N_8088);
or U8490 (N_8490,N_8110,N_8224);
xor U8491 (N_8491,N_8055,N_8036);
xor U8492 (N_8492,N_8164,N_8141);
nor U8493 (N_8493,N_8247,N_8010);
nand U8494 (N_8494,N_8014,N_8153);
or U8495 (N_8495,N_8065,N_8166);
or U8496 (N_8496,N_8202,N_8130);
and U8497 (N_8497,N_8212,N_8077);
nand U8498 (N_8498,N_8211,N_8081);
and U8499 (N_8499,N_8207,N_8172);
nor U8500 (N_8500,N_8494,N_8283);
nor U8501 (N_8501,N_8383,N_8466);
nand U8502 (N_8502,N_8352,N_8322);
or U8503 (N_8503,N_8476,N_8330);
xor U8504 (N_8504,N_8270,N_8405);
xor U8505 (N_8505,N_8473,N_8376);
xnor U8506 (N_8506,N_8347,N_8412);
and U8507 (N_8507,N_8321,N_8271);
xor U8508 (N_8508,N_8419,N_8447);
and U8509 (N_8509,N_8395,N_8257);
nand U8510 (N_8510,N_8492,N_8278);
xnor U8511 (N_8511,N_8478,N_8329);
and U8512 (N_8512,N_8420,N_8438);
xor U8513 (N_8513,N_8470,N_8307);
or U8514 (N_8514,N_8454,N_8315);
nand U8515 (N_8515,N_8264,N_8333);
nand U8516 (N_8516,N_8382,N_8289);
nor U8517 (N_8517,N_8432,N_8305);
nand U8518 (N_8518,N_8430,N_8427);
and U8519 (N_8519,N_8325,N_8442);
and U8520 (N_8520,N_8387,N_8403);
xnor U8521 (N_8521,N_8274,N_8444);
nor U8522 (N_8522,N_8313,N_8407);
and U8523 (N_8523,N_8413,N_8388);
and U8524 (N_8524,N_8471,N_8378);
nand U8525 (N_8525,N_8287,N_8256);
nor U8526 (N_8526,N_8421,N_8269);
nor U8527 (N_8527,N_8469,N_8304);
nor U8528 (N_8528,N_8255,N_8448);
nor U8529 (N_8529,N_8360,N_8439);
xor U8530 (N_8530,N_8346,N_8362);
xnor U8531 (N_8531,N_8331,N_8295);
nor U8532 (N_8532,N_8385,N_8277);
nor U8533 (N_8533,N_8401,N_8349);
xor U8534 (N_8534,N_8497,N_8338);
nand U8535 (N_8535,N_8493,N_8279);
and U8536 (N_8536,N_8417,N_8293);
nor U8537 (N_8537,N_8446,N_8273);
xnor U8538 (N_8538,N_8299,N_8288);
and U8539 (N_8539,N_8353,N_8339);
nand U8540 (N_8540,N_8328,N_8296);
nor U8541 (N_8541,N_8400,N_8272);
and U8542 (N_8542,N_8443,N_8480);
nor U8543 (N_8543,N_8266,N_8397);
nor U8544 (N_8544,N_8286,N_8425);
and U8545 (N_8545,N_8404,N_8357);
nor U8546 (N_8546,N_8457,N_8459);
xor U8547 (N_8547,N_8379,N_8458);
and U8548 (N_8548,N_8391,N_8265);
nand U8549 (N_8549,N_8474,N_8250);
xnor U8550 (N_8550,N_8365,N_8341);
xor U8551 (N_8551,N_8298,N_8259);
or U8552 (N_8552,N_8260,N_8336);
and U8553 (N_8553,N_8472,N_8496);
nand U8554 (N_8554,N_8275,N_8377);
nor U8555 (N_8555,N_8462,N_8491);
or U8556 (N_8556,N_8344,N_8488);
nor U8557 (N_8557,N_8253,N_8441);
nand U8558 (N_8558,N_8453,N_8426);
or U8559 (N_8559,N_8418,N_8334);
or U8560 (N_8560,N_8402,N_8440);
or U8561 (N_8561,N_8369,N_8487);
or U8562 (N_8562,N_8258,N_8316);
xnor U8563 (N_8563,N_8399,N_8381);
nor U8564 (N_8564,N_8414,N_8386);
xnor U8565 (N_8565,N_8319,N_8340);
nor U8566 (N_8566,N_8428,N_8364);
xnor U8567 (N_8567,N_8375,N_8398);
or U8568 (N_8568,N_8300,N_8498);
nor U8569 (N_8569,N_8394,N_8261);
and U8570 (N_8570,N_8485,N_8396);
and U8571 (N_8571,N_8429,N_8436);
xnor U8572 (N_8572,N_8371,N_8358);
and U8573 (N_8573,N_8351,N_8252);
xnor U8574 (N_8574,N_8366,N_8433);
nor U8575 (N_8575,N_8373,N_8354);
xnor U8576 (N_8576,N_8481,N_8372);
nand U8577 (N_8577,N_8356,N_8499);
and U8578 (N_8578,N_8456,N_8348);
xor U8579 (N_8579,N_8370,N_8276);
nand U8580 (N_8580,N_8363,N_8312);
nor U8581 (N_8581,N_8445,N_8464);
and U8582 (N_8582,N_8455,N_8406);
xnor U8583 (N_8583,N_8326,N_8342);
and U8584 (N_8584,N_8380,N_8297);
and U8585 (N_8585,N_8477,N_8318);
and U8586 (N_8586,N_8280,N_8251);
or U8587 (N_8587,N_8311,N_8465);
or U8588 (N_8588,N_8343,N_8282);
nand U8589 (N_8589,N_8415,N_8408);
nand U8590 (N_8590,N_8451,N_8332);
nor U8591 (N_8591,N_8483,N_8324);
and U8592 (N_8592,N_8263,N_8392);
nor U8593 (N_8593,N_8337,N_8450);
or U8594 (N_8594,N_8489,N_8422);
nor U8595 (N_8595,N_8317,N_8320);
or U8596 (N_8596,N_8367,N_8285);
nor U8597 (N_8597,N_8467,N_8490);
or U8598 (N_8598,N_8424,N_8461);
nand U8599 (N_8599,N_8294,N_8292);
and U8600 (N_8600,N_8301,N_8262);
and U8601 (N_8601,N_8460,N_8374);
and U8602 (N_8602,N_8423,N_8479);
nor U8603 (N_8603,N_8361,N_8486);
nor U8604 (N_8604,N_8310,N_8449);
xor U8605 (N_8605,N_8308,N_8350);
or U8606 (N_8606,N_8268,N_8384);
nand U8607 (N_8607,N_8495,N_8345);
or U8608 (N_8608,N_8359,N_8303);
nor U8609 (N_8609,N_8267,N_8431);
and U8610 (N_8610,N_8389,N_8393);
xor U8611 (N_8611,N_8452,N_8409);
nor U8612 (N_8612,N_8355,N_8435);
and U8613 (N_8613,N_8368,N_8434);
nor U8614 (N_8614,N_8390,N_8327);
or U8615 (N_8615,N_8314,N_8410);
xnor U8616 (N_8616,N_8309,N_8290);
or U8617 (N_8617,N_8468,N_8475);
xnor U8618 (N_8618,N_8482,N_8323);
xor U8619 (N_8619,N_8302,N_8254);
or U8620 (N_8620,N_8306,N_8411);
nand U8621 (N_8621,N_8484,N_8284);
nor U8622 (N_8622,N_8335,N_8281);
or U8623 (N_8623,N_8437,N_8416);
nand U8624 (N_8624,N_8291,N_8463);
xnor U8625 (N_8625,N_8369,N_8310);
nor U8626 (N_8626,N_8385,N_8479);
and U8627 (N_8627,N_8365,N_8325);
and U8628 (N_8628,N_8268,N_8417);
nand U8629 (N_8629,N_8253,N_8255);
nand U8630 (N_8630,N_8264,N_8375);
and U8631 (N_8631,N_8462,N_8381);
xnor U8632 (N_8632,N_8301,N_8473);
xor U8633 (N_8633,N_8421,N_8348);
or U8634 (N_8634,N_8258,N_8426);
and U8635 (N_8635,N_8251,N_8263);
xnor U8636 (N_8636,N_8311,N_8398);
xor U8637 (N_8637,N_8429,N_8283);
nor U8638 (N_8638,N_8452,N_8314);
or U8639 (N_8639,N_8432,N_8271);
xnor U8640 (N_8640,N_8342,N_8328);
nand U8641 (N_8641,N_8328,N_8363);
xnor U8642 (N_8642,N_8328,N_8335);
nor U8643 (N_8643,N_8427,N_8388);
or U8644 (N_8644,N_8315,N_8474);
or U8645 (N_8645,N_8391,N_8411);
nand U8646 (N_8646,N_8430,N_8305);
xnor U8647 (N_8647,N_8484,N_8412);
nand U8648 (N_8648,N_8276,N_8319);
xor U8649 (N_8649,N_8302,N_8463);
and U8650 (N_8650,N_8303,N_8395);
and U8651 (N_8651,N_8461,N_8402);
and U8652 (N_8652,N_8379,N_8301);
nor U8653 (N_8653,N_8362,N_8295);
or U8654 (N_8654,N_8412,N_8318);
or U8655 (N_8655,N_8405,N_8394);
xor U8656 (N_8656,N_8355,N_8383);
nand U8657 (N_8657,N_8324,N_8424);
nor U8658 (N_8658,N_8373,N_8405);
xor U8659 (N_8659,N_8452,N_8381);
xor U8660 (N_8660,N_8492,N_8328);
and U8661 (N_8661,N_8370,N_8268);
nand U8662 (N_8662,N_8337,N_8486);
xnor U8663 (N_8663,N_8483,N_8306);
nor U8664 (N_8664,N_8414,N_8278);
xnor U8665 (N_8665,N_8473,N_8406);
and U8666 (N_8666,N_8317,N_8457);
nand U8667 (N_8667,N_8309,N_8474);
and U8668 (N_8668,N_8406,N_8367);
or U8669 (N_8669,N_8254,N_8259);
nor U8670 (N_8670,N_8458,N_8373);
xor U8671 (N_8671,N_8413,N_8351);
xnor U8672 (N_8672,N_8364,N_8352);
and U8673 (N_8673,N_8290,N_8469);
xnor U8674 (N_8674,N_8304,N_8498);
nand U8675 (N_8675,N_8370,N_8421);
and U8676 (N_8676,N_8434,N_8260);
nor U8677 (N_8677,N_8395,N_8317);
nor U8678 (N_8678,N_8439,N_8465);
xnor U8679 (N_8679,N_8376,N_8299);
nand U8680 (N_8680,N_8363,N_8426);
nor U8681 (N_8681,N_8416,N_8308);
and U8682 (N_8682,N_8347,N_8441);
and U8683 (N_8683,N_8425,N_8457);
nor U8684 (N_8684,N_8278,N_8265);
nand U8685 (N_8685,N_8408,N_8317);
nor U8686 (N_8686,N_8365,N_8412);
or U8687 (N_8687,N_8376,N_8445);
nor U8688 (N_8688,N_8319,N_8448);
or U8689 (N_8689,N_8282,N_8436);
or U8690 (N_8690,N_8258,N_8370);
or U8691 (N_8691,N_8276,N_8401);
and U8692 (N_8692,N_8444,N_8357);
nor U8693 (N_8693,N_8348,N_8315);
xnor U8694 (N_8694,N_8257,N_8453);
or U8695 (N_8695,N_8449,N_8282);
xnor U8696 (N_8696,N_8293,N_8445);
or U8697 (N_8697,N_8426,N_8458);
or U8698 (N_8698,N_8354,N_8334);
and U8699 (N_8699,N_8346,N_8365);
nand U8700 (N_8700,N_8322,N_8368);
nand U8701 (N_8701,N_8460,N_8358);
or U8702 (N_8702,N_8258,N_8255);
nor U8703 (N_8703,N_8385,N_8290);
and U8704 (N_8704,N_8479,N_8411);
or U8705 (N_8705,N_8295,N_8484);
and U8706 (N_8706,N_8323,N_8357);
or U8707 (N_8707,N_8481,N_8295);
nand U8708 (N_8708,N_8444,N_8370);
and U8709 (N_8709,N_8420,N_8353);
and U8710 (N_8710,N_8299,N_8429);
nor U8711 (N_8711,N_8260,N_8476);
nand U8712 (N_8712,N_8470,N_8486);
and U8713 (N_8713,N_8332,N_8350);
xor U8714 (N_8714,N_8326,N_8436);
or U8715 (N_8715,N_8462,N_8268);
nand U8716 (N_8716,N_8354,N_8363);
and U8717 (N_8717,N_8491,N_8333);
nand U8718 (N_8718,N_8421,N_8380);
xor U8719 (N_8719,N_8445,N_8465);
and U8720 (N_8720,N_8327,N_8402);
and U8721 (N_8721,N_8444,N_8253);
nor U8722 (N_8722,N_8489,N_8463);
xnor U8723 (N_8723,N_8320,N_8476);
and U8724 (N_8724,N_8352,N_8405);
nand U8725 (N_8725,N_8454,N_8348);
nand U8726 (N_8726,N_8316,N_8312);
nand U8727 (N_8727,N_8438,N_8317);
and U8728 (N_8728,N_8278,N_8334);
xor U8729 (N_8729,N_8430,N_8338);
nor U8730 (N_8730,N_8264,N_8340);
or U8731 (N_8731,N_8498,N_8478);
xnor U8732 (N_8732,N_8471,N_8341);
xor U8733 (N_8733,N_8303,N_8389);
and U8734 (N_8734,N_8366,N_8384);
xnor U8735 (N_8735,N_8390,N_8422);
and U8736 (N_8736,N_8490,N_8491);
nor U8737 (N_8737,N_8253,N_8288);
xor U8738 (N_8738,N_8393,N_8361);
and U8739 (N_8739,N_8288,N_8312);
xor U8740 (N_8740,N_8470,N_8361);
xor U8741 (N_8741,N_8338,N_8494);
nand U8742 (N_8742,N_8274,N_8303);
or U8743 (N_8743,N_8429,N_8492);
and U8744 (N_8744,N_8389,N_8490);
and U8745 (N_8745,N_8352,N_8287);
xor U8746 (N_8746,N_8437,N_8474);
or U8747 (N_8747,N_8264,N_8266);
and U8748 (N_8748,N_8297,N_8340);
nand U8749 (N_8749,N_8447,N_8310);
xnor U8750 (N_8750,N_8711,N_8511);
nor U8751 (N_8751,N_8618,N_8748);
xnor U8752 (N_8752,N_8684,N_8653);
or U8753 (N_8753,N_8551,N_8547);
or U8754 (N_8754,N_8508,N_8506);
and U8755 (N_8755,N_8616,N_8633);
nand U8756 (N_8756,N_8699,N_8580);
nor U8757 (N_8757,N_8589,N_8505);
nor U8758 (N_8758,N_8529,N_8715);
and U8759 (N_8759,N_8746,N_8563);
xor U8760 (N_8760,N_8738,N_8745);
and U8761 (N_8761,N_8526,N_8610);
or U8762 (N_8762,N_8562,N_8736);
or U8763 (N_8763,N_8577,N_8679);
nand U8764 (N_8764,N_8724,N_8701);
nor U8765 (N_8765,N_8624,N_8688);
nor U8766 (N_8766,N_8602,N_8625);
xnor U8767 (N_8767,N_8622,N_8587);
nor U8768 (N_8768,N_8564,N_8513);
and U8769 (N_8769,N_8667,N_8716);
or U8770 (N_8770,N_8594,N_8747);
nand U8771 (N_8771,N_8559,N_8663);
nor U8772 (N_8772,N_8552,N_8630);
or U8773 (N_8773,N_8517,N_8582);
or U8774 (N_8774,N_8648,N_8600);
xor U8775 (N_8775,N_8675,N_8540);
and U8776 (N_8776,N_8612,N_8601);
nor U8777 (N_8777,N_8742,N_8683);
and U8778 (N_8778,N_8635,N_8509);
or U8779 (N_8779,N_8689,N_8717);
xnor U8780 (N_8780,N_8514,N_8703);
and U8781 (N_8781,N_8696,N_8518);
nand U8782 (N_8782,N_8500,N_8568);
nor U8783 (N_8783,N_8678,N_8671);
nand U8784 (N_8784,N_8535,N_8634);
nor U8785 (N_8785,N_8645,N_8655);
or U8786 (N_8786,N_8729,N_8673);
nand U8787 (N_8787,N_8543,N_8669);
nand U8788 (N_8788,N_8657,N_8569);
xnor U8789 (N_8789,N_8578,N_8520);
or U8790 (N_8790,N_8515,N_8672);
and U8791 (N_8791,N_8579,N_8565);
nand U8792 (N_8792,N_8640,N_8609);
or U8793 (N_8793,N_8560,N_8687);
or U8794 (N_8794,N_8694,N_8642);
xor U8795 (N_8795,N_8650,N_8607);
xnor U8796 (N_8796,N_8718,N_8593);
xor U8797 (N_8797,N_8561,N_8702);
or U8798 (N_8798,N_8503,N_8501);
or U8799 (N_8799,N_8712,N_8735);
nor U8800 (N_8800,N_8744,N_8682);
nor U8801 (N_8801,N_8660,N_8581);
nor U8802 (N_8802,N_8668,N_8629);
nor U8803 (N_8803,N_8659,N_8698);
or U8804 (N_8804,N_8725,N_8662);
or U8805 (N_8805,N_8544,N_8628);
xor U8806 (N_8806,N_8710,N_8567);
nor U8807 (N_8807,N_8566,N_8597);
nor U8808 (N_8808,N_8636,N_8727);
and U8809 (N_8809,N_8549,N_8697);
or U8810 (N_8810,N_8538,N_8583);
nand U8811 (N_8811,N_8680,N_8700);
nor U8812 (N_8812,N_8525,N_8739);
and U8813 (N_8813,N_8686,N_8615);
and U8814 (N_8814,N_8656,N_8714);
and U8815 (N_8815,N_8548,N_8627);
xor U8816 (N_8816,N_8596,N_8521);
and U8817 (N_8817,N_8510,N_8608);
nand U8818 (N_8818,N_8614,N_8741);
and U8819 (N_8819,N_8522,N_8644);
nor U8820 (N_8820,N_8732,N_8570);
or U8821 (N_8821,N_8512,N_8664);
or U8822 (N_8822,N_8652,N_8524);
nand U8823 (N_8823,N_8595,N_8527);
nand U8824 (N_8824,N_8626,N_8575);
xnor U8825 (N_8825,N_8558,N_8731);
nor U8826 (N_8826,N_8557,N_8542);
xor U8827 (N_8827,N_8619,N_8709);
xnor U8828 (N_8828,N_8692,N_8572);
nand U8829 (N_8829,N_8666,N_8553);
nand U8830 (N_8830,N_8523,N_8654);
xor U8831 (N_8831,N_8516,N_8533);
nor U8832 (N_8832,N_8705,N_8706);
and U8833 (N_8833,N_8685,N_8643);
and U8834 (N_8834,N_8519,N_8605);
or U8835 (N_8835,N_8591,N_8649);
and U8836 (N_8836,N_8647,N_8611);
and U8837 (N_8837,N_8658,N_8532);
or U8838 (N_8838,N_8599,N_8690);
nand U8839 (N_8839,N_8528,N_8681);
and U8840 (N_8840,N_8670,N_8720);
or U8841 (N_8841,N_8631,N_8584);
nor U8842 (N_8842,N_8740,N_8677);
or U8843 (N_8843,N_8555,N_8586);
nand U8844 (N_8844,N_8554,N_8545);
nor U8845 (N_8845,N_8536,N_8728);
nor U8846 (N_8846,N_8651,N_8691);
nor U8847 (N_8847,N_8620,N_8502);
nor U8848 (N_8848,N_8576,N_8541);
xnor U8849 (N_8849,N_8556,N_8623);
or U8850 (N_8850,N_8613,N_8638);
nand U8851 (N_8851,N_8530,N_8721);
and U8852 (N_8852,N_8598,N_8719);
or U8853 (N_8853,N_8639,N_8734);
or U8854 (N_8854,N_8621,N_8504);
xor U8855 (N_8855,N_8637,N_8585);
and U8856 (N_8856,N_8661,N_8592);
xor U8857 (N_8857,N_8507,N_8743);
xnor U8858 (N_8858,N_8604,N_8641);
and U8859 (N_8859,N_8606,N_8617);
xnor U8860 (N_8860,N_8588,N_8632);
and U8861 (N_8861,N_8574,N_8749);
nor U8862 (N_8862,N_8590,N_8546);
and U8863 (N_8863,N_8704,N_8707);
xnor U8864 (N_8864,N_8726,N_8730);
or U8865 (N_8865,N_8713,N_8573);
nor U8866 (N_8866,N_8693,N_8733);
and U8867 (N_8867,N_8646,N_8537);
nor U8868 (N_8868,N_8722,N_8571);
or U8869 (N_8869,N_8737,N_8676);
nor U8870 (N_8870,N_8674,N_8665);
or U8871 (N_8871,N_8539,N_8603);
and U8872 (N_8872,N_8531,N_8695);
nor U8873 (N_8873,N_8550,N_8723);
nor U8874 (N_8874,N_8708,N_8534);
or U8875 (N_8875,N_8652,N_8555);
or U8876 (N_8876,N_8611,N_8506);
nor U8877 (N_8877,N_8581,N_8545);
or U8878 (N_8878,N_8606,N_8519);
nor U8879 (N_8879,N_8506,N_8517);
xnor U8880 (N_8880,N_8596,N_8642);
xor U8881 (N_8881,N_8620,N_8611);
and U8882 (N_8882,N_8530,N_8685);
nor U8883 (N_8883,N_8551,N_8687);
nand U8884 (N_8884,N_8569,N_8580);
or U8885 (N_8885,N_8722,N_8584);
or U8886 (N_8886,N_8565,N_8668);
or U8887 (N_8887,N_8695,N_8742);
nor U8888 (N_8888,N_8732,N_8613);
and U8889 (N_8889,N_8744,N_8620);
xor U8890 (N_8890,N_8697,N_8552);
nand U8891 (N_8891,N_8723,N_8520);
nand U8892 (N_8892,N_8605,N_8647);
or U8893 (N_8893,N_8620,N_8683);
nor U8894 (N_8894,N_8699,N_8554);
nand U8895 (N_8895,N_8596,N_8639);
nand U8896 (N_8896,N_8635,N_8630);
xnor U8897 (N_8897,N_8674,N_8637);
nor U8898 (N_8898,N_8629,N_8735);
nand U8899 (N_8899,N_8556,N_8513);
xor U8900 (N_8900,N_8546,N_8663);
or U8901 (N_8901,N_8720,N_8507);
nor U8902 (N_8902,N_8683,N_8646);
nor U8903 (N_8903,N_8613,N_8560);
and U8904 (N_8904,N_8651,N_8537);
nor U8905 (N_8905,N_8649,N_8630);
nand U8906 (N_8906,N_8564,N_8537);
nand U8907 (N_8907,N_8585,N_8706);
or U8908 (N_8908,N_8612,N_8606);
xor U8909 (N_8909,N_8698,N_8600);
and U8910 (N_8910,N_8640,N_8568);
nor U8911 (N_8911,N_8500,N_8734);
and U8912 (N_8912,N_8503,N_8706);
nor U8913 (N_8913,N_8701,N_8715);
nor U8914 (N_8914,N_8589,N_8724);
and U8915 (N_8915,N_8545,N_8600);
nand U8916 (N_8916,N_8559,N_8582);
nor U8917 (N_8917,N_8655,N_8641);
nand U8918 (N_8918,N_8591,N_8734);
xor U8919 (N_8919,N_8648,N_8578);
nor U8920 (N_8920,N_8646,N_8651);
and U8921 (N_8921,N_8542,N_8720);
nand U8922 (N_8922,N_8589,N_8556);
nor U8923 (N_8923,N_8712,N_8556);
nor U8924 (N_8924,N_8629,N_8747);
and U8925 (N_8925,N_8618,N_8650);
xnor U8926 (N_8926,N_8516,N_8654);
nand U8927 (N_8927,N_8719,N_8572);
nand U8928 (N_8928,N_8532,N_8721);
nor U8929 (N_8929,N_8506,N_8521);
and U8930 (N_8930,N_8550,N_8503);
or U8931 (N_8931,N_8654,N_8717);
and U8932 (N_8932,N_8554,N_8510);
nor U8933 (N_8933,N_8735,N_8626);
nand U8934 (N_8934,N_8745,N_8731);
xor U8935 (N_8935,N_8612,N_8717);
and U8936 (N_8936,N_8709,N_8719);
or U8937 (N_8937,N_8502,N_8722);
and U8938 (N_8938,N_8549,N_8622);
and U8939 (N_8939,N_8628,N_8585);
nand U8940 (N_8940,N_8717,N_8500);
or U8941 (N_8941,N_8722,N_8564);
nand U8942 (N_8942,N_8734,N_8718);
nor U8943 (N_8943,N_8692,N_8641);
nand U8944 (N_8944,N_8547,N_8511);
xnor U8945 (N_8945,N_8711,N_8690);
nand U8946 (N_8946,N_8679,N_8747);
and U8947 (N_8947,N_8581,N_8594);
or U8948 (N_8948,N_8626,N_8660);
nand U8949 (N_8949,N_8723,N_8615);
nor U8950 (N_8950,N_8621,N_8573);
xor U8951 (N_8951,N_8678,N_8642);
nand U8952 (N_8952,N_8743,N_8500);
and U8953 (N_8953,N_8557,N_8735);
xor U8954 (N_8954,N_8731,N_8703);
xor U8955 (N_8955,N_8645,N_8609);
nor U8956 (N_8956,N_8652,N_8515);
and U8957 (N_8957,N_8539,N_8618);
or U8958 (N_8958,N_8672,N_8530);
or U8959 (N_8959,N_8687,N_8746);
nand U8960 (N_8960,N_8648,N_8634);
nand U8961 (N_8961,N_8632,N_8542);
and U8962 (N_8962,N_8736,N_8507);
nor U8963 (N_8963,N_8608,N_8670);
xnor U8964 (N_8964,N_8673,N_8508);
and U8965 (N_8965,N_8711,N_8633);
nor U8966 (N_8966,N_8529,N_8675);
nand U8967 (N_8967,N_8629,N_8647);
or U8968 (N_8968,N_8643,N_8519);
xnor U8969 (N_8969,N_8630,N_8507);
xor U8970 (N_8970,N_8571,N_8668);
and U8971 (N_8971,N_8665,N_8673);
nand U8972 (N_8972,N_8714,N_8557);
xor U8973 (N_8973,N_8514,N_8657);
and U8974 (N_8974,N_8715,N_8625);
or U8975 (N_8975,N_8543,N_8626);
nand U8976 (N_8976,N_8705,N_8555);
nor U8977 (N_8977,N_8547,N_8561);
and U8978 (N_8978,N_8561,N_8674);
nand U8979 (N_8979,N_8626,N_8711);
nand U8980 (N_8980,N_8647,N_8669);
and U8981 (N_8981,N_8567,N_8706);
xnor U8982 (N_8982,N_8658,N_8701);
nor U8983 (N_8983,N_8552,N_8521);
nand U8984 (N_8984,N_8569,N_8661);
nor U8985 (N_8985,N_8575,N_8514);
xnor U8986 (N_8986,N_8730,N_8646);
xor U8987 (N_8987,N_8720,N_8561);
and U8988 (N_8988,N_8710,N_8602);
and U8989 (N_8989,N_8660,N_8680);
xnor U8990 (N_8990,N_8541,N_8650);
and U8991 (N_8991,N_8545,N_8744);
or U8992 (N_8992,N_8565,N_8740);
nand U8993 (N_8993,N_8624,N_8617);
xnor U8994 (N_8994,N_8726,N_8665);
xnor U8995 (N_8995,N_8660,N_8745);
nand U8996 (N_8996,N_8528,N_8603);
nor U8997 (N_8997,N_8711,N_8532);
or U8998 (N_8998,N_8573,N_8633);
nand U8999 (N_8999,N_8614,N_8602);
and U9000 (N_9000,N_8787,N_8900);
or U9001 (N_9001,N_8825,N_8805);
nor U9002 (N_9002,N_8903,N_8797);
nor U9003 (N_9003,N_8931,N_8830);
nand U9004 (N_9004,N_8909,N_8885);
nand U9005 (N_9005,N_8881,N_8906);
or U9006 (N_9006,N_8877,N_8939);
or U9007 (N_9007,N_8803,N_8934);
nor U9008 (N_9008,N_8936,N_8827);
and U9009 (N_9009,N_8769,N_8995);
nand U9010 (N_9010,N_8776,N_8879);
nor U9011 (N_9011,N_8831,N_8937);
or U9012 (N_9012,N_8772,N_8821);
and U9013 (N_9013,N_8959,N_8976);
and U9014 (N_9014,N_8948,N_8849);
xor U9015 (N_9015,N_8893,N_8818);
or U9016 (N_9016,N_8897,N_8929);
nor U9017 (N_9017,N_8910,N_8895);
and U9018 (N_9018,N_8800,N_8779);
and U9019 (N_9019,N_8832,N_8771);
xnor U9020 (N_9020,N_8853,N_8971);
nor U9021 (N_9021,N_8878,N_8850);
xor U9022 (N_9022,N_8894,N_8997);
nor U9023 (N_9023,N_8943,N_8819);
and U9024 (N_9024,N_8915,N_8801);
xor U9025 (N_9025,N_8998,N_8784);
xnor U9026 (N_9026,N_8980,N_8880);
or U9027 (N_9027,N_8780,N_8923);
and U9028 (N_9028,N_8872,N_8814);
and U9029 (N_9029,N_8911,N_8858);
nor U9030 (N_9030,N_8761,N_8945);
nand U9031 (N_9031,N_8927,N_8951);
xnor U9032 (N_9032,N_8925,N_8790);
nor U9033 (N_9033,N_8773,N_8802);
and U9034 (N_9034,N_8975,N_8752);
nor U9035 (N_9035,N_8846,N_8826);
nor U9036 (N_9036,N_8969,N_8992);
nand U9037 (N_9037,N_8860,N_8989);
nor U9038 (N_9038,N_8793,N_8766);
or U9039 (N_9039,N_8755,N_8857);
xor U9040 (N_9040,N_8875,N_8839);
xor U9041 (N_9041,N_8926,N_8918);
xnor U9042 (N_9042,N_8843,N_8859);
nor U9043 (N_9043,N_8938,N_8847);
and U9044 (N_9044,N_8952,N_8987);
nand U9045 (N_9045,N_8891,N_8774);
xor U9046 (N_9046,N_8810,N_8892);
nor U9047 (N_9047,N_8941,N_8977);
or U9048 (N_9048,N_8753,N_8956);
or U9049 (N_9049,N_8901,N_8867);
or U9050 (N_9050,N_8795,N_8981);
xnor U9051 (N_9051,N_8905,N_8777);
nor U9052 (N_9052,N_8794,N_8796);
nor U9053 (N_9053,N_8986,N_8838);
xnor U9054 (N_9054,N_8770,N_8913);
and U9055 (N_9055,N_8815,N_8767);
nand U9056 (N_9056,N_8882,N_8865);
nor U9057 (N_9057,N_8807,N_8876);
nand U9058 (N_9058,N_8829,N_8778);
and U9059 (N_9059,N_8908,N_8788);
nand U9060 (N_9060,N_8984,N_8896);
or U9061 (N_9061,N_8904,N_8965);
nor U9062 (N_9062,N_8811,N_8841);
xnor U9063 (N_9063,N_8874,N_8845);
nor U9064 (N_9064,N_8763,N_8968);
nor U9065 (N_9065,N_8791,N_8933);
xnor U9066 (N_9066,N_8883,N_8957);
xor U9067 (N_9067,N_8963,N_8994);
nor U9068 (N_9068,N_8768,N_8823);
nand U9069 (N_9069,N_8862,N_8828);
xor U9070 (N_9070,N_8789,N_8835);
xnor U9071 (N_9071,N_8960,N_8855);
and U9072 (N_9072,N_8961,N_8754);
or U9073 (N_9073,N_8804,N_8886);
xor U9074 (N_9074,N_8983,N_8812);
nor U9075 (N_9075,N_8813,N_8889);
xnor U9076 (N_9076,N_8912,N_8928);
nor U9077 (N_9077,N_8873,N_8834);
nor U9078 (N_9078,N_8944,N_8757);
nor U9079 (N_9079,N_8820,N_8932);
nor U9080 (N_9080,N_8982,N_8864);
or U9081 (N_9081,N_8851,N_8863);
or U9082 (N_9082,N_8848,N_8781);
or U9083 (N_9083,N_8840,N_8852);
nor U9084 (N_9084,N_8972,N_8762);
nor U9085 (N_9085,N_8954,N_8868);
nor U9086 (N_9086,N_8764,N_8887);
and U9087 (N_9087,N_8988,N_8884);
nor U9088 (N_9088,N_8962,N_8782);
and U9089 (N_9089,N_8817,N_8899);
nor U9090 (N_9090,N_8760,N_8970);
nand U9091 (N_9091,N_8833,N_8750);
or U9092 (N_9092,N_8898,N_8861);
nand U9093 (N_9093,N_8870,N_8759);
and U9094 (N_9094,N_8783,N_8964);
xnor U9095 (N_9095,N_8775,N_8993);
or U9096 (N_9096,N_8888,N_8955);
xor U9097 (N_9097,N_8974,N_8999);
xnor U9098 (N_9098,N_8798,N_8990);
or U9099 (N_9099,N_8914,N_8949);
xnor U9100 (N_9100,N_8921,N_8917);
xor U9101 (N_9101,N_8940,N_8942);
and U9102 (N_9102,N_8996,N_8924);
nand U9103 (N_9103,N_8935,N_8785);
nand U9104 (N_9104,N_8973,N_8946);
or U9105 (N_9105,N_8837,N_8966);
xor U9106 (N_9106,N_8958,N_8919);
nor U9107 (N_9107,N_8922,N_8786);
xnor U9108 (N_9108,N_8842,N_8758);
or U9109 (N_9109,N_8751,N_8808);
nor U9110 (N_9110,N_8950,N_8916);
and U9111 (N_9111,N_8856,N_8869);
and U9112 (N_9112,N_8866,N_8978);
xnor U9113 (N_9113,N_8902,N_8836);
or U9114 (N_9114,N_8756,N_8967);
nor U9115 (N_9115,N_8871,N_8947);
xnor U9116 (N_9116,N_8806,N_8822);
and U9117 (N_9117,N_8930,N_8907);
xor U9118 (N_9118,N_8792,N_8824);
and U9119 (N_9119,N_8890,N_8799);
nand U9120 (N_9120,N_8979,N_8765);
and U9121 (N_9121,N_8816,N_8953);
xnor U9122 (N_9122,N_8844,N_8985);
or U9123 (N_9123,N_8920,N_8809);
or U9124 (N_9124,N_8991,N_8854);
xnor U9125 (N_9125,N_8750,N_8807);
nand U9126 (N_9126,N_8798,N_8789);
or U9127 (N_9127,N_8839,N_8829);
or U9128 (N_9128,N_8750,N_8765);
nand U9129 (N_9129,N_8862,N_8779);
xor U9130 (N_9130,N_8824,N_8944);
nand U9131 (N_9131,N_8900,N_8990);
nor U9132 (N_9132,N_8875,N_8794);
or U9133 (N_9133,N_8827,N_8901);
and U9134 (N_9134,N_8811,N_8761);
xnor U9135 (N_9135,N_8908,N_8930);
and U9136 (N_9136,N_8914,N_8894);
nand U9137 (N_9137,N_8996,N_8794);
nor U9138 (N_9138,N_8778,N_8815);
nand U9139 (N_9139,N_8891,N_8804);
and U9140 (N_9140,N_8981,N_8909);
xor U9141 (N_9141,N_8835,N_8898);
xnor U9142 (N_9142,N_8836,N_8800);
nand U9143 (N_9143,N_8989,N_8809);
xnor U9144 (N_9144,N_8751,N_8901);
nand U9145 (N_9145,N_8841,N_8789);
nand U9146 (N_9146,N_8928,N_8821);
or U9147 (N_9147,N_8751,N_8989);
and U9148 (N_9148,N_8867,N_8955);
nor U9149 (N_9149,N_8949,N_8807);
xor U9150 (N_9150,N_8803,N_8859);
nand U9151 (N_9151,N_8768,N_8829);
or U9152 (N_9152,N_8776,N_8892);
or U9153 (N_9153,N_8943,N_8790);
nor U9154 (N_9154,N_8876,N_8988);
and U9155 (N_9155,N_8764,N_8804);
or U9156 (N_9156,N_8888,N_8943);
xor U9157 (N_9157,N_8848,N_8962);
nand U9158 (N_9158,N_8777,N_8768);
xnor U9159 (N_9159,N_8922,N_8857);
xor U9160 (N_9160,N_8952,N_8906);
nor U9161 (N_9161,N_8858,N_8820);
and U9162 (N_9162,N_8751,N_8972);
or U9163 (N_9163,N_8989,N_8879);
nand U9164 (N_9164,N_8861,N_8970);
xor U9165 (N_9165,N_8966,N_8962);
and U9166 (N_9166,N_8757,N_8824);
xnor U9167 (N_9167,N_8991,N_8793);
nor U9168 (N_9168,N_8787,N_8959);
nor U9169 (N_9169,N_8943,N_8863);
and U9170 (N_9170,N_8917,N_8894);
and U9171 (N_9171,N_8961,N_8765);
or U9172 (N_9172,N_8833,N_8782);
nand U9173 (N_9173,N_8923,N_8791);
or U9174 (N_9174,N_8998,N_8839);
and U9175 (N_9175,N_8803,N_8879);
xnor U9176 (N_9176,N_8868,N_8929);
or U9177 (N_9177,N_8938,N_8884);
and U9178 (N_9178,N_8845,N_8974);
or U9179 (N_9179,N_8781,N_8963);
and U9180 (N_9180,N_8859,N_8801);
nor U9181 (N_9181,N_8808,N_8987);
xnor U9182 (N_9182,N_8881,N_8761);
xnor U9183 (N_9183,N_8837,N_8893);
or U9184 (N_9184,N_8785,N_8817);
and U9185 (N_9185,N_8865,N_8794);
nand U9186 (N_9186,N_8792,N_8754);
xor U9187 (N_9187,N_8805,N_8965);
nor U9188 (N_9188,N_8999,N_8947);
xnor U9189 (N_9189,N_8910,N_8937);
and U9190 (N_9190,N_8929,N_8845);
nor U9191 (N_9191,N_8879,N_8823);
and U9192 (N_9192,N_8859,N_8766);
or U9193 (N_9193,N_8998,N_8840);
or U9194 (N_9194,N_8780,N_8993);
or U9195 (N_9195,N_8956,N_8995);
nand U9196 (N_9196,N_8892,N_8954);
nor U9197 (N_9197,N_8927,N_8785);
xnor U9198 (N_9198,N_8852,N_8853);
xnor U9199 (N_9199,N_8878,N_8796);
or U9200 (N_9200,N_8921,N_8939);
nor U9201 (N_9201,N_8967,N_8947);
nand U9202 (N_9202,N_8778,N_8949);
or U9203 (N_9203,N_8914,N_8934);
nor U9204 (N_9204,N_8757,N_8765);
nor U9205 (N_9205,N_8955,N_8851);
xor U9206 (N_9206,N_8977,N_8938);
nand U9207 (N_9207,N_8792,N_8804);
and U9208 (N_9208,N_8965,N_8897);
nand U9209 (N_9209,N_8873,N_8837);
nand U9210 (N_9210,N_8917,N_8829);
xor U9211 (N_9211,N_8815,N_8930);
xnor U9212 (N_9212,N_8931,N_8929);
xor U9213 (N_9213,N_8906,N_8962);
and U9214 (N_9214,N_8939,N_8858);
nor U9215 (N_9215,N_8753,N_8830);
or U9216 (N_9216,N_8842,N_8893);
and U9217 (N_9217,N_8969,N_8829);
and U9218 (N_9218,N_8920,N_8848);
or U9219 (N_9219,N_8913,N_8763);
nand U9220 (N_9220,N_8892,N_8804);
xor U9221 (N_9221,N_8750,N_8788);
or U9222 (N_9222,N_8844,N_8819);
or U9223 (N_9223,N_8890,N_8911);
nand U9224 (N_9224,N_8890,N_8931);
and U9225 (N_9225,N_8910,N_8815);
or U9226 (N_9226,N_8756,N_8968);
and U9227 (N_9227,N_8791,N_8938);
xor U9228 (N_9228,N_8945,N_8785);
or U9229 (N_9229,N_8840,N_8809);
nand U9230 (N_9230,N_8788,N_8886);
xor U9231 (N_9231,N_8783,N_8891);
or U9232 (N_9232,N_8864,N_8914);
nor U9233 (N_9233,N_8947,N_8905);
or U9234 (N_9234,N_8797,N_8994);
nand U9235 (N_9235,N_8936,N_8759);
and U9236 (N_9236,N_8887,N_8821);
nor U9237 (N_9237,N_8874,N_8972);
and U9238 (N_9238,N_8763,N_8975);
xnor U9239 (N_9239,N_8982,N_8847);
nand U9240 (N_9240,N_8839,N_8906);
nand U9241 (N_9241,N_8994,N_8810);
nand U9242 (N_9242,N_8991,N_8770);
nand U9243 (N_9243,N_8798,N_8833);
and U9244 (N_9244,N_8985,N_8924);
nor U9245 (N_9245,N_8961,N_8785);
nor U9246 (N_9246,N_8795,N_8847);
xnor U9247 (N_9247,N_8970,N_8851);
nand U9248 (N_9248,N_8954,N_8983);
nor U9249 (N_9249,N_8756,N_8777);
nand U9250 (N_9250,N_9045,N_9104);
and U9251 (N_9251,N_9096,N_9042);
or U9252 (N_9252,N_9224,N_9161);
and U9253 (N_9253,N_9182,N_9032);
or U9254 (N_9254,N_9015,N_9158);
nand U9255 (N_9255,N_9036,N_9072);
nand U9256 (N_9256,N_9165,N_9085);
or U9257 (N_9257,N_9133,N_9120);
xor U9258 (N_9258,N_9092,N_9172);
nor U9259 (N_9259,N_9209,N_9213);
or U9260 (N_9260,N_9138,N_9014);
and U9261 (N_9261,N_9047,N_9062);
nand U9262 (N_9262,N_9013,N_9060);
or U9263 (N_9263,N_9073,N_9067);
nand U9264 (N_9264,N_9169,N_9126);
xor U9265 (N_9265,N_9152,N_9191);
nor U9266 (N_9266,N_9123,N_9214);
and U9267 (N_9267,N_9043,N_9156);
nand U9268 (N_9268,N_9184,N_9210);
or U9269 (N_9269,N_9022,N_9219);
nand U9270 (N_9270,N_9054,N_9121);
nand U9271 (N_9271,N_9241,N_9141);
or U9272 (N_9272,N_9239,N_9159);
nand U9273 (N_9273,N_9164,N_9175);
nand U9274 (N_9274,N_9140,N_9134);
nor U9275 (N_9275,N_9094,N_9147);
or U9276 (N_9276,N_9245,N_9232);
and U9277 (N_9277,N_9129,N_9021);
xor U9278 (N_9278,N_9075,N_9144);
xnor U9279 (N_9279,N_9160,N_9145);
nor U9280 (N_9280,N_9052,N_9176);
and U9281 (N_9281,N_9193,N_9207);
nor U9282 (N_9282,N_9248,N_9227);
or U9283 (N_9283,N_9098,N_9171);
and U9284 (N_9284,N_9064,N_9105);
nand U9285 (N_9285,N_9007,N_9202);
nand U9286 (N_9286,N_9135,N_9142);
nor U9287 (N_9287,N_9058,N_9185);
or U9288 (N_9288,N_9137,N_9153);
xor U9289 (N_9289,N_9222,N_9003);
nor U9290 (N_9290,N_9183,N_9076);
nand U9291 (N_9291,N_9125,N_9243);
nor U9292 (N_9292,N_9132,N_9055);
nor U9293 (N_9293,N_9034,N_9056);
and U9294 (N_9294,N_9107,N_9231);
and U9295 (N_9295,N_9100,N_9217);
and U9296 (N_9296,N_9151,N_9087);
or U9297 (N_9297,N_9127,N_9012);
nand U9298 (N_9298,N_9017,N_9074);
nand U9299 (N_9299,N_9097,N_9167);
and U9300 (N_9300,N_9106,N_9149);
and U9301 (N_9301,N_9061,N_9068);
or U9302 (N_9302,N_9208,N_9101);
and U9303 (N_9303,N_9095,N_9071);
nor U9304 (N_9304,N_9069,N_9089);
xnor U9305 (N_9305,N_9242,N_9001);
nor U9306 (N_9306,N_9238,N_9166);
or U9307 (N_9307,N_9008,N_9006);
nand U9308 (N_9308,N_9139,N_9170);
and U9309 (N_9309,N_9025,N_9240);
xor U9310 (N_9310,N_9016,N_9244);
or U9311 (N_9311,N_9024,N_9011);
nand U9312 (N_9312,N_9163,N_9146);
nor U9313 (N_9313,N_9143,N_9118);
nand U9314 (N_9314,N_9004,N_9028);
and U9315 (N_9315,N_9194,N_9044);
and U9316 (N_9316,N_9178,N_9131);
nand U9317 (N_9317,N_9122,N_9216);
nand U9318 (N_9318,N_9057,N_9174);
and U9319 (N_9319,N_9198,N_9203);
nor U9320 (N_9320,N_9093,N_9235);
nand U9321 (N_9321,N_9080,N_9115);
and U9322 (N_9322,N_9037,N_9220);
xnor U9323 (N_9323,N_9188,N_9030);
nor U9324 (N_9324,N_9070,N_9031);
xor U9325 (N_9325,N_9005,N_9078);
nor U9326 (N_9326,N_9228,N_9099);
nand U9327 (N_9327,N_9090,N_9002);
nand U9328 (N_9328,N_9181,N_9212);
or U9329 (N_9329,N_9130,N_9082);
nor U9330 (N_9330,N_9218,N_9205);
xnor U9331 (N_9331,N_9091,N_9223);
or U9332 (N_9332,N_9000,N_9230);
nor U9333 (N_9333,N_9081,N_9050);
nor U9334 (N_9334,N_9117,N_9150);
xnor U9335 (N_9335,N_9168,N_9204);
nand U9336 (N_9336,N_9136,N_9112);
and U9337 (N_9337,N_9116,N_9221);
or U9338 (N_9338,N_9103,N_9211);
xnor U9339 (N_9339,N_9053,N_9246);
or U9340 (N_9340,N_9051,N_9083);
nand U9341 (N_9341,N_9110,N_9111);
and U9342 (N_9342,N_9079,N_9088);
and U9343 (N_9343,N_9019,N_9148);
or U9344 (N_9344,N_9114,N_9086);
nand U9345 (N_9345,N_9234,N_9201);
xnor U9346 (N_9346,N_9236,N_9084);
xnor U9347 (N_9347,N_9187,N_9066);
and U9348 (N_9348,N_9010,N_9195);
xnor U9349 (N_9349,N_9077,N_9200);
or U9350 (N_9350,N_9197,N_9109);
nor U9351 (N_9351,N_9196,N_9237);
nand U9352 (N_9352,N_9018,N_9199);
xnor U9353 (N_9353,N_9046,N_9038);
or U9354 (N_9354,N_9128,N_9226);
and U9355 (N_9355,N_9177,N_9192);
nand U9356 (N_9356,N_9040,N_9225);
nor U9357 (N_9357,N_9119,N_9155);
or U9358 (N_9358,N_9059,N_9157);
nor U9359 (N_9359,N_9039,N_9162);
xnor U9360 (N_9360,N_9154,N_9180);
nor U9361 (N_9361,N_9065,N_9108);
or U9362 (N_9362,N_9215,N_9189);
nand U9363 (N_9363,N_9049,N_9033);
and U9364 (N_9364,N_9035,N_9029);
xnor U9365 (N_9365,N_9190,N_9041);
nand U9366 (N_9366,N_9113,N_9186);
or U9367 (N_9367,N_9048,N_9124);
and U9368 (N_9368,N_9027,N_9247);
nand U9369 (N_9369,N_9063,N_9173);
or U9370 (N_9370,N_9229,N_9023);
nand U9371 (N_9371,N_9206,N_9249);
nand U9372 (N_9372,N_9102,N_9020);
nor U9373 (N_9373,N_9179,N_9026);
xnor U9374 (N_9374,N_9233,N_9009);
nand U9375 (N_9375,N_9085,N_9083);
xnor U9376 (N_9376,N_9127,N_9083);
nand U9377 (N_9377,N_9056,N_9040);
or U9378 (N_9378,N_9148,N_9048);
or U9379 (N_9379,N_9029,N_9207);
and U9380 (N_9380,N_9243,N_9120);
nor U9381 (N_9381,N_9238,N_9173);
nor U9382 (N_9382,N_9009,N_9131);
and U9383 (N_9383,N_9140,N_9215);
nand U9384 (N_9384,N_9198,N_9020);
and U9385 (N_9385,N_9002,N_9156);
xnor U9386 (N_9386,N_9174,N_9185);
or U9387 (N_9387,N_9113,N_9220);
or U9388 (N_9388,N_9240,N_9201);
nand U9389 (N_9389,N_9057,N_9082);
nor U9390 (N_9390,N_9056,N_9038);
nor U9391 (N_9391,N_9175,N_9024);
xnor U9392 (N_9392,N_9200,N_9171);
and U9393 (N_9393,N_9245,N_9200);
nor U9394 (N_9394,N_9082,N_9247);
nand U9395 (N_9395,N_9074,N_9122);
nand U9396 (N_9396,N_9094,N_9231);
xor U9397 (N_9397,N_9121,N_9128);
nand U9398 (N_9398,N_9191,N_9200);
and U9399 (N_9399,N_9219,N_9009);
xor U9400 (N_9400,N_9103,N_9075);
or U9401 (N_9401,N_9019,N_9196);
and U9402 (N_9402,N_9035,N_9161);
nor U9403 (N_9403,N_9103,N_9021);
or U9404 (N_9404,N_9061,N_9182);
or U9405 (N_9405,N_9245,N_9167);
xor U9406 (N_9406,N_9113,N_9233);
nor U9407 (N_9407,N_9084,N_9058);
and U9408 (N_9408,N_9083,N_9055);
or U9409 (N_9409,N_9031,N_9162);
nand U9410 (N_9410,N_9189,N_9137);
xnor U9411 (N_9411,N_9141,N_9077);
nor U9412 (N_9412,N_9073,N_9064);
nand U9413 (N_9413,N_9180,N_9106);
nor U9414 (N_9414,N_9156,N_9206);
nor U9415 (N_9415,N_9227,N_9107);
nand U9416 (N_9416,N_9115,N_9150);
nor U9417 (N_9417,N_9071,N_9195);
nand U9418 (N_9418,N_9088,N_9248);
nor U9419 (N_9419,N_9084,N_9182);
and U9420 (N_9420,N_9110,N_9218);
nand U9421 (N_9421,N_9207,N_9140);
or U9422 (N_9422,N_9242,N_9137);
nor U9423 (N_9423,N_9173,N_9016);
or U9424 (N_9424,N_9013,N_9221);
and U9425 (N_9425,N_9107,N_9061);
or U9426 (N_9426,N_9009,N_9170);
nand U9427 (N_9427,N_9169,N_9172);
or U9428 (N_9428,N_9163,N_9178);
or U9429 (N_9429,N_9222,N_9086);
or U9430 (N_9430,N_9195,N_9024);
xnor U9431 (N_9431,N_9112,N_9148);
and U9432 (N_9432,N_9118,N_9049);
xnor U9433 (N_9433,N_9164,N_9160);
nor U9434 (N_9434,N_9134,N_9190);
nor U9435 (N_9435,N_9125,N_9215);
nor U9436 (N_9436,N_9167,N_9240);
and U9437 (N_9437,N_9085,N_9011);
nand U9438 (N_9438,N_9068,N_9156);
xor U9439 (N_9439,N_9225,N_9223);
and U9440 (N_9440,N_9033,N_9108);
nand U9441 (N_9441,N_9205,N_9128);
xnor U9442 (N_9442,N_9235,N_9106);
or U9443 (N_9443,N_9017,N_9090);
and U9444 (N_9444,N_9123,N_9022);
xor U9445 (N_9445,N_9045,N_9059);
xnor U9446 (N_9446,N_9233,N_9100);
nand U9447 (N_9447,N_9084,N_9033);
nand U9448 (N_9448,N_9224,N_9009);
and U9449 (N_9449,N_9218,N_9189);
nor U9450 (N_9450,N_9236,N_9119);
xor U9451 (N_9451,N_9084,N_9080);
or U9452 (N_9452,N_9001,N_9012);
xnor U9453 (N_9453,N_9162,N_9134);
or U9454 (N_9454,N_9164,N_9052);
or U9455 (N_9455,N_9123,N_9176);
and U9456 (N_9456,N_9248,N_9027);
nand U9457 (N_9457,N_9153,N_9218);
xor U9458 (N_9458,N_9025,N_9097);
and U9459 (N_9459,N_9245,N_9078);
nand U9460 (N_9460,N_9073,N_9128);
and U9461 (N_9461,N_9072,N_9234);
xnor U9462 (N_9462,N_9118,N_9195);
nor U9463 (N_9463,N_9025,N_9022);
nand U9464 (N_9464,N_9178,N_9165);
nand U9465 (N_9465,N_9052,N_9214);
xor U9466 (N_9466,N_9229,N_9039);
or U9467 (N_9467,N_9128,N_9002);
nand U9468 (N_9468,N_9084,N_9094);
nand U9469 (N_9469,N_9184,N_9153);
and U9470 (N_9470,N_9073,N_9124);
nor U9471 (N_9471,N_9035,N_9220);
or U9472 (N_9472,N_9035,N_9247);
xor U9473 (N_9473,N_9184,N_9171);
xnor U9474 (N_9474,N_9100,N_9017);
nor U9475 (N_9475,N_9113,N_9079);
nor U9476 (N_9476,N_9226,N_9161);
nor U9477 (N_9477,N_9139,N_9093);
or U9478 (N_9478,N_9045,N_9216);
or U9479 (N_9479,N_9018,N_9017);
nand U9480 (N_9480,N_9085,N_9088);
and U9481 (N_9481,N_9206,N_9237);
xor U9482 (N_9482,N_9162,N_9237);
or U9483 (N_9483,N_9182,N_9108);
xnor U9484 (N_9484,N_9225,N_9074);
nor U9485 (N_9485,N_9184,N_9015);
and U9486 (N_9486,N_9009,N_9207);
xor U9487 (N_9487,N_9162,N_9087);
and U9488 (N_9488,N_9074,N_9045);
xor U9489 (N_9489,N_9044,N_9033);
and U9490 (N_9490,N_9147,N_9050);
or U9491 (N_9491,N_9049,N_9028);
xor U9492 (N_9492,N_9062,N_9201);
and U9493 (N_9493,N_9070,N_9086);
and U9494 (N_9494,N_9025,N_9149);
or U9495 (N_9495,N_9032,N_9185);
nor U9496 (N_9496,N_9087,N_9126);
nand U9497 (N_9497,N_9072,N_9070);
and U9498 (N_9498,N_9206,N_9178);
nand U9499 (N_9499,N_9143,N_9240);
nand U9500 (N_9500,N_9354,N_9384);
xnor U9501 (N_9501,N_9256,N_9334);
xnor U9502 (N_9502,N_9411,N_9376);
and U9503 (N_9503,N_9355,N_9497);
and U9504 (N_9504,N_9313,N_9358);
and U9505 (N_9505,N_9270,N_9438);
and U9506 (N_9506,N_9476,N_9449);
and U9507 (N_9507,N_9262,N_9283);
nor U9508 (N_9508,N_9275,N_9265);
and U9509 (N_9509,N_9378,N_9442);
and U9510 (N_9510,N_9474,N_9401);
or U9511 (N_9511,N_9272,N_9302);
nor U9512 (N_9512,N_9426,N_9499);
nand U9513 (N_9513,N_9435,N_9261);
nand U9514 (N_9514,N_9319,N_9407);
and U9515 (N_9515,N_9306,N_9473);
or U9516 (N_9516,N_9260,N_9255);
xor U9517 (N_9517,N_9338,N_9316);
or U9518 (N_9518,N_9364,N_9361);
nand U9519 (N_9519,N_9267,N_9429);
nor U9520 (N_9520,N_9370,N_9408);
or U9521 (N_9521,N_9336,N_9337);
nand U9522 (N_9522,N_9252,N_9277);
or U9523 (N_9523,N_9397,N_9367);
and U9524 (N_9524,N_9259,N_9434);
nor U9525 (N_9525,N_9314,N_9431);
nor U9526 (N_9526,N_9460,N_9420);
nand U9527 (N_9527,N_9415,N_9357);
or U9528 (N_9528,N_9375,N_9471);
xor U9529 (N_9529,N_9414,N_9379);
nor U9530 (N_9530,N_9341,N_9463);
or U9531 (N_9531,N_9305,N_9496);
and U9532 (N_9532,N_9482,N_9441);
nor U9533 (N_9533,N_9383,N_9391);
nand U9534 (N_9534,N_9273,N_9439);
nor U9535 (N_9535,N_9263,N_9294);
and U9536 (N_9536,N_9444,N_9381);
or U9537 (N_9537,N_9393,N_9394);
nor U9538 (N_9538,N_9349,N_9284);
and U9539 (N_9539,N_9418,N_9369);
nor U9540 (N_9540,N_9345,N_9329);
xnor U9541 (N_9541,N_9488,N_9390);
or U9542 (N_9542,N_9322,N_9455);
and U9543 (N_9543,N_9288,N_9350);
xor U9544 (N_9544,N_9328,N_9333);
and U9545 (N_9545,N_9368,N_9347);
nand U9546 (N_9546,N_9320,N_9484);
nand U9547 (N_9547,N_9392,N_9280);
or U9548 (N_9548,N_9312,N_9366);
nor U9549 (N_9549,N_9400,N_9303);
nor U9550 (N_9550,N_9459,N_9486);
nand U9551 (N_9551,N_9469,N_9371);
and U9552 (N_9552,N_9396,N_9282);
and U9553 (N_9553,N_9290,N_9285);
nand U9554 (N_9554,N_9492,N_9413);
xor U9555 (N_9555,N_9352,N_9271);
nor U9556 (N_9556,N_9300,N_9268);
nor U9557 (N_9557,N_9296,N_9462);
and U9558 (N_9558,N_9250,N_9385);
and U9559 (N_9559,N_9377,N_9477);
or U9560 (N_9560,N_9269,N_9495);
xnor U9561 (N_9561,N_9339,N_9453);
or U9562 (N_9562,N_9398,N_9490);
nor U9563 (N_9563,N_9436,N_9382);
or U9564 (N_9564,N_9421,N_9363);
or U9565 (N_9565,N_9342,N_9351);
or U9566 (N_9566,N_9399,N_9325);
nand U9567 (N_9567,N_9359,N_9362);
or U9568 (N_9568,N_9257,N_9389);
xor U9569 (N_9569,N_9278,N_9409);
nand U9570 (N_9570,N_9326,N_9419);
nand U9571 (N_9571,N_9321,N_9481);
and U9572 (N_9572,N_9472,N_9340);
xor U9573 (N_9573,N_9372,N_9251);
and U9574 (N_9574,N_9478,N_9348);
and U9575 (N_9575,N_9299,N_9447);
or U9576 (N_9576,N_9388,N_9346);
xor U9577 (N_9577,N_9307,N_9254);
xor U9578 (N_9578,N_9432,N_9417);
and U9579 (N_9579,N_9406,N_9446);
nor U9580 (N_9580,N_9485,N_9308);
nand U9581 (N_9581,N_9445,N_9468);
or U9582 (N_9582,N_9323,N_9423);
or U9583 (N_9583,N_9464,N_9493);
and U9584 (N_9584,N_9309,N_9343);
nor U9585 (N_9585,N_9301,N_9311);
or U9586 (N_9586,N_9458,N_9365);
xnor U9587 (N_9587,N_9467,N_9487);
and U9588 (N_9588,N_9412,N_9466);
xnor U9589 (N_9589,N_9479,N_9292);
xor U9590 (N_9590,N_9483,N_9279);
xnor U9591 (N_9591,N_9451,N_9425);
and U9592 (N_9592,N_9266,N_9295);
nor U9593 (N_9593,N_9494,N_9274);
and U9594 (N_9594,N_9498,N_9374);
nor U9595 (N_9595,N_9291,N_9470);
xnor U9596 (N_9596,N_9491,N_9310);
xnor U9597 (N_9597,N_9264,N_9331);
and U9598 (N_9598,N_9403,N_9448);
nand U9599 (N_9599,N_9258,N_9410);
and U9600 (N_9600,N_9298,N_9289);
or U9601 (N_9601,N_9454,N_9433);
or U9602 (N_9602,N_9395,N_9344);
xnor U9603 (N_9603,N_9356,N_9335);
nor U9604 (N_9604,N_9324,N_9405);
nand U9605 (N_9605,N_9452,N_9456);
nor U9606 (N_9606,N_9297,N_9430);
or U9607 (N_9607,N_9427,N_9387);
and U9608 (N_9608,N_9293,N_9480);
or U9609 (N_9609,N_9443,N_9360);
nor U9610 (N_9610,N_9450,N_9457);
or U9611 (N_9611,N_9315,N_9402);
or U9612 (N_9612,N_9440,N_9437);
xnor U9613 (N_9613,N_9253,N_9276);
or U9614 (N_9614,N_9318,N_9332);
or U9615 (N_9615,N_9373,N_9304);
xnor U9616 (N_9616,N_9353,N_9461);
nand U9617 (N_9617,N_9416,N_9475);
nor U9618 (N_9618,N_9287,N_9489);
nor U9619 (N_9619,N_9404,N_9327);
nor U9620 (N_9620,N_9428,N_9317);
and U9621 (N_9621,N_9424,N_9281);
nor U9622 (N_9622,N_9386,N_9422);
or U9623 (N_9623,N_9330,N_9465);
nand U9624 (N_9624,N_9380,N_9286);
nor U9625 (N_9625,N_9464,N_9424);
xor U9626 (N_9626,N_9285,N_9312);
nor U9627 (N_9627,N_9408,N_9353);
and U9628 (N_9628,N_9388,N_9455);
nand U9629 (N_9629,N_9431,N_9384);
nor U9630 (N_9630,N_9310,N_9480);
and U9631 (N_9631,N_9333,N_9311);
or U9632 (N_9632,N_9271,N_9453);
xnor U9633 (N_9633,N_9480,N_9485);
xnor U9634 (N_9634,N_9405,N_9374);
nor U9635 (N_9635,N_9365,N_9276);
or U9636 (N_9636,N_9490,N_9494);
or U9637 (N_9637,N_9266,N_9470);
and U9638 (N_9638,N_9426,N_9436);
nor U9639 (N_9639,N_9262,N_9261);
or U9640 (N_9640,N_9420,N_9411);
xor U9641 (N_9641,N_9478,N_9350);
nand U9642 (N_9642,N_9436,N_9434);
xnor U9643 (N_9643,N_9304,N_9390);
nand U9644 (N_9644,N_9467,N_9446);
xnor U9645 (N_9645,N_9271,N_9418);
and U9646 (N_9646,N_9294,N_9285);
nand U9647 (N_9647,N_9313,N_9364);
nor U9648 (N_9648,N_9254,N_9354);
or U9649 (N_9649,N_9356,N_9491);
xnor U9650 (N_9650,N_9377,N_9343);
xor U9651 (N_9651,N_9312,N_9304);
nor U9652 (N_9652,N_9325,N_9360);
xor U9653 (N_9653,N_9266,N_9280);
nand U9654 (N_9654,N_9286,N_9497);
xor U9655 (N_9655,N_9463,N_9423);
nand U9656 (N_9656,N_9309,N_9427);
nand U9657 (N_9657,N_9382,N_9317);
nor U9658 (N_9658,N_9253,N_9274);
xnor U9659 (N_9659,N_9463,N_9352);
nand U9660 (N_9660,N_9384,N_9401);
or U9661 (N_9661,N_9364,N_9263);
nand U9662 (N_9662,N_9252,N_9399);
nand U9663 (N_9663,N_9295,N_9404);
nand U9664 (N_9664,N_9443,N_9356);
nor U9665 (N_9665,N_9314,N_9299);
or U9666 (N_9666,N_9351,N_9472);
and U9667 (N_9667,N_9477,N_9418);
xor U9668 (N_9668,N_9497,N_9390);
and U9669 (N_9669,N_9370,N_9436);
and U9670 (N_9670,N_9347,N_9286);
and U9671 (N_9671,N_9297,N_9472);
nor U9672 (N_9672,N_9332,N_9290);
or U9673 (N_9673,N_9394,N_9450);
xnor U9674 (N_9674,N_9289,N_9352);
and U9675 (N_9675,N_9370,N_9379);
xor U9676 (N_9676,N_9268,N_9323);
nand U9677 (N_9677,N_9472,N_9312);
nor U9678 (N_9678,N_9398,N_9337);
nor U9679 (N_9679,N_9313,N_9373);
nand U9680 (N_9680,N_9372,N_9498);
and U9681 (N_9681,N_9308,N_9408);
nand U9682 (N_9682,N_9463,N_9479);
xnor U9683 (N_9683,N_9276,N_9264);
nand U9684 (N_9684,N_9388,N_9359);
nand U9685 (N_9685,N_9325,N_9354);
or U9686 (N_9686,N_9393,N_9405);
nor U9687 (N_9687,N_9478,N_9472);
xor U9688 (N_9688,N_9330,N_9414);
and U9689 (N_9689,N_9323,N_9452);
or U9690 (N_9690,N_9456,N_9359);
or U9691 (N_9691,N_9277,N_9294);
nor U9692 (N_9692,N_9489,N_9493);
nand U9693 (N_9693,N_9413,N_9483);
nor U9694 (N_9694,N_9318,N_9251);
nand U9695 (N_9695,N_9452,N_9354);
nand U9696 (N_9696,N_9489,N_9307);
and U9697 (N_9697,N_9351,N_9313);
and U9698 (N_9698,N_9409,N_9332);
and U9699 (N_9699,N_9272,N_9384);
xor U9700 (N_9700,N_9322,N_9304);
or U9701 (N_9701,N_9480,N_9257);
and U9702 (N_9702,N_9419,N_9356);
and U9703 (N_9703,N_9253,N_9387);
nand U9704 (N_9704,N_9451,N_9457);
nor U9705 (N_9705,N_9415,N_9272);
and U9706 (N_9706,N_9439,N_9292);
xnor U9707 (N_9707,N_9315,N_9354);
xnor U9708 (N_9708,N_9351,N_9362);
or U9709 (N_9709,N_9385,N_9277);
nor U9710 (N_9710,N_9337,N_9295);
and U9711 (N_9711,N_9345,N_9367);
or U9712 (N_9712,N_9295,N_9335);
nor U9713 (N_9713,N_9344,N_9460);
nand U9714 (N_9714,N_9281,N_9363);
and U9715 (N_9715,N_9309,N_9405);
xor U9716 (N_9716,N_9307,N_9267);
nor U9717 (N_9717,N_9462,N_9282);
or U9718 (N_9718,N_9326,N_9253);
or U9719 (N_9719,N_9347,N_9360);
and U9720 (N_9720,N_9357,N_9360);
nor U9721 (N_9721,N_9263,N_9491);
xnor U9722 (N_9722,N_9338,N_9415);
or U9723 (N_9723,N_9318,N_9421);
xor U9724 (N_9724,N_9370,N_9280);
nor U9725 (N_9725,N_9444,N_9376);
nand U9726 (N_9726,N_9320,N_9419);
nor U9727 (N_9727,N_9306,N_9254);
nand U9728 (N_9728,N_9314,N_9404);
nor U9729 (N_9729,N_9305,N_9296);
or U9730 (N_9730,N_9368,N_9446);
and U9731 (N_9731,N_9399,N_9290);
nand U9732 (N_9732,N_9411,N_9457);
xor U9733 (N_9733,N_9262,N_9321);
nand U9734 (N_9734,N_9303,N_9489);
nor U9735 (N_9735,N_9289,N_9369);
xnor U9736 (N_9736,N_9347,N_9350);
nor U9737 (N_9737,N_9290,N_9360);
or U9738 (N_9738,N_9331,N_9300);
nand U9739 (N_9739,N_9393,N_9492);
xor U9740 (N_9740,N_9476,N_9313);
and U9741 (N_9741,N_9466,N_9414);
or U9742 (N_9742,N_9371,N_9492);
and U9743 (N_9743,N_9415,N_9438);
nand U9744 (N_9744,N_9479,N_9324);
xnor U9745 (N_9745,N_9349,N_9467);
xnor U9746 (N_9746,N_9321,N_9390);
nand U9747 (N_9747,N_9262,N_9490);
nor U9748 (N_9748,N_9296,N_9270);
nand U9749 (N_9749,N_9281,N_9337);
nor U9750 (N_9750,N_9565,N_9606);
nand U9751 (N_9751,N_9641,N_9642);
xor U9752 (N_9752,N_9744,N_9590);
nor U9753 (N_9753,N_9734,N_9612);
and U9754 (N_9754,N_9598,N_9675);
nand U9755 (N_9755,N_9657,N_9634);
or U9756 (N_9756,N_9595,N_9672);
or U9757 (N_9757,N_9702,N_9738);
nand U9758 (N_9758,N_9706,N_9669);
nor U9759 (N_9759,N_9736,N_9639);
nand U9760 (N_9760,N_9503,N_9609);
or U9761 (N_9761,N_9514,N_9599);
nand U9762 (N_9762,N_9714,N_9589);
and U9763 (N_9763,N_9645,N_9695);
nor U9764 (N_9764,N_9660,N_9517);
and U9765 (N_9765,N_9532,N_9650);
and U9766 (N_9766,N_9741,N_9525);
xnor U9767 (N_9767,N_9518,N_9647);
nor U9768 (N_9768,N_9524,N_9501);
nor U9769 (N_9769,N_9577,N_9563);
and U9770 (N_9770,N_9731,N_9694);
xnor U9771 (N_9771,N_9547,N_9723);
and U9772 (N_9772,N_9516,N_9560);
or U9773 (N_9773,N_9586,N_9666);
nor U9774 (N_9774,N_9730,N_9504);
nand U9775 (N_9775,N_9570,N_9554);
xnor U9776 (N_9776,N_9604,N_9584);
xnor U9777 (N_9777,N_9626,N_9515);
and U9778 (N_9778,N_9637,N_9538);
or U9779 (N_9779,N_9636,N_9557);
or U9780 (N_9780,N_9581,N_9739);
xor U9781 (N_9781,N_9566,N_9594);
or U9782 (N_9782,N_9630,N_9659);
xnor U9783 (N_9783,N_9733,N_9740);
xnor U9784 (N_9784,N_9511,N_9726);
nor U9785 (N_9785,N_9638,N_9541);
and U9786 (N_9786,N_9673,N_9545);
nor U9787 (N_9787,N_9713,N_9686);
nand U9788 (N_9788,N_9572,N_9663);
nor U9789 (N_9789,N_9704,N_9749);
xor U9790 (N_9790,N_9664,N_9549);
nand U9791 (N_9791,N_9512,N_9725);
nor U9792 (N_9792,N_9658,N_9597);
or U9793 (N_9793,N_9519,N_9613);
nand U9794 (N_9794,N_9536,N_9632);
nand U9795 (N_9795,N_9717,N_9722);
or U9796 (N_9796,N_9593,N_9521);
or U9797 (N_9797,N_9601,N_9643);
nor U9798 (N_9798,N_9543,N_9729);
nor U9799 (N_9799,N_9537,N_9656);
nor U9800 (N_9800,N_9627,N_9746);
xnor U9801 (N_9801,N_9665,N_9710);
nand U9802 (N_9802,N_9558,N_9608);
nand U9803 (N_9803,N_9576,N_9569);
xnor U9804 (N_9804,N_9742,N_9587);
nor U9805 (N_9805,N_9678,N_9591);
nor U9806 (N_9806,N_9596,N_9644);
or U9807 (N_9807,N_9700,N_9534);
xnor U9808 (N_9808,N_9715,N_9683);
nor U9809 (N_9809,N_9564,N_9691);
xnor U9810 (N_9810,N_9507,N_9509);
and U9811 (N_9811,N_9625,N_9708);
nor U9812 (N_9812,N_9535,N_9531);
and U9813 (N_9813,N_9711,N_9703);
nor U9814 (N_9814,N_9724,N_9668);
and U9815 (N_9815,N_9667,N_9561);
or U9816 (N_9816,N_9677,N_9533);
and U9817 (N_9817,N_9611,N_9747);
or U9818 (N_9818,N_9548,N_9640);
nand U9819 (N_9819,N_9692,N_9559);
xnor U9820 (N_9820,N_9651,N_9629);
and U9821 (N_9821,N_9748,N_9633);
and U9822 (N_9822,N_9684,N_9567);
or U9823 (N_9823,N_9624,N_9552);
nand U9824 (N_9824,N_9701,N_9529);
nor U9825 (N_9825,N_9592,N_9648);
xor U9826 (N_9826,N_9690,N_9674);
or U9827 (N_9827,N_9614,N_9737);
nand U9828 (N_9828,N_9522,N_9520);
and U9829 (N_9829,N_9631,N_9681);
or U9830 (N_9830,N_9693,N_9688);
and U9831 (N_9831,N_9699,N_9680);
or U9832 (N_9832,N_9618,N_9732);
xnor U9833 (N_9833,N_9583,N_9513);
xor U9834 (N_9834,N_9575,N_9528);
or U9835 (N_9835,N_9628,N_9661);
xor U9836 (N_9836,N_9506,N_9696);
nand U9837 (N_9837,N_9670,N_9574);
and U9838 (N_9838,N_9743,N_9662);
or U9839 (N_9839,N_9600,N_9655);
or U9840 (N_9840,N_9556,N_9620);
or U9841 (N_9841,N_9588,N_9579);
xor U9842 (N_9842,N_9530,N_9526);
nor U9843 (N_9843,N_9709,N_9697);
xor U9844 (N_9844,N_9505,N_9735);
and U9845 (N_9845,N_9540,N_9653);
or U9846 (N_9846,N_9544,N_9510);
or U9847 (N_9847,N_9698,N_9500);
or U9848 (N_9848,N_9745,N_9502);
xor U9849 (N_9849,N_9687,N_9649);
and U9850 (N_9850,N_9602,N_9728);
nand U9851 (N_9851,N_9562,N_9635);
xnor U9852 (N_9852,N_9539,N_9721);
nor U9853 (N_9853,N_9623,N_9603);
or U9854 (N_9854,N_9542,N_9707);
or U9855 (N_9855,N_9585,N_9716);
nor U9856 (N_9856,N_9616,N_9568);
nor U9857 (N_9857,N_9573,N_9527);
or U9858 (N_9858,N_9550,N_9580);
or U9859 (N_9859,N_9508,N_9646);
and U9860 (N_9860,N_9619,N_9685);
xnor U9861 (N_9861,N_9727,N_9705);
or U9862 (N_9862,N_9546,N_9679);
xnor U9863 (N_9863,N_9671,N_9551);
and U9864 (N_9864,N_9523,N_9718);
or U9865 (N_9865,N_9553,N_9621);
nor U9866 (N_9866,N_9622,N_9607);
or U9867 (N_9867,N_9719,N_9676);
and U9868 (N_9868,N_9582,N_9615);
nand U9869 (N_9869,N_9605,N_9652);
or U9870 (N_9870,N_9720,N_9617);
xor U9871 (N_9871,N_9689,N_9682);
or U9872 (N_9872,N_9712,N_9654);
nand U9873 (N_9873,N_9571,N_9610);
or U9874 (N_9874,N_9578,N_9555);
nand U9875 (N_9875,N_9663,N_9716);
or U9876 (N_9876,N_9691,N_9628);
nand U9877 (N_9877,N_9722,N_9593);
nor U9878 (N_9878,N_9725,N_9672);
nand U9879 (N_9879,N_9634,N_9531);
nor U9880 (N_9880,N_9742,N_9589);
and U9881 (N_9881,N_9526,N_9699);
nand U9882 (N_9882,N_9562,N_9612);
nand U9883 (N_9883,N_9653,N_9538);
and U9884 (N_9884,N_9540,N_9611);
or U9885 (N_9885,N_9715,N_9599);
xnor U9886 (N_9886,N_9591,N_9551);
nor U9887 (N_9887,N_9680,N_9615);
and U9888 (N_9888,N_9649,N_9730);
or U9889 (N_9889,N_9728,N_9718);
nand U9890 (N_9890,N_9720,N_9706);
or U9891 (N_9891,N_9630,N_9530);
nor U9892 (N_9892,N_9650,N_9692);
xnor U9893 (N_9893,N_9545,N_9577);
or U9894 (N_9894,N_9659,N_9677);
nor U9895 (N_9895,N_9605,N_9626);
or U9896 (N_9896,N_9640,N_9735);
nand U9897 (N_9897,N_9623,N_9649);
and U9898 (N_9898,N_9672,N_9512);
xor U9899 (N_9899,N_9523,N_9704);
xor U9900 (N_9900,N_9533,N_9530);
xor U9901 (N_9901,N_9623,N_9733);
and U9902 (N_9902,N_9664,N_9721);
nor U9903 (N_9903,N_9557,N_9626);
and U9904 (N_9904,N_9547,N_9606);
nor U9905 (N_9905,N_9528,N_9539);
and U9906 (N_9906,N_9685,N_9726);
xor U9907 (N_9907,N_9686,N_9538);
xor U9908 (N_9908,N_9542,N_9730);
xor U9909 (N_9909,N_9561,N_9553);
and U9910 (N_9910,N_9510,N_9545);
nand U9911 (N_9911,N_9679,N_9644);
and U9912 (N_9912,N_9724,N_9567);
and U9913 (N_9913,N_9744,N_9594);
and U9914 (N_9914,N_9529,N_9706);
xnor U9915 (N_9915,N_9701,N_9532);
and U9916 (N_9916,N_9698,N_9667);
nand U9917 (N_9917,N_9618,N_9533);
xor U9918 (N_9918,N_9707,N_9747);
and U9919 (N_9919,N_9572,N_9527);
and U9920 (N_9920,N_9711,N_9673);
and U9921 (N_9921,N_9528,N_9521);
or U9922 (N_9922,N_9511,N_9533);
nor U9923 (N_9923,N_9705,N_9701);
or U9924 (N_9924,N_9668,N_9597);
and U9925 (N_9925,N_9547,N_9634);
and U9926 (N_9926,N_9620,N_9652);
or U9927 (N_9927,N_9686,N_9597);
or U9928 (N_9928,N_9747,N_9691);
or U9929 (N_9929,N_9622,N_9655);
nor U9930 (N_9930,N_9512,N_9611);
xor U9931 (N_9931,N_9652,N_9646);
xor U9932 (N_9932,N_9599,N_9521);
or U9933 (N_9933,N_9715,N_9711);
or U9934 (N_9934,N_9569,N_9541);
or U9935 (N_9935,N_9722,N_9521);
xor U9936 (N_9936,N_9531,N_9514);
or U9937 (N_9937,N_9586,N_9604);
nor U9938 (N_9938,N_9539,N_9730);
nand U9939 (N_9939,N_9726,N_9638);
or U9940 (N_9940,N_9550,N_9693);
xor U9941 (N_9941,N_9699,N_9698);
and U9942 (N_9942,N_9728,N_9639);
and U9943 (N_9943,N_9634,N_9694);
xor U9944 (N_9944,N_9620,N_9544);
and U9945 (N_9945,N_9644,N_9641);
or U9946 (N_9946,N_9659,N_9742);
or U9947 (N_9947,N_9534,N_9676);
nand U9948 (N_9948,N_9540,N_9620);
or U9949 (N_9949,N_9572,N_9724);
and U9950 (N_9950,N_9605,N_9723);
xnor U9951 (N_9951,N_9695,N_9519);
nand U9952 (N_9952,N_9607,N_9595);
xnor U9953 (N_9953,N_9695,N_9624);
nor U9954 (N_9954,N_9594,N_9608);
or U9955 (N_9955,N_9583,N_9528);
nor U9956 (N_9956,N_9585,N_9594);
xor U9957 (N_9957,N_9529,N_9667);
xnor U9958 (N_9958,N_9691,N_9511);
and U9959 (N_9959,N_9510,N_9709);
nand U9960 (N_9960,N_9675,N_9506);
and U9961 (N_9961,N_9690,N_9531);
or U9962 (N_9962,N_9735,N_9603);
nand U9963 (N_9963,N_9722,N_9590);
and U9964 (N_9964,N_9542,N_9719);
xor U9965 (N_9965,N_9736,N_9566);
xor U9966 (N_9966,N_9557,N_9573);
nand U9967 (N_9967,N_9530,N_9560);
xor U9968 (N_9968,N_9607,N_9570);
nand U9969 (N_9969,N_9633,N_9657);
nand U9970 (N_9970,N_9620,N_9619);
nor U9971 (N_9971,N_9682,N_9687);
nor U9972 (N_9972,N_9550,N_9675);
and U9973 (N_9973,N_9642,N_9538);
or U9974 (N_9974,N_9645,N_9574);
xor U9975 (N_9975,N_9649,N_9545);
nand U9976 (N_9976,N_9544,N_9524);
nor U9977 (N_9977,N_9557,N_9628);
and U9978 (N_9978,N_9639,N_9542);
nand U9979 (N_9979,N_9541,N_9667);
nor U9980 (N_9980,N_9666,N_9676);
nor U9981 (N_9981,N_9513,N_9672);
nor U9982 (N_9982,N_9550,N_9508);
or U9983 (N_9983,N_9578,N_9579);
or U9984 (N_9984,N_9681,N_9669);
xor U9985 (N_9985,N_9652,N_9564);
nand U9986 (N_9986,N_9602,N_9514);
xor U9987 (N_9987,N_9718,N_9668);
xnor U9988 (N_9988,N_9713,N_9605);
nand U9989 (N_9989,N_9524,N_9674);
xnor U9990 (N_9990,N_9527,N_9721);
nor U9991 (N_9991,N_9611,N_9690);
or U9992 (N_9992,N_9679,N_9639);
nand U9993 (N_9993,N_9681,N_9593);
nand U9994 (N_9994,N_9579,N_9642);
and U9995 (N_9995,N_9591,N_9514);
nor U9996 (N_9996,N_9548,N_9526);
and U9997 (N_9997,N_9721,N_9585);
xnor U9998 (N_9998,N_9637,N_9547);
and U9999 (N_9999,N_9716,N_9741);
nand U10000 (N_10000,N_9883,N_9987);
nand U10001 (N_10001,N_9807,N_9887);
and U10002 (N_10002,N_9834,N_9928);
or U10003 (N_10003,N_9878,N_9773);
nand U10004 (N_10004,N_9752,N_9828);
nand U10005 (N_10005,N_9798,N_9952);
nand U10006 (N_10006,N_9983,N_9939);
or U10007 (N_10007,N_9940,N_9758);
and U10008 (N_10008,N_9818,N_9995);
or U10009 (N_10009,N_9962,N_9930);
xnor U10010 (N_10010,N_9801,N_9862);
and U10011 (N_10011,N_9922,N_9902);
nand U10012 (N_10012,N_9994,N_9757);
nand U10013 (N_10013,N_9786,N_9869);
nor U10014 (N_10014,N_9776,N_9965);
xnor U10015 (N_10015,N_9949,N_9796);
nand U10016 (N_10016,N_9899,N_9825);
nor U10017 (N_10017,N_9919,N_9882);
or U10018 (N_10018,N_9859,N_9893);
xnor U10019 (N_10019,N_9783,N_9840);
and U10020 (N_10020,N_9836,N_9992);
nor U10021 (N_10021,N_9875,N_9936);
xor U10022 (N_10022,N_9872,N_9830);
and U10023 (N_10023,N_9966,N_9866);
and U10024 (N_10024,N_9898,N_9890);
nand U10025 (N_10025,N_9993,N_9754);
nor U10026 (N_10026,N_9946,N_9876);
xor U10027 (N_10027,N_9802,N_9809);
nor U10028 (N_10028,N_9756,N_9907);
nand U10029 (N_10029,N_9920,N_9864);
xnor U10030 (N_10030,N_9774,N_9751);
and U10031 (N_10031,N_9850,N_9944);
xnor U10032 (N_10032,N_9925,N_9941);
and U10033 (N_10033,N_9951,N_9981);
and U10034 (N_10034,N_9874,N_9979);
and U10035 (N_10035,N_9942,N_9811);
or U10036 (N_10036,N_9963,N_9891);
nand U10037 (N_10037,N_9770,N_9917);
nand U10038 (N_10038,N_9845,N_9842);
and U10039 (N_10039,N_9915,N_9847);
nor U10040 (N_10040,N_9817,N_9999);
nand U10041 (N_10041,N_9892,N_9932);
and U10042 (N_10042,N_9856,N_9781);
xor U10043 (N_10043,N_9977,N_9950);
and U10044 (N_10044,N_9797,N_9903);
xnor U10045 (N_10045,N_9775,N_9894);
and U10046 (N_10046,N_9832,N_9820);
xnor U10047 (N_10047,N_9986,N_9881);
or U10048 (N_10048,N_9923,N_9769);
nor U10049 (N_10049,N_9823,N_9763);
nand U10050 (N_10050,N_9918,N_9897);
and U10051 (N_10051,N_9810,N_9961);
or U10052 (N_10052,N_9762,N_9974);
nand U10053 (N_10053,N_9867,N_9889);
or U10054 (N_10054,N_9985,N_9844);
xor U10055 (N_10055,N_9997,N_9848);
and U10056 (N_10056,N_9764,N_9831);
xnor U10057 (N_10057,N_9771,N_9821);
nor U10058 (N_10058,N_9849,N_9795);
xnor U10059 (N_10059,N_9971,N_9901);
nand U10060 (N_10060,N_9860,N_9793);
nor U10061 (N_10061,N_9970,N_9865);
nor U10062 (N_10062,N_9838,N_9779);
and U10063 (N_10063,N_9826,N_9855);
nand U10064 (N_10064,N_9908,N_9800);
or U10065 (N_10065,N_9753,N_9822);
xor U10066 (N_10066,N_9768,N_9964);
xnor U10067 (N_10067,N_9789,N_9976);
or U10068 (N_10068,N_9996,N_9759);
xor U10069 (N_10069,N_9955,N_9824);
and U10070 (N_10070,N_9788,N_9905);
nand U10071 (N_10071,N_9837,N_9861);
nand U10072 (N_10072,N_9948,N_9792);
or U10073 (N_10073,N_9814,N_9806);
nor U10074 (N_10074,N_9868,N_9841);
and U10075 (N_10075,N_9765,N_9808);
nor U10076 (N_10076,N_9953,N_9787);
xor U10077 (N_10077,N_9880,N_9960);
or U10078 (N_10078,N_9988,N_9959);
or U10079 (N_10079,N_9895,N_9916);
xor U10080 (N_10080,N_9816,N_9854);
nand U10081 (N_10081,N_9835,N_9921);
nand U10082 (N_10082,N_9782,N_9982);
or U10083 (N_10083,N_9791,N_9934);
nor U10084 (N_10084,N_9896,N_9794);
xor U10085 (N_10085,N_9761,N_9888);
and U10086 (N_10086,N_9913,N_9829);
xnor U10087 (N_10087,N_9935,N_9760);
xor U10088 (N_10088,N_9772,N_9805);
or U10089 (N_10089,N_9975,N_9978);
and U10090 (N_10090,N_9937,N_9857);
nand U10091 (N_10091,N_9815,N_9813);
nand U10092 (N_10092,N_9900,N_9873);
or U10093 (N_10093,N_9968,N_9933);
nor U10094 (N_10094,N_9885,N_9750);
nor U10095 (N_10095,N_9780,N_9973);
nor U10096 (N_10096,N_9767,N_9906);
or U10097 (N_10097,N_9804,N_9927);
and U10098 (N_10098,N_9909,N_9863);
xor U10099 (N_10099,N_9910,N_9991);
xnor U10100 (N_10100,N_9755,N_9998);
nand U10101 (N_10101,N_9877,N_9943);
and U10102 (N_10102,N_9957,N_9871);
and U10103 (N_10103,N_9777,N_9853);
nor U10104 (N_10104,N_9969,N_9839);
and U10105 (N_10105,N_9947,N_9954);
nand U10106 (N_10106,N_9972,N_9967);
nor U10107 (N_10107,N_9980,N_9904);
and U10108 (N_10108,N_9912,N_9884);
or U10109 (N_10109,N_9803,N_9812);
nand U10110 (N_10110,N_9851,N_9956);
and U10111 (N_10111,N_9945,N_9984);
nor U10112 (N_10112,N_9785,N_9858);
or U10113 (N_10113,N_9852,N_9886);
xnor U10114 (N_10114,N_9958,N_9931);
nor U10115 (N_10115,N_9870,N_9827);
xnor U10116 (N_10116,N_9784,N_9833);
or U10117 (N_10117,N_9926,N_9843);
xor U10118 (N_10118,N_9846,N_9914);
and U10119 (N_10119,N_9938,N_9778);
nor U10120 (N_10120,N_9766,N_9799);
xor U10121 (N_10121,N_9990,N_9924);
and U10122 (N_10122,N_9819,N_9911);
or U10123 (N_10123,N_9989,N_9790);
nor U10124 (N_10124,N_9879,N_9929);
nor U10125 (N_10125,N_9867,N_9811);
nand U10126 (N_10126,N_9988,N_9907);
nand U10127 (N_10127,N_9802,N_9835);
and U10128 (N_10128,N_9761,N_9818);
nand U10129 (N_10129,N_9759,N_9921);
or U10130 (N_10130,N_9775,N_9922);
and U10131 (N_10131,N_9959,N_9981);
nand U10132 (N_10132,N_9775,N_9779);
xor U10133 (N_10133,N_9960,N_9819);
or U10134 (N_10134,N_9932,N_9900);
xor U10135 (N_10135,N_9927,N_9781);
and U10136 (N_10136,N_9897,N_9931);
nor U10137 (N_10137,N_9908,N_9927);
or U10138 (N_10138,N_9959,N_9754);
xnor U10139 (N_10139,N_9824,N_9848);
nand U10140 (N_10140,N_9942,N_9945);
nor U10141 (N_10141,N_9870,N_9848);
or U10142 (N_10142,N_9796,N_9843);
and U10143 (N_10143,N_9778,N_9828);
nand U10144 (N_10144,N_9916,N_9993);
nand U10145 (N_10145,N_9934,N_9870);
nor U10146 (N_10146,N_9806,N_9970);
and U10147 (N_10147,N_9841,N_9857);
xnor U10148 (N_10148,N_9858,N_9841);
nand U10149 (N_10149,N_9897,N_9895);
and U10150 (N_10150,N_9816,N_9889);
nor U10151 (N_10151,N_9868,N_9850);
nand U10152 (N_10152,N_9822,N_9838);
xor U10153 (N_10153,N_9841,N_9862);
xor U10154 (N_10154,N_9877,N_9981);
nand U10155 (N_10155,N_9985,N_9945);
or U10156 (N_10156,N_9932,N_9991);
or U10157 (N_10157,N_9792,N_9852);
or U10158 (N_10158,N_9951,N_9856);
nor U10159 (N_10159,N_9853,N_9752);
and U10160 (N_10160,N_9978,N_9797);
nor U10161 (N_10161,N_9919,N_9872);
nor U10162 (N_10162,N_9790,N_9938);
nor U10163 (N_10163,N_9952,N_9860);
nor U10164 (N_10164,N_9940,N_9952);
nor U10165 (N_10165,N_9862,N_9931);
nor U10166 (N_10166,N_9841,N_9780);
xnor U10167 (N_10167,N_9955,N_9796);
nand U10168 (N_10168,N_9946,N_9752);
or U10169 (N_10169,N_9961,N_9830);
and U10170 (N_10170,N_9903,N_9832);
and U10171 (N_10171,N_9902,N_9824);
nor U10172 (N_10172,N_9995,N_9923);
or U10173 (N_10173,N_9979,N_9784);
and U10174 (N_10174,N_9887,N_9773);
or U10175 (N_10175,N_9850,N_9884);
xnor U10176 (N_10176,N_9913,N_9891);
nor U10177 (N_10177,N_9954,N_9752);
and U10178 (N_10178,N_9924,N_9813);
nor U10179 (N_10179,N_9977,N_9767);
xnor U10180 (N_10180,N_9875,N_9871);
or U10181 (N_10181,N_9803,N_9920);
xnor U10182 (N_10182,N_9920,N_9794);
and U10183 (N_10183,N_9892,N_9816);
or U10184 (N_10184,N_9830,N_9809);
or U10185 (N_10185,N_9815,N_9857);
nand U10186 (N_10186,N_9998,N_9821);
and U10187 (N_10187,N_9974,N_9910);
and U10188 (N_10188,N_9994,N_9797);
and U10189 (N_10189,N_9759,N_9997);
and U10190 (N_10190,N_9895,N_9872);
or U10191 (N_10191,N_9960,N_9810);
xor U10192 (N_10192,N_9812,N_9864);
nor U10193 (N_10193,N_9817,N_9950);
and U10194 (N_10194,N_9840,N_9797);
and U10195 (N_10195,N_9892,N_9802);
and U10196 (N_10196,N_9769,N_9996);
or U10197 (N_10197,N_9842,N_9756);
xnor U10198 (N_10198,N_9880,N_9975);
xnor U10199 (N_10199,N_9936,N_9993);
nor U10200 (N_10200,N_9871,N_9905);
nor U10201 (N_10201,N_9901,N_9773);
nor U10202 (N_10202,N_9963,N_9932);
xnor U10203 (N_10203,N_9814,N_9992);
nand U10204 (N_10204,N_9944,N_9881);
nor U10205 (N_10205,N_9823,N_9919);
or U10206 (N_10206,N_9797,N_9839);
or U10207 (N_10207,N_9921,N_9963);
nor U10208 (N_10208,N_9770,N_9759);
or U10209 (N_10209,N_9787,N_9802);
and U10210 (N_10210,N_9916,N_9927);
xnor U10211 (N_10211,N_9766,N_9932);
nand U10212 (N_10212,N_9947,N_9851);
and U10213 (N_10213,N_9978,N_9992);
nand U10214 (N_10214,N_9815,N_9780);
nor U10215 (N_10215,N_9754,N_9881);
or U10216 (N_10216,N_9953,N_9859);
nor U10217 (N_10217,N_9757,N_9936);
or U10218 (N_10218,N_9851,N_9777);
or U10219 (N_10219,N_9756,N_9783);
nor U10220 (N_10220,N_9791,N_9976);
nand U10221 (N_10221,N_9914,N_9783);
nand U10222 (N_10222,N_9969,N_9840);
nand U10223 (N_10223,N_9930,N_9942);
or U10224 (N_10224,N_9974,N_9961);
or U10225 (N_10225,N_9921,N_9788);
xor U10226 (N_10226,N_9751,N_9794);
nor U10227 (N_10227,N_9819,N_9902);
nor U10228 (N_10228,N_9958,N_9762);
xnor U10229 (N_10229,N_9755,N_9888);
and U10230 (N_10230,N_9777,N_9824);
and U10231 (N_10231,N_9905,N_9887);
nand U10232 (N_10232,N_9756,N_9990);
nand U10233 (N_10233,N_9792,N_9945);
xor U10234 (N_10234,N_9763,N_9753);
and U10235 (N_10235,N_9952,N_9814);
and U10236 (N_10236,N_9956,N_9904);
nor U10237 (N_10237,N_9939,N_9978);
and U10238 (N_10238,N_9904,N_9803);
or U10239 (N_10239,N_9770,N_9890);
nand U10240 (N_10240,N_9794,N_9836);
nor U10241 (N_10241,N_9903,N_9764);
nand U10242 (N_10242,N_9784,N_9969);
xor U10243 (N_10243,N_9953,N_9822);
and U10244 (N_10244,N_9808,N_9754);
and U10245 (N_10245,N_9945,N_9857);
and U10246 (N_10246,N_9968,N_9884);
xnor U10247 (N_10247,N_9751,N_9812);
nand U10248 (N_10248,N_9898,N_9919);
nand U10249 (N_10249,N_9968,N_9975);
or U10250 (N_10250,N_10031,N_10238);
and U10251 (N_10251,N_10036,N_10218);
nand U10252 (N_10252,N_10005,N_10090);
nor U10253 (N_10253,N_10185,N_10158);
xor U10254 (N_10254,N_10242,N_10084);
xor U10255 (N_10255,N_10108,N_10067);
and U10256 (N_10256,N_10065,N_10081);
nor U10257 (N_10257,N_10012,N_10190);
or U10258 (N_10258,N_10011,N_10162);
and U10259 (N_10259,N_10069,N_10038);
and U10260 (N_10260,N_10114,N_10153);
nand U10261 (N_10261,N_10040,N_10004);
or U10262 (N_10262,N_10023,N_10175);
or U10263 (N_10263,N_10187,N_10174);
nand U10264 (N_10264,N_10091,N_10182);
nor U10265 (N_10265,N_10127,N_10247);
xnor U10266 (N_10266,N_10056,N_10053);
xnor U10267 (N_10267,N_10100,N_10070);
xor U10268 (N_10268,N_10024,N_10246);
nor U10269 (N_10269,N_10019,N_10121);
and U10270 (N_10270,N_10200,N_10214);
or U10271 (N_10271,N_10155,N_10112);
xor U10272 (N_10272,N_10119,N_10229);
nor U10273 (N_10273,N_10022,N_10054);
nand U10274 (N_10274,N_10248,N_10183);
or U10275 (N_10275,N_10195,N_10220);
or U10276 (N_10276,N_10046,N_10064);
or U10277 (N_10277,N_10192,N_10222);
xnor U10278 (N_10278,N_10223,N_10126);
nor U10279 (N_10279,N_10008,N_10191);
nor U10280 (N_10280,N_10082,N_10140);
nand U10281 (N_10281,N_10129,N_10102);
or U10282 (N_10282,N_10093,N_10203);
nor U10283 (N_10283,N_10186,N_10132);
nor U10284 (N_10284,N_10213,N_10156);
nor U10285 (N_10285,N_10124,N_10197);
and U10286 (N_10286,N_10166,N_10151);
nor U10287 (N_10287,N_10060,N_10078);
and U10288 (N_10288,N_10225,N_10131);
and U10289 (N_10289,N_10048,N_10017);
nor U10290 (N_10290,N_10176,N_10167);
and U10291 (N_10291,N_10179,N_10116);
nand U10292 (N_10292,N_10075,N_10105);
nand U10293 (N_10293,N_10111,N_10142);
and U10294 (N_10294,N_10130,N_10122);
nand U10295 (N_10295,N_10106,N_10107);
and U10296 (N_10296,N_10210,N_10049);
nand U10297 (N_10297,N_10224,N_10184);
and U10298 (N_10298,N_10208,N_10232);
and U10299 (N_10299,N_10094,N_10120);
xor U10300 (N_10300,N_10128,N_10103);
xnor U10301 (N_10301,N_10139,N_10165);
nor U10302 (N_10302,N_10086,N_10228);
and U10303 (N_10303,N_10180,N_10085);
nor U10304 (N_10304,N_10144,N_10079);
or U10305 (N_10305,N_10147,N_10217);
nand U10306 (N_10306,N_10115,N_10039);
xor U10307 (N_10307,N_10006,N_10020);
nand U10308 (N_10308,N_10194,N_10138);
and U10309 (N_10309,N_10073,N_10101);
xnor U10310 (N_10310,N_10014,N_10193);
or U10311 (N_10311,N_10118,N_10087);
and U10312 (N_10312,N_10041,N_10146);
and U10313 (N_10313,N_10010,N_10149);
xor U10314 (N_10314,N_10161,N_10168);
nor U10315 (N_10315,N_10009,N_10234);
or U10316 (N_10316,N_10032,N_10050);
nor U10317 (N_10317,N_10063,N_10237);
nor U10318 (N_10318,N_10033,N_10235);
and U10319 (N_10319,N_10042,N_10123);
nor U10320 (N_10320,N_10002,N_10001);
xor U10321 (N_10321,N_10052,N_10216);
and U10322 (N_10322,N_10212,N_10249);
or U10323 (N_10323,N_10134,N_10071);
and U10324 (N_10324,N_10034,N_10072);
nand U10325 (N_10325,N_10000,N_10177);
or U10326 (N_10326,N_10205,N_10241);
xor U10327 (N_10327,N_10169,N_10188);
or U10328 (N_10328,N_10150,N_10037);
nor U10329 (N_10329,N_10051,N_10154);
and U10330 (N_10330,N_10021,N_10136);
nand U10331 (N_10331,N_10089,N_10148);
and U10332 (N_10332,N_10074,N_10080);
nand U10333 (N_10333,N_10025,N_10061);
nand U10334 (N_10334,N_10178,N_10152);
xor U10335 (N_10335,N_10230,N_10059);
or U10336 (N_10336,N_10239,N_10233);
nand U10337 (N_10337,N_10215,N_10104);
nand U10338 (N_10338,N_10027,N_10245);
nor U10339 (N_10339,N_10170,N_10219);
nand U10340 (N_10340,N_10207,N_10141);
xnor U10341 (N_10341,N_10029,N_10206);
or U10342 (N_10342,N_10173,N_10083);
nand U10343 (N_10343,N_10226,N_10244);
and U10344 (N_10344,N_10135,N_10198);
nor U10345 (N_10345,N_10055,N_10015);
and U10346 (N_10346,N_10202,N_10236);
nand U10347 (N_10347,N_10204,N_10221);
or U10348 (N_10348,N_10013,N_10227);
xnor U10349 (N_10349,N_10243,N_10189);
nand U10350 (N_10350,N_10095,N_10076);
or U10351 (N_10351,N_10099,N_10018);
xor U10352 (N_10352,N_10181,N_10109);
nor U10353 (N_10353,N_10199,N_10163);
and U10354 (N_10354,N_10211,N_10047);
or U10355 (N_10355,N_10231,N_10117);
or U10356 (N_10356,N_10172,N_10030);
and U10357 (N_10357,N_10159,N_10137);
xor U10358 (N_10358,N_10016,N_10145);
nand U10359 (N_10359,N_10133,N_10043);
nand U10360 (N_10360,N_10077,N_10201);
nor U10361 (N_10361,N_10057,N_10164);
xor U10362 (N_10362,N_10171,N_10098);
and U10363 (N_10363,N_10125,N_10110);
or U10364 (N_10364,N_10058,N_10160);
nand U10365 (N_10365,N_10143,N_10196);
nand U10366 (N_10366,N_10066,N_10209);
or U10367 (N_10367,N_10028,N_10007);
or U10368 (N_10368,N_10062,N_10044);
xor U10369 (N_10369,N_10035,N_10240);
nor U10370 (N_10370,N_10157,N_10003);
nor U10371 (N_10371,N_10113,N_10096);
nor U10372 (N_10372,N_10068,N_10045);
or U10373 (N_10373,N_10026,N_10088);
and U10374 (N_10374,N_10092,N_10097);
and U10375 (N_10375,N_10090,N_10043);
xor U10376 (N_10376,N_10031,N_10145);
and U10377 (N_10377,N_10228,N_10248);
xor U10378 (N_10378,N_10017,N_10161);
nand U10379 (N_10379,N_10104,N_10098);
nor U10380 (N_10380,N_10131,N_10182);
nor U10381 (N_10381,N_10207,N_10093);
xnor U10382 (N_10382,N_10180,N_10146);
nor U10383 (N_10383,N_10217,N_10213);
and U10384 (N_10384,N_10220,N_10223);
nand U10385 (N_10385,N_10128,N_10139);
and U10386 (N_10386,N_10216,N_10206);
or U10387 (N_10387,N_10050,N_10192);
and U10388 (N_10388,N_10095,N_10077);
xnor U10389 (N_10389,N_10173,N_10000);
or U10390 (N_10390,N_10054,N_10084);
xor U10391 (N_10391,N_10112,N_10015);
xor U10392 (N_10392,N_10197,N_10109);
nor U10393 (N_10393,N_10166,N_10028);
nor U10394 (N_10394,N_10243,N_10131);
nand U10395 (N_10395,N_10143,N_10016);
and U10396 (N_10396,N_10116,N_10238);
nand U10397 (N_10397,N_10143,N_10078);
nand U10398 (N_10398,N_10187,N_10242);
and U10399 (N_10399,N_10055,N_10091);
or U10400 (N_10400,N_10101,N_10214);
xnor U10401 (N_10401,N_10128,N_10037);
nor U10402 (N_10402,N_10167,N_10126);
and U10403 (N_10403,N_10025,N_10152);
xnor U10404 (N_10404,N_10096,N_10040);
xor U10405 (N_10405,N_10151,N_10206);
nand U10406 (N_10406,N_10053,N_10130);
nor U10407 (N_10407,N_10005,N_10164);
or U10408 (N_10408,N_10071,N_10060);
nor U10409 (N_10409,N_10140,N_10229);
nand U10410 (N_10410,N_10154,N_10140);
nand U10411 (N_10411,N_10111,N_10103);
and U10412 (N_10412,N_10156,N_10011);
xnor U10413 (N_10413,N_10209,N_10056);
and U10414 (N_10414,N_10071,N_10084);
and U10415 (N_10415,N_10107,N_10108);
xor U10416 (N_10416,N_10013,N_10138);
nor U10417 (N_10417,N_10067,N_10090);
and U10418 (N_10418,N_10225,N_10065);
xnor U10419 (N_10419,N_10057,N_10128);
xnor U10420 (N_10420,N_10188,N_10092);
and U10421 (N_10421,N_10049,N_10146);
nand U10422 (N_10422,N_10024,N_10191);
and U10423 (N_10423,N_10022,N_10030);
nand U10424 (N_10424,N_10011,N_10212);
nand U10425 (N_10425,N_10185,N_10071);
nand U10426 (N_10426,N_10240,N_10180);
nand U10427 (N_10427,N_10249,N_10071);
nor U10428 (N_10428,N_10011,N_10207);
nand U10429 (N_10429,N_10245,N_10185);
or U10430 (N_10430,N_10161,N_10203);
nor U10431 (N_10431,N_10014,N_10159);
and U10432 (N_10432,N_10094,N_10132);
or U10433 (N_10433,N_10199,N_10070);
nand U10434 (N_10434,N_10032,N_10026);
xnor U10435 (N_10435,N_10242,N_10189);
and U10436 (N_10436,N_10127,N_10089);
and U10437 (N_10437,N_10227,N_10142);
xor U10438 (N_10438,N_10061,N_10173);
nand U10439 (N_10439,N_10094,N_10143);
or U10440 (N_10440,N_10145,N_10132);
xor U10441 (N_10441,N_10063,N_10164);
nor U10442 (N_10442,N_10185,N_10020);
nand U10443 (N_10443,N_10230,N_10030);
and U10444 (N_10444,N_10088,N_10247);
nand U10445 (N_10445,N_10103,N_10245);
nor U10446 (N_10446,N_10050,N_10179);
xor U10447 (N_10447,N_10173,N_10228);
xor U10448 (N_10448,N_10157,N_10005);
and U10449 (N_10449,N_10104,N_10195);
and U10450 (N_10450,N_10034,N_10187);
nand U10451 (N_10451,N_10085,N_10218);
or U10452 (N_10452,N_10078,N_10184);
nand U10453 (N_10453,N_10190,N_10166);
nand U10454 (N_10454,N_10117,N_10018);
nand U10455 (N_10455,N_10103,N_10059);
xor U10456 (N_10456,N_10123,N_10097);
nor U10457 (N_10457,N_10240,N_10011);
nand U10458 (N_10458,N_10145,N_10160);
nor U10459 (N_10459,N_10140,N_10022);
nand U10460 (N_10460,N_10052,N_10055);
and U10461 (N_10461,N_10062,N_10158);
nor U10462 (N_10462,N_10084,N_10137);
and U10463 (N_10463,N_10009,N_10069);
nor U10464 (N_10464,N_10085,N_10151);
nor U10465 (N_10465,N_10142,N_10017);
nand U10466 (N_10466,N_10220,N_10023);
and U10467 (N_10467,N_10221,N_10105);
nor U10468 (N_10468,N_10221,N_10095);
nor U10469 (N_10469,N_10103,N_10104);
nor U10470 (N_10470,N_10067,N_10017);
xnor U10471 (N_10471,N_10018,N_10132);
nand U10472 (N_10472,N_10186,N_10100);
nand U10473 (N_10473,N_10126,N_10114);
xnor U10474 (N_10474,N_10198,N_10160);
or U10475 (N_10475,N_10031,N_10067);
nand U10476 (N_10476,N_10214,N_10135);
xor U10477 (N_10477,N_10186,N_10181);
or U10478 (N_10478,N_10021,N_10154);
nor U10479 (N_10479,N_10084,N_10231);
or U10480 (N_10480,N_10131,N_10244);
xnor U10481 (N_10481,N_10201,N_10058);
nor U10482 (N_10482,N_10021,N_10083);
nand U10483 (N_10483,N_10249,N_10055);
or U10484 (N_10484,N_10016,N_10243);
and U10485 (N_10485,N_10113,N_10183);
xor U10486 (N_10486,N_10104,N_10173);
nor U10487 (N_10487,N_10113,N_10195);
or U10488 (N_10488,N_10016,N_10052);
nor U10489 (N_10489,N_10149,N_10001);
and U10490 (N_10490,N_10141,N_10219);
and U10491 (N_10491,N_10047,N_10159);
xor U10492 (N_10492,N_10047,N_10223);
and U10493 (N_10493,N_10222,N_10046);
or U10494 (N_10494,N_10075,N_10141);
nor U10495 (N_10495,N_10118,N_10224);
nand U10496 (N_10496,N_10001,N_10236);
xnor U10497 (N_10497,N_10183,N_10047);
xnor U10498 (N_10498,N_10178,N_10093);
nand U10499 (N_10499,N_10167,N_10188);
nor U10500 (N_10500,N_10389,N_10313);
or U10501 (N_10501,N_10476,N_10408);
or U10502 (N_10502,N_10457,N_10287);
and U10503 (N_10503,N_10473,N_10449);
xnor U10504 (N_10504,N_10467,N_10442);
or U10505 (N_10505,N_10370,N_10355);
nand U10506 (N_10506,N_10298,N_10263);
nand U10507 (N_10507,N_10391,N_10266);
nor U10508 (N_10508,N_10260,N_10361);
nor U10509 (N_10509,N_10375,N_10279);
xnor U10510 (N_10510,N_10397,N_10407);
nor U10511 (N_10511,N_10431,N_10258);
and U10512 (N_10512,N_10265,N_10455);
nor U10513 (N_10513,N_10338,N_10403);
xor U10514 (N_10514,N_10489,N_10444);
nand U10515 (N_10515,N_10435,N_10418);
nor U10516 (N_10516,N_10339,N_10477);
and U10517 (N_10517,N_10302,N_10463);
nand U10518 (N_10518,N_10280,N_10417);
and U10519 (N_10519,N_10494,N_10464);
xor U10520 (N_10520,N_10354,N_10255);
and U10521 (N_10521,N_10459,N_10433);
or U10522 (N_10522,N_10336,N_10323);
nand U10523 (N_10523,N_10469,N_10289);
xor U10524 (N_10524,N_10350,N_10496);
or U10525 (N_10525,N_10380,N_10286);
nand U10526 (N_10526,N_10371,N_10458);
xnor U10527 (N_10527,N_10275,N_10365);
or U10528 (N_10528,N_10471,N_10429);
or U10529 (N_10529,N_10267,N_10337);
and U10530 (N_10530,N_10251,N_10368);
nor U10531 (N_10531,N_10297,N_10330);
nor U10532 (N_10532,N_10383,N_10493);
nand U10533 (N_10533,N_10411,N_10331);
xor U10534 (N_10534,N_10474,N_10293);
and U10535 (N_10535,N_10386,N_10405);
xor U10536 (N_10536,N_10490,N_10396);
and U10537 (N_10537,N_10308,N_10475);
nand U10538 (N_10538,N_10443,N_10281);
nor U10539 (N_10539,N_10438,N_10273);
xnor U10540 (N_10540,N_10349,N_10398);
and U10541 (N_10541,N_10470,N_10420);
nor U10542 (N_10542,N_10479,N_10432);
or U10543 (N_10543,N_10421,N_10282);
nand U10544 (N_10544,N_10310,N_10283);
nand U10545 (N_10545,N_10482,N_10448);
nand U10546 (N_10546,N_10326,N_10352);
or U10547 (N_10547,N_10402,N_10440);
and U10548 (N_10548,N_10484,N_10300);
or U10549 (N_10549,N_10285,N_10306);
nand U10550 (N_10550,N_10364,N_10445);
xor U10551 (N_10551,N_10462,N_10343);
nor U10552 (N_10552,N_10325,N_10413);
nand U10553 (N_10553,N_10498,N_10393);
nor U10554 (N_10554,N_10276,N_10357);
or U10555 (N_10555,N_10264,N_10478);
and U10556 (N_10556,N_10495,N_10472);
xor U10557 (N_10557,N_10390,N_10384);
xor U10558 (N_10558,N_10404,N_10394);
and U10559 (N_10559,N_10410,N_10299);
nor U10560 (N_10560,N_10372,N_10346);
nand U10561 (N_10561,N_10342,N_10486);
nand U10562 (N_10562,N_10428,N_10288);
nand U10563 (N_10563,N_10454,N_10378);
and U10564 (N_10564,N_10318,N_10284);
nand U10565 (N_10565,N_10274,N_10292);
xor U10566 (N_10566,N_10452,N_10319);
and U10567 (N_10567,N_10460,N_10328);
xor U10568 (N_10568,N_10422,N_10291);
and U10569 (N_10569,N_10304,N_10252);
nor U10570 (N_10570,N_10480,N_10362);
nor U10571 (N_10571,N_10468,N_10340);
nand U10572 (N_10572,N_10409,N_10345);
nor U10573 (N_10573,N_10447,N_10312);
and U10574 (N_10574,N_10307,N_10415);
xnor U10575 (N_10575,N_10359,N_10363);
nor U10576 (N_10576,N_10314,N_10395);
xor U10577 (N_10577,N_10483,N_10257);
nor U10578 (N_10578,N_10385,N_10436);
xor U10579 (N_10579,N_10256,N_10412);
nand U10580 (N_10580,N_10369,N_10382);
or U10581 (N_10581,N_10253,N_10358);
xnor U10582 (N_10582,N_10466,N_10488);
nand U10583 (N_10583,N_10269,N_10262);
xor U10584 (N_10584,N_10261,N_10491);
nor U10585 (N_10585,N_10430,N_10414);
nor U10586 (N_10586,N_10426,N_10465);
or U10587 (N_10587,N_10450,N_10499);
nor U10588 (N_10588,N_10356,N_10254);
and U10589 (N_10589,N_10311,N_10296);
nor U10590 (N_10590,N_10316,N_10439);
nor U10591 (N_10591,N_10392,N_10320);
and U10592 (N_10592,N_10333,N_10272);
and U10593 (N_10593,N_10324,N_10381);
nor U10594 (N_10594,N_10353,N_10301);
and U10595 (N_10595,N_10481,N_10374);
xnor U10596 (N_10596,N_10268,N_10367);
nand U10597 (N_10597,N_10423,N_10387);
and U10598 (N_10598,N_10425,N_10377);
xor U10599 (N_10599,N_10379,N_10347);
nor U10600 (N_10600,N_10321,N_10332);
xor U10601 (N_10601,N_10309,N_10388);
xor U10602 (N_10602,N_10487,N_10366);
nand U10603 (N_10603,N_10348,N_10295);
or U10604 (N_10604,N_10427,N_10334);
and U10605 (N_10605,N_10315,N_10434);
or U10606 (N_10606,N_10322,N_10335);
nor U10607 (N_10607,N_10401,N_10376);
or U10608 (N_10608,N_10446,N_10461);
nor U10609 (N_10609,N_10406,N_10294);
xor U10610 (N_10610,N_10437,N_10277);
xor U10611 (N_10611,N_10453,N_10259);
xnor U10612 (N_10612,N_10399,N_10303);
nand U10613 (N_10613,N_10441,N_10485);
or U10614 (N_10614,N_10317,N_10327);
or U10615 (N_10615,N_10351,N_10329);
or U10616 (N_10616,N_10344,N_10290);
nor U10617 (N_10617,N_10250,N_10416);
nand U10618 (N_10618,N_10271,N_10424);
or U10619 (N_10619,N_10497,N_10492);
nand U10620 (N_10620,N_10456,N_10373);
nor U10621 (N_10621,N_10278,N_10451);
nand U10622 (N_10622,N_10419,N_10400);
nor U10623 (N_10623,N_10305,N_10341);
nor U10624 (N_10624,N_10270,N_10360);
nand U10625 (N_10625,N_10423,N_10372);
xnor U10626 (N_10626,N_10392,N_10467);
or U10627 (N_10627,N_10350,N_10433);
nand U10628 (N_10628,N_10312,N_10416);
and U10629 (N_10629,N_10363,N_10468);
or U10630 (N_10630,N_10277,N_10465);
nand U10631 (N_10631,N_10483,N_10318);
nand U10632 (N_10632,N_10423,N_10264);
xor U10633 (N_10633,N_10286,N_10348);
nand U10634 (N_10634,N_10479,N_10271);
xor U10635 (N_10635,N_10433,N_10329);
xor U10636 (N_10636,N_10329,N_10391);
xnor U10637 (N_10637,N_10316,N_10321);
nand U10638 (N_10638,N_10481,N_10376);
and U10639 (N_10639,N_10400,N_10425);
nor U10640 (N_10640,N_10340,N_10321);
and U10641 (N_10641,N_10482,N_10379);
and U10642 (N_10642,N_10264,N_10458);
nor U10643 (N_10643,N_10433,N_10361);
xnor U10644 (N_10644,N_10418,N_10329);
and U10645 (N_10645,N_10318,N_10299);
or U10646 (N_10646,N_10461,N_10351);
nor U10647 (N_10647,N_10252,N_10303);
nand U10648 (N_10648,N_10442,N_10366);
or U10649 (N_10649,N_10484,N_10469);
nand U10650 (N_10650,N_10350,N_10441);
nor U10651 (N_10651,N_10274,N_10332);
nand U10652 (N_10652,N_10380,N_10460);
or U10653 (N_10653,N_10423,N_10332);
xor U10654 (N_10654,N_10351,N_10427);
nor U10655 (N_10655,N_10350,N_10336);
or U10656 (N_10656,N_10431,N_10429);
or U10657 (N_10657,N_10358,N_10493);
nor U10658 (N_10658,N_10267,N_10250);
nor U10659 (N_10659,N_10372,N_10410);
and U10660 (N_10660,N_10394,N_10488);
or U10661 (N_10661,N_10343,N_10346);
nand U10662 (N_10662,N_10485,N_10338);
nand U10663 (N_10663,N_10286,N_10478);
nor U10664 (N_10664,N_10315,N_10485);
and U10665 (N_10665,N_10318,N_10463);
nand U10666 (N_10666,N_10322,N_10370);
or U10667 (N_10667,N_10471,N_10457);
and U10668 (N_10668,N_10425,N_10375);
or U10669 (N_10669,N_10413,N_10398);
xor U10670 (N_10670,N_10343,N_10365);
nand U10671 (N_10671,N_10413,N_10421);
or U10672 (N_10672,N_10472,N_10360);
or U10673 (N_10673,N_10431,N_10259);
or U10674 (N_10674,N_10499,N_10404);
nor U10675 (N_10675,N_10280,N_10336);
nand U10676 (N_10676,N_10414,N_10333);
xnor U10677 (N_10677,N_10496,N_10321);
nand U10678 (N_10678,N_10404,N_10445);
nand U10679 (N_10679,N_10346,N_10353);
nor U10680 (N_10680,N_10317,N_10443);
or U10681 (N_10681,N_10364,N_10321);
nor U10682 (N_10682,N_10486,N_10288);
nand U10683 (N_10683,N_10389,N_10291);
xor U10684 (N_10684,N_10364,N_10338);
and U10685 (N_10685,N_10291,N_10250);
or U10686 (N_10686,N_10317,N_10438);
xor U10687 (N_10687,N_10344,N_10309);
nor U10688 (N_10688,N_10459,N_10271);
or U10689 (N_10689,N_10418,N_10346);
or U10690 (N_10690,N_10477,N_10345);
nand U10691 (N_10691,N_10317,N_10390);
nor U10692 (N_10692,N_10489,N_10285);
or U10693 (N_10693,N_10366,N_10447);
nor U10694 (N_10694,N_10292,N_10387);
nand U10695 (N_10695,N_10438,N_10473);
or U10696 (N_10696,N_10441,N_10335);
nor U10697 (N_10697,N_10476,N_10447);
and U10698 (N_10698,N_10285,N_10427);
nor U10699 (N_10699,N_10395,N_10393);
nand U10700 (N_10700,N_10443,N_10276);
xnor U10701 (N_10701,N_10305,N_10431);
nand U10702 (N_10702,N_10274,N_10319);
xor U10703 (N_10703,N_10461,N_10489);
nand U10704 (N_10704,N_10357,N_10286);
xnor U10705 (N_10705,N_10388,N_10472);
and U10706 (N_10706,N_10488,N_10481);
nand U10707 (N_10707,N_10455,N_10270);
nor U10708 (N_10708,N_10439,N_10499);
or U10709 (N_10709,N_10400,N_10472);
nand U10710 (N_10710,N_10378,N_10323);
nor U10711 (N_10711,N_10284,N_10278);
or U10712 (N_10712,N_10489,N_10441);
or U10713 (N_10713,N_10471,N_10493);
and U10714 (N_10714,N_10280,N_10359);
nor U10715 (N_10715,N_10258,N_10350);
nand U10716 (N_10716,N_10374,N_10468);
xnor U10717 (N_10717,N_10342,N_10272);
nor U10718 (N_10718,N_10269,N_10287);
and U10719 (N_10719,N_10361,N_10347);
or U10720 (N_10720,N_10284,N_10465);
nand U10721 (N_10721,N_10315,N_10468);
xnor U10722 (N_10722,N_10330,N_10457);
nand U10723 (N_10723,N_10277,N_10417);
nor U10724 (N_10724,N_10440,N_10346);
and U10725 (N_10725,N_10431,N_10393);
xnor U10726 (N_10726,N_10349,N_10341);
nor U10727 (N_10727,N_10463,N_10328);
or U10728 (N_10728,N_10321,N_10305);
and U10729 (N_10729,N_10375,N_10424);
and U10730 (N_10730,N_10349,N_10383);
xnor U10731 (N_10731,N_10460,N_10439);
xor U10732 (N_10732,N_10317,N_10393);
and U10733 (N_10733,N_10486,N_10408);
or U10734 (N_10734,N_10418,N_10405);
and U10735 (N_10735,N_10306,N_10469);
xor U10736 (N_10736,N_10378,N_10345);
or U10737 (N_10737,N_10494,N_10405);
nor U10738 (N_10738,N_10346,N_10473);
xnor U10739 (N_10739,N_10464,N_10301);
nor U10740 (N_10740,N_10473,N_10434);
nor U10741 (N_10741,N_10312,N_10361);
nor U10742 (N_10742,N_10398,N_10446);
xor U10743 (N_10743,N_10294,N_10479);
and U10744 (N_10744,N_10441,N_10298);
nand U10745 (N_10745,N_10309,N_10314);
xnor U10746 (N_10746,N_10320,N_10294);
nor U10747 (N_10747,N_10397,N_10367);
nor U10748 (N_10748,N_10317,N_10346);
and U10749 (N_10749,N_10439,N_10362);
xor U10750 (N_10750,N_10587,N_10593);
nand U10751 (N_10751,N_10543,N_10722);
nor U10752 (N_10752,N_10630,N_10512);
nor U10753 (N_10753,N_10605,N_10572);
nor U10754 (N_10754,N_10507,N_10730);
nor U10755 (N_10755,N_10599,N_10579);
and U10756 (N_10756,N_10668,N_10501);
or U10757 (N_10757,N_10651,N_10694);
or U10758 (N_10758,N_10531,N_10533);
or U10759 (N_10759,N_10746,N_10739);
or U10760 (N_10760,N_10703,N_10621);
xor U10761 (N_10761,N_10734,N_10673);
nand U10762 (N_10762,N_10596,N_10608);
and U10763 (N_10763,N_10625,N_10679);
and U10764 (N_10764,N_10548,N_10671);
and U10765 (N_10765,N_10697,N_10657);
or U10766 (N_10766,N_10513,N_10591);
nand U10767 (N_10767,N_10552,N_10562);
and U10768 (N_10768,N_10502,N_10615);
or U10769 (N_10769,N_10616,N_10623);
nor U10770 (N_10770,N_10558,N_10660);
nor U10771 (N_10771,N_10690,N_10565);
or U10772 (N_10772,N_10567,N_10656);
and U10773 (N_10773,N_10725,N_10662);
or U10774 (N_10774,N_10546,N_10529);
or U10775 (N_10775,N_10612,N_10652);
or U10776 (N_10776,N_10631,N_10555);
and U10777 (N_10777,N_10653,N_10738);
and U10778 (N_10778,N_10607,N_10594);
nor U10779 (N_10779,N_10520,N_10744);
nand U10780 (N_10780,N_10540,N_10573);
and U10781 (N_10781,N_10667,N_10584);
nor U10782 (N_10782,N_10721,N_10559);
nand U10783 (N_10783,N_10748,N_10505);
and U10784 (N_10784,N_10648,N_10570);
xor U10785 (N_10785,N_10649,N_10664);
or U10786 (N_10786,N_10696,N_10698);
nor U10787 (N_10787,N_10569,N_10613);
nand U10788 (N_10788,N_10692,N_10589);
or U10789 (N_10789,N_10709,N_10655);
or U10790 (N_10790,N_10702,N_10729);
or U10791 (N_10791,N_10586,N_10715);
and U10792 (N_10792,N_10672,N_10574);
xor U10793 (N_10793,N_10609,N_10724);
nor U10794 (N_10794,N_10723,N_10614);
nor U10795 (N_10795,N_10583,N_10517);
or U10796 (N_10796,N_10603,N_10699);
nand U10797 (N_10797,N_10633,N_10598);
and U10798 (N_10798,N_10627,N_10658);
nand U10799 (N_10799,N_10665,N_10522);
nand U10800 (N_10800,N_10680,N_10553);
and U10801 (N_10801,N_10669,N_10560);
or U10802 (N_10802,N_10720,N_10578);
and U10803 (N_10803,N_10708,N_10537);
xor U10804 (N_10804,N_10606,N_10563);
nor U10805 (N_10805,N_10726,N_10564);
or U10806 (N_10806,N_10557,N_10530);
and U10807 (N_10807,N_10595,N_10639);
and U10808 (N_10808,N_10597,N_10687);
or U10809 (N_10809,N_10521,N_10674);
or U10810 (N_10810,N_10685,N_10646);
xor U10811 (N_10811,N_10650,N_10528);
or U10812 (N_10812,N_10618,N_10617);
or U10813 (N_10813,N_10632,N_10727);
nor U10814 (N_10814,N_10515,N_10706);
or U10815 (N_10815,N_10527,N_10740);
or U10816 (N_10816,N_10514,N_10532);
xnor U10817 (N_10817,N_10571,N_10619);
or U10818 (N_10818,N_10675,N_10733);
nand U10819 (N_10819,N_10509,N_10549);
nor U10820 (N_10820,N_10745,N_10535);
nand U10821 (N_10821,N_10676,N_10686);
or U10822 (N_10822,N_10647,N_10731);
or U10823 (N_10823,N_10511,N_10610);
xnor U10824 (N_10824,N_10636,N_10503);
nor U10825 (N_10825,N_10682,N_10714);
or U10826 (N_10826,N_10550,N_10576);
or U10827 (N_10827,N_10622,N_10523);
xor U10828 (N_10828,N_10566,N_10626);
nor U10829 (N_10829,N_10519,N_10749);
or U10830 (N_10830,N_10742,N_10635);
or U10831 (N_10831,N_10638,N_10624);
nor U10832 (N_10832,N_10504,N_10735);
nand U10833 (N_10833,N_10683,N_10666);
nor U10834 (N_10834,N_10604,N_10684);
xnor U10835 (N_10835,N_10590,N_10737);
nor U10836 (N_10836,N_10510,N_10719);
and U10837 (N_10837,N_10732,N_10691);
xnor U10838 (N_10838,N_10556,N_10516);
nor U10839 (N_10839,N_10585,N_10743);
nand U10840 (N_10840,N_10580,N_10678);
xnor U10841 (N_10841,N_10506,N_10701);
and U10842 (N_10842,N_10693,N_10736);
or U10843 (N_10843,N_10539,N_10547);
nor U10844 (N_10844,N_10536,N_10545);
and U10845 (N_10845,N_10641,N_10538);
and U10846 (N_10846,N_10542,N_10601);
and U10847 (N_10847,N_10554,N_10602);
nand U10848 (N_10848,N_10534,N_10654);
and U10849 (N_10849,N_10551,N_10707);
nor U10850 (N_10850,N_10508,N_10541);
nand U10851 (N_10851,N_10592,N_10677);
and U10852 (N_10852,N_10640,N_10718);
nor U10853 (N_10853,N_10561,N_10642);
and U10854 (N_10854,N_10710,N_10500);
or U10855 (N_10855,N_10611,N_10524);
and U10856 (N_10856,N_10645,N_10643);
and U10857 (N_10857,N_10544,N_10689);
nor U10858 (N_10858,N_10600,N_10741);
nand U10859 (N_10859,N_10575,N_10713);
nor U10860 (N_10860,N_10620,N_10568);
and U10861 (N_10861,N_10577,N_10712);
nor U10862 (N_10862,N_10526,N_10628);
xnor U10863 (N_10863,N_10634,N_10629);
and U10864 (N_10864,N_10582,N_10525);
and U10865 (N_10865,N_10663,N_10588);
or U10866 (N_10866,N_10728,N_10695);
and U10867 (N_10867,N_10716,N_10705);
and U10868 (N_10868,N_10659,N_10644);
or U10869 (N_10869,N_10717,N_10637);
xor U10870 (N_10870,N_10518,N_10581);
and U10871 (N_10871,N_10670,N_10661);
and U10872 (N_10872,N_10711,N_10688);
or U10873 (N_10873,N_10747,N_10704);
xnor U10874 (N_10874,N_10681,N_10700);
or U10875 (N_10875,N_10677,N_10729);
or U10876 (N_10876,N_10514,N_10558);
or U10877 (N_10877,N_10715,N_10722);
and U10878 (N_10878,N_10569,N_10741);
nand U10879 (N_10879,N_10555,N_10664);
or U10880 (N_10880,N_10680,N_10606);
or U10881 (N_10881,N_10686,N_10730);
or U10882 (N_10882,N_10733,N_10635);
xor U10883 (N_10883,N_10675,N_10630);
xnor U10884 (N_10884,N_10746,N_10709);
xor U10885 (N_10885,N_10540,N_10517);
nor U10886 (N_10886,N_10681,N_10732);
nand U10887 (N_10887,N_10722,N_10606);
xor U10888 (N_10888,N_10507,N_10505);
xor U10889 (N_10889,N_10618,N_10592);
xnor U10890 (N_10890,N_10694,N_10745);
and U10891 (N_10891,N_10543,N_10639);
or U10892 (N_10892,N_10530,N_10719);
and U10893 (N_10893,N_10684,N_10697);
and U10894 (N_10894,N_10559,N_10526);
or U10895 (N_10895,N_10515,N_10605);
nand U10896 (N_10896,N_10522,N_10655);
xor U10897 (N_10897,N_10555,N_10667);
xor U10898 (N_10898,N_10630,N_10641);
xor U10899 (N_10899,N_10551,N_10733);
and U10900 (N_10900,N_10735,N_10653);
or U10901 (N_10901,N_10640,N_10726);
xor U10902 (N_10902,N_10708,N_10737);
and U10903 (N_10903,N_10697,N_10524);
or U10904 (N_10904,N_10730,N_10671);
and U10905 (N_10905,N_10614,N_10724);
nand U10906 (N_10906,N_10590,N_10502);
xor U10907 (N_10907,N_10506,N_10708);
and U10908 (N_10908,N_10689,N_10659);
or U10909 (N_10909,N_10642,N_10747);
and U10910 (N_10910,N_10504,N_10631);
and U10911 (N_10911,N_10510,N_10566);
or U10912 (N_10912,N_10685,N_10678);
xor U10913 (N_10913,N_10707,N_10569);
nand U10914 (N_10914,N_10747,N_10607);
nor U10915 (N_10915,N_10556,N_10695);
and U10916 (N_10916,N_10657,N_10561);
nand U10917 (N_10917,N_10559,N_10622);
nor U10918 (N_10918,N_10613,N_10658);
xor U10919 (N_10919,N_10650,N_10590);
xnor U10920 (N_10920,N_10731,N_10508);
and U10921 (N_10921,N_10597,N_10622);
nor U10922 (N_10922,N_10700,N_10676);
nor U10923 (N_10923,N_10613,N_10668);
and U10924 (N_10924,N_10505,N_10725);
nand U10925 (N_10925,N_10573,N_10695);
or U10926 (N_10926,N_10656,N_10717);
nor U10927 (N_10927,N_10539,N_10579);
or U10928 (N_10928,N_10536,N_10527);
nand U10929 (N_10929,N_10706,N_10731);
nor U10930 (N_10930,N_10668,N_10718);
or U10931 (N_10931,N_10704,N_10514);
or U10932 (N_10932,N_10635,N_10684);
and U10933 (N_10933,N_10594,N_10529);
nor U10934 (N_10934,N_10697,N_10680);
and U10935 (N_10935,N_10738,N_10582);
xor U10936 (N_10936,N_10523,N_10520);
nor U10937 (N_10937,N_10679,N_10635);
nand U10938 (N_10938,N_10666,N_10623);
or U10939 (N_10939,N_10686,N_10619);
and U10940 (N_10940,N_10529,N_10744);
nor U10941 (N_10941,N_10518,N_10614);
nand U10942 (N_10942,N_10605,N_10665);
nor U10943 (N_10943,N_10540,N_10660);
or U10944 (N_10944,N_10541,N_10719);
nand U10945 (N_10945,N_10620,N_10535);
or U10946 (N_10946,N_10596,N_10638);
or U10947 (N_10947,N_10510,N_10732);
or U10948 (N_10948,N_10622,N_10567);
xor U10949 (N_10949,N_10733,N_10749);
xor U10950 (N_10950,N_10527,N_10721);
nor U10951 (N_10951,N_10703,N_10586);
and U10952 (N_10952,N_10585,N_10660);
xor U10953 (N_10953,N_10529,N_10509);
and U10954 (N_10954,N_10590,N_10655);
nand U10955 (N_10955,N_10633,N_10655);
and U10956 (N_10956,N_10582,N_10675);
nand U10957 (N_10957,N_10564,N_10669);
nor U10958 (N_10958,N_10599,N_10573);
nand U10959 (N_10959,N_10667,N_10621);
or U10960 (N_10960,N_10542,N_10707);
nand U10961 (N_10961,N_10595,N_10590);
xor U10962 (N_10962,N_10530,N_10502);
nand U10963 (N_10963,N_10658,N_10531);
and U10964 (N_10964,N_10621,N_10593);
nand U10965 (N_10965,N_10604,N_10554);
nand U10966 (N_10966,N_10614,N_10662);
nor U10967 (N_10967,N_10695,N_10583);
nor U10968 (N_10968,N_10607,N_10606);
nor U10969 (N_10969,N_10594,N_10698);
xnor U10970 (N_10970,N_10541,N_10545);
nand U10971 (N_10971,N_10599,N_10745);
xor U10972 (N_10972,N_10700,N_10523);
and U10973 (N_10973,N_10559,N_10656);
xor U10974 (N_10974,N_10710,N_10747);
xnor U10975 (N_10975,N_10666,N_10592);
nor U10976 (N_10976,N_10749,N_10534);
nor U10977 (N_10977,N_10743,N_10536);
nor U10978 (N_10978,N_10629,N_10740);
xnor U10979 (N_10979,N_10696,N_10624);
or U10980 (N_10980,N_10527,N_10629);
and U10981 (N_10981,N_10717,N_10721);
xor U10982 (N_10982,N_10698,N_10565);
nand U10983 (N_10983,N_10619,N_10706);
and U10984 (N_10984,N_10589,N_10511);
nand U10985 (N_10985,N_10529,N_10725);
and U10986 (N_10986,N_10745,N_10645);
xnor U10987 (N_10987,N_10714,N_10695);
nand U10988 (N_10988,N_10502,N_10611);
nor U10989 (N_10989,N_10613,N_10575);
nor U10990 (N_10990,N_10723,N_10556);
nor U10991 (N_10991,N_10616,N_10520);
or U10992 (N_10992,N_10747,N_10715);
nand U10993 (N_10993,N_10711,N_10742);
nand U10994 (N_10994,N_10565,N_10563);
and U10995 (N_10995,N_10746,N_10527);
nand U10996 (N_10996,N_10695,N_10699);
nand U10997 (N_10997,N_10509,N_10552);
and U10998 (N_10998,N_10707,N_10608);
and U10999 (N_10999,N_10663,N_10597);
and U11000 (N_11000,N_10755,N_10975);
nor U11001 (N_11001,N_10992,N_10839);
xnor U11002 (N_11002,N_10811,N_10929);
nand U11003 (N_11003,N_10916,N_10955);
and U11004 (N_11004,N_10984,N_10849);
or U11005 (N_11005,N_10863,N_10959);
or U11006 (N_11006,N_10936,N_10951);
and U11007 (N_11007,N_10878,N_10753);
nand U11008 (N_11008,N_10952,N_10870);
or U11009 (N_11009,N_10902,N_10911);
nand U11010 (N_11010,N_10773,N_10832);
nand U11011 (N_11011,N_10901,N_10893);
xnor U11012 (N_11012,N_10971,N_10814);
or U11013 (N_11013,N_10816,N_10809);
and U11014 (N_11014,N_10977,N_10801);
nor U11015 (N_11015,N_10821,N_10833);
xor U11016 (N_11016,N_10790,N_10986);
or U11017 (N_11017,N_10835,N_10912);
xor U11018 (N_11018,N_10909,N_10823);
nor U11019 (N_11019,N_10907,N_10824);
and U11020 (N_11020,N_10879,N_10787);
xor U11021 (N_11021,N_10890,N_10886);
and U11022 (N_11022,N_10953,N_10758);
xor U11023 (N_11023,N_10900,N_10923);
and U11024 (N_11024,N_10813,N_10922);
and U11025 (N_11025,N_10750,N_10966);
nand U11026 (N_11026,N_10976,N_10892);
xor U11027 (N_11027,N_10974,N_10856);
or U11028 (N_11028,N_10874,N_10961);
nor U11029 (N_11029,N_10882,N_10777);
and U11030 (N_11030,N_10838,N_10967);
nand U11031 (N_11031,N_10990,N_10830);
nand U11032 (N_11032,N_10941,N_10866);
xor U11033 (N_11033,N_10931,N_10751);
nand U11034 (N_11034,N_10897,N_10972);
xor U11035 (N_11035,N_10895,N_10978);
and U11036 (N_11036,N_10855,N_10829);
nor U11037 (N_11037,N_10812,N_10915);
nor U11038 (N_11038,N_10857,N_10919);
nor U11039 (N_11039,N_10944,N_10793);
nor U11040 (N_11040,N_10756,N_10840);
xnor U11041 (N_11041,N_10752,N_10780);
and U11042 (N_11042,N_10965,N_10876);
nor U11043 (N_11043,N_10917,N_10921);
or U11044 (N_11044,N_10940,N_10935);
or U11045 (N_11045,N_10846,N_10881);
nor U11046 (N_11046,N_10904,N_10837);
nor U11047 (N_11047,N_10760,N_10864);
xor U11048 (N_11048,N_10762,N_10989);
xor U11049 (N_11049,N_10981,N_10873);
and U11050 (N_11050,N_10920,N_10867);
nand U11051 (N_11051,N_10774,N_10903);
or U11052 (N_11052,N_10898,N_10982);
or U11053 (N_11053,N_10754,N_10788);
and U11054 (N_11054,N_10905,N_10943);
and U11055 (N_11055,N_10791,N_10785);
nand U11056 (N_11056,N_10875,N_10843);
xor U11057 (N_11057,N_10766,N_10947);
nand U11058 (N_11058,N_10808,N_10850);
xnor U11059 (N_11059,N_10815,N_10805);
or U11060 (N_11060,N_10862,N_10995);
nand U11061 (N_11061,N_10980,N_10770);
nor U11062 (N_11062,N_10871,N_10860);
and U11063 (N_11063,N_10759,N_10767);
nor U11064 (N_11064,N_10776,N_10956);
xor U11065 (N_11065,N_10988,N_10768);
nor U11066 (N_11066,N_10970,N_10964);
and U11067 (N_11067,N_10819,N_10845);
xnor U11068 (N_11068,N_10854,N_10769);
nand U11069 (N_11069,N_10859,N_10868);
nand U11070 (N_11070,N_10872,N_10851);
xnor U11071 (N_11071,N_10834,N_10979);
nand U11072 (N_11072,N_10803,N_10925);
and U11073 (N_11073,N_10884,N_10764);
nand U11074 (N_11074,N_10927,N_10889);
nor U11075 (N_11075,N_10782,N_10847);
nand U11076 (N_11076,N_10877,N_10945);
xor U11077 (N_11077,N_10786,N_10858);
or U11078 (N_11078,N_10896,N_10985);
or U11079 (N_11079,N_10825,N_10963);
nand U11080 (N_11080,N_10802,N_10761);
or U11081 (N_11081,N_10796,N_10807);
nand U11082 (N_11082,N_10842,N_10998);
nor U11083 (N_11083,N_10810,N_10932);
nor U11084 (N_11084,N_10831,N_10918);
nor U11085 (N_11085,N_10894,N_10983);
and U11086 (N_11086,N_10910,N_10869);
and U11087 (N_11087,N_10844,N_10954);
nand U11088 (N_11088,N_10775,N_10899);
nand U11089 (N_11089,N_10934,N_10827);
nor U11090 (N_11090,N_10926,N_10973);
and U11091 (N_11091,N_10933,N_10960);
nor U11092 (N_11092,N_10993,N_10930);
or U11093 (N_11093,N_10861,N_10928);
nand U11094 (N_11094,N_10772,N_10853);
nor U11095 (N_11095,N_10883,N_10778);
xor U11096 (N_11096,N_10997,N_10800);
or U11097 (N_11097,N_10942,N_10820);
and U11098 (N_11098,N_10783,N_10806);
nor U11099 (N_11099,N_10924,N_10996);
or U11100 (N_11100,N_10987,N_10913);
or U11101 (N_11101,N_10962,N_10880);
nor U11102 (N_11102,N_10999,N_10958);
nor U11103 (N_11103,N_10781,N_10799);
nor U11104 (N_11104,N_10957,N_10949);
and U11105 (N_11105,N_10784,N_10822);
nand U11106 (N_11106,N_10795,N_10826);
nand U11107 (N_11107,N_10771,N_10779);
xnor U11108 (N_11108,N_10797,N_10804);
nor U11109 (N_11109,N_10938,N_10757);
or U11110 (N_11110,N_10969,N_10836);
nor U11111 (N_11111,N_10937,N_10906);
or U11112 (N_11112,N_10794,N_10885);
and U11113 (N_11113,N_10789,N_10828);
and U11114 (N_11114,N_10818,N_10765);
or U11115 (N_11115,N_10968,N_10841);
nand U11116 (N_11116,N_10991,N_10763);
xor U11117 (N_11117,N_10888,N_10939);
nand U11118 (N_11118,N_10994,N_10891);
nor U11119 (N_11119,N_10908,N_10817);
xnor U11120 (N_11120,N_10792,N_10887);
and U11121 (N_11121,N_10948,N_10914);
or U11122 (N_11122,N_10798,N_10852);
or U11123 (N_11123,N_10950,N_10865);
xnor U11124 (N_11124,N_10946,N_10848);
nand U11125 (N_11125,N_10908,N_10988);
nor U11126 (N_11126,N_10878,N_10797);
nand U11127 (N_11127,N_10814,N_10893);
or U11128 (N_11128,N_10869,N_10928);
nor U11129 (N_11129,N_10778,N_10801);
nand U11130 (N_11130,N_10994,N_10956);
xor U11131 (N_11131,N_10827,N_10817);
xor U11132 (N_11132,N_10903,N_10759);
xnor U11133 (N_11133,N_10936,N_10847);
and U11134 (N_11134,N_10951,N_10938);
and U11135 (N_11135,N_10958,N_10916);
or U11136 (N_11136,N_10779,N_10960);
xnor U11137 (N_11137,N_10908,N_10957);
and U11138 (N_11138,N_10885,N_10970);
and U11139 (N_11139,N_10882,N_10865);
and U11140 (N_11140,N_10918,N_10993);
nor U11141 (N_11141,N_10813,N_10892);
or U11142 (N_11142,N_10796,N_10922);
xnor U11143 (N_11143,N_10941,N_10909);
xor U11144 (N_11144,N_10834,N_10896);
and U11145 (N_11145,N_10926,N_10772);
nand U11146 (N_11146,N_10827,N_10942);
and U11147 (N_11147,N_10887,N_10910);
and U11148 (N_11148,N_10869,N_10904);
nand U11149 (N_11149,N_10806,N_10921);
and U11150 (N_11150,N_10882,N_10845);
nor U11151 (N_11151,N_10909,N_10906);
and U11152 (N_11152,N_10989,N_10831);
or U11153 (N_11153,N_10904,N_10846);
nand U11154 (N_11154,N_10923,N_10991);
or U11155 (N_11155,N_10809,N_10837);
nor U11156 (N_11156,N_10819,N_10818);
nand U11157 (N_11157,N_10773,N_10924);
nand U11158 (N_11158,N_10878,N_10824);
nand U11159 (N_11159,N_10787,N_10925);
or U11160 (N_11160,N_10944,N_10970);
nor U11161 (N_11161,N_10911,N_10824);
or U11162 (N_11162,N_10940,N_10878);
xnor U11163 (N_11163,N_10915,N_10868);
and U11164 (N_11164,N_10851,N_10856);
and U11165 (N_11165,N_10795,N_10981);
xor U11166 (N_11166,N_10816,N_10946);
nor U11167 (N_11167,N_10822,N_10813);
and U11168 (N_11168,N_10862,N_10883);
nor U11169 (N_11169,N_10811,N_10829);
nand U11170 (N_11170,N_10994,N_10864);
and U11171 (N_11171,N_10845,N_10901);
or U11172 (N_11172,N_10924,N_10829);
nor U11173 (N_11173,N_10900,N_10958);
and U11174 (N_11174,N_10868,N_10910);
or U11175 (N_11175,N_10879,N_10851);
nor U11176 (N_11176,N_10814,N_10983);
nand U11177 (N_11177,N_10864,N_10940);
and U11178 (N_11178,N_10882,N_10775);
nand U11179 (N_11179,N_10788,N_10965);
nand U11180 (N_11180,N_10808,N_10901);
or U11181 (N_11181,N_10793,N_10838);
nand U11182 (N_11182,N_10804,N_10815);
xnor U11183 (N_11183,N_10928,N_10935);
xnor U11184 (N_11184,N_10858,N_10888);
or U11185 (N_11185,N_10792,N_10775);
or U11186 (N_11186,N_10866,N_10933);
or U11187 (N_11187,N_10919,N_10849);
nand U11188 (N_11188,N_10764,N_10983);
xor U11189 (N_11189,N_10828,N_10762);
xnor U11190 (N_11190,N_10993,N_10834);
nor U11191 (N_11191,N_10926,N_10756);
xnor U11192 (N_11192,N_10924,N_10902);
and U11193 (N_11193,N_10936,N_10809);
and U11194 (N_11194,N_10786,N_10813);
xnor U11195 (N_11195,N_10865,N_10768);
nand U11196 (N_11196,N_10788,N_10791);
and U11197 (N_11197,N_10848,N_10884);
xor U11198 (N_11198,N_10775,N_10881);
nand U11199 (N_11199,N_10771,N_10809);
nand U11200 (N_11200,N_10953,N_10934);
and U11201 (N_11201,N_10982,N_10853);
and U11202 (N_11202,N_10855,N_10843);
nor U11203 (N_11203,N_10911,N_10785);
nor U11204 (N_11204,N_10823,N_10967);
xnor U11205 (N_11205,N_10788,N_10847);
nand U11206 (N_11206,N_10834,N_10903);
or U11207 (N_11207,N_10806,N_10983);
or U11208 (N_11208,N_10847,N_10931);
nor U11209 (N_11209,N_10790,N_10847);
and U11210 (N_11210,N_10805,N_10947);
nand U11211 (N_11211,N_10759,N_10799);
or U11212 (N_11212,N_10968,N_10982);
xor U11213 (N_11213,N_10974,N_10801);
nor U11214 (N_11214,N_10982,N_10790);
xnor U11215 (N_11215,N_10850,N_10822);
or U11216 (N_11216,N_10898,N_10806);
or U11217 (N_11217,N_10865,N_10911);
nand U11218 (N_11218,N_10848,N_10833);
xor U11219 (N_11219,N_10950,N_10837);
nand U11220 (N_11220,N_10944,N_10882);
nand U11221 (N_11221,N_10964,N_10887);
xnor U11222 (N_11222,N_10798,N_10860);
xnor U11223 (N_11223,N_10812,N_10806);
nand U11224 (N_11224,N_10754,N_10897);
xor U11225 (N_11225,N_10916,N_10925);
nand U11226 (N_11226,N_10756,N_10908);
nor U11227 (N_11227,N_10784,N_10754);
xor U11228 (N_11228,N_10857,N_10778);
nor U11229 (N_11229,N_10808,N_10803);
nor U11230 (N_11230,N_10843,N_10799);
xnor U11231 (N_11231,N_10990,N_10906);
and U11232 (N_11232,N_10877,N_10776);
xnor U11233 (N_11233,N_10847,N_10764);
and U11234 (N_11234,N_10818,N_10837);
and U11235 (N_11235,N_10902,N_10941);
and U11236 (N_11236,N_10814,N_10999);
or U11237 (N_11237,N_10833,N_10964);
or U11238 (N_11238,N_10852,N_10903);
and U11239 (N_11239,N_10836,N_10895);
or U11240 (N_11240,N_10925,N_10790);
or U11241 (N_11241,N_10835,N_10901);
and U11242 (N_11242,N_10955,N_10825);
xor U11243 (N_11243,N_10815,N_10934);
xor U11244 (N_11244,N_10919,N_10909);
nand U11245 (N_11245,N_10997,N_10974);
xor U11246 (N_11246,N_10779,N_10961);
or U11247 (N_11247,N_10988,N_10984);
nand U11248 (N_11248,N_10845,N_10970);
or U11249 (N_11249,N_10994,N_10768);
xor U11250 (N_11250,N_11094,N_11069);
or U11251 (N_11251,N_11011,N_11140);
or U11252 (N_11252,N_11249,N_11233);
nor U11253 (N_11253,N_11131,N_11063);
and U11254 (N_11254,N_11203,N_11006);
nand U11255 (N_11255,N_11231,N_11126);
nor U11256 (N_11256,N_11236,N_11220);
and U11257 (N_11257,N_11205,N_11034);
or U11258 (N_11258,N_11056,N_11244);
nor U11259 (N_11259,N_11014,N_11246);
xnor U11260 (N_11260,N_11076,N_11208);
or U11261 (N_11261,N_11184,N_11122);
xor U11262 (N_11262,N_11241,N_11147);
nor U11263 (N_11263,N_11234,N_11007);
or U11264 (N_11264,N_11017,N_11188);
nor U11265 (N_11265,N_11004,N_11186);
and U11266 (N_11266,N_11127,N_11087);
nor U11267 (N_11267,N_11105,N_11039);
and U11268 (N_11268,N_11030,N_11154);
xnor U11269 (N_11269,N_11183,N_11120);
or U11270 (N_11270,N_11042,N_11185);
and U11271 (N_11271,N_11061,N_11035);
nand U11272 (N_11272,N_11202,N_11070);
xnor U11273 (N_11273,N_11113,N_11168);
nor U11274 (N_11274,N_11060,N_11074);
and U11275 (N_11275,N_11090,N_11083);
nand U11276 (N_11276,N_11046,N_11098);
or U11277 (N_11277,N_11107,N_11193);
or U11278 (N_11278,N_11002,N_11165);
nand U11279 (N_11279,N_11163,N_11081);
nor U11280 (N_11280,N_11211,N_11102);
or U11281 (N_11281,N_11169,N_11027);
or U11282 (N_11282,N_11130,N_11172);
or U11283 (N_11283,N_11104,N_11100);
and U11284 (N_11284,N_11182,N_11155);
and U11285 (N_11285,N_11103,N_11020);
or U11286 (N_11286,N_11051,N_11111);
nand U11287 (N_11287,N_11162,N_11115);
or U11288 (N_11288,N_11174,N_11239);
xor U11289 (N_11289,N_11093,N_11227);
and U11290 (N_11290,N_11071,N_11065);
nand U11291 (N_11291,N_11114,N_11134);
nand U11292 (N_11292,N_11116,N_11132);
or U11293 (N_11293,N_11024,N_11119);
and U11294 (N_11294,N_11009,N_11232);
xnor U11295 (N_11295,N_11237,N_11179);
and U11296 (N_11296,N_11075,N_11175);
and U11297 (N_11297,N_11044,N_11156);
or U11298 (N_11298,N_11078,N_11141);
and U11299 (N_11299,N_11243,N_11040);
nand U11300 (N_11300,N_11230,N_11146);
and U11301 (N_11301,N_11021,N_11109);
or U11302 (N_11302,N_11229,N_11047);
nand U11303 (N_11303,N_11137,N_11041);
xor U11304 (N_11304,N_11150,N_11158);
xor U11305 (N_11305,N_11210,N_11072);
and U11306 (N_11306,N_11191,N_11173);
nor U11307 (N_11307,N_11110,N_11023);
xnor U11308 (N_11308,N_11057,N_11053);
xor U11309 (N_11309,N_11187,N_11050);
xor U11310 (N_11310,N_11149,N_11048);
xor U11311 (N_11311,N_11095,N_11031);
xor U11312 (N_11312,N_11003,N_11022);
nand U11313 (N_11313,N_11223,N_11121);
and U11314 (N_11314,N_11153,N_11089);
or U11315 (N_11315,N_11190,N_11088);
nor U11316 (N_11316,N_11008,N_11224);
nor U11317 (N_11317,N_11189,N_11062);
xnor U11318 (N_11318,N_11079,N_11195);
or U11319 (N_11319,N_11219,N_11038);
nand U11320 (N_11320,N_11215,N_11178);
nand U11321 (N_11321,N_11043,N_11036);
xnor U11322 (N_11322,N_11181,N_11240);
nand U11323 (N_11323,N_11054,N_11139);
or U11324 (N_11324,N_11064,N_11026);
nand U11325 (N_11325,N_11018,N_11029);
nand U11326 (N_11326,N_11108,N_11001);
nor U11327 (N_11327,N_11016,N_11217);
and U11328 (N_11328,N_11086,N_11222);
nand U11329 (N_11329,N_11138,N_11013);
nand U11330 (N_11330,N_11037,N_11199);
and U11331 (N_11331,N_11144,N_11052);
or U11332 (N_11332,N_11152,N_11067);
and U11333 (N_11333,N_11133,N_11209);
or U11334 (N_11334,N_11101,N_11025);
xor U11335 (N_11335,N_11012,N_11032);
nor U11336 (N_11336,N_11245,N_11143);
xor U11337 (N_11337,N_11207,N_11160);
nand U11338 (N_11338,N_11055,N_11212);
nand U11339 (N_11339,N_11148,N_11015);
nand U11340 (N_11340,N_11028,N_11091);
nand U11341 (N_11341,N_11176,N_11033);
nor U11342 (N_11342,N_11082,N_11180);
and U11343 (N_11343,N_11198,N_11005);
xnor U11344 (N_11344,N_11106,N_11068);
nor U11345 (N_11345,N_11196,N_11092);
nand U11346 (N_11346,N_11213,N_11096);
nand U11347 (N_11347,N_11216,N_11214);
nor U11348 (N_11348,N_11010,N_11226);
or U11349 (N_11349,N_11118,N_11161);
xor U11350 (N_11350,N_11200,N_11049);
or U11351 (N_11351,N_11084,N_11097);
xnor U11352 (N_11352,N_11170,N_11123);
nor U11353 (N_11353,N_11228,N_11000);
nor U11354 (N_11354,N_11166,N_11066);
nor U11355 (N_11355,N_11059,N_11077);
or U11356 (N_11356,N_11019,N_11225);
xor U11357 (N_11357,N_11073,N_11204);
and U11358 (N_11358,N_11197,N_11080);
nand U11359 (N_11359,N_11221,N_11248);
nand U11360 (N_11360,N_11117,N_11124);
nor U11361 (N_11361,N_11128,N_11099);
xor U11362 (N_11362,N_11247,N_11159);
and U11363 (N_11363,N_11242,N_11218);
xor U11364 (N_11364,N_11145,N_11136);
or U11365 (N_11365,N_11167,N_11157);
xnor U11366 (N_11366,N_11192,N_11085);
xor U11367 (N_11367,N_11125,N_11238);
and U11368 (N_11368,N_11045,N_11171);
nand U11369 (N_11369,N_11206,N_11235);
and U11370 (N_11370,N_11177,N_11151);
and U11371 (N_11371,N_11112,N_11129);
nand U11372 (N_11372,N_11164,N_11201);
and U11373 (N_11373,N_11058,N_11135);
nand U11374 (N_11374,N_11194,N_11142);
nor U11375 (N_11375,N_11049,N_11096);
xnor U11376 (N_11376,N_11051,N_11105);
nor U11377 (N_11377,N_11078,N_11139);
and U11378 (N_11378,N_11113,N_11167);
or U11379 (N_11379,N_11186,N_11023);
and U11380 (N_11380,N_11124,N_11227);
nor U11381 (N_11381,N_11117,N_11004);
nor U11382 (N_11382,N_11043,N_11195);
nand U11383 (N_11383,N_11143,N_11249);
and U11384 (N_11384,N_11176,N_11186);
or U11385 (N_11385,N_11027,N_11077);
nor U11386 (N_11386,N_11057,N_11003);
xor U11387 (N_11387,N_11192,N_11150);
nand U11388 (N_11388,N_11154,N_11200);
xnor U11389 (N_11389,N_11018,N_11176);
xnor U11390 (N_11390,N_11226,N_11100);
and U11391 (N_11391,N_11047,N_11038);
xnor U11392 (N_11392,N_11016,N_11035);
and U11393 (N_11393,N_11127,N_11149);
nand U11394 (N_11394,N_11110,N_11025);
or U11395 (N_11395,N_11219,N_11199);
nand U11396 (N_11396,N_11044,N_11023);
nor U11397 (N_11397,N_11006,N_11130);
xnor U11398 (N_11398,N_11160,N_11235);
nor U11399 (N_11399,N_11207,N_11235);
nand U11400 (N_11400,N_11222,N_11133);
nor U11401 (N_11401,N_11101,N_11042);
or U11402 (N_11402,N_11249,N_11139);
nor U11403 (N_11403,N_11235,N_11094);
nand U11404 (N_11404,N_11159,N_11214);
xor U11405 (N_11405,N_11243,N_11027);
nor U11406 (N_11406,N_11072,N_11190);
xnor U11407 (N_11407,N_11071,N_11012);
nor U11408 (N_11408,N_11236,N_11192);
or U11409 (N_11409,N_11084,N_11017);
and U11410 (N_11410,N_11152,N_11009);
nand U11411 (N_11411,N_11152,N_11241);
and U11412 (N_11412,N_11232,N_11211);
nand U11413 (N_11413,N_11175,N_11118);
or U11414 (N_11414,N_11081,N_11039);
nand U11415 (N_11415,N_11014,N_11189);
nor U11416 (N_11416,N_11039,N_11192);
nand U11417 (N_11417,N_11162,N_11133);
nand U11418 (N_11418,N_11223,N_11111);
nand U11419 (N_11419,N_11212,N_11245);
or U11420 (N_11420,N_11068,N_11180);
and U11421 (N_11421,N_11167,N_11112);
nor U11422 (N_11422,N_11092,N_11225);
or U11423 (N_11423,N_11086,N_11154);
xnor U11424 (N_11424,N_11202,N_11133);
nor U11425 (N_11425,N_11028,N_11217);
or U11426 (N_11426,N_11005,N_11075);
or U11427 (N_11427,N_11149,N_11179);
xor U11428 (N_11428,N_11048,N_11229);
nor U11429 (N_11429,N_11228,N_11038);
xor U11430 (N_11430,N_11092,N_11173);
nand U11431 (N_11431,N_11051,N_11036);
nor U11432 (N_11432,N_11209,N_11005);
and U11433 (N_11433,N_11074,N_11109);
nor U11434 (N_11434,N_11201,N_11072);
and U11435 (N_11435,N_11175,N_11064);
xor U11436 (N_11436,N_11235,N_11111);
nand U11437 (N_11437,N_11099,N_11045);
nand U11438 (N_11438,N_11069,N_11210);
nand U11439 (N_11439,N_11089,N_11104);
nor U11440 (N_11440,N_11202,N_11062);
or U11441 (N_11441,N_11067,N_11089);
nor U11442 (N_11442,N_11037,N_11029);
or U11443 (N_11443,N_11170,N_11030);
and U11444 (N_11444,N_11093,N_11137);
nor U11445 (N_11445,N_11106,N_11230);
or U11446 (N_11446,N_11127,N_11004);
or U11447 (N_11447,N_11185,N_11074);
or U11448 (N_11448,N_11012,N_11067);
and U11449 (N_11449,N_11130,N_11242);
nand U11450 (N_11450,N_11047,N_11008);
and U11451 (N_11451,N_11224,N_11213);
nand U11452 (N_11452,N_11111,N_11069);
nor U11453 (N_11453,N_11127,N_11058);
xor U11454 (N_11454,N_11095,N_11042);
and U11455 (N_11455,N_11230,N_11165);
and U11456 (N_11456,N_11136,N_11106);
and U11457 (N_11457,N_11111,N_11201);
xnor U11458 (N_11458,N_11020,N_11230);
and U11459 (N_11459,N_11026,N_11020);
or U11460 (N_11460,N_11218,N_11160);
or U11461 (N_11461,N_11022,N_11119);
and U11462 (N_11462,N_11057,N_11099);
nor U11463 (N_11463,N_11064,N_11156);
xor U11464 (N_11464,N_11145,N_11241);
xnor U11465 (N_11465,N_11147,N_11221);
xor U11466 (N_11466,N_11094,N_11028);
and U11467 (N_11467,N_11219,N_11225);
nor U11468 (N_11468,N_11145,N_11215);
nor U11469 (N_11469,N_11194,N_11003);
and U11470 (N_11470,N_11195,N_11232);
nand U11471 (N_11471,N_11182,N_11004);
xor U11472 (N_11472,N_11212,N_11153);
and U11473 (N_11473,N_11144,N_11089);
xnor U11474 (N_11474,N_11199,N_11059);
nand U11475 (N_11475,N_11004,N_11073);
xor U11476 (N_11476,N_11043,N_11141);
xnor U11477 (N_11477,N_11181,N_11180);
or U11478 (N_11478,N_11131,N_11068);
or U11479 (N_11479,N_11131,N_11247);
nor U11480 (N_11480,N_11166,N_11032);
xnor U11481 (N_11481,N_11234,N_11135);
xor U11482 (N_11482,N_11186,N_11225);
or U11483 (N_11483,N_11210,N_11126);
nor U11484 (N_11484,N_11067,N_11191);
or U11485 (N_11485,N_11050,N_11146);
xor U11486 (N_11486,N_11193,N_11146);
xnor U11487 (N_11487,N_11182,N_11160);
xnor U11488 (N_11488,N_11149,N_11067);
nand U11489 (N_11489,N_11245,N_11185);
or U11490 (N_11490,N_11012,N_11222);
nor U11491 (N_11491,N_11144,N_11245);
xor U11492 (N_11492,N_11092,N_11205);
or U11493 (N_11493,N_11223,N_11138);
or U11494 (N_11494,N_11142,N_11092);
and U11495 (N_11495,N_11101,N_11097);
and U11496 (N_11496,N_11151,N_11223);
nor U11497 (N_11497,N_11000,N_11056);
xnor U11498 (N_11498,N_11094,N_11089);
and U11499 (N_11499,N_11211,N_11161);
or U11500 (N_11500,N_11297,N_11478);
nor U11501 (N_11501,N_11488,N_11349);
nor U11502 (N_11502,N_11359,N_11264);
and U11503 (N_11503,N_11282,N_11269);
nor U11504 (N_11504,N_11321,N_11270);
nand U11505 (N_11505,N_11430,N_11258);
xnor U11506 (N_11506,N_11473,N_11303);
nand U11507 (N_11507,N_11437,N_11362);
and U11508 (N_11508,N_11479,N_11256);
nand U11509 (N_11509,N_11317,N_11419);
xnor U11510 (N_11510,N_11277,N_11391);
or U11511 (N_11511,N_11443,N_11475);
and U11512 (N_11512,N_11451,N_11330);
xor U11513 (N_11513,N_11375,N_11319);
or U11514 (N_11514,N_11352,N_11260);
nor U11515 (N_11515,N_11315,N_11445);
and U11516 (N_11516,N_11374,N_11403);
nand U11517 (N_11517,N_11275,N_11448);
xnor U11518 (N_11518,N_11398,N_11407);
or U11519 (N_11519,N_11386,N_11463);
xnor U11520 (N_11520,N_11265,N_11369);
and U11521 (N_11521,N_11438,N_11339);
or U11522 (N_11522,N_11356,N_11471);
nor U11523 (N_11523,N_11468,N_11323);
and U11524 (N_11524,N_11484,N_11287);
or U11525 (N_11525,N_11461,N_11395);
or U11526 (N_11526,N_11472,N_11279);
or U11527 (N_11527,N_11316,N_11253);
nor U11528 (N_11528,N_11283,N_11465);
xor U11529 (N_11529,N_11254,N_11492);
or U11530 (N_11530,N_11347,N_11299);
or U11531 (N_11531,N_11425,N_11250);
xor U11532 (N_11532,N_11336,N_11453);
nand U11533 (N_11533,N_11482,N_11309);
or U11534 (N_11534,N_11284,N_11289);
nor U11535 (N_11535,N_11450,N_11285);
or U11536 (N_11536,N_11385,N_11298);
xnor U11537 (N_11537,N_11392,N_11486);
nand U11538 (N_11538,N_11312,N_11344);
nor U11539 (N_11539,N_11380,N_11435);
and U11540 (N_11540,N_11459,N_11396);
nand U11541 (N_11541,N_11372,N_11367);
nor U11542 (N_11542,N_11333,N_11263);
nor U11543 (N_11543,N_11278,N_11497);
nand U11544 (N_11544,N_11409,N_11365);
or U11545 (N_11545,N_11257,N_11410);
nor U11546 (N_11546,N_11268,N_11259);
nor U11547 (N_11547,N_11329,N_11480);
xor U11548 (N_11548,N_11308,N_11417);
or U11549 (N_11549,N_11304,N_11255);
nor U11550 (N_11550,N_11483,N_11360);
or U11551 (N_11551,N_11357,N_11455);
nor U11552 (N_11552,N_11481,N_11301);
and U11553 (N_11553,N_11293,N_11324);
or U11554 (N_11554,N_11311,N_11320);
nand U11555 (N_11555,N_11427,N_11408);
or U11556 (N_11556,N_11335,N_11322);
xor U11557 (N_11557,N_11341,N_11383);
xor U11558 (N_11558,N_11251,N_11397);
and U11559 (N_11559,N_11416,N_11426);
or U11560 (N_11560,N_11389,N_11456);
nand U11561 (N_11561,N_11373,N_11272);
xnor U11562 (N_11562,N_11493,N_11495);
xor U11563 (N_11563,N_11280,N_11305);
or U11564 (N_11564,N_11420,N_11345);
nor U11565 (N_11565,N_11469,N_11368);
and U11566 (N_11566,N_11381,N_11432);
xnor U11567 (N_11567,N_11325,N_11418);
xor U11568 (N_11568,N_11262,N_11485);
nand U11569 (N_11569,N_11387,N_11370);
nor U11570 (N_11570,N_11444,N_11252);
nand U11571 (N_11571,N_11400,N_11464);
and U11572 (N_11572,N_11394,N_11361);
nor U11573 (N_11573,N_11494,N_11490);
or U11574 (N_11574,N_11292,N_11281);
and U11575 (N_11575,N_11348,N_11328);
nand U11576 (N_11576,N_11466,N_11449);
or U11577 (N_11577,N_11390,N_11261);
or U11578 (N_11578,N_11379,N_11428);
and U11579 (N_11579,N_11286,N_11405);
or U11580 (N_11580,N_11441,N_11306);
and U11581 (N_11581,N_11295,N_11462);
nor U11582 (N_11582,N_11440,N_11499);
and U11583 (N_11583,N_11291,N_11331);
xor U11584 (N_11584,N_11267,N_11354);
nand U11585 (N_11585,N_11414,N_11489);
nor U11586 (N_11586,N_11477,N_11366);
xnor U11587 (N_11587,N_11431,N_11314);
or U11588 (N_11588,N_11340,N_11274);
nand U11589 (N_11589,N_11326,N_11351);
or U11590 (N_11590,N_11288,N_11327);
or U11591 (N_11591,N_11310,N_11415);
nand U11592 (N_11592,N_11377,N_11358);
nand U11593 (N_11593,N_11439,N_11364);
and U11594 (N_11594,N_11470,N_11302);
or U11595 (N_11595,N_11434,N_11436);
or U11596 (N_11596,N_11457,N_11424);
xor U11597 (N_11597,N_11353,N_11307);
or U11598 (N_11598,N_11423,N_11313);
and U11599 (N_11599,N_11447,N_11371);
nand U11600 (N_11600,N_11266,N_11346);
nand U11601 (N_11601,N_11446,N_11402);
nor U11602 (N_11602,N_11296,N_11496);
and U11603 (N_11603,N_11337,N_11384);
nand U11604 (N_11604,N_11452,N_11338);
or U11605 (N_11605,N_11498,N_11388);
nor U11606 (N_11606,N_11382,N_11454);
nand U11607 (N_11607,N_11294,N_11290);
and U11608 (N_11608,N_11378,N_11276);
xor U11609 (N_11609,N_11491,N_11442);
xor U11610 (N_11610,N_11411,N_11355);
nor U11611 (N_11611,N_11476,N_11332);
nor U11612 (N_11612,N_11467,N_11460);
or U11613 (N_11613,N_11433,N_11404);
and U11614 (N_11614,N_11273,N_11406);
nor U11615 (N_11615,N_11421,N_11458);
or U11616 (N_11616,N_11318,N_11401);
nand U11617 (N_11617,N_11343,N_11393);
xor U11618 (N_11618,N_11399,N_11363);
nand U11619 (N_11619,N_11487,N_11474);
nand U11620 (N_11620,N_11334,N_11376);
or U11621 (N_11621,N_11350,N_11271);
and U11622 (N_11622,N_11412,N_11429);
xor U11623 (N_11623,N_11342,N_11422);
and U11624 (N_11624,N_11413,N_11300);
nand U11625 (N_11625,N_11452,N_11268);
nand U11626 (N_11626,N_11398,N_11490);
nand U11627 (N_11627,N_11273,N_11356);
nand U11628 (N_11628,N_11394,N_11342);
xor U11629 (N_11629,N_11356,N_11306);
nor U11630 (N_11630,N_11315,N_11374);
xor U11631 (N_11631,N_11478,N_11492);
nor U11632 (N_11632,N_11257,N_11363);
or U11633 (N_11633,N_11437,N_11285);
xor U11634 (N_11634,N_11357,N_11264);
and U11635 (N_11635,N_11327,N_11392);
and U11636 (N_11636,N_11266,N_11414);
xor U11637 (N_11637,N_11261,N_11311);
or U11638 (N_11638,N_11280,N_11456);
nand U11639 (N_11639,N_11310,N_11357);
or U11640 (N_11640,N_11278,N_11474);
or U11641 (N_11641,N_11316,N_11461);
or U11642 (N_11642,N_11299,N_11260);
xor U11643 (N_11643,N_11403,N_11370);
or U11644 (N_11644,N_11269,N_11303);
nor U11645 (N_11645,N_11332,N_11316);
nand U11646 (N_11646,N_11338,N_11260);
or U11647 (N_11647,N_11293,N_11475);
or U11648 (N_11648,N_11375,N_11326);
xor U11649 (N_11649,N_11424,N_11493);
and U11650 (N_11650,N_11343,N_11350);
or U11651 (N_11651,N_11454,N_11316);
nor U11652 (N_11652,N_11389,N_11305);
nor U11653 (N_11653,N_11261,N_11279);
or U11654 (N_11654,N_11441,N_11413);
or U11655 (N_11655,N_11360,N_11369);
or U11656 (N_11656,N_11472,N_11354);
or U11657 (N_11657,N_11364,N_11320);
and U11658 (N_11658,N_11439,N_11360);
nor U11659 (N_11659,N_11366,N_11294);
xnor U11660 (N_11660,N_11303,N_11328);
and U11661 (N_11661,N_11372,N_11312);
nor U11662 (N_11662,N_11372,N_11465);
xnor U11663 (N_11663,N_11423,N_11333);
or U11664 (N_11664,N_11468,N_11303);
or U11665 (N_11665,N_11350,N_11356);
and U11666 (N_11666,N_11408,N_11303);
or U11667 (N_11667,N_11469,N_11448);
xnor U11668 (N_11668,N_11480,N_11408);
nor U11669 (N_11669,N_11404,N_11291);
nor U11670 (N_11670,N_11499,N_11330);
xor U11671 (N_11671,N_11418,N_11403);
xor U11672 (N_11672,N_11399,N_11334);
nor U11673 (N_11673,N_11489,N_11303);
or U11674 (N_11674,N_11383,N_11413);
or U11675 (N_11675,N_11441,N_11416);
and U11676 (N_11676,N_11322,N_11256);
xor U11677 (N_11677,N_11406,N_11383);
nor U11678 (N_11678,N_11343,N_11456);
or U11679 (N_11679,N_11456,N_11403);
nor U11680 (N_11680,N_11302,N_11447);
or U11681 (N_11681,N_11303,N_11480);
xnor U11682 (N_11682,N_11412,N_11339);
xor U11683 (N_11683,N_11484,N_11268);
nand U11684 (N_11684,N_11479,N_11306);
or U11685 (N_11685,N_11490,N_11356);
or U11686 (N_11686,N_11342,N_11293);
xor U11687 (N_11687,N_11282,N_11294);
or U11688 (N_11688,N_11314,N_11251);
and U11689 (N_11689,N_11326,N_11457);
and U11690 (N_11690,N_11284,N_11408);
and U11691 (N_11691,N_11257,N_11300);
nand U11692 (N_11692,N_11263,N_11423);
or U11693 (N_11693,N_11280,N_11390);
or U11694 (N_11694,N_11384,N_11451);
and U11695 (N_11695,N_11403,N_11476);
nor U11696 (N_11696,N_11351,N_11284);
or U11697 (N_11697,N_11329,N_11302);
nand U11698 (N_11698,N_11258,N_11439);
nand U11699 (N_11699,N_11351,N_11261);
and U11700 (N_11700,N_11282,N_11471);
or U11701 (N_11701,N_11470,N_11321);
nor U11702 (N_11702,N_11351,N_11419);
or U11703 (N_11703,N_11304,N_11466);
xnor U11704 (N_11704,N_11452,N_11283);
nand U11705 (N_11705,N_11263,N_11342);
and U11706 (N_11706,N_11364,N_11279);
nor U11707 (N_11707,N_11367,N_11459);
and U11708 (N_11708,N_11445,N_11420);
or U11709 (N_11709,N_11406,N_11468);
nand U11710 (N_11710,N_11440,N_11267);
nor U11711 (N_11711,N_11322,N_11442);
nor U11712 (N_11712,N_11271,N_11320);
xor U11713 (N_11713,N_11448,N_11430);
or U11714 (N_11714,N_11374,N_11453);
nor U11715 (N_11715,N_11398,N_11480);
xor U11716 (N_11716,N_11263,N_11481);
or U11717 (N_11717,N_11251,N_11362);
xnor U11718 (N_11718,N_11344,N_11482);
nand U11719 (N_11719,N_11295,N_11473);
xnor U11720 (N_11720,N_11288,N_11483);
nand U11721 (N_11721,N_11484,N_11274);
or U11722 (N_11722,N_11279,N_11287);
or U11723 (N_11723,N_11430,N_11339);
and U11724 (N_11724,N_11316,N_11301);
or U11725 (N_11725,N_11265,N_11330);
xnor U11726 (N_11726,N_11377,N_11412);
nand U11727 (N_11727,N_11483,N_11335);
and U11728 (N_11728,N_11479,N_11387);
or U11729 (N_11729,N_11306,N_11312);
xnor U11730 (N_11730,N_11353,N_11285);
nand U11731 (N_11731,N_11482,N_11424);
xor U11732 (N_11732,N_11459,N_11257);
xor U11733 (N_11733,N_11297,N_11257);
nor U11734 (N_11734,N_11307,N_11483);
and U11735 (N_11735,N_11264,N_11338);
or U11736 (N_11736,N_11372,N_11306);
xnor U11737 (N_11737,N_11344,N_11279);
nand U11738 (N_11738,N_11252,N_11363);
and U11739 (N_11739,N_11376,N_11451);
or U11740 (N_11740,N_11315,N_11334);
or U11741 (N_11741,N_11459,N_11284);
or U11742 (N_11742,N_11304,N_11387);
xnor U11743 (N_11743,N_11358,N_11462);
nand U11744 (N_11744,N_11453,N_11399);
nand U11745 (N_11745,N_11274,N_11287);
and U11746 (N_11746,N_11475,N_11456);
nand U11747 (N_11747,N_11373,N_11477);
and U11748 (N_11748,N_11411,N_11346);
nor U11749 (N_11749,N_11333,N_11267);
xor U11750 (N_11750,N_11556,N_11692);
or U11751 (N_11751,N_11548,N_11673);
nor U11752 (N_11752,N_11735,N_11642);
nand U11753 (N_11753,N_11658,N_11524);
nand U11754 (N_11754,N_11716,N_11573);
nor U11755 (N_11755,N_11676,N_11688);
or U11756 (N_11756,N_11592,N_11696);
nand U11757 (N_11757,N_11677,N_11749);
xor U11758 (N_11758,N_11547,N_11501);
and U11759 (N_11759,N_11517,N_11715);
nand U11760 (N_11760,N_11578,N_11685);
nand U11761 (N_11761,N_11671,N_11509);
nor U11762 (N_11762,N_11670,N_11657);
and U11763 (N_11763,N_11510,N_11589);
or U11764 (N_11764,N_11698,N_11582);
nor U11765 (N_11765,N_11527,N_11544);
and U11766 (N_11766,N_11551,N_11745);
nor U11767 (N_11767,N_11615,N_11746);
and U11768 (N_11768,N_11555,N_11534);
xor U11769 (N_11769,N_11566,N_11744);
and U11770 (N_11770,N_11617,N_11726);
and U11771 (N_11771,N_11683,N_11631);
xnor U11772 (N_11772,N_11662,N_11741);
or U11773 (N_11773,N_11655,N_11733);
nand U11774 (N_11774,N_11740,N_11525);
nor U11775 (N_11775,N_11540,N_11559);
xnor U11776 (N_11776,N_11674,N_11633);
nand U11777 (N_11777,N_11554,N_11652);
and U11778 (N_11778,N_11634,N_11514);
or U11779 (N_11779,N_11624,N_11699);
nand U11780 (N_11780,N_11668,N_11546);
xor U11781 (N_11781,N_11706,N_11639);
or U11782 (N_11782,N_11563,N_11637);
xor U11783 (N_11783,N_11653,N_11586);
nand U11784 (N_11784,N_11585,N_11604);
nor U11785 (N_11785,N_11650,N_11616);
or U11786 (N_11786,N_11581,N_11576);
or U11787 (N_11787,N_11700,N_11720);
nand U11788 (N_11788,N_11601,N_11721);
nand U11789 (N_11789,N_11623,N_11538);
nand U11790 (N_11790,N_11602,N_11553);
or U11791 (N_11791,N_11739,N_11504);
or U11792 (N_11792,N_11607,N_11738);
xnor U11793 (N_11793,N_11507,N_11505);
or U11794 (N_11794,N_11622,N_11513);
and U11795 (N_11795,N_11728,N_11691);
nor U11796 (N_11796,N_11612,N_11545);
nor U11797 (N_11797,N_11725,N_11594);
and U11798 (N_11798,N_11552,N_11702);
xnor U11799 (N_11799,N_11568,N_11695);
xnor U11800 (N_11800,N_11729,N_11506);
or U11801 (N_11801,N_11532,N_11656);
nor U11802 (N_11802,N_11579,N_11610);
or U11803 (N_11803,N_11743,N_11742);
xnor U11804 (N_11804,N_11694,N_11647);
nor U11805 (N_11805,N_11533,N_11584);
nor U11806 (N_11806,N_11645,N_11502);
and U11807 (N_11807,N_11543,N_11710);
and U11808 (N_11808,N_11638,N_11669);
nor U11809 (N_11809,N_11675,N_11665);
and U11810 (N_11810,N_11569,N_11521);
or U11811 (N_11811,N_11666,N_11736);
xor U11812 (N_11812,N_11549,N_11709);
nand U11813 (N_11813,N_11664,N_11500);
and U11814 (N_11814,N_11574,N_11718);
or U11815 (N_11815,N_11714,N_11618);
nand U11816 (N_11816,N_11705,N_11723);
or U11817 (N_11817,N_11708,N_11678);
nor U11818 (N_11818,N_11711,N_11595);
xnor U11819 (N_11819,N_11689,N_11599);
nand U11820 (N_11820,N_11636,N_11680);
or U11821 (N_11821,N_11590,N_11606);
or U11822 (N_11822,N_11648,N_11522);
and U11823 (N_11823,N_11528,N_11518);
nor U11824 (N_11824,N_11719,N_11619);
xnor U11825 (N_11825,N_11603,N_11508);
and U11826 (N_11826,N_11580,N_11632);
nor U11827 (N_11827,N_11597,N_11526);
and U11828 (N_11828,N_11724,N_11596);
nand U11829 (N_11829,N_11747,N_11503);
nand U11830 (N_11830,N_11542,N_11535);
xor U11831 (N_11831,N_11593,N_11681);
nand U11832 (N_11832,N_11529,N_11613);
xnor U11833 (N_11833,N_11697,N_11516);
nor U11834 (N_11834,N_11734,N_11686);
nor U11835 (N_11835,N_11541,N_11651);
or U11836 (N_11836,N_11609,N_11727);
nor U11837 (N_11837,N_11560,N_11536);
and U11838 (N_11838,N_11539,N_11628);
nor U11839 (N_11839,N_11682,N_11512);
nand U11840 (N_11840,N_11591,N_11620);
or U11841 (N_11841,N_11731,N_11570);
nor U11842 (N_11842,N_11672,N_11565);
nand U11843 (N_11843,N_11667,N_11564);
xor U11844 (N_11844,N_11614,N_11713);
nor U11845 (N_11845,N_11635,N_11572);
nor U11846 (N_11846,N_11701,N_11660);
xor U11847 (N_11847,N_11608,N_11712);
nand U11848 (N_11848,N_11690,N_11703);
xnor U11849 (N_11849,N_11629,N_11707);
and U11850 (N_11850,N_11693,N_11679);
or U11851 (N_11851,N_11537,N_11625);
nand U11852 (N_11852,N_11626,N_11732);
xor U11853 (N_11853,N_11567,N_11588);
nand U11854 (N_11854,N_11611,N_11558);
nor U11855 (N_11855,N_11704,N_11644);
and U11856 (N_11856,N_11643,N_11519);
or U11857 (N_11857,N_11515,N_11621);
xnor U11858 (N_11858,N_11640,N_11730);
xor U11859 (N_11859,N_11661,N_11562);
nand U11860 (N_11860,N_11577,N_11659);
xor U11861 (N_11861,N_11684,N_11605);
nor U11862 (N_11862,N_11550,N_11687);
xor U11863 (N_11863,N_11531,N_11641);
nor U11864 (N_11864,N_11663,N_11649);
nand U11865 (N_11865,N_11561,N_11571);
and U11866 (N_11866,N_11737,N_11722);
xor U11867 (N_11867,N_11587,N_11630);
nand U11868 (N_11868,N_11748,N_11654);
or U11869 (N_11869,N_11598,N_11557);
or U11870 (N_11870,N_11520,N_11511);
or U11871 (N_11871,N_11627,N_11583);
xor U11872 (N_11872,N_11646,N_11523);
or U11873 (N_11873,N_11717,N_11575);
nor U11874 (N_11874,N_11530,N_11600);
or U11875 (N_11875,N_11748,N_11557);
and U11876 (N_11876,N_11685,N_11660);
or U11877 (N_11877,N_11584,N_11618);
nor U11878 (N_11878,N_11601,N_11652);
xor U11879 (N_11879,N_11573,N_11600);
or U11880 (N_11880,N_11709,N_11576);
or U11881 (N_11881,N_11683,N_11706);
nand U11882 (N_11882,N_11743,N_11701);
xnor U11883 (N_11883,N_11641,N_11606);
nor U11884 (N_11884,N_11730,N_11614);
nand U11885 (N_11885,N_11664,N_11720);
nand U11886 (N_11886,N_11575,N_11583);
or U11887 (N_11887,N_11738,N_11530);
xor U11888 (N_11888,N_11694,N_11719);
xnor U11889 (N_11889,N_11503,N_11604);
nand U11890 (N_11890,N_11747,N_11723);
and U11891 (N_11891,N_11594,N_11562);
xor U11892 (N_11892,N_11530,N_11613);
and U11893 (N_11893,N_11526,N_11679);
and U11894 (N_11894,N_11731,N_11739);
or U11895 (N_11895,N_11539,N_11699);
xor U11896 (N_11896,N_11696,N_11637);
nor U11897 (N_11897,N_11509,N_11690);
or U11898 (N_11898,N_11608,N_11593);
or U11899 (N_11899,N_11660,N_11688);
xnor U11900 (N_11900,N_11622,N_11564);
and U11901 (N_11901,N_11542,N_11513);
xor U11902 (N_11902,N_11713,N_11555);
and U11903 (N_11903,N_11682,N_11687);
nand U11904 (N_11904,N_11732,N_11630);
xnor U11905 (N_11905,N_11721,N_11610);
xnor U11906 (N_11906,N_11500,N_11653);
or U11907 (N_11907,N_11657,N_11559);
nand U11908 (N_11908,N_11647,N_11707);
and U11909 (N_11909,N_11620,N_11640);
and U11910 (N_11910,N_11703,N_11717);
nor U11911 (N_11911,N_11560,N_11625);
xnor U11912 (N_11912,N_11535,N_11630);
nand U11913 (N_11913,N_11561,N_11678);
xor U11914 (N_11914,N_11644,N_11597);
and U11915 (N_11915,N_11747,N_11615);
or U11916 (N_11916,N_11693,N_11574);
xor U11917 (N_11917,N_11514,N_11601);
and U11918 (N_11918,N_11618,N_11666);
xor U11919 (N_11919,N_11735,N_11624);
or U11920 (N_11920,N_11676,N_11569);
or U11921 (N_11921,N_11707,N_11706);
nor U11922 (N_11922,N_11701,N_11538);
xor U11923 (N_11923,N_11744,N_11668);
nand U11924 (N_11924,N_11556,N_11700);
or U11925 (N_11925,N_11534,N_11661);
nand U11926 (N_11926,N_11648,N_11744);
nor U11927 (N_11927,N_11688,N_11561);
nor U11928 (N_11928,N_11705,N_11606);
and U11929 (N_11929,N_11625,N_11616);
or U11930 (N_11930,N_11744,N_11706);
xnor U11931 (N_11931,N_11676,N_11504);
or U11932 (N_11932,N_11567,N_11744);
nand U11933 (N_11933,N_11681,N_11562);
and U11934 (N_11934,N_11696,N_11542);
and U11935 (N_11935,N_11628,N_11533);
and U11936 (N_11936,N_11706,N_11613);
nand U11937 (N_11937,N_11610,N_11674);
nor U11938 (N_11938,N_11748,N_11540);
nand U11939 (N_11939,N_11635,N_11731);
nand U11940 (N_11940,N_11591,N_11534);
nand U11941 (N_11941,N_11701,N_11516);
nor U11942 (N_11942,N_11749,N_11552);
and U11943 (N_11943,N_11666,N_11602);
nor U11944 (N_11944,N_11647,N_11573);
xor U11945 (N_11945,N_11646,N_11629);
nor U11946 (N_11946,N_11674,N_11727);
nand U11947 (N_11947,N_11710,N_11684);
or U11948 (N_11948,N_11672,N_11676);
nor U11949 (N_11949,N_11704,N_11676);
or U11950 (N_11950,N_11617,N_11519);
nand U11951 (N_11951,N_11560,N_11748);
or U11952 (N_11952,N_11519,N_11707);
and U11953 (N_11953,N_11718,N_11547);
or U11954 (N_11954,N_11650,N_11671);
nand U11955 (N_11955,N_11518,N_11592);
nor U11956 (N_11956,N_11507,N_11535);
xor U11957 (N_11957,N_11736,N_11521);
nand U11958 (N_11958,N_11504,N_11613);
nand U11959 (N_11959,N_11593,N_11626);
nor U11960 (N_11960,N_11562,N_11687);
and U11961 (N_11961,N_11576,N_11726);
xor U11962 (N_11962,N_11569,N_11724);
and U11963 (N_11963,N_11629,N_11729);
or U11964 (N_11964,N_11703,N_11585);
and U11965 (N_11965,N_11614,N_11710);
xor U11966 (N_11966,N_11665,N_11686);
and U11967 (N_11967,N_11647,N_11617);
nand U11968 (N_11968,N_11737,N_11543);
nor U11969 (N_11969,N_11602,N_11722);
and U11970 (N_11970,N_11509,N_11656);
xor U11971 (N_11971,N_11603,N_11533);
nand U11972 (N_11972,N_11691,N_11554);
xor U11973 (N_11973,N_11602,N_11711);
nor U11974 (N_11974,N_11737,N_11645);
xnor U11975 (N_11975,N_11600,N_11715);
nand U11976 (N_11976,N_11719,N_11576);
nand U11977 (N_11977,N_11660,N_11508);
or U11978 (N_11978,N_11595,N_11660);
or U11979 (N_11979,N_11677,N_11723);
xnor U11980 (N_11980,N_11561,N_11709);
xor U11981 (N_11981,N_11731,N_11692);
nor U11982 (N_11982,N_11638,N_11539);
and U11983 (N_11983,N_11688,N_11567);
and U11984 (N_11984,N_11674,N_11596);
xor U11985 (N_11985,N_11517,N_11712);
and U11986 (N_11986,N_11640,N_11687);
xnor U11987 (N_11987,N_11605,N_11690);
nand U11988 (N_11988,N_11565,N_11590);
xor U11989 (N_11989,N_11633,N_11516);
nand U11990 (N_11990,N_11646,N_11704);
nor U11991 (N_11991,N_11542,N_11628);
or U11992 (N_11992,N_11660,N_11501);
nor U11993 (N_11993,N_11685,N_11609);
nand U11994 (N_11994,N_11593,N_11546);
nor U11995 (N_11995,N_11724,N_11653);
xnor U11996 (N_11996,N_11612,N_11505);
or U11997 (N_11997,N_11644,N_11739);
nor U11998 (N_11998,N_11572,N_11655);
and U11999 (N_11999,N_11671,N_11552);
nor U12000 (N_12000,N_11976,N_11928);
and U12001 (N_12001,N_11968,N_11931);
nand U12002 (N_12002,N_11990,N_11960);
nand U12003 (N_12003,N_11998,N_11800);
nand U12004 (N_12004,N_11835,N_11818);
nor U12005 (N_12005,N_11858,N_11946);
xor U12006 (N_12006,N_11839,N_11861);
xnor U12007 (N_12007,N_11804,N_11954);
nand U12008 (N_12008,N_11788,N_11805);
nor U12009 (N_12009,N_11905,N_11843);
nor U12010 (N_12010,N_11810,N_11852);
nor U12011 (N_12011,N_11914,N_11897);
xor U12012 (N_12012,N_11876,N_11951);
nand U12013 (N_12013,N_11992,N_11957);
nor U12014 (N_12014,N_11791,N_11765);
or U12015 (N_12015,N_11823,N_11831);
xnor U12016 (N_12016,N_11873,N_11851);
nand U12017 (N_12017,N_11772,N_11838);
or U12018 (N_12018,N_11942,N_11774);
or U12019 (N_12019,N_11881,N_11987);
or U12020 (N_12020,N_11811,N_11926);
xor U12021 (N_12021,N_11803,N_11848);
or U12022 (N_12022,N_11939,N_11947);
xnor U12023 (N_12023,N_11763,N_11773);
xnor U12024 (N_12024,N_11904,N_11948);
or U12025 (N_12025,N_11920,N_11780);
and U12026 (N_12026,N_11909,N_11925);
nor U12027 (N_12027,N_11941,N_11880);
or U12028 (N_12028,N_11883,N_11991);
nand U12029 (N_12029,N_11761,N_11824);
xnor U12030 (N_12030,N_11967,N_11859);
nor U12031 (N_12031,N_11817,N_11875);
or U12032 (N_12032,N_11902,N_11844);
nor U12033 (N_12033,N_11979,N_11837);
nand U12034 (N_12034,N_11940,N_11955);
xor U12035 (N_12035,N_11985,N_11945);
and U12036 (N_12036,N_11972,N_11783);
nand U12037 (N_12037,N_11965,N_11898);
and U12038 (N_12038,N_11980,N_11950);
nand U12039 (N_12039,N_11785,N_11997);
nand U12040 (N_12040,N_11799,N_11860);
nand U12041 (N_12041,N_11878,N_11994);
nor U12042 (N_12042,N_11962,N_11892);
nand U12043 (N_12043,N_11944,N_11770);
nor U12044 (N_12044,N_11751,N_11934);
nand U12045 (N_12045,N_11850,N_11961);
and U12046 (N_12046,N_11777,N_11753);
nand U12047 (N_12047,N_11787,N_11993);
xnor U12048 (N_12048,N_11906,N_11958);
xnor U12049 (N_12049,N_11999,N_11879);
xnor U12050 (N_12050,N_11973,N_11932);
or U12051 (N_12051,N_11825,N_11866);
xor U12052 (N_12052,N_11807,N_11828);
and U12053 (N_12053,N_11927,N_11963);
xor U12054 (N_12054,N_11830,N_11755);
and U12055 (N_12055,N_11794,N_11943);
xnor U12056 (N_12056,N_11845,N_11863);
or U12057 (N_12057,N_11870,N_11907);
or U12058 (N_12058,N_11801,N_11933);
or U12059 (N_12059,N_11750,N_11857);
nand U12060 (N_12060,N_11891,N_11816);
nand U12061 (N_12061,N_11969,N_11856);
or U12062 (N_12062,N_11834,N_11793);
nand U12063 (N_12063,N_11759,N_11841);
nand U12064 (N_12064,N_11869,N_11929);
xor U12065 (N_12065,N_11923,N_11890);
nand U12066 (N_12066,N_11796,N_11970);
nor U12067 (N_12067,N_11918,N_11836);
xnor U12068 (N_12068,N_11952,N_11995);
nor U12069 (N_12069,N_11819,N_11978);
nand U12070 (N_12070,N_11762,N_11809);
or U12071 (N_12071,N_11986,N_11829);
xor U12072 (N_12072,N_11886,N_11826);
or U12073 (N_12073,N_11754,N_11867);
xnor U12074 (N_12074,N_11849,N_11853);
or U12075 (N_12075,N_11833,N_11862);
nand U12076 (N_12076,N_11885,N_11781);
nor U12077 (N_12077,N_11922,N_11908);
or U12078 (N_12078,N_11840,N_11893);
or U12079 (N_12079,N_11792,N_11956);
xor U12080 (N_12080,N_11903,N_11864);
nand U12081 (N_12081,N_11868,N_11822);
and U12082 (N_12082,N_11798,N_11789);
xnor U12083 (N_12083,N_11854,N_11784);
xnor U12084 (N_12084,N_11916,N_11764);
and U12085 (N_12085,N_11975,N_11821);
or U12086 (N_12086,N_11808,N_11775);
nand U12087 (N_12087,N_11981,N_11756);
or U12088 (N_12088,N_11971,N_11937);
xor U12089 (N_12089,N_11855,N_11894);
and U12090 (N_12090,N_11806,N_11769);
nor U12091 (N_12091,N_11884,N_11887);
xnor U12092 (N_12092,N_11779,N_11871);
or U12093 (N_12093,N_11896,N_11771);
nand U12094 (N_12094,N_11872,N_11786);
xnor U12095 (N_12095,N_11874,N_11911);
nand U12096 (N_12096,N_11984,N_11912);
nor U12097 (N_12097,N_11996,N_11752);
and U12098 (N_12098,N_11974,N_11767);
nor U12099 (N_12099,N_11813,N_11865);
xnor U12100 (N_12100,N_11949,N_11846);
nor U12101 (N_12101,N_11812,N_11847);
nand U12102 (N_12102,N_11758,N_11782);
xnor U12103 (N_12103,N_11921,N_11827);
or U12104 (N_12104,N_11988,N_11795);
nand U12105 (N_12105,N_11760,N_11953);
and U12106 (N_12106,N_11982,N_11778);
or U12107 (N_12107,N_11842,N_11889);
nand U12108 (N_12108,N_11901,N_11935);
nand U12109 (N_12109,N_11919,N_11938);
nor U12110 (N_12110,N_11977,N_11966);
or U12111 (N_12111,N_11820,N_11832);
or U12112 (N_12112,N_11900,N_11899);
and U12113 (N_12113,N_11888,N_11913);
xor U12114 (N_12114,N_11882,N_11814);
and U12115 (N_12115,N_11917,N_11910);
and U12116 (N_12116,N_11983,N_11815);
nand U12117 (N_12117,N_11924,N_11936);
nor U12118 (N_12118,N_11797,N_11989);
xor U12119 (N_12119,N_11959,N_11757);
xor U12120 (N_12120,N_11766,N_11895);
and U12121 (N_12121,N_11776,N_11768);
or U12122 (N_12122,N_11790,N_11964);
nor U12123 (N_12123,N_11802,N_11930);
and U12124 (N_12124,N_11877,N_11915);
nor U12125 (N_12125,N_11924,N_11947);
nand U12126 (N_12126,N_11823,N_11788);
nand U12127 (N_12127,N_11969,N_11824);
xnor U12128 (N_12128,N_11806,N_11950);
nor U12129 (N_12129,N_11872,N_11775);
nor U12130 (N_12130,N_11929,N_11783);
nand U12131 (N_12131,N_11933,N_11988);
nor U12132 (N_12132,N_11853,N_11847);
xnor U12133 (N_12133,N_11770,N_11822);
xnor U12134 (N_12134,N_11902,N_11750);
and U12135 (N_12135,N_11893,N_11823);
nor U12136 (N_12136,N_11867,N_11855);
and U12137 (N_12137,N_11988,N_11870);
or U12138 (N_12138,N_11775,N_11786);
xor U12139 (N_12139,N_11983,N_11792);
or U12140 (N_12140,N_11961,N_11819);
nand U12141 (N_12141,N_11936,N_11912);
nand U12142 (N_12142,N_11945,N_11953);
and U12143 (N_12143,N_11808,N_11877);
or U12144 (N_12144,N_11799,N_11833);
nand U12145 (N_12145,N_11921,N_11855);
nor U12146 (N_12146,N_11817,N_11771);
xnor U12147 (N_12147,N_11820,N_11960);
xor U12148 (N_12148,N_11873,N_11864);
nor U12149 (N_12149,N_11985,N_11951);
and U12150 (N_12150,N_11906,N_11895);
and U12151 (N_12151,N_11755,N_11928);
xnor U12152 (N_12152,N_11968,N_11934);
and U12153 (N_12153,N_11975,N_11802);
xnor U12154 (N_12154,N_11823,N_11811);
nor U12155 (N_12155,N_11793,N_11786);
and U12156 (N_12156,N_11859,N_11837);
nand U12157 (N_12157,N_11948,N_11805);
or U12158 (N_12158,N_11890,N_11866);
and U12159 (N_12159,N_11785,N_11750);
nor U12160 (N_12160,N_11902,N_11800);
nor U12161 (N_12161,N_11955,N_11792);
and U12162 (N_12162,N_11908,N_11918);
nor U12163 (N_12163,N_11872,N_11766);
nand U12164 (N_12164,N_11807,N_11857);
xnor U12165 (N_12165,N_11922,N_11913);
xor U12166 (N_12166,N_11851,N_11932);
or U12167 (N_12167,N_11964,N_11766);
nor U12168 (N_12168,N_11856,N_11975);
xnor U12169 (N_12169,N_11907,N_11989);
or U12170 (N_12170,N_11975,N_11868);
and U12171 (N_12171,N_11778,N_11808);
xnor U12172 (N_12172,N_11806,N_11793);
or U12173 (N_12173,N_11997,N_11762);
and U12174 (N_12174,N_11861,N_11831);
or U12175 (N_12175,N_11751,N_11964);
xor U12176 (N_12176,N_11810,N_11941);
nor U12177 (N_12177,N_11855,N_11817);
or U12178 (N_12178,N_11839,N_11963);
xor U12179 (N_12179,N_11847,N_11940);
nor U12180 (N_12180,N_11774,N_11935);
nor U12181 (N_12181,N_11939,N_11827);
and U12182 (N_12182,N_11883,N_11760);
nor U12183 (N_12183,N_11890,N_11761);
and U12184 (N_12184,N_11860,N_11820);
nand U12185 (N_12185,N_11987,N_11992);
xnor U12186 (N_12186,N_11934,N_11826);
nand U12187 (N_12187,N_11959,N_11921);
nand U12188 (N_12188,N_11764,N_11863);
nand U12189 (N_12189,N_11846,N_11820);
and U12190 (N_12190,N_11836,N_11757);
or U12191 (N_12191,N_11773,N_11870);
nor U12192 (N_12192,N_11813,N_11773);
nor U12193 (N_12193,N_11870,N_11834);
or U12194 (N_12194,N_11989,N_11960);
or U12195 (N_12195,N_11793,N_11935);
nand U12196 (N_12196,N_11927,N_11993);
and U12197 (N_12197,N_11788,N_11972);
xor U12198 (N_12198,N_11761,N_11822);
nand U12199 (N_12199,N_11902,N_11901);
nor U12200 (N_12200,N_11985,N_11879);
and U12201 (N_12201,N_11954,N_11853);
xor U12202 (N_12202,N_11908,N_11752);
or U12203 (N_12203,N_11786,N_11869);
or U12204 (N_12204,N_11948,N_11829);
nand U12205 (N_12205,N_11812,N_11771);
nand U12206 (N_12206,N_11903,N_11949);
nor U12207 (N_12207,N_11923,N_11830);
or U12208 (N_12208,N_11880,N_11954);
nand U12209 (N_12209,N_11792,N_11862);
xor U12210 (N_12210,N_11948,N_11847);
and U12211 (N_12211,N_11937,N_11780);
and U12212 (N_12212,N_11887,N_11969);
xor U12213 (N_12213,N_11829,N_11953);
and U12214 (N_12214,N_11767,N_11831);
nor U12215 (N_12215,N_11821,N_11926);
and U12216 (N_12216,N_11787,N_11862);
nor U12217 (N_12217,N_11867,N_11995);
or U12218 (N_12218,N_11807,N_11776);
nor U12219 (N_12219,N_11877,N_11896);
or U12220 (N_12220,N_11918,N_11784);
and U12221 (N_12221,N_11993,N_11971);
nand U12222 (N_12222,N_11849,N_11960);
nor U12223 (N_12223,N_11840,N_11816);
nand U12224 (N_12224,N_11814,N_11899);
nand U12225 (N_12225,N_11991,N_11766);
nand U12226 (N_12226,N_11892,N_11846);
xnor U12227 (N_12227,N_11804,N_11827);
nor U12228 (N_12228,N_11750,N_11961);
or U12229 (N_12229,N_11899,N_11824);
and U12230 (N_12230,N_11825,N_11936);
and U12231 (N_12231,N_11948,N_11962);
nor U12232 (N_12232,N_11751,N_11835);
nand U12233 (N_12233,N_11919,N_11908);
nor U12234 (N_12234,N_11908,N_11865);
nand U12235 (N_12235,N_11847,N_11858);
xor U12236 (N_12236,N_11914,N_11882);
or U12237 (N_12237,N_11831,N_11816);
xor U12238 (N_12238,N_11956,N_11844);
nor U12239 (N_12239,N_11773,N_11778);
nor U12240 (N_12240,N_11962,N_11970);
or U12241 (N_12241,N_11830,N_11985);
nand U12242 (N_12242,N_11986,N_11850);
nor U12243 (N_12243,N_11797,N_11770);
and U12244 (N_12244,N_11925,N_11821);
nor U12245 (N_12245,N_11979,N_11911);
and U12246 (N_12246,N_11855,N_11958);
xor U12247 (N_12247,N_11853,N_11822);
and U12248 (N_12248,N_11825,N_11811);
and U12249 (N_12249,N_11945,N_11947);
nand U12250 (N_12250,N_12245,N_12190);
or U12251 (N_12251,N_12220,N_12194);
nand U12252 (N_12252,N_12093,N_12149);
nor U12253 (N_12253,N_12001,N_12085);
or U12254 (N_12254,N_12117,N_12089);
nand U12255 (N_12255,N_12243,N_12121);
nand U12256 (N_12256,N_12102,N_12237);
xnor U12257 (N_12257,N_12208,N_12173);
or U12258 (N_12258,N_12054,N_12109);
nor U12259 (N_12259,N_12071,N_12123);
xor U12260 (N_12260,N_12185,N_12215);
xnor U12261 (N_12261,N_12087,N_12045);
nor U12262 (N_12262,N_12053,N_12193);
nor U12263 (N_12263,N_12078,N_12004);
or U12264 (N_12264,N_12161,N_12095);
or U12265 (N_12265,N_12118,N_12189);
xor U12266 (N_12266,N_12012,N_12120);
xnor U12267 (N_12267,N_12157,N_12076);
nand U12268 (N_12268,N_12113,N_12147);
xor U12269 (N_12269,N_12130,N_12209);
nand U12270 (N_12270,N_12204,N_12198);
or U12271 (N_12271,N_12009,N_12145);
nor U12272 (N_12272,N_12031,N_12143);
nor U12273 (N_12273,N_12063,N_12138);
or U12274 (N_12274,N_12154,N_12036);
nor U12275 (N_12275,N_12224,N_12119);
or U12276 (N_12276,N_12229,N_12035);
xnor U12277 (N_12277,N_12065,N_12034);
and U12278 (N_12278,N_12216,N_12195);
nor U12279 (N_12279,N_12210,N_12079);
nand U12280 (N_12280,N_12021,N_12013);
or U12281 (N_12281,N_12142,N_12181);
or U12282 (N_12282,N_12165,N_12169);
nand U12283 (N_12283,N_12104,N_12062);
or U12284 (N_12284,N_12170,N_12186);
or U12285 (N_12285,N_12082,N_12188);
xor U12286 (N_12286,N_12105,N_12177);
or U12287 (N_12287,N_12155,N_12151);
or U12288 (N_12288,N_12249,N_12213);
xor U12289 (N_12289,N_12112,N_12039);
nor U12290 (N_12290,N_12111,N_12074);
nor U12291 (N_12291,N_12097,N_12050);
nand U12292 (N_12292,N_12131,N_12196);
and U12293 (N_12293,N_12146,N_12152);
or U12294 (N_12294,N_12060,N_12038);
or U12295 (N_12295,N_12235,N_12160);
or U12296 (N_12296,N_12136,N_12172);
xor U12297 (N_12297,N_12137,N_12067);
xor U12298 (N_12298,N_12070,N_12128);
xor U12299 (N_12299,N_12217,N_12010);
xor U12300 (N_12300,N_12125,N_12134);
nor U12301 (N_12301,N_12099,N_12230);
xor U12302 (N_12302,N_12098,N_12005);
nand U12303 (N_12303,N_12066,N_12014);
xor U12304 (N_12304,N_12044,N_12207);
xnor U12305 (N_12305,N_12124,N_12094);
nor U12306 (N_12306,N_12025,N_12020);
or U12307 (N_12307,N_12200,N_12046);
nor U12308 (N_12308,N_12233,N_12096);
and U12309 (N_12309,N_12016,N_12000);
and U12310 (N_12310,N_12027,N_12234);
or U12311 (N_12311,N_12068,N_12159);
and U12312 (N_12312,N_12199,N_12212);
or U12313 (N_12313,N_12168,N_12037);
xnor U12314 (N_12314,N_12158,N_12006);
nand U12315 (N_12315,N_12144,N_12041);
xnor U12316 (N_12316,N_12248,N_12040);
and U12317 (N_12317,N_12205,N_12116);
nand U12318 (N_12318,N_12231,N_12103);
nand U12319 (N_12319,N_12226,N_12129);
and U12320 (N_12320,N_12140,N_12055);
and U12321 (N_12321,N_12197,N_12135);
and U12322 (N_12322,N_12156,N_12081);
nor U12323 (N_12323,N_12202,N_12176);
xnor U12324 (N_12324,N_12191,N_12242);
and U12325 (N_12325,N_12163,N_12122);
nor U12326 (N_12326,N_12174,N_12241);
or U12327 (N_12327,N_12227,N_12171);
xnor U12328 (N_12328,N_12222,N_12106);
and U12329 (N_12329,N_12030,N_12033);
nand U12330 (N_12330,N_12083,N_12127);
and U12331 (N_12331,N_12084,N_12043);
xnor U12332 (N_12332,N_12028,N_12192);
nor U12333 (N_12333,N_12064,N_12166);
xor U12334 (N_12334,N_12080,N_12139);
and U12335 (N_12335,N_12107,N_12141);
and U12336 (N_12336,N_12240,N_12100);
or U12337 (N_12337,N_12047,N_12187);
and U12338 (N_12338,N_12072,N_12164);
and U12339 (N_12339,N_12017,N_12225);
nor U12340 (N_12340,N_12075,N_12018);
nand U12341 (N_12341,N_12003,N_12029);
and U12342 (N_12342,N_12223,N_12178);
nor U12343 (N_12343,N_12101,N_12077);
xor U12344 (N_12344,N_12049,N_12180);
and U12345 (N_12345,N_12184,N_12232);
or U12346 (N_12346,N_12059,N_12182);
xnor U12347 (N_12347,N_12011,N_12048);
nand U12348 (N_12348,N_12115,N_12150);
xor U12349 (N_12349,N_12132,N_12008);
nor U12350 (N_12350,N_12214,N_12092);
xnor U12351 (N_12351,N_12022,N_12058);
xnor U12352 (N_12352,N_12024,N_12206);
nand U12353 (N_12353,N_12007,N_12179);
xor U12354 (N_12354,N_12175,N_12246);
and U12355 (N_12355,N_12073,N_12057);
and U12356 (N_12356,N_12239,N_12203);
or U12357 (N_12357,N_12148,N_12167);
and U12358 (N_12358,N_12026,N_12211);
nor U12359 (N_12359,N_12088,N_12218);
nand U12360 (N_12360,N_12023,N_12236);
xor U12361 (N_12361,N_12090,N_12052);
xor U12362 (N_12362,N_12162,N_12032);
xor U12363 (N_12363,N_12086,N_12183);
xnor U12364 (N_12364,N_12019,N_12244);
nor U12365 (N_12365,N_12114,N_12091);
and U12366 (N_12366,N_12153,N_12201);
nor U12367 (N_12367,N_12042,N_12069);
and U12368 (N_12368,N_12110,N_12219);
xnor U12369 (N_12369,N_12002,N_12108);
nand U12370 (N_12370,N_12126,N_12247);
nor U12371 (N_12371,N_12228,N_12238);
nand U12372 (N_12372,N_12051,N_12056);
and U12373 (N_12373,N_12015,N_12061);
xor U12374 (N_12374,N_12133,N_12221);
xnor U12375 (N_12375,N_12203,N_12142);
nand U12376 (N_12376,N_12016,N_12059);
or U12377 (N_12377,N_12136,N_12014);
and U12378 (N_12378,N_12070,N_12248);
and U12379 (N_12379,N_12224,N_12202);
xor U12380 (N_12380,N_12199,N_12236);
nand U12381 (N_12381,N_12049,N_12201);
nand U12382 (N_12382,N_12099,N_12054);
nor U12383 (N_12383,N_12098,N_12037);
or U12384 (N_12384,N_12205,N_12130);
or U12385 (N_12385,N_12017,N_12139);
nand U12386 (N_12386,N_12122,N_12180);
and U12387 (N_12387,N_12083,N_12085);
and U12388 (N_12388,N_12001,N_12168);
nor U12389 (N_12389,N_12172,N_12128);
nor U12390 (N_12390,N_12199,N_12055);
xnor U12391 (N_12391,N_12022,N_12108);
and U12392 (N_12392,N_12085,N_12158);
or U12393 (N_12393,N_12106,N_12022);
xor U12394 (N_12394,N_12135,N_12198);
nand U12395 (N_12395,N_12145,N_12205);
nand U12396 (N_12396,N_12002,N_12202);
xnor U12397 (N_12397,N_12183,N_12024);
nand U12398 (N_12398,N_12046,N_12115);
xnor U12399 (N_12399,N_12137,N_12114);
or U12400 (N_12400,N_12016,N_12151);
nor U12401 (N_12401,N_12188,N_12175);
nand U12402 (N_12402,N_12089,N_12169);
nor U12403 (N_12403,N_12003,N_12218);
and U12404 (N_12404,N_12194,N_12243);
or U12405 (N_12405,N_12119,N_12173);
nor U12406 (N_12406,N_12196,N_12245);
nor U12407 (N_12407,N_12004,N_12193);
xor U12408 (N_12408,N_12072,N_12135);
and U12409 (N_12409,N_12231,N_12151);
or U12410 (N_12410,N_12212,N_12043);
nor U12411 (N_12411,N_12057,N_12165);
nand U12412 (N_12412,N_12126,N_12224);
nor U12413 (N_12413,N_12042,N_12172);
xnor U12414 (N_12414,N_12129,N_12212);
and U12415 (N_12415,N_12222,N_12196);
or U12416 (N_12416,N_12090,N_12058);
xor U12417 (N_12417,N_12080,N_12056);
and U12418 (N_12418,N_12016,N_12185);
or U12419 (N_12419,N_12159,N_12087);
or U12420 (N_12420,N_12185,N_12118);
xnor U12421 (N_12421,N_12172,N_12062);
nor U12422 (N_12422,N_12125,N_12101);
and U12423 (N_12423,N_12226,N_12104);
nand U12424 (N_12424,N_12089,N_12161);
or U12425 (N_12425,N_12114,N_12026);
nor U12426 (N_12426,N_12114,N_12230);
or U12427 (N_12427,N_12020,N_12231);
xor U12428 (N_12428,N_12006,N_12245);
and U12429 (N_12429,N_12076,N_12115);
xor U12430 (N_12430,N_12122,N_12183);
or U12431 (N_12431,N_12178,N_12133);
nor U12432 (N_12432,N_12029,N_12091);
nor U12433 (N_12433,N_12149,N_12025);
nor U12434 (N_12434,N_12065,N_12141);
and U12435 (N_12435,N_12076,N_12033);
and U12436 (N_12436,N_12024,N_12012);
nand U12437 (N_12437,N_12021,N_12036);
nor U12438 (N_12438,N_12118,N_12188);
nand U12439 (N_12439,N_12239,N_12191);
nand U12440 (N_12440,N_12194,N_12071);
xor U12441 (N_12441,N_12063,N_12121);
and U12442 (N_12442,N_12123,N_12107);
or U12443 (N_12443,N_12025,N_12146);
xnor U12444 (N_12444,N_12224,N_12145);
or U12445 (N_12445,N_12006,N_12057);
and U12446 (N_12446,N_12138,N_12072);
nor U12447 (N_12447,N_12224,N_12097);
nor U12448 (N_12448,N_12019,N_12071);
nand U12449 (N_12449,N_12117,N_12240);
nand U12450 (N_12450,N_12053,N_12146);
nand U12451 (N_12451,N_12059,N_12121);
or U12452 (N_12452,N_12079,N_12246);
and U12453 (N_12453,N_12000,N_12176);
xor U12454 (N_12454,N_12028,N_12132);
xnor U12455 (N_12455,N_12248,N_12111);
nand U12456 (N_12456,N_12095,N_12093);
or U12457 (N_12457,N_12102,N_12001);
nor U12458 (N_12458,N_12160,N_12098);
or U12459 (N_12459,N_12008,N_12012);
xnor U12460 (N_12460,N_12201,N_12182);
or U12461 (N_12461,N_12106,N_12010);
nor U12462 (N_12462,N_12238,N_12068);
nand U12463 (N_12463,N_12097,N_12116);
nor U12464 (N_12464,N_12163,N_12101);
nor U12465 (N_12465,N_12045,N_12232);
or U12466 (N_12466,N_12122,N_12243);
xor U12467 (N_12467,N_12245,N_12110);
xnor U12468 (N_12468,N_12134,N_12242);
xnor U12469 (N_12469,N_12132,N_12229);
nand U12470 (N_12470,N_12082,N_12056);
and U12471 (N_12471,N_12015,N_12145);
and U12472 (N_12472,N_12231,N_12081);
xnor U12473 (N_12473,N_12051,N_12207);
or U12474 (N_12474,N_12214,N_12178);
or U12475 (N_12475,N_12158,N_12012);
nor U12476 (N_12476,N_12037,N_12018);
nor U12477 (N_12477,N_12101,N_12222);
or U12478 (N_12478,N_12130,N_12193);
xnor U12479 (N_12479,N_12026,N_12083);
and U12480 (N_12480,N_12134,N_12143);
xnor U12481 (N_12481,N_12083,N_12153);
nand U12482 (N_12482,N_12210,N_12063);
xnor U12483 (N_12483,N_12036,N_12145);
nand U12484 (N_12484,N_12055,N_12235);
xnor U12485 (N_12485,N_12166,N_12084);
xnor U12486 (N_12486,N_12035,N_12153);
nor U12487 (N_12487,N_12223,N_12119);
xnor U12488 (N_12488,N_12194,N_12209);
and U12489 (N_12489,N_12246,N_12112);
and U12490 (N_12490,N_12051,N_12205);
or U12491 (N_12491,N_12121,N_12244);
and U12492 (N_12492,N_12061,N_12142);
nand U12493 (N_12493,N_12019,N_12120);
nor U12494 (N_12494,N_12052,N_12225);
or U12495 (N_12495,N_12176,N_12214);
nor U12496 (N_12496,N_12153,N_12080);
nand U12497 (N_12497,N_12111,N_12078);
nand U12498 (N_12498,N_12016,N_12152);
nor U12499 (N_12499,N_12101,N_12083);
nand U12500 (N_12500,N_12277,N_12278);
nor U12501 (N_12501,N_12474,N_12316);
nor U12502 (N_12502,N_12310,N_12482);
nor U12503 (N_12503,N_12335,N_12375);
nor U12504 (N_12504,N_12493,N_12410);
nor U12505 (N_12505,N_12487,N_12328);
nand U12506 (N_12506,N_12450,N_12349);
and U12507 (N_12507,N_12284,N_12368);
xor U12508 (N_12508,N_12313,N_12299);
xnor U12509 (N_12509,N_12398,N_12281);
nor U12510 (N_12510,N_12403,N_12257);
nand U12511 (N_12511,N_12466,N_12460);
nor U12512 (N_12512,N_12388,N_12418);
and U12513 (N_12513,N_12414,N_12424);
nand U12514 (N_12514,N_12434,N_12304);
xor U12515 (N_12515,N_12491,N_12321);
xor U12516 (N_12516,N_12295,N_12290);
nor U12517 (N_12517,N_12324,N_12279);
nand U12518 (N_12518,N_12417,N_12308);
and U12519 (N_12519,N_12261,N_12339);
and U12520 (N_12520,N_12400,N_12371);
xnor U12521 (N_12521,N_12392,N_12325);
or U12522 (N_12522,N_12486,N_12382);
xor U12523 (N_12523,N_12262,N_12370);
nand U12524 (N_12524,N_12383,N_12444);
and U12525 (N_12525,N_12285,N_12344);
or U12526 (N_12526,N_12471,N_12397);
and U12527 (N_12527,N_12301,N_12439);
nor U12528 (N_12528,N_12399,N_12468);
nor U12529 (N_12529,N_12440,N_12459);
nand U12530 (N_12530,N_12276,N_12307);
xor U12531 (N_12531,N_12275,N_12435);
or U12532 (N_12532,N_12427,N_12391);
xnor U12533 (N_12533,N_12350,N_12378);
nand U12534 (N_12534,N_12258,N_12489);
xor U12535 (N_12535,N_12413,N_12393);
nand U12536 (N_12536,N_12374,N_12320);
xor U12537 (N_12537,N_12409,N_12360);
xnor U12538 (N_12538,N_12488,N_12467);
xor U12539 (N_12539,N_12300,N_12351);
xnor U12540 (N_12540,N_12494,N_12363);
or U12541 (N_12541,N_12446,N_12454);
or U12542 (N_12542,N_12408,N_12411);
xnor U12543 (N_12543,N_12379,N_12340);
and U12544 (N_12544,N_12437,N_12296);
nand U12545 (N_12545,N_12390,N_12432);
xor U12546 (N_12546,N_12469,N_12356);
nand U12547 (N_12547,N_12254,N_12260);
xor U12548 (N_12548,N_12481,N_12354);
and U12549 (N_12549,N_12438,N_12425);
nand U12550 (N_12550,N_12298,N_12449);
nor U12551 (N_12551,N_12426,N_12365);
or U12552 (N_12552,N_12431,N_12381);
nor U12553 (N_12553,N_12452,N_12401);
nand U12554 (N_12554,N_12266,N_12362);
xor U12555 (N_12555,N_12259,N_12492);
or U12556 (N_12556,N_12280,N_12480);
and U12557 (N_12557,N_12359,N_12343);
and U12558 (N_12558,N_12376,N_12357);
nor U12559 (N_12559,N_12463,N_12263);
or U12560 (N_12560,N_12282,N_12289);
and U12561 (N_12561,N_12421,N_12317);
xnor U12562 (N_12562,N_12384,N_12334);
xnor U12563 (N_12563,N_12380,N_12430);
xnor U12564 (N_12564,N_12485,N_12457);
nand U12565 (N_12565,N_12297,N_12332);
or U12566 (N_12566,N_12353,N_12346);
nor U12567 (N_12567,N_12271,N_12287);
nand U12568 (N_12568,N_12322,N_12419);
xor U12569 (N_12569,N_12473,N_12273);
or U12570 (N_12570,N_12477,N_12270);
and U12571 (N_12571,N_12367,N_12406);
or U12572 (N_12572,N_12269,N_12436);
and U12573 (N_12573,N_12445,N_12288);
nand U12574 (N_12574,N_12472,N_12373);
or U12575 (N_12575,N_12441,N_12336);
nor U12576 (N_12576,N_12323,N_12361);
and U12577 (N_12577,N_12420,N_12305);
and U12578 (N_12578,N_12448,N_12293);
xor U12579 (N_12579,N_12291,N_12302);
xor U12580 (N_12580,N_12267,N_12428);
and U12581 (N_12581,N_12462,N_12451);
or U12582 (N_12582,N_12333,N_12264);
and U12583 (N_12583,N_12348,N_12352);
nor U12584 (N_12584,N_12318,N_12498);
xnor U12585 (N_12585,N_12345,N_12475);
and U12586 (N_12586,N_12478,N_12395);
nand U12587 (N_12587,N_12465,N_12292);
and U12588 (N_12588,N_12455,N_12252);
xnor U12589 (N_12589,N_12274,N_12326);
or U12590 (N_12590,N_12364,N_12294);
nand U12591 (N_12591,N_12484,N_12433);
and U12592 (N_12592,N_12256,N_12355);
xnor U12593 (N_12593,N_12423,N_12458);
xnor U12594 (N_12594,N_12312,N_12347);
nor U12595 (N_12595,N_12404,N_12422);
and U12596 (N_12596,N_12309,N_12464);
or U12597 (N_12597,N_12314,N_12396);
and U12598 (N_12598,N_12315,N_12272);
and U12599 (N_12599,N_12470,N_12415);
or U12600 (N_12600,N_12255,N_12453);
xnor U12601 (N_12601,N_12442,N_12483);
and U12602 (N_12602,N_12416,N_12496);
xor U12603 (N_12603,N_12495,N_12461);
nor U12604 (N_12604,N_12394,N_12479);
nand U12605 (N_12605,N_12265,N_12330);
or U12606 (N_12606,N_12377,N_12329);
and U12607 (N_12607,N_12476,N_12286);
nor U12608 (N_12608,N_12319,N_12303);
or U12609 (N_12609,N_12447,N_12372);
or U12610 (N_12610,N_12253,N_12402);
xor U12611 (N_12611,N_12497,N_12358);
nor U12612 (N_12612,N_12311,N_12456);
or U12613 (N_12613,N_12386,N_12443);
xor U12614 (N_12614,N_12331,N_12306);
xnor U12615 (N_12615,N_12412,N_12389);
nand U12616 (N_12616,N_12429,N_12342);
nor U12617 (N_12617,N_12341,N_12327);
xor U12618 (N_12618,N_12337,N_12369);
xnor U12619 (N_12619,N_12387,N_12268);
xnor U12620 (N_12620,N_12366,N_12490);
nor U12621 (N_12621,N_12407,N_12338);
or U12622 (N_12622,N_12251,N_12250);
nor U12623 (N_12623,N_12283,N_12499);
and U12624 (N_12624,N_12405,N_12385);
nor U12625 (N_12625,N_12339,N_12473);
or U12626 (N_12626,N_12425,N_12439);
or U12627 (N_12627,N_12429,N_12431);
or U12628 (N_12628,N_12468,N_12424);
or U12629 (N_12629,N_12470,N_12455);
nand U12630 (N_12630,N_12272,N_12371);
nor U12631 (N_12631,N_12373,N_12329);
xnor U12632 (N_12632,N_12469,N_12437);
or U12633 (N_12633,N_12494,N_12482);
and U12634 (N_12634,N_12265,N_12461);
nand U12635 (N_12635,N_12375,N_12343);
and U12636 (N_12636,N_12300,N_12373);
nand U12637 (N_12637,N_12362,N_12259);
xor U12638 (N_12638,N_12498,N_12428);
nand U12639 (N_12639,N_12348,N_12345);
and U12640 (N_12640,N_12437,N_12329);
nor U12641 (N_12641,N_12342,N_12267);
xnor U12642 (N_12642,N_12390,N_12426);
or U12643 (N_12643,N_12367,N_12359);
nor U12644 (N_12644,N_12338,N_12370);
and U12645 (N_12645,N_12480,N_12466);
and U12646 (N_12646,N_12260,N_12386);
nand U12647 (N_12647,N_12312,N_12380);
and U12648 (N_12648,N_12380,N_12402);
and U12649 (N_12649,N_12335,N_12492);
and U12650 (N_12650,N_12267,N_12251);
or U12651 (N_12651,N_12499,N_12490);
nor U12652 (N_12652,N_12262,N_12440);
and U12653 (N_12653,N_12436,N_12261);
and U12654 (N_12654,N_12469,N_12273);
and U12655 (N_12655,N_12354,N_12329);
or U12656 (N_12656,N_12341,N_12435);
nor U12657 (N_12657,N_12408,N_12322);
xnor U12658 (N_12658,N_12464,N_12314);
nand U12659 (N_12659,N_12340,N_12281);
or U12660 (N_12660,N_12344,N_12497);
xor U12661 (N_12661,N_12499,N_12427);
nor U12662 (N_12662,N_12330,N_12357);
nand U12663 (N_12663,N_12298,N_12339);
or U12664 (N_12664,N_12432,N_12275);
nor U12665 (N_12665,N_12449,N_12338);
or U12666 (N_12666,N_12343,N_12422);
xor U12667 (N_12667,N_12268,N_12435);
nor U12668 (N_12668,N_12400,N_12290);
and U12669 (N_12669,N_12365,N_12484);
nor U12670 (N_12670,N_12252,N_12383);
nand U12671 (N_12671,N_12458,N_12451);
xor U12672 (N_12672,N_12253,N_12311);
or U12673 (N_12673,N_12408,N_12297);
and U12674 (N_12674,N_12328,N_12443);
or U12675 (N_12675,N_12309,N_12287);
nor U12676 (N_12676,N_12287,N_12386);
or U12677 (N_12677,N_12474,N_12265);
or U12678 (N_12678,N_12293,N_12325);
xnor U12679 (N_12679,N_12365,N_12433);
or U12680 (N_12680,N_12369,N_12269);
or U12681 (N_12681,N_12374,N_12343);
nor U12682 (N_12682,N_12432,N_12324);
nor U12683 (N_12683,N_12322,N_12290);
or U12684 (N_12684,N_12332,N_12418);
or U12685 (N_12685,N_12309,N_12441);
nand U12686 (N_12686,N_12325,N_12481);
nor U12687 (N_12687,N_12261,N_12444);
or U12688 (N_12688,N_12307,N_12454);
xor U12689 (N_12689,N_12253,N_12332);
and U12690 (N_12690,N_12446,N_12253);
xnor U12691 (N_12691,N_12260,N_12414);
xor U12692 (N_12692,N_12443,N_12424);
and U12693 (N_12693,N_12310,N_12417);
nand U12694 (N_12694,N_12305,N_12470);
or U12695 (N_12695,N_12448,N_12426);
xor U12696 (N_12696,N_12271,N_12474);
or U12697 (N_12697,N_12494,N_12486);
or U12698 (N_12698,N_12344,N_12316);
nand U12699 (N_12699,N_12374,N_12288);
nand U12700 (N_12700,N_12367,N_12494);
xnor U12701 (N_12701,N_12384,N_12495);
xnor U12702 (N_12702,N_12387,N_12453);
xnor U12703 (N_12703,N_12400,N_12359);
nor U12704 (N_12704,N_12499,N_12318);
xor U12705 (N_12705,N_12351,N_12299);
and U12706 (N_12706,N_12404,N_12398);
or U12707 (N_12707,N_12383,N_12404);
or U12708 (N_12708,N_12439,N_12436);
nor U12709 (N_12709,N_12340,N_12286);
nand U12710 (N_12710,N_12390,N_12308);
xor U12711 (N_12711,N_12444,N_12301);
or U12712 (N_12712,N_12473,N_12424);
nand U12713 (N_12713,N_12342,N_12337);
nand U12714 (N_12714,N_12265,N_12266);
or U12715 (N_12715,N_12489,N_12388);
xor U12716 (N_12716,N_12359,N_12487);
and U12717 (N_12717,N_12497,N_12416);
nor U12718 (N_12718,N_12455,N_12350);
nor U12719 (N_12719,N_12395,N_12250);
nor U12720 (N_12720,N_12366,N_12462);
nand U12721 (N_12721,N_12437,N_12353);
nand U12722 (N_12722,N_12473,N_12324);
xnor U12723 (N_12723,N_12430,N_12410);
nor U12724 (N_12724,N_12498,N_12471);
and U12725 (N_12725,N_12481,N_12433);
nor U12726 (N_12726,N_12481,N_12437);
nor U12727 (N_12727,N_12492,N_12489);
nor U12728 (N_12728,N_12461,N_12485);
and U12729 (N_12729,N_12299,N_12338);
nor U12730 (N_12730,N_12468,N_12330);
and U12731 (N_12731,N_12253,N_12251);
nand U12732 (N_12732,N_12268,N_12395);
and U12733 (N_12733,N_12350,N_12453);
nand U12734 (N_12734,N_12290,N_12470);
xnor U12735 (N_12735,N_12396,N_12274);
and U12736 (N_12736,N_12277,N_12413);
and U12737 (N_12737,N_12473,N_12362);
xnor U12738 (N_12738,N_12359,N_12309);
or U12739 (N_12739,N_12273,N_12284);
nor U12740 (N_12740,N_12285,N_12476);
xor U12741 (N_12741,N_12481,N_12284);
or U12742 (N_12742,N_12258,N_12351);
or U12743 (N_12743,N_12379,N_12462);
xor U12744 (N_12744,N_12270,N_12451);
or U12745 (N_12745,N_12391,N_12466);
nor U12746 (N_12746,N_12460,N_12497);
or U12747 (N_12747,N_12291,N_12411);
and U12748 (N_12748,N_12355,N_12266);
nand U12749 (N_12749,N_12306,N_12467);
nor U12750 (N_12750,N_12591,N_12548);
nand U12751 (N_12751,N_12647,N_12612);
xnor U12752 (N_12752,N_12708,N_12524);
or U12753 (N_12753,N_12570,N_12707);
and U12754 (N_12754,N_12597,N_12526);
nor U12755 (N_12755,N_12571,N_12628);
nand U12756 (N_12756,N_12550,N_12648);
and U12757 (N_12757,N_12692,N_12511);
or U12758 (N_12758,N_12711,N_12653);
xnor U12759 (N_12759,N_12660,N_12603);
nor U12760 (N_12760,N_12697,N_12616);
xnor U12761 (N_12761,N_12741,N_12541);
nand U12762 (N_12762,N_12639,N_12558);
or U12763 (N_12763,N_12572,N_12677);
nand U12764 (N_12764,N_12670,N_12688);
xnor U12765 (N_12765,N_12720,N_12632);
nand U12766 (N_12766,N_12503,N_12587);
or U12767 (N_12767,N_12536,N_12540);
and U12768 (N_12768,N_12557,N_12695);
xor U12769 (N_12769,N_12620,N_12615);
or U12770 (N_12770,N_12694,N_12722);
or U12771 (N_12771,N_12740,N_12748);
and U12772 (N_12772,N_12621,N_12568);
and U12773 (N_12773,N_12631,N_12714);
nand U12774 (N_12774,N_12658,N_12641);
nor U12775 (N_12775,N_12627,N_12706);
and U12776 (N_12776,N_12516,N_12687);
nor U12777 (N_12777,N_12517,N_12691);
nand U12778 (N_12778,N_12736,N_12640);
and U12779 (N_12779,N_12574,N_12683);
and U12780 (N_12780,N_12651,N_12563);
and U12781 (N_12781,N_12607,N_12745);
xor U12782 (N_12782,N_12732,N_12680);
nor U12783 (N_12783,N_12674,N_12724);
nand U12784 (N_12784,N_12643,N_12525);
and U12785 (N_12785,N_12601,N_12617);
nand U12786 (N_12786,N_12712,N_12522);
xor U12787 (N_12787,N_12638,N_12567);
and U12788 (N_12788,N_12537,N_12730);
and U12789 (N_12789,N_12704,N_12595);
or U12790 (N_12790,N_12609,N_12645);
xnor U12791 (N_12791,N_12553,N_12593);
nor U12792 (N_12792,N_12657,N_12698);
nand U12793 (N_12793,N_12713,N_12676);
nand U12794 (N_12794,N_12715,N_12555);
xnor U12795 (N_12795,N_12596,N_12652);
xor U12796 (N_12796,N_12738,N_12661);
or U12797 (N_12797,N_12605,N_12725);
and U12798 (N_12798,N_12678,N_12733);
nand U12799 (N_12799,N_12510,N_12662);
and U12800 (N_12800,N_12659,N_12644);
xor U12801 (N_12801,N_12635,N_12565);
xor U12802 (N_12802,N_12646,N_12602);
nor U12803 (N_12803,N_12686,N_12531);
and U12804 (N_12804,N_12669,N_12577);
xnor U12805 (N_12805,N_12664,N_12727);
and U12806 (N_12806,N_12671,N_12513);
nand U12807 (N_12807,N_12705,N_12668);
nand U12808 (N_12808,N_12501,N_12505);
nor U12809 (N_12809,N_12560,N_12625);
nor U12810 (N_12810,N_12578,N_12527);
nor U12811 (N_12811,N_12518,N_12598);
nor U12812 (N_12812,N_12702,N_12693);
nand U12813 (N_12813,N_12729,N_12533);
or U12814 (N_12814,N_12504,N_12746);
xor U12815 (N_12815,N_12543,N_12690);
and U12816 (N_12816,N_12590,N_12588);
or U12817 (N_12817,N_12728,N_12564);
and U12818 (N_12818,N_12675,N_12703);
nand U12819 (N_12819,N_12608,N_12726);
nand U12820 (N_12820,N_12606,N_12610);
and U12821 (N_12821,N_12542,N_12585);
xor U12822 (N_12822,N_12656,N_12731);
nand U12823 (N_12823,N_12684,N_12559);
and U12824 (N_12824,N_12681,N_12519);
or U12825 (N_12825,N_12534,N_12636);
or U12826 (N_12826,N_12600,N_12619);
nand U12827 (N_12827,N_12624,N_12663);
or U12828 (N_12828,N_12575,N_12583);
nor U12829 (N_12829,N_12744,N_12586);
xnor U12830 (N_12830,N_12637,N_12584);
nand U12831 (N_12831,N_12710,N_12515);
nor U12832 (N_12832,N_12665,N_12734);
nand U12833 (N_12833,N_12573,N_12580);
nor U12834 (N_12834,N_12672,N_12629);
nor U12835 (N_12835,N_12654,N_12523);
xor U12836 (N_12836,N_12554,N_12633);
or U12837 (N_12837,N_12514,N_12630);
nand U12838 (N_12838,N_12599,N_12545);
xor U12839 (N_12839,N_12626,N_12581);
and U12840 (N_12840,N_12649,N_12569);
xor U12841 (N_12841,N_12502,N_12614);
or U12842 (N_12842,N_12561,N_12666);
nand U12843 (N_12843,N_12579,N_12566);
nor U12844 (N_12844,N_12592,N_12549);
xor U12845 (N_12845,N_12589,N_12655);
or U12846 (N_12846,N_12512,N_12700);
or U12847 (N_12847,N_12622,N_12749);
or U12848 (N_12848,N_12613,N_12538);
xor U12849 (N_12849,N_12667,N_12539);
xnor U12850 (N_12850,N_12546,N_12642);
nand U12851 (N_12851,N_12650,N_12735);
xor U12852 (N_12852,N_12506,N_12618);
xor U12853 (N_12853,N_12737,N_12500);
nor U12854 (N_12854,N_12582,N_12719);
xor U12855 (N_12855,N_12747,N_12528);
and U12856 (N_12856,N_12521,N_12556);
xor U12857 (N_12857,N_12551,N_12716);
and U12858 (N_12858,N_12679,N_12717);
xor U12859 (N_12859,N_12594,N_12743);
xnor U12860 (N_12860,N_12699,N_12552);
or U12861 (N_12861,N_12718,N_12508);
xnor U12862 (N_12862,N_12689,N_12682);
nor U12863 (N_12863,N_12723,N_12544);
xnor U12864 (N_12864,N_12685,N_12739);
or U12865 (N_12865,N_12547,N_12634);
or U12866 (N_12866,N_12562,N_12709);
or U12867 (N_12867,N_12623,N_12532);
xor U12868 (N_12868,N_12696,N_12535);
nor U12869 (N_12869,N_12520,N_12611);
xor U12870 (N_12870,N_12701,N_12529);
and U12871 (N_12871,N_12507,N_12673);
xnor U12872 (N_12872,N_12509,N_12576);
xnor U12873 (N_12873,N_12530,N_12604);
or U12874 (N_12874,N_12742,N_12721);
xor U12875 (N_12875,N_12739,N_12728);
or U12876 (N_12876,N_12592,N_12684);
or U12877 (N_12877,N_12696,N_12531);
nor U12878 (N_12878,N_12638,N_12584);
or U12879 (N_12879,N_12625,N_12690);
and U12880 (N_12880,N_12550,N_12749);
xnor U12881 (N_12881,N_12627,N_12544);
nand U12882 (N_12882,N_12609,N_12716);
nor U12883 (N_12883,N_12738,N_12507);
or U12884 (N_12884,N_12713,N_12545);
nor U12885 (N_12885,N_12503,N_12545);
xor U12886 (N_12886,N_12590,N_12675);
xor U12887 (N_12887,N_12659,N_12575);
nor U12888 (N_12888,N_12565,N_12717);
or U12889 (N_12889,N_12661,N_12534);
nand U12890 (N_12890,N_12593,N_12508);
nor U12891 (N_12891,N_12716,N_12550);
or U12892 (N_12892,N_12672,N_12620);
xnor U12893 (N_12893,N_12729,N_12513);
nand U12894 (N_12894,N_12578,N_12642);
nor U12895 (N_12895,N_12572,N_12508);
xnor U12896 (N_12896,N_12718,N_12528);
xnor U12897 (N_12897,N_12623,N_12667);
nor U12898 (N_12898,N_12566,N_12600);
xor U12899 (N_12899,N_12719,N_12740);
or U12900 (N_12900,N_12663,N_12733);
and U12901 (N_12901,N_12737,N_12675);
xnor U12902 (N_12902,N_12509,N_12506);
nor U12903 (N_12903,N_12709,N_12636);
xor U12904 (N_12904,N_12699,N_12635);
nand U12905 (N_12905,N_12703,N_12603);
and U12906 (N_12906,N_12545,N_12649);
nor U12907 (N_12907,N_12748,N_12559);
and U12908 (N_12908,N_12550,N_12530);
or U12909 (N_12909,N_12572,N_12611);
xnor U12910 (N_12910,N_12619,N_12655);
and U12911 (N_12911,N_12630,N_12589);
or U12912 (N_12912,N_12509,N_12529);
and U12913 (N_12913,N_12726,N_12688);
nand U12914 (N_12914,N_12521,N_12592);
xor U12915 (N_12915,N_12677,N_12536);
nor U12916 (N_12916,N_12625,N_12656);
or U12917 (N_12917,N_12546,N_12573);
and U12918 (N_12918,N_12671,N_12530);
nor U12919 (N_12919,N_12713,N_12536);
xor U12920 (N_12920,N_12731,N_12507);
xor U12921 (N_12921,N_12691,N_12717);
nand U12922 (N_12922,N_12622,N_12678);
and U12923 (N_12923,N_12633,N_12564);
or U12924 (N_12924,N_12684,N_12544);
or U12925 (N_12925,N_12737,N_12648);
and U12926 (N_12926,N_12738,N_12591);
or U12927 (N_12927,N_12559,N_12711);
or U12928 (N_12928,N_12585,N_12699);
xnor U12929 (N_12929,N_12734,N_12741);
and U12930 (N_12930,N_12683,N_12635);
nor U12931 (N_12931,N_12729,N_12538);
or U12932 (N_12932,N_12508,N_12539);
xnor U12933 (N_12933,N_12666,N_12575);
and U12934 (N_12934,N_12557,N_12535);
or U12935 (N_12935,N_12718,N_12500);
nand U12936 (N_12936,N_12589,N_12638);
xnor U12937 (N_12937,N_12575,N_12573);
nand U12938 (N_12938,N_12720,N_12715);
and U12939 (N_12939,N_12648,N_12740);
or U12940 (N_12940,N_12591,N_12578);
and U12941 (N_12941,N_12525,N_12659);
xor U12942 (N_12942,N_12716,N_12668);
or U12943 (N_12943,N_12682,N_12728);
or U12944 (N_12944,N_12635,N_12706);
or U12945 (N_12945,N_12605,N_12607);
nand U12946 (N_12946,N_12626,N_12587);
or U12947 (N_12947,N_12743,N_12551);
xnor U12948 (N_12948,N_12503,N_12722);
xnor U12949 (N_12949,N_12540,N_12585);
xnor U12950 (N_12950,N_12667,N_12742);
and U12951 (N_12951,N_12723,N_12532);
and U12952 (N_12952,N_12607,N_12691);
nor U12953 (N_12953,N_12520,N_12534);
nand U12954 (N_12954,N_12523,N_12501);
or U12955 (N_12955,N_12747,N_12640);
xnor U12956 (N_12956,N_12625,N_12574);
xnor U12957 (N_12957,N_12516,N_12608);
or U12958 (N_12958,N_12562,N_12688);
nor U12959 (N_12959,N_12696,N_12729);
nor U12960 (N_12960,N_12525,N_12717);
or U12961 (N_12961,N_12635,N_12572);
xor U12962 (N_12962,N_12521,N_12598);
nor U12963 (N_12963,N_12563,N_12630);
nor U12964 (N_12964,N_12716,N_12616);
xnor U12965 (N_12965,N_12575,N_12610);
nor U12966 (N_12966,N_12734,N_12573);
nand U12967 (N_12967,N_12728,N_12711);
and U12968 (N_12968,N_12594,N_12744);
nand U12969 (N_12969,N_12716,N_12712);
nand U12970 (N_12970,N_12509,N_12726);
nor U12971 (N_12971,N_12603,N_12743);
nand U12972 (N_12972,N_12572,N_12586);
xor U12973 (N_12973,N_12606,N_12687);
xor U12974 (N_12974,N_12573,N_12558);
nor U12975 (N_12975,N_12678,N_12715);
and U12976 (N_12976,N_12519,N_12696);
xnor U12977 (N_12977,N_12622,N_12542);
and U12978 (N_12978,N_12505,N_12636);
xor U12979 (N_12979,N_12539,N_12698);
xor U12980 (N_12980,N_12588,N_12568);
xor U12981 (N_12981,N_12681,N_12667);
xnor U12982 (N_12982,N_12676,N_12700);
xnor U12983 (N_12983,N_12733,N_12605);
xnor U12984 (N_12984,N_12609,N_12698);
or U12985 (N_12985,N_12740,N_12683);
nor U12986 (N_12986,N_12679,N_12533);
xor U12987 (N_12987,N_12566,N_12534);
and U12988 (N_12988,N_12679,N_12726);
nor U12989 (N_12989,N_12518,N_12740);
nor U12990 (N_12990,N_12643,N_12688);
and U12991 (N_12991,N_12525,N_12737);
and U12992 (N_12992,N_12708,N_12601);
nor U12993 (N_12993,N_12512,N_12702);
and U12994 (N_12994,N_12513,N_12742);
and U12995 (N_12995,N_12689,N_12638);
nor U12996 (N_12996,N_12739,N_12673);
xor U12997 (N_12997,N_12569,N_12681);
nand U12998 (N_12998,N_12502,N_12696);
or U12999 (N_12999,N_12741,N_12624);
and U13000 (N_13000,N_12880,N_12818);
nor U13001 (N_13001,N_12866,N_12838);
or U13002 (N_13002,N_12924,N_12931);
xnor U13003 (N_13003,N_12884,N_12830);
and U13004 (N_13004,N_12815,N_12959);
nor U13005 (N_13005,N_12782,N_12810);
nor U13006 (N_13006,N_12992,N_12907);
or U13007 (N_13007,N_12820,N_12977);
or U13008 (N_13008,N_12895,N_12811);
xor U13009 (N_13009,N_12845,N_12856);
nor U13010 (N_13010,N_12971,N_12787);
nand U13011 (N_13011,N_12836,N_12763);
or U13012 (N_13012,N_12869,N_12934);
xor U13013 (N_13013,N_12808,N_12842);
nor U13014 (N_13014,N_12751,N_12939);
nand U13015 (N_13015,N_12802,N_12860);
or U13016 (N_13016,N_12864,N_12926);
nand U13017 (N_13017,N_12968,N_12991);
xor U13018 (N_13018,N_12755,N_12862);
and U13019 (N_13019,N_12908,N_12803);
or U13020 (N_13020,N_12916,N_12790);
nor U13021 (N_13021,N_12897,N_12874);
nand U13022 (N_13022,N_12919,N_12982);
nor U13023 (N_13023,N_12767,N_12921);
or U13024 (N_13024,N_12956,N_12758);
nand U13025 (N_13025,N_12909,N_12910);
or U13026 (N_13026,N_12801,N_12792);
and U13027 (N_13027,N_12998,N_12843);
and U13028 (N_13028,N_12891,N_12817);
and U13029 (N_13029,N_12796,N_12976);
nand U13030 (N_13030,N_12964,N_12783);
nand U13031 (N_13031,N_12881,N_12816);
and U13032 (N_13032,N_12943,N_12806);
nand U13033 (N_13033,N_12775,N_12993);
nor U13034 (N_13034,N_12784,N_12904);
or U13035 (N_13035,N_12954,N_12872);
and U13036 (N_13036,N_12854,N_12839);
nor U13037 (N_13037,N_12788,N_12994);
or U13038 (N_13038,N_12821,N_12987);
nor U13039 (N_13039,N_12957,N_12835);
or U13040 (N_13040,N_12868,N_12940);
nor U13041 (N_13041,N_12911,N_12963);
xor U13042 (N_13042,N_12780,N_12804);
xor U13043 (N_13043,N_12958,N_12932);
xnor U13044 (N_13044,N_12899,N_12847);
or U13045 (N_13045,N_12955,N_12915);
nand U13046 (N_13046,N_12850,N_12844);
or U13047 (N_13047,N_12773,N_12826);
nand U13048 (N_13048,N_12873,N_12795);
or U13049 (N_13049,N_12781,N_12990);
or U13050 (N_13050,N_12805,N_12876);
or U13051 (N_13051,N_12985,N_12950);
nor U13052 (N_13052,N_12962,N_12861);
nor U13053 (N_13053,N_12834,N_12886);
or U13054 (N_13054,N_12917,N_12807);
nor U13055 (N_13055,N_12814,N_12969);
or U13056 (N_13056,N_12945,N_12942);
xor U13057 (N_13057,N_12999,N_12941);
and U13058 (N_13058,N_12892,N_12898);
nor U13059 (N_13059,N_12809,N_12831);
nor U13060 (N_13060,N_12966,N_12827);
and U13061 (N_13061,N_12879,N_12825);
nor U13062 (N_13062,N_12865,N_12833);
and U13063 (N_13063,N_12829,N_12851);
xnor U13064 (N_13064,N_12855,N_12766);
nand U13065 (N_13065,N_12756,N_12961);
nor U13066 (N_13066,N_12846,N_12785);
or U13067 (N_13067,N_12912,N_12770);
nor U13068 (N_13068,N_12936,N_12761);
or U13069 (N_13069,N_12914,N_12885);
nand U13070 (N_13070,N_12970,N_12894);
and U13071 (N_13071,N_12857,N_12798);
xor U13072 (N_13072,N_12822,N_12965);
nor U13073 (N_13073,N_12887,N_12757);
or U13074 (N_13074,N_12824,N_12975);
or U13075 (N_13075,N_12774,N_12753);
xor U13076 (N_13076,N_12776,N_12989);
xor U13077 (N_13077,N_12901,N_12933);
or U13078 (N_13078,N_12896,N_12949);
nand U13079 (N_13079,N_12759,N_12800);
and U13080 (N_13080,N_12799,N_12980);
or U13081 (N_13081,N_12973,N_12867);
nand U13082 (N_13082,N_12967,N_12797);
xor U13083 (N_13083,N_12832,N_12922);
xor U13084 (N_13084,N_12750,N_12819);
xor U13085 (N_13085,N_12925,N_12972);
nand U13086 (N_13086,N_12841,N_12794);
nor U13087 (N_13087,N_12900,N_12764);
xor U13088 (N_13088,N_12870,N_12920);
and U13089 (N_13089,N_12983,N_12938);
nor U13090 (N_13090,N_12979,N_12840);
or U13091 (N_13091,N_12765,N_12984);
nand U13092 (N_13092,N_12863,N_12877);
and U13093 (N_13093,N_12890,N_12848);
xor U13094 (N_13094,N_12889,N_12883);
nor U13095 (N_13095,N_12929,N_12978);
and U13096 (N_13096,N_12859,N_12947);
or U13097 (N_13097,N_12918,N_12762);
and U13098 (N_13098,N_12760,N_12813);
or U13099 (N_13099,N_12944,N_12905);
nand U13100 (N_13100,N_12952,N_12754);
xor U13101 (N_13101,N_12997,N_12812);
or U13102 (N_13102,N_12913,N_12778);
xnor U13103 (N_13103,N_12779,N_12882);
and U13104 (N_13104,N_12902,N_12893);
and U13105 (N_13105,N_12995,N_12903);
nor U13106 (N_13106,N_12772,N_12777);
and U13107 (N_13107,N_12771,N_12752);
and U13108 (N_13108,N_12852,N_12974);
or U13109 (N_13109,N_12937,N_12981);
xor U13110 (N_13110,N_12789,N_12930);
nor U13111 (N_13111,N_12948,N_12986);
nor U13112 (N_13112,N_12996,N_12828);
nand U13113 (N_13113,N_12951,N_12791);
and U13114 (N_13114,N_12960,N_12871);
nor U13115 (N_13115,N_12793,N_12946);
or U13116 (N_13116,N_12888,N_12858);
xor U13117 (N_13117,N_12786,N_12837);
xor U13118 (N_13118,N_12823,N_12878);
or U13119 (N_13119,N_12849,N_12935);
nor U13120 (N_13120,N_12923,N_12953);
xor U13121 (N_13121,N_12768,N_12906);
or U13122 (N_13122,N_12853,N_12928);
nor U13123 (N_13123,N_12927,N_12988);
nand U13124 (N_13124,N_12769,N_12875);
nor U13125 (N_13125,N_12791,N_12971);
nor U13126 (N_13126,N_12861,N_12947);
xor U13127 (N_13127,N_12908,N_12893);
and U13128 (N_13128,N_12940,N_12820);
xnor U13129 (N_13129,N_12842,N_12995);
nor U13130 (N_13130,N_12882,N_12820);
or U13131 (N_13131,N_12784,N_12952);
or U13132 (N_13132,N_12839,N_12935);
nand U13133 (N_13133,N_12992,N_12983);
and U13134 (N_13134,N_12884,N_12788);
and U13135 (N_13135,N_12952,N_12913);
xor U13136 (N_13136,N_12921,N_12924);
and U13137 (N_13137,N_12757,N_12889);
nor U13138 (N_13138,N_12854,N_12752);
and U13139 (N_13139,N_12781,N_12891);
nand U13140 (N_13140,N_12818,N_12775);
nor U13141 (N_13141,N_12926,N_12896);
or U13142 (N_13142,N_12774,N_12842);
nand U13143 (N_13143,N_12956,N_12807);
nand U13144 (N_13144,N_12859,N_12835);
nand U13145 (N_13145,N_12772,N_12894);
nand U13146 (N_13146,N_12758,N_12944);
nor U13147 (N_13147,N_12834,N_12791);
or U13148 (N_13148,N_12876,N_12968);
xnor U13149 (N_13149,N_12842,N_12908);
or U13150 (N_13150,N_12865,N_12925);
xnor U13151 (N_13151,N_12817,N_12811);
or U13152 (N_13152,N_12766,N_12956);
nor U13153 (N_13153,N_12907,N_12764);
nor U13154 (N_13154,N_12988,N_12785);
or U13155 (N_13155,N_12884,N_12790);
or U13156 (N_13156,N_12978,N_12867);
nor U13157 (N_13157,N_12865,N_12973);
nand U13158 (N_13158,N_12821,N_12910);
or U13159 (N_13159,N_12870,N_12898);
and U13160 (N_13160,N_12859,N_12910);
nand U13161 (N_13161,N_12862,N_12945);
nor U13162 (N_13162,N_12811,N_12853);
nand U13163 (N_13163,N_12848,N_12974);
xnor U13164 (N_13164,N_12821,N_12900);
nand U13165 (N_13165,N_12943,N_12787);
nor U13166 (N_13166,N_12888,N_12841);
xor U13167 (N_13167,N_12829,N_12951);
nor U13168 (N_13168,N_12800,N_12835);
or U13169 (N_13169,N_12994,N_12757);
or U13170 (N_13170,N_12844,N_12949);
nand U13171 (N_13171,N_12838,N_12908);
nor U13172 (N_13172,N_12754,N_12872);
xnor U13173 (N_13173,N_12821,N_12983);
and U13174 (N_13174,N_12989,N_12865);
nand U13175 (N_13175,N_12845,N_12906);
xnor U13176 (N_13176,N_12926,N_12991);
xnor U13177 (N_13177,N_12991,N_12851);
xor U13178 (N_13178,N_12989,N_12977);
nor U13179 (N_13179,N_12857,N_12762);
or U13180 (N_13180,N_12783,N_12981);
xnor U13181 (N_13181,N_12870,N_12933);
xnor U13182 (N_13182,N_12787,N_12851);
and U13183 (N_13183,N_12835,N_12789);
and U13184 (N_13184,N_12992,N_12895);
and U13185 (N_13185,N_12828,N_12824);
nor U13186 (N_13186,N_12891,N_12830);
and U13187 (N_13187,N_12883,N_12922);
or U13188 (N_13188,N_12911,N_12943);
or U13189 (N_13189,N_12815,N_12862);
or U13190 (N_13190,N_12997,N_12962);
nand U13191 (N_13191,N_12893,N_12778);
nor U13192 (N_13192,N_12846,N_12967);
nor U13193 (N_13193,N_12937,N_12891);
and U13194 (N_13194,N_12780,N_12871);
nand U13195 (N_13195,N_12751,N_12973);
and U13196 (N_13196,N_12850,N_12959);
or U13197 (N_13197,N_12759,N_12919);
nor U13198 (N_13198,N_12963,N_12969);
xnor U13199 (N_13199,N_12958,N_12850);
xor U13200 (N_13200,N_12917,N_12971);
or U13201 (N_13201,N_12832,N_12991);
or U13202 (N_13202,N_12843,N_12862);
xnor U13203 (N_13203,N_12774,N_12888);
nand U13204 (N_13204,N_12845,N_12772);
and U13205 (N_13205,N_12812,N_12762);
or U13206 (N_13206,N_12843,N_12782);
and U13207 (N_13207,N_12877,N_12861);
or U13208 (N_13208,N_12961,N_12909);
nor U13209 (N_13209,N_12983,N_12968);
xor U13210 (N_13210,N_12915,N_12756);
nor U13211 (N_13211,N_12928,N_12774);
or U13212 (N_13212,N_12819,N_12832);
xnor U13213 (N_13213,N_12760,N_12762);
and U13214 (N_13214,N_12826,N_12769);
nand U13215 (N_13215,N_12812,N_12822);
or U13216 (N_13216,N_12758,N_12975);
nand U13217 (N_13217,N_12783,N_12863);
nor U13218 (N_13218,N_12988,N_12944);
nand U13219 (N_13219,N_12755,N_12770);
xor U13220 (N_13220,N_12873,N_12920);
and U13221 (N_13221,N_12905,N_12820);
and U13222 (N_13222,N_12832,N_12826);
nor U13223 (N_13223,N_12893,N_12981);
and U13224 (N_13224,N_12894,N_12863);
xor U13225 (N_13225,N_12902,N_12941);
xnor U13226 (N_13226,N_12849,N_12913);
xor U13227 (N_13227,N_12984,N_12909);
or U13228 (N_13228,N_12971,N_12766);
xor U13229 (N_13229,N_12817,N_12915);
or U13230 (N_13230,N_12841,N_12917);
nand U13231 (N_13231,N_12756,N_12840);
and U13232 (N_13232,N_12781,N_12890);
and U13233 (N_13233,N_12826,N_12950);
and U13234 (N_13234,N_12826,N_12983);
xnor U13235 (N_13235,N_12783,N_12880);
nand U13236 (N_13236,N_12980,N_12848);
nand U13237 (N_13237,N_12870,N_12769);
xor U13238 (N_13238,N_12791,N_12955);
nor U13239 (N_13239,N_12890,N_12873);
and U13240 (N_13240,N_12795,N_12973);
xnor U13241 (N_13241,N_12899,N_12895);
nor U13242 (N_13242,N_12876,N_12902);
xnor U13243 (N_13243,N_12782,N_12827);
or U13244 (N_13244,N_12933,N_12924);
nor U13245 (N_13245,N_12987,N_12993);
and U13246 (N_13246,N_12772,N_12910);
nor U13247 (N_13247,N_12842,N_12761);
and U13248 (N_13248,N_12905,N_12868);
and U13249 (N_13249,N_12885,N_12939);
xnor U13250 (N_13250,N_13174,N_13108);
nand U13251 (N_13251,N_13217,N_13194);
nand U13252 (N_13252,N_13042,N_13131);
nand U13253 (N_13253,N_13197,N_13113);
or U13254 (N_13254,N_13187,N_13009);
nor U13255 (N_13255,N_13040,N_13204);
and U13256 (N_13256,N_13230,N_13125);
and U13257 (N_13257,N_13126,N_13192);
xor U13258 (N_13258,N_13136,N_13201);
nand U13259 (N_13259,N_13248,N_13015);
or U13260 (N_13260,N_13013,N_13026);
and U13261 (N_13261,N_13016,N_13143);
xnor U13262 (N_13262,N_13072,N_13082);
xor U13263 (N_13263,N_13024,N_13055);
and U13264 (N_13264,N_13068,N_13019);
xnor U13265 (N_13265,N_13021,N_13229);
xor U13266 (N_13266,N_13234,N_13039);
xnor U13267 (N_13267,N_13169,N_13062);
or U13268 (N_13268,N_13132,N_13018);
nand U13269 (N_13269,N_13077,N_13209);
xnor U13270 (N_13270,N_13138,N_13227);
xor U13271 (N_13271,N_13189,N_13109);
nand U13272 (N_13272,N_13249,N_13215);
or U13273 (N_13273,N_13045,N_13036);
and U13274 (N_13274,N_13076,N_13180);
and U13275 (N_13275,N_13065,N_13218);
nor U13276 (N_13276,N_13089,N_13154);
and U13277 (N_13277,N_13128,N_13142);
and U13278 (N_13278,N_13231,N_13107);
nand U13279 (N_13279,N_13175,N_13239);
nor U13280 (N_13280,N_13228,N_13149);
xnor U13281 (N_13281,N_13240,N_13033);
and U13282 (N_13282,N_13099,N_13202);
xnor U13283 (N_13283,N_13027,N_13245);
or U13284 (N_13284,N_13014,N_13117);
nor U13285 (N_13285,N_13145,N_13114);
xnor U13286 (N_13286,N_13166,N_13066);
xnor U13287 (N_13287,N_13195,N_13071);
or U13288 (N_13288,N_13199,N_13102);
nor U13289 (N_13289,N_13012,N_13105);
nor U13290 (N_13290,N_13122,N_13073);
nand U13291 (N_13291,N_13165,N_13130);
or U13292 (N_13292,N_13177,N_13101);
nor U13293 (N_13293,N_13184,N_13002);
or U13294 (N_13294,N_13241,N_13060);
nand U13295 (N_13295,N_13119,N_13236);
nor U13296 (N_13296,N_13111,N_13148);
and U13297 (N_13297,N_13163,N_13146);
and U13298 (N_13298,N_13008,N_13235);
xor U13299 (N_13299,N_13124,N_13020);
xor U13300 (N_13300,N_13196,N_13216);
or U13301 (N_13301,N_13049,N_13147);
nor U13302 (N_13302,N_13158,N_13244);
xor U13303 (N_13303,N_13162,N_13023);
or U13304 (N_13304,N_13246,N_13211);
xnor U13305 (N_13305,N_13198,N_13170);
or U13306 (N_13306,N_13046,N_13185);
or U13307 (N_13307,N_13096,N_13004);
nor U13308 (N_13308,N_13050,N_13086);
nand U13309 (N_13309,N_13176,N_13193);
nor U13310 (N_13310,N_13074,N_13092);
and U13311 (N_13311,N_13220,N_13210);
or U13312 (N_13312,N_13080,N_13100);
or U13313 (N_13313,N_13135,N_13129);
xor U13314 (N_13314,N_13094,N_13063);
and U13315 (N_13315,N_13078,N_13153);
and U13316 (N_13316,N_13173,N_13075);
or U13317 (N_13317,N_13051,N_13161);
and U13318 (N_13318,N_13150,N_13043);
nand U13319 (N_13319,N_13121,N_13186);
and U13320 (N_13320,N_13041,N_13237);
nor U13321 (N_13321,N_13106,N_13031);
nor U13322 (N_13322,N_13067,N_13118);
or U13323 (N_13323,N_13144,N_13238);
xnor U13324 (N_13324,N_13053,N_13047);
and U13325 (N_13325,N_13167,N_13133);
nand U13326 (N_13326,N_13214,N_13242);
nand U13327 (N_13327,N_13152,N_13090);
nand U13328 (N_13328,N_13134,N_13178);
xnor U13329 (N_13329,N_13035,N_13059);
nand U13330 (N_13330,N_13182,N_13213);
and U13331 (N_13331,N_13123,N_13205);
nand U13332 (N_13332,N_13001,N_13110);
nand U13333 (N_13333,N_13091,N_13159);
xnor U13334 (N_13334,N_13093,N_13222);
nand U13335 (N_13335,N_13200,N_13140);
and U13336 (N_13336,N_13168,N_13037);
nand U13337 (N_13337,N_13069,N_13172);
or U13338 (N_13338,N_13017,N_13005);
xor U13339 (N_13339,N_13225,N_13137);
nand U13340 (N_13340,N_13083,N_13155);
xnor U13341 (N_13341,N_13183,N_13156);
nand U13342 (N_13342,N_13103,N_13219);
and U13343 (N_13343,N_13000,N_13056);
and U13344 (N_13344,N_13007,N_13104);
and U13345 (N_13345,N_13233,N_13098);
nor U13346 (N_13346,N_13188,N_13029);
nand U13347 (N_13347,N_13243,N_13203);
xor U13348 (N_13348,N_13088,N_13157);
nand U13349 (N_13349,N_13116,N_13171);
nor U13350 (N_13350,N_13207,N_13006);
nand U13351 (N_13351,N_13087,N_13224);
nand U13352 (N_13352,N_13160,N_13044);
nand U13353 (N_13353,N_13191,N_13003);
or U13354 (N_13354,N_13151,N_13212);
and U13355 (N_13355,N_13048,N_13070);
or U13356 (N_13356,N_13221,N_13064);
nand U13357 (N_13357,N_13223,N_13232);
or U13358 (N_13358,N_13085,N_13097);
nor U13359 (N_13359,N_13247,N_13226);
nand U13360 (N_13360,N_13127,N_13057);
xor U13361 (N_13361,N_13022,N_13115);
and U13362 (N_13362,N_13139,N_13079);
xor U13363 (N_13363,N_13120,N_13034);
nor U13364 (N_13364,N_13179,N_13030);
or U13365 (N_13365,N_13181,N_13081);
nand U13366 (N_13366,N_13010,N_13032);
nor U13367 (N_13367,N_13025,N_13084);
xor U13368 (N_13368,N_13206,N_13054);
nor U13369 (N_13369,N_13028,N_13190);
nand U13370 (N_13370,N_13038,N_13052);
or U13371 (N_13371,N_13141,N_13061);
xnor U13372 (N_13372,N_13095,N_13208);
or U13373 (N_13373,N_13112,N_13011);
and U13374 (N_13374,N_13164,N_13058);
nor U13375 (N_13375,N_13167,N_13044);
nor U13376 (N_13376,N_13039,N_13035);
and U13377 (N_13377,N_13017,N_13126);
nand U13378 (N_13378,N_13249,N_13143);
xor U13379 (N_13379,N_13091,N_13161);
and U13380 (N_13380,N_13086,N_13071);
and U13381 (N_13381,N_13032,N_13168);
and U13382 (N_13382,N_13069,N_13039);
or U13383 (N_13383,N_13179,N_13245);
nor U13384 (N_13384,N_13174,N_13241);
xnor U13385 (N_13385,N_13110,N_13012);
xnor U13386 (N_13386,N_13025,N_13217);
nor U13387 (N_13387,N_13146,N_13166);
xor U13388 (N_13388,N_13012,N_13005);
xor U13389 (N_13389,N_13046,N_13029);
nor U13390 (N_13390,N_13107,N_13105);
nor U13391 (N_13391,N_13142,N_13147);
xnor U13392 (N_13392,N_13099,N_13019);
nand U13393 (N_13393,N_13192,N_13018);
nor U13394 (N_13394,N_13178,N_13019);
xnor U13395 (N_13395,N_13119,N_13114);
nand U13396 (N_13396,N_13060,N_13171);
nor U13397 (N_13397,N_13198,N_13233);
nor U13398 (N_13398,N_13199,N_13200);
nand U13399 (N_13399,N_13150,N_13086);
xnor U13400 (N_13400,N_13135,N_13236);
and U13401 (N_13401,N_13019,N_13006);
nand U13402 (N_13402,N_13016,N_13183);
nor U13403 (N_13403,N_13140,N_13043);
nand U13404 (N_13404,N_13129,N_13131);
or U13405 (N_13405,N_13022,N_13189);
nand U13406 (N_13406,N_13107,N_13039);
and U13407 (N_13407,N_13240,N_13050);
nand U13408 (N_13408,N_13181,N_13060);
xor U13409 (N_13409,N_13217,N_13162);
and U13410 (N_13410,N_13142,N_13032);
nand U13411 (N_13411,N_13155,N_13026);
nor U13412 (N_13412,N_13049,N_13199);
nor U13413 (N_13413,N_13017,N_13217);
or U13414 (N_13414,N_13005,N_13022);
or U13415 (N_13415,N_13168,N_13019);
nand U13416 (N_13416,N_13073,N_13028);
and U13417 (N_13417,N_13182,N_13187);
nor U13418 (N_13418,N_13127,N_13134);
nor U13419 (N_13419,N_13210,N_13106);
xor U13420 (N_13420,N_13078,N_13209);
nor U13421 (N_13421,N_13228,N_13205);
xnor U13422 (N_13422,N_13116,N_13216);
nor U13423 (N_13423,N_13083,N_13116);
and U13424 (N_13424,N_13116,N_13010);
nand U13425 (N_13425,N_13064,N_13033);
nor U13426 (N_13426,N_13023,N_13157);
xor U13427 (N_13427,N_13036,N_13221);
or U13428 (N_13428,N_13162,N_13239);
xnor U13429 (N_13429,N_13244,N_13003);
or U13430 (N_13430,N_13082,N_13118);
nor U13431 (N_13431,N_13122,N_13128);
nand U13432 (N_13432,N_13121,N_13063);
and U13433 (N_13433,N_13012,N_13176);
or U13434 (N_13434,N_13051,N_13143);
and U13435 (N_13435,N_13128,N_13118);
xnor U13436 (N_13436,N_13035,N_13131);
nand U13437 (N_13437,N_13032,N_13161);
and U13438 (N_13438,N_13178,N_13080);
and U13439 (N_13439,N_13051,N_13159);
or U13440 (N_13440,N_13209,N_13105);
xnor U13441 (N_13441,N_13054,N_13015);
or U13442 (N_13442,N_13115,N_13178);
xnor U13443 (N_13443,N_13012,N_13232);
and U13444 (N_13444,N_13081,N_13043);
xnor U13445 (N_13445,N_13034,N_13042);
and U13446 (N_13446,N_13226,N_13075);
nand U13447 (N_13447,N_13047,N_13175);
xnor U13448 (N_13448,N_13117,N_13247);
nand U13449 (N_13449,N_13100,N_13178);
or U13450 (N_13450,N_13247,N_13209);
and U13451 (N_13451,N_13027,N_13219);
or U13452 (N_13452,N_13141,N_13081);
or U13453 (N_13453,N_13010,N_13197);
and U13454 (N_13454,N_13014,N_13063);
xor U13455 (N_13455,N_13159,N_13025);
xnor U13456 (N_13456,N_13109,N_13152);
nand U13457 (N_13457,N_13222,N_13248);
nor U13458 (N_13458,N_13126,N_13224);
nand U13459 (N_13459,N_13073,N_13230);
or U13460 (N_13460,N_13185,N_13129);
or U13461 (N_13461,N_13248,N_13035);
xnor U13462 (N_13462,N_13204,N_13064);
nand U13463 (N_13463,N_13144,N_13167);
and U13464 (N_13464,N_13172,N_13035);
xor U13465 (N_13465,N_13184,N_13007);
xor U13466 (N_13466,N_13051,N_13201);
xnor U13467 (N_13467,N_13020,N_13138);
xnor U13468 (N_13468,N_13078,N_13243);
nand U13469 (N_13469,N_13125,N_13184);
nand U13470 (N_13470,N_13141,N_13019);
and U13471 (N_13471,N_13169,N_13159);
nor U13472 (N_13472,N_13209,N_13180);
nor U13473 (N_13473,N_13104,N_13123);
and U13474 (N_13474,N_13034,N_13040);
xnor U13475 (N_13475,N_13125,N_13191);
nor U13476 (N_13476,N_13177,N_13039);
or U13477 (N_13477,N_13159,N_13037);
nor U13478 (N_13478,N_13191,N_13226);
xor U13479 (N_13479,N_13018,N_13106);
or U13480 (N_13480,N_13016,N_13063);
nor U13481 (N_13481,N_13142,N_13208);
nand U13482 (N_13482,N_13119,N_13089);
nor U13483 (N_13483,N_13054,N_13119);
and U13484 (N_13484,N_13059,N_13167);
nor U13485 (N_13485,N_13082,N_13237);
or U13486 (N_13486,N_13165,N_13170);
nor U13487 (N_13487,N_13033,N_13124);
xnor U13488 (N_13488,N_13043,N_13240);
nand U13489 (N_13489,N_13219,N_13045);
xor U13490 (N_13490,N_13234,N_13048);
xor U13491 (N_13491,N_13142,N_13233);
nand U13492 (N_13492,N_13190,N_13229);
or U13493 (N_13493,N_13236,N_13155);
nor U13494 (N_13494,N_13143,N_13141);
xor U13495 (N_13495,N_13046,N_13242);
or U13496 (N_13496,N_13219,N_13206);
or U13497 (N_13497,N_13026,N_13060);
or U13498 (N_13498,N_13206,N_13202);
or U13499 (N_13499,N_13088,N_13104);
or U13500 (N_13500,N_13284,N_13404);
nand U13501 (N_13501,N_13487,N_13292);
or U13502 (N_13502,N_13288,N_13299);
and U13503 (N_13503,N_13477,N_13462);
nand U13504 (N_13504,N_13301,N_13260);
and U13505 (N_13505,N_13371,N_13403);
xor U13506 (N_13506,N_13412,N_13359);
or U13507 (N_13507,N_13428,N_13431);
nor U13508 (N_13508,N_13256,N_13420);
xor U13509 (N_13509,N_13258,N_13336);
nor U13510 (N_13510,N_13330,N_13360);
nor U13511 (N_13511,N_13480,N_13463);
and U13512 (N_13512,N_13343,N_13375);
xnor U13513 (N_13513,N_13255,N_13282);
or U13514 (N_13514,N_13277,N_13281);
or U13515 (N_13515,N_13278,N_13347);
and U13516 (N_13516,N_13468,N_13352);
xnor U13517 (N_13517,N_13400,N_13493);
and U13518 (N_13518,N_13327,N_13322);
or U13519 (N_13519,N_13443,N_13422);
nand U13520 (N_13520,N_13460,N_13426);
and U13521 (N_13521,N_13419,N_13435);
and U13522 (N_13522,N_13449,N_13250);
nand U13523 (N_13523,N_13318,N_13483);
or U13524 (N_13524,N_13499,N_13251);
nor U13525 (N_13525,N_13309,N_13459);
or U13526 (N_13526,N_13399,N_13302);
xor U13527 (N_13527,N_13490,N_13466);
xor U13528 (N_13528,N_13437,N_13384);
xor U13529 (N_13529,N_13446,N_13316);
and U13530 (N_13530,N_13315,N_13286);
and U13531 (N_13531,N_13252,N_13409);
nand U13532 (N_13532,N_13464,N_13311);
and U13533 (N_13533,N_13436,N_13323);
nor U13534 (N_13534,N_13484,N_13355);
and U13535 (N_13535,N_13314,N_13313);
nand U13536 (N_13536,N_13306,N_13398);
or U13537 (N_13537,N_13329,N_13310);
or U13538 (N_13538,N_13442,N_13401);
nor U13539 (N_13539,N_13396,N_13351);
or U13540 (N_13540,N_13290,N_13394);
nor U13541 (N_13541,N_13391,N_13357);
nand U13542 (N_13542,N_13332,N_13272);
nand U13543 (N_13543,N_13317,N_13274);
nand U13544 (N_13544,N_13273,N_13312);
and U13545 (N_13545,N_13358,N_13334);
nor U13546 (N_13546,N_13319,N_13366);
nor U13547 (N_13547,N_13455,N_13451);
nor U13548 (N_13548,N_13485,N_13433);
xor U13549 (N_13549,N_13370,N_13305);
nor U13550 (N_13550,N_13498,N_13430);
and U13551 (N_13551,N_13265,N_13264);
nand U13552 (N_13552,N_13349,N_13254);
or U13553 (N_13553,N_13440,N_13388);
nand U13554 (N_13554,N_13425,N_13478);
or U13555 (N_13555,N_13479,N_13297);
xnor U13556 (N_13556,N_13296,N_13368);
nor U13557 (N_13557,N_13465,N_13450);
or U13558 (N_13558,N_13467,N_13365);
or U13559 (N_13559,N_13331,N_13476);
nand U13560 (N_13560,N_13362,N_13488);
nand U13561 (N_13561,N_13275,N_13339);
and U13562 (N_13562,N_13387,N_13304);
nand U13563 (N_13563,N_13432,N_13452);
xor U13564 (N_13564,N_13494,N_13389);
xnor U13565 (N_13565,N_13390,N_13453);
or U13566 (N_13566,N_13475,N_13376);
and U13567 (N_13567,N_13456,N_13356);
nand U13568 (N_13568,N_13324,N_13289);
xnor U13569 (N_13569,N_13427,N_13361);
nand U13570 (N_13570,N_13374,N_13364);
nand U13571 (N_13571,N_13378,N_13385);
nor U13572 (N_13572,N_13441,N_13344);
nand U13573 (N_13573,N_13495,N_13380);
and U13574 (N_13574,N_13262,N_13406);
or U13575 (N_13575,N_13345,N_13280);
nor U13576 (N_13576,N_13393,N_13413);
nand U13577 (N_13577,N_13285,N_13335);
and U13578 (N_13578,N_13342,N_13461);
nor U13579 (N_13579,N_13328,N_13397);
or U13580 (N_13580,N_13259,N_13271);
and U13581 (N_13581,N_13307,N_13372);
and U13582 (N_13582,N_13300,N_13482);
or U13583 (N_13583,N_13382,N_13270);
nor U13584 (N_13584,N_13408,N_13353);
and U13585 (N_13585,N_13407,N_13333);
nand U13586 (N_13586,N_13350,N_13373);
xor U13587 (N_13587,N_13415,N_13308);
or U13588 (N_13588,N_13445,N_13392);
and U13589 (N_13589,N_13411,N_13421);
nor U13590 (N_13590,N_13253,N_13269);
xor U13591 (N_13591,N_13377,N_13473);
nand U13592 (N_13592,N_13448,N_13447);
nor U13593 (N_13593,N_13418,N_13386);
nor U13594 (N_13594,N_13291,N_13303);
and U13595 (N_13595,N_13439,N_13348);
xor U13596 (N_13596,N_13423,N_13325);
or U13597 (N_13597,N_13492,N_13268);
xor U13598 (N_13598,N_13321,N_13454);
nand U13599 (N_13599,N_13486,N_13474);
nand U13600 (N_13600,N_13497,N_13276);
nor U13601 (N_13601,N_13295,N_13341);
and U13602 (N_13602,N_13402,N_13491);
nand U13603 (N_13603,N_13424,N_13266);
nand U13604 (N_13604,N_13340,N_13414);
and U13605 (N_13605,N_13444,N_13410);
nor U13606 (N_13606,N_13472,N_13294);
and U13607 (N_13607,N_13326,N_13458);
nand U13608 (N_13608,N_13369,N_13416);
or U13609 (N_13609,N_13257,N_13470);
nand U13610 (N_13610,N_13383,N_13429);
nor U13611 (N_13611,N_13279,N_13263);
nor U13612 (N_13612,N_13346,N_13489);
or U13613 (N_13613,N_13367,N_13267);
and U13614 (N_13614,N_13261,N_13338);
nor U13615 (N_13615,N_13379,N_13438);
and U13616 (N_13616,N_13354,N_13457);
and U13617 (N_13617,N_13481,N_13405);
and U13618 (N_13618,N_13287,N_13298);
and U13619 (N_13619,N_13320,N_13496);
and U13620 (N_13620,N_13283,N_13471);
nor U13621 (N_13621,N_13417,N_13395);
or U13622 (N_13622,N_13469,N_13363);
or U13623 (N_13623,N_13293,N_13434);
xnor U13624 (N_13624,N_13337,N_13381);
xnor U13625 (N_13625,N_13408,N_13299);
nor U13626 (N_13626,N_13426,N_13497);
nand U13627 (N_13627,N_13472,N_13486);
nor U13628 (N_13628,N_13359,N_13279);
or U13629 (N_13629,N_13317,N_13294);
nand U13630 (N_13630,N_13476,N_13335);
and U13631 (N_13631,N_13365,N_13435);
nor U13632 (N_13632,N_13334,N_13318);
nor U13633 (N_13633,N_13372,N_13495);
nor U13634 (N_13634,N_13476,N_13330);
nor U13635 (N_13635,N_13358,N_13377);
xor U13636 (N_13636,N_13415,N_13391);
nor U13637 (N_13637,N_13394,N_13364);
or U13638 (N_13638,N_13353,N_13377);
and U13639 (N_13639,N_13317,N_13431);
xnor U13640 (N_13640,N_13417,N_13483);
and U13641 (N_13641,N_13405,N_13331);
or U13642 (N_13642,N_13293,N_13273);
nand U13643 (N_13643,N_13494,N_13295);
and U13644 (N_13644,N_13379,N_13308);
xor U13645 (N_13645,N_13408,N_13295);
nor U13646 (N_13646,N_13427,N_13481);
nand U13647 (N_13647,N_13334,N_13290);
xnor U13648 (N_13648,N_13263,N_13457);
or U13649 (N_13649,N_13447,N_13259);
or U13650 (N_13650,N_13403,N_13359);
nor U13651 (N_13651,N_13473,N_13346);
xnor U13652 (N_13652,N_13309,N_13327);
or U13653 (N_13653,N_13354,N_13475);
and U13654 (N_13654,N_13492,N_13274);
nor U13655 (N_13655,N_13368,N_13461);
xnor U13656 (N_13656,N_13346,N_13480);
nor U13657 (N_13657,N_13490,N_13440);
nand U13658 (N_13658,N_13309,N_13388);
nand U13659 (N_13659,N_13255,N_13362);
or U13660 (N_13660,N_13422,N_13478);
nand U13661 (N_13661,N_13348,N_13370);
or U13662 (N_13662,N_13379,N_13448);
and U13663 (N_13663,N_13439,N_13448);
nand U13664 (N_13664,N_13256,N_13252);
xor U13665 (N_13665,N_13289,N_13490);
xor U13666 (N_13666,N_13461,N_13275);
and U13667 (N_13667,N_13381,N_13302);
nand U13668 (N_13668,N_13348,N_13426);
nand U13669 (N_13669,N_13294,N_13460);
xor U13670 (N_13670,N_13364,N_13393);
xor U13671 (N_13671,N_13446,N_13250);
xor U13672 (N_13672,N_13431,N_13360);
xor U13673 (N_13673,N_13453,N_13338);
nand U13674 (N_13674,N_13315,N_13271);
xnor U13675 (N_13675,N_13374,N_13401);
and U13676 (N_13676,N_13393,N_13300);
or U13677 (N_13677,N_13442,N_13355);
nor U13678 (N_13678,N_13352,N_13255);
or U13679 (N_13679,N_13288,N_13471);
and U13680 (N_13680,N_13446,N_13430);
and U13681 (N_13681,N_13341,N_13371);
and U13682 (N_13682,N_13357,N_13457);
nand U13683 (N_13683,N_13328,N_13287);
or U13684 (N_13684,N_13337,N_13365);
nand U13685 (N_13685,N_13479,N_13426);
nor U13686 (N_13686,N_13412,N_13283);
nor U13687 (N_13687,N_13480,N_13386);
xnor U13688 (N_13688,N_13356,N_13281);
xor U13689 (N_13689,N_13311,N_13322);
xnor U13690 (N_13690,N_13451,N_13476);
nor U13691 (N_13691,N_13282,N_13489);
or U13692 (N_13692,N_13343,N_13424);
or U13693 (N_13693,N_13257,N_13342);
and U13694 (N_13694,N_13384,N_13450);
and U13695 (N_13695,N_13251,N_13386);
nor U13696 (N_13696,N_13397,N_13429);
nand U13697 (N_13697,N_13447,N_13306);
nand U13698 (N_13698,N_13487,N_13498);
or U13699 (N_13699,N_13357,N_13272);
nor U13700 (N_13700,N_13402,N_13438);
or U13701 (N_13701,N_13292,N_13474);
or U13702 (N_13702,N_13317,N_13445);
nor U13703 (N_13703,N_13253,N_13487);
nand U13704 (N_13704,N_13305,N_13253);
xor U13705 (N_13705,N_13438,N_13399);
or U13706 (N_13706,N_13437,N_13275);
xor U13707 (N_13707,N_13353,N_13280);
xor U13708 (N_13708,N_13491,N_13326);
or U13709 (N_13709,N_13284,N_13377);
and U13710 (N_13710,N_13378,N_13418);
xnor U13711 (N_13711,N_13384,N_13419);
and U13712 (N_13712,N_13451,N_13292);
or U13713 (N_13713,N_13307,N_13314);
and U13714 (N_13714,N_13429,N_13279);
nand U13715 (N_13715,N_13376,N_13377);
and U13716 (N_13716,N_13410,N_13294);
nor U13717 (N_13717,N_13345,N_13407);
or U13718 (N_13718,N_13285,N_13261);
or U13719 (N_13719,N_13303,N_13438);
or U13720 (N_13720,N_13475,N_13463);
nor U13721 (N_13721,N_13463,N_13434);
xor U13722 (N_13722,N_13432,N_13271);
nand U13723 (N_13723,N_13405,N_13369);
xor U13724 (N_13724,N_13454,N_13405);
nand U13725 (N_13725,N_13417,N_13376);
xor U13726 (N_13726,N_13315,N_13391);
nor U13727 (N_13727,N_13324,N_13385);
or U13728 (N_13728,N_13354,N_13343);
and U13729 (N_13729,N_13422,N_13474);
nor U13730 (N_13730,N_13401,N_13356);
xnor U13731 (N_13731,N_13429,N_13280);
nor U13732 (N_13732,N_13399,N_13295);
and U13733 (N_13733,N_13293,N_13320);
nor U13734 (N_13734,N_13269,N_13382);
or U13735 (N_13735,N_13363,N_13481);
or U13736 (N_13736,N_13467,N_13419);
or U13737 (N_13737,N_13319,N_13490);
and U13738 (N_13738,N_13385,N_13313);
and U13739 (N_13739,N_13268,N_13451);
and U13740 (N_13740,N_13340,N_13434);
xnor U13741 (N_13741,N_13289,N_13475);
xnor U13742 (N_13742,N_13451,N_13428);
nand U13743 (N_13743,N_13305,N_13333);
nand U13744 (N_13744,N_13495,N_13423);
nor U13745 (N_13745,N_13264,N_13313);
or U13746 (N_13746,N_13351,N_13266);
or U13747 (N_13747,N_13393,N_13319);
and U13748 (N_13748,N_13444,N_13293);
xor U13749 (N_13749,N_13333,N_13459);
xor U13750 (N_13750,N_13552,N_13646);
xnor U13751 (N_13751,N_13650,N_13538);
and U13752 (N_13752,N_13508,N_13642);
or U13753 (N_13753,N_13676,N_13608);
nor U13754 (N_13754,N_13560,N_13717);
nor U13755 (N_13755,N_13696,N_13692);
or U13756 (N_13756,N_13701,N_13574);
nand U13757 (N_13757,N_13592,N_13689);
nor U13758 (N_13758,N_13669,N_13513);
and U13759 (N_13759,N_13655,N_13584);
and U13760 (N_13760,N_13688,N_13607);
and U13761 (N_13761,N_13520,N_13534);
and U13762 (N_13762,N_13525,N_13599);
nor U13763 (N_13763,N_13517,N_13622);
nor U13764 (N_13764,N_13714,N_13531);
and U13765 (N_13765,N_13743,N_13734);
and U13766 (N_13766,N_13524,N_13647);
nor U13767 (N_13767,N_13710,N_13548);
and U13768 (N_13768,N_13736,N_13621);
or U13769 (N_13769,N_13747,N_13549);
or U13770 (N_13770,N_13526,N_13562);
and U13771 (N_13771,N_13609,N_13698);
nand U13772 (N_13772,N_13519,N_13542);
nand U13773 (N_13773,N_13545,N_13648);
nor U13774 (N_13774,N_13706,N_13658);
nand U13775 (N_13775,N_13652,N_13606);
nor U13776 (N_13776,N_13656,N_13615);
nor U13777 (N_13777,N_13687,N_13539);
or U13778 (N_13778,N_13677,N_13675);
nand U13779 (N_13779,N_13521,N_13708);
nand U13780 (N_13780,N_13505,N_13593);
nor U13781 (N_13781,N_13641,N_13620);
or U13782 (N_13782,N_13566,N_13724);
nor U13783 (N_13783,N_13651,N_13554);
nand U13784 (N_13784,N_13674,N_13564);
nor U13785 (N_13785,N_13719,N_13604);
nand U13786 (N_13786,N_13600,N_13516);
or U13787 (N_13787,N_13636,N_13660);
nor U13788 (N_13788,N_13661,N_13618);
nand U13789 (N_13789,N_13718,N_13720);
xor U13790 (N_13790,N_13594,N_13684);
nand U13791 (N_13791,N_13670,N_13640);
nand U13792 (N_13792,N_13553,N_13630);
nor U13793 (N_13793,N_13536,N_13707);
nand U13794 (N_13794,N_13523,N_13738);
xor U13795 (N_13795,N_13711,N_13702);
xor U13796 (N_13796,N_13737,N_13697);
nor U13797 (N_13797,N_13629,N_13537);
nor U13798 (N_13798,N_13581,N_13597);
nand U13799 (N_13799,N_13511,N_13590);
or U13800 (N_13800,N_13579,N_13583);
nor U13801 (N_13801,N_13506,N_13569);
and U13802 (N_13802,N_13632,N_13682);
and U13803 (N_13803,N_13730,N_13735);
nand U13804 (N_13804,N_13644,N_13625);
and U13805 (N_13805,N_13741,N_13654);
or U13806 (N_13806,N_13703,N_13673);
xnor U13807 (N_13807,N_13598,N_13572);
nand U13808 (N_13808,N_13712,N_13504);
xor U13809 (N_13809,N_13726,N_13685);
nand U13810 (N_13810,N_13613,N_13510);
nand U13811 (N_13811,N_13605,N_13589);
nor U13812 (N_13812,N_13699,N_13602);
nand U13813 (N_13813,N_13666,N_13623);
and U13814 (N_13814,N_13663,N_13507);
xnor U13815 (N_13815,N_13722,N_13515);
and U13816 (N_13816,N_13619,N_13561);
nor U13817 (N_13817,N_13700,N_13540);
nand U13818 (N_13818,N_13558,N_13500);
nand U13819 (N_13819,N_13533,N_13631);
nand U13820 (N_13820,N_13638,N_13744);
nand U13821 (N_13821,N_13679,N_13628);
xor U13822 (N_13822,N_13749,N_13532);
xor U13823 (N_13823,N_13691,N_13501);
nand U13824 (N_13824,N_13727,N_13530);
nor U13825 (N_13825,N_13657,N_13614);
nand U13826 (N_13826,N_13695,N_13627);
nand U13827 (N_13827,N_13535,N_13585);
or U13828 (N_13828,N_13728,N_13528);
xor U13829 (N_13829,N_13557,N_13509);
or U13830 (N_13830,N_13616,N_13514);
and U13831 (N_13831,N_13704,N_13643);
nand U13832 (N_13832,N_13740,N_13716);
and U13833 (N_13833,N_13576,N_13543);
and U13834 (N_13834,N_13522,N_13649);
and U13835 (N_13835,N_13551,N_13550);
nor U13836 (N_13836,N_13575,N_13731);
xor U13837 (N_13837,N_13596,N_13659);
or U13838 (N_13838,N_13635,N_13665);
and U13839 (N_13839,N_13544,N_13681);
nand U13840 (N_13840,N_13748,N_13586);
nor U13841 (N_13841,N_13577,N_13746);
nor U13842 (N_13842,N_13555,N_13678);
and U13843 (N_13843,N_13527,N_13693);
and U13844 (N_13844,N_13603,N_13683);
nor U13845 (N_13845,N_13729,N_13742);
nand U13846 (N_13846,N_13588,N_13694);
xnor U13847 (N_13847,N_13671,N_13745);
and U13848 (N_13848,N_13582,N_13723);
xor U13849 (N_13849,N_13591,N_13612);
nor U13850 (N_13850,N_13617,N_13637);
and U13851 (N_13851,N_13667,N_13578);
and U13852 (N_13852,N_13653,N_13705);
xnor U13853 (N_13853,N_13611,N_13664);
nand U13854 (N_13854,N_13709,N_13668);
and U13855 (N_13855,N_13512,N_13645);
xor U13856 (N_13856,N_13601,N_13721);
nor U13857 (N_13857,N_13732,N_13518);
nand U13858 (N_13858,N_13541,N_13686);
or U13859 (N_13859,N_13547,N_13680);
and U13860 (N_13860,N_13595,N_13610);
nand U13861 (N_13861,N_13624,N_13587);
or U13862 (N_13862,N_13556,N_13502);
and U13863 (N_13863,N_13563,N_13739);
and U13864 (N_13864,N_13672,N_13733);
nor U13865 (N_13865,N_13529,N_13570);
and U13866 (N_13866,N_13559,N_13662);
nor U13867 (N_13867,N_13565,N_13713);
xnor U13868 (N_13868,N_13567,N_13573);
nor U13869 (N_13869,N_13639,N_13690);
nor U13870 (N_13870,N_13546,N_13715);
or U13871 (N_13871,N_13580,N_13634);
nor U13872 (N_13872,N_13503,N_13633);
nor U13873 (N_13873,N_13626,N_13571);
nor U13874 (N_13874,N_13568,N_13725);
nor U13875 (N_13875,N_13599,N_13522);
nor U13876 (N_13876,N_13576,N_13734);
and U13877 (N_13877,N_13677,N_13673);
nand U13878 (N_13878,N_13599,N_13717);
and U13879 (N_13879,N_13571,N_13733);
nand U13880 (N_13880,N_13615,N_13736);
nand U13881 (N_13881,N_13717,N_13671);
xor U13882 (N_13882,N_13671,N_13560);
nand U13883 (N_13883,N_13515,N_13571);
and U13884 (N_13884,N_13735,N_13737);
nand U13885 (N_13885,N_13613,N_13624);
and U13886 (N_13886,N_13722,N_13683);
and U13887 (N_13887,N_13702,N_13544);
xnor U13888 (N_13888,N_13641,N_13747);
nand U13889 (N_13889,N_13685,N_13707);
and U13890 (N_13890,N_13521,N_13589);
or U13891 (N_13891,N_13550,N_13665);
or U13892 (N_13892,N_13720,N_13651);
and U13893 (N_13893,N_13666,N_13637);
xor U13894 (N_13894,N_13642,N_13514);
and U13895 (N_13895,N_13648,N_13623);
and U13896 (N_13896,N_13568,N_13682);
xor U13897 (N_13897,N_13703,N_13674);
nor U13898 (N_13898,N_13727,N_13673);
nand U13899 (N_13899,N_13722,N_13583);
xor U13900 (N_13900,N_13634,N_13706);
or U13901 (N_13901,N_13740,N_13726);
and U13902 (N_13902,N_13587,N_13647);
nand U13903 (N_13903,N_13668,N_13502);
and U13904 (N_13904,N_13629,N_13743);
xor U13905 (N_13905,N_13598,N_13715);
xnor U13906 (N_13906,N_13650,N_13508);
nand U13907 (N_13907,N_13671,N_13652);
nor U13908 (N_13908,N_13518,N_13602);
nand U13909 (N_13909,N_13615,N_13599);
xnor U13910 (N_13910,N_13578,N_13574);
nand U13911 (N_13911,N_13672,N_13552);
and U13912 (N_13912,N_13662,N_13697);
xor U13913 (N_13913,N_13529,N_13678);
and U13914 (N_13914,N_13632,N_13511);
nand U13915 (N_13915,N_13513,N_13530);
and U13916 (N_13916,N_13636,N_13746);
or U13917 (N_13917,N_13579,N_13694);
nand U13918 (N_13918,N_13628,N_13630);
nand U13919 (N_13919,N_13530,N_13614);
xnor U13920 (N_13920,N_13749,N_13710);
or U13921 (N_13921,N_13740,N_13615);
xor U13922 (N_13922,N_13540,N_13562);
or U13923 (N_13923,N_13668,N_13659);
or U13924 (N_13924,N_13655,N_13598);
nor U13925 (N_13925,N_13730,N_13573);
and U13926 (N_13926,N_13527,N_13591);
nand U13927 (N_13927,N_13595,N_13547);
nand U13928 (N_13928,N_13609,N_13661);
or U13929 (N_13929,N_13520,N_13554);
xor U13930 (N_13930,N_13686,N_13588);
nand U13931 (N_13931,N_13742,N_13672);
and U13932 (N_13932,N_13648,N_13506);
nor U13933 (N_13933,N_13582,N_13722);
nand U13934 (N_13934,N_13525,N_13700);
nand U13935 (N_13935,N_13535,N_13711);
xnor U13936 (N_13936,N_13592,N_13728);
and U13937 (N_13937,N_13687,N_13515);
nor U13938 (N_13938,N_13601,N_13622);
xor U13939 (N_13939,N_13685,N_13630);
nand U13940 (N_13940,N_13743,N_13567);
and U13941 (N_13941,N_13685,N_13631);
xor U13942 (N_13942,N_13697,N_13634);
and U13943 (N_13943,N_13554,N_13666);
nor U13944 (N_13944,N_13647,N_13711);
xor U13945 (N_13945,N_13564,N_13631);
xor U13946 (N_13946,N_13696,N_13698);
and U13947 (N_13947,N_13506,N_13567);
xor U13948 (N_13948,N_13569,N_13743);
and U13949 (N_13949,N_13522,N_13576);
or U13950 (N_13950,N_13617,N_13674);
xnor U13951 (N_13951,N_13714,N_13579);
nor U13952 (N_13952,N_13602,N_13722);
nand U13953 (N_13953,N_13598,N_13563);
and U13954 (N_13954,N_13691,N_13504);
and U13955 (N_13955,N_13690,N_13679);
or U13956 (N_13956,N_13657,N_13601);
xor U13957 (N_13957,N_13730,N_13557);
or U13958 (N_13958,N_13637,N_13675);
nor U13959 (N_13959,N_13659,N_13551);
nand U13960 (N_13960,N_13719,N_13732);
nand U13961 (N_13961,N_13625,N_13740);
nor U13962 (N_13962,N_13624,N_13635);
nor U13963 (N_13963,N_13575,N_13645);
and U13964 (N_13964,N_13629,N_13643);
or U13965 (N_13965,N_13640,N_13742);
and U13966 (N_13966,N_13560,N_13683);
and U13967 (N_13967,N_13702,N_13560);
or U13968 (N_13968,N_13501,N_13607);
or U13969 (N_13969,N_13623,N_13528);
nand U13970 (N_13970,N_13720,N_13650);
xnor U13971 (N_13971,N_13626,N_13698);
xnor U13972 (N_13972,N_13689,N_13513);
and U13973 (N_13973,N_13664,N_13689);
nor U13974 (N_13974,N_13560,N_13681);
and U13975 (N_13975,N_13681,N_13508);
nor U13976 (N_13976,N_13592,N_13540);
nor U13977 (N_13977,N_13506,N_13546);
and U13978 (N_13978,N_13598,N_13589);
nor U13979 (N_13979,N_13713,N_13684);
or U13980 (N_13980,N_13605,N_13685);
xor U13981 (N_13981,N_13589,N_13553);
and U13982 (N_13982,N_13680,N_13559);
nand U13983 (N_13983,N_13667,N_13643);
or U13984 (N_13984,N_13622,N_13602);
nor U13985 (N_13985,N_13733,N_13557);
or U13986 (N_13986,N_13606,N_13698);
or U13987 (N_13987,N_13529,N_13669);
xnor U13988 (N_13988,N_13644,N_13528);
or U13989 (N_13989,N_13662,N_13748);
nand U13990 (N_13990,N_13632,N_13743);
nand U13991 (N_13991,N_13620,N_13688);
and U13992 (N_13992,N_13682,N_13696);
xnor U13993 (N_13993,N_13553,N_13646);
or U13994 (N_13994,N_13577,N_13563);
nor U13995 (N_13995,N_13557,N_13632);
or U13996 (N_13996,N_13723,N_13513);
and U13997 (N_13997,N_13583,N_13597);
xor U13998 (N_13998,N_13510,N_13508);
nor U13999 (N_13999,N_13638,N_13615);
or U14000 (N_14000,N_13776,N_13777);
nor U14001 (N_14001,N_13768,N_13881);
nor U14002 (N_14002,N_13950,N_13868);
and U14003 (N_14003,N_13965,N_13767);
nand U14004 (N_14004,N_13949,N_13864);
nand U14005 (N_14005,N_13945,N_13972);
or U14006 (N_14006,N_13880,N_13981);
nand U14007 (N_14007,N_13826,N_13982);
xor U14008 (N_14008,N_13919,N_13835);
xor U14009 (N_14009,N_13855,N_13967);
or U14010 (N_14010,N_13993,N_13874);
xor U14011 (N_14011,N_13805,N_13912);
nand U14012 (N_14012,N_13947,N_13812);
xor U14013 (N_14013,N_13964,N_13936);
nand U14014 (N_14014,N_13802,N_13778);
nand U14015 (N_14015,N_13848,N_13910);
nand U14016 (N_14016,N_13951,N_13896);
nor U14017 (N_14017,N_13895,N_13761);
xnor U14018 (N_14018,N_13774,N_13992);
or U14019 (N_14019,N_13892,N_13760);
or U14020 (N_14020,N_13833,N_13997);
and U14021 (N_14021,N_13753,N_13819);
nand U14022 (N_14022,N_13754,N_13946);
xnor U14023 (N_14023,N_13983,N_13773);
or U14024 (N_14024,N_13934,N_13929);
and U14025 (N_14025,N_13762,N_13764);
and U14026 (N_14026,N_13884,N_13822);
xnor U14027 (N_14027,N_13867,N_13901);
nand U14028 (N_14028,N_13834,N_13963);
nand U14029 (N_14029,N_13861,N_13968);
or U14030 (N_14030,N_13866,N_13783);
nor U14031 (N_14031,N_13841,N_13932);
or U14032 (N_14032,N_13844,N_13978);
nor U14033 (N_14033,N_13837,N_13926);
nand U14034 (N_14034,N_13839,N_13890);
xnor U14035 (N_14035,N_13820,N_13853);
nor U14036 (N_14036,N_13869,N_13821);
or U14037 (N_14037,N_13977,N_13914);
and U14038 (N_14038,N_13898,N_13921);
nor U14039 (N_14039,N_13860,N_13856);
xor U14040 (N_14040,N_13800,N_13911);
or U14041 (N_14041,N_13976,N_13799);
nand U14042 (N_14042,N_13899,N_13902);
or U14043 (N_14043,N_13924,N_13813);
nor U14044 (N_14044,N_13918,N_13888);
or U14045 (N_14045,N_13958,N_13771);
and U14046 (N_14046,N_13938,N_13830);
and U14047 (N_14047,N_13999,N_13765);
xor U14048 (N_14048,N_13883,N_13779);
xor U14049 (N_14049,N_13859,N_13757);
or U14050 (N_14050,N_13996,N_13810);
nand U14051 (N_14051,N_13956,N_13786);
nand U14052 (N_14052,N_13877,N_13785);
and U14053 (N_14053,N_13903,N_13980);
nor U14054 (N_14054,N_13940,N_13916);
xnor U14055 (N_14055,N_13900,N_13782);
xor U14056 (N_14056,N_13935,N_13905);
xor U14057 (N_14057,N_13792,N_13970);
and U14058 (N_14058,N_13758,N_13876);
and U14059 (N_14059,N_13960,N_13751);
and U14060 (N_14060,N_13770,N_13807);
nand U14061 (N_14061,N_13991,N_13794);
xor U14062 (N_14062,N_13811,N_13838);
nand U14063 (N_14063,N_13781,N_13897);
nor U14064 (N_14064,N_13763,N_13878);
or U14065 (N_14065,N_13939,N_13825);
nand U14066 (N_14066,N_13818,N_13986);
nor U14067 (N_14067,N_13942,N_13827);
and U14068 (N_14068,N_13840,N_13941);
nand U14069 (N_14069,N_13850,N_13784);
or U14070 (N_14070,N_13831,N_13962);
and U14071 (N_14071,N_13790,N_13974);
or U14072 (N_14072,N_13985,N_13971);
and U14073 (N_14073,N_13828,N_13804);
and U14074 (N_14074,N_13930,N_13922);
nand U14075 (N_14075,N_13766,N_13843);
nor U14076 (N_14076,N_13824,N_13961);
xor U14077 (N_14077,N_13882,N_13927);
nor U14078 (N_14078,N_13858,N_13920);
nor U14079 (N_14079,N_13873,N_13943);
xor U14080 (N_14080,N_13886,N_13852);
and U14081 (N_14081,N_13787,N_13756);
nand U14082 (N_14082,N_13775,N_13988);
xor U14083 (N_14083,N_13772,N_13979);
xor U14084 (N_14084,N_13798,N_13891);
and U14085 (N_14085,N_13832,N_13944);
and U14086 (N_14086,N_13955,N_13809);
or U14087 (N_14087,N_13925,N_13842);
and U14088 (N_14088,N_13803,N_13863);
and U14089 (N_14089,N_13928,N_13788);
or U14090 (N_14090,N_13917,N_13847);
xor U14091 (N_14091,N_13857,N_13865);
and U14092 (N_14092,N_13854,N_13937);
nand U14093 (N_14093,N_13814,N_13871);
and U14094 (N_14094,N_13795,N_13875);
nor U14095 (N_14095,N_13849,N_13987);
nor U14096 (N_14096,N_13904,N_13801);
xnor U14097 (N_14097,N_13957,N_13894);
nand U14098 (N_14098,N_13907,N_13879);
nor U14099 (N_14099,N_13923,N_13984);
or U14100 (N_14100,N_13780,N_13887);
and U14101 (N_14101,N_13906,N_13952);
or U14102 (N_14102,N_13889,N_13908);
and U14103 (N_14103,N_13969,N_13829);
nand U14104 (N_14104,N_13870,N_13851);
nor U14105 (N_14105,N_13793,N_13750);
nand U14106 (N_14106,N_13846,N_13862);
and U14107 (N_14107,N_13759,N_13975);
nor U14108 (N_14108,N_13959,N_13808);
and U14109 (N_14109,N_13994,N_13933);
or U14110 (N_14110,N_13872,N_13796);
nor U14111 (N_14111,N_13752,N_13948);
nor U14112 (N_14112,N_13806,N_13954);
or U14113 (N_14113,N_13990,N_13953);
nand U14114 (N_14114,N_13769,N_13995);
and U14115 (N_14115,N_13797,N_13915);
nor U14116 (N_14116,N_13817,N_13913);
nand U14117 (N_14117,N_13885,N_13791);
and U14118 (N_14118,N_13931,N_13823);
and U14119 (N_14119,N_13816,N_13755);
xor U14120 (N_14120,N_13815,N_13998);
or U14121 (N_14121,N_13973,N_13789);
or U14122 (N_14122,N_13845,N_13989);
nor U14123 (N_14123,N_13836,N_13893);
nor U14124 (N_14124,N_13966,N_13909);
nand U14125 (N_14125,N_13860,N_13813);
nand U14126 (N_14126,N_13810,N_13891);
or U14127 (N_14127,N_13911,N_13966);
nor U14128 (N_14128,N_13888,N_13922);
and U14129 (N_14129,N_13897,N_13983);
nand U14130 (N_14130,N_13777,N_13786);
xor U14131 (N_14131,N_13908,N_13904);
xor U14132 (N_14132,N_13771,N_13907);
or U14133 (N_14133,N_13833,N_13882);
xor U14134 (N_14134,N_13922,N_13829);
or U14135 (N_14135,N_13937,N_13812);
and U14136 (N_14136,N_13753,N_13944);
or U14137 (N_14137,N_13891,N_13953);
and U14138 (N_14138,N_13873,N_13888);
and U14139 (N_14139,N_13996,N_13778);
nor U14140 (N_14140,N_13883,N_13896);
xor U14141 (N_14141,N_13771,N_13879);
and U14142 (N_14142,N_13790,N_13883);
or U14143 (N_14143,N_13851,N_13947);
xor U14144 (N_14144,N_13859,N_13753);
nand U14145 (N_14145,N_13984,N_13960);
and U14146 (N_14146,N_13814,N_13950);
xor U14147 (N_14147,N_13977,N_13786);
and U14148 (N_14148,N_13815,N_13867);
nor U14149 (N_14149,N_13894,N_13832);
nor U14150 (N_14150,N_13815,N_13767);
and U14151 (N_14151,N_13897,N_13993);
nor U14152 (N_14152,N_13978,N_13899);
nand U14153 (N_14153,N_13943,N_13871);
nand U14154 (N_14154,N_13778,N_13936);
nor U14155 (N_14155,N_13927,N_13982);
or U14156 (N_14156,N_13858,N_13950);
nand U14157 (N_14157,N_13983,N_13799);
or U14158 (N_14158,N_13973,N_13935);
nand U14159 (N_14159,N_13826,N_13781);
xor U14160 (N_14160,N_13961,N_13778);
or U14161 (N_14161,N_13956,N_13990);
and U14162 (N_14162,N_13878,N_13816);
xnor U14163 (N_14163,N_13815,N_13770);
xor U14164 (N_14164,N_13863,N_13887);
or U14165 (N_14165,N_13995,N_13806);
xnor U14166 (N_14166,N_13855,N_13960);
xnor U14167 (N_14167,N_13757,N_13788);
xor U14168 (N_14168,N_13934,N_13943);
or U14169 (N_14169,N_13979,N_13753);
nand U14170 (N_14170,N_13762,N_13952);
nor U14171 (N_14171,N_13865,N_13793);
or U14172 (N_14172,N_13921,N_13938);
or U14173 (N_14173,N_13909,N_13888);
xor U14174 (N_14174,N_13921,N_13776);
nor U14175 (N_14175,N_13751,N_13769);
xor U14176 (N_14176,N_13961,N_13991);
or U14177 (N_14177,N_13854,N_13840);
nor U14178 (N_14178,N_13824,N_13766);
or U14179 (N_14179,N_13991,N_13811);
or U14180 (N_14180,N_13965,N_13927);
xor U14181 (N_14181,N_13929,N_13768);
xnor U14182 (N_14182,N_13829,N_13906);
nor U14183 (N_14183,N_13921,N_13992);
xor U14184 (N_14184,N_13765,N_13861);
nand U14185 (N_14185,N_13852,N_13844);
nand U14186 (N_14186,N_13981,N_13865);
xnor U14187 (N_14187,N_13782,N_13901);
nand U14188 (N_14188,N_13774,N_13896);
nor U14189 (N_14189,N_13958,N_13825);
or U14190 (N_14190,N_13949,N_13836);
nand U14191 (N_14191,N_13753,N_13758);
and U14192 (N_14192,N_13852,N_13825);
and U14193 (N_14193,N_13833,N_13853);
nor U14194 (N_14194,N_13758,N_13844);
nand U14195 (N_14195,N_13855,N_13790);
nor U14196 (N_14196,N_13934,N_13766);
nor U14197 (N_14197,N_13988,N_13925);
or U14198 (N_14198,N_13835,N_13804);
and U14199 (N_14199,N_13821,N_13835);
nand U14200 (N_14200,N_13958,N_13965);
xnor U14201 (N_14201,N_13964,N_13999);
xnor U14202 (N_14202,N_13937,N_13813);
nor U14203 (N_14203,N_13781,N_13866);
or U14204 (N_14204,N_13854,N_13908);
or U14205 (N_14205,N_13939,N_13984);
and U14206 (N_14206,N_13768,N_13998);
or U14207 (N_14207,N_13975,N_13785);
or U14208 (N_14208,N_13989,N_13898);
nor U14209 (N_14209,N_13884,N_13976);
nand U14210 (N_14210,N_13786,N_13779);
nor U14211 (N_14211,N_13765,N_13777);
nor U14212 (N_14212,N_13907,N_13913);
or U14213 (N_14213,N_13862,N_13883);
nand U14214 (N_14214,N_13843,N_13847);
nand U14215 (N_14215,N_13859,N_13766);
or U14216 (N_14216,N_13766,N_13975);
nand U14217 (N_14217,N_13993,N_13986);
and U14218 (N_14218,N_13756,N_13882);
nand U14219 (N_14219,N_13770,N_13840);
and U14220 (N_14220,N_13856,N_13983);
or U14221 (N_14221,N_13812,N_13929);
nor U14222 (N_14222,N_13984,N_13891);
and U14223 (N_14223,N_13952,N_13880);
nand U14224 (N_14224,N_13854,N_13912);
and U14225 (N_14225,N_13929,N_13833);
nand U14226 (N_14226,N_13853,N_13985);
xnor U14227 (N_14227,N_13820,N_13904);
and U14228 (N_14228,N_13846,N_13910);
xnor U14229 (N_14229,N_13756,N_13975);
and U14230 (N_14230,N_13799,N_13906);
nand U14231 (N_14231,N_13969,N_13830);
nand U14232 (N_14232,N_13943,N_13872);
or U14233 (N_14233,N_13811,N_13954);
or U14234 (N_14234,N_13822,N_13781);
and U14235 (N_14235,N_13901,N_13768);
and U14236 (N_14236,N_13776,N_13981);
nand U14237 (N_14237,N_13754,N_13855);
nand U14238 (N_14238,N_13797,N_13765);
nor U14239 (N_14239,N_13899,N_13805);
and U14240 (N_14240,N_13999,N_13797);
or U14241 (N_14241,N_13971,N_13901);
nand U14242 (N_14242,N_13838,N_13978);
xor U14243 (N_14243,N_13920,N_13998);
or U14244 (N_14244,N_13841,N_13826);
or U14245 (N_14245,N_13891,N_13955);
or U14246 (N_14246,N_13879,N_13857);
and U14247 (N_14247,N_13979,N_13822);
or U14248 (N_14248,N_13776,N_13928);
xnor U14249 (N_14249,N_13841,N_13772);
or U14250 (N_14250,N_14039,N_14207);
nand U14251 (N_14251,N_14075,N_14077);
xor U14252 (N_14252,N_14240,N_14153);
or U14253 (N_14253,N_14095,N_14034);
nand U14254 (N_14254,N_14029,N_14194);
or U14255 (N_14255,N_14241,N_14027);
nor U14256 (N_14256,N_14135,N_14148);
or U14257 (N_14257,N_14230,N_14249);
nand U14258 (N_14258,N_14166,N_14118);
xor U14259 (N_14259,N_14214,N_14035);
xnor U14260 (N_14260,N_14147,N_14248);
nand U14261 (N_14261,N_14141,N_14164);
nor U14262 (N_14262,N_14043,N_14036);
or U14263 (N_14263,N_14012,N_14102);
or U14264 (N_14264,N_14126,N_14243);
or U14265 (N_14265,N_14080,N_14183);
or U14266 (N_14266,N_14023,N_14111);
xor U14267 (N_14267,N_14074,N_14178);
xnor U14268 (N_14268,N_14070,N_14206);
or U14269 (N_14269,N_14175,N_14200);
and U14270 (N_14270,N_14052,N_14062);
nor U14271 (N_14271,N_14142,N_14218);
and U14272 (N_14272,N_14203,N_14184);
or U14273 (N_14273,N_14127,N_14065);
nor U14274 (N_14274,N_14197,N_14071);
xor U14275 (N_14275,N_14172,N_14238);
nand U14276 (N_14276,N_14140,N_14022);
and U14277 (N_14277,N_14201,N_14193);
nor U14278 (N_14278,N_14190,N_14100);
nor U14279 (N_14279,N_14128,N_14056);
nand U14280 (N_14280,N_14078,N_14168);
or U14281 (N_14281,N_14046,N_14146);
or U14282 (N_14282,N_14231,N_14092);
nor U14283 (N_14283,N_14109,N_14158);
nor U14284 (N_14284,N_14076,N_14167);
and U14285 (N_14285,N_14173,N_14122);
xor U14286 (N_14286,N_14234,N_14038);
nand U14287 (N_14287,N_14138,N_14124);
or U14288 (N_14288,N_14223,N_14087);
xor U14289 (N_14289,N_14139,N_14120);
nor U14290 (N_14290,N_14055,N_14174);
and U14291 (N_14291,N_14099,N_14058);
xor U14292 (N_14292,N_14053,N_14179);
nand U14293 (N_14293,N_14073,N_14208);
xor U14294 (N_14294,N_14216,N_14067);
xnor U14295 (N_14295,N_14017,N_14176);
xor U14296 (N_14296,N_14125,N_14050);
and U14297 (N_14297,N_14066,N_14025);
nor U14298 (N_14298,N_14145,N_14237);
or U14299 (N_14299,N_14181,N_14103);
xnor U14300 (N_14300,N_14180,N_14239);
xor U14301 (N_14301,N_14170,N_14221);
or U14302 (N_14302,N_14217,N_14090);
or U14303 (N_14303,N_14032,N_14060);
xnor U14304 (N_14304,N_14160,N_14199);
xor U14305 (N_14305,N_14165,N_14048);
xnor U14306 (N_14306,N_14051,N_14117);
xor U14307 (N_14307,N_14205,N_14169);
nor U14308 (N_14308,N_14245,N_14011);
xor U14309 (N_14309,N_14098,N_14112);
nand U14310 (N_14310,N_14185,N_14150);
or U14311 (N_14311,N_14202,N_14009);
and U14312 (N_14312,N_14049,N_14026);
nand U14313 (N_14313,N_14013,N_14162);
or U14314 (N_14314,N_14123,N_14163);
or U14315 (N_14315,N_14091,N_14044);
nand U14316 (N_14316,N_14161,N_14064);
nand U14317 (N_14317,N_14089,N_14079);
or U14318 (N_14318,N_14024,N_14191);
and U14319 (N_14319,N_14136,N_14041);
xor U14320 (N_14320,N_14008,N_14083);
or U14321 (N_14321,N_14233,N_14110);
and U14322 (N_14322,N_14014,N_14182);
and U14323 (N_14323,N_14229,N_14211);
nand U14324 (N_14324,N_14037,N_14155);
nand U14325 (N_14325,N_14085,N_14005);
nor U14326 (N_14326,N_14000,N_14045);
xor U14327 (N_14327,N_14104,N_14068);
nand U14328 (N_14328,N_14133,N_14059);
nor U14329 (N_14329,N_14131,N_14119);
and U14330 (N_14330,N_14069,N_14016);
nor U14331 (N_14331,N_14130,N_14086);
and U14332 (N_14332,N_14159,N_14084);
or U14333 (N_14333,N_14116,N_14033);
and U14334 (N_14334,N_14219,N_14002);
xor U14335 (N_14335,N_14143,N_14018);
xor U14336 (N_14336,N_14226,N_14157);
nand U14337 (N_14337,N_14031,N_14061);
xor U14338 (N_14338,N_14082,N_14232);
xor U14339 (N_14339,N_14210,N_14105);
or U14340 (N_14340,N_14003,N_14224);
and U14341 (N_14341,N_14154,N_14236);
nand U14342 (N_14342,N_14047,N_14115);
nand U14343 (N_14343,N_14220,N_14187);
nand U14344 (N_14344,N_14010,N_14189);
nor U14345 (N_14345,N_14004,N_14101);
and U14346 (N_14346,N_14088,N_14209);
or U14347 (N_14347,N_14188,N_14129);
nor U14348 (N_14348,N_14212,N_14151);
nand U14349 (N_14349,N_14177,N_14081);
nor U14350 (N_14350,N_14020,N_14108);
nand U14351 (N_14351,N_14192,N_14235);
or U14352 (N_14352,N_14195,N_14096);
or U14353 (N_14353,N_14106,N_14144);
or U14354 (N_14354,N_14019,N_14134);
xor U14355 (N_14355,N_14198,N_14196);
or U14356 (N_14356,N_14006,N_14121);
or U14357 (N_14357,N_14215,N_14152);
and U14358 (N_14358,N_14040,N_14227);
or U14359 (N_14359,N_14007,N_14107);
or U14360 (N_14360,N_14001,N_14042);
xnor U14361 (N_14361,N_14244,N_14030);
xnor U14362 (N_14362,N_14132,N_14093);
and U14363 (N_14363,N_14186,N_14225);
nand U14364 (N_14364,N_14072,N_14213);
and U14365 (N_14365,N_14028,N_14113);
xnor U14366 (N_14366,N_14246,N_14054);
or U14367 (N_14367,N_14242,N_14228);
nor U14368 (N_14368,N_14247,N_14097);
nor U14369 (N_14369,N_14063,N_14204);
xor U14370 (N_14370,N_14057,N_14015);
xor U14371 (N_14371,N_14149,N_14222);
and U14372 (N_14372,N_14156,N_14094);
or U14373 (N_14373,N_14137,N_14171);
and U14374 (N_14374,N_14114,N_14021);
xnor U14375 (N_14375,N_14011,N_14003);
or U14376 (N_14376,N_14157,N_14084);
nand U14377 (N_14377,N_14013,N_14149);
nor U14378 (N_14378,N_14123,N_14138);
nor U14379 (N_14379,N_14012,N_14247);
or U14380 (N_14380,N_14241,N_14066);
or U14381 (N_14381,N_14181,N_14135);
and U14382 (N_14382,N_14159,N_14245);
xnor U14383 (N_14383,N_14212,N_14198);
and U14384 (N_14384,N_14213,N_14107);
and U14385 (N_14385,N_14040,N_14068);
and U14386 (N_14386,N_14065,N_14157);
nand U14387 (N_14387,N_14033,N_14175);
and U14388 (N_14388,N_14170,N_14061);
or U14389 (N_14389,N_14000,N_14227);
and U14390 (N_14390,N_14010,N_14229);
nand U14391 (N_14391,N_14188,N_14091);
nor U14392 (N_14392,N_14099,N_14248);
and U14393 (N_14393,N_14243,N_14010);
and U14394 (N_14394,N_14019,N_14012);
nor U14395 (N_14395,N_14075,N_14047);
or U14396 (N_14396,N_14231,N_14170);
and U14397 (N_14397,N_14016,N_14100);
and U14398 (N_14398,N_14123,N_14050);
and U14399 (N_14399,N_14069,N_14188);
nand U14400 (N_14400,N_14048,N_14191);
nand U14401 (N_14401,N_14249,N_14189);
or U14402 (N_14402,N_14023,N_14186);
xnor U14403 (N_14403,N_14187,N_14188);
or U14404 (N_14404,N_14125,N_14182);
nand U14405 (N_14405,N_14132,N_14029);
or U14406 (N_14406,N_14128,N_14052);
nand U14407 (N_14407,N_14180,N_14086);
nand U14408 (N_14408,N_14138,N_14025);
xnor U14409 (N_14409,N_14205,N_14125);
nor U14410 (N_14410,N_14149,N_14052);
nor U14411 (N_14411,N_14122,N_14045);
nand U14412 (N_14412,N_14133,N_14132);
nand U14413 (N_14413,N_14176,N_14233);
nand U14414 (N_14414,N_14204,N_14228);
nor U14415 (N_14415,N_14130,N_14001);
nor U14416 (N_14416,N_14029,N_14108);
and U14417 (N_14417,N_14239,N_14205);
and U14418 (N_14418,N_14204,N_14173);
and U14419 (N_14419,N_14124,N_14132);
xnor U14420 (N_14420,N_14080,N_14228);
xnor U14421 (N_14421,N_14213,N_14123);
nor U14422 (N_14422,N_14208,N_14151);
nor U14423 (N_14423,N_14162,N_14190);
and U14424 (N_14424,N_14117,N_14098);
xnor U14425 (N_14425,N_14065,N_14130);
or U14426 (N_14426,N_14102,N_14122);
and U14427 (N_14427,N_14053,N_14075);
xor U14428 (N_14428,N_14115,N_14055);
xor U14429 (N_14429,N_14168,N_14217);
xnor U14430 (N_14430,N_14154,N_14129);
nand U14431 (N_14431,N_14247,N_14085);
or U14432 (N_14432,N_14005,N_14089);
nor U14433 (N_14433,N_14088,N_14052);
xor U14434 (N_14434,N_14223,N_14188);
xnor U14435 (N_14435,N_14175,N_14191);
or U14436 (N_14436,N_14243,N_14217);
nor U14437 (N_14437,N_14001,N_14111);
and U14438 (N_14438,N_14069,N_14072);
xor U14439 (N_14439,N_14207,N_14232);
nand U14440 (N_14440,N_14067,N_14171);
nand U14441 (N_14441,N_14199,N_14195);
nor U14442 (N_14442,N_14107,N_14055);
nand U14443 (N_14443,N_14068,N_14114);
and U14444 (N_14444,N_14130,N_14057);
nand U14445 (N_14445,N_14222,N_14096);
xnor U14446 (N_14446,N_14086,N_14136);
xnor U14447 (N_14447,N_14216,N_14093);
and U14448 (N_14448,N_14091,N_14085);
or U14449 (N_14449,N_14109,N_14027);
and U14450 (N_14450,N_14202,N_14195);
nand U14451 (N_14451,N_14115,N_14013);
xor U14452 (N_14452,N_14193,N_14237);
nor U14453 (N_14453,N_14237,N_14115);
xor U14454 (N_14454,N_14092,N_14062);
nor U14455 (N_14455,N_14112,N_14246);
nand U14456 (N_14456,N_14021,N_14231);
and U14457 (N_14457,N_14167,N_14056);
nand U14458 (N_14458,N_14178,N_14087);
or U14459 (N_14459,N_14174,N_14185);
nand U14460 (N_14460,N_14190,N_14231);
nand U14461 (N_14461,N_14234,N_14246);
and U14462 (N_14462,N_14155,N_14237);
nand U14463 (N_14463,N_14072,N_14190);
or U14464 (N_14464,N_14151,N_14190);
and U14465 (N_14465,N_14013,N_14125);
xor U14466 (N_14466,N_14065,N_14114);
or U14467 (N_14467,N_14095,N_14051);
nor U14468 (N_14468,N_14062,N_14226);
and U14469 (N_14469,N_14012,N_14036);
xor U14470 (N_14470,N_14174,N_14067);
nand U14471 (N_14471,N_14195,N_14240);
and U14472 (N_14472,N_14067,N_14166);
nor U14473 (N_14473,N_14146,N_14114);
nand U14474 (N_14474,N_14094,N_14095);
and U14475 (N_14475,N_14039,N_14176);
or U14476 (N_14476,N_14178,N_14133);
nand U14477 (N_14477,N_14178,N_14226);
xnor U14478 (N_14478,N_14007,N_14124);
and U14479 (N_14479,N_14191,N_14147);
xor U14480 (N_14480,N_14030,N_14167);
and U14481 (N_14481,N_14063,N_14108);
or U14482 (N_14482,N_14023,N_14126);
nand U14483 (N_14483,N_14176,N_14201);
xor U14484 (N_14484,N_14016,N_14127);
xnor U14485 (N_14485,N_14103,N_14011);
nand U14486 (N_14486,N_14111,N_14014);
and U14487 (N_14487,N_14027,N_14097);
nand U14488 (N_14488,N_14013,N_14072);
xor U14489 (N_14489,N_14042,N_14043);
or U14490 (N_14490,N_14206,N_14073);
xor U14491 (N_14491,N_14246,N_14057);
nor U14492 (N_14492,N_14231,N_14019);
nor U14493 (N_14493,N_14150,N_14072);
nor U14494 (N_14494,N_14245,N_14089);
xnor U14495 (N_14495,N_14075,N_14202);
xor U14496 (N_14496,N_14148,N_14117);
or U14497 (N_14497,N_14074,N_14029);
xnor U14498 (N_14498,N_14129,N_14193);
or U14499 (N_14499,N_14131,N_14234);
nand U14500 (N_14500,N_14453,N_14332);
xor U14501 (N_14501,N_14283,N_14304);
and U14502 (N_14502,N_14279,N_14340);
nor U14503 (N_14503,N_14345,N_14309);
and U14504 (N_14504,N_14342,N_14413);
nand U14505 (N_14505,N_14465,N_14344);
nand U14506 (N_14506,N_14468,N_14299);
xor U14507 (N_14507,N_14323,N_14356);
nand U14508 (N_14508,N_14321,N_14372);
and U14509 (N_14509,N_14290,N_14254);
nand U14510 (N_14510,N_14302,N_14359);
or U14511 (N_14511,N_14445,N_14261);
xor U14512 (N_14512,N_14423,N_14441);
xnor U14513 (N_14513,N_14449,N_14410);
xnor U14514 (N_14514,N_14466,N_14292);
nor U14515 (N_14515,N_14409,N_14471);
nand U14516 (N_14516,N_14310,N_14399);
xnor U14517 (N_14517,N_14333,N_14252);
or U14518 (N_14518,N_14262,N_14335);
nor U14519 (N_14519,N_14434,N_14398);
xnor U14520 (N_14520,N_14438,N_14381);
or U14521 (N_14521,N_14319,N_14388);
nor U14522 (N_14522,N_14464,N_14357);
nor U14523 (N_14523,N_14426,N_14267);
nor U14524 (N_14524,N_14336,N_14461);
nor U14525 (N_14525,N_14355,N_14295);
and U14526 (N_14526,N_14311,N_14322);
nand U14527 (N_14527,N_14324,N_14286);
nor U14528 (N_14528,N_14268,N_14258);
nand U14529 (N_14529,N_14493,N_14264);
or U14530 (N_14530,N_14462,N_14368);
and U14531 (N_14531,N_14376,N_14492);
xnor U14532 (N_14532,N_14424,N_14451);
xnor U14533 (N_14533,N_14288,N_14430);
nand U14534 (N_14534,N_14411,N_14259);
nand U14535 (N_14535,N_14384,N_14421);
xnor U14536 (N_14536,N_14369,N_14488);
xor U14537 (N_14537,N_14425,N_14494);
or U14538 (N_14538,N_14270,N_14379);
xnor U14539 (N_14539,N_14457,N_14330);
nand U14540 (N_14540,N_14337,N_14275);
or U14541 (N_14541,N_14392,N_14354);
and U14542 (N_14542,N_14440,N_14377);
or U14543 (N_14543,N_14469,N_14452);
nor U14544 (N_14544,N_14325,N_14403);
nand U14545 (N_14545,N_14467,N_14269);
xor U14546 (N_14546,N_14484,N_14439);
xor U14547 (N_14547,N_14300,N_14414);
xor U14548 (N_14548,N_14273,N_14334);
and U14549 (N_14549,N_14412,N_14459);
and U14550 (N_14550,N_14408,N_14393);
nand U14551 (N_14551,N_14478,N_14378);
xor U14552 (N_14552,N_14437,N_14353);
or U14553 (N_14553,N_14455,N_14475);
xnor U14554 (N_14554,N_14301,N_14317);
nand U14555 (N_14555,N_14266,N_14431);
or U14556 (N_14556,N_14397,N_14297);
or U14557 (N_14557,N_14497,N_14479);
xor U14558 (N_14558,N_14486,N_14447);
xnor U14559 (N_14559,N_14442,N_14489);
nor U14560 (N_14560,N_14362,N_14390);
and U14561 (N_14561,N_14422,N_14443);
nor U14562 (N_14562,N_14343,N_14260);
or U14563 (N_14563,N_14482,N_14491);
and U14564 (N_14564,N_14281,N_14418);
and U14565 (N_14565,N_14305,N_14473);
nand U14566 (N_14566,N_14320,N_14396);
and U14567 (N_14567,N_14298,N_14276);
nand U14568 (N_14568,N_14285,N_14278);
nand U14569 (N_14569,N_14394,N_14454);
and U14570 (N_14570,N_14307,N_14282);
or U14571 (N_14571,N_14406,N_14402);
or U14572 (N_14572,N_14389,N_14327);
or U14573 (N_14573,N_14253,N_14433);
nor U14574 (N_14574,N_14487,N_14428);
or U14575 (N_14575,N_14289,N_14458);
nor U14576 (N_14576,N_14280,N_14456);
and U14577 (N_14577,N_14374,N_14287);
and U14578 (N_14578,N_14460,N_14367);
and U14579 (N_14579,N_14271,N_14407);
and U14580 (N_14580,N_14485,N_14293);
and U14581 (N_14581,N_14348,N_14391);
nand U14582 (N_14582,N_14251,N_14315);
or U14583 (N_14583,N_14498,N_14364);
or U14584 (N_14584,N_14395,N_14387);
or U14585 (N_14585,N_14417,N_14480);
nand U14586 (N_14586,N_14339,N_14420);
nand U14587 (N_14587,N_14366,N_14470);
nand U14588 (N_14588,N_14419,N_14274);
nand U14589 (N_14589,N_14306,N_14316);
xnor U14590 (N_14590,N_14415,N_14263);
nand U14591 (N_14591,N_14256,N_14435);
nor U14592 (N_14592,N_14477,N_14463);
nor U14593 (N_14593,N_14446,N_14382);
xnor U14594 (N_14594,N_14352,N_14296);
nor U14595 (N_14595,N_14350,N_14481);
and U14596 (N_14596,N_14404,N_14351);
xnor U14597 (N_14597,N_14432,N_14483);
nand U14598 (N_14598,N_14294,N_14265);
and U14599 (N_14599,N_14429,N_14401);
nor U14600 (N_14600,N_14318,N_14365);
or U14601 (N_14601,N_14371,N_14346);
nor U14602 (N_14602,N_14328,N_14495);
nand U14603 (N_14603,N_14284,N_14448);
or U14604 (N_14604,N_14370,N_14326);
nor U14605 (N_14605,N_14312,N_14380);
and U14606 (N_14606,N_14331,N_14375);
nand U14607 (N_14607,N_14361,N_14386);
nor U14608 (N_14608,N_14474,N_14250);
nor U14609 (N_14609,N_14363,N_14405);
xnor U14610 (N_14610,N_14476,N_14303);
and U14611 (N_14611,N_14329,N_14313);
xor U14612 (N_14612,N_14450,N_14490);
nor U14613 (N_14613,N_14496,N_14349);
nor U14614 (N_14614,N_14291,N_14255);
or U14615 (N_14615,N_14277,N_14338);
nor U14616 (N_14616,N_14358,N_14499);
or U14617 (N_14617,N_14308,N_14436);
or U14618 (N_14618,N_14341,N_14272);
xnor U14619 (N_14619,N_14257,N_14383);
and U14620 (N_14620,N_14385,N_14472);
nor U14621 (N_14621,N_14444,N_14416);
and U14622 (N_14622,N_14314,N_14360);
nor U14623 (N_14623,N_14400,N_14427);
nor U14624 (N_14624,N_14373,N_14347);
xor U14625 (N_14625,N_14315,N_14472);
nor U14626 (N_14626,N_14436,N_14278);
nand U14627 (N_14627,N_14331,N_14389);
or U14628 (N_14628,N_14488,N_14442);
xnor U14629 (N_14629,N_14295,N_14367);
nand U14630 (N_14630,N_14457,N_14420);
xor U14631 (N_14631,N_14333,N_14338);
and U14632 (N_14632,N_14350,N_14478);
nand U14633 (N_14633,N_14461,N_14311);
or U14634 (N_14634,N_14267,N_14470);
xnor U14635 (N_14635,N_14330,N_14322);
xor U14636 (N_14636,N_14311,N_14389);
xnor U14637 (N_14637,N_14324,N_14469);
nand U14638 (N_14638,N_14385,N_14486);
nor U14639 (N_14639,N_14392,N_14424);
and U14640 (N_14640,N_14323,N_14272);
and U14641 (N_14641,N_14341,N_14444);
nand U14642 (N_14642,N_14406,N_14467);
xor U14643 (N_14643,N_14429,N_14456);
xnor U14644 (N_14644,N_14389,N_14399);
or U14645 (N_14645,N_14341,N_14450);
nor U14646 (N_14646,N_14273,N_14365);
nor U14647 (N_14647,N_14436,N_14335);
nand U14648 (N_14648,N_14334,N_14264);
xor U14649 (N_14649,N_14358,N_14451);
or U14650 (N_14650,N_14444,N_14347);
xor U14651 (N_14651,N_14451,N_14492);
and U14652 (N_14652,N_14469,N_14387);
nor U14653 (N_14653,N_14404,N_14378);
nand U14654 (N_14654,N_14419,N_14476);
xnor U14655 (N_14655,N_14277,N_14380);
and U14656 (N_14656,N_14444,N_14337);
or U14657 (N_14657,N_14305,N_14477);
xnor U14658 (N_14658,N_14327,N_14344);
and U14659 (N_14659,N_14378,N_14332);
nand U14660 (N_14660,N_14475,N_14331);
and U14661 (N_14661,N_14274,N_14424);
nor U14662 (N_14662,N_14277,N_14254);
nor U14663 (N_14663,N_14396,N_14499);
or U14664 (N_14664,N_14404,N_14402);
xnor U14665 (N_14665,N_14437,N_14362);
and U14666 (N_14666,N_14483,N_14479);
nor U14667 (N_14667,N_14487,N_14291);
xor U14668 (N_14668,N_14330,N_14417);
or U14669 (N_14669,N_14376,N_14496);
nor U14670 (N_14670,N_14491,N_14286);
xnor U14671 (N_14671,N_14289,N_14435);
nor U14672 (N_14672,N_14252,N_14458);
nand U14673 (N_14673,N_14386,N_14339);
xnor U14674 (N_14674,N_14426,N_14341);
xor U14675 (N_14675,N_14376,N_14401);
and U14676 (N_14676,N_14269,N_14443);
xnor U14677 (N_14677,N_14391,N_14401);
nand U14678 (N_14678,N_14381,N_14337);
and U14679 (N_14679,N_14425,N_14291);
or U14680 (N_14680,N_14304,N_14295);
xnor U14681 (N_14681,N_14366,N_14323);
and U14682 (N_14682,N_14422,N_14458);
and U14683 (N_14683,N_14370,N_14404);
nand U14684 (N_14684,N_14441,N_14321);
nand U14685 (N_14685,N_14284,N_14476);
xor U14686 (N_14686,N_14402,N_14382);
nand U14687 (N_14687,N_14339,N_14361);
or U14688 (N_14688,N_14439,N_14348);
nor U14689 (N_14689,N_14410,N_14373);
nor U14690 (N_14690,N_14313,N_14285);
or U14691 (N_14691,N_14316,N_14494);
nand U14692 (N_14692,N_14292,N_14296);
or U14693 (N_14693,N_14357,N_14250);
xor U14694 (N_14694,N_14427,N_14279);
nor U14695 (N_14695,N_14260,N_14251);
and U14696 (N_14696,N_14421,N_14460);
or U14697 (N_14697,N_14481,N_14290);
nand U14698 (N_14698,N_14278,N_14262);
nor U14699 (N_14699,N_14250,N_14251);
or U14700 (N_14700,N_14372,N_14423);
and U14701 (N_14701,N_14419,N_14282);
xor U14702 (N_14702,N_14342,N_14365);
nand U14703 (N_14703,N_14303,N_14285);
nand U14704 (N_14704,N_14411,N_14289);
nand U14705 (N_14705,N_14382,N_14406);
xnor U14706 (N_14706,N_14462,N_14372);
xnor U14707 (N_14707,N_14427,N_14422);
xor U14708 (N_14708,N_14370,N_14491);
nor U14709 (N_14709,N_14436,N_14371);
or U14710 (N_14710,N_14445,N_14258);
and U14711 (N_14711,N_14443,N_14365);
or U14712 (N_14712,N_14495,N_14410);
or U14713 (N_14713,N_14461,N_14329);
xnor U14714 (N_14714,N_14390,N_14345);
nand U14715 (N_14715,N_14367,N_14457);
and U14716 (N_14716,N_14433,N_14332);
or U14717 (N_14717,N_14269,N_14398);
nand U14718 (N_14718,N_14356,N_14284);
xor U14719 (N_14719,N_14449,N_14432);
xnor U14720 (N_14720,N_14342,N_14309);
or U14721 (N_14721,N_14481,N_14440);
and U14722 (N_14722,N_14267,N_14266);
and U14723 (N_14723,N_14276,N_14337);
nand U14724 (N_14724,N_14394,N_14267);
nand U14725 (N_14725,N_14288,N_14484);
nand U14726 (N_14726,N_14464,N_14458);
and U14727 (N_14727,N_14395,N_14319);
or U14728 (N_14728,N_14273,N_14497);
nand U14729 (N_14729,N_14285,N_14389);
and U14730 (N_14730,N_14428,N_14380);
nor U14731 (N_14731,N_14406,N_14253);
xor U14732 (N_14732,N_14464,N_14309);
nand U14733 (N_14733,N_14328,N_14471);
nor U14734 (N_14734,N_14342,N_14337);
nand U14735 (N_14735,N_14487,N_14446);
or U14736 (N_14736,N_14378,N_14483);
nand U14737 (N_14737,N_14468,N_14339);
xnor U14738 (N_14738,N_14411,N_14276);
or U14739 (N_14739,N_14332,N_14350);
or U14740 (N_14740,N_14366,N_14428);
nor U14741 (N_14741,N_14296,N_14471);
and U14742 (N_14742,N_14464,N_14362);
xnor U14743 (N_14743,N_14354,N_14403);
xnor U14744 (N_14744,N_14262,N_14449);
nor U14745 (N_14745,N_14471,N_14417);
xnor U14746 (N_14746,N_14499,N_14280);
xor U14747 (N_14747,N_14303,N_14320);
nor U14748 (N_14748,N_14482,N_14287);
and U14749 (N_14749,N_14262,N_14434);
nor U14750 (N_14750,N_14708,N_14705);
nand U14751 (N_14751,N_14687,N_14656);
nand U14752 (N_14752,N_14574,N_14552);
and U14753 (N_14753,N_14589,N_14738);
nor U14754 (N_14754,N_14633,N_14704);
xor U14755 (N_14755,N_14565,N_14606);
nand U14756 (N_14756,N_14679,N_14509);
or U14757 (N_14757,N_14542,N_14570);
nor U14758 (N_14758,N_14683,N_14594);
nand U14759 (N_14759,N_14528,N_14666);
nand U14760 (N_14760,N_14616,N_14518);
nor U14761 (N_14761,N_14661,N_14722);
and U14762 (N_14762,N_14662,N_14619);
or U14763 (N_14763,N_14506,N_14676);
xnor U14764 (N_14764,N_14572,N_14688);
nor U14765 (N_14765,N_14669,N_14527);
nand U14766 (N_14766,N_14733,N_14674);
nand U14767 (N_14767,N_14573,N_14747);
xor U14768 (N_14768,N_14595,N_14627);
and U14769 (N_14769,N_14699,N_14504);
nor U14770 (N_14770,N_14582,N_14678);
and U14771 (N_14771,N_14701,N_14710);
nor U14772 (N_14772,N_14618,N_14569);
xor U14773 (N_14773,N_14501,N_14728);
nand U14774 (N_14774,N_14653,N_14588);
and U14775 (N_14775,N_14671,N_14713);
nor U14776 (N_14776,N_14717,N_14643);
nand U14777 (N_14777,N_14673,N_14514);
or U14778 (N_14778,N_14657,N_14607);
or U14779 (N_14779,N_14742,N_14736);
xnor U14780 (N_14780,N_14567,N_14651);
nor U14781 (N_14781,N_14608,N_14693);
and U14782 (N_14782,N_14591,N_14700);
and U14783 (N_14783,N_14571,N_14744);
and U14784 (N_14784,N_14556,N_14706);
and U14785 (N_14785,N_14525,N_14500);
or U14786 (N_14786,N_14549,N_14531);
nor U14787 (N_14787,N_14642,N_14630);
xor U14788 (N_14788,N_14536,N_14603);
and U14789 (N_14789,N_14548,N_14545);
xnor U14790 (N_14790,N_14614,N_14557);
xor U14791 (N_14791,N_14602,N_14513);
or U14792 (N_14792,N_14696,N_14709);
nor U14793 (N_14793,N_14748,N_14597);
nor U14794 (N_14794,N_14724,N_14519);
xor U14795 (N_14795,N_14664,N_14625);
nor U14796 (N_14796,N_14532,N_14732);
or U14797 (N_14797,N_14530,N_14712);
nor U14798 (N_14798,N_14741,N_14659);
xor U14799 (N_14799,N_14655,N_14621);
and U14800 (N_14800,N_14521,N_14533);
xnor U14801 (N_14801,N_14635,N_14730);
nand U14802 (N_14802,N_14576,N_14707);
nor U14803 (N_14803,N_14507,N_14610);
or U14804 (N_14804,N_14586,N_14613);
xor U14805 (N_14805,N_14541,N_14740);
xor U14806 (N_14806,N_14640,N_14714);
nor U14807 (N_14807,N_14539,N_14590);
xor U14808 (N_14808,N_14604,N_14680);
and U14809 (N_14809,N_14677,N_14524);
nor U14810 (N_14810,N_14537,N_14681);
nand U14811 (N_14811,N_14638,N_14660);
or U14812 (N_14812,N_14534,N_14727);
and U14813 (N_14813,N_14526,N_14502);
xor U14814 (N_14814,N_14726,N_14566);
nand U14815 (N_14815,N_14652,N_14617);
and U14816 (N_14816,N_14550,N_14731);
or U14817 (N_14817,N_14670,N_14698);
xnor U14818 (N_14818,N_14682,N_14596);
nand U14819 (N_14819,N_14649,N_14538);
nand U14820 (N_14820,N_14592,N_14675);
nand U14821 (N_14821,N_14644,N_14515);
nor U14822 (N_14822,N_14721,N_14665);
nor U14823 (N_14823,N_14720,N_14637);
and U14824 (N_14824,N_14559,N_14739);
nand U14825 (N_14825,N_14737,N_14568);
and U14826 (N_14826,N_14612,N_14563);
or U14827 (N_14827,N_14690,N_14746);
or U14828 (N_14828,N_14689,N_14650);
nand U14829 (N_14829,N_14697,N_14729);
or U14830 (N_14830,N_14648,N_14555);
or U14831 (N_14831,N_14646,N_14522);
xnor U14832 (N_14832,N_14749,N_14520);
nor U14833 (N_14833,N_14641,N_14562);
and U14834 (N_14834,N_14702,N_14654);
nand U14835 (N_14835,N_14624,N_14577);
or U14836 (N_14836,N_14636,N_14584);
nand U14837 (N_14837,N_14523,N_14535);
or U14838 (N_14838,N_14719,N_14672);
nand U14839 (N_14839,N_14626,N_14658);
nand U14840 (N_14840,N_14743,N_14685);
nor U14841 (N_14841,N_14516,N_14735);
xnor U14842 (N_14842,N_14579,N_14547);
and U14843 (N_14843,N_14623,N_14718);
xnor U14844 (N_14844,N_14628,N_14723);
nor U14845 (N_14845,N_14543,N_14622);
nand U14846 (N_14846,N_14629,N_14560);
xor U14847 (N_14847,N_14605,N_14734);
xnor U14848 (N_14848,N_14715,N_14575);
and U14849 (N_14849,N_14598,N_14580);
xnor U14850 (N_14850,N_14599,N_14716);
or U14851 (N_14851,N_14554,N_14578);
and U14852 (N_14852,N_14540,N_14564);
nor U14853 (N_14853,N_14551,N_14711);
and U14854 (N_14854,N_14691,N_14645);
nand U14855 (N_14855,N_14600,N_14601);
or U14856 (N_14856,N_14632,N_14695);
or U14857 (N_14857,N_14667,N_14745);
nor U14858 (N_14858,N_14684,N_14544);
xor U14859 (N_14859,N_14692,N_14663);
or U14860 (N_14860,N_14634,N_14611);
nand U14861 (N_14861,N_14503,N_14631);
nor U14862 (N_14862,N_14581,N_14512);
and U14863 (N_14863,N_14615,N_14583);
nand U14864 (N_14864,N_14593,N_14558);
or U14865 (N_14865,N_14620,N_14668);
nor U14866 (N_14866,N_14511,N_14561);
or U14867 (N_14867,N_14639,N_14553);
and U14868 (N_14868,N_14686,N_14703);
nor U14869 (N_14869,N_14587,N_14585);
and U14870 (N_14870,N_14529,N_14694);
or U14871 (N_14871,N_14517,N_14609);
xnor U14872 (N_14872,N_14725,N_14505);
xnor U14873 (N_14873,N_14508,N_14510);
nor U14874 (N_14874,N_14546,N_14647);
xor U14875 (N_14875,N_14520,N_14651);
xor U14876 (N_14876,N_14507,N_14702);
xor U14877 (N_14877,N_14510,N_14589);
or U14878 (N_14878,N_14591,N_14583);
nand U14879 (N_14879,N_14735,N_14691);
nand U14880 (N_14880,N_14518,N_14687);
nor U14881 (N_14881,N_14535,N_14677);
nor U14882 (N_14882,N_14587,N_14739);
or U14883 (N_14883,N_14707,N_14580);
nor U14884 (N_14884,N_14504,N_14651);
nand U14885 (N_14885,N_14608,N_14665);
nand U14886 (N_14886,N_14585,N_14590);
nand U14887 (N_14887,N_14710,N_14711);
xnor U14888 (N_14888,N_14577,N_14500);
or U14889 (N_14889,N_14687,N_14556);
xor U14890 (N_14890,N_14689,N_14710);
nor U14891 (N_14891,N_14642,N_14500);
nor U14892 (N_14892,N_14620,N_14565);
nor U14893 (N_14893,N_14668,N_14533);
nor U14894 (N_14894,N_14592,N_14702);
and U14895 (N_14895,N_14570,N_14704);
nor U14896 (N_14896,N_14515,N_14625);
nor U14897 (N_14897,N_14722,N_14514);
xor U14898 (N_14898,N_14579,N_14552);
nand U14899 (N_14899,N_14666,N_14698);
and U14900 (N_14900,N_14728,N_14571);
nand U14901 (N_14901,N_14694,N_14567);
nor U14902 (N_14902,N_14695,N_14561);
nor U14903 (N_14903,N_14622,N_14693);
and U14904 (N_14904,N_14696,N_14501);
nand U14905 (N_14905,N_14565,N_14733);
and U14906 (N_14906,N_14670,N_14501);
or U14907 (N_14907,N_14528,N_14630);
nor U14908 (N_14908,N_14538,N_14559);
and U14909 (N_14909,N_14547,N_14571);
or U14910 (N_14910,N_14710,N_14523);
and U14911 (N_14911,N_14740,N_14697);
nor U14912 (N_14912,N_14603,N_14722);
and U14913 (N_14913,N_14659,N_14596);
xnor U14914 (N_14914,N_14616,N_14626);
or U14915 (N_14915,N_14679,N_14688);
nand U14916 (N_14916,N_14558,N_14710);
nor U14917 (N_14917,N_14700,N_14542);
nor U14918 (N_14918,N_14519,N_14636);
and U14919 (N_14919,N_14534,N_14528);
nor U14920 (N_14920,N_14662,N_14514);
nand U14921 (N_14921,N_14706,N_14530);
or U14922 (N_14922,N_14557,N_14700);
nand U14923 (N_14923,N_14508,N_14573);
and U14924 (N_14924,N_14507,N_14667);
nor U14925 (N_14925,N_14717,N_14577);
nand U14926 (N_14926,N_14500,N_14734);
xor U14927 (N_14927,N_14628,N_14560);
nand U14928 (N_14928,N_14739,N_14660);
or U14929 (N_14929,N_14675,N_14658);
and U14930 (N_14930,N_14586,N_14572);
and U14931 (N_14931,N_14568,N_14624);
nand U14932 (N_14932,N_14650,N_14708);
or U14933 (N_14933,N_14709,N_14607);
xnor U14934 (N_14934,N_14639,N_14658);
nand U14935 (N_14935,N_14669,N_14660);
nand U14936 (N_14936,N_14586,N_14549);
and U14937 (N_14937,N_14505,N_14635);
xnor U14938 (N_14938,N_14610,N_14506);
or U14939 (N_14939,N_14661,N_14716);
or U14940 (N_14940,N_14701,N_14732);
and U14941 (N_14941,N_14684,N_14600);
or U14942 (N_14942,N_14526,N_14618);
nand U14943 (N_14943,N_14665,N_14613);
and U14944 (N_14944,N_14688,N_14550);
xnor U14945 (N_14945,N_14541,N_14589);
nand U14946 (N_14946,N_14552,N_14503);
xnor U14947 (N_14947,N_14502,N_14567);
and U14948 (N_14948,N_14611,N_14594);
nor U14949 (N_14949,N_14590,N_14717);
nor U14950 (N_14950,N_14536,N_14665);
xor U14951 (N_14951,N_14706,N_14678);
nand U14952 (N_14952,N_14535,N_14582);
and U14953 (N_14953,N_14505,N_14681);
or U14954 (N_14954,N_14739,N_14503);
nand U14955 (N_14955,N_14691,N_14506);
or U14956 (N_14956,N_14665,N_14634);
or U14957 (N_14957,N_14732,N_14594);
nand U14958 (N_14958,N_14638,N_14684);
and U14959 (N_14959,N_14579,N_14524);
or U14960 (N_14960,N_14743,N_14674);
xnor U14961 (N_14961,N_14667,N_14516);
xnor U14962 (N_14962,N_14647,N_14601);
nor U14963 (N_14963,N_14705,N_14737);
nor U14964 (N_14964,N_14523,N_14705);
nand U14965 (N_14965,N_14544,N_14717);
xnor U14966 (N_14966,N_14678,N_14587);
or U14967 (N_14967,N_14580,N_14569);
nor U14968 (N_14968,N_14528,N_14722);
xor U14969 (N_14969,N_14574,N_14686);
nand U14970 (N_14970,N_14731,N_14614);
xor U14971 (N_14971,N_14666,N_14622);
xor U14972 (N_14972,N_14584,N_14579);
nand U14973 (N_14973,N_14653,N_14665);
nand U14974 (N_14974,N_14600,N_14580);
nor U14975 (N_14975,N_14564,N_14500);
nand U14976 (N_14976,N_14680,N_14501);
and U14977 (N_14977,N_14582,N_14590);
nand U14978 (N_14978,N_14694,N_14691);
xnor U14979 (N_14979,N_14510,N_14590);
nor U14980 (N_14980,N_14687,N_14580);
nand U14981 (N_14981,N_14744,N_14652);
xor U14982 (N_14982,N_14514,N_14560);
nor U14983 (N_14983,N_14561,N_14562);
nand U14984 (N_14984,N_14680,N_14639);
and U14985 (N_14985,N_14720,N_14658);
or U14986 (N_14986,N_14598,N_14720);
or U14987 (N_14987,N_14576,N_14593);
nand U14988 (N_14988,N_14698,N_14530);
and U14989 (N_14989,N_14614,N_14747);
xor U14990 (N_14990,N_14675,N_14525);
nand U14991 (N_14991,N_14717,N_14673);
xor U14992 (N_14992,N_14647,N_14748);
nor U14993 (N_14993,N_14723,N_14547);
nand U14994 (N_14994,N_14519,N_14552);
nor U14995 (N_14995,N_14698,N_14652);
xnor U14996 (N_14996,N_14556,N_14664);
and U14997 (N_14997,N_14515,N_14604);
or U14998 (N_14998,N_14667,N_14683);
nor U14999 (N_14999,N_14501,N_14593);
xnor UO_0 (O_0,N_14793,N_14848);
xor UO_1 (O_1,N_14830,N_14949);
nor UO_2 (O_2,N_14814,N_14854);
nand UO_3 (O_3,N_14826,N_14787);
and UO_4 (O_4,N_14803,N_14795);
or UO_5 (O_5,N_14886,N_14956);
xnor UO_6 (O_6,N_14918,N_14768);
or UO_7 (O_7,N_14978,N_14895);
and UO_8 (O_8,N_14836,N_14766);
nor UO_9 (O_9,N_14917,N_14801);
nor UO_10 (O_10,N_14948,N_14792);
nor UO_11 (O_11,N_14817,N_14852);
or UO_12 (O_12,N_14868,N_14984);
xor UO_13 (O_13,N_14955,N_14977);
xor UO_14 (O_14,N_14820,N_14783);
or UO_15 (O_15,N_14763,N_14858);
xor UO_16 (O_16,N_14941,N_14937);
nand UO_17 (O_17,N_14780,N_14804);
nand UO_18 (O_18,N_14876,N_14981);
and UO_19 (O_19,N_14930,N_14775);
and UO_20 (O_20,N_14965,N_14844);
nand UO_21 (O_21,N_14771,N_14944);
xor UO_22 (O_22,N_14811,N_14791);
nor UO_23 (O_23,N_14901,N_14878);
or UO_24 (O_24,N_14913,N_14750);
nand UO_25 (O_25,N_14823,N_14983);
nor UO_26 (O_26,N_14778,N_14967);
nor UO_27 (O_27,N_14921,N_14943);
xor UO_28 (O_28,N_14985,N_14888);
xor UO_29 (O_29,N_14924,N_14890);
nor UO_30 (O_30,N_14782,N_14831);
and UO_31 (O_31,N_14935,N_14964);
nor UO_32 (O_32,N_14767,N_14860);
and UO_33 (O_33,N_14870,N_14970);
or UO_34 (O_34,N_14899,N_14845);
or UO_35 (O_35,N_14821,N_14797);
nand UO_36 (O_36,N_14798,N_14954);
or UO_37 (O_37,N_14754,N_14835);
xnor UO_38 (O_38,N_14927,N_14802);
xnor UO_39 (O_39,N_14769,N_14786);
xnor UO_40 (O_40,N_14796,N_14806);
xnor UO_41 (O_41,N_14968,N_14887);
nor UO_42 (O_42,N_14907,N_14963);
or UO_43 (O_43,N_14946,N_14897);
or UO_44 (O_44,N_14997,N_14859);
nand UO_45 (O_45,N_14986,N_14815);
and UO_46 (O_46,N_14822,N_14829);
and UO_47 (O_47,N_14837,N_14961);
nand UO_48 (O_48,N_14816,N_14932);
and UO_49 (O_49,N_14863,N_14862);
and UO_50 (O_50,N_14973,N_14996);
xnor UO_51 (O_51,N_14923,N_14936);
or UO_52 (O_52,N_14819,N_14869);
nand UO_53 (O_53,N_14951,N_14885);
and UO_54 (O_54,N_14893,N_14753);
nor UO_55 (O_55,N_14812,N_14942);
xor UO_56 (O_56,N_14762,N_14914);
and UO_57 (O_57,N_14827,N_14759);
xor UO_58 (O_58,N_14898,N_14853);
nand UO_59 (O_59,N_14980,N_14889);
xor UO_60 (O_60,N_14999,N_14912);
nor UO_61 (O_61,N_14777,N_14785);
and UO_62 (O_62,N_14872,N_14883);
nand UO_63 (O_63,N_14765,N_14903);
nand UO_64 (O_64,N_14906,N_14789);
and UO_65 (O_65,N_14784,N_14857);
and UO_66 (O_66,N_14843,N_14866);
xor UO_67 (O_67,N_14894,N_14969);
or UO_68 (O_68,N_14755,N_14904);
nand UO_69 (O_69,N_14781,N_14877);
and UO_70 (O_70,N_14947,N_14865);
and UO_71 (O_71,N_14756,N_14884);
nor UO_72 (O_72,N_14770,N_14879);
xor UO_73 (O_73,N_14752,N_14988);
nor UO_74 (O_74,N_14991,N_14851);
or UO_75 (O_75,N_14794,N_14881);
or UO_76 (O_76,N_14842,N_14774);
nor UO_77 (O_77,N_14875,N_14995);
nor UO_78 (O_78,N_14779,N_14920);
nor UO_79 (O_79,N_14758,N_14846);
nor UO_80 (O_80,N_14925,N_14790);
nor UO_81 (O_81,N_14761,N_14849);
or UO_82 (O_82,N_14864,N_14805);
xnor UO_83 (O_83,N_14873,N_14922);
and UO_84 (O_84,N_14909,N_14976);
nor UO_85 (O_85,N_14838,N_14957);
and UO_86 (O_86,N_14840,N_14994);
nor UO_87 (O_87,N_14799,N_14861);
and UO_88 (O_88,N_14828,N_14962);
xor UO_89 (O_89,N_14807,N_14952);
xor UO_90 (O_90,N_14919,N_14833);
and UO_91 (O_91,N_14929,N_14834);
nand UO_92 (O_92,N_14867,N_14931);
nand UO_93 (O_93,N_14841,N_14800);
xor UO_94 (O_94,N_14900,N_14891);
xnor UO_95 (O_95,N_14809,N_14751);
nor UO_96 (O_96,N_14832,N_14975);
xor UO_97 (O_97,N_14908,N_14953);
and UO_98 (O_98,N_14773,N_14938);
nor UO_99 (O_99,N_14971,N_14982);
nor UO_100 (O_100,N_14998,N_14989);
nand UO_101 (O_101,N_14966,N_14772);
and UO_102 (O_102,N_14990,N_14915);
nand UO_103 (O_103,N_14939,N_14979);
xnor UO_104 (O_104,N_14850,N_14950);
xnor UO_105 (O_105,N_14825,N_14757);
and UO_106 (O_106,N_14776,N_14910);
xnor UO_107 (O_107,N_14839,N_14874);
nor UO_108 (O_108,N_14824,N_14959);
nor UO_109 (O_109,N_14960,N_14880);
xor UO_110 (O_110,N_14788,N_14760);
or UO_111 (O_111,N_14856,N_14871);
xnor UO_112 (O_112,N_14958,N_14896);
nor UO_113 (O_113,N_14987,N_14916);
and UO_114 (O_114,N_14764,N_14905);
and UO_115 (O_115,N_14902,N_14892);
xnor UO_116 (O_116,N_14855,N_14810);
and UO_117 (O_117,N_14882,N_14813);
or UO_118 (O_118,N_14926,N_14847);
and UO_119 (O_119,N_14818,N_14945);
and UO_120 (O_120,N_14940,N_14808);
or UO_121 (O_121,N_14972,N_14992);
nor UO_122 (O_122,N_14934,N_14933);
or UO_123 (O_123,N_14928,N_14974);
xor UO_124 (O_124,N_14993,N_14911);
xnor UO_125 (O_125,N_14838,N_14814);
xor UO_126 (O_126,N_14876,N_14832);
and UO_127 (O_127,N_14960,N_14867);
or UO_128 (O_128,N_14984,N_14902);
nand UO_129 (O_129,N_14781,N_14951);
and UO_130 (O_130,N_14783,N_14947);
and UO_131 (O_131,N_14903,N_14761);
nor UO_132 (O_132,N_14940,N_14998);
nor UO_133 (O_133,N_14861,N_14915);
or UO_134 (O_134,N_14887,N_14980);
and UO_135 (O_135,N_14787,N_14964);
xor UO_136 (O_136,N_14783,N_14846);
nor UO_137 (O_137,N_14979,N_14955);
nand UO_138 (O_138,N_14985,N_14987);
or UO_139 (O_139,N_14967,N_14790);
nor UO_140 (O_140,N_14784,N_14878);
or UO_141 (O_141,N_14873,N_14809);
and UO_142 (O_142,N_14814,N_14903);
xnor UO_143 (O_143,N_14856,N_14986);
nor UO_144 (O_144,N_14913,N_14914);
nand UO_145 (O_145,N_14834,N_14823);
and UO_146 (O_146,N_14911,N_14753);
and UO_147 (O_147,N_14896,N_14979);
or UO_148 (O_148,N_14762,N_14810);
and UO_149 (O_149,N_14865,N_14915);
or UO_150 (O_150,N_14961,N_14754);
nor UO_151 (O_151,N_14922,N_14760);
nand UO_152 (O_152,N_14990,N_14783);
nor UO_153 (O_153,N_14977,N_14960);
nand UO_154 (O_154,N_14920,N_14915);
or UO_155 (O_155,N_14784,N_14902);
and UO_156 (O_156,N_14831,N_14792);
nor UO_157 (O_157,N_14757,N_14794);
nor UO_158 (O_158,N_14768,N_14854);
or UO_159 (O_159,N_14786,N_14904);
xnor UO_160 (O_160,N_14852,N_14993);
or UO_161 (O_161,N_14804,N_14823);
nor UO_162 (O_162,N_14868,N_14894);
nor UO_163 (O_163,N_14996,N_14966);
xor UO_164 (O_164,N_14920,N_14857);
nor UO_165 (O_165,N_14981,N_14825);
nand UO_166 (O_166,N_14928,N_14948);
nand UO_167 (O_167,N_14921,N_14808);
nand UO_168 (O_168,N_14899,N_14881);
nand UO_169 (O_169,N_14963,N_14820);
nor UO_170 (O_170,N_14892,N_14765);
nor UO_171 (O_171,N_14861,N_14966);
xnor UO_172 (O_172,N_14809,N_14888);
or UO_173 (O_173,N_14761,N_14887);
or UO_174 (O_174,N_14980,N_14862);
nor UO_175 (O_175,N_14756,N_14936);
nand UO_176 (O_176,N_14957,N_14936);
or UO_177 (O_177,N_14793,N_14821);
nor UO_178 (O_178,N_14940,N_14987);
and UO_179 (O_179,N_14907,N_14948);
and UO_180 (O_180,N_14778,N_14849);
nor UO_181 (O_181,N_14799,N_14800);
xor UO_182 (O_182,N_14766,N_14955);
xnor UO_183 (O_183,N_14878,N_14929);
and UO_184 (O_184,N_14755,N_14786);
nand UO_185 (O_185,N_14944,N_14790);
xnor UO_186 (O_186,N_14765,N_14913);
nor UO_187 (O_187,N_14850,N_14843);
or UO_188 (O_188,N_14835,N_14872);
nand UO_189 (O_189,N_14857,N_14823);
nor UO_190 (O_190,N_14852,N_14899);
nand UO_191 (O_191,N_14942,N_14843);
nand UO_192 (O_192,N_14889,N_14896);
xnor UO_193 (O_193,N_14780,N_14932);
or UO_194 (O_194,N_14981,N_14997);
xor UO_195 (O_195,N_14866,N_14902);
nand UO_196 (O_196,N_14849,N_14979);
and UO_197 (O_197,N_14914,N_14880);
xnor UO_198 (O_198,N_14897,N_14754);
nor UO_199 (O_199,N_14973,N_14914);
nor UO_200 (O_200,N_14799,N_14896);
nor UO_201 (O_201,N_14939,N_14857);
xnor UO_202 (O_202,N_14975,N_14754);
nand UO_203 (O_203,N_14863,N_14796);
xor UO_204 (O_204,N_14843,N_14903);
or UO_205 (O_205,N_14837,N_14950);
xor UO_206 (O_206,N_14830,N_14984);
nor UO_207 (O_207,N_14848,N_14755);
or UO_208 (O_208,N_14888,N_14873);
nor UO_209 (O_209,N_14897,N_14883);
nor UO_210 (O_210,N_14836,N_14904);
and UO_211 (O_211,N_14913,N_14897);
nand UO_212 (O_212,N_14856,N_14755);
xor UO_213 (O_213,N_14786,N_14963);
or UO_214 (O_214,N_14761,N_14785);
nor UO_215 (O_215,N_14767,N_14959);
or UO_216 (O_216,N_14997,N_14791);
and UO_217 (O_217,N_14754,N_14852);
or UO_218 (O_218,N_14843,N_14853);
or UO_219 (O_219,N_14812,N_14782);
nand UO_220 (O_220,N_14815,N_14855);
or UO_221 (O_221,N_14918,N_14826);
nand UO_222 (O_222,N_14970,N_14822);
or UO_223 (O_223,N_14771,N_14827);
or UO_224 (O_224,N_14788,N_14798);
nand UO_225 (O_225,N_14752,N_14919);
nand UO_226 (O_226,N_14859,N_14926);
nand UO_227 (O_227,N_14943,N_14754);
nor UO_228 (O_228,N_14750,N_14814);
or UO_229 (O_229,N_14810,N_14808);
nand UO_230 (O_230,N_14951,N_14876);
and UO_231 (O_231,N_14948,N_14786);
nand UO_232 (O_232,N_14798,N_14933);
nor UO_233 (O_233,N_14920,N_14755);
or UO_234 (O_234,N_14811,N_14775);
or UO_235 (O_235,N_14840,N_14896);
and UO_236 (O_236,N_14896,N_14931);
nor UO_237 (O_237,N_14918,N_14803);
nor UO_238 (O_238,N_14897,N_14925);
nor UO_239 (O_239,N_14758,N_14784);
or UO_240 (O_240,N_14978,N_14826);
nand UO_241 (O_241,N_14964,N_14868);
nand UO_242 (O_242,N_14914,N_14831);
xnor UO_243 (O_243,N_14757,N_14898);
or UO_244 (O_244,N_14869,N_14919);
and UO_245 (O_245,N_14819,N_14829);
nor UO_246 (O_246,N_14750,N_14915);
and UO_247 (O_247,N_14980,N_14947);
nand UO_248 (O_248,N_14819,N_14913);
xor UO_249 (O_249,N_14888,N_14829);
or UO_250 (O_250,N_14807,N_14987);
or UO_251 (O_251,N_14893,N_14807);
nand UO_252 (O_252,N_14983,N_14993);
or UO_253 (O_253,N_14932,N_14853);
nor UO_254 (O_254,N_14868,N_14885);
and UO_255 (O_255,N_14780,N_14867);
and UO_256 (O_256,N_14752,N_14887);
nand UO_257 (O_257,N_14911,N_14803);
and UO_258 (O_258,N_14834,N_14977);
xnor UO_259 (O_259,N_14961,N_14859);
nand UO_260 (O_260,N_14917,N_14988);
or UO_261 (O_261,N_14870,N_14862);
nand UO_262 (O_262,N_14993,N_14782);
or UO_263 (O_263,N_14953,N_14779);
xor UO_264 (O_264,N_14894,N_14783);
xnor UO_265 (O_265,N_14823,N_14788);
nor UO_266 (O_266,N_14876,N_14980);
xnor UO_267 (O_267,N_14859,N_14970);
and UO_268 (O_268,N_14874,N_14913);
nand UO_269 (O_269,N_14985,N_14950);
and UO_270 (O_270,N_14852,N_14834);
nor UO_271 (O_271,N_14907,N_14836);
xor UO_272 (O_272,N_14786,N_14875);
or UO_273 (O_273,N_14853,N_14863);
xor UO_274 (O_274,N_14900,N_14852);
and UO_275 (O_275,N_14898,N_14759);
nand UO_276 (O_276,N_14838,N_14850);
or UO_277 (O_277,N_14780,N_14762);
nand UO_278 (O_278,N_14938,N_14852);
or UO_279 (O_279,N_14977,N_14813);
xor UO_280 (O_280,N_14934,N_14811);
and UO_281 (O_281,N_14807,N_14813);
and UO_282 (O_282,N_14933,N_14812);
nor UO_283 (O_283,N_14927,N_14873);
nor UO_284 (O_284,N_14883,N_14972);
xor UO_285 (O_285,N_14871,N_14829);
and UO_286 (O_286,N_14812,N_14854);
xnor UO_287 (O_287,N_14918,N_14860);
or UO_288 (O_288,N_14999,N_14977);
nor UO_289 (O_289,N_14955,N_14764);
xor UO_290 (O_290,N_14972,N_14819);
and UO_291 (O_291,N_14835,N_14924);
nand UO_292 (O_292,N_14816,N_14996);
and UO_293 (O_293,N_14935,N_14868);
nand UO_294 (O_294,N_14897,N_14911);
nand UO_295 (O_295,N_14884,N_14752);
nor UO_296 (O_296,N_14985,N_14956);
or UO_297 (O_297,N_14776,N_14855);
xor UO_298 (O_298,N_14927,N_14913);
xnor UO_299 (O_299,N_14955,N_14933);
nand UO_300 (O_300,N_14955,N_14818);
and UO_301 (O_301,N_14949,N_14857);
and UO_302 (O_302,N_14772,N_14882);
xor UO_303 (O_303,N_14922,N_14753);
or UO_304 (O_304,N_14902,N_14756);
xor UO_305 (O_305,N_14871,N_14869);
xor UO_306 (O_306,N_14808,N_14928);
or UO_307 (O_307,N_14780,N_14876);
xor UO_308 (O_308,N_14768,N_14793);
or UO_309 (O_309,N_14974,N_14943);
and UO_310 (O_310,N_14897,N_14974);
and UO_311 (O_311,N_14867,N_14889);
xor UO_312 (O_312,N_14840,N_14845);
or UO_313 (O_313,N_14805,N_14824);
and UO_314 (O_314,N_14810,N_14875);
and UO_315 (O_315,N_14876,N_14978);
and UO_316 (O_316,N_14831,N_14827);
or UO_317 (O_317,N_14845,N_14989);
nor UO_318 (O_318,N_14923,N_14856);
or UO_319 (O_319,N_14871,N_14860);
or UO_320 (O_320,N_14805,N_14902);
nor UO_321 (O_321,N_14902,N_14793);
and UO_322 (O_322,N_14780,N_14837);
nor UO_323 (O_323,N_14798,N_14764);
nand UO_324 (O_324,N_14896,N_14830);
xor UO_325 (O_325,N_14901,N_14926);
or UO_326 (O_326,N_14994,N_14905);
nor UO_327 (O_327,N_14893,N_14935);
and UO_328 (O_328,N_14765,N_14904);
or UO_329 (O_329,N_14911,N_14862);
nor UO_330 (O_330,N_14877,N_14943);
and UO_331 (O_331,N_14948,N_14837);
xor UO_332 (O_332,N_14802,N_14806);
nand UO_333 (O_333,N_14780,N_14824);
nand UO_334 (O_334,N_14750,N_14838);
or UO_335 (O_335,N_14905,N_14936);
and UO_336 (O_336,N_14954,N_14935);
or UO_337 (O_337,N_14760,N_14928);
and UO_338 (O_338,N_14756,N_14876);
xnor UO_339 (O_339,N_14754,N_14829);
nor UO_340 (O_340,N_14962,N_14775);
or UO_341 (O_341,N_14845,N_14847);
nor UO_342 (O_342,N_14820,N_14906);
or UO_343 (O_343,N_14854,N_14894);
nor UO_344 (O_344,N_14870,N_14840);
nor UO_345 (O_345,N_14806,N_14919);
or UO_346 (O_346,N_14994,N_14752);
and UO_347 (O_347,N_14870,N_14883);
nor UO_348 (O_348,N_14838,N_14770);
nor UO_349 (O_349,N_14805,N_14781);
nand UO_350 (O_350,N_14757,N_14886);
or UO_351 (O_351,N_14979,N_14819);
or UO_352 (O_352,N_14782,N_14762);
nand UO_353 (O_353,N_14956,N_14955);
nor UO_354 (O_354,N_14974,N_14936);
nor UO_355 (O_355,N_14983,N_14816);
nand UO_356 (O_356,N_14764,N_14823);
xor UO_357 (O_357,N_14787,N_14784);
xor UO_358 (O_358,N_14799,N_14775);
nand UO_359 (O_359,N_14842,N_14986);
and UO_360 (O_360,N_14833,N_14798);
or UO_361 (O_361,N_14819,N_14879);
nand UO_362 (O_362,N_14849,N_14928);
xor UO_363 (O_363,N_14785,N_14844);
nand UO_364 (O_364,N_14913,N_14835);
and UO_365 (O_365,N_14750,N_14775);
or UO_366 (O_366,N_14890,N_14867);
and UO_367 (O_367,N_14847,N_14890);
nand UO_368 (O_368,N_14877,N_14999);
and UO_369 (O_369,N_14823,N_14887);
nor UO_370 (O_370,N_14982,N_14831);
nand UO_371 (O_371,N_14899,N_14875);
nand UO_372 (O_372,N_14940,N_14972);
and UO_373 (O_373,N_14997,N_14980);
xnor UO_374 (O_374,N_14778,N_14772);
and UO_375 (O_375,N_14857,N_14951);
nor UO_376 (O_376,N_14844,N_14750);
nand UO_377 (O_377,N_14838,N_14794);
or UO_378 (O_378,N_14821,N_14901);
and UO_379 (O_379,N_14894,N_14774);
nand UO_380 (O_380,N_14951,N_14839);
nand UO_381 (O_381,N_14848,N_14859);
nor UO_382 (O_382,N_14871,N_14815);
nand UO_383 (O_383,N_14834,N_14840);
nand UO_384 (O_384,N_14808,N_14862);
xnor UO_385 (O_385,N_14898,N_14784);
or UO_386 (O_386,N_14809,N_14928);
nand UO_387 (O_387,N_14928,N_14888);
and UO_388 (O_388,N_14836,N_14821);
or UO_389 (O_389,N_14958,N_14798);
or UO_390 (O_390,N_14756,N_14840);
xor UO_391 (O_391,N_14987,N_14766);
and UO_392 (O_392,N_14776,N_14757);
xnor UO_393 (O_393,N_14922,N_14823);
nor UO_394 (O_394,N_14997,N_14852);
nor UO_395 (O_395,N_14860,N_14945);
xor UO_396 (O_396,N_14885,N_14960);
or UO_397 (O_397,N_14949,N_14897);
or UO_398 (O_398,N_14843,N_14778);
xnor UO_399 (O_399,N_14879,N_14924);
nor UO_400 (O_400,N_14929,N_14846);
nor UO_401 (O_401,N_14881,N_14940);
xor UO_402 (O_402,N_14771,N_14866);
nand UO_403 (O_403,N_14897,N_14794);
and UO_404 (O_404,N_14881,N_14968);
and UO_405 (O_405,N_14841,N_14848);
or UO_406 (O_406,N_14902,N_14868);
xnor UO_407 (O_407,N_14817,N_14790);
and UO_408 (O_408,N_14901,N_14960);
and UO_409 (O_409,N_14955,N_14799);
or UO_410 (O_410,N_14818,N_14960);
xnor UO_411 (O_411,N_14784,N_14949);
nand UO_412 (O_412,N_14837,N_14929);
and UO_413 (O_413,N_14854,N_14989);
or UO_414 (O_414,N_14782,N_14878);
and UO_415 (O_415,N_14827,N_14800);
xnor UO_416 (O_416,N_14931,N_14884);
xnor UO_417 (O_417,N_14938,N_14963);
nor UO_418 (O_418,N_14973,N_14793);
and UO_419 (O_419,N_14944,N_14840);
xor UO_420 (O_420,N_14926,N_14992);
nand UO_421 (O_421,N_14794,N_14850);
xnor UO_422 (O_422,N_14759,N_14905);
and UO_423 (O_423,N_14901,N_14758);
and UO_424 (O_424,N_14993,N_14991);
and UO_425 (O_425,N_14846,N_14961);
and UO_426 (O_426,N_14958,N_14949);
and UO_427 (O_427,N_14909,N_14877);
nand UO_428 (O_428,N_14923,N_14906);
nor UO_429 (O_429,N_14905,N_14827);
xnor UO_430 (O_430,N_14772,N_14847);
nor UO_431 (O_431,N_14925,N_14901);
xnor UO_432 (O_432,N_14872,N_14772);
and UO_433 (O_433,N_14756,N_14919);
or UO_434 (O_434,N_14945,N_14891);
xnor UO_435 (O_435,N_14823,N_14967);
nor UO_436 (O_436,N_14806,N_14859);
nand UO_437 (O_437,N_14901,N_14889);
nor UO_438 (O_438,N_14826,N_14900);
and UO_439 (O_439,N_14971,N_14901);
nand UO_440 (O_440,N_14939,N_14913);
and UO_441 (O_441,N_14941,N_14770);
or UO_442 (O_442,N_14832,N_14849);
nor UO_443 (O_443,N_14984,N_14838);
and UO_444 (O_444,N_14864,N_14816);
xor UO_445 (O_445,N_14774,N_14998);
nand UO_446 (O_446,N_14767,N_14785);
and UO_447 (O_447,N_14762,N_14959);
nand UO_448 (O_448,N_14973,N_14866);
nor UO_449 (O_449,N_14801,N_14835);
nand UO_450 (O_450,N_14976,N_14768);
or UO_451 (O_451,N_14948,N_14986);
nor UO_452 (O_452,N_14899,N_14916);
nor UO_453 (O_453,N_14803,N_14822);
and UO_454 (O_454,N_14871,N_14933);
nor UO_455 (O_455,N_14767,N_14993);
nand UO_456 (O_456,N_14837,N_14849);
or UO_457 (O_457,N_14926,N_14954);
nor UO_458 (O_458,N_14772,N_14792);
nand UO_459 (O_459,N_14816,N_14802);
nor UO_460 (O_460,N_14880,N_14859);
xnor UO_461 (O_461,N_14966,N_14858);
xnor UO_462 (O_462,N_14876,N_14838);
nand UO_463 (O_463,N_14868,N_14838);
nor UO_464 (O_464,N_14916,N_14889);
or UO_465 (O_465,N_14974,N_14766);
nand UO_466 (O_466,N_14848,N_14993);
and UO_467 (O_467,N_14994,N_14965);
nand UO_468 (O_468,N_14860,N_14855);
xnor UO_469 (O_469,N_14827,N_14990);
nand UO_470 (O_470,N_14978,N_14782);
xnor UO_471 (O_471,N_14919,N_14831);
xnor UO_472 (O_472,N_14786,N_14759);
nand UO_473 (O_473,N_14938,N_14793);
nand UO_474 (O_474,N_14753,N_14984);
xor UO_475 (O_475,N_14800,N_14985);
nand UO_476 (O_476,N_14772,N_14893);
nor UO_477 (O_477,N_14758,N_14783);
nand UO_478 (O_478,N_14770,N_14809);
nor UO_479 (O_479,N_14864,N_14775);
nor UO_480 (O_480,N_14900,N_14804);
nand UO_481 (O_481,N_14807,N_14963);
and UO_482 (O_482,N_14762,N_14787);
nand UO_483 (O_483,N_14758,N_14971);
xnor UO_484 (O_484,N_14933,N_14806);
and UO_485 (O_485,N_14946,N_14843);
xnor UO_486 (O_486,N_14823,N_14795);
and UO_487 (O_487,N_14910,N_14913);
xnor UO_488 (O_488,N_14801,N_14932);
nand UO_489 (O_489,N_14847,N_14842);
and UO_490 (O_490,N_14819,N_14811);
or UO_491 (O_491,N_14769,N_14868);
xor UO_492 (O_492,N_14876,N_14884);
and UO_493 (O_493,N_14786,N_14814);
nor UO_494 (O_494,N_14771,N_14967);
nand UO_495 (O_495,N_14788,N_14881);
nor UO_496 (O_496,N_14914,N_14844);
and UO_497 (O_497,N_14774,N_14796);
nor UO_498 (O_498,N_14767,N_14947);
and UO_499 (O_499,N_14765,N_14893);
nand UO_500 (O_500,N_14963,N_14940);
or UO_501 (O_501,N_14909,N_14979);
nor UO_502 (O_502,N_14771,N_14901);
and UO_503 (O_503,N_14961,N_14769);
nand UO_504 (O_504,N_14817,N_14761);
and UO_505 (O_505,N_14791,N_14935);
nand UO_506 (O_506,N_14776,N_14917);
nor UO_507 (O_507,N_14773,N_14976);
xnor UO_508 (O_508,N_14977,N_14929);
or UO_509 (O_509,N_14819,N_14778);
nor UO_510 (O_510,N_14938,N_14826);
and UO_511 (O_511,N_14756,N_14813);
xnor UO_512 (O_512,N_14899,N_14870);
nor UO_513 (O_513,N_14942,N_14939);
xor UO_514 (O_514,N_14821,N_14953);
or UO_515 (O_515,N_14843,N_14779);
nand UO_516 (O_516,N_14858,N_14932);
nand UO_517 (O_517,N_14881,N_14822);
xnor UO_518 (O_518,N_14934,N_14836);
and UO_519 (O_519,N_14828,N_14815);
xor UO_520 (O_520,N_14881,N_14780);
nand UO_521 (O_521,N_14977,N_14907);
xor UO_522 (O_522,N_14928,N_14912);
and UO_523 (O_523,N_14970,N_14909);
nor UO_524 (O_524,N_14904,N_14801);
xor UO_525 (O_525,N_14849,N_14935);
xnor UO_526 (O_526,N_14954,N_14961);
nand UO_527 (O_527,N_14903,N_14780);
or UO_528 (O_528,N_14961,N_14755);
nor UO_529 (O_529,N_14893,N_14917);
nor UO_530 (O_530,N_14937,N_14936);
xnor UO_531 (O_531,N_14931,N_14935);
and UO_532 (O_532,N_14985,N_14946);
or UO_533 (O_533,N_14961,N_14895);
xnor UO_534 (O_534,N_14968,N_14827);
nor UO_535 (O_535,N_14952,N_14855);
or UO_536 (O_536,N_14777,N_14817);
and UO_537 (O_537,N_14940,N_14911);
nand UO_538 (O_538,N_14808,N_14837);
nand UO_539 (O_539,N_14929,N_14820);
xor UO_540 (O_540,N_14996,N_14767);
xor UO_541 (O_541,N_14816,N_14942);
nand UO_542 (O_542,N_14853,N_14948);
or UO_543 (O_543,N_14909,N_14772);
or UO_544 (O_544,N_14793,N_14874);
nor UO_545 (O_545,N_14957,N_14839);
xnor UO_546 (O_546,N_14978,N_14796);
xnor UO_547 (O_547,N_14787,N_14847);
or UO_548 (O_548,N_14819,N_14974);
nor UO_549 (O_549,N_14873,N_14994);
nor UO_550 (O_550,N_14864,N_14838);
or UO_551 (O_551,N_14789,N_14902);
xnor UO_552 (O_552,N_14885,N_14828);
nor UO_553 (O_553,N_14767,N_14916);
or UO_554 (O_554,N_14946,N_14914);
nand UO_555 (O_555,N_14932,N_14883);
xnor UO_556 (O_556,N_14901,N_14855);
nand UO_557 (O_557,N_14913,N_14877);
nor UO_558 (O_558,N_14792,N_14965);
nor UO_559 (O_559,N_14764,N_14820);
or UO_560 (O_560,N_14952,N_14980);
nor UO_561 (O_561,N_14877,N_14942);
nand UO_562 (O_562,N_14857,N_14776);
nand UO_563 (O_563,N_14862,N_14895);
and UO_564 (O_564,N_14982,N_14804);
nand UO_565 (O_565,N_14970,N_14961);
nand UO_566 (O_566,N_14802,N_14817);
nand UO_567 (O_567,N_14884,N_14862);
xor UO_568 (O_568,N_14951,N_14804);
xor UO_569 (O_569,N_14919,N_14876);
nor UO_570 (O_570,N_14988,N_14841);
xnor UO_571 (O_571,N_14798,N_14872);
nor UO_572 (O_572,N_14949,N_14890);
nand UO_573 (O_573,N_14803,N_14785);
nand UO_574 (O_574,N_14926,N_14771);
or UO_575 (O_575,N_14789,N_14846);
xnor UO_576 (O_576,N_14832,N_14961);
and UO_577 (O_577,N_14906,N_14753);
nor UO_578 (O_578,N_14981,N_14964);
and UO_579 (O_579,N_14990,N_14841);
nor UO_580 (O_580,N_14799,N_14753);
and UO_581 (O_581,N_14826,N_14991);
xor UO_582 (O_582,N_14764,N_14804);
xor UO_583 (O_583,N_14930,N_14968);
or UO_584 (O_584,N_14872,N_14930);
xor UO_585 (O_585,N_14901,N_14853);
nor UO_586 (O_586,N_14979,N_14897);
nor UO_587 (O_587,N_14899,N_14891);
xnor UO_588 (O_588,N_14859,N_14972);
and UO_589 (O_589,N_14820,N_14926);
nand UO_590 (O_590,N_14801,N_14982);
xor UO_591 (O_591,N_14831,N_14833);
or UO_592 (O_592,N_14797,N_14933);
or UO_593 (O_593,N_14827,N_14958);
or UO_594 (O_594,N_14984,N_14944);
nand UO_595 (O_595,N_14850,N_14909);
xor UO_596 (O_596,N_14781,N_14785);
nand UO_597 (O_597,N_14841,N_14820);
xor UO_598 (O_598,N_14957,N_14987);
and UO_599 (O_599,N_14971,N_14883);
or UO_600 (O_600,N_14894,N_14770);
nor UO_601 (O_601,N_14924,N_14947);
and UO_602 (O_602,N_14794,N_14916);
nand UO_603 (O_603,N_14756,N_14754);
nor UO_604 (O_604,N_14927,N_14761);
nand UO_605 (O_605,N_14852,N_14847);
and UO_606 (O_606,N_14965,N_14845);
nor UO_607 (O_607,N_14978,N_14847);
nor UO_608 (O_608,N_14978,N_14911);
nor UO_609 (O_609,N_14999,N_14913);
nor UO_610 (O_610,N_14853,N_14791);
nor UO_611 (O_611,N_14783,N_14952);
nor UO_612 (O_612,N_14829,N_14913);
or UO_613 (O_613,N_14967,N_14905);
nand UO_614 (O_614,N_14909,N_14930);
or UO_615 (O_615,N_14784,N_14854);
xnor UO_616 (O_616,N_14769,N_14917);
and UO_617 (O_617,N_14955,N_14992);
nor UO_618 (O_618,N_14830,N_14857);
xor UO_619 (O_619,N_14929,N_14779);
nor UO_620 (O_620,N_14969,N_14917);
nor UO_621 (O_621,N_14816,N_14926);
xor UO_622 (O_622,N_14990,N_14895);
xor UO_623 (O_623,N_14776,N_14779);
or UO_624 (O_624,N_14765,N_14837);
nor UO_625 (O_625,N_14838,N_14849);
xor UO_626 (O_626,N_14904,N_14879);
and UO_627 (O_627,N_14845,N_14887);
and UO_628 (O_628,N_14916,N_14820);
or UO_629 (O_629,N_14828,N_14912);
and UO_630 (O_630,N_14808,N_14986);
xor UO_631 (O_631,N_14901,N_14804);
and UO_632 (O_632,N_14797,N_14886);
or UO_633 (O_633,N_14840,N_14885);
or UO_634 (O_634,N_14830,N_14871);
nand UO_635 (O_635,N_14782,N_14825);
xor UO_636 (O_636,N_14757,N_14889);
and UO_637 (O_637,N_14755,N_14923);
or UO_638 (O_638,N_14972,N_14867);
nand UO_639 (O_639,N_14885,N_14802);
nand UO_640 (O_640,N_14779,N_14931);
nor UO_641 (O_641,N_14758,N_14923);
nand UO_642 (O_642,N_14780,N_14869);
nor UO_643 (O_643,N_14821,N_14885);
nor UO_644 (O_644,N_14826,N_14793);
nor UO_645 (O_645,N_14974,N_14864);
or UO_646 (O_646,N_14819,N_14878);
xnor UO_647 (O_647,N_14986,N_14972);
nand UO_648 (O_648,N_14990,N_14959);
and UO_649 (O_649,N_14839,N_14831);
and UO_650 (O_650,N_14750,N_14773);
and UO_651 (O_651,N_14922,N_14757);
nand UO_652 (O_652,N_14946,N_14953);
nand UO_653 (O_653,N_14983,N_14830);
or UO_654 (O_654,N_14942,N_14844);
or UO_655 (O_655,N_14962,N_14798);
or UO_656 (O_656,N_14977,N_14823);
or UO_657 (O_657,N_14917,N_14867);
or UO_658 (O_658,N_14896,N_14793);
nand UO_659 (O_659,N_14791,N_14855);
xor UO_660 (O_660,N_14765,N_14786);
xor UO_661 (O_661,N_14898,N_14955);
and UO_662 (O_662,N_14857,N_14865);
nor UO_663 (O_663,N_14781,N_14998);
and UO_664 (O_664,N_14874,N_14877);
xor UO_665 (O_665,N_14855,N_14891);
nor UO_666 (O_666,N_14890,N_14879);
or UO_667 (O_667,N_14878,N_14809);
or UO_668 (O_668,N_14908,N_14967);
nor UO_669 (O_669,N_14957,N_14974);
xnor UO_670 (O_670,N_14956,N_14868);
nand UO_671 (O_671,N_14785,N_14980);
xor UO_672 (O_672,N_14904,N_14906);
nor UO_673 (O_673,N_14890,N_14755);
or UO_674 (O_674,N_14924,N_14762);
or UO_675 (O_675,N_14916,N_14915);
nor UO_676 (O_676,N_14860,N_14977);
nor UO_677 (O_677,N_14782,N_14961);
xnor UO_678 (O_678,N_14800,N_14977);
nand UO_679 (O_679,N_14796,N_14800);
or UO_680 (O_680,N_14866,N_14854);
nand UO_681 (O_681,N_14886,N_14904);
and UO_682 (O_682,N_14913,N_14810);
nor UO_683 (O_683,N_14851,N_14937);
and UO_684 (O_684,N_14928,N_14851);
and UO_685 (O_685,N_14949,N_14871);
nand UO_686 (O_686,N_14802,N_14760);
nor UO_687 (O_687,N_14876,N_14750);
nor UO_688 (O_688,N_14999,N_14854);
nand UO_689 (O_689,N_14896,N_14888);
or UO_690 (O_690,N_14931,N_14871);
nor UO_691 (O_691,N_14879,N_14920);
nand UO_692 (O_692,N_14871,N_14813);
xor UO_693 (O_693,N_14771,N_14766);
nor UO_694 (O_694,N_14798,N_14864);
nand UO_695 (O_695,N_14781,N_14811);
or UO_696 (O_696,N_14990,N_14786);
and UO_697 (O_697,N_14871,N_14837);
xnor UO_698 (O_698,N_14971,N_14911);
and UO_699 (O_699,N_14873,N_14889);
or UO_700 (O_700,N_14996,N_14881);
and UO_701 (O_701,N_14810,N_14884);
or UO_702 (O_702,N_14983,N_14836);
xnor UO_703 (O_703,N_14890,N_14881);
xnor UO_704 (O_704,N_14900,N_14950);
xor UO_705 (O_705,N_14874,N_14778);
and UO_706 (O_706,N_14978,N_14910);
nand UO_707 (O_707,N_14865,N_14808);
nor UO_708 (O_708,N_14877,N_14776);
and UO_709 (O_709,N_14859,N_14895);
nand UO_710 (O_710,N_14989,N_14786);
and UO_711 (O_711,N_14980,N_14849);
nor UO_712 (O_712,N_14909,N_14974);
nor UO_713 (O_713,N_14795,N_14769);
nand UO_714 (O_714,N_14952,N_14771);
nand UO_715 (O_715,N_14961,N_14858);
nor UO_716 (O_716,N_14822,N_14775);
nand UO_717 (O_717,N_14785,N_14784);
or UO_718 (O_718,N_14754,N_14939);
nor UO_719 (O_719,N_14782,N_14946);
nor UO_720 (O_720,N_14888,N_14810);
nand UO_721 (O_721,N_14977,N_14973);
nor UO_722 (O_722,N_14985,N_14772);
and UO_723 (O_723,N_14912,N_14960);
nor UO_724 (O_724,N_14773,N_14913);
or UO_725 (O_725,N_14923,N_14882);
xor UO_726 (O_726,N_14881,N_14768);
nand UO_727 (O_727,N_14783,N_14797);
xnor UO_728 (O_728,N_14900,N_14979);
xor UO_729 (O_729,N_14968,N_14855);
and UO_730 (O_730,N_14890,N_14975);
nand UO_731 (O_731,N_14834,N_14854);
nor UO_732 (O_732,N_14778,N_14780);
nand UO_733 (O_733,N_14951,N_14909);
xnor UO_734 (O_734,N_14799,N_14971);
and UO_735 (O_735,N_14894,N_14769);
nor UO_736 (O_736,N_14967,N_14825);
and UO_737 (O_737,N_14863,N_14871);
or UO_738 (O_738,N_14828,N_14855);
nand UO_739 (O_739,N_14763,N_14918);
and UO_740 (O_740,N_14985,N_14785);
nor UO_741 (O_741,N_14856,N_14905);
nor UO_742 (O_742,N_14761,N_14987);
or UO_743 (O_743,N_14949,N_14826);
nand UO_744 (O_744,N_14822,N_14810);
or UO_745 (O_745,N_14965,N_14846);
nand UO_746 (O_746,N_14861,N_14910);
nand UO_747 (O_747,N_14767,N_14986);
and UO_748 (O_748,N_14884,N_14815);
or UO_749 (O_749,N_14892,N_14932);
nand UO_750 (O_750,N_14856,N_14922);
or UO_751 (O_751,N_14807,N_14808);
nand UO_752 (O_752,N_14780,N_14801);
nor UO_753 (O_753,N_14850,N_14888);
xor UO_754 (O_754,N_14880,N_14988);
nand UO_755 (O_755,N_14757,N_14766);
nand UO_756 (O_756,N_14987,N_14907);
nor UO_757 (O_757,N_14946,N_14768);
and UO_758 (O_758,N_14912,N_14934);
or UO_759 (O_759,N_14880,N_14978);
nand UO_760 (O_760,N_14836,N_14751);
nor UO_761 (O_761,N_14900,N_14751);
or UO_762 (O_762,N_14987,N_14950);
and UO_763 (O_763,N_14859,N_14782);
nand UO_764 (O_764,N_14794,N_14966);
xor UO_765 (O_765,N_14950,N_14929);
nor UO_766 (O_766,N_14925,N_14860);
and UO_767 (O_767,N_14926,N_14762);
xor UO_768 (O_768,N_14773,N_14836);
nor UO_769 (O_769,N_14920,N_14847);
or UO_770 (O_770,N_14795,N_14979);
and UO_771 (O_771,N_14914,N_14883);
and UO_772 (O_772,N_14825,N_14940);
nor UO_773 (O_773,N_14854,N_14828);
or UO_774 (O_774,N_14962,N_14778);
nor UO_775 (O_775,N_14877,N_14810);
nand UO_776 (O_776,N_14901,N_14847);
or UO_777 (O_777,N_14841,N_14897);
xnor UO_778 (O_778,N_14886,N_14781);
nor UO_779 (O_779,N_14984,N_14872);
or UO_780 (O_780,N_14889,N_14917);
and UO_781 (O_781,N_14884,N_14994);
xnor UO_782 (O_782,N_14899,N_14871);
and UO_783 (O_783,N_14802,N_14952);
and UO_784 (O_784,N_14857,N_14872);
nand UO_785 (O_785,N_14838,N_14844);
nor UO_786 (O_786,N_14913,N_14826);
nand UO_787 (O_787,N_14820,N_14895);
nand UO_788 (O_788,N_14985,N_14902);
and UO_789 (O_789,N_14786,N_14850);
nand UO_790 (O_790,N_14983,N_14881);
and UO_791 (O_791,N_14996,N_14935);
and UO_792 (O_792,N_14910,N_14827);
or UO_793 (O_793,N_14859,N_14897);
and UO_794 (O_794,N_14943,N_14806);
xnor UO_795 (O_795,N_14976,N_14831);
xnor UO_796 (O_796,N_14928,N_14905);
xor UO_797 (O_797,N_14856,N_14907);
nor UO_798 (O_798,N_14888,N_14886);
nand UO_799 (O_799,N_14779,N_14752);
nand UO_800 (O_800,N_14884,N_14985);
xor UO_801 (O_801,N_14832,N_14865);
nor UO_802 (O_802,N_14960,N_14994);
nand UO_803 (O_803,N_14958,N_14766);
nand UO_804 (O_804,N_14985,N_14780);
nor UO_805 (O_805,N_14865,N_14957);
xor UO_806 (O_806,N_14823,N_14962);
or UO_807 (O_807,N_14827,N_14776);
nand UO_808 (O_808,N_14838,N_14966);
nor UO_809 (O_809,N_14759,N_14791);
nor UO_810 (O_810,N_14918,N_14751);
and UO_811 (O_811,N_14995,N_14931);
nor UO_812 (O_812,N_14888,N_14902);
and UO_813 (O_813,N_14780,N_14842);
or UO_814 (O_814,N_14865,N_14846);
nand UO_815 (O_815,N_14945,N_14815);
or UO_816 (O_816,N_14897,N_14916);
xor UO_817 (O_817,N_14776,N_14894);
nor UO_818 (O_818,N_14971,N_14940);
xnor UO_819 (O_819,N_14985,N_14750);
nand UO_820 (O_820,N_14930,N_14829);
and UO_821 (O_821,N_14974,N_14870);
or UO_822 (O_822,N_14849,N_14963);
xor UO_823 (O_823,N_14931,N_14899);
nor UO_824 (O_824,N_14844,N_14908);
nand UO_825 (O_825,N_14787,N_14862);
nand UO_826 (O_826,N_14797,N_14950);
or UO_827 (O_827,N_14782,N_14811);
or UO_828 (O_828,N_14776,N_14772);
xnor UO_829 (O_829,N_14768,N_14987);
or UO_830 (O_830,N_14891,N_14812);
or UO_831 (O_831,N_14829,N_14780);
xnor UO_832 (O_832,N_14951,N_14814);
nand UO_833 (O_833,N_14977,N_14810);
or UO_834 (O_834,N_14917,N_14794);
or UO_835 (O_835,N_14972,N_14851);
nor UO_836 (O_836,N_14980,N_14912);
or UO_837 (O_837,N_14780,N_14800);
xnor UO_838 (O_838,N_14768,N_14831);
or UO_839 (O_839,N_14946,N_14956);
or UO_840 (O_840,N_14985,N_14978);
and UO_841 (O_841,N_14942,N_14904);
nand UO_842 (O_842,N_14828,N_14904);
xnor UO_843 (O_843,N_14968,N_14987);
nand UO_844 (O_844,N_14920,N_14767);
nand UO_845 (O_845,N_14871,N_14785);
and UO_846 (O_846,N_14877,N_14840);
or UO_847 (O_847,N_14986,N_14981);
or UO_848 (O_848,N_14792,N_14879);
xnor UO_849 (O_849,N_14964,N_14793);
nand UO_850 (O_850,N_14986,N_14890);
or UO_851 (O_851,N_14929,N_14751);
nor UO_852 (O_852,N_14856,N_14769);
nand UO_853 (O_853,N_14786,N_14775);
nand UO_854 (O_854,N_14855,N_14797);
and UO_855 (O_855,N_14870,N_14964);
and UO_856 (O_856,N_14852,N_14751);
nand UO_857 (O_857,N_14996,N_14808);
nor UO_858 (O_858,N_14849,N_14788);
and UO_859 (O_859,N_14865,N_14814);
nand UO_860 (O_860,N_14821,N_14878);
or UO_861 (O_861,N_14780,N_14755);
nor UO_862 (O_862,N_14797,N_14815);
or UO_863 (O_863,N_14750,N_14954);
xnor UO_864 (O_864,N_14927,N_14750);
or UO_865 (O_865,N_14991,N_14945);
and UO_866 (O_866,N_14998,N_14912);
nor UO_867 (O_867,N_14839,N_14807);
xnor UO_868 (O_868,N_14777,N_14977);
xnor UO_869 (O_869,N_14921,N_14774);
nor UO_870 (O_870,N_14758,N_14983);
xor UO_871 (O_871,N_14809,N_14959);
and UO_872 (O_872,N_14822,N_14937);
and UO_873 (O_873,N_14943,N_14924);
or UO_874 (O_874,N_14782,N_14948);
nand UO_875 (O_875,N_14964,N_14980);
nor UO_876 (O_876,N_14944,N_14779);
or UO_877 (O_877,N_14840,N_14992);
xor UO_878 (O_878,N_14817,N_14765);
nand UO_879 (O_879,N_14827,N_14811);
or UO_880 (O_880,N_14863,N_14869);
nor UO_881 (O_881,N_14829,N_14859);
and UO_882 (O_882,N_14908,N_14933);
nor UO_883 (O_883,N_14883,N_14988);
xnor UO_884 (O_884,N_14794,N_14980);
and UO_885 (O_885,N_14783,N_14845);
nand UO_886 (O_886,N_14923,N_14796);
xnor UO_887 (O_887,N_14833,N_14969);
nor UO_888 (O_888,N_14795,N_14845);
nor UO_889 (O_889,N_14764,N_14810);
nor UO_890 (O_890,N_14927,N_14763);
or UO_891 (O_891,N_14781,N_14896);
nor UO_892 (O_892,N_14785,N_14954);
nor UO_893 (O_893,N_14862,N_14890);
nand UO_894 (O_894,N_14797,N_14957);
or UO_895 (O_895,N_14966,N_14866);
nor UO_896 (O_896,N_14964,N_14847);
xnor UO_897 (O_897,N_14956,N_14818);
or UO_898 (O_898,N_14970,N_14803);
xnor UO_899 (O_899,N_14829,N_14853);
xnor UO_900 (O_900,N_14826,N_14878);
xnor UO_901 (O_901,N_14912,N_14982);
nand UO_902 (O_902,N_14852,N_14949);
nand UO_903 (O_903,N_14939,N_14998);
and UO_904 (O_904,N_14792,N_14921);
xor UO_905 (O_905,N_14912,N_14907);
and UO_906 (O_906,N_14845,N_14936);
xnor UO_907 (O_907,N_14923,N_14835);
xnor UO_908 (O_908,N_14851,N_14915);
nor UO_909 (O_909,N_14871,N_14866);
xnor UO_910 (O_910,N_14870,N_14849);
nand UO_911 (O_911,N_14911,N_14871);
xnor UO_912 (O_912,N_14816,N_14767);
or UO_913 (O_913,N_14888,N_14803);
nor UO_914 (O_914,N_14780,N_14786);
or UO_915 (O_915,N_14985,N_14898);
xor UO_916 (O_916,N_14878,N_14800);
and UO_917 (O_917,N_14832,N_14866);
nor UO_918 (O_918,N_14985,N_14961);
and UO_919 (O_919,N_14904,N_14932);
nor UO_920 (O_920,N_14974,N_14924);
nor UO_921 (O_921,N_14796,N_14982);
nand UO_922 (O_922,N_14951,N_14979);
nand UO_923 (O_923,N_14903,N_14789);
and UO_924 (O_924,N_14759,N_14806);
or UO_925 (O_925,N_14965,N_14939);
nand UO_926 (O_926,N_14894,N_14785);
nor UO_927 (O_927,N_14788,N_14864);
or UO_928 (O_928,N_14815,N_14776);
or UO_929 (O_929,N_14759,N_14875);
xor UO_930 (O_930,N_14873,N_14872);
or UO_931 (O_931,N_14921,N_14938);
xnor UO_932 (O_932,N_14935,N_14827);
nor UO_933 (O_933,N_14998,N_14966);
nor UO_934 (O_934,N_14790,N_14799);
xor UO_935 (O_935,N_14841,N_14903);
nand UO_936 (O_936,N_14885,N_14872);
and UO_937 (O_937,N_14790,N_14796);
nand UO_938 (O_938,N_14970,N_14762);
and UO_939 (O_939,N_14959,N_14812);
nor UO_940 (O_940,N_14863,N_14784);
and UO_941 (O_941,N_14848,N_14823);
xor UO_942 (O_942,N_14848,N_14873);
nor UO_943 (O_943,N_14884,N_14817);
nor UO_944 (O_944,N_14875,N_14907);
and UO_945 (O_945,N_14986,N_14780);
and UO_946 (O_946,N_14956,N_14881);
or UO_947 (O_947,N_14824,N_14905);
or UO_948 (O_948,N_14757,N_14755);
and UO_949 (O_949,N_14800,N_14921);
nor UO_950 (O_950,N_14784,N_14962);
and UO_951 (O_951,N_14864,N_14750);
xor UO_952 (O_952,N_14827,N_14788);
nand UO_953 (O_953,N_14830,N_14844);
and UO_954 (O_954,N_14949,N_14986);
or UO_955 (O_955,N_14861,N_14827);
and UO_956 (O_956,N_14945,N_14912);
and UO_957 (O_957,N_14942,N_14973);
and UO_958 (O_958,N_14935,N_14825);
nor UO_959 (O_959,N_14758,N_14920);
or UO_960 (O_960,N_14955,N_14797);
or UO_961 (O_961,N_14892,N_14921);
nor UO_962 (O_962,N_14905,N_14786);
nor UO_963 (O_963,N_14918,N_14812);
and UO_964 (O_964,N_14929,N_14970);
and UO_965 (O_965,N_14992,N_14847);
or UO_966 (O_966,N_14786,N_14958);
or UO_967 (O_967,N_14918,N_14946);
and UO_968 (O_968,N_14778,N_14909);
xnor UO_969 (O_969,N_14831,N_14798);
and UO_970 (O_970,N_14968,N_14918);
nor UO_971 (O_971,N_14832,N_14838);
nor UO_972 (O_972,N_14905,N_14920);
nor UO_973 (O_973,N_14938,N_14813);
or UO_974 (O_974,N_14815,N_14844);
nand UO_975 (O_975,N_14806,N_14758);
xor UO_976 (O_976,N_14889,N_14774);
and UO_977 (O_977,N_14884,N_14968);
xnor UO_978 (O_978,N_14827,N_14779);
or UO_979 (O_979,N_14869,N_14795);
nand UO_980 (O_980,N_14946,N_14875);
nor UO_981 (O_981,N_14958,N_14984);
xor UO_982 (O_982,N_14937,N_14968);
nand UO_983 (O_983,N_14873,N_14936);
and UO_984 (O_984,N_14876,N_14921);
xor UO_985 (O_985,N_14998,N_14769);
and UO_986 (O_986,N_14755,N_14801);
and UO_987 (O_987,N_14949,N_14907);
nand UO_988 (O_988,N_14788,N_14983);
or UO_989 (O_989,N_14784,N_14800);
xor UO_990 (O_990,N_14967,N_14811);
xnor UO_991 (O_991,N_14814,N_14850);
nand UO_992 (O_992,N_14790,N_14869);
nor UO_993 (O_993,N_14840,N_14968);
or UO_994 (O_994,N_14930,N_14831);
nand UO_995 (O_995,N_14752,N_14971);
nor UO_996 (O_996,N_14957,N_14872);
nor UO_997 (O_997,N_14826,N_14795);
xor UO_998 (O_998,N_14804,N_14773);
and UO_999 (O_999,N_14993,N_14837);
xor UO_1000 (O_1000,N_14795,N_14993);
or UO_1001 (O_1001,N_14899,N_14820);
xnor UO_1002 (O_1002,N_14764,N_14756);
and UO_1003 (O_1003,N_14751,N_14875);
and UO_1004 (O_1004,N_14973,N_14911);
nand UO_1005 (O_1005,N_14830,N_14939);
nor UO_1006 (O_1006,N_14948,N_14934);
and UO_1007 (O_1007,N_14762,N_14945);
and UO_1008 (O_1008,N_14976,N_14792);
or UO_1009 (O_1009,N_14898,N_14870);
and UO_1010 (O_1010,N_14938,N_14949);
xnor UO_1011 (O_1011,N_14910,N_14825);
nor UO_1012 (O_1012,N_14817,N_14984);
and UO_1013 (O_1013,N_14930,N_14810);
xor UO_1014 (O_1014,N_14844,N_14752);
or UO_1015 (O_1015,N_14760,N_14874);
nand UO_1016 (O_1016,N_14923,N_14895);
and UO_1017 (O_1017,N_14905,N_14938);
xor UO_1018 (O_1018,N_14855,N_14796);
or UO_1019 (O_1019,N_14998,N_14947);
xor UO_1020 (O_1020,N_14799,N_14866);
and UO_1021 (O_1021,N_14787,N_14854);
nor UO_1022 (O_1022,N_14957,N_14857);
xnor UO_1023 (O_1023,N_14925,N_14900);
or UO_1024 (O_1024,N_14972,N_14901);
and UO_1025 (O_1025,N_14858,N_14938);
nor UO_1026 (O_1026,N_14768,N_14876);
nand UO_1027 (O_1027,N_14848,N_14830);
nand UO_1028 (O_1028,N_14869,N_14804);
and UO_1029 (O_1029,N_14751,N_14948);
or UO_1030 (O_1030,N_14813,N_14947);
nor UO_1031 (O_1031,N_14832,N_14954);
or UO_1032 (O_1032,N_14778,N_14913);
xnor UO_1033 (O_1033,N_14783,N_14945);
nor UO_1034 (O_1034,N_14758,N_14814);
xor UO_1035 (O_1035,N_14758,N_14937);
xor UO_1036 (O_1036,N_14864,N_14874);
and UO_1037 (O_1037,N_14894,N_14759);
nand UO_1038 (O_1038,N_14977,N_14805);
nor UO_1039 (O_1039,N_14782,N_14976);
nand UO_1040 (O_1040,N_14921,N_14910);
and UO_1041 (O_1041,N_14939,N_14825);
xnor UO_1042 (O_1042,N_14989,N_14783);
nand UO_1043 (O_1043,N_14966,N_14755);
nor UO_1044 (O_1044,N_14924,N_14872);
xor UO_1045 (O_1045,N_14886,N_14877);
nand UO_1046 (O_1046,N_14805,N_14818);
and UO_1047 (O_1047,N_14787,N_14837);
xnor UO_1048 (O_1048,N_14859,N_14934);
or UO_1049 (O_1049,N_14860,N_14936);
or UO_1050 (O_1050,N_14930,N_14894);
and UO_1051 (O_1051,N_14871,N_14926);
nor UO_1052 (O_1052,N_14929,N_14853);
or UO_1053 (O_1053,N_14886,N_14934);
and UO_1054 (O_1054,N_14860,N_14857);
nand UO_1055 (O_1055,N_14935,N_14806);
nand UO_1056 (O_1056,N_14950,N_14769);
nor UO_1057 (O_1057,N_14829,N_14933);
nand UO_1058 (O_1058,N_14937,N_14871);
xor UO_1059 (O_1059,N_14774,N_14833);
and UO_1060 (O_1060,N_14861,N_14818);
xnor UO_1061 (O_1061,N_14795,N_14879);
or UO_1062 (O_1062,N_14886,N_14805);
or UO_1063 (O_1063,N_14796,N_14785);
xnor UO_1064 (O_1064,N_14836,N_14894);
or UO_1065 (O_1065,N_14906,N_14961);
nor UO_1066 (O_1066,N_14803,N_14995);
xnor UO_1067 (O_1067,N_14885,N_14754);
xnor UO_1068 (O_1068,N_14895,N_14905);
and UO_1069 (O_1069,N_14884,N_14757);
nand UO_1070 (O_1070,N_14874,N_14934);
or UO_1071 (O_1071,N_14906,N_14761);
nor UO_1072 (O_1072,N_14809,N_14942);
or UO_1073 (O_1073,N_14778,N_14770);
xnor UO_1074 (O_1074,N_14875,N_14813);
xor UO_1075 (O_1075,N_14915,N_14991);
xor UO_1076 (O_1076,N_14782,N_14915);
xnor UO_1077 (O_1077,N_14897,N_14938);
nor UO_1078 (O_1078,N_14868,N_14854);
xor UO_1079 (O_1079,N_14972,N_14941);
xnor UO_1080 (O_1080,N_14920,N_14923);
nand UO_1081 (O_1081,N_14900,N_14827);
nand UO_1082 (O_1082,N_14968,N_14843);
nor UO_1083 (O_1083,N_14903,N_14952);
xnor UO_1084 (O_1084,N_14765,N_14886);
nor UO_1085 (O_1085,N_14880,N_14889);
or UO_1086 (O_1086,N_14865,N_14788);
xor UO_1087 (O_1087,N_14894,N_14908);
nand UO_1088 (O_1088,N_14925,N_14766);
nor UO_1089 (O_1089,N_14882,N_14921);
nor UO_1090 (O_1090,N_14826,N_14755);
or UO_1091 (O_1091,N_14924,N_14970);
and UO_1092 (O_1092,N_14858,N_14860);
nor UO_1093 (O_1093,N_14995,N_14909);
nor UO_1094 (O_1094,N_14948,N_14756);
xor UO_1095 (O_1095,N_14791,N_14932);
or UO_1096 (O_1096,N_14831,N_14855);
and UO_1097 (O_1097,N_14817,N_14766);
nand UO_1098 (O_1098,N_14796,N_14973);
xnor UO_1099 (O_1099,N_14934,N_14835);
nor UO_1100 (O_1100,N_14845,N_14864);
nor UO_1101 (O_1101,N_14933,N_14897);
xor UO_1102 (O_1102,N_14765,N_14994);
nor UO_1103 (O_1103,N_14890,N_14766);
or UO_1104 (O_1104,N_14810,N_14835);
xnor UO_1105 (O_1105,N_14875,N_14828);
nand UO_1106 (O_1106,N_14951,N_14806);
xnor UO_1107 (O_1107,N_14900,N_14767);
nand UO_1108 (O_1108,N_14875,N_14891);
and UO_1109 (O_1109,N_14978,N_14875);
xor UO_1110 (O_1110,N_14890,N_14806);
and UO_1111 (O_1111,N_14851,N_14987);
or UO_1112 (O_1112,N_14875,N_14939);
and UO_1113 (O_1113,N_14753,N_14890);
and UO_1114 (O_1114,N_14986,N_14783);
or UO_1115 (O_1115,N_14998,N_14987);
nor UO_1116 (O_1116,N_14951,N_14904);
or UO_1117 (O_1117,N_14839,N_14907);
xor UO_1118 (O_1118,N_14879,N_14942);
nor UO_1119 (O_1119,N_14996,N_14850);
nand UO_1120 (O_1120,N_14850,N_14970);
and UO_1121 (O_1121,N_14973,N_14810);
nor UO_1122 (O_1122,N_14790,N_14825);
and UO_1123 (O_1123,N_14820,N_14810);
xor UO_1124 (O_1124,N_14841,N_14936);
nand UO_1125 (O_1125,N_14946,N_14911);
or UO_1126 (O_1126,N_14801,N_14833);
xnor UO_1127 (O_1127,N_14890,N_14788);
or UO_1128 (O_1128,N_14770,N_14869);
nor UO_1129 (O_1129,N_14959,N_14943);
or UO_1130 (O_1130,N_14944,N_14880);
nand UO_1131 (O_1131,N_14779,N_14774);
nand UO_1132 (O_1132,N_14882,N_14852);
or UO_1133 (O_1133,N_14945,N_14950);
and UO_1134 (O_1134,N_14778,N_14906);
and UO_1135 (O_1135,N_14802,N_14914);
nor UO_1136 (O_1136,N_14872,N_14886);
nor UO_1137 (O_1137,N_14987,N_14803);
or UO_1138 (O_1138,N_14869,N_14797);
and UO_1139 (O_1139,N_14816,N_14763);
xor UO_1140 (O_1140,N_14968,N_14891);
nand UO_1141 (O_1141,N_14767,N_14895);
nand UO_1142 (O_1142,N_14795,N_14896);
or UO_1143 (O_1143,N_14855,N_14786);
or UO_1144 (O_1144,N_14809,N_14753);
xor UO_1145 (O_1145,N_14888,N_14780);
nand UO_1146 (O_1146,N_14857,N_14893);
or UO_1147 (O_1147,N_14872,N_14796);
nor UO_1148 (O_1148,N_14753,N_14773);
nand UO_1149 (O_1149,N_14776,N_14897);
xnor UO_1150 (O_1150,N_14872,N_14862);
nand UO_1151 (O_1151,N_14873,N_14952);
xor UO_1152 (O_1152,N_14940,N_14946);
xor UO_1153 (O_1153,N_14907,N_14942);
or UO_1154 (O_1154,N_14752,N_14912);
nand UO_1155 (O_1155,N_14963,N_14969);
nor UO_1156 (O_1156,N_14774,N_14971);
nand UO_1157 (O_1157,N_14989,N_14837);
and UO_1158 (O_1158,N_14829,N_14811);
nor UO_1159 (O_1159,N_14940,N_14788);
nand UO_1160 (O_1160,N_14869,N_14791);
and UO_1161 (O_1161,N_14892,N_14984);
and UO_1162 (O_1162,N_14857,N_14827);
and UO_1163 (O_1163,N_14756,N_14896);
nor UO_1164 (O_1164,N_14845,N_14925);
or UO_1165 (O_1165,N_14974,N_14896);
xnor UO_1166 (O_1166,N_14848,N_14996);
xor UO_1167 (O_1167,N_14904,N_14989);
or UO_1168 (O_1168,N_14853,N_14889);
and UO_1169 (O_1169,N_14753,N_14788);
nor UO_1170 (O_1170,N_14883,N_14911);
and UO_1171 (O_1171,N_14870,N_14904);
or UO_1172 (O_1172,N_14893,N_14865);
and UO_1173 (O_1173,N_14804,N_14948);
and UO_1174 (O_1174,N_14866,N_14784);
nor UO_1175 (O_1175,N_14861,N_14968);
and UO_1176 (O_1176,N_14926,N_14920);
or UO_1177 (O_1177,N_14850,N_14766);
nor UO_1178 (O_1178,N_14828,N_14922);
nor UO_1179 (O_1179,N_14751,N_14932);
or UO_1180 (O_1180,N_14755,N_14869);
nor UO_1181 (O_1181,N_14913,N_14873);
nor UO_1182 (O_1182,N_14805,N_14903);
or UO_1183 (O_1183,N_14767,N_14921);
and UO_1184 (O_1184,N_14975,N_14830);
and UO_1185 (O_1185,N_14830,N_14751);
and UO_1186 (O_1186,N_14779,N_14880);
and UO_1187 (O_1187,N_14943,N_14874);
nor UO_1188 (O_1188,N_14822,N_14930);
xnor UO_1189 (O_1189,N_14999,N_14872);
xnor UO_1190 (O_1190,N_14930,N_14823);
xor UO_1191 (O_1191,N_14885,N_14777);
nand UO_1192 (O_1192,N_14903,N_14828);
or UO_1193 (O_1193,N_14803,N_14793);
and UO_1194 (O_1194,N_14976,N_14974);
nor UO_1195 (O_1195,N_14781,N_14807);
or UO_1196 (O_1196,N_14955,N_14864);
nand UO_1197 (O_1197,N_14872,N_14905);
nand UO_1198 (O_1198,N_14867,N_14804);
or UO_1199 (O_1199,N_14921,N_14878);
nor UO_1200 (O_1200,N_14888,N_14872);
and UO_1201 (O_1201,N_14936,N_14824);
and UO_1202 (O_1202,N_14831,N_14894);
or UO_1203 (O_1203,N_14991,N_14810);
and UO_1204 (O_1204,N_14869,N_14902);
nand UO_1205 (O_1205,N_14932,N_14948);
or UO_1206 (O_1206,N_14947,N_14810);
or UO_1207 (O_1207,N_14831,N_14871);
or UO_1208 (O_1208,N_14782,N_14795);
and UO_1209 (O_1209,N_14831,N_14971);
or UO_1210 (O_1210,N_14864,N_14782);
and UO_1211 (O_1211,N_14913,N_14752);
or UO_1212 (O_1212,N_14991,N_14972);
nand UO_1213 (O_1213,N_14774,N_14855);
or UO_1214 (O_1214,N_14889,N_14890);
xor UO_1215 (O_1215,N_14821,N_14952);
xor UO_1216 (O_1216,N_14863,N_14889);
or UO_1217 (O_1217,N_14956,N_14826);
and UO_1218 (O_1218,N_14773,N_14992);
nor UO_1219 (O_1219,N_14905,N_14780);
nor UO_1220 (O_1220,N_14881,N_14999);
or UO_1221 (O_1221,N_14816,N_14933);
nand UO_1222 (O_1222,N_14983,N_14822);
nor UO_1223 (O_1223,N_14966,N_14890);
or UO_1224 (O_1224,N_14812,N_14825);
nor UO_1225 (O_1225,N_14986,N_14768);
nor UO_1226 (O_1226,N_14947,N_14886);
nand UO_1227 (O_1227,N_14978,N_14897);
nand UO_1228 (O_1228,N_14778,N_14756);
nand UO_1229 (O_1229,N_14985,N_14782);
xor UO_1230 (O_1230,N_14894,N_14935);
and UO_1231 (O_1231,N_14955,N_14774);
nand UO_1232 (O_1232,N_14815,N_14875);
xnor UO_1233 (O_1233,N_14903,N_14923);
or UO_1234 (O_1234,N_14981,N_14790);
or UO_1235 (O_1235,N_14846,N_14880);
or UO_1236 (O_1236,N_14777,N_14884);
nand UO_1237 (O_1237,N_14962,N_14901);
and UO_1238 (O_1238,N_14795,N_14956);
and UO_1239 (O_1239,N_14795,N_14754);
nand UO_1240 (O_1240,N_14802,N_14750);
or UO_1241 (O_1241,N_14787,N_14985);
nand UO_1242 (O_1242,N_14779,N_14977);
or UO_1243 (O_1243,N_14922,N_14871);
or UO_1244 (O_1244,N_14776,N_14891);
and UO_1245 (O_1245,N_14835,N_14883);
and UO_1246 (O_1246,N_14966,N_14983);
nor UO_1247 (O_1247,N_14907,N_14755);
and UO_1248 (O_1248,N_14973,N_14974);
nand UO_1249 (O_1249,N_14827,N_14883);
nand UO_1250 (O_1250,N_14802,N_14920);
or UO_1251 (O_1251,N_14774,N_14886);
and UO_1252 (O_1252,N_14957,N_14984);
xor UO_1253 (O_1253,N_14981,N_14818);
nor UO_1254 (O_1254,N_14972,N_14879);
or UO_1255 (O_1255,N_14998,N_14877);
xnor UO_1256 (O_1256,N_14785,N_14968);
or UO_1257 (O_1257,N_14902,N_14996);
and UO_1258 (O_1258,N_14865,N_14930);
or UO_1259 (O_1259,N_14806,N_14813);
nand UO_1260 (O_1260,N_14945,N_14770);
or UO_1261 (O_1261,N_14973,N_14852);
and UO_1262 (O_1262,N_14883,N_14767);
nand UO_1263 (O_1263,N_14798,N_14977);
and UO_1264 (O_1264,N_14902,N_14918);
and UO_1265 (O_1265,N_14753,N_14778);
xnor UO_1266 (O_1266,N_14948,N_14952);
or UO_1267 (O_1267,N_14821,N_14894);
and UO_1268 (O_1268,N_14897,N_14798);
and UO_1269 (O_1269,N_14837,N_14940);
xnor UO_1270 (O_1270,N_14758,N_14839);
or UO_1271 (O_1271,N_14915,N_14826);
nor UO_1272 (O_1272,N_14769,N_14919);
or UO_1273 (O_1273,N_14966,N_14934);
nor UO_1274 (O_1274,N_14866,N_14880);
xnor UO_1275 (O_1275,N_14930,N_14951);
and UO_1276 (O_1276,N_14953,N_14995);
and UO_1277 (O_1277,N_14798,N_14753);
or UO_1278 (O_1278,N_14911,N_14998);
xnor UO_1279 (O_1279,N_14878,N_14854);
nand UO_1280 (O_1280,N_14808,N_14953);
and UO_1281 (O_1281,N_14873,N_14807);
xor UO_1282 (O_1282,N_14849,N_14821);
xor UO_1283 (O_1283,N_14962,N_14816);
nand UO_1284 (O_1284,N_14753,N_14938);
xnor UO_1285 (O_1285,N_14921,N_14916);
and UO_1286 (O_1286,N_14921,N_14852);
nand UO_1287 (O_1287,N_14987,N_14788);
xnor UO_1288 (O_1288,N_14823,N_14873);
nor UO_1289 (O_1289,N_14784,N_14786);
and UO_1290 (O_1290,N_14769,N_14962);
and UO_1291 (O_1291,N_14899,N_14877);
or UO_1292 (O_1292,N_14791,N_14911);
nand UO_1293 (O_1293,N_14922,N_14751);
and UO_1294 (O_1294,N_14908,N_14892);
and UO_1295 (O_1295,N_14868,N_14905);
or UO_1296 (O_1296,N_14766,N_14999);
or UO_1297 (O_1297,N_14964,N_14820);
nand UO_1298 (O_1298,N_14942,N_14917);
nor UO_1299 (O_1299,N_14826,N_14950);
nor UO_1300 (O_1300,N_14967,N_14815);
nand UO_1301 (O_1301,N_14979,N_14922);
nor UO_1302 (O_1302,N_14833,N_14915);
nand UO_1303 (O_1303,N_14859,N_14757);
nor UO_1304 (O_1304,N_14992,N_14875);
nor UO_1305 (O_1305,N_14832,N_14763);
and UO_1306 (O_1306,N_14883,N_14886);
xor UO_1307 (O_1307,N_14945,N_14947);
and UO_1308 (O_1308,N_14947,N_14801);
nor UO_1309 (O_1309,N_14922,N_14780);
or UO_1310 (O_1310,N_14957,N_14758);
xnor UO_1311 (O_1311,N_14889,N_14956);
or UO_1312 (O_1312,N_14989,N_14808);
nand UO_1313 (O_1313,N_14809,N_14962);
nand UO_1314 (O_1314,N_14977,N_14965);
nand UO_1315 (O_1315,N_14899,N_14778);
nand UO_1316 (O_1316,N_14852,N_14827);
nor UO_1317 (O_1317,N_14763,N_14752);
nand UO_1318 (O_1318,N_14893,N_14970);
nand UO_1319 (O_1319,N_14760,N_14936);
nand UO_1320 (O_1320,N_14874,N_14939);
or UO_1321 (O_1321,N_14933,N_14776);
nor UO_1322 (O_1322,N_14915,N_14756);
nand UO_1323 (O_1323,N_14883,N_14948);
xnor UO_1324 (O_1324,N_14916,N_14906);
or UO_1325 (O_1325,N_14915,N_14908);
nand UO_1326 (O_1326,N_14852,N_14881);
or UO_1327 (O_1327,N_14802,N_14918);
or UO_1328 (O_1328,N_14980,N_14801);
and UO_1329 (O_1329,N_14901,N_14862);
nand UO_1330 (O_1330,N_14767,N_14819);
or UO_1331 (O_1331,N_14876,N_14971);
xnor UO_1332 (O_1332,N_14909,N_14936);
nor UO_1333 (O_1333,N_14757,N_14988);
nor UO_1334 (O_1334,N_14958,N_14935);
nand UO_1335 (O_1335,N_14913,N_14931);
or UO_1336 (O_1336,N_14895,N_14944);
and UO_1337 (O_1337,N_14916,N_14968);
nor UO_1338 (O_1338,N_14799,N_14780);
nor UO_1339 (O_1339,N_14915,N_14891);
xnor UO_1340 (O_1340,N_14985,N_14964);
or UO_1341 (O_1341,N_14815,N_14891);
nor UO_1342 (O_1342,N_14759,N_14764);
or UO_1343 (O_1343,N_14826,N_14836);
nor UO_1344 (O_1344,N_14980,N_14978);
nand UO_1345 (O_1345,N_14963,N_14843);
nor UO_1346 (O_1346,N_14908,N_14796);
and UO_1347 (O_1347,N_14939,N_14783);
and UO_1348 (O_1348,N_14975,N_14951);
nor UO_1349 (O_1349,N_14856,N_14887);
nand UO_1350 (O_1350,N_14942,N_14815);
xor UO_1351 (O_1351,N_14857,N_14923);
or UO_1352 (O_1352,N_14872,N_14821);
and UO_1353 (O_1353,N_14916,N_14853);
and UO_1354 (O_1354,N_14773,N_14916);
nor UO_1355 (O_1355,N_14832,N_14791);
nand UO_1356 (O_1356,N_14997,N_14769);
nand UO_1357 (O_1357,N_14833,N_14900);
xnor UO_1358 (O_1358,N_14913,N_14885);
or UO_1359 (O_1359,N_14863,N_14880);
or UO_1360 (O_1360,N_14756,N_14867);
xnor UO_1361 (O_1361,N_14786,N_14992);
xor UO_1362 (O_1362,N_14769,N_14875);
nor UO_1363 (O_1363,N_14846,N_14994);
or UO_1364 (O_1364,N_14995,N_14902);
nand UO_1365 (O_1365,N_14889,N_14850);
and UO_1366 (O_1366,N_14847,N_14903);
nor UO_1367 (O_1367,N_14924,N_14766);
nor UO_1368 (O_1368,N_14856,N_14838);
or UO_1369 (O_1369,N_14909,N_14804);
or UO_1370 (O_1370,N_14755,N_14779);
xor UO_1371 (O_1371,N_14833,N_14757);
and UO_1372 (O_1372,N_14914,N_14835);
xnor UO_1373 (O_1373,N_14868,N_14873);
nor UO_1374 (O_1374,N_14769,N_14851);
nand UO_1375 (O_1375,N_14779,N_14895);
xnor UO_1376 (O_1376,N_14766,N_14946);
and UO_1377 (O_1377,N_14796,N_14940);
and UO_1378 (O_1378,N_14980,N_14818);
or UO_1379 (O_1379,N_14850,N_14886);
and UO_1380 (O_1380,N_14836,N_14814);
or UO_1381 (O_1381,N_14906,N_14948);
nand UO_1382 (O_1382,N_14797,N_14990);
and UO_1383 (O_1383,N_14964,N_14896);
or UO_1384 (O_1384,N_14941,N_14919);
xor UO_1385 (O_1385,N_14882,N_14914);
or UO_1386 (O_1386,N_14962,N_14818);
nand UO_1387 (O_1387,N_14832,N_14837);
nor UO_1388 (O_1388,N_14945,N_14972);
xnor UO_1389 (O_1389,N_14911,N_14933);
nand UO_1390 (O_1390,N_14972,N_14880);
nor UO_1391 (O_1391,N_14795,N_14772);
xor UO_1392 (O_1392,N_14919,N_14751);
and UO_1393 (O_1393,N_14921,N_14821);
xnor UO_1394 (O_1394,N_14844,N_14778);
xnor UO_1395 (O_1395,N_14825,N_14945);
and UO_1396 (O_1396,N_14753,N_14970);
xor UO_1397 (O_1397,N_14820,N_14784);
or UO_1398 (O_1398,N_14777,N_14989);
or UO_1399 (O_1399,N_14818,N_14966);
and UO_1400 (O_1400,N_14998,N_14825);
nand UO_1401 (O_1401,N_14974,N_14952);
nand UO_1402 (O_1402,N_14869,N_14874);
or UO_1403 (O_1403,N_14835,N_14951);
nor UO_1404 (O_1404,N_14886,N_14855);
nand UO_1405 (O_1405,N_14910,N_14867);
xnor UO_1406 (O_1406,N_14965,N_14755);
xnor UO_1407 (O_1407,N_14763,N_14874);
xor UO_1408 (O_1408,N_14975,N_14821);
and UO_1409 (O_1409,N_14989,N_14891);
nor UO_1410 (O_1410,N_14957,N_14855);
or UO_1411 (O_1411,N_14944,N_14857);
nor UO_1412 (O_1412,N_14902,N_14951);
xor UO_1413 (O_1413,N_14962,N_14892);
nor UO_1414 (O_1414,N_14969,N_14792);
nor UO_1415 (O_1415,N_14983,N_14907);
and UO_1416 (O_1416,N_14882,N_14958);
nor UO_1417 (O_1417,N_14934,N_14860);
nand UO_1418 (O_1418,N_14815,N_14938);
xor UO_1419 (O_1419,N_14954,N_14883);
xor UO_1420 (O_1420,N_14987,N_14865);
and UO_1421 (O_1421,N_14974,N_14889);
and UO_1422 (O_1422,N_14819,N_14984);
nand UO_1423 (O_1423,N_14822,N_14927);
or UO_1424 (O_1424,N_14868,N_14845);
nand UO_1425 (O_1425,N_14808,N_14870);
and UO_1426 (O_1426,N_14802,N_14784);
and UO_1427 (O_1427,N_14999,N_14800);
nor UO_1428 (O_1428,N_14872,N_14837);
nand UO_1429 (O_1429,N_14889,N_14966);
xnor UO_1430 (O_1430,N_14828,N_14870);
nand UO_1431 (O_1431,N_14881,N_14991);
and UO_1432 (O_1432,N_14873,N_14810);
or UO_1433 (O_1433,N_14898,N_14918);
nand UO_1434 (O_1434,N_14888,N_14753);
nor UO_1435 (O_1435,N_14897,N_14900);
nor UO_1436 (O_1436,N_14935,N_14907);
and UO_1437 (O_1437,N_14964,N_14959);
nand UO_1438 (O_1438,N_14758,N_14886);
nor UO_1439 (O_1439,N_14981,N_14821);
xor UO_1440 (O_1440,N_14896,N_14930);
and UO_1441 (O_1441,N_14947,N_14990);
nor UO_1442 (O_1442,N_14994,N_14774);
nor UO_1443 (O_1443,N_14798,N_14761);
and UO_1444 (O_1444,N_14914,N_14783);
nor UO_1445 (O_1445,N_14872,N_14818);
and UO_1446 (O_1446,N_14988,N_14992);
and UO_1447 (O_1447,N_14925,N_14975);
xnor UO_1448 (O_1448,N_14752,N_14920);
or UO_1449 (O_1449,N_14855,N_14966);
nand UO_1450 (O_1450,N_14936,N_14785);
or UO_1451 (O_1451,N_14797,N_14959);
nand UO_1452 (O_1452,N_14966,N_14767);
nand UO_1453 (O_1453,N_14781,N_14859);
or UO_1454 (O_1454,N_14888,N_14922);
nor UO_1455 (O_1455,N_14767,N_14864);
nand UO_1456 (O_1456,N_14897,N_14998);
and UO_1457 (O_1457,N_14801,N_14778);
or UO_1458 (O_1458,N_14831,N_14969);
xor UO_1459 (O_1459,N_14861,N_14938);
and UO_1460 (O_1460,N_14900,N_14830);
nor UO_1461 (O_1461,N_14995,N_14844);
nand UO_1462 (O_1462,N_14978,N_14757);
and UO_1463 (O_1463,N_14916,N_14839);
xor UO_1464 (O_1464,N_14999,N_14996);
nor UO_1465 (O_1465,N_14881,N_14790);
and UO_1466 (O_1466,N_14987,N_14868);
xor UO_1467 (O_1467,N_14811,N_14911);
or UO_1468 (O_1468,N_14864,N_14795);
nor UO_1469 (O_1469,N_14757,N_14981);
xnor UO_1470 (O_1470,N_14848,N_14831);
xor UO_1471 (O_1471,N_14887,N_14807);
nand UO_1472 (O_1472,N_14812,N_14926);
or UO_1473 (O_1473,N_14948,N_14847);
nor UO_1474 (O_1474,N_14964,N_14815);
or UO_1475 (O_1475,N_14756,N_14769);
xnor UO_1476 (O_1476,N_14843,N_14854);
xor UO_1477 (O_1477,N_14977,N_14790);
nor UO_1478 (O_1478,N_14757,N_14890);
and UO_1479 (O_1479,N_14793,N_14883);
nor UO_1480 (O_1480,N_14832,N_14879);
nand UO_1481 (O_1481,N_14873,N_14763);
and UO_1482 (O_1482,N_14908,N_14912);
or UO_1483 (O_1483,N_14785,N_14863);
xnor UO_1484 (O_1484,N_14921,N_14762);
xor UO_1485 (O_1485,N_14976,N_14828);
nor UO_1486 (O_1486,N_14855,N_14889);
xor UO_1487 (O_1487,N_14821,N_14822);
or UO_1488 (O_1488,N_14949,N_14809);
nor UO_1489 (O_1489,N_14976,N_14829);
xnor UO_1490 (O_1490,N_14918,N_14862);
xnor UO_1491 (O_1491,N_14915,N_14911);
xor UO_1492 (O_1492,N_14882,N_14971);
nand UO_1493 (O_1493,N_14944,N_14911);
and UO_1494 (O_1494,N_14835,N_14966);
nor UO_1495 (O_1495,N_14804,N_14973);
nand UO_1496 (O_1496,N_14850,N_14868);
xor UO_1497 (O_1497,N_14908,N_14891);
and UO_1498 (O_1498,N_14757,N_14751);
or UO_1499 (O_1499,N_14767,N_14754);
nor UO_1500 (O_1500,N_14858,N_14918);
or UO_1501 (O_1501,N_14955,N_14755);
or UO_1502 (O_1502,N_14943,N_14847);
nor UO_1503 (O_1503,N_14975,N_14972);
and UO_1504 (O_1504,N_14867,N_14817);
xnor UO_1505 (O_1505,N_14875,N_14954);
and UO_1506 (O_1506,N_14906,N_14838);
and UO_1507 (O_1507,N_14908,N_14904);
nand UO_1508 (O_1508,N_14986,N_14757);
and UO_1509 (O_1509,N_14814,N_14770);
nor UO_1510 (O_1510,N_14780,N_14832);
or UO_1511 (O_1511,N_14829,N_14894);
nand UO_1512 (O_1512,N_14879,N_14831);
xor UO_1513 (O_1513,N_14891,N_14918);
and UO_1514 (O_1514,N_14923,N_14978);
and UO_1515 (O_1515,N_14769,N_14816);
nor UO_1516 (O_1516,N_14826,N_14777);
nor UO_1517 (O_1517,N_14932,N_14922);
and UO_1518 (O_1518,N_14986,N_14777);
or UO_1519 (O_1519,N_14870,N_14938);
nor UO_1520 (O_1520,N_14925,N_14818);
nand UO_1521 (O_1521,N_14764,N_14952);
and UO_1522 (O_1522,N_14901,N_14958);
nor UO_1523 (O_1523,N_14882,N_14811);
xnor UO_1524 (O_1524,N_14891,N_14932);
nor UO_1525 (O_1525,N_14990,N_14810);
nor UO_1526 (O_1526,N_14812,N_14841);
or UO_1527 (O_1527,N_14915,N_14771);
and UO_1528 (O_1528,N_14774,N_14789);
nand UO_1529 (O_1529,N_14991,N_14952);
nor UO_1530 (O_1530,N_14880,N_14796);
or UO_1531 (O_1531,N_14892,N_14993);
xnor UO_1532 (O_1532,N_14923,N_14799);
xnor UO_1533 (O_1533,N_14811,N_14871);
nor UO_1534 (O_1534,N_14946,N_14912);
xor UO_1535 (O_1535,N_14772,N_14841);
nor UO_1536 (O_1536,N_14868,N_14932);
xor UO_1537 (O_1537,N_14824,N_14904);
xnor UO_1538 (O_1538,N_14911,N_14817);
nor UO_1539 (O_1539,N_14823,N_14806);
xnor UO_1540 (O_1540,N_14975,N_14787);
nor UO_1541 (O_1541,N_14898,N_14908);
nor UO_1542 (O_1542,N_14815,N_14834);
and UO_1543 (O_1543,N_14758,N_14928);
xor UO_1544 (O_1544,N_14959,N_14930);
or UO_1545 (O_1545,N_14936,N_14975);
xnor UO_1546 (O_1546,N_14814,N_14752);
xnor UO_1547 (O_1547,N_14776,N_14949);
or UO_1548 (O_1548,N_14898,N_14810);
xor UO_1549 (O_1549,N_14889,N_14808);
and UO_1550 (O_1550,N_14922,N_14755);
and UO_1551 (O_1551,N_14996,N_14920);
nand UO_1552 (O_1552,N_14755,N_14876);
nor UO_1553 (O_1553,N_14817,N_14809);
xor UO_1554 (O_1554,N_14901,N_14952);
nand UO_1555 (O_1555,N_14859,N_14933);
nand UO_1556 (O_1556,N_14976,N_14913);
and UO_1557 (O_1557,N_14790,N_14909);
nand UO_1558 (O_1558,N_14880,N_14770);
nand UO_1559 (O_1559,N_14888,N_14789);
xor UO_1560 (O_1560,N_14922,N_14936);
xor UO_1561 (O_1561,N_14971,N_14779);
xor UO_1562 (O_1562,N_14889,N_14913);
nor UO_1563 (O_1563,N_14895,N_14848);
nand UO_1564 (O_1564,N_14999,N_14867);
or UO_1565 (O_1565,N_14997,N_14830);
nand UO_1566 (O_1566,N_14847,N_14856);
nor UO_1567 (O_1567,N_14904,N_14900);
xor UO_1568 (O_1568,N_14944,N_14791);
or UO_1569 (O_1569,N_14981,N_14830);
xor UO_1570 (O_1570,N_14783,N_14998);
nand UO_1571 (O_1571,N_14982,N_14775);
and UO_1572 (O_1572,N_14988,N_14846);
nand UO_1573 (O_1573,N_14968,N_14774);
nand UO_1574 (O_1574,N_14782,N_14956);
xnor UO_1575 (O_1575,N_14960,N_14933);
nor UO_1576 (O_1576,N_14992,N_14768);
or UO_1577 (O_1577,N_14924,N_14927);
and UO_1578 (O_1578,N_14878,N_14823);
and UO_1579 (O_1579,N_14888,N_14899);
xor UO_1580 (O_1580,N_14844,N_14954);
nor UO_1581 (O_1581,N_14762,N_14857);
xnor UO_1582 (O_1582,N_14946,N_14902);
nor UO_1583 (O_1583,N_14937,N_14922);
and UO_1584 (O_1584,N_14957,N_14879);
or UO_1585 (O_1585,N_14883,N_14903);
and UO_1586 (O_1586,N_14825,N_14911);
nor UO_1587 (O_1587,N_14812,N_14884);
xor UO_1588 (O_1588,N_14968,N_14953);
or UO_1589 (O_1589,N_14926,N_14947);
and UO_1590 (O_1590,N_14897,N_14788);
nand UO_1591 (O_1591,N_14888,N_14778);
nand UO_1592 (O_1592,N_14765,N_14939);
nand UO_1593 (O_1593,N_14988,N_14767);
or UO_1594 (O_1594,N_14765,N_14965);
nor UO_1595 (O_1595,N_14958,N_14810);
nand UO_1596 (O_1596,N_14791,N_14862);
nor UO_1597 (O_1597,N_14953,N_14900);
or UO_1598 (O_1598,N_14801,N_14805);
nor UO_1599 (O_1599,N_14862,N_14991);
and UO_1600 (O_1600,N_14892,N_14822);
or UO_1601 (O_1601,N_14861,N_14979);
nor UO_1602 (O_1602,N_14951,N_14970);
and UO_1603 (O_1603,N_14882,N_14774);
xor UO_1604 (O_1604,N_14942,N_14874);
nor UO_1605 (O_1605,N_14942,N_14757);
or UO_1606 (O_1606,N_14808,N_14919);
and UO_1607 (O_1607,N_14887,N_14780);
xnor UO_1608 (O_1608,N_14961,N_14805);
or UO_1609 (O_1609,N_14979,N_14792);
or UO_1610 (O_1610,N_14994,N_14768);
or UO_1611 (O_1611,N_14974,N_14764);
nand UO_1612 (O_1612,N_14852,N_14815);
or UO_1613 (O_1613,N_14757,N_14837);
nor UO_1614 (O_1614,N_14773,N_14824);
and UO_1615 (O_1615,N_14836,N_14935);
nor UO_1616 (O_1616,N_14804,N_14996);
or UO_1617 (O_1617,N_14923,N_14950);
xnor UO_1618 (O_1618,N_14825,N_14916);
nor UO_1619 (O_1619,N_14859,N_14813);
xnor UO_1620 (O_1620,N_14958,N_14936);
and UO_1621 (O_1621,N_14865,N_14991);
and UO_1622 (O_1622,N_14753,N_14800);
and UO_1623 (O_1623,N_14917,N_14752);
or UO_1624 (O_1624,N_14864,N_14862);
xnor UO_1625 (O_1625,N_14755,N_14773);
nand UO_1626 (O_1626,N_14973,N_14969);
xnor UO_1627 (O_1627,N_14911,N_14773);
or UO_1628 (O_1628,N_14772,N_14840);
nor UO_1629 (O_1629,N_14902,N_14967);
nor UO_1630 (O_1630,N_14937,N_14995);
and UO_1631 (O_1631,N_14963,N_14958);
and UO_1632 (O_1632,N_14796,N_14983);
and UO_1633 (O_1633,N_14786,N_14869);
or UO_1634 (O_1634,N_14968,N_14761);
xnor UO_1635 (O_1635,N_14840,N_14911);
nand UO_1636 (O_1636,N_14812,N_14840);
nand UO_1637 (O_1637,N_14989,N_14896);
nor UO_1638 (O_1638,N_14832,N_14765);
or UO_1639 (O_1639,N_14754,N_14881);
xnor UO_1640 (O_1640,N_14761,N_14873);
or UO_1641 (O_1641,N_14812,N_14936);
xnor UO_1642 (O_1642,N_14945,N_14896);
xor UO_1643 (O_1643,N_14904,N_14928);
and UO_1644 (O_1644,N_14755,N_14827);
nor UO_1645 (O_1645,N_14771,N_14808);
nor UO_1646 (O_1646,N_14982,N_14916);
or UO_1647 (O_1647,N_14774,N_14870);
nand UO_1648 (O_1648,N_14941,N_14948);
and UO_1649 (O_1649,N_14750,N_14986);
and UO_1650 (O_1650,N_14952,N_14878);
nand UO_1651 (O_1651,N_14772,N_14958);
xnor UO_1652 (O_1652,N_14989,N_14981);
nand UO_1653 (O_1653,N_14950,N_14795);
xnor UO_1654 (O_1654,N_14875,N_14909);
nand UO_1655 (O_1655,N_14934,N_14828);
nand UO_1656 (O_1656,N_14993,N_14927);
or UO_1657 (O_1657,N_14791,N_14846);
or UO_1658 (O_1658,N_14952,N_14907);
nand UO_1659 (O_1659,N_14792,N_14750);
xnor UO_1660 (O_1660,N_14803,N_14973);
nor UO_1661 (O_1661,N_14974,N_14930);
and UO_1662 (O_1662,N_14868,N_14787);
nand UO_1663 (O_1663,N_14920,N_14993);
and UO_1664 (O_1664,N_14958,N_14820);
xnor UO_1665 (O_1665,N_14761,N_14989);
and UO_1666 (O_1666,N_14829,N_14885);
and UO_1667 (O_1667,N_14848,N_14913);
and UO_1668 (O_1668,N_14862,N_14886);
nor UO_1669 (O_1669,N_14879,N_14973);
and UO_1670 (O_1670,N_14962,N_14834);
nor UO_1671 (O_1671,N_14968,N_14836);
xnor UO_1672 (O_1672,N_14802,N_14832);
or UO_1673 (O_1673,N_14992,N_14757);
and UO_1674 (O_1674,N_14880,N_14896);
or UO_1675 (O_1675,N_14754,N_14808);
xnor UO_1676 (O_1676,N_14761,N_14911);
nor UO_1677 (O_1677,N_14920,N_14919);
nor UO_1678 (O_1678,N_14904,N_14933);
or UO_1679 (O_1679,N_14841,N_14934);
nor UO_1680 (O_1680,N_14750,N_14774);
or UO_1681 (O_1681,N_14873,N_14867);
and UO_1682 (O_1682,N_14800,N_14994);
xnor UO_1683 (O_1683,N_14994,N_14834);
nand UO_1684 (O_1684,N_14970,N_14908);
xnor UO_1685 (O_1685,N_14844,N_14851);
or UO_1686 (O_1686,N_14792,N_14799);
nand UO_1687 (O_1687,N_14958,N_14904);
xnor UO_1688 (O_1688,N_14847,N_14892);
and UO_1689 (O_1689,N_14884,N_14988);
and UO_1690 (O_1690,N_14773,N_14778);
or UO_1691 (O_1691,N_14791,N_14966);
nor UO_1692 (O_1692,N_14866,N_14935);
and UO_1693 (O_1693,N_14784,N_14795);
nor UO_1694 (O_1694,N_14997,N_14823);
nand UO_1695 (O_1695,N_14862,N_14825);
nand UO_1696 (O_1696,N_14963,N_14996);
xor UO_1697 (O_1697,N_14929,N_14873);
nor UO_1698 (O_1698,N_14783,N_14887);
xnor UO_1699 (O_1699,N_14845,N_14820);
nand UO_1700 (O_1700,N_14812,N_14991);
xor UO_1701 (O_1701,N_14757,N_14861);
nor UO_1702 (O_1702,N_14872,N_14950);
and UO_1703 (O_1703,N_14861,N_14862);
nor UO_1704 (O_1704,N_14905,N_14807);
and UO_1705 (O_1705,N_14751,N_14886);
nor UO_1706 (O_1706,N_14950,N_14875);
or UO_1707 (O_1707,N_14848,N_14953);
nor UO_1708 (O_1708,N_14957,N_14991);
and UO_1709 (O_1709,N_14798,N_14969);
and UO_1710 (O_1710,N_14894,N_14826);
or UO_1711 (O_1711,N_14880,N_14771);
nor UO_1712 (O_1712,N_14988,N_14958);
nor UO_1713 (O_1713,N_14821,N_14934);
or UO_1714 (O_1714,N_14876,N_14812);
nand UO_1715 (O_1715,N_14853,N_14763);
nor UO_1716 (O_1716,N_14775,N_14768);
nor UO_1717 (O_1717,N_14754,N_14868);
and UO_1718 (O_1718,N_14970,N_14815);
nand UO_1719 (O_1719,N_14878,N_14955);
or UO_1720 (O_1720,N_14878,N_14890);
and UO_1721 (O_1721,N_14787,N_14873);
or UO_1722 (O_1722,N_14860,N_14779);
or UO_1723 (O_1723,N_14915,N_14952);
nor UO_1724 (O_1724,N_14871,N_14868);
nand UO_1725 (O_1725,N_14935,N_14959);
nor UO_1726 (O_1726,N_14842,N_14969);
and UO_1727 (O_1727,N_14904,N_14913);
or UO_1728 (O_1728,N_14775,N_14774);
and UO_1729 (O_1729,N_14967,N_14972);
xor UO_1730 (O_1730,N_14964,N_14908);
nand UO_1731 (O_1731,N_14792,N_14826);
nand UO_1732 (O_1732,N_14797,N_14984);
nand UO_1733 (O_1733,N_14764,N_14771);
and UO_1734 (O_1734,N_14964,N_14755);
xor UO_1735 (O_1735,N_14827,N_14841);
xnor UO_1736 (O_1736,N_14759,N_14766);
xnor UO_1737 (O_1737,N_14814,N_14970);
nor UO_1738 (O_1738,N_14996,N_14979);
nand UO_1739 (O_1739,N_14910,N_14916);
nor UO_1740 (O_1740,N_14790,N_14892);
nor UO_1741 (O_1741,N_14917,N_14978);
nand UO_1742 (O_1742,N_14967,N_14857);
and UO_1743 (O_1743,N_14919,N_14784);
xnor UO_1744 (O_1744,N_14944,N_14851);
and UO_1745 (O_1745,N_14885,N_14794);
or UO_1746 (O_1746,N_14961,N_14937);
xnor UO_1747 (O_1747,N_14897,N_14804);
and UO_1748 (O_1748,N_14874,N_14941);
or UO_1749 (O_1749,N_14860,N_14753);
nand UO_1750 (O_1750,N_14756,N_14967);
xor UO_1751 (O_1751,N_14934,N_14950);
and UO_1752 (O_1752,N_14888,N_14801);
nand UO_1753 (O_1753,N_14979,N_14774);
nand UO_1754 (O_1754,N_14932,N_14786);
nor UO_1755 (O_1755,N_14892,N_14800);
nor UO_1756 (O_1756,N_14795,N_14940);
or UO_1757 (O_1757,N_14817,N_14769);
nor UO_1758 (O_1758,N_14791,N_14804);
or UO_1759 (O_1759,N_14910,N_14954);
nand UO_1760 (O_1760,N_14993,N_14919);
xnor UO_1761 (O_1761,N_14882,N_14784);
or UO_1762 (O_1762,N_14784,N_14936);
and UO_1763 (O_1763,N_14853,N_14775);
nand UO_1764 (O_1764,N_14778,N_14761);
xor UO_1765 (O_1765,N_14980,N_14760);
nand UO_1766 (O_1766,N_14953,N_14884);
xnor UO_1767 (O_1767,N_14874,N_14806);
and UO_1768 (O_1768,N_14919,N_14889);
or UO_1769 (O_1769,N_14978,N_14805);
nor UO_1770 (O_1770,N_14774,N_14890);
or UO_1771 (O_1771,N_14885,N_14832);
or UO_1772 (O_1772,N_14813,N_14881);
nand UO_1773 (O_1773,N_14893,N_14878);
nand UO_1774 (O_1774,N_14928,N_14973);
nand UO_1775 (O_1775,N_14796,N_14823);
nor UO_1776 (O_1776,N_14849,N_14896);
nor UO_1777 (O_1777,N_14815,N_14851);
and UO_1778 (O_1778,N_14840,N_14915);
nand UO_1779 (O_1779,N_14803,N_14750);
or UO_1780 (O_1780,N_14786,N_14952);
xnor UO_1781 (O_1781,N_14909,N_14969);
nand UO_1782 (O_1782,N_14879,N_14980);
nor UO_1783 (O_1783,N_14953,N_14927);
or UO_1784 (O_1784,N_14824,N_14827);
nor UO_1785 (O_1785,N_14775,N_14994);
or UO_1786 (O_1786,N_14993,N_14955);
or UO_1787 (O_1787,N_14984,N_14842);
or UO_1788 (O_1788,N_14878,N_14936);
nand UO_1789 (O_1789,N_14917,N_14828);
xor UO_1790 (O_1790,N_14944,N_14903);
or UO_1791 (O_1791,N_14875,N_14784);
or UO_1792 (O_1792,N_14838,N_14797);
or UO_1793 (O_1793,N_14789,N_14777);
xor UO_1794 (O_1794,N_14817,N_14781);
nand UO_1795 (O_1795,N_14988,N_14765);
and UO_1796 (O_1796,N_14978,N_14800);
or UO_1797 (O_1797,N_14836,N_14796);
xnor UO_1798 (O_1798,N_14835,N_14850);
or UO_1799 (O_1799,N_14773,N_14921);
and UO_1800 (O_1800,N_14909,N_14956);
nor UO_1801 (O_1801,N_14981,N_14826);
nand UO_1802 (O_1802,N_14774,N_14854);
and UO_1803 (O_1803,N_14914,N_14984);
nand UO_1804 (O_1804,N_14950,N_14786);
xor UO_1805 (O_1805,N_14890,N_14839);
nor UO_1806 (O_1806,N_14766,N_14809);
xor UO_1807 (O_1807,N_14916,N_14807);
nand UO_1808 (O_1808,N_14845,N_14775);
or UO_1809 (O_1809,N_14919,N_14811);
and UO_1810 (O_1810,N_14908,N_14761);
nor UO_1811 (O_1811,N_14880,N_14783);
and UO_1812 (O_1812,N_14791,N_14984);
nand UO_1813 (O_1813,N_14879,N_14913);
and UO_1814 (O_1814,N_14846,N_14756);
xor UO_1815 (O_1815,N_14931,N_14900);
nand UO_1816 (O_1816,N_14974,N_14959);
nand UO_1817 (O_1817,N_14840,N_14923);
and UO_1818 (O_1818,N_14904,N_14927);
or UO_1819 (O_1819,N_14859,N_14823);
xor UO_1820 (O_1820,N_14977,N_14825);
and UO_1821 (O_1821,N_14941,N_14871);
nor UO_1822 (O_1822,N_14890,N_14796);
and UO_1823 (O_1823,N_14879,N_14886);
and UO_1824 (O_1824,N_14934,N_14909);
nor UO_1825 (O_1825,N_14777,N_14945);
xor UO_1826 (O_1826,N_14980,N_14934);
or UO_1827 (O_1827,N_14858,N_14831);
and UO_1828 (O_1828,N_14751,N_14813);
and UO_1829 (O_1829,N_14822,N_14888);
and UO_1830 (O_1830,N_14905,N_14861);
nor UO_1831 (O_1831,N_14860,N_14786);
and UO_1832 (O_1832,N_14863,N_14962);
nand UO_1833 (O_1833,N_14975,N_14990);
xnor UO_1834 (O_1834,N_14784,N_14764);
and UO_1835 (O_1835,N_14942,N_14823);
xnor UO_1836 (O_1836,N_14919,N_14910);
xnor UO_1837 (O_1837,N_14987,N_14828);
and UO_1838 (O_1838,N_14988,N_14779);
nand UO_1839 (O_1839,N_14838,N_14792);
or UO_1840 (O_1840,N_14968,N_14757);
or UO_1841 (O_1841,N_14922,N_14782);
xnor UO_1842 (O_1842,N_14750,N_14917);
and UO_1843 (O_1843,N_14930,N_14821);
nand UO_1844 (O_1844,N_14880,N_14975);
xor UO_1845 (O_1845,N_14858,N_14975);
nor UO_1846 (O_1846,N_14806,N_14946);
xor UO_1847 (O_1847,N_14989,N_14869);
or UO_1848 (O_1848,N_14947,N_14771);
and UO_1849 (O_1849,N_14894,N_14867);
xnor UO_1850 (O_1850,N_14752,N_14968);
xnor UO_1851 (O_1851,N_14961,N_14771);
xnor UO_1852 (O_1852,N_14772,N_14973);
nand UO_1853 (O_1853,N_14928,N_14759);
nor UO_1854 (O_1854,N_14999,N_14919);
nor UO_1855 (O_1855,N_14798,N_14913);
and UO_1856 (O_1856,N_14816,N_14778);
and UO_1857 (O_1857,N_14874,N_14987);
and UO_1858 (O_1858,N_14915,N_14789);
or UO_1859 (O_1859,N_14943,N_14809);
and UO_1860 (O_1860,N_14819,N_14893);
nor UO_1861 (O_1861,N_14888,N_14879);
nand UO_1862 (O_1862,N_14759,N_14811);
xnor UO_1863 (O_1863,N_14799,N_14917);
xnor UO_1864 (O_1864,N_14972,N_14848);
nand UO_1865 (O_1865,N_14943,N_14827);
and UO_1866 (O_1866,N_14918,N_14917);
xor UO_1867 (O_1867,N_14942,N_14957);
xor UO_1868 (O_1868,N_14762,N_14948);
xnor UO_1869 (O_1869,N_14848,N_14910);
xnor UO_1870 (O_1870,N_14884,N_14944);
and UO_1871 (O_1871,N_14891,N_14814);
or UO_1872 (O_1872,N_14927,N_14875);
nand UO_1873 (O_1873,N_14795,N_14796);
xor UO_1874 (O_1874,N_14905,N_14849);
xor UO_1875 (O_1875,N_14845,N_14949);
nand UO_1876 (O_1876,N_14849,N_14750);
nand UO_1877 (O_1877,N_14779,N_14826);
and UO_1878 (O_1878,N_14941,N_14960);
xor UO_1879 (O_1879,N_14998,N_14941);
or UO_1880 (O_1880,N_14814,N_14807);
and UO_1881 (O_1881,N_14839,N_14857);
xnor UO_1882 (O_1882,N_14869,N_14798);
nor UO_1883 (O_1883,N_14818,N_14800);
and UO_1884 (O_1884,N_14870,N_14931);
nand UO_1885 (O_1885,N_14886,N_14990);
nand UO_1886 (O_1886,N_14990,N_14881);
nor UO_1887 (O_1887,N_14981,N_14786);
or UO_1888 (O_1888,N_14929,N_14805);
nand UO_1889 (O_1889,N_14796,N_14972);
or UO_1890 (O_1890,N_14816,N_14885);
or UO_1891 (O_1891,N_14911,N_14868);
xnor UO_1892 (O_1892,N_14825,N_14934);
and UO_1893 (O_1893,N_14875,N_14771);
nor UO_1894 (O_1894,N_14789,N_14761);
and UO_1895 (O_1895,N_14920,N_14911);
nor UO_1896 (O_1896,N_14867,N_14847);
xor UO_1897 (O_1897,N_14919,N_14829);
and UO_1898 (O_1898,N_14819,N_14773);
xor UO_1899 (O_1899,N_14970,N_14833);
nand UO_1900 (O_1900,N_14965,N_14975);
xor UO_1901 (O_1901,N_14999,N_14752);
or UO_1902 (O_1902,N_14886,N_14799);
nand UO_1903 (O_1903,N_14933,N_14991);
xnor UO_1904 (O_1904,N_14933,N_14932);
xor UO_1905 (O_1905,N_14916,N_14907);
xor UO_1906 (O_1906,N_14767,N_14773);
or UO_1907 (O_1907,N_14778,N_14940);
nor UO_1908 (O_1908,N_14965,N_14875);
nand UO_1909 (O_1909,N_14948,N_14865);
xor UO_1910 (O_1910,N_14921,N_14755);
xnor UO_1911 (O_1911,N_14931,N_14967);
and UO_1912 (O_1912,N_14854,N_14995);
nor UO_1913 (O_1913,N_14794,N_14870);
xor UO_1914 (O_1914,N_14941,N_14962);
and UO_1915 (O_1915,N_14994,N_14810);
nor UO_1916 (O_1916,N_14824,N_14937);
or UO_1917 (O_1917,N_14932,N_14981);
xor UO_1918 (O_1918,N_14806,N_14940);
nor UO_1919 (O_1919,N_14919,N_14790);
nor UO_1920 (O_1920,N_14946,N_14834);
and UO_1921 (O_1921,N_14753,N_14766);
xnor UO_1922 (O_1922,N_14844,N_14891);
and UO_1923 (O_1923,N_14799,N_14909);
and UO_1924 (O_1924,N_14929,N_14789);
or UO_1925 (O_1925,N_14958,N_14948);
and UO_1926 (O_1926,N_14828,N_14774);
xor UO_1927 (O_1927,N_14911,N_14774);
or UO_1928 (O_1928,N_14768,N_14865);
and UO_1929 (O_1929,N_14892,N_14899);
and UO_1930 (O_1930,N_14870,N_14752);
nor UO_1931 (O_1931,N_14847,N_14973);
and UO_1932 (O_1932,N_14909,N_14753);
xor UO_1933 (O_1933,N_14771,N_14801);
and UO_1934 (O_1934,N_14991,N_14771);
nand UO_1935 (O_1935,N_14867,N_14849);
or UO_1936 (O_1936,N_14849,N_14929);
or UO_1937 (O_1937,N_14776,N_14781);
nand UO_1938 (O_1938,N_14843,N_14938);
xnor UO_1939 (O_1939,N_14968,N_14860);
nor UO_1940 (O_1940,N_14851,N_14834);
nor UO_1941 (O_1941,N_14869,N_14896);
nand UO_1942 (O_1942,N_14864,N_14831);
or UO_1943 (O_1943,N_14856,N_14978);
nor UO_1944 (O_1944,N_14918,N_14916);
nor UO_1945 (O_1945,N_14855,N_14913);
nor UO_1946 (O_1946,N_14790,N_14920);
xor UO_1947 (O_1947,N_14838,N_14782);
and UO_1948 (O_1948,N_14980,N_14836);
nor UO_1949 (O_1949,N_14832,N_14766);
nand UO_1950 (O_1950,N_14806,N_14875);
nor UO_1951 (O_1951,N_14753,N_14929);
and UO_1952 (O_1952,N_14778,N_14971);
or UO_1953 (O_1953,N_14975,N_14852);
nand UO_1954 (O_1954,N_14865,N_14880);
xor UO_1955 (O_1955,N_14880,N_14856);
xor UO_1956 (O_1956,N_14899,N_14813);
nor UO_1957 (O_1957,N_14930,N_14911);
or UO_1958 (O_1958,N_14822,N_14879);
nor UO_1959 (O_1959,N_14983,N_14905);
or UO_1960 (O_1960,N_14839,N_14879);
or UO_1961 (O_1961,N_14894,N_14775);
xnor UO_1962 (O_1962,N_14936,N_14775);
nor UO_1963 (O_1963,N_14751,N_14766);
nor UO_1964 (O_1964,N_14948,N_14911);
xnor UO_1965 (O_1965,N_14845,N_14831);
nor UO_1966 (O_1966,N_14877,N_14861);
nand UO_1967 (O_1967,N_14967,N_14899);
and UO_1968 (O_1968,N_14842,N_14804);
and UO_1969 (O_1969,N_14958,N_14759);
nor UO_1970 (O_1970,N_14915,N_14817);
nor UO_1971 (O_1971,N_14874,N_14781);
xnor UO_1972 (O_1972,N_14932,N_14909);
nand UO_1973 (O_1973,N_14989,N_14864);
nor UO_1974 (O_1974,N_14776,N_14789);
xnor UO_1975 (O_1975,N_14904,N_14947);
nand UO_1976 (O_1976,N_14907,N_14810);
nand UO_1977 (O_1977,N_14942,N_14946);
and UO_1978 (O_1978,N_14960,N_14983);
and UO_1979 (O_1979,N_14979,N_14841);
nor UO_1980 (O_1980,N_14867,N_14791);
nand UO_1981 (O_1981,N_14984,N_14835);
nand UO_1982 (O_1982,N_14805,N_14975);
nor UO_1983 (O_1983,N_14820,N_14803);
nor UO_1984 (O_1984,N_14970,N_14941);
or UO_1985 (O_1985,N_14793,N_14812);
nand UO_1986 (O_1986,N_14780,N_14841);
xnor UO_1987 (O_1987,N_14984,N_14899);
and UO_1988 (O_1988,N_14769,N_14907);
xor UO_1989 (O_1989,N_14952,N_14921);
or UO_1990 (O_1990,N_14876,N_14995);
or UO_1991 (O_1991,N_14955,N_14855);
and UO_1992 (O_1992,N_14972,N_14950);
and UO_1993 (O_1993,N_14769,N_14923);
and UO_1994 (O_1994,N_14932,N_14837);
nor UO_1995 (O_1995,N_14935,N_14929);
nor UO_1996 (O_1996,N_14981,N_14956);
nor UO_1997 (O_1997,N_14791,N_14844);
nor UO_1998 (O_1998,N_14949,N_14822);
and UO_1999 (O_1999,N_14819,N_14820);
endmodule